

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9726, n9727, n9728,
         n9729, n9730, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131;

  BUF_X1 U11160 ( .A(n12819), .Z(n14377) );
  NAND2_X1 U11161 ( .A1(n11037), .A2(n19015), .ZN(n11038) );
  INV_X2 U11162 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11980) );
  CLKBUF_X1 U11163 ( .A(n10748), .Z(n10756) );
  AND2_X1 U11164 ( .A1(n10987), .A2(n9778), .ZN(n11047) );
  AOI211_X2 U11165 ( .C1(n17159), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n10266), .B(n10265), .ZN(n17366) );
  AND2_X2 U11167 ( .A1(n14125), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10970) );
  INV_X1 U11168 ( .A(n17031), .ZN(n17188) );
  INV_X1 U11169 ( .A(n10334), .ZN(n10464) );
  AND2_X1 U11170 ( .A1(n14115), .A2(n10804), .ZN(n14153) );
  CLKBUF_X2 U11171 ( .A(n11898), .Z(n12514) );
  INV_X1 U11172 ( .A(n10221), .ZN(n17156) );
  INV_X1 U11173 ( .A(n14099), .ZN(n14135) );
  CLKBUF_X1 U11175 ( .A(n12010), .Z(n11899) );
  CLKBUF_X2 U11176 ( .A(n11876), .Z(n12515) );
  CLKBUF_X2 U11177 ( .A(n11917), .Z(n13351) );
  OR2_X2 U11178 ( .A1(n20165), .A2(n20144), .ZN(n13141) );
  CLKBUF_X1 U11179 ( .A(n10609), .Z(n19230) );
  INV_X1 U11180 ( .A(n20144), .ZN(n12593) );
  AOI21_X1 U11181 ( .B1(n12520), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n11831), .ZN(n11832) );
  INV_X2 U11182 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15527) );
  AND2_X2 U11183 ( .A1(n18878), .A2(n19884), .ZN(n19029) );
  CLKBUF_X1 U11184 ( .A(n18582), .Z(n9716) );
  NOR2_X1 U11185 ( .A1(n18205), .A2(n18521), .ZN(n18582) );
  AND2_X1 U11186 ( .A1(n14115), .A2(n10788), .ZN(n14137) );
  AND2_X1 U11187 ( .A1(n10691), .A2(n10227), .ZN(n9742) );
  INV_X2 U11190 ( .A(n10742), .ZN(n11361) );
  AND2_X1 U11191 ( .A1(n14115), .A2(n10789), .ZN(n14138) );
  INV_X1 U11192 ( .A(n14165), .ZN(n10796) );
  AND2_X1 U11193 ( .A1(n11890), .A2(n11888), .ZN(n11875) );
  AND2_X1 U11194 ( .A1(n10911), .A2(n10907), .ZN(n10903) );
  AND2_X1 U11195 ( .A1(n11135), .A2(n11134), .ZN(n16107) );
  INV_X1 U11196 ( .A(n9800), .ZN(n16998) );
  INV_X1 U11197 ( .A(n9794), .ZN(n17104) );
  INV_X1 U11198 ( .A(n17121), .ZN(n17155) );
  AND3_X1 U11199 ( .A1(n12114), .A2(n12115), .A3(n9854), .ZN(n13643) );
  AND2_X1 U11200 ( .A1(n14652), .A2(n9898), .ZN(n14630) );
  AOI21_X1 U11201 ( .B1(n15130), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n9817), .ZN(n9911) );
  INV_X1 U11202 ( .A(n17581), .ZN(n17999) );
  INV_X1 U11203 ( .A(n12619), .ZN(n12609) );
  INV_X1 U11204 ( .A(n19052), .ZN(n19032) );
  XNOR2_X1 U11205 ( .A(n9912), .B(n14046), .ZN(n15130) );
  INV_X1 U11206 ( .A(n16525), .ZN(n16841) );
  INV_X2 U11207 ( .A(n17121), .ZN(n9722) );
  INV_X1 U11208 ( .A(n17861), .ZN(n17847) );
  NAND2_X1 U11209 ( .A1(n18068), .A2(n18670), .ZN(n18088) );
  INV_X1 U11210 ( .A(n19982), .ZN(n19992) );
  OR2_X1 U11211 ( .A1(n15048), .A2(n15047), .ZN(n15274) );
  INV_X1 U11212 ( .A(n9795), .ZN(n10268) );
  INV_X2 U11213 ( .A(n17679), .ZN(n17765) );
  OAI21_X1 U11215 ( .B1(n13371), .B2(n12740), .A(n12725), .ZN(n13395) );
  INV_X1 U11216 ( .A(n14165), .ZN(n9717) );
  AND2_X4 U11217 ( .A1(n11191), .A2(n10802), .ZN(n10795) );
  OAI22_X2 U11218 ( .A1(n13058), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n12741), 
        .B2(n12009), .ZN(n11974) );
  AND2_X1 U11219 ( .A1(n10787), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9718) );
  INV_X2 U11221 ( .A(n11419), .ZN(n10699) );
  OR2_X2 U11222 ( .A1(n16867), .A2(n10247), .ZN(n9800) );
  AND2_X1 U11223 ( .A1(n13344), .A2(n11720), .ZN(n9720) );
  AND2_X2 U11224 ( .A1(n13344), .A2(n11720), .ZN(n9721) );
  AND2_X1 U11225 ( .A1(n13344), .A2(n11720), .ZN(n9757) );
  AND2_X1 U11226 ( .A1(n13344), .A2(n11720), .ZN(n11960) );
  AND3_X4 U11227 ( .A1(n9981), .A2(n9884), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10639) );
  NOR2_X2 U11228 ( .A1(n18185), .A2(n17951), .ZN(n17992) );
  NAND2_X4 U11229 ( .A1(n10188), .A2(n10187), .ZN(n10688) );
  OR2_X2 U11230 ( .A1(n15224), .A2(n15225), .ZN(n9874) );
  AND2_X4 U11231 ( .A1(n11729), .A2(n11731), .ZN(n11900) );
  NOR2_X2 U11235 ( .A1(n15191), .A2(n15190), .ZN(n15192) );
  NOR2_X2 U11236 ( .A1(n17754), .A2(n17974), .ZN(n17637) );
  XNOR2_X2 U11237 ( .A(n11038), .B(n15483), .ZN(n15255) );
  AND2_X1 U11239 ( .A1(n15327), .A2(n9933), .ZN(n15126) );
  AND2_X1 U11240 ( .A1(n9883), .A2(n15419), .ZN(n16133) );
  OAI21_X1 U11241 ( .B1(n15415), .B2(n15433), .A(n14024), .ZN(n9883) );
  AOI21_X1 U11243 ( .B1(n10006), .B2(n10112), .A(n9901), .ZN(n9893) );
  INV_X1 U11244 ( .A(n13504), .ZN(n12115) );
  NOR2_X2 U11245 ( .A1(n15084), .A2(n15074), .ZN(n15076) );
  OAI21_X1 U11246 ( .B1(n13600), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13601), .ZN(n9880) );
  NAND2_X1 U11247 ( .A1(n9738), .A2(n14734), .ZN(n14735) );
  CLKBUF_X1 U11248 ( .A(n13371), .Z(n13372) );
  OAI211_X1 U11249 ( .C1(n13371), .C2(n12220), .A(n11983), .B(n11982), .ZN(
        n11984) );
  AND2_X1 U11250 ( .A1(n14541), .A2(n9788), .ZN(n14508) );
  NOR2_X1 U11251 ( .A1(n15451), .A2(n15450), .ZN(n13465) );
  AND2_X1 U11252 ( .A1(n10761), .A2(n10780), .ZN(n13539) );
  NOR2_X1 U11253 ( .A1(n10772), .A2(n10776), .ZN(n19374) );
  CLKBUF_X2 U11254 ( .A(n10762), .Z(n15517) );
  CLKBUF_X1 U11255 ( .A(n14059), .Z(n20521) );
  AND2_X1 U11256 ( .A1(n10753), .A2(n10752), .ZN(n19170) );
  OR2_X1 U11257 ( .A1(n12588), .A2(n12587), .ZN(n14351) );
  XNOR2_X1 U11258 ( .A(n11890), .B(n11889), .ZN(n11995) );
  NAND2_X1 U11259 ( .A1(n17808), .A2(n17809), .ZN(n17807) );
  NAND4_X1 U11260 ( .A1(n9820), .A2(n9887), .A3(n9886), .A4(n9890), .ZN(n9889)
         );
  INV_X1 U11261 ( .A(n18210), .ZN(n18855) );
  INV_X1 U11262 ( .A(n18227), .ZN(n17238) );
  AOI211_X2 U11263 ( .C1(n17159), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n10404), .B(n10403), .ZN(n18210) );
  OAI211_X1 U11264 ( .C1(n10298), .C2(n20961), .A(n10414), .B(n10413), .ZN(
        n10537) );
  INV_X2 U11265 ( .A(n12907), .ZN(n10702) );
  OR3_X1 U11266 ( .A1(n10296), .A2(n10295), .A3(n10294), .ZN(n10508) );
  NAND2_X1 U11267 ( .A1(n14257), .A2(n9730), .ZN(n11381) );
  CLKBUF_X1 U11268 ( .A(n12863), .Z(n9740) );
  NAND2_X1 U11269 ( .A1(n10657), .A2(n11034), .ZN(n10680) );
  NAND2_X2 U11270 ( .A1(n19883), .A2(n10688), .ZN(n12907) );
  INV_X2 U11271 ( .A(n20155), .ZN(n12606) );
  INV_X1 U11272 ( .A(n11034), .ZN(n14042) );
  BUF_X1 U11273 ( .A(n10672), .Z(n10711) );
  INV_X1 U11274 ( .A(n19224), .ZN(n9726) );
  MUX2_X1 U11275 ( .A(n10655), .B(n10654), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10672) );
  INV_X4 U11276 ( .A(n10275), .ZN(n9727) );
  INV_X2 U11277 ( .A(n10298), .ZN(n17182) );
  CLKBUF_X2 U11278 ( .A(n12015), .Z(n11903) );
  CLKBUF_X3 U11279 ( .A(n10287), .Z(n9733) );
  CLKBUF_X2 U11280 ( .A(n11958), .Z(n12522) );
  CLKBUF_X2 U11282 ( .A(n10301), .Z(n17143) );
  CLKBUF_X2 U11283 ( .A(n10965), .Z(n14143) );
  BUF_X2 U11285 ( .A(n10801), .Z(n14315) );
  BUF_X2 U11286 ( .A(n10639), .Z(n10038) );
  INV_X2 U11287 ( .A(n14309), .ZN(n14125) );
  NAND2_X1 U11288 ( .A1(n21016), .A2(n18834), .ZN(n16867) );
  XNOR2_X1 U11289 ( .A(n14377), .B(n12818), .ZN(n14629) );
  AND2_X1 U11290 ( .A1(n14403), .A2(n14499), .ZN(n15656) );
  NAND2_X1 U11291 ( .A1(n10049), .A2(n10050), .ZN(n15119) );
  NOR2_X1 U11292 ( .A1(n9899), .A2(n9872), .ZN(n9898) );
  NAND2_X1 U11293 ( .A1(n15217), .A2(n15214), .ZN(n15204) );
  AND2_X1 U11294 ( .A1(n9749), .A2(n9750), .ZN(n15191) );
  NAND2_X1 U11295 ( .A1(n9874), .A2(n15176), .ZN(n15217) );
  OAI21_X1 U11296 ( .B1(n11717), .B2(n19196), .A(n9816), .ZN(n9931) );
  OR2_X1 U11297 ( .A1(n10104), .A2(n10103), .ZN(n12807) );
  NAND2_X1 U11298 ( .A1(n9960), .A2(n14685), .ZN(n14642) );
  NAND2_X1 U11299 ( .A1(n14970), .A2(n10136), .ZN(n10141) );
  AOI21_X1 U11300 ( .B1(n10138), .B2(n14970), .A(n10137), .ZN(n10139) );
  NAND2_X1 U11301 ( .A1(n15464), .A2(n11701), .ZN(n16109) );
  NAND2_X1 U11303 ( .A1(n14744), .A2(n12794), .ZN(n14705) );
  NOR2_X1 U11304 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15547), .ZN(
        n10389) );
  AND2_X1 U11305 ( .A1(n14040), .A2(n10048), .ZN(n10050) );
  INV_X1 U11306 ( .A(n16390), .ZN(n17521) );
  OAI21_X1 U11307 ( .B1(n17532), .B2(n9958), .A(n9957), .ZN(n17522) );
  AOI21_X1 U11308 ( .B1(n10145), .B2(n10146), .A(n15470), .ZN(n10143) );
  AND2_X1 U11309 ( .A1(n11039), .A2(n9848), .ZN(n9984) );
  AND2_X1 U11310 ( .A1(n15057), .A2(n15056), .ZN(n16020) );
  NAND2_X1 U11311 ( .A1(n10158), .A2(n9856), .ZN(n10157) );
  OR2_X1 U11312 ( .A1(n10383), .A2(n10382), .ZN(n10384) );
  AOI21_X1 U11313 ( .B1(n10147), .B2(n15243), .A(n9818), .ZN(n10145) );
  OR2_X1 U11314 ( .A1(n10992), .A2(n13781), .ZN(n10226) );
  NOR2_X1 U11315 ( .A1(n14999), .A2(n14998), .ZN(n14997) );
  NAND2_X1 U11316 ( .A1(n9915), .A2(n9810), .ZN(n9918) );
  NAND2_X1 U11317 ( .A1(n15076), .A2(n15065), .ZN(n15067) );
  AOI211_X1 U11318 ( .C1(n14374), .C2(n14373), .A(n14372), .B(n14371), .ZN(
        n14375) );
  NAND2_X1 U11319 ( .A1(n10913), .A2(n9880), .ZN(n19157) );
  OR2_X1 U11320 ( .A1(n17765), .A2(n17559), .ZN(n17549) );
  NAND2_X1 U11321 ( .A1(n11153), .A2(n11152), .ZN(n14044) );
  OR2_X1 U11322 ( .A1(n12800), .A2(n10114), .ZN(n10113) );
  AND2_X1 U11323 ( .A1(n10093), .A2(n12775), .ZN(n10092) );
  AND2_X1 U11324 ( .A1(n11662), .A2(n11661), .ZN(n11691) );
  INV_X1 U11325 ( .A(n10074), .ZN(n17559) );
  AND2_X1 U11326 ( .A1(n12793), .A2(n10230), .ZN(n10119) );
  OR2_X1 U11327 ( .A1(n11684), .A2(n13781), .ZN(n13775) );
  INV_X1 U11328 ( .A(n14701), .ZN(n9901) );
  NAND2_X1 U11329 ( .A1(n10983), .A2(n9799), .ZN(n11661) );
  NAND2_X1 U11330 ( .A1(n10983), .A2(n10982), .ZN(n11663) );
  AND2_X1 U11331 ( .A1(n13403), .A2(n13404), .ZN(n13438) );
  NOR2_X2 U11332 ( .A1(n13528), .A2(n13519), .ZN(n13558) );
  INV_X1 U11333 ( .A(n10981), .ZN(n10983) );
  NAND2_X1 U11334 ( .A1(n10235), .A2(n13486), .ZN(n13528) );
  NAND2_X1 U11335 ( .A1(n16246), .A2(n10181), .ZN(n15391) );
  AND2_X1 U11336 ( .A1(n10153), .A2(n9852), .ZN(n10235) );
  NAND2_X1 U11337 ( .A1(n10011), .A2(n10012), .ZN(n12789) );
  NAND2_X1 U11338 ( .A1(n10534), .A2(n17755), .ZN(n18056) );
  AND2_X1 U11339 ( .A1(n10979), .A2(n10978), .ZN(n10982) );
  INV_X1 U11340 ( .A(n9744), .ZN(n10380) );
  AND2_X1 U11341 ( .A1(n10370), .A2(n17679), .ZN(n17650) );
  NAND2_X1 U11342 ( .A1(n9744), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9949) );
  NOR2_X2 U11343 ( .A1(n17857), .A2(n17850), .ZN(n17708) );
  INV_X1 U11344 ( .A(n15202), .ZN(n9728) );
  NAND2_X1 U11345 ( .A1(n11032), .A2(n11031), .ZN(n11686) );
  NAND2_X1 U11346 ( .A1(n12051), .A2(n9843), .ZN(n12106) );
  NAND2_X1 U11347 ( .A1(n13309), .A2(n13308), .ZN(n13380) );
  NAND2_X1 U11348 ( .A1(n13307), .A2(n13306), .ZN(n13308) );
  NAND2_X1 U11349 ( .A1(n12025), .A2(n11977), .ZN(n13371) );
  NAND2_X1 U11350 ( .A1(n10007), .A2(n10008), .ZN(n12025) );
  AND2_X1 U11351 ( .A1(n13305), .A2(n13385), .ZN(n13309) );
  INV_X1 U11352 ( .A(n19374), .ZN(n10946) );
  NAND2_X1 U11353 ( .A1(n11987), .A2(n11986), .ZN(n20223) );
  OR2_X1 U11354 ( .A1(n13381), .A2(n13304), .ZN(n13305) );
  INV_X1 U11355 ( .A(n9765), .ZN(n9766) );
  NAND2_X1 U11356 ( .A1(n10781), .A2(n10777), .ZN(n10994) );
  NAND2_X1 U11357 ( .A1(n13303), .A2(n13302), .ZN(n13381) );
  AND2_X1 U11358 ( .A1(n10781), .A2(n10780), .ZN(n19559) );
  AND2_X1 U11359 ( .A1(n9903), .A2(n10781), .ZN(n19472) );
  CLKBUF_X1 U11360 ( .A(n12864), .Z(n14619) );
  NAND2_X1 U11361 ( .A1(n13218), .A2(n13217), .ZN(n13306) );
  OR2_X1 U11362 ( .A1(n13218), .A2(n13217), .ZN(n13219) );
  NAND2_X1 U11363 ( .A1(n13076), .A2(n13075), .ZN(n13223) );
  NAND2_X1 U11364 ( .A1(n13216), .A2(n13215), .ZN(n13218) );
  NAND2_X1 U11365 ( .A1(n10528), .A2(n17782), .ZN(n17776) );
  NAND2_X1 U11366 ( .A1(n11940), .A2(n11939), .ZN(n11942) );
  NAND2_X1 U11367 ( .A1(n9896), .A2(n12023), .ZN(n13373) );
  NOR2_X1 U11368 ( .A1(n15937), .A2(n13727), .ZN(n15758) );
  NAND2_X1 U11369 ( .A1(n13778), .A2(n11444), .ZN(n13109) );
  XNOR2_X1 U11370 ( .A(n13220), .B(n13221), .ZN(n13076) );
  NAND2_X1 U11371 ( .A1(n13104), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13103) );
  NAND2_X1 U11372 ( .A1(n13015), .A2(n13014), .ZN(n13220) );
  NOR2_X1 U11373 ( .A1(n18240), .A2(n17383), .ZN(n17353) );
  NAND2_X1 U11374 ( .A1(n10003), .A2(n11932), .ZN(n11938) );
  CLKBUF_X1 U11375 ( .A(n12729), .Z(n20222) );
  NOR2_X1 U11376 ( .A1(n13478), .A2(n11439), .ZN(n13566) );
  OR2_X1 U11377 ( .A1(n13078), .A2(n19170), .ZN(n10760) );
  NAND2_X1 U11379 ( .A1(n10734), .A2(n10733), .ZN(n10735) );
  CLKBUF_X1 U11380 ( .A(n11995), .Z(n20256) );
  AND2_X1 U11381 ( .A1(n9956), .A2(n17785), .ZN(n9954) );
  NOR2_X1 U11382 ( .A1(n13429), .A2(n11429), .ZN(n13476) );
  XNOR2_X1 U11383 ( .A(n11264), .B(n11263), .ZN(n11261) );
  OAI21_X1 U11384 ( .B1(n17807), .B2(n9951), .A(n9950), .ZN(n9955) );
  XNOR2_X1 U11385 ( .A(n11857), .B(n11943), .ZN(n20257) );
  NAND2_X1 U11386 ( .A1(n11145), .A2(n11048), .ZN(n11050) );
  OR2_X1 U11387 ( .A1(n11429), .A2(n11427), .ZN(n13428) );
  AND2_X1 U11388 ( .A1(n10014), .A2(n10013), .ZN(n13443) );
  OAI21_X1 U11389 ( .B1(n16297), .B2(n10741), .A(n10745), .ZN(n11263) );
  AOI21_X1 U11390 ( .B1(n13082), .B2(n11426), .A(n11425), .ZN(n11429) );
  INV_X1 U11391 ( .A(n11888), .ZN(n11889) );
  NAND2_X1 U11392 ( .A1(n17824), .A2(n10358), .ZN(n17808) );
  NAND2_X1 U11393 ( .A1(n9889), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U11394 ( .A1(n17825), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17824) );
  OR2_X1 U11395 ( .A1(n11872), .A2(n13145), .ZN(n11888) );
  INV_X1 U11396 ( .A(n10364), .ZN(n16394) );
  NAND2_X1 U11397 ( .A1(n10904), .A2(n10903), .ZN(n10985) );
  INV_X2 U11398 ( .A(n17500), .ZN(n9729) );
  AND2_X1 U11399 ( .A1(n10709), .A2(n10708), .ZN(n10710) );
  AND2_X1 U11400 ( .A1(n9797), .A2(n11840), .ZN(n9887) );
  AND2_X1 U11401 ( .A1(n13041), .A2(n13042), .ZN(n13040) );
  AOI21_X1 U11402 ( .B1(n10100), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n9775), 
        .ZN(n10098) );
  NAND2_X1 U11403 ( .A1(n10044), .A2(n10043), .ZN(n10911) );
  CLKBUF_X1 U11404 ( .A(n11197), .Z(n13033) );
  NAND2_X1 U11405 ( .A1(n17837), .A2(n17836), .ZN(n17835) );
  NAND2_X1 U11406 ( .A1(n10703), .A2(n11643), .ZN(n13319) );
  INV_X1 U11407 ( .A(n18204), .ZN(n17392) );
  NOR2_X1 U11408 ( .A1(n11993), .A2(n11924), .ZN(n10100) );
  NAND2_X1 U11409 ( .A1(n12613), .A2(n12612), .ZN(n10019) );
  NAND2_X1 U11410 ( .A1(n10682), .A2(n10681), .ZN(n11206) );
  NOR3_X1 U11411 ( .A1(n10537), .A2(n17231), .A3(n13906), .ZN(n10544) );
  AND2_X1 U11412 ( .A1(n11376), .A2(n10696), .ZN(n10703) );
  AND2_X1 U11413 ( .A1(n11846), .A2(n12606), .ZN(n13353) );
  AND2_X1 U11414 ( .A1(n11851), .A2(n11850), .ZN(n12816) );
  AND2_X1 U11415 ( .A1(n10282), .A2(n10281), .ZN(n17373) );
  AND2_X1 U11416 ( .A1(n12603), .A2(n20144), .ZN(n11846) );
  AOI211_X2 U11417 ( .C1(n9727), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n10452), .B(n10451), .ZN(n18227) );
  AND2_X1 U11418 ( .A1(n10702), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11228) );
  INV_X1 U11419 ( .A(n11848), .ZN(n12595) );
  OAI211_X1 U11420 ( .C1(n17170), .C2(n10425), .A(n10424), .B(n10423), .ZN(
        n17231) );
  AOI211_X1 U11421 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n10412), .B(n10411), .ZN(n10413) );
  BUF_X4 U11423 ( .A(n14042), .Z(n9755) );
  OR2_X2 U11424 ( .A1(n12606), .A2(n20144), .ZN(n12610) );
  NAND3_X1 U11425 ( .A1(n9944), .A2(n9945), .A3(n9812), .ZN(n10348) );
  OR2_X1 U11426 ( .A1(n11029), .A2(n11028), .ZN(n11443) );
  NOR2_X1 U11427 ( .A1(n10672), .A2(n9726), .ZN(n10676) );
  OR2_X1 U11428 ( .A1(n10810), .A2(n10809), .ZN(n11430) );
  OR2_X1 U11429 ( .A1(n10930), .A2(n10929), .ZN(n11435) );
  INV_X1 U11430 ( .A(n12551), .ZN(n12817) );
  NAND2_X1 U11431 ( .A1(n11034), .A2(n19230), .ZN(n11419) );
  AND3_X1 U11432 ( .A1(n10310), .A2(n10305), .A3(n10308), .ZN(n9944) );
  NAND2_X1 U11433 ( .A1(n12009), .A2(n12008), .ZN(n12585) );
  NAND2_X1 U11434 ( .A1(n20188), .A2(n20181), .ZN(n12863) );
  CLKBUF_X1 U11435 ( .A(n11841), .Z(n20160) );
  NAND2_X2 U11436 ( .A1(n10630), .A2(n10629), .ZN(n19224) );
  NAND2_X2 U11437 ( .A1(n10185), .A2(n10184), .ZN(n11034) );
  NAND2_X2 U11438 ( .A1(n9802), .A2(n10237), .ZN(n20181) );
  NAND2_X1 U11440 ( .A1(n10580), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10184) );
  NAND2_X1 U11441 ( .A1(n10597), .A2(n10596), .ZN(n10609) );
  AND3_X1 U11443 ( .A1(n11833), .A2(n11821), .A3(n11834), .ZN(n10015) );
  NAND2_X1 U11444 ( .A1(n10585), .A2(n10614), .ZN(n10185) );
  INV_X2 U11445 ( .A(n19883), .ZN(n9730) );
  OR2_X2 U11446 ( .A1(n11793), .A2(n11792), .ZN(n20188) );
  NAND2_X2 U11447 ( .A1(n18869), .A2(n21050), .ZN(n18791) );
  AND4_X1 U11448 ( .A1(n11797), .A2(n11796), .A3(n11795), .A4(n11794), .ZN(
        n11813) );
  AND4_X1 U11449 ( .A1(n11805), .A2(n11804), .A3(n11803), .A4(n11802), .ZN(
        n11811) );
  AND4_X1 U11450 ( .A1(n11809), .A2(n11808), .A3(n11807), .A4(n11806), .ZN(
        n11810) );
  AND4_X1 U11451 ( .A1(n11801), .A2(n11800), .A3(n11799), .A4(n11798), .ZN(
        n11812) );
  NAND2_X2 U11452 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19805), .ZN(n19813) );
  AND4_X1 U11453 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n11815), .ZN(
        n11834) );
  AND2_X2 U11454 ( .A1(n14302), .A2(n13326), .ZN(n14150) );
  AND4_X1 U11455 ( .A1(n11827), .A2(n11826), .A3(n11825), .A4(n11824), .ZN(
        n11833) );
  AND4_X1 U11456 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11762) );
  INV_X2 U11457 ( .A(n16481), .ZN(U215) );
  AND4_X1 U11458 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n10238) );
  AND4_X1 U11459 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(
        n11763) );
  NAND2_X2 U11461 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18869), .ZN(n18794) );
  NAND2_X2 U11462 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10241), .ZN(
        n10298) );
  INV_X2 U11463 ( .A(n18179), .ZN(n9732) );
  BUF_X2 U11464 ( .A(n11916), .Z(n11893) );
  INV_X2 U11465 ( .A(n20107), .ZN(n13397) );
  CLKBUF_X1 U11466 ( .A(n13811), .Z(n13550) );
  INV_X4 U11467 ( .A(n10234), .ZN(n17162) );
  AND3_X1 U11468 ( .A1(n10638), .A2(n10637), .A3(n10614), .ZN(n10643) );
  AND3_X1 U11469 ( .A1(n10632), .A2(n10631), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10636) );
  INV_X2 U11470 ( .A(n10287), .ZN(n17170) );
  CLKBUF_X1 U11471 ( .A(n9798), .Z(n17118) );
  INV_X2 U11472 ( .A(n16483), .ZN(n16485) );
  BUF_X2 U11473 ( .A(n11901), .Z(n11911) );
  OR2_X2 U11474 ( .A1(n10245), .A2(n16867), .ZN(n10221) );
  OAI221_X1 U11475 ( .B1(n20990), .B2(keyinput122), .C1(n13461), .C2(
        keyinput103), .A(n20989), .ZN(n20991) );
  NOR3_X2 U11476 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n16867), .ZN(n10334) );
  BUF_X2 U11477 ( .A(n12016), .Z(n12521) );
  OR2_X2 U11478 ( .A1(n18685), .A2(n10247), .ZN(n10234) );
  OR2_X1 U11479 ( .A1(n10246), .A2(n10245), .ZN(n17121) );
  INV_X1 U11480 ( .A(n14309), .ZN(n9763) );
  AND2_X2 U11481 ( .A1(n11730), .A2(n13345), .ZN(n11958) );
  AND2_X2 U11482 ( .A1(n11732), .A2(n13361), .ZN(n11898) );
  INV_X2 U11483 ( .A(n19891), .ZN(n19805) );
  NAND2_X1 U11484 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18826), .ZN(
        n10245) );
  NAND2_X1 U11485 ( .A1(n21016), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10246) );
  INV_X2 U11486 ( .A(n20800), .ZN(n9734) );
  NAND2_X1 U11487 ( .A1(n18819), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10247) );
  AND2_X2 U11488 ( .A1(n11952), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11732) );
  NAND3_X2 U11489 ( .A1(n15505), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14309) );
  AND2_X1 U11490 ( .A1(n11191), .A2(n10802), .ZN(n9761) );
  NOR2_X1 U11491 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11853), .ZN(
        n11730) );
  BUF_X2 U11492 ( .A(n11723), .Z(n13345) );
  NOR2_X2 U11493 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10789) );
  INV_X1 U11494 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18819) );
  INV_X2 U11495 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21016) );
  NAND2_X2 U11496 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18685) );
  INV_X1 U11497 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15505) );
  INV_X4 U11499 ( .A(n11619), .ZN(n11635) );
  NAND2_X1 U11501 ( .A1(n11206), .A2(n13814), .ZN(n9735) );
  NAND2_X1 U11502 ( .A1(n12806), .A2(n9738), .ZN(n9736) );
  AND2_X2 U11503 ( .A1(n9736), .A2(n9737), .ZN(n14669) );
  OR2_X1 U11504 ( .A1(n15794), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9737) );
  INV_X1 U11507 ( .A(n13324), .ZN(n9741) );
  OR2_X2 U11508 ( .A1(n11646), .A2(n9742), .ZN(n10695) );
  AND2_X1 U11509 ( .A1(n9743), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10241) );
  AND2_X1 U11510 ( .A1(n18834), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9743) );
  OR2_X2 U11511 ( .A1(n17974), .A2(n17696), .ZN(n9744) );
  NAND2_X1 U11512 ( .A1(n14631), .A2(n10111), .ZN(n12811) );
  OAI21_X1 U11513 ( .B1(n9735), .B2(n19218), .A(n10683), .ZN(n9745) );
  OAI21_X1 U11514 ( .B1(n11371), .B2(n19218), .A(n10683), .ZN(n10720) );
  AND2_X2 U11517 ( .A1(n14412), .A2(n12407), .ZN(n14413) );
  BUF_X8 U11518 ( .A(n11900), .Z(n12520) );
  XNOR2_X1 U11519 ( .A(n10736), .B(n10735), .ZN(n10746) );
  NOR2_X2 U11520 ( .A1(n14551), .A2(n14550), .ZN(n14552) );
  NAND2_X1 U11521 ( .A1(n11243), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10741) );
  INV_X1 U11522 ( .A(n11952), .ZN(n9746) );
  NOR2_X1 U11523 ( .A1(n14692), .A2(n9747), .ZN(n10103) );
  OR2_X1 U11524 ( .A1(n9871), .A2(n14687), .ZN(n9747) );
  XNOR2_X1 U11525 ( .A(n12747), .B(n20101), .ZN(n9748) );
  INV_X4 U11526 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11952) );
  XNOR2_X1 U11527 ( .A(n12747), .B(n20101), .ZN(n13411) );
  NAND2_X1 U11528 ( .A1(n9874), .A2(n15176), .ZN(n9749) );
  AND2_X1 U11529 ( .A1(n9728), .A2(n15214), .ZN(n9750) );
  NAND2_X1 U11530 ( .A1(n10938), .A2(n10937), .ZN(n13772) );
  NAND2_X1 U11531 ( .A1(n12808), .A2(n9900), .ZN(n14652) );
  OAI22_X1 U11532 ( .A1(n14626), .A2(n9738), .B1(n12811), .B2(n14783), .ZN(
        n12812) );
  NAND2_X1 U11533 ( .A1(n13314), .A2(n12737), .ZN(n12738) );
  OAI21_X1 U11534 ( .B1(n15191), .B2(n15178), .A(n15188), .ZN(n15179) );
  XNOR2_X1 U11535 ( .A(n9751), .B(n15179), .ZN(n15363) );
  AND2_X1 U11536 ( .A1(n15170), .A2(n15169), .ZN(n9751) );
  XNOR2_X1 U11537 ( .A(n10756), .B(n10749), .ZN(n13078) );
  NAND2_X1 U11538 ( .A1(n11243), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U11539 ( .A1(n11243), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9753) );
  BUF_X1 U11540 ( .A(n9753), .Z(n11355) );
  AND4_X1 U11541 ( .A1(n10622), .A2(n10621), .A3(n10620), .A4(n10619), .ZN(
        n10623) );
  AOI211_X2 U11542 ( .C1(n17972), .C2(n18058), .A(n17971), .B(n17970), .ZN(
        n17982) );
  NOR2_X2 U11544 ( .A1(n14451), .A2(n14452), .ZN(n14438) );
  OAI211_X2 U11545 ( .C1(n9983), .C2(n15254), .A(n10215), .B(n9913), .ZN(
        n16160) );
  NAND2_X2 U11546 ( .A1(n10993), .A2(n10226), .ZN(n15254) );
  NOR2_X1 U11547 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U11548 ( .A1(n10623), .A2(n10614), .ZN(n10630) );
  AND2_X1 U11549 ( .A1(n13344), .A2(n11720), .ZN(n9756) );
  OR2_X1 U11550 ( .A1(n10720), .A2(n10712), .ZN(n10684) );
  NAND2_X1 U11551 ( .A1(n10707), .A2(n10706), .ZN(n10742) );
  NOR2_X2 U11552 ( .A1(n16391), .A2(n17860), .ZN(n17767) );
  NOR2_X1 U11553 ( .A1(n10768), .A2(n10760), .ZN(n19590) );
  NAND2_X1 U11554 ( .A1(n10685), .A2(n10684), .ZN(n10728) );
  AND2_X1 U11555 ( .A1(n11732), .A2(n13361), .ZN(n9758) );
  INV_X1 U11556 ( .A(n10741), .ZN(n9759) );
  AND2_X1 U11557 ( .A1(n11191), .A2(n10802), .ZN(n9760) );
  NOR2_X4 U11558 ( .A1(n16129), .A2(n16251), .ZN(n10168) );
  OAI21_X2 U11559 ( .B1(n16117), .B2(n14026), .A(n16119), .ZN(n15174) );
  INV_X1 U11560 ( .A(n10663), .ZN(n9762) );
  INV_X4 U11561 ( .A(n14275), .ZN(n10663) );
  NAND2_X1 U11562 ( .A1(n9982), .A2(n9981), .ZN(n14275) );
  INV_X2 U11563 ( .A(n19313), .ZN(n10950) );
  NOR2_X2 U11564 ( .A1(n10779), .A2(n10778), .ZN(n19313) );
  INV_X2 U11565 ( .A(n14309), .ZN(n9764) );
  INV_X1 U11566 ( .A(n18645), .ZN(n9765) );
  AND2_X4 U11567 ( .A1(n11729), .A2(n11728), .ZN(n12015) );
  OAI21_X1 U11568 ( .B1(n10702), .B2(n10701), .A(n10700), .ZN(n11643) );
  NAND2_X1 U11569 ( .A1(n10699), .A2(n10711), .ZN(n10700) );
  NAND2_X1 U11570 ( .A1(n10698), .A2(n19218), .ZN(n10701) );
  INV_X1 U11571 ( .A(n10697), .ZN(n10698) );
  INV_X1 U11572 ( .A(n9939), .ZN(n9938) );
  OAI211_X1 U11573 ( .C1(n10268), .C2(n9942), .A(n9941), .B(n9940), .ZN(n9939)
         );
  INV_X1 U11574 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n9942) );
  NAND2_X1 U11575 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n9941) );
  INV_X1 U11576 ( .A(n12105), .ZN(n10012) );
  INV_X1 U11577 ( .A(n12106), .ZN(n10011) );
  INV_X1 U11578 ( .A(n13071), .ZN(n14207) );
  NAND2_X1 U11579 ( .A1(n10603), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10188) );
  NAND2_X1 U11580 ( .A1(n10608), .A2(n10614), .ZN(n10187) );
  NAND2_X1 U11581 ( .A1(n9759), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10734) );
  NAND2_X1 U11582 ( .A1(n13539), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10759) );
  INV_X1 U11583 ( .A(n13539), .ZN(n11008) );
  AND2_X1 U11584 ( .A1(n12096), .A2(n12095), .ZN(n12105) );
  NAND2_X1 U11585 ( .A1(n11931), .A2(n11930), .ZN(n11993) );
  AND3_X1 U11586 ( .A1(n11929), .A2(n11928), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11930) );
  NAND2_X1 U11587 ( .A1(n20171), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12009) );
  AND2_X2 U11588 ( .A1(n10038), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14136) );
  INV_X1 U11590 ( .A(n14404), .ZN(n10131) );
  AND2_X1 U11591 ( .A1(n14498), .A2(n14510), .ZN(n10132) );
  INV_X1 U11592 ( .A(n12780), .ZN(n12790) );
  AND2_X1 U11593 ( .A1(n14207), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13304) );
  INV_X1 U11594 ( .A(n15021), .ZN(n10202) );
  NAND2_X1 U11595 ( .A1(n9910), .A2(n15149), .ZN(n11151) );
  NAND2_X1 U11596 ( .A1(n15150), .A2(n15152), .ZN(n9910) );
  AND4_X1 U11597 ( .A1(n10879), .A2(n10878), .A3(n10877), .A4(n10876), .ZN(
        n10892) );
  NOR2_X1 U11598 ( .A1(n13071), .A2(n9730), .ZN(n10707) );
  AND2_X1 U11599 ( .A1(n13814), .A2(n19871), .ZN(n11418) );
  AND4_X1 U11600 ( .A1(n13814), .A2(n10689), .A3(n19218), .A4(n9726), .ZN(
        n10696) );
  INV_X1 U11601 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9884) );
  NAND2_X1 U11602 ( .A1(n21016), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10089) );
  NOR2_X1 U11603 ( .A1(n18240), .A2(n18219), .ZN(n10552) );
  NAND2_X1 U11604 ( .A1(n13411), .A2(n13410), .ZN(n13409) );
  NAND2_X1 U11605 ( .A1(n13141), .A2(n12619), .ZN(n14354) );
  NAND2_X1 U11607 ( .A1(n14685), .A2(n10105), .ZN(n10104) );
  AND2_X1 U11608 ( .A1(n10107), .A2(n10106), .ZN(n10105) );
  INV_X1 U11609 ( .A(n13150), .ZN(n13149) );
  NAND2_X1 U11610 ( .A1(n10092), .A2(n10095), .ZN(n10090) );
  NAND2_X1 U11611 ( .A1(n13443), .A2(n9804), .ZN(n15967) );
  OR2_X1 U11612 ( .A1(n20077), .A2(n20092), .ZN(n10117) );
  NOR2_X1 U11613 ( .A1(n11370), .A2(n11369), .ZN(n16316) );
  NOR2_X1 U11614 ( .A1(n13382), .A2(n10155), .ZN(n10154) );
  INV_X1 U11615 ( .A(n13379), .ZN(n10155) );
  AND2_X1 U11616 ( .A1(n13381), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13382) );
  XNOR2_X1 U11617 ( .A(n11712), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12896) );
  NAND2_X1 U11618 ( .A1(n15121), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11712) );
  NAND2_X1 U11619 ( .A1(n14039), .A2(n14040), .ZN(n9912) );
  AND2_X1 U11620 ( .A1(n11241), .A2(n19737), .ZN(n11704) );
  NAND2_X1 U11621 ( .A1(n13219), .A2(n13306), .ZN(n13226) );
  NAND2_X1 U11622 ( .A1(n19282), .A2(n19848), .ZN(n19438) );
  AND2_X1 U11623 ( .A1(n19282), .A2(n19281), .ZN(n19369) );
  NAND2_X1 U11624 ( .A1(n17522), .A2(n9959), .ZN(n15547) );
  NOR2_X1 U11625 ( .A1(n17765), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9959) );
  NOR2_X1 U11626 ( .A1(n17650), .A2(n10223), .ZN(n10374) );
  NAND2_X1 U11627 ( .A1(n9949), .A2(n9948), .ZN(n17645) );
  AND2_X1 U11628 ( .A1(n10374), .A2(n17981), .ZN(n9948) );
  XNOR2_X1 U11629 ( .A(n11367), .B(n11366), .ZN(n11715) );
  OR2_X1 U11630 ( .A1(n14950), .A2(n11360), .ZN(n11367) );
  INV_X1 U11631 ( .A(n12564), .ZN(n12541) );
  OR2_X1 U11632 ( .A1(n12554), .A2(n12555), .ZN(n12556) );
  OAI21_X1 U11633 ( .B1(n19409), .B2(n14084), .A(n9877), .ZN(n10957) );
  NAND2_X1 U11634 ( .A1(n9904), .A2(n9902), .ZN(n10828) );
  NAND2_X1 U11635 ( .A1(n19590), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n9904) );
  NAND2_X1 U11636 ( .A1(n19472), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n9902) );
  AND2_X1 U11637 ( .A1(n12049), .A2(n12048), .ZN(n12052) );
  NAND2_X1 U11638 ( .A1(n12051), .A2(n12050), .ZN(n12082) );
  INV_X1 U11639 ( .A(n11976), .ZN(n10007) );
  NAND2_X1 U11640 ( .A1(n20171), .A2(n20176), .ZN(n12551) );
  NAND2_X1 U11641 ( .A1(n9891), .A2(n11855), .ZN(n11857) );
  NOR2_X1 U11642 ( .A1(n11092), .A2(n11071), .ZN(n11076) );
  NAND2_X1 U11643 ( .A1(n15415), .A2(n9920), .ZN(n9919) );
  INV_X1 U11644 ( .A(n9917), .ZN(n9916) );
  OAI21_X1 U11645 ( .B1(n9918), .B2(n11109), .A(n9921), .ZN(n9917) );
  AND2_X1 U11646 ( .A1(n16107), .A2(n15158), .ZN(n9921) );
  OAI21_X1 U11647 ( .B1(n19409), .B2(n11570), .A(n9876), .ZN(n11011) );
  AND2_X2 U11648 ( .A1(n9906), .A2(n10812), .ZN(n10212) );
  NAND2_X1 U11649 ( .A1(n10811), .A2(n14257), .ZN(n10812) );
  AND2_X1 U11650 ( .A1(n10755), .A2(n19170), .ZN(n10780) );
  NOR2_X1 U11651 ( .A1(n17366), .A2(n10333), .ZN(n10332) );
  NOR2_X1 U11652 ( .A1(n17373), .A2(n10354), .ZN(n10359) );
  NAND2_X1 U11653 ( .A1(n10508), .A2(n10348), .ZN(n10354) );
  AND2_X1 U11654 ( .A1(n12813), .A2(n11845), .ZN(n12603) );
  NAND2_X1 U11655 ( .A1(n13352), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12509) );
  INV_X1 U11656 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12101) );
  INV_X1 U11657 ( .A(n11988), .ZN(n12534) );
  INV_X1 U11658 ( .A(n12765), .ZN(n10094) );
  NOR2_X1 U11659 ( .A1(n12610), .A2(n12609), .ZN(n12692) );
  NOR2_X1 U11660 ( .A1(n10101), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10097) );
  INV_X1 U11661 ( .A(n11993), .ZN(n10101) );
  NAND2_X1 U11662 ( .A1(n10004), .A2(n11993), .ZN(n10003) );
  NAND2_X1 U11663 ( .A1(n10102), .A2(n11925), .ZN(n10004) );
  OR2_X1 U11664 ( .A1(n11937), .A2(n12009), .ZN(n11887) );
  NAND2_X1 U11666 ( .A1(n20399), .A2(n20708), .ZN(n9896) );
  AOI21_X1 U11667 ( .B1(n11145), .B2(n11125), .A(n11126), .ZN(n11137) );
  NAND2_X1 U11668 ( .A1(n11076), .A2(n11105), .ZN(n11104) );
  INV_X1 U11669 ( .A(n10051), .ZN(n11083) );
  NAND2_X1 U11670 ( .A1(n9755), .A2(n10901), .ZN(n10043) );
  NOR2_X1 U11671 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14115) );
  OR2_X1 U11672 ( .A1(n14274), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14141) );
  NAND2_X1 U11673 ( .A1(n10694), .A2(n10693), .ZN(n10725) );
  CLKBUF_X1 U11674 ( .A(n10663), .Z(n14236) );
  NAND2_X1 U11675 ( .A1(n9856), .A2(n14986), .ZN(n10156) );
  AND2_X1 U11676 ( .A1(n10162), .A2(n10161), .ZN(n10160) );
  INV_X1 U11677 ( .A(n15015), .ZN(n10161) );
  AND2_X1 U11678 ( .A1(n13532), .A2(n13520), .ZN(n10205) );
  NAND2_X1 U11679 ( .A1(n10191), .A2(n13416), .ZN(n10190) );
  INV_X1 U11680 ( .A(n13389), .ZN(n10191) );
  XNOR2_X1 U11681 ( .A(n10725), .B(n10726), .ZN(n10748) );
  INV_X1 U11682 ( .A(n14973), .ZN(n10207) );
  INV_X1 U11683 ( .A(n14980), .ZN(n10208) );
  OR3_X1 U11684 ( .A1(n16041), .A2(n14045), .A3(n15317), .ZN(n11156) );
  INV_X1 U11685 ( .A(n14940), .ZN(n10201) );
  NOR2_X1 U11686 ( .A1(n14015), .A2(n10183), .ZN(n10182) );
  INV_X1 U11687 ( .A(n12911), .ZN(n10183) );
  AND2_X1 U11688 ( .A1(n10205), .A2(n10204), .ZN(n10203) );
  INV_X1 U11689 ( .A(n13648), .ZN(n10204) );
  INV_X1 U11690 ( .A(n15255), .ZN(n9914) );
  NOR2_X1 U11691 ( .A1(n10217), .A2(n15460), .ZN(n10216) );
  INV_X1 U11692 ( .A(n11045), .ZN(n10217) );
  NOR2_X1 U11693 ( .A1(n10173), .A2(n11469), .ZN(n10172) );
  INV_X1 U11694 ( .A(n13160), .ZN(n10173) );
  INV_X1 U11695 ( .A(n16185), .ZN(n10148) );
  NOR2_X1 U11696 ( .A1(n10190), .A2(n13456), .ZN(n10192) );
  AOI21_X1 U11697 ( .B1(n10740), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10729), .ZN(n10736) );
  NAND2_X1 U11698 ( .A1(n9928), .A2(n9730), .ZN(n9927) );
  NAND2_X1 U11699 ( .A1(n19218), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9882) );
  OR2_X1 U11700 ( .A1(n10857), .A2(n10856), .ZN(n11665) );
  INV_X1 U11701 ( .A(n11588), .ZN(n11608) );
  AND2_X1 U11702 ( .A1(n11181), .A2(n11180), .ZN(n11232) );
  NOR2_X1 U11703 ( .A1(n9796), .A2(n10283), .ZN(n10284) );
  NAND2_X1 U11704 ( .A1(n10309), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n9947) );
  NOR2_X1 U11705 ( .A1(n10304), .A2(n10303), .ZN(n10305) );
  OAI21_X1 U11706 ( .B1(n10301), .B2(n20876), .A(n10302), .ZN(n10303) );
  NOR3_X1 U11707 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n18685), .ZN(n10395) );
  NAND2_X1 U11708 ( .A1(n9769), .A2(n9999), .ZN(n9998) );
  AND2_X1 U11709 ( .A1(n10001), .A2(n10000), .ZN(n9999) );
  INV_X1 U11710 ( .A(n17655), .ZN(n10000) );
  INV_X1 U11711 ( .A(n10361), .ZN(n9953) );
  NAND2_X1 U11712 ( .A1(n10332), .A2(n17362), .ZN(n10364) );
  NAND2_X1 U11713 ( .A1(n17570), .A2(n9814), .ZN(n10074) );
  NAND2_X1 U11714 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n10372), .ZN(
        n18053) );
  AOI21_X1 U11715 ( .B1(n17358), .B2(n10364), .A(n17765), .ZN(n10367) );
  OAI21_X1 U11716 ( .B1(n10502), .B2(n10482), .A(n10501), .ZN(n12707) );
  INV_X1 U11717 ( .A(n9977), .ZN(n9976) );
  NAND2_X1 U11718 ( .A1(n20798), .A2(n13614), .ZN(n14417) );
  NAND2_X1 U11719 ( .A1(n14417), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14475) );
  INV_X1 U11720 ( .A(n12273), .ZN(n12820) );
  AND2_X1 U11721 ( .A1(n12489), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12490) );
  AND2_X1 U11722 ( .A1(n9841), .A2(n14389), .ZN(n10130) );
  NAND2_X1 U11723 ( .A1(n12452), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12488) );
  NAND2_X1 U11724 ( .A1(n12341), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12362) );
  NOR2_X1 U11725 ( .A1(n10125), .A2(n10124), .ZN(n10123) );
  NAND2_X1 U11726 ( .A1(n9894), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12793) );
  INV_X1 U11727 ( .A(n13737), .ZN(n9894) );
  NAND2_X1 U11728 ( .A1(n13739), .A2(n12792), .ZN(n10120) );
  NAND2_X1 U11729 ( .A1(n13438), .A2(n13439), .ZN(n13468) );
  NOR2_X1 U11730 ( .A1(n10030), .A2(n14380), .ZN(n10027) );
  NAND2_X1 U11731 ( .A1(n10031), .A2(n14353), .ZN(n10030) );
  INV_X1 U11732 ( .A(n14391), .ZN(n10031) );
  NAND2_X1 U11733 ( .A1(n10024), .A2(n12688), .ZN(n10023) );
  AND2_X1 U11734 ( .A1(n10026), .A2(n14401), .ZN(n10025) );
  INV_X1 U11735 ( .A(n10028), .ZN(n10026) );
  OR2_X1 U11737 ( .A1(n14838), .A2(n14844), .ZN(n14819) );
  INV_X1 U11738 ( .A(n10107), .ZN(n9961) );
  AND2_X1 U11739 ( .A1(n12772), .A2(n12771), .ZN(n15838) );
  INV_X1 U11740 ( .A(n15846), .ZN(n12762) );
  NAND2_X1 U11741 ( .A1(n20077), .A2(n20092), .ZN(n10118) );
  INV_X1 U11742 ( .A(n13445), .ZN(n10013) );
  INV_X1 U11743 ( .A(n13444), .ZN(n10014) );
  NOR2_X1 U11744 ( .A1(n13150), .A2(n14343), .ZN(n20086) );
  OAI221_X1 U11745 ( .B1(n15602), .B2(n15976), .C1(n15602), .C2(n15981), .A(
        n20708), .ZN(n20294) );
  INV_X1 U11746 ( .A(n19894), .ZN(n13129) );
  NAND2_X1 U11747 ( .A1(n13374), .A2(n13373), .ZN(n20651) );
  AND2_X1 U11748 ( .A1(n11147), .A2(n14984), .ZN(n11149) );
  AND2_X1 U11749 ( .A1(n11139), .A2(n11138), .ZN(n11147) );
  AND2_X1 U11750 ( .A1(n11345), .A2(n11344), .ZN(n14967) );
  AND2_X1 U11751 ( .A1(n14207), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13383) );
  OAI21_X1 U11752 ( .B1(n10748), .B2(n10749), .A(n10727), .ZN(n9923) );
  OR2_X1 U11753 ( .A1(n10726), .A2(n10725), .ZN(n10727) );
  NOR2_X1 U11754 ( .A1(n10688), .A2(n11034), .ZN(n10186) );
  NAND2_X1 U11755 ( .A1(n10135), .A2(n14254), .ZN(n14957) );
  NAND2_X1 U11756 ( .A1(n14970), .A2(n10228), .ZN(n10135) );
  NAND2_X1 U11757 ( .A1(n9987), .A2(n10614), .ZN(n9986) );
  NAND2_X1 U11758 ( .A1(n9989), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9988) );
  NOR2_X1 U11759 ( .A1(n10657), .A2(n19884), .ZN(n13017) );
  INV_X1 U11760 ( .A(n13811), .ZN(n13812) );
  OR2_X1 U11761 ( .A1(n14993), .A2(n14994), .ZN(n14996) );
  AND2_X1 U11762 ( .A1(n13493), .A2(n13492), .ZN(n13533) );
  AOI21_X1 U11763 ( .B1(n10050), .B2(n9767), .A(n10046), .ZN(n10045) );
  INV_X1 U11764 ( .A(n14047), .ZN(n14046) );
  AND2_X1 U11765 ( .A1(n11320), .A2(n11319), .ZN(n14925) );
  NOR2_X1 U11766 ( .A1(n13639), .A2(n13640), .ZN(n13638) );
  NAND2_X1 U11767 ( .A1(n13465), .A2(n13464), .ZN(n13472) );
  AND2_X1 U11768 ( .A1(n11060), .A2(n15470), .ZN(n15460) );
  AND2_X1 U11769 ( .A1(n11046), .A2(n10216), .ZN(n15458) );
  INV_X1 U11770 ( .A(n15246), .ZN(n10151) );
  NOR2_X1 U11771 ( .A1(n13487), .A2(n13488), .ZN(n13492) );
  NAND2_X1 U11772 ( .A1(n16347), .A2(n9929), .ZN(n11645) );
  CLKBUF_X1 U11773 ( .A(n11646), .Z(n11647) );
  NAND2_X1 U11774 ( .A1(n19170), .A2(n16345), .ZN(n13015) );
  INV_X1 U11775 ( .A(n19472), .ZN(n19469) );
  INV_X1 U11776 ( .A(n16352), .ZN(n13542) );
  INV_X1 U11777 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19871) );
  NAND2_X1 U11778 ( .A1(n11234), .A2(n11233), .ZN(n16315) );
  NAND2_X1 U11779 ( .A1(n11232), .A2(n12937), .ZN(n11233) );
  AND2_X1 U11780 ( .A1(n19884), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16345) );
  INV_X1 U11781 ( .A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n20841) );
  INV_X2 U11782 ( .A(n9794), .ZN(n17180) );
  INV_X1 U11783 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n20882) );
  NOR2_X1 U11784 ( .A1(n13910), .A2(n15537), .ZN(n15641) );
  NOR3_X1 U11785 ( .A1(n13907), .A2(n13906), .A3(n17218), .ZN(n13910) );
  AOI21_X1 U11786 ( .B1(n16507), .B2(n9807), .A(n15539), .ZN(n15643) );
  NOR2_X1 U11787 ( .A1(n17513), .A2(n17514), .ZN(n12713) );
  NOR2_X1 U11788 ( .A1(n17625), .A2(n9860), .ZN(n17608) );
  NOR2_X1 U11789 ( .A1(n9998), .A2(n17746), .ZN(n17640) );
  NAND2_X1 U11790 ( .A1(n17680), .A2(n10369), .ZN(n10370) );
  AND2_X1 U11791 ( .A1(n17731), .A2(n10082), .ZN(n10081) );
  NOR2_X1 U11792 ( .A1(n18227), .A2(n10537), .ZN(n10545) );
  INV_X1 U11793 ( .A(n12707), .ZN(n18649) );
  NAND2_X1 U11794 ( .A1(n18656), .A2(n18657), .ZN(n16507) );
  NOR2_X1 U11795 ( .A1(n10431), .A2(n9936), .ZN(n18204) );
  OR2_X1 U11796 ( .A1(n10432), .A2(n9937), .ZN(n9936) );
  AND2_X1 U11797 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n9937) );
  INV_X1 U11798 ( .A(n18713), .ZN(n18862) );
  INV_X1 U11799 ( .A(n20015), .ZN(n15768) );
  XNOR2_X1 U11800 ( .A(n14655), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14814) );
  NAND2_X1 U11801 ( .A1(n13149), .A2(n13138), .ZN(n20109) );
  OR2_X1 U11802 ( .A1(n11707), .A2(n11706), .ZN(n12928) );
  OR2_X1 U11803 ( .A1(n19148), .A2(n19144), .ZN(n19150) );
  NAND2_X1 U11804 ( .A1(n10236), .A2(n10197), .ZN(n10196) );
  AOI21_X1 U11805 ( .B1(n12896), .B2(n16198), .A(n10198), .ZN(n10197) );
  NAND2_X1 U11806 ( .A1(n11713), .A2(n11714), .ZN(n10198) );
  INV_X1 U11807 ( .A(n15403), .ZN(n10167) );
  AND2_X1 U11808 ( .A1(n16204), .A2(n19847), .ZN(n19171) );
  AOI21_X1 U11809 ( .B1(n15993), .B2(n19192), .A(n10170), .ZN(n10169) );
  NAND2_X1 U11810 ( .A1(n15992), .A2(n19186), .ZN(n9932) );
  OR2_X1 U11811 ( .A1(n11660), .A2(n10171), .ZN(n10170) );
  INV_X1 U11812 ( .A(n19186), .ZN(n16289) );
  INV_X1 U11813 ( .A(n16305), .ZN(n19187) );
  INV_X1 U11814 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19872) );
  INV_X1 U11815 ( .A(n19248), .ZN(n19857) );
  NAND2_X1 U11816 ( .A1(n13223), .A2(n13077), .ZN(n19848) );
  OR2_X1 U11817 ( .A1(n13076), .A2(n13075), .ZN(n13077) );
  AND2_X1 U11818 ( .A1(n13307), .A2(n13227), .ZN(n19282) );
  INV_X1 U11819 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19884) );
  NAND2_X1 U11820 ( .A1(n16667), .A2(n10002), .ZN(n16638) );
  NAND2_X1 U11821 ( .A1(n16525), .A2(n9860), .ZN(n10002) );
  NOR2_X1 U11822 ( .A1(n16995), .A2(n16994), .ZN(n16979) );
  NAND2_X1 U11823 ( .A1(n17330), .A2(P3_EAX_REG_15__SCAN_IN), .ZN(n17321) );
  XNOR2_X1 U11824 ( .A(n15549), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16383) );
  OAI21_X1 U11825 ( .B1(n16382), .B2(n16381), .A(n10085), .ZN(n10084) );
  AOI22_X1 U11826 ( .A1(n10087), .A2(n10086), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16385), .ZN(n10085) );
  NAND2_X1 U11827 ( .A1(n16386), .A2(n16387), .ZN(n10086) );
  NOR2_X2 U11828 ( .A1(n17358), .A2(n17860), .ZN(n17766) );
  AND2_X1 U11829 ( .A1(n12556), .A2(n12538), .ZN(n12564) );
  INV_X1 U11830 ( .A(n12565), .ZN(n12542) );
  NOR2_X1 U11831 ( .A1(n12573), .A2(n12574), .ZN(n12572) );
  AND2_X1 U11832 ( .A1(n12597), .A2(n13136), .ZN(n11861) );
  NOR2_X1 U11833 ( .A1(n11861), .A2(n11870), .ZN(n11852) );
  NOR2_X1 U11834 ( .A1(n11853), .A2(n20708), .ZN(n9888) );
  INV_X1 U11835 ( .A(n19559), .ZN(n10995) );
  NAND3_X1 U11836 ( .A1(n10212), .A2(n10213), .A3(n11435), .ZN(n10981) );
  AOI22_X1 U11837 ( .A1(n19559), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10781), .B2(n9924), .ZN(n10826) );
  AND2_X1 U11838 ( .A1(n10763), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9924) );
  NAND2_X1 U11839 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n9940) );
  AOI21_X1 U11840 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20488), .A(
        n12572), .ZN(n12544) );
  AND3_X1 U11841 ( .A1(n12571), .A2(n12570), .A3(n12569), .ZN(n12578) );
  OR2_X1 U11842 ( .A1(n12072), .A2(n12071), .ZN(n12768) );
  OR2_X1 U11843 ( .A1(n11923), .A2(n11922), .ZN(n12730) );
  OR2_X1 U11844 ( .A1(n11886), .A2(n11885), .ZN(n12731) );
  INV_X1 U11845 ( .A(n11975), .ZN(n10008) );
  AND2_X1 U11846 ( .A1(n11978), .A2(n20176), .ZN(n11848) );
  AOI22_X1 U11848 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14290) );
  AOI22_X1 U11849 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14283) );
  AOI22_X1 U11850 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14249) );
  AOI22_X1 U11851 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14242) );
  AOI22_X1 U11852 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14219) );
  INV_X1 U11853 ( .A(n14163), .ZN(n10158) );
  AOI22_X1 U11854 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14203) );
  AOI22_X1 U11855 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14196) );
  AOI22_X1 U11856 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14179) );
  AOI22_X1 U11857 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14172) );
  AOI21_X1 U11858 ( .B1(n14236), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A(n9864), .ZN(n14124) );
  AOI22_X1 U11859 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U11860 ( .A1(n11663), .A2(n11686), .ZN(n11662) );
  NOR2_X1 U11861 ( .A1(n10673), .A2(n10689), .ZN(n10674) );
  NAND2_X1 U11862 ( .A1(n10699), .A2(n9726), .ZN(n10681) );
  NOR2_X1 U11863 ( .A1(n10657), .A2(n11034), .ZN(n10679) );
  OR2_X1 U11864 ( .A1(n10483), .A2(n10486), .ZN(n10502) );
  OAI211_X1 U11865 ( .C1(n17170), .C2(n17120), .A(n9979), .B(n9978), .ZN(n9977) );
  NAND2_X1 U11866 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n9978) );
  AOI21_X1 U11867 ( .B1(n9722), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(n9980), .ZN(n9979) );
  NOR2_X1 U11868 ( .A1(n17188), .A2(n20882), .ZN(n9980) );
  AND2_X1 U11869 ( .A1(n12582), .A2(n12786), .ZN(n12586) );
  INV_X1 U11870 ( .A(n14531), .ZN(n10126) );
  NOR2_X1 U11871 ( .A1(n14542), .A2(n10128), .ZN(n10127) );
  INV_X1 U11872 ( .A(n14546), .ZN(n10128) );
  NAND2_X1 U11873 ( .A1(n9786), .A2(n9846), .ZN(n10125) );
  NAND2_X1 U11874 ( .A1(n10122), .A2(n12165), .ZN(n13862) );
  INV_X1 U11875 ( .A(n13719), .ZN(n10129) );
  INV_X1 U11876 ( .A(n13609), .ZN(n12130) );
  XNOR2_X1 U11877 ( .A(n12789), .B(n12109), .ZN(n12776) );
  INV_X1 U11878 ( .A(n13503), .ZN(n12114) );
  NOR2_X1 U11879 ( .A1(n11971), .A2(n11970), .ZN(n12741) );
  OR2_X1 U11880 ( .A1(n14380), .A2(n14391), .ZN(n10028) );
  INV_X1 U11881 ( .A(n14644), .ZN(n10106) );
  OR2_X1 U11882 ( .A1(n9738), .A2(n14687), .ZN(n10107) );
  INV_X1 U11883 ( .A(n14517), .ZN(n10032) );
  NAND2_X1 U11884 ( .A1(n14707), .A2(n14708), .ZN(n10005) );
  INV_X1 U11885 ( .A(n13894), .ZN(n10020) );
  NOR2_X1 U11886 ( .A1(n13875), .A2(n10022), .ZN(n10021) );
  INV_X1 U11887 ( .A(n13886), .ZN(n10022) );
  OR2_X1 U11888 ( .A1(n12047), .A2(n12046), .ZN(n12756) );
  INV_X1 U11889 ( .A(n13141), .ZN(n12670) );
  NAND2_X1 U11890 ( .A1(n12670), .A2(n12610), .ZN(n12673) );
  INV_X1 U11891 ( .A(n12730), .ZN(n12727) );
  INV_X1 U11892 ( .A(n12582), .ZN(n12568) );
  INV_X1 U11893 ( .A(n11938), .ZN(n11939) );
  AND2_X1 U11894 ( .A1(n12813), .A2(n20144), .ZN(n9962) );
  OAI211_X1 U11895 ( .C1(n20146), .C2(n12831), .A(n11954), .B(n11953), .ZN(
        n11955) );
  NAND2_X1 U11896 ( .A1(n11874), .A2(n11873), .ZN(n20197) );
  NAND2_X1 U11897 ( .A1(n11822), .A2(n11823), .ZN(n10017) );
  AND2_X1 U11898 ( .A1(n11764), .A2(n11765), .ZN(n11768) );
  INV_X1 U11899 ( .A(n20803), .ZN(n13117) );
  NAND2_X1 U11900 ( .A1(n11145), .A2(n14041), .ZN(n11153) );
  NAND2_X1 U11901 ( .A1(n11050), .A2(n13495), .ZN(n11053) );
  NAND2_X1 U11902 ( .A1(n10987), .A2(n9768), .ZN(n11042) );
  INV_X1 U11903 ( .A(n10935), .ZN(n10984) );
  NAND2_X1 U11904 ( .A1(n11272), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U11905 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14270) );
  AOI22_X1 U11906 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14263) );
  NOR2_X1 U11907 ( .A1(n15343), .A2(n10180), .ZN(n10179) );
  INV_X1 U11908 ( .A(n14921), .ZN(n10180) );
  NAND2_X1 U11909 ( .A1(n13635), .A2(n9845), .ZN(n15004) );
  AND2_X1 U11910 ( .A1(n13850), .A2(n13634), .ZN(n10162) );
  AND2_X1 U11911 ( .A1(n13851), .A2(n13849), .ZN(n13850) );
  AOI22_X1 U11912 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9764), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10613) );
  OR2_X1 U11913 ( .A1(n10976), .A2(n10975), .ZN(n11440) );
  NOR2_X1 U11914 ( .A1(n15133), .A2(n10062), .ZN(n10061) );
  INV_X1 U11915 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U11916 ( .A1(n15182), .A2(n10059), .ZN(n10058) );
  INV_X1 U11917 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10059) );
  NOR2_X1 U11918 ( .A1(n16146), .A2(n10055), .ZN(n10054) );
  INV_X1 U11919 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U11920 ( .A1(n16205), .A2(n10069), .ZN(n10072) );
  NOR2_X1 U11921 ( .A1(n15317), .A2(n15335), .ZN(n9935) );
  AND2_X1 U11922 ( .A1(n10179), .A2(n15091), .ZN(n10178) );
  NAND2_X1 U11923 ( .A1(n10035), .A2(n10034), .ZN(n9990) );
  AOI21_X1 U11924 ( .B1(n16107), .B2(n10037), .A(n10036), .ZN(n10034) );
  NAND2_X1 U11925 ( .A1(n9919), .A2(n9916), .ZN(n10035) );
  INV_X1 U11926 ( .A(n11639), .ZN(n11632) );
  NOR2_X1 U11927 ( .A1(n13814), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11404) );
  INV_X1 U11928 ( .A(n9928), .ZN(n10719) );
  NAND2_X1 U11929 ( .A1(n11195), .A2(n9808), .ZN(n9929) );
  NAND2_X1 U11930 ( .A1(n13013), .A2(n19871), .ZN(n13301) );
  AND2_X1 U11931 ( .A1(n14207), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13217) );
  OR2_X1 U11932 ( .A1(n13071), .A2(n13072), .ZN(n13221) );
  NOR2_X1 U11933 ( .A1(n10779), .A2(n10776), .ZN(n19249) );
  NAND2_X1 U11934 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10637) );
  NAND2_X1 U11935 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10631) );
  INV_X1 U11936 ( .A(n10768), .ZN(n10761) );
  NAND3_X1 U11937 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19825), .A3(n19651), 
        .ZN(n13551) );
  AND2_X1 U11938 ( .A1(n19861), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11184) );
  NAND2_X1 U11939 ( .A1(n11230), .A2(n11229), .ZN(n11234) );
  NOR3_X2 U11940 ( .A1(n18826), .A2(n18819), .A3(n16867), .ZN(n10287) );
  INV_X1 U11941 ( .A(n16647), .ZN(n10001) );
  INV_X1 U11942 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10079) );
  NOR2_X1 U11943 ( .A1(n17775), .A2(n18106), .ZN(n10529) );
  OR2_X1 U11944 ( .A1(n18240), .A2(n17392), .ZN(n10497) );
  NAND2_X1 U11945 ( .A1(n17454), .A2(n10550), .ZN(n16508) );
  AOI21_X1 U11946 ( .B1(n10548), .B2(n10547), .A(n10546), .ZN(n10551) );
  NOR4_X1 U11947 ( .A1(n10548), .A2(n13906), .A3(n10497), .A4(n10496), .ZN(
        n10549) );
  INV_X1 U11948 ( .A(n10429), .ZN(n9943) );
  NOR2_X1 U11949 ( .A1(n10489), .A2(n10498), .ZN(n16392) );
  NAND2_X1 U11950 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18666) );
  OR2_X1 U11951 ( .A1(n14882), .A2(n12601), .ZN(n14343) );
  INV_X1 U11952 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15722) );
  NAND2_X1 U11953 ( .A1(n12131), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12156) );
  INV_X1 U11954 ( .A(n19989), .ZN(n15647) );
  NOR2_X1 U11955 ( .A1(n14390), .A2(n10028), .ZN(n14379) );
  OR2_X1 U11956 ( .A1(n14458), .A2(n14442), .ZN(n14551) );
  NAND2_X1 U11957 ( .A1(n13097), .A2(n13162), .ZN(n10018) );
  AOI21_X1 U11958 ( .B1(n12754), .B2(n12231), .A(n12081), .ZN(n13467) );
  OAI21_X1 U11959 ( .B1(n12055), .B2(n14634), .A(n12511), .ZN(n14378) );
  NOR2_X1 U11960 ( .A1(n12451), .A2(n15650), .ZN(n12452) );
  OAI21_X1 U11961 ( .B1(n12055), .B2(n14657), .A(n12471), .ZN(n14404) );
  AOI21_X1 U11962 ( .B1(n12450), .B2(n12449), .A(n12448), .ZN(n14498) );
  AND2_X1 U11963 ( .A1(n12431), .A2(n12430), .ZN(n14510) );
  OR2_X1 U11964 ( .A1(n15672), .A2(n12055), .ZN(n12430) );
  INV_X1 U11965 ( .A(n14414), .ZN(n12407) );
  NOR2_X1 U11966 ( .A1(n12362), .A2(n12361), .ZN(n12363) );
  NAND2_X1 U11967 ( .A1(n12363), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12424) );
  AOI21_X1 U11968 ( .B1(n12360), .B2(n12359), .A(n12358), .ZN(n14524) );
  AND2_X1 U11969 ( .A1(n13611), .A2(n15681), .ZN(n12358) );
  CLKBUF_X1 U11970 ( .A(n14522), .Z(n14523) );
  AND2_X1 U11971 ( .A1(n12306), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12307) );
  NAND2_X1 U11972 ( .A1(n12307), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12340) );
  NAND2_X1 U11973 ( .A1(n14547), .A2(n14546), .ZN(n14549) );
  NAND2_X1 U11974 ( .A1(n12261), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12262) );
  NOR2_X1 U11975 ( .A1(n20990), .A2(n12262), .ZN(n12306) );
  NOR2_X1 U11976 ( .A1(n12241), .A2(n15722), .ZN(n12261) );
  OR2_X1 U11977 ( .A1(n12222), .A2(n15730), .ZN(n12241) );
  INV_X1 U11978 ( .A(n13900), .ZN(n12239) );
  NAND2_X1 U11979 ( .A1(n12217), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12222) );
  INV_X1 U11980 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n21034) );
  NOR2_X1 U11981 ( .A1(n21034), .A2(n12191), .ZN(n12217) );
  AND2_X1 U11982 ( .A1(n12160), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12161) );
  NAND2_X1 U11983 ( .A1(n12161), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12191) );
  NOR2_X1 U11984 ( .A1(n12156), .A2(n19919), .ZN(n12160) );
  NAND2_X1 U11985 ( .A1(n12110), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12126) );
  NOR2_X1 U11986 ( .A1(n12097), .A2(n12101), .ZN(n12110) );
  NOR2_X2 U11987 ( .A1(n13468), .A2(n13467), .ZN(n13499) );
  NAND2_X1 U11988 ( .A1(n12104), .A2(n12103), .ZN(n13498) );
  NAND2_X1 U11989 ( .A1(n12077), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12097) );
  INV_X1 U11990 ( .A(n12076), .ZN(n12077) );
  NAND2_X1 U11991 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12029) );
  NOR2_X1 U11992 ( .A1(n12029), .A2(n12028), .ZN(n12054) );
  INV_X1 U11993 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12028) );
  NAND2_X1 U11994 ( .A1(n12027), .A2(n12231), .ZN(n12036) );
  NAND2_X1 U11995 ( .A1(n12003), .A2(n12002), .ZN(n13334) );
  INV_X1 U11996 ( .A(n13336), .ZN(n12002) );
  INV_X1 U11997 ( .A(n13337), .ZN(n12003) );
  NOR2_X1 U11998 ( .A1(n15794), .A2(n14795), .ZN(n10111) );
  NAND2_X1 U11999 ( .A1(n9885), .A2(n14783), .ZN(n14626) );
  INV_X1 U12000 ( .A(n14662), .ZN(n9899) );
  OR2_X1 U12001 ( .A1(n14390), .A2(n14391), .ZN(n14393) );
  NAND2_X1 U12002 ( .A1(n14541), .A2(n9781), .ZN(n14519) );
  NAND2_X1 U12003 ( .A1(n14541), .A2(n9835), .ZN(n14528) );
  NAND2_X1 U12004 ( .A1(n10110), .A2(n10109), .ZN(n10108) );
  NOR3_X1 U12005 ( .A1(n15607), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U12006 ( .A1(n10005), .A2(n9770), .ZN(n15792) );
  OR2_X1 U12007 ( .A1(n14560), .A2(n14456), .ZN(n14458) );
  NOR2_X1 U12008 ( .A1(n15805), .A2(n15804), .ZN(n14708) );
  AND2_X1 U12009 ( .A1(n15893), .A2(n14761), .ZN(n14857) );
  AND2_X1 U12010 ( .A1(n15794), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15804) );
  NAND2_X1 U12011 ( .A1(n15760), .A2(n10021), .ZN(n13895) );
  NAND2_X1 U12012 ( .A1(n15760), .A2(n13886), .ZN(n13888) );
  AND2_X1 U12013 ( .A1(n15758), .A2(n15757), .ZN(n15760) );
  AND2_X1 U12014 ( .A1(n12641), .A2(n12640), .ZN(n13727) );
  CLKBUF_X1 U12015 ( .A(n14705), .Z(n14706) );
  OR2_X1 U12016 ( .A1(n15935), .A2(n15934), .ZN(n15937) );
  OR2_X1 U12017 ( .A1(n13506), .A2(n13621), .ZN(n15935) );
  NOR2_X1 U12018 ( .A1(n15794), .A2(n9840), .ZN(n13737) );
  NOR2_X1 U12019 ( .A1(n15967), .A2(n13500), .ZN(n13508) );
  AND2_X1 U12020 ( .A1(n12632), .A2(n12631), .ZN(n13507) );
  NAND2_X1 U12021 ( .A1(n12773), .A2(n10094), .ZN(n10093) );
  INV_X1 U12022 ( .A(n12773), .ZN(n10095) );
  NOR2_X1 U12023 ( .A1(n13339), .A2(n13338), .ZN(n13406) );
  AND2_X1 U12024 ( .A1(n13120), .A2(n11849), .ZN(n11838) );
  NAND2_X1 U12025 ( .A1(n13130), .A2(n13129), .ZN(n13150) );
  INV_X1 U12026 ( .A(n10100), .ZN(n10099) );
  INV_X1 U12027 ( .A(n13372), .ZN(n13374) );
  NAND2_X1 U12028 ( .A1(n12007), .A2(n12006), .ZN(n20288) );
  OR2_X1 U12029 ( .A1(n11951), .A2(n12543), .ZN(n12007) );
  CLKBUF_X1 U12030 ( .A(n11728), .Z(n14884) );
  INV_X1 U12031 ( .A(n14879), .ZN(n13352) );
  NAND2_X1 U12032 ( .A1(n20137), .A2(n13372), .ZN(n20262) );
  NOR2_X1 U12033 ( .A1(n13372), .A2(n13373), .ZN(n20370) );
  NAND2_X1 U12034 ( .A1(n20223), .A2(n20222), .ZN(n20455) );
  INV_X1 U12035 ( .A(n20493), .ZN(n20487) );
  INV_X1 U12036 ( .A(n20294), .ZN(n20185) );
  INV_X1 U12037 ( .A(n20170), .ZN(n20187) );
  AND2_X1 U12038 ( .A1(n14351), .A2(n13131), .ZN(n15590) );
  INV_X1 U12039 ( .A(n14351), .ZN(n14342) );
  NAND2_X1 U12040 ( .A1(n10871), .A2(n10702), .ZN(n10041) );
  NAND2_X1 U12041 ( .A1(n10042), .A2(n10702), .ZN(n10040) );
  AND2_X1 U12042 ( .A1(n11137), .A2(n11136), .ZN(n11139) );
  NAND2_X1 U12043 ( .A1(n10066), .A2(n9815), .ZN(n15560) );
  NOR2_X1 U12044 ( .A1(n10064), .A2(n10068), .ZN(n10063) );
  NAND2_X1 U12045 ( .A1(n11124), .A2(n15013), .ZN(n11125) );
  INV_X1 U12046 ( .A(n11123), .ZN(n11124) );
  AND2_X1 U12047 ( .A1(n10066), .A2(n9776), .ZN(n14935) );
  NOR2_X1 U12048 ( .A1(n14900), .A2(n18924), .ZN(n14904) );
  NAND2_X1 U12049 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n14901), .ZN(
        n14900) );
  NAND2_X1 U12050 ( .A1(n10051), .A2(n9844), .ZN(n11092) );
  AND2_X1 U12051 ( .A1(n11085), .A2(n11084), .ZN(n18949) );
  NAND2_X1 U12052 ( .A1(n11062), .A2(n11063), .ZN(n11089) );
  NAND2_X1 U12053 ( .A1(n11145), .A2(n11064), .ZN(n11062) );
  AND2_X1 U12054 ( .A1(n10987), .A2(n10986), .ZN(n11036) );
  NAND2_X1 U12055 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12884) );
  AND2_X1 U12056 ( .A1(n11312), .A2(n11311), .ZN(n15021) );
  OR2_X1 U12057 ( .A1(n11486), .A2(n11485), .ZN(n13518) );
  AND2_X1 U12058 ( .A1(n13383), .A2(n9868), .ZN(n10152) );
  NOR2_X1 U12059 ( .A1(n15067), .A2(n9789), .ZN(n15048) );
  NOR3_X1 U12060 ( .A1(n10176), .A2(n9789), .A3(n10177), .ZN(n10175) );
  INV_X1 U12061 ( .A(n15065), .ZN(n10176) );
  AOI21_X1 U12062 ( .B1(n14236), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A(n9870), .ZN(n14317) );
  AOI22_X1 U12063 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10038), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14301) );
  NAND2_X1 U12064 ( .A1(n10139), .A2(n10141), .ZN(n14953) );
  OAI21_X1 U12065 ( .B1(n14254), .B2(n10140), .A(n14958), .ZN(n10137) );
  NOR2_X1 U12066 ( .A1(n10134), .A2(n10140), .ZN(n10138) );
  XNOR2_X1 U12067 ( .A(n14213), .B(n14209), .ZN(n14979) );
  NAND2_X1 U12068 ( .A1(n13635), .A2(n10162), .ZN(n15016) );
  INV_X1 U12069 ( .A(n11231), .ZN(n12937) );
  NAND2_X1 U12070 ( .A1(n15985), .A2(n9790), .ZN(n15122) );
  AND2_X1 U12071 ( .A1(n15985), .A2(n10060), .ZN(n15121) );
  AND2_X1 U12072 ( .A1(n9790), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10060) );
  NAND2_X1 U12073 ( .A1(n15985), .A2(n10061), .ZN(n15131) );
  NAND2_X1 U12074 ( .A1(n15985), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15144) );
  NOR3_X1 U12075 ( .A1(n14996), .A2(n10208), .A3(n14909), .ZN(n14983) );
  NOR2_X1 U12076 ( .A1(n15986), .A2(n16097), .ZN(n15985) );
  NAND2_X1 U12077 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n14896), .ZN(
        n15986) );
  NOR2_X1 U12078 ( .A1(n14996), .A2(n14909), .ZN(n14981) );
  AND2_X1 U12079 ( .A1(n14906), .A2(n10057), .ZN(n14896) );
  AND2_X1 U12080 ( .A1(n9791), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10057) );
  NAND2_X1 U12081 ( .A1(n14906), .A2(n9791), .ZN(n14907) );
  AND2_X1 U12082 ( .A1(n11316), .A2(n11315), .ZN(n14940) );
  NAND2_X1 U12083 ( .A1(n15038), .A2(n9836), .ZN(n15023) );
  NAND2_X1 U12084 ( .A1(n14906), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14905) );
  AND2_X1 U12085 ( .A1(n14904), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14902) );
  AND2_X1 U12086 ( .A1(n14902), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14906) );
  AND2_X1 U12087 ( .A1(n12894), .A2(n10053), .ZN(n14901) );
  AND2_X1 U12088 ( .A1(n9783), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10053) );
  NAND2_X1 U12089 ( .A1(n12894), .A2(n9783), .ZN(n12895) );
  NAND2_X1 U12090 ( .A1(n12894), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12893) );
  AND2_X1 U12091 ( .A1(n11252), .A2(n11251), .ZN(n13648) );
  NAND2_X1 U12092 ( .A1(n13533), .A2(n10205), .ZN(n13647) );
  NOR2_X1 U12093 ( .A1(n16170), .A2(n12891), .ZN(n12894) );
  NAND2_X1 U12094 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n12892), .ZN(
        n12891) );
  AND2_X1 U12095 ( .A1(n13533), .A2(n13532), .ZN(n13535) );
  NOR2_X1 U12096 ( .A1(n21003), .A2(n12889), .ZN(n12892) );
  NAND2_X1 U12097 ( .A1(n10071), .A2(n10070), .ZN(n12889) );
  AND2_X1 U12098 ( .A1(n9785), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10070) );
  AND2_X1 U12099 ( .A1(n10071), .A2(n9785), .ZN(n12890) );
  NAND2_X1 U12100 ( .A1(n10071), .A2(n10072), .ZN(n12887) );
  NOR2_X1 U12101 ( .A1(n12885), .A2(n16205), .ZN(n12888) );
  NAND2_X1 U12102 ( .A1(n10193), .A2(n10194), .ZN(n13455) );
  INV_X1 U12103 ( .A(n10190), .ZN(n10194) );
  NOR2_X1 U12104 ( .A1(n12884), .A2(n13661), .ZN(n12886) );
  NAND2_X1 U12105 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12886), .ZN(
        n12885) );
  AND2_X1 U12106 ( .A1(n11271), .A2(n11270), .ZN(n13389) );
  NAND2_X1 U12107 ( .A1(n11651), .A2(n11714), .ZN(n10171) );
  OR2_X1 U12108 ( .A1(n14948), .A2(n14947), .ZN(n14950) );
  NOR2_X1 U12109 ( .A1(n9934), .A2(n15267), .ZN(n9933) );
  INV_X1 U12110 ( .A(n9935), .ZN(n9934) );
  NAND2_X1 U12111 ( .A1(n10210), .A2(n9873), .ZN(n10048) );
  NAND2_X1 U12112 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U12113 ( .A1(n14996), .A2(n9862), .ZN(n14051) );
  AND2_X1 U12114 ( .A1(n15336), .A2(n11401), .ZN(n15302) );
  NOR2_X1 U12115 ( .A1(n15142), .A2(n15301), .ZN(n15136) );
  NAND2_X1 U12116 ( .A1(n15327), .A2(n9935), .ZN(n15142) );
  NAND2_X1 U12117 ( .A1(n15327), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15329) );
  INV_X1 U12118 ( .A(n11151), .ZN(n15326) );
  AND2_X1 U12119 ( .A1(n14934), .A2(n10178), .ZN(n15093) );
  NAND2_X1 U12120 ( .A1(n9990), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15149) );
  NAND2_X1 U12121 ( .A1(n14934), .A2(n14921), .ZN(n15342) );
  AND2_X1 U12122 ( .A1(n15038), .A2(n9851), .ZN(n15003) );
  INV_X1 U12123 ( .A(n14925), .ZN(n10200) );
  NAND2_X1 U12124 ( .A1(n15038), .A2(n9837), .ZN(n14942) );
  AND2_X1 U12125 ( .A1(n9782), .A2(n11615), .ZN(n10181) );
  NAND2_X1 U12126 ( .A1(n16246), .A2(n9782), .ZN(n15389) );
  AND2_X1 U12127 ( .A1(n11303), .A2(n11302), .ZN(n15036) );
  NOR2_X1 U12128 ( .A1(n15037), .A2(n15036), .ZN(n15038) );
  NAND2_X1 U12129 ( .A1(n13764), .A2(n13763), .ZN(n15037) );
  AND2_X1 U12130 ( .A1(n16246), .A2(n10182), .ZN(n14018) );
  NAND2_X1 U12131 ( .A1(n16246), .A2(n12911), .ZN(n14016) );
  AND2_X1 U12132 ( .A1(n12913), .A2(n13638), .ZN(n13764) );
  NAND2_X1 U12133 ( .A1(n13533), .A2(n9773), .ZN(n13639) );
  AND2_X1 U12134 ( .A1(n15447), .A2(n10216), .ZN(n10215) );
  NAND2_X1 U12135 ( .A1(n9984), .A2(n9914), .ZN(n9913) );
  AND2_X1 U12136 ( .A1(n11067), .A2(n16152), .ZN(n16162) );
  NAND2_X1 U12137 ( .A1(n13161), .A2(n9771), .ZN(n15451) );
  NAND2_X1 U12138 ( .A1(n15246), .A2(n10147), .ZN(n9925) );
  INV_X1 U12139 ( .A(n10145), .ZN(n10144) );
  AND2_X1 U12140 ( .A1(n10192), .A2(n13448), .ZN(n10189) );
  NAND2_X1 U12141 ( .A1(n9985), .A2(n11039), .ZN(n16191) );
  NAND2_X1 U12142 ( .A1(n10209), .A2(n10738), .ZN(n11262) );
  NAND2_X1 U12143 ( .A1(n11678), .A2(n14045), .ZN(n9879) );
  INV_X1 U12144 ( .A(n10875), .ZN(n9878) );
  OAI22_X1 U12145 ( .A1(n10728), .A2(n10713), .B1(n11272), .B2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10133) );
  XNOR2_X1 U12146 ( .A(n13040), .B(n11416), .ZN(n13084) );
  AND2_X1 U12147 ( .A1(n11421), .A2(n11420), .ZN(n13083) );
  NAND2_X1 U12148 ( .A1(n10066), .A2(n10065), .ZN(n19052) );
  CLKBUF_X1 U12149 ( .A(n10787), .Z(n10788) );
  NOR2_X1 U12150 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10033) );
  NAND2_X1 U12151 ( .A1(n10142), .A2(n13224), .ZN(n13307) );
  INV_X1 U12152 ( .A(n10760), .ZN(n9903) );
  INV_X1 U12153 ( .A(n19368), .ZN(n19434) );
  INV_X1 U12154 ( .A(n19590), .ZN(n19593) );
  INV_X1 U12155 ( .A(n19567), .ZN(n13580) );
  INV_X1 U12156 ( .A(n19438), .ZN(n13552) );
  INV_X1 U12157 ( .A(n19235), .ZN(n19236) );
  INV_X1 U12158 ( .A(n19234), .ZN(n19238) );
  NAND2_X1 U12159 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19651), .ZN(n19240) );
  OR3_X1 U12160 ( .A1(n13539), .A2(n19727), .A3(n19872), .ZN(n13548) );
  NOR2_X2 U12161 ( .A1(n13812), .A2(n13551), .ZN(n19235) );
  NOR2_X2 U12162 ( .A1(n13550), .A2(n13551), .ZN(n19234) );
  NOR2_X1 U12163 ( .A1(n16547), .A2(n16546), .ZN(n16545) );
  NOR2_X1 U12164 ( .A1(n17504), .A2(n16560), .ZN(n16559) );
  NOR2_X1 U12165 ( .A1(n16603), .A2(n16602), .ZN(n16601) );
  NOR2_X1 U12166 ( .A1(n17584), .A2(n16622), .ZN(n16621) );
  NOR2_X1 U12167 ( .A1(n17718), .A2(n12710), .ZN(n16753) );
  AND2_X1 U12168 ( .A1(n9967), .A2(P3_EBX_REG_23__SCAN_IN), .ZN(n9966) );
  NAND2_X1 U12169 ( .A1(n16979), .A2(n9966), .ZN(n16945) );
  NOR2_X1 U12170 ( .A1(n16681), .A2(n9970), .ZN(n9969) );
  INV_X1 U12171 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n9970) );
  NOR2_X1 U12172 ( .A1(n17083), .A2(n17114), .ZN(n17080) );
  INV_X1 U12173 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17179) );
  INV_X1 U12174 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n20858) );
  OAI211_X1 U12175 ( .C1(n10275), .C2(n20841), .A(n10321), .B(n10320), .ZN(
        n10522) );
  NOR2_X1 U12176 ( .A1(n10311), .A2(n9946), .ZN(n9945) );
  NAND4_X1 U12177 ( .A1(n10552), .A2(n18227), .A3(n10544), .A4(n17392), .ZN(
        n17454) );
  NOR2_X1 U12178 ( .A1(n12714), .A2(n17848), .ZN(n16374) );
  INV_X1 U12179 ( .A(n16388), .ZN(n10087) );
  AND2_X1 U12180 ( .A1(n17608), .A2(n9850), .ZN(n17533) );
  INV_X1 U12181 ( .A(n17545), .ZN(n9991) );
  NOR2_X1 U12182 ( .A1(n17586), .A2(n9993), .ZN(n9992) );
  INV_X1 U12183 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U12184 ( .A1(n17608), .A2(n9784), .ZN(n17544) );
  NAND2_X1 U12185 ( .A1(n17608), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17585) );
  NOR2_X1 U12186 ( .A1(n17746), .A2(n9996), .ZN(n9995) );
  INV_X1 U12187 ( .A(n9998), .ZN(n9997) );
  INV_X1 U12188 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20927) );
  AOI21_X1 U12189 ( .B1(n12712), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n18241), .ZN(n17691) );
  INV_X1 U12190 ( .A(n18053), .ZN(n17726) );
  NAND2_X1 U12191 ( .A1(n17807), .A2(n9952), .ZN(n9956) );
  NOR2_X1 U12192 ( .A1(n9953), .A2(n17799), .ZN(n9952) );
  INV_X1 U12193 ( .A(n17799), .ZN(n9951) );
  AOI21_X1 U12194 ( .B1(n9953), .B2(n17799), .A(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9950) );
  NOR2_X1 U12195 ( .A1(n17797), .A2(n20943), .ZN(n17790) );
  AND2_X1 U12196 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17815) );
  NOR2_X1 U12197 ( .A1(n18654), .A2(n18713), .ZN(n12719) );
  INV_X1 U12198 ( .A(n17358), .ZN(n16391) );
  NOR2_X1 U12199 ( .A1(n10384), .A2(n10076), .ZN(n10075) );
  NAND2_X1 U12200 ( .A1(n10377), .A2(n10232), .ZN(n10378) );
  NAND2_X1 U12201 ( .A1(n10380), .A2(n17558), .ZN(n10377) );
  NOR2_X1 U12202 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n10376), .ZN(
        n17601) );
  INV_X1 U12203 ( .A(n10556), .ZN(n17974) );
  NAND2_X1 U12204 ( .A1(n10080), .A2(n10078), .ZN(n17662) );
  AND2_X1 U12205 ( .A1(n9792), .A2(n20895), .ZN(n10078) );
  NAND2_X1 U12206 ( .A1(n17764), .A2(n10373), .ZN(n17696) );
  OAI21_X1 U12207 ( .B1(n10552), .B2(n15534), .A(n10551), .ZN(n18660) );
  NOR2_X1 U12208 ( .A1(n10548), .A2(n10537), .ZN(n18661) );
  NAND2_X1 U12209 ( .A1(n18093), .A2(n17765), .ZN(n17764) );
  NOR2_X1 U12210 ( .A1(n17777), .A2(n17776), .ZN(n17775) );
  NAND2_X1 U12211 ( .A1(n17771), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17770) );
  NOR2_X1 U12212 ( .A1(n18855), .A2(n18088), .ZN(n18645) );
  AOI21_X1 U12213 ( .B1(n10542), .B2(n10541), .A(n16508), .ZN(n18656) );
  INV_X1 U12214 ( .A(n10497), .ZN(n10542) );
  NOR2_X1 U12215 ( .A1(n18855), .A2(n13907), .ZN(n10541) );
  AND2_X1 U12216 ( .A1(n10551), .A2(n10549), .ZN(n18657) );
  INV_X1 U12217 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18675) );
  NOR4_X2 U12218 ( .A1(n10470), .A2(n10468), .A3(n9975), .A4(n9974), .ZN(
        n18219) );
  INV_X1 U12219 ( .A(n10469), .ZN(n9974) );
  OAI21_X1 U12220 ( .B1(n12882), .B2(n12881), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13811) );
  INV_X1 U12221 ( .A(n15662), .ZN(n19985) );
  NAND2_X1 U12222 ( .A1(n13626), .A2(n13625), .ZN(n19946) );
  NAND2_X1 U12223 ( .A1(n13626), .A2(n13624), .ZN(n15662) );
  INV_X1 U12224 ( .A(n19975), .ZN(n19993) );
  INV_X1 U12225 ( .A(n19946), .ZN(n19994) );
  AND2_X1 U12226 ( .A1(n15751), .A2(n14473), .ZN(n19999) );
  INV_X1 U12227 ( .A(n14612), .ZN(n14617) );
  OAI211_X2 U12228 ( .C1(n12956), .C2(n12849), .A(n12848), .B(n12847), .ZN(
        n20015) );
  NAND2_X1 U12229 ( .A1(n14351), .A2(n12980), .ZN(n20051) );
  INV_X2 U12230 ( .A(n20044), .ZN(n20049) );
  XNOR2_X1 U12231 ( .A(n12830), .B(n14362), .ZN(n13616) );
  OAI21_X1 U12232 ( .B1(n14388), .B2(n14389), .A(n14376), .ZN(n14651) );
  AND2_X1 U12233 ( .A1(n15784), .A2(n12828), .ZN(n15820) );
  INV_X1 U12234 ( .A(n15784), .ZN(n20076) );
  INV_X1 U12235 ( .A(n20081), .ZN(n19900) );
  INV_X1 U12236 ( .A(n14666), .ZN(n20142) );
  XNOR2_X1 U12237 ( .A(n14356), .B(n14355), .ZN(n14756) );
  NAND2_X1 U12238 ( .A1(n14502), .A2(n9861), .ZN(n10029) );
  NAND2_X1 U12239 ( .A1(n13149), .A2(n14031), .ZN(n15893) );
  NAND2_X1 U12240 ( .A1(n15843), .A2(n12765), .ZN(n15840) );
  OR2_X1 U12241 ( .A1(n13443), .A2(n9804), .ZN(n15966) );
  OAI21_X1 U12242 ( .B1(n20079), .B2(n10116), .A(n10118), .ZN(n15845) );
  INV_X1 U12243 ( .A(n10117), .ZN(n10116) );
  NOR2_X1 U12244 ( .A1(n20111), .A2(n15915), .ZN(n20098) );
  NAND2_X1 U12245 ( .A1(n13163), .A2(n13162), .ZN(n13165) );
  XNOR2_X1 U12246 ( .A(n10019), .B(n13097), .ZN(n13163) );
  INV_X1 U12247 ( .A(n20109), .ZN(n20126) );
  INV_X1 U12248 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20488) );
  INV_X1 U12249 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12975) );
  OR2_X1 U12250 ( .A1(n20651), .A2(n20369), .ZN(n20656) );
  INV_X1 U12251 ( .A(n20267), .ZN(n20284) );
  NOR2_X2 U12252 ( .A1(n20493), .A2(n20455), .ZN(n20512) );
  OAI211_X1 U12253 ( .C1(n20634), .C2(n20606), .A(n20605), .B(n20604), .ZN(
        n20638) );
  INV_X1 U12254 ( .A(n20525), .ZN(n20645) );
  INV_X1 U12255 ( .A(n20536), .ZN(n20646) );
  INV_X1 U12256 ( .A(n20541), .ZN(n20662) );
  INV_X1 U12257 ( .A(n20546), .ZN(n20668) );
  AND2_X1 U12258 ( .A1(n20165), .A2(n20187), .ZN(n20673) );
  INV_X1 U12259 ( .A(n20551), .ZN(n20674) );
  INV_X1 U12260 ( .A(n20552), .ZN(n20679) );
  INV_X1 U12261 ( .A(n20556), .ZN(n20680) );
  INV_X1 U12262 ( .A(n20561), .ZN(n20686) );
  AND2_X1 U12263 ( .A1(n20181), .A2(n20187), .ZN(n20691) );
  INV_X1 U12264 ( .A(n21074), .ZN(n20692) );
  INV_X1 U12265 ( .A(n20656), .ZN(n20701) );
  INV_X1 U12266 ( .A(n20567), .ZN(n20698) );
  NOR2_X1 U12267 ( .A1(n14342), .A2(n20532), .ZN(n15602) );
  AND2_X1 U12268 ( .A1(n13156), .A2(n19049), .ZN(n19875) );
  INV_X1 U12269 ( .A(n19067), .ZN(n19041) );
  INV_X1 U12270 ( .A(n19741), .ZN(n19036) );
  INV_X1 U12271 ( .A(n19047), .ZN(n19070) );
  OR2_X1 U12272 ( .A1(n11585), .A2(n11584), .ZN(n13636) );
  OR2_X1 U12273 ( .A1(n11526), .A2(n11525), .ZN(n13652) );
  OR2_X1 U12274 ( .A1(n11505), .A2(n11504), .ZN(n13530) );
  INV_X1 U12275 ( .A(n15026), .ZN(n15007) );
  INV_X1 U12276 ( .A(n19848), .ZN(n19281) );
  INV_X2 U12277 ( .A(n14992), .ZN(n15040) );
  NOR2_X1 U12278 ( .A1(n14964), .A2(n14963), .ZN(n14962) );
  NAND2_X1 U12279 ( .A1(n10141), .A2(n14957), .ZN(n14964) );
  NOR2_X1 U12280 ( .A1(n14997), .A2(n14163), .ZN(n14987) );
  AND2_X1 U12281 ( .A1(n13813), .A2(n13811), .ZN(n19084) );
  AND2_X1 U12282 ( .A1(n13813), .A2(n13812), .ZN(n19083) );
  AND2_X1 U12283 ( .A1(n19103), .A2(n13815), .ZN(n19082) );
  AND2_X1 U12284 ( .A1(n19107), .A2(n16092), .ZN(n19113) );
  NAND2_X1 U12285 ( .A1(n13380), .A2(n13379), .ZN(n13387) );
  NOR2_X1 U12286 ( .A1(n13220), .A2(n13018), .ZN(n19248) );
  INV_X1 U12287 ( .A(n16092), .ZN(n19087) );
  INV_X1 U12288 ( .A(n19103), .ZN(n19104) );
  AOI21_X1 U12289 ( .B1(n12936), .B2(n13294), .A(n19881), .ZN(n19148) );
  NAND2_X1 U12290 ( .A1(n16108), .A2(n16107), .ZN(n16106) );
  NAND2_X1 U12291 ( .A1(n10214), .A2(n15159), .ZN(n16108) );
  INV_X1 U12292 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21003) );
  INV_X1 U12293 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16205) );
  INV_X1 U12294 ( .A(n16198), .ZN(n19167) );
  NAND2_X1 U12295 ( .A1(n12928), .A2(n11709), .ZN(n16204) );
  AND2_X1 U12296 ( .A1(n16204), .A2(n19168), .ZN(n16198) );
  XNOR2_X1 U12297 ( .A(n15111), .B(n15110), .ZN(n15263) );
  XNOR2_X1 U12298 ( .A(n14950), .B(n14331), .ZN(n15999) );
  XNOR2_X1 U12299 ( .A(n9911), .B(n14049), .ZN(n15285) );
  OR2_X1 U12300 ( .A1(n15353), .A2(n15181), .ZN(n16224) );
  NAND2_X1 U12301 ( .A1(n19196), .A2(n14013), .ZN(n10165) );
  INV_X1 U12302 ( .A(n10164), .ZN(n10163) );
  AOI21_X1 U12303 ( .B1(n15237), .B2(n14014), .A(n16240), .ZN(n10164) );
  NAND2_X1 U12304 ( .A1(n11046), .A2(n11045), .ZN(n15459) );
  NOR3_X1 U12305 ( .A1(n11696), .A2(n16285), .A3(n16272), .ZN(n15471) );
  NAND2_X1 U12306 ( .A1(n10149), .A2(n15242), .ZN(n16184) );
  NAND2_X1 U12307 ( .A1(n10151), .A2(n10150), .ZN(n10149) );
  OR2_X1 U12308 ( .A1(n16309), .A2(n11654), .ZN(n16298) );
  AND2_X1 U12309 ( .A1(n14013), .A2(n13992), .ZN(n16309) );
  AND2_X1 U12310 ( .A1(n11704), .A2(n11650), .ZN(n19186) );
  INV_X1 U12311 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19861) );
  INV_X1 U12312 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19845) );
  INV_X1 U12313 ( .A(n19256), .ZN(n19273) );
  OAI21_X1 U12314 ( .B1(n19347), .B2(n19346), .A(n19345), .ZN(n19365) );
  AND2_X1 U12315 ( .A1(n19408), .A2(n19407), .ZN(n19415) );
  NOR2_X1 U12316 ( .A1(n19434), .A2(n19370), .ZN(n19412) );
  INV_X1 U12317 ( .A(n19415), .ZN(n19430) );
  NOR2_X2 U12318 ( .A1(n19400), .A2(n19438), .ZN(n19459) );
  INV_X1 U12319 ( .A(n19443), .ZN(n19460) );
  INV_X1 U12320 ( .A(n19516), .ZN(n19522) );
  OAI21_X1 U12321 ( .B1(n19535), .B2(n19550), .A(n19651), .ZN(n19553) );
  INV_X1 U12322 ( .A(n19667), .ZN(n19602) );
  OAI22_X1 U12323 ( .A1(n19223), .A2(n19238), .B1(n19222), .B2(n19236), .ZN(
        n19610) );
  INV_X1 U12324 ( .A(n19643), .ZN(n19630) );
  INV_X1 U12325 ( .A(n19699), .ZN(n19668) );
  OAI21_X1 U12326 ( .B1(n19657), .B2(n19656), .A(n19655), .ZN(n19687) );
  INV_X1 U12327 ( .A(n19730), .ZN(n19692) );
  INV_X1 U12328 ( .A(n19661), .ZN(n19598) );
  AND2_X1 U12329 ( .A1(n10757), .A2(n13586), .ZN(n19662) );
  INV_X1 U12330 ( .A(n19675), .ZN(n19702) );
  NAND2_X1 U12331 ( .A1(n19527), .A2(n13552), .ZN(n19724) );
  INV_X1 U12332 ( .A(n19735), .ZN(n19721) );
  INV_X1 U12333 ( .A(n19724), .ZN(n19731) );
  AND2_X1 U12334 ( .A1(n16346), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19737) );
  NOR3_X1 U12335 ( .A1(n16351), .A2(n19873), .A3(n16350), .ZN(n19743) );
  INV_X1 U12336 ( .A(n18873), .ZN(n18872) );
  NAND2_X1 U12337 ( .A1(n17454), .A2(n10539), .ZN(n16492) );
  NAND2_X1 U12338 ( .A1(n18862), .A2(n18649), .ZN(n17455) );
  NOR2_X1 U12339 ( .A1(n18648), .A2(n17455), .ZN(n18873) );
  INV_X1 U12340 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18859) );
  INV_X1 U12341 ( .A(n12719), .ZN(n16493) );
  NOR2_X1 U12342 ( .A1(n17537), .A2(n16580), .ZN(n16579) );
  NOR2_X1 U12343 ( .A1(n17612), .A2(n16638), .ZN(n16637) );
  NAND2_X1 U12344 ( .A1(n16525), .A2(n9847), .ZN(n16667) );
  NOR2_X1 U12345 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16727), .ZN(n16709) );
  NAND2_X1 U12346 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16884), .ZN(n16870) );
  INV_X1 U12347 ( .A(n16884), .ZN(n16868) );
  INV_X1 U12348 ( .A(n16881), .ZN(n16880) );
  NAND4_X1 U12349 ( .A1(n18179), .A2(n18872), .A3(n18721), .A4(n18711), .ZN(
        n16884) );
  AND2_X1 U12350 ( .A1(n9966), .A2(n9965), .ZN(n9964) );
  NOR2_X1 U12351 ( .A1(n16940), .A2(n16888), .ZN(n9965) );
  NOR2_X1 U12352 ( .A1(n13911), .A2(n16981), .ZN(n9967) );
  AND2_X1 U12353 ( .A1(n17066), .A2(n9968), .ZN(n17010) );
  AND2_X1 U12354 ( .A1(n9793), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n9968) );
  NAND2_X1 U12355 ( .A1(n17066), .A2(n9793), .ZN(n16997) );
  NAND2_X1 U12356 ( .A1(n17066), .A2(P3_EBX_REG_16__SCAN_IN), .ZN(n17049) );
  NOR2_X1 U12357 ( .A1(n21047), .A2(n17051), .ZN(n17066) );
  NAND2_X1 U12358 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17135), .ZN(n17114) );
  NOR2_X1 U12359 ( .A1(n17204), .A2(n17081), .ZN(n17135) );
  NAND2_X1 U12360 ( .A1(n17211), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n17204) );
  NAND2_X1 U12361 ( .A1(n17230), .A2(n9972), .ZN(n17208) );
  AND2_X1 U12362 ( .A1(n17205), .A2(P3_EBX_REG_4__SCAN_IN), .ZN(n9972) );
  NOR2_X1 U12363 ( .A1(n17208), .A2(n16822), .ZN(n17211) );
  NOR2_X1 U12364 ( .A1(n15641), .A2(n9973), .ZN(n17230) );
  OR3_X1 U12365 ( .A1(n18204), .A2(n18210), .A3(n18713), .ZN(n9973) );
  NOR2_X1 U12366 ( .A1(n17397), .A2(n17257), .ZN(n17250) );
  NAND2_X1 U12367 ( .A1(n17261), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n17257) );
  NOR2_X1 U12368 ( .A1(n17266), .A2(n17400), .ZN(n17261) );
  NOR2_X1 U12369 ( .A1(n17270), .A2(n17404), .ZN(n17271) );
  NAND2_X1 U12370 ( .A1(n17271), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17266) );
  NOR2_X1 U12371 ( .A1(n17406), .A2(n17278), .ZN(n17277) );
  INV_X1 U12372 ( .A(n17294), .ZN(n17290) );
  INV_X1 U12373 ( .A(n17304), .ZN(n17309) );
  NOR2_X1 U12374 ( .A1(n17321), .A2(n17420), .ZN(n17316) );
  INV_X1 U12375 ( .A(n17283), .ZN(n17314) );
  NOR2_X1 U12376 ( .A1(n17354), .A2(n9867), .ZN(n17330) );
  NAND2_X1 U12377 ( .A1(n17233), .A2(n17325), .ZN(n17354) );
  AND2_X1 U12378 ( .A1(n17325), .A2(n17386), .ZN(n17360) );
  OAI211_X1 U12379 ( .C1(n10464), .C2(n17068), .A(n10331), .B(n10330), .ZN(
        n17362) );
  NOR2_X1 U12380 ( .A1(n10280), .A2(n10279), .ZN(n10281) );
  INV_X1 U12381 ( .A(n10508), .ZN(n17379) );
  NAND2_X1 U12382 ( .A1(n17353), .A2(n18669), .ZN(n17382) );
  INV_X1 U12383 ( .A(n17353), .ZN(n17378) );
  INV_X1 U12384 ( .A(n10348), .ZN(n10350) );
  OAI21_X1 U12385 ( .B1(n15643), .B2(n15642), .A(n18862), .ZN(n17383) );
  NAND2_X1 U12386 ( .A1(n15644), .A2(n17233), .ZN(n17389) );
  INV_X1 U12387 ( .A(n17383), .ZN(n17233) );
  INV_X1 U12388 ( .A(n17389), .ZN(n17344) );
  INV_X1 U12389 ( .A(n17382), .ZN(n17384) );
  INV_X1 U12390 ( .A(n17444), .ZN(n17426) );
  NOR2_X1 U12391 ( .A1(n17455), .A2(n17390), .ZN(n17447) );
  OR2_X1 U12392 ( .A1(n17455), .A2(n18705), .ZN(n17500) );
  INV_X1 U12393 ( .A(n17495), .ZN(n17498) );
  NOR2_X1 U12394 ( .A1(n9719), .A2(n17726), .ZN(n18093) );
  NAND2_X1 U12395 ( .A1(n17815), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17797) );
  INV_X1 U12396 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20943) );
  INV_X1 U12397 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17826) );
  INV_X1 U12398 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17841) );
  NAND2_X1 U12399 ( .A1(n17855), .A2(n17822), .ZN(n17850) );
  OAI21_X1 U12400 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18861), .A(n16493), 
        .ZN(n17855) );
  NAND2_X1 U12401 ( .A1(n10076), .A2(n17876), .ZN(n9958) );
  INV_X1 U12402 ( .A(n18094), .ZN(n18023) );
  AND2_X1 U12403 ( .A1(n9949), .A2(n10374), .ZN(n17646) );
  NOR2_X1 U12404 ( .A1(n18658), .A2(n18673), .ZN(n18068) );
  NAND2_X1 U12405 ( .A1(n10080), .A2(n10081), .ZN(n17716) );
  INV_X1 U12406 ( .A(n18099), .ZN(n18072) );
  NOR2_X1 U12407 ( .A1(n17743), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17729) );
  AOI21_X2 U12408 ( .B1(n18661), .B2(n18656), .A(n18660), .ZN(n18670) );
  NAND2_X1 U12409 ( .A1(n17800), .A2(n17799), .ZN(n17798) );
  NAND2_X1 U12410 ( .A1(n17807), .A2(n10361), .ZN(n17800) );
  NOR2_X2 U12411 ( .A1(n18871), .A2(n13908), .ZN(n18658) );
  AOI21_X2 U12412 ( .B1(n10507), .B2(n10506), .A(n18713), .ZN(n18163) );
  NOR2_X1 U12413 ( .A1(n9732), .A2(n18163), .ZN(n18164) );
  NAND2_X1 U12414 ( .A1(n18656), .A2(n15535), .ZN(n18673) );
  INV_X1 U12415 ( .A(n18657), .ZN(n15535) );
  INV_X1 U12416 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18674) );
  INV_X1 U12417 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18197) );
  NOR2_X1 U12418 ( .A1(n18203), .A2(n15540), .ZN(n18841) );
  INV_X1 U12419 ( .A(n18841), .ZN(n18839) );
  INV_X1 U12420 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20831) );
  INV_X1 U12421 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18222) );
  INV_X1 U12422 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n21001) );
  INV_X1 U12423 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18810) );
  OAI21_X1 U12425 ( .B1(n14814), .B2(n15913), .A(n10009), .ZN(P1_U3004) );
  NOR2_X1 U12426 ( .A1(n14815), .A2(n10010), .ZN(n10009) );
  AND2_X1 U12427 ( .A1(n14817), .A2(n14816), .ZN(n10010) );
  NOR2_X1 U12428 ( .A1(n10199), .A2(n10196), .ZN(n11718) );
  NOR2_X1 U12429 ( .A1(n11715), .A2(n16158), .ZN(n10199) );
  NAND2_X1 U12430 ( .A1(n11705), .A2(n9930), .ZN(P2_U3015) );
  INV_X1 U12431 ( .A(n9931), .ZN(n9930) );
  NAND2_X1 U12432 ( .A1(n16979), .A2(P3_EBX_REG_21__SCAN_IN), .ZN(n16966) );
  NAND2_X1 U12433 ( .A1(n10088), .A2(n10083), .ZN(P3_U2801) );
  NOR2_X1 U12434 ( .A1(n16384), .A2(n10084), .ZN(n10083) );
  OR2_X1 U12435 ( .A1(n16383), .A2(n17741), .ZN(n10088) );
  INV_X1 U12436 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13326) );
  CLKBUF_X3 U12437 ( .A(n10395), .Z(n17139) );
  OR3_X2 U12438 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n10246), .ZN(n9796) );
  AND2_X1 U12439 ( .A1(n14048), .A2(n10211), .ZN(n9767) );
  NAND2_X2 U12440 ( .A1(n10645), .A2(n10644), .ZN(n10689) );
  AND2_X1 U12441 ( .A1(n11035), .A2(n10986), .ZN(n9768) );
  NAND2_X1 U12442 ( .A1(n14547), .A2(n9832), .ZN(n14426) );
  AND2_X1 U12443 ( .A1(n17692), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9769) );
  AND2_X1 U12444 ( .A1(n15802), .A2(n14711), .ZN(n9770) );
  AND2_X1 U12445 ( .A1(n14413), .A2(n9841), .ZN(n14388) );
  AND2_X1 U12446 ( .A1(n10172), .A2(n13317), .ZN(n9771) );
  INV_X1 U12447 ( .A(n15243), .ZN(n10150) );
  AND2_X1 U12448 ( .A1(n11695), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15243) );
  AND2_X1 U12449 ( .A1(n12817), .A2(n9962), .ZN(n9772) );
  AND2_X1 U12450 ( .A1(n10203), .A2(n13559), .ZN(n9773) );
  AND4_X1 U12451 ( .A1(n11781), .A2(n11780), .A3(n11779), .A4(n11778), .ZN(
        n9774) );
  AND2_X1 U12452 ( .A1(n11924), .A2(n11993), .ZN(n9775) );
  NOR2_X1 U12453 ( .A1(n10067), .A2(n10068), .ZN(n9776) );
  AND4_X1 U12454 ( .A1(n10870), .A2(n10869), .A3(n10868), .A4(n10867), .ZN(
        n9777) );
  AND2_X1 U12455 ( .A1(n9768), .A2(n10052), .ZN(n9778) );
  AND2_X1 U12456 ( .A1(n9797), .A2(n12591), .ZN(n9779) );
  NAND2_X1 U12457 ( .A1(n10688), .A2(n19871), .ZN(n11619) );
  NAND2_X1 U12458 ( .A1(n10153), .A2(n13383), .ZN(n13447) );
  OR2_X1 U12459 ( .A1(n13644), .A2(n10125), .ZN(n9780) );
  AND2_X1 U12460 ( .A1(n9835), .A2(n10032), .ZN(n9781) );
  AND2_X1 U12461 ( .A1(n10182), .A2(n13808), .ZN(n9782) );
  AND2_X1 U12462 ( .A1(n10054), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9783) );
  AND2_X1 U12463 ( .A1(n9992), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9784) );
  AND2_X1 U12464 ( .A1(n10072), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9785) );
  INV_X1 U12465 ( .A(n10159), .ZN(n15010) );
  AND2_X1 U12466 ( .A1(n13863), .A2(n13889), .ZN(n9786) );
  AND2_X1 U12467 ( .A1(n10021), .A2(n10020), .ZN(n9787) );
  AND2_X1 U12468 ( .A1(n9781), .A2(n9863), .ZN(n9788) );
  INV_X1 U12469 ( .A(n10795), .ZN(n14165) );
  OR2_X1 U12470 ( .A1(n15055), .A2(n15046), .ZN(n9789) );
  AND2_X1 U12471 ( .A1(n10061), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9790) );
  AND2_X1 U12472 ( .A1(n10058), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9791) );
  INV_X1 U12473 ( .A(n14963), .ZN(n10140) );
  AND2_X1 U12474 ( .A1(n10081), .A2(n10079), .ZN(n9792) );
  AND2_X1 U12475 ( .A1(n9969), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n9793) );
  OR2_X1 U12476 ( .A1(n10246), .A2(n10247), .ZN(n9794) );
  INV_X1 U12477 ( .A(n11820), .ZN(n11819) );
  NAND2_X1 U12478 ( .A1(n11723), .A2(n11728), .ZN(n11820) );
  INV_X2 U12479 ( .A(n11820), .ZN(n12243) );
  AND4_X1 U12480 ( .A1(n18819), .A2(n18826), .A3(n18834), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9795) );
  INV_X1 U12481 ( .A(n10742), .ZN(n11248) );
  OR2_X1 U12482 ( .A1(n14348), .A2(n12606), .ZN(n9797) );
  OR3_X1 U12483 ( .A1(n18826), .A2(n18819), .A3(n18685), .ZN(n9798) );
  AND2_X1 U12484 ( .A1(n14547), .A2(n10127), .ZN(n14425) );
  INV_X1 U12485 ( .A(n10168), .ZN(n16122) );
  INV_X1 U12486 ( .A(n11272), .ZN(n11341) );
  AND2_X1 U12487 ( .A1(n10705), .A2(n9881), .ZN(n11272) );
  INV_X1 U12488 ( .A(n9918), .ZN(n9920) );
  INV_X1 U12489 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14035) );
  AND2_X1 U12490 ( .A1(n11033), .A2(n10982), .ZN(n9799) );
  AND4_X1 U12491 ( .A1(n11739), .A2(n11738), .A3(n11737), .A4(n11736), .ZN(
        n9801) );
  AND4_X1 U12492 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n9802) );
  INV_X1 U12494 ( .A(n14048), .ZN(n10210) );
  AND2_X1 U12495 ( .A1(n13078), .A2(n13021), .ZN(n10763) );
  OAI21_X1 U12496 ( .B1(n15415), .B2(n9922), .A(n9920), .ZN(n15160) );
  AND2_X1 U12497 ( .A1(n12626), .A2(n12625), .ZN(n9804) );
  INV_X1 U12498 ( .A(n9895), .ZN(n12051) );
  INV_X1 U12499 ( .A(n20176), .ZN(n11849) );
  NAND2_X1 U12500 ( .A1(n15076), .A2(n10175), .ZN(n9805) );
  AND3_X1 U12501 ( .A1(n10767), .A2(n10766), .A3(n10782), .ZN(n9806) );
  OR2_X1 U12502 ( .A1(n17454), .A2(n18210), .ZN(n9807) );
  AND2_X1 U12503 ( .A1(n10689), .A2(n10688), .ZN(n9808) );
  AND2_X1 U12504 ( .A1(n15793), .A2(n10113), .ZN(n10112) );
  OAI21_X1 U12505 ( .B1(n14705), .B2(n10006), .A(n10112), .ZN(n14702) );
  NOR2_X1 U12506 ( .A1(n14987), .A2(n14986), .ZN(n9809) );
  NOR2_X1 U12507 ( .A1(n11122), .A2(n15202), .ZN(n9810) );
  AND2_X1 U12508 ( .A1(n9778), .A2(n11034), .ZN(n9811) );
  OR2_X1 U12509 ( .A1(n10275), .A2(n17158), .ZN(n9812) );
  AND4_X1 U12510 ( .A1(n10427), .A2(n9943), .A3(n10428), .A4(n9938), .ZN(n9813) );
  AND2_X1 U12511 ( .A1(n10378), .A2(n17904), .ZN(n9814) );
  OR2_X1 U12512 ( .A1(n9776), .A2(n10063), .ZN(n9815) );
  INV_X1 U12513 ( .A(n10039), .ZN(n11672) );
  OR2_X1 U12514 ( .A1(n10042), .A2(n10871), .ZN(n10039) );
  INV_X1 U12515 ( .A(n12802), .ZN(n10114) );
  INV_X1 U12516 ( .A(n10147), .ZN(n10146) );
  AND2_X1 U12517 ( .A1(n15242), .A2(n10148), .ZN(n10147) );
  INV_X1 U12518 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n20881) );
  AND2_X1 U12519 ( .A1(n10169), .A2(n9932), .ZN(n9816) );
  AND2_X1 U12520 ( .A1(n9912), .A2(n14047), .ZN(n9817) );
  INV_X1 U12521 ( .A(n10833), .ZN(n14105) );
  AND2_X1 U12522 ( .A1(n11700), .A2(n11699), .ZN(n9818) );
  NAND2_X1 U12523 ( .A1(n11870), .A2(n20155), .ZN(n9819) );
  INV_X1 U12524 ( .A(n10166), .ZN(n15235) );
  NAND2_X1 U12525 ( .A1(n10168), .A2(n10167), .ZN(n10166) );
  INV_X2 U12526 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18834) );
  AND2_X1 U12527 ( .A1(n11852), .A2(n11871), .ZN(n9820) );
  AND2_X1 U12528 ( .A1(n14413), .A2(n14510), .ZN(n14497) );
  OR2_X1 U12529 ( .A1(n14235), .A2(n14234), .ZN(n10228) );
  INV_X1 U12530 ( .A(n10228), .ZN(n10134) );
  AND2_X1 U12531 ( .A1(n10862), .A2(n10859), .ZN(n9821) );
  AND2_X1 U12532 ( .A1(n11776), .A2(n11777), .ZN(n9822) );
  AND2_X1 U12533 ( .A1(n20160), .A2(n12551), .ZN(n9823) );
  NAND2_X1 U12534 ( .A1(n9803), .A2(n10239), .ZN(n11841) );
  AND2_X1 U12535 ( .A1(n11840), .A2(n13137), .ZN(n9824) );
  AND2_X1 U12536 ( .A1(n9770), .A2(n12802), .ZN(n9825) );
  INV_X1 U12537 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10614) );
  INV_X1 U12538 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U12539 ( .A1(n15760), .A2(n15759), .ZN(n9826) );
  NAND2_X1 U12540 ( .A1(n11383), .A2(n10705), .ZN(n9827) );
  NAND2_X1 U12541 ( .A1(n13380), .A2(n10154), .ZN(n10153) );
  INV_X1 U12542 ( .A(n12885), .ZN(n10071) );
  NAND2_X1 U12543 ( .A1(n13017), .A2(n10688), .ZN(n13071) );
  AND2_X1 U12544 ( .A1(n16979), .A2(n9964), .ZN(n9828) );
  AND2_X1 U12545 ( .A1(n17066), .A2(n9969), .ZN(n9829) );
  NAND2_X1 U12546 ( .A1(n15038), .A2(n15032), .ZN(n15020) );
  AND2_X1 U12547 ( .A1(n14934), .A2(n10179), .ZN(n9830) );
  AND2_X1 U12548 ( .A1(n14906), .A2(n10058), .ZN(n9831) );
  AND2_X1 U12549 ( .A1(n10127), .A2(n10233), .ZN(n9832) );
  AND2_X1 U12550 ( .A1(n10080), .A2(n9792), .ZN(n9833) );
  AND2_X1 U12551 ( .A1(n12894), .A2(n10054), .ZN(n9834) );
  INV_X1 U12552 ( .A(n14045), .ZN(n11694) );
  AND2_X1 U12553 ( .A1(n12676), .A2(n14526), .ZN(n9835) );
  AND2_X1 U12554 ( .A1(n10202), .A2(n15032), .ZN(n9836) );
  AND2_X1 U12555 ( .A1(n9836), .A2(n10201), .ZN(n9837) );
  NAND2_X1 U12556 ( .A1(n12114), .A2(n12115), .ZN(n13502) );
  INV_X1 U12557 ( .A(n14257), .ZN(n10757) );
  AND2_X1 U12558 ( .A1(n13558), .A2(n13557), .ZN(n13635) );
  OAI21_X1 U12559 ( .B1(n15843), .B2(n10095), .A(n10092), .ZN(n15831) );
  INV_X1 U12560 ( .A(n11041), .ZN(n10052) );
  NAND2_X1 U12561 ( .A1(n10120), .A2(n12793), .ZN(n13766) );
  AND2_X1 U12562 ( .A1(n13635), .A2(n13634), .ZN(n9838) );
  AND2_X1 U12563 ( .A1(n15760), .A2(n9787), .ZN(n9839) );
  NOR3_X1 U12564 ( .A1(n12791), .A2(n12790), .A3(n20803), .ZN(n9840) );
  INV_X1 U12565 ( .A(n20181), .ZN(n11978) );
  NAND2_X1 U12566 ( .A1(n17645), .A2(n17679), .ZN(n17570) );
  AND2_X1 U12567 ( .A1(n10132), .A2(n10131), .ZN(n9841) );
  AND2_X1 U12568 ( .A1(n16979), .A2(n9967), .ZN(n9842) );
  AND2_X1 U12569 ( .A1(n12050), .A2(n12083), .ZN(n9843) );
  NAND2_X1 U12570 ( .A1(n9755), .A2(n11068), .ZN(n9844) );
  AND2_X1 U12571 ( .A1(n10160), .A2(n15012), .ZN(n9845) );
  OR2_X1 U12572 ( .A1(n12165), .A2(n12177), .ZN(n9846) );
  OR2_X1 U12573 ( .A1(n16674), .A2(n9996), .ZN(n9847) );
  INV_X1 U12574 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15248) );
  NAND2_X1 U12575 ( .A1(n13635), .A2(n10160), .ZN(n10159) );
  AND2_X1 U12576 ( .A1(n20176), .A2(n20155), .ZN(n12786) );
  INV_X1 U12577 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20708) );
  AND2_X1 U12578 ( .A1(n14541), .A2(n12676), .ZN(n14525) );
  AND2_X1 U12579 ( .A1(n16186), .A2(n16188), .ZN(n9848) );
  NAND3_X1 U12580 ( .A1(n16159), .A2(n15416), .A3(n16161), .ZN(n9849) );
  AND2_X1 U12581 ( .A1(n9784), .A2(n9991), .ZN(n9850) );
  AND2_X1 U12582 ( .A1(n9837), .A2(n10200), .ZN(n9851) );
  AND2_X1 U12583 ( .A1(n10152), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9852) );
  AND2_X1 U12584 ( .A1(n10126), .A2(n9832), .ZN(n9853) );
  AND2_X1 U12585 ( .A1(n12130), .A2(n10129), .ZN(n9854) );
  AND2_X1 U12586 ( .A1(n9787), .A2(n14558), .ZN(n9855) );
  NAND2_X1 U12587 ( .A1(n14188), .A2(n14187), .ZN(n9856) );
  NAND2_X1 U12588 ( .A1(n11447), .A2(n11446), .ZN(n13161) );
  INV_X1 U12589 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9996) );
  AND2_X1 U12590 ( .A1(n10153), .A2(n10152), .ZN(n13485) );
  AND2_X1 U12591 ( .A1(n10781), .A2(n10763), .ZN(n19528) );
  AND2_X1 U12592 ( .A1(n17608), .A2(n9992), .ZN(n9857) );
  OR2_X1 U12593 ( .A1(n13390), .A2(n13389), .ZN(n9858) );
  NAND2_X1 U12594 ( .A1(n13334), .A2(n12004), .ZN(n13403) );
  OR2_X1 U12595 ( .A1(n14909), .A2(n10207), .ZN(n9859) );
  OR2_X1 U12596 ( .A1(n17635), .A2(n16654), .ZN(n9860) );
  AND2_X1 U12597 ( .A1(n14401), .A2(n10027), .ZN(n9861) );
  OR2_X1 U12598 ( .A1(n12896), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10066) );
  OR3_X1 U12599 ( .A1(n9859), .A2(n10208), .A3(n14967), .ZN(n9862) );
  AND2_X1 U12600 ( .A1(n14505), .A2(n14506), .ZN(n9863) );
  NAND2_X1 U12601 ( .A1(n9895), .A2(n12026), .ZN(n20137) );
  NAND2_X1 U12602 ( .A1(n10193), .A2(n10192), .ZN(n10195) );
  AND2_X1 U12603 ( .A1(n10038), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n9864) );
  AND2_X1 U12604 ( .A1(n13161), .A2(n13160), .ZN(n9865) );
  NAND2_X1 U12605 ( .A1(n13533), .A2(n10203), .ZN(n10206) );
  NAND2_X1 U12606 ( .A1(n13161), .A2(n10172), .ZN(n10174) );
  AND2_X1 U12607 ( .A1(n10178), .A2(n14911), .ZN(n9866) );
  INV_X1 U12608 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9994) );
  INV_X1 U12609 ( .A(n14325), .ZN(n10177) );
  INV_X1 U12610 ( .A(n13881), .ZN(n10124) );
  NAND2_X1 U12611 ( .A1(n12962), .A2(n11814), .ZN(n14348) );
  INV_X1 U12612 ( .A(n14348), .ZN(n11839) );
  INV_X1 U12613 ( .A(n15184), .ZN(n10064) );
  OR2_X1 U12614 ( .A1(n17326), .A2(n17423), .ZN(n9867) );
  AND2_X1 U12615 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9868) );
  INV_X1 U12616 ( .A(n10068), .ZN(n10065) );
  NOR2_X1 U12617 ( .A1(n19884), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10068) );
  INV_X1 U12618 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10056) );
  OR2_X1 U12619 ( .A1(n17746), .A2(n16647), .ZN(n9869) );
  INV_X1 U12620 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9963) );
  AND2_X1 U12621 ( .A1(n10038), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n9870) );
  NAND2_X1 U12622 ( .A1(n17790), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17746) );
  OR2_X1 U12623 ( .A1(n12805), .A2(n12804), .ZN(n9871) );
  INV_X1 U12624 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10076) );
  OR2_X1 U12625 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9872) );
  INV_X1 U12626 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10069) );
  INV_X1 U12627 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n9971) );
  INV_X1 U12628 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10082) );
  OR2_X1 U12629 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9873) );
  OR2_X1 U12630 ( .A1(n19251), .A2(n19857), .ZN(n19567) );
  NOR2_X1 U12631 ( .A1(n19251), .A2(n19248), .ZN(n19527) );
  NOR3_X2 U12632 ( .A1(n18548), .A2(n18498), .A3(n18471), .ZN(n18465) );
  OAI21_X1 U12633 ( .B1(n15174), .B2(n15173), .A(n15172), .ZN(n15224) );
  OAI21_X1 U12634 ( .B1(n19409), .B2(n11511), .A(n9875), .ZN(n10754) );
  NAND2_X1 U12635 ( .A1(n19338), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n9875) );
  NAND2_X1 U12636 ( .A1(n19338), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n9876) );
  NAND2_X1 U12637 ( .A1(n19338), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n9877) );
  OAI21_X2 U12638 ( .B1(n9879), .B2(n9878), .A(n13666), .ZN(n13600) );
  NAND2_X1 U12639 ( .A1(n10875), .A2(n11678), .ZN(n13599) );
  NOR2_X2 U12640 ( .A1(n11374), .A2(n10711), .ZN(n11383) );
  NOR2_X1 U12641 ( .A1(n11374), .A2(n9882), .ZN(n9881) );
  AND2_X2 U12642 ( .A1(n16133), .A2(n16131), .ZN(n16117) );
  NAND2_X2 U12643 ( .A1(n11059), .A2(n11058), .ZN(n15415) );
  OAI21_X1 U12644 ( .B1(n14783), .B2(n9885), .A(n14626), .ZN(n14779) );
  NAND2_X1 U12646 ( .A1(n9824), .A2(n9779), .ZN(n11856) );
  NAND2_X1 U12647 ( .A1(n9889), .A2(n9888), .ZN(n9891) );
  NOR2_X1 U12648 ( .A1(n11847), .A2(n12589), .ZN(n9890) );
  OR2_X2 U12649 ( .A1(n14692), .A2(n9871), .ZN(n12806) );
  INV_X2 U12651 ( .A(n15794), .ZN(n9738) );
  INV_X2 U12652 ( .A(n12813), .ZN(n20165) );
  AND2_X2 U12654 ( .A1(n12809), .A2(n14796), .ZN(n14631) );
  NAND3_X1 U12655 ( .A1(n10007), .A2(n10008), .A3(n13373), .ZN(n9895) );
  XNOR2_X2 U12656 ( .A(n9897), .B(n20288), .ZN(n20399) );
  OR2_X1 U12657 ( .A1(n9897), .A2(n20519), .ZN(n12972) );
  NAND2_X1 U12658 ( .A1(n11957), .A2(n9897), .ZN(n13058) );
  NAND2_X1 U12659 ( .A1(n11956), .A2(n11955), .ZN(n9897) );
  OAI21_X1 U12660 ( .B1(n11842), .B2(n9823), .A(n20144), .ZN(n11844) );
  INV_X1 U12661 ( .A(n12809), .ZN(n14653) );
  AND2_X4 U12662 ( .A1(n12789), .A2(n12788), .ZN(n15794) );
  AND3_X4 U12663 ( .A1(n15527), .A2(n10802), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10801) );
  INV_X2 U12664 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10802) );
  AND2_X2 U12665 ( .A1(n13678), .A2(n13296), .ZN(n10781) );
  INV_X1 U12666 ( .A(n10212), .ZN(n10874) );
  INV_X1 U12667 ( .A(n10213), .ZN(n10873) );
  AND2_X2 U12668 ( .A1(n9905), .A2(n10872), .ZN(n10213) );
  NAND4_X1 U12669 ( .A1(n10829), .A2(n10832), .A3(n10831), .A4(n10830), .ZN(
        n9905) );
  NAND2_X1 U12670 ( .A1(n9907), .A2(n9806), .ZN(n9906) );
  NOR2_X1 U12671 ( .A1(n9909), .A2(n9908), .ZN(n9907) );
  NAND2_X1 U12672 ( .A1(n10783), .A2(n10785), .ZN(n9908) );
  NAND3_X1 U12673 ( .A1(n10784), .A2(n10764), .A3(n10765), .ZN(n9909) );
  OR2_X2 U12674 ( .A1(n9990), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15150) );
  NAND2_X1 U12675 ( .A1(n11109), .A2(n9849), .ZN(n9915) );
  INV_X1 U12676 ( .A(n11109), .ZN(n9922) );
  NAND3_X1 U12677 ( .A1(n11662), .A2(n11661), .A3(n14045), .ZN(n11037) );
  NAND2_X1 U12678 ( .A1(n9923), .A2(n10746), .ZN(n10209) );
  XNOR2_X1 U12679 ( .A(n9923), .B(n10746), .ZN(n10762) );
  XNOR2_X2 U12680 ( .A(n11262), .B(n11261), .ZN(n13296) );
  INV_X1 U12681 ( .A(n15517), .ZN(n13678) );
  NAND2_X2 U12682 ( .A1(n9925), .A2(n10145), .ZN(n15464) );
  NAND2_X2 U12683 ( .A1(n15256), .A2(n11693), .ZN(n15246) );
  INV_X1 U12684 ( .A(n10706), .ZN(n16347) );
  NAND2_X1 U12685 ( .A1(n11373), .A2(n11374), .ZN(n9928) );
  NAND4_X1 U12686 ( .A1(n19241), .A2(n10657), .A3(n10680), .A4(n19224), .ZN(
        n11374) );
  NAND3_X1 U12687 ( .A1(n11385), .A2(n9927), .A3(n9926), .ZN(n10721) );
  NAND3_X1 U12688 ( .A1(n16347), .A2(n9929), .A3(n19883), .ZN(n9926) );
  NAND2_X1 U12689 ( .A1(n15126), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11702) );
  INV_X2 U12690 ( .A(n10268), .ZN(n17183) );
  XNOR2_X2 U12691 ( .A(n10356), .B(n10355), .ZN(n17825) );
  NAND2_X2 U12692 ( .A1(n17835), .A2(n10353), .ZN(n10356) );
  NAND2_X1 U12693 ( .A1(n17844), .A2(n10349), .ZN(n17836) );
  XNOR2_X1 U12694 ( .A(n10352), .B(n10351), .ZN(n17837) );
  NAND3_X1 U12695 ( .A1(n10306), .A2(n10307), .A3(n9947), .ZN(n9946) );
  NAND2_X1 U12696 ( .A1(n9954), .A2(n9955), .ZN(n17784) );
  AND2_X1 U12697 ( .A1(n9955), .A2(n9956), .ZN(n17786) );
  NAND2_X1 U12698 ( .A1(n10384), .A2(n10076), .ZN(n9957) );
  NOR2_X2 U12699 ( .A1(n17532), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17531) );
  INV_X2 U12700 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18826) );
  NAND2_X1 U12701 ( .A1(n14642), .A2(n14643), .ZN(n12808) );
  NOR2_X1 U12702 ( .A1(n10103), .A2(n9961), .ZN(n9960) );
  XNOR2_X1 U12703 ( .A(n15794), .B(n9963), .ZN(n14711) );
  NAND3_X1 U12704 ( .A1(n10466), .A2(n10467), .A3(n9976), .ZN(n9975) );
  NAND2_X1 U12705 ( .A1(n9985), .A2(n9984), .ZN(n11046) );
  NAND2_X1 U12706 ( .A1(n15254), .A2(n15255), .ZN(n9985) );
  INV_X1 U12707 ( .A(n9984), .ZN(n9983) );
  INV_X2 U12708 ( .A(n13814), .ZN(n19241) );
  NAND4_X1 U12709 ( .A1(n10613), .A2(n10610), .A3(n10612), .A4(n10611), .ZN(
        n9987) );
  NAND4_X1 U12710 ( .A1(n10618), .A2(n10617), .A3(n10615), .A4(n10616), .ZN(
        n9989) );
  NAND2_X1 U12711 ( .A1(n9997), .A2(n9995), .ZN(n17625) );
  NAND3_X1 U12712 ( .A1(n17757), .A2(n9769), .A3(n10001), .ZN(n17654) );
  XNOR2_X2 U12713 ( .A(n12711), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16525) );
  AND2_X2 U12714 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11728) );
  AOI21_X1 U12715 ( .B1(n12734), .B2(n11938), .A(n11985), .ZN(n11941) );
  OAI21_X2 U12716 ( .B1(n14059), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11887), 
        .ZN(n12734) );
  NAND2_X1 U12717 ( .A1(n20197), .A2(n10121), .ZN(n14059) );
  NAND2_X1 U12718 ( .A1(n20257), .A2(n11875), .ZN(n10121) );
  NAND2_X1 U12719 ( .A1(n10005), .A2(n9825), .ZN(n10006) );
  NAND2_X1 U12720 ( .A1(n15794), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14719) );
  NAND3_X4 U12721 ( .A1(n10015), .A2(n10016), .A3(n11832), .ZN(n20155) );
  NAND2_X1 U12722 ( .A1(n10019), .A2(n10018), .ZN(n13339) );
  NAND2_X1 U12723 ( .A1(n15760), .A2(n9855), .ZN(n14560) );
  NAND2_X1 U12724 ( .A1(n14502), .A2(n10025), .ZN(n10024) );
  NAND2_X1 U12725 ( .A1(n14502), .A2(n14401), .ZN(n14390) );
  NAND2_X1 U12726 ( .A1(n10029), .A2(n10023), .ZN(n14356) );
  NOR2_X1 U12727 ( .A1(n11191), .A2(n10033), .ZN(n15519) );
  INV_X1 U12728 ( .A(n11135), .ZN(n10036) );
  INV_X1 U12729 ( .A(n15159), .ZN(n10037) );
  NAND3_X1 U12730 ( .A1(n10041), .A2(n10040), .A3(n11221), .ZN(n11173) );
  NAND4_X1 U12731 ( .A1(n9777), .A2(n10860), .A3(n10861), .A4(n9821), .ZN(
        n10042) );
  NAND2_X1 U12732 ( .A1(n11173), .A2(n11034), .ZN(n10044) );
  NAND2_X1 U12733 ( .A1(n10047), .A2(n10045), .ZN(n15106) );
  INV_X1 U12734 ( .A(n15118), .ZN(n10046) );
  NAND2_X1 U12735 ( .A1(n14039), .A2(n10050), .ZN(n10047) );
  OR2_X1 U12736 ( .A1(n14039), .A2(n9767), .ZN(n10049) );
  NOR2_X2 U12737 ( .A1(n11089), .A2(n11087), .ZN(n10051) );
  NAND2_X2 U12738 ( .A1(n10987), .A2(n9811), .ZN(n11145) );
  AND2_X1 U12739 ( .A1(n14936), .A2(n15198), .ZN(n10067) );
  XNOR2_X1 U12740 ( .A(n10350), .B(n10508), .ZN(n10352) );
  NAND2_X1 U12741 ( .A1(n17570), .A2(n10378), .ZN(n17560) );
  NOR2_X2 U12742 ( .A1(n17571), .A2(n10073), .ZN(n17550) );
  NAND2_X1 U12743 ( .A1(n10074), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10073) );
  NAND2_X1 U12744 ( .A1(n10077), .A2(n10075), .ZN(n16390) );
  INV_X1 U12745 ( .A(n17531), .ZN(n10077) );
  INV_X1 U12746 ( .A(n17743), .ZN(n10080) );
  NOR2_X2 U12747 ( .A1(n18666), .A2(n10089), .ZN(n17031) );
  NAND3_X1 U12748 ( .A1(n10091), .A2(n15833), .A3(n10090), .ZN(n12785) );
  NAND2_X1 U12749 ( .A1(n15843), .A2(n10092), .ZN(n10091) );
  NAND2_X1 U12750 ( .A1(n11995), .A2(n10097), .ZN(n10096) );
  OAI211_X1 U12751 ( .C1(n11995), .C2(n10099), .A(n10096), .B(n10098), .ZN(
        n12729) );
  NAND2_X1 U12752 ( .A1(n11995), .A2(n20708), .ZN(n10102) );
  NAND2_X1 U12753 ( .A1(n12806), .A2(n9738), .ZN(n14686) );
  INV_X1 U12754 ( .A(n14702), .ZN(n10110) );
  NAND2_X1 U12755 ( .A1(n20079), .A2(n10118), .ZN(n10115) );
  NAND2_X1 U12756 ( .A1(n10115), .A2(n10117), .ZN(n12763) );
  NAND2_X1 U12757 ( .A1(n10121), .A2(n11947), .ZN(n11956) );
  INV_X2 U12758 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11853) );
  INV_X1 U12759 ( .A(n13644), .ZN(n10122) );
  NAND2_X1 U12760 ( .A1(n10122), .A2(n10123), .ZN(n13882) );
  AND2_X2 U12761 ( .A1(n14547), .A2(n9853), .ZN(n14522) );
  NAND3_X1 U12762 ( .A1(n12114), .A2(n12115), .A3(n12130), .ZN(n13607) );
  NAND2_X1 U12763 ( .A1(n14413), .A2(n10130), .ZN(n14376) );
  NAND2_X1 U12764 ( .A1(n14413), .A2(n10132), .ZN(n14403) );
  NAND2_X1 U12765 ( .A1(n10133), .A2(n10715), .ZN(n10751) );
  AND2_X2 U12766 ( .A1(n10751), .A2(n10750), .ZN(n10749) );
  NOR2_X1 U12767 ( .A1(n10134), .A2(n14254), .ZN(n10136) );
  INV_X1 U12768 ( .A(n13226), .ZN(n10142) );
  OAI21_X2 U12769 ( .B1(n15246), .B2(n10144), .A(n10143), .ZN(n16154) );
  OAI21_X2 U12770 ( .B1(n14997), .B2(n10157), .A(n10156), .ZN(n14213) );
  NAND2_X2 U12771 ( .A1(n10213), .A2(n10212), .ZN(n11678) );
  AOI21_X2 U12772 ( .B1(n10166), .B2(n10165), .A(n10163), .ZN(n15402) );
  INV_X1 U12773 ( .A(n10174), .ZN(n16275) );
  OR2_X2 U12774 ( .A1(n15067), .A2(n15055), .ZN(n15057) );
  NAND2_X1 U12775 ( .A1(n14934), .A2(n9866), .ZN(n15082) );
  NAND2_X2 U12776 ( .A1(n11418), .A2(n10186), .ZN(n11639) );
  INV_X4 U12777 ( .A(n10688), .ZN(n14257) );
  INV_X1 U12778 ( .A(n13390), .ZN(n10193) );
  NAND2_X1 U12779 ( .A1(n10193), .A2(n10189), .ZN(n13487) );
  INV_X1 U12780 ( .A(n10195), .ZN(n13457) );
  INV_X1 U12781 ( .A(n10206), .ZN(n13649) );
  OR3_X1 U12782 ( .A1(n14996), .A2(n10208), .A3(n9859), .ZN(n14966) );
  NAND2_X2 U12783 ( .A1(n11151), .A2(n11150), .ZN(n14039) );
  NAND2_X1 U12784 ( .A1(n15160), .A2(n15158), .ZN(n10214) );
  INV_X1 U12785 ( .A(n16160), .ZN(n11059) );
  OAI21_X1 U12788 ( .B1(n13309), .B2(n13308), .A(n13380), .ZN(n19251) );
  OR2_X1 U12789 ( .A1(n12254), .A2(n12595), .ZN(n14879) );
  NAND2_X1 U12790 ( .A1(n11839), .A2(n10231), .ZN(n11840) );
  AND2_X1 U12791 ( .A1(n11926), .A2(n13136), .ZN(n12582) );
  CLKBUF_X1 U12792 ( .A(n13058), .Z(n20520) );
  NAND2_X1 U12793 ( .A1(n12785), .A2(n15832), .ZN(n13739) );
  NAND2_X1 U12794 ( .A1(n11856), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11943) );
  CLKBUF_X1 U12795 ( .A(n15004), .Z(n15011) );
  OR2_X2 U12796 ( .A1(n10779), .A2(n10771), .ZN(n10941) );
  INV_X1 U12797 ( .A(n12863), .ZN(n13120) );
  CLKBUF_X1 U12798 ( .A(n13643), .Z(n13721) );
  NAND2_X1 U12799 ( .A1(n13643), .A2(n13645), .ZN(n13644) );
  AND2_X1 U12800 ( .A1(n15005), .A2(n14188), .ZN(n14163) );
  NAND2_X1 U12801 ( .A1(n15003), .A2(n15002), .ZN(n14993) );
  NAND2_X1 U12802 ( .A1(n13539), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10820) );
  AOI22_X1 U12803 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10633) );
  AND2_X2 U12804 ( .A1(n11730), .A2(n11732), .ZN(n11876) );
  NAND2_X1 U12805 ( .A1(n11267), .A2(n11266), .ZN(n13390) );
  OR2_X1 U12806 ( .A1(n11956), .A2(n11955), .ZN(n11957) );
  OR2_X1 U12807 ( .A1(n12899), .A2(n12900), .ZN(n13156) );
  NAND2_X1 U12808 ( .A1(n12899), .A2(n11197), .ZN(n11646) );
  NAND2_X1 U12809 ( .A1(n14522), .A2(n14524), .ZN(n14513) );
  AND2_X4 U12810 ( .A1(n11729), .A2(n13361), .ZN(n11891) );
  INV_X1 U12811 ( .A(n10786), .ZN(n14274) );
  OR2_X1 U12812 ( .A1(n12720), .A2(n17861), .ZN(n10218) );
  AND3_X1 U12813 ( .A1(n12722), .A2(n12721), .A3(n10218), .ZN(n10219) );
  AND2_X1 U12814 ( .A1(n17230), .A2(n17218), .ZN(n17227) );
  NOR2_X1 U12815 ( .A1(n20457), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10220) );
  NAND2_X1 U12816 ( .A1(n20012), .A2(n14345), .ZN(n20001) );
  OR4_X1 U12817 ( .A1(n15305), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15276), .A4(n15301), .ZN(n10222) );
  AND2_X1 U12818 ( .A1(n17765), .A2(n17967), .ZN(n10223) );
  AND2_X1 U12819 ( .A1(n10342), .A2(n10341), .ZN(n10224) );
  INV_X1 U12820 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13036) );
  OR2_X1 U12821 ( .A1(n19068), .A2(n16301), .ZN(n10225) );
  AND3_X1 U12822 ( .A1(n14042), .A2(n10690), .A3(n13810), .ZN(n10227) );
  INV_X1 U12823 ( .A(n18800), .ZN(n18868) );
  INV_X1 U12824 ( .A(n18868), .ZN(n18869) );
  NAND2_X1 U12825 ( .A1(n10697), .A2(n10680), .ZN(n11199) );
  OR2_X1 U12826 ( .A1(n20012), .A2(n14370), .ZN(n10229) );
  OR2_X1 U12827 ( .A1(n9738), .A2(n15943), .ZN(n10230) );
  XOR2_X1 U12828 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .Z(n10231) );
  OR2_X1 U12829 ( .A1(n15040), .A2(n19241), .ZN(n15026) );
  INV_X1 U12830 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n20990) );
  OR3_X1 U12831 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17579), .ZN(n10232) );
  AND2_X1 U12832 ( .A1(n12325), .A2(n12324), .ZN(n10233) );
  NAND2_X1 U12833 ( .A1(n17689), .A2(n17855), .ZN(n17607) );
  INV_X1 U12834 ( .A(n17607), .ZN(n12712) );
  OR2_X1 U12835 ( .A1(n11465), .A2(n11464), .ZN(n13486) );
  INV_X1 U12836 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13299) );
  INV_X1 U12837 ( .A(n20654), .ZN(n20644) );
  NAND2_X1 U12838 ( .A1(n11978), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12220) );
  INV_X1 U12839 ( .A(n11404), .ZN(n11620) );
  OR2_X1 U12840 ( .A1(n11717), .A2(n19177), .ZN(n10236) );
  AND4_X1 U12841 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n10237) );
  AND3_X1 U12842 ( .A1(n11735), .A2(n11734), .A3(n11733), .ZN(n10239) );
  NOR2_X1 U12843 ( .A1(n20188), .A2(n11980), .ZN(n12075) );
  INV_X1 U12844 ( .A(n12075), .ZN(n11988) );
  AND2_X1 U12845 ( .A1(n11844), .A2(n11843), .ZN(n11871) );
  NAND2_X1 U12846 ( .A1(n20524), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12538) );
  OAI21_X1 U12847 ( .B1(n19409), .B2(n11471), .A(n10820), .ZN(n10821) );
  AOI21_X1 U12848 ( .B1(n19374), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n14257), .ZN(n10758) );
  INV_X1 U12849 ( .A(n10982), .ZN(n10980) );
  INV_X1 U12850 ( .A(n12563), .ZN(n12540) );
  NAND2_X1 U12851 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20568), .ZN(
        n12555) );
  OR2_X1 U12852 ( .A1(n12568), .A2(n12037), .ZN(n12049) );
  INV_X1 U12853 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10893) );
  AND2_X1 U12854 ( .A1(n10744), .A2(n10743), .ZN(n10745) );
  AND2_X1 U12855 ( .A1(n10759), .A2(n10758), .ZN(n10766) );
  AND2_X1 U12856 ( .A1(n11419), .A2(n14257), .ZN(n11373) );
  NAND2_X1 U12857 ( .A1(n17031), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10302) );
  NAND2_X1 U12858 ( .A1(n12541), .A2(n12540), .ZN(n12565) );
  AOI21_X1 U12859 ( .B1(n12539), .B2(n9746), .A(n12542), .ZN(n12573) );
  OR2_X1 U12860 ( .A1(n12094), .A2(n12093), .ZN(n12778) );
  AND2_X1 U12861 ( .A1(n11722), .A2(n11721), .ZN(n11727) );
  AND2_X1 U12862 ( .A1(n10732), .A2(n10731), .ZN(n10733) );
  NAND2_X1 U12863 ( .A1(n10795), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10632) );
  NOR2_X1 U12864 ( .A1(n10234), .A2(n20856), .ZN(n10340) );
  AND2_X1 U12865 ( .A1(n12975), .A2(n12544), .ZN(n12545) );
  AND2_X1 U12866 ( .A1(n11867), .A2(n11866), .ZN(n13142) );
  AOI22_X1 U12867 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11898), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11773) );
  INV_X1 U12868 ( .A(n14307), .ZN(n14277) );
  AOI21_X1 U12869 ( .B1(n10740), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10739), .ZN(n11264) );
  OR2_X1 U12870 ( .A1(n13040), .A2(n11422), .ZN(n11426) );
  INV_X1 U12871 ( .A(n17864), .ZN(n10381) );
  INV_X1 U12872 ( .A(n10299), .ZN(n10307) );
  NAND2_X1 U12873 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12545), .ZN(
        n12841) );
  AND2_X1 U12874 ( .A1(n15655), .A2(n13611), .ZN(n12448) );
  INV_X1 U12875 ( .A(n15753), .ZN(n12177) );
  AND3_X1 U12876 ( .A1(n12816), .A2(n12815), .A3(n12814), .ZN(n12965) );
  NAND2_X1 U12878 ( .A1(n13353), .A2(n11838), .ZN(n13137) );
  INV_X1 U12879 ( .A(n12731), .ZN(n11937) );
  NAND2_X1 U12880 ( .A1(n9819), .A2(n11871), .ZN(n13145) );
  OR2_X1 U12881 ( .A1(n12022), .A2(n12021), .ZN(n12755) );
  AOI22_X1 U12882 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11775) );
  NAND2_X1 U12883 ( .A1(n11149), .A2(n11340), .ZN(n14041) );
  NAND2_X1 U12884 ( .A1(n11055), .A2(n13521), .ZN(n11064) );
  INV_X2 U12885 ( .A(n11341), .ZN(n11362) );
  INV_X1 U12886 ( .A(n14105), .ZN(n14155) );
  NAND2_X1 U12887 ( .A1(n13296), .A2(n16345), .ZN(n13303) );
  INV_X1 U12888 ( .A(n14136), .ZN(n14089) );
  INV_X1 U12889 ( .A(n10689), .ZN(n11380) );
  AND2_X1 U12890 ( .A1(n16130), .A2(n16118), .ZN(n14025) );
  NAND2_X1 U12891 ( .A1(n11406), .A2(n14257), .ZN(n11588) );
  INV_X1 U12892 ( .A(n11435), .ZN(n11679) );
  NOR2_X1 U12893 ( .A1(n18232), .A2(n17238), .ZN(n10538) );
  INV_X1 U12894 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12710) );
  NOR2_X1 U12895 ( .A1(n17679), .A2(n10381), .ZN(n10382) );
  AND2_X1 U12896 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10311) );
  AND2_X1 U12897 ( .A1(n20188), .A2(n12593), .ZN(n11814) );
  INV_X1 U12898 ( .A(n12424), .ZN(n12425) );
  OR2_X1 U12899 ( .A1(n12829), .A2(n14623), .ZN(n12830) );
  NOR2_X1 U12900 ( .A1(n12340), .A2(n14428), .ZN(n12341) );
  INV_X1 U12901 ( .A(n12220), .ZN(n12231) );
  AND2_X1 U12902 ( .A1(n14708), .A2(n14718), .ZN(n15793) );
  INV_X1 U12903 ( .A(n14354), .ZN(n13096) );
  INV_X1 U12904 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12539) );
  AND2_X1 U12905 ( .A1(n10657), .A2(n11034), .ZN(n10675) );
  AND2_X1 U12906 ( .A1(n11260), .A2(n11259), .ZN(n13456) );
  INV_X1 U12907 ( .A(n13225), .ZN(n13224) );
  OR2_X1 U12908 ( .A1(n14213), .A2(n14212), .ZN(n14214) );
  INV_X1 U12909 ( .A(n11620), .ZN(n11637) );
  AND2_X1 U12910 ( .A1(n16315), .A2(n10757), .ZN(n13025) );
  AND2_X1 U12911 ( .A1(n11333), .A2(n11332), .ZN(n14909) );
  OAI211_X1 U12912 ( .C1(n16266), .C2(n16012), .A(n15277), .B(n10222), .ZN(
        n15278) );
  AND2_X1 U12913 ( .A1(n11154), .A2(n15335), .ZN(n15323) );
  NOR2_X1 U12914 ( .A1(n10890), .A2(n10889), .ZN(n10891) );
  AND2_X1 U12915 ( .A1(n11121), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15202) );
  NOR2_X1 U12916 ( .A1(n13428), .A2(n13427), .ZN(n13429) );
  AOI21_X1 U12917 ( .B1(n13078), .B2(n16345), .A(n13074), .ZN(n13075) );
  AOI21_X1 U12918 ( .B1(n17159), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n10276), .ZN(n10277) );
  NOR2_X1 U12919 ( .A1(n18651), .A2(n16391), .ZN(n18094) );
  INV_X1 U12920 ( .A(n18224), .ZN(n13906) );
  NAND2_X1 U12921 ( .A1(n20165), .A2(n20155), .ZN(n12619) );
  AND2_X1 U12922 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12425), .ZN(
        n12426) );
  AND2_X1 U12923 ( .A1(n12665), .A2(n12664), .ZN(n14550) );
  INV_X1 U12924 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15730) );
  INV_X1 U12925 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19919) );
  AND2_X1 U12926 ( .A1(n13616), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13615) );
  INV_X1 U12927 ( .A(n13620), .ZN(n13626) );
  NAND2_X1 U12928 ( .A1(n12490), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12829) );
  INV_X1 U12929 ( .A(n12055), .ZN(n13611) );
  INV_X1 U12930 ( .A(n14425), .ZN(n14544) );
  AND3_X1 U12931 ( .A1(n12129), .A2(n12128), .A3(n12127), .ZN(n13609) );
  INV_X1 U12932 ( .A(n20644), .ZN(n20649) );
  AOI21_X1 U12933 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n15627), .A(
        n15852), .ZN(n15875) );
  OR2_X1 U12934 ( .A1(n15816), .A2(n15815), .ZN(n15813) );
  INV_X1 U12935 ( .A(n20086), .ZN(n20114) );
  NAND2_X1 U12936 ( .A1(n11941), .A2(n11942), .ZN(n11987) );
  INV_X1 U12937 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20524) );
  OR2_X1 U12938 ( .A1(n20137), .A2(n13374), .ZN(n20493) );
  AND2_X1 U12939 ( .A1(n20489), .A2(n11950), .ZN(n20146) );
  INV_X1 U12940 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20568) );
  OR2_X1 U12941 ( .A1(n19030), .A2(n19871), .ZN(n19072) );
  AND2_X1 U12942 ( .A1(n11329), .A2(n11328), .ZN(n14994) );
  OR2_X1 U12943 ( .A1(n11546), .A2(n11545), .ZN(n13651) );
  NAND2_X1 U12944 ( .A1(n14977), .A2(n14214), .ZN(n14233) );
  INV_X1 U12945 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13661) );
  AND2_X1 U12946 ( .A1(n15322), .A2(n11156), .ZN(n14040) );
  OR2_X1 U12947 ( .A1(n16298), .A2(n11655), .ZN(n16272) );
  NAND2_X1 U12948 ( .A1(n13542), .A2(n13541), .ZN(n13543) );
  INV_X1 U12949 ( .A(n19826), .ZN(n19566) );
  INV_X1 U12950 ( .A(n19651), .ZN(n19498) );
  NOR2_X1 U12951 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16794), .ZN(n16777) );
  NAND2_X1 U12952 ( .A1(n18873), .A2(n17392), .ZN(n16512) );
  NOR2_X1 U12953 ( .A1(n13909), .A2(n13908), .ZN(n15537) );
  INV_X1 U12954 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20961) );
  INV_X1 U12955 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17101) );
  INV_X1 U12956 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17158) );
  INV_X1 U12957 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20968) );
  NOR2_X1 U12958 ( .A1(n17581), .A2(n17862), .ZN(n17506) );
  NOR2_X1 U12959 ( .A1(n17974), .A2(n18053), .ZN(n18000) );
  NOR2_X1 U12960 ( .A1(n20927), .A2(n17693), .ZN(n17692) );
  NAND2_X1 U12961 ( .A1(n17601), .A2(n17934), .ZN(n17579) );
  NOR2_X1 U12962 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17765), .ZN(
        n17629) );
  INV_X1 U12963 ( .A(n10367), .ZN(n10365) );
  AOI21_X1 U12964 ( .B1(n18649), .B2(n10500), .A(n15536), .ZN(n10507) );
  INV_X1 U12965 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10351) );
  NOR2_X1 U12966 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18201), .ZN(n18554) );
  AOI22_X1 U12967 ( .A1(n18646), .A2(n18645), .B1(n18650), .B2(n16392), .ZN(
        n18654) );
  NAND2_X1 U12968 ( .A1(n12426), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12451) );
  AND2_X1 U12969 ( .A1(n14417), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19975) );
  INV_X1 U12970 ( .A(n12126), .ZN(n12131) );
  AND2_X1 U12971 ( .A1(n14417), .A2(n13617), .ZN(n19949) );
  AND2_X1 U12972 ( .A1(n14417), .A2(n13615), .ZN(n19982) );
  INV_X1 U12973 ( .A(n20001), .ZN(n20007) );
  AND2_X1 U12974 ( .A1(n20015), .A2(n13112), .ZN(n15771) );
  INV_X1 U12975 ( .A(n13051), .ZN(n20060) );
  AND2_X1 U12976 ( .A1(n13890), .A2(n13889), .ZN(n13892) );
  NAND2_X1 U12977 ( .A1(n12054), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12076) );
  AND2_X1 U12978 ( .A1(n15590), .A2(n13129), .ZN(n20081) );
  AND2_X1 U12979 ( .A1(n20649), .A2(n12824), .ZN(n14666) );
  AND2_X1 U12980 ( .A1(n14393), .A2(n14392), .ZN(n14805) );
  INV_X1 U12981 ( .A(n14819), .ZN(n15859) );
  INV_X1 U12982 ( .A(n14857), .ZN(n20123) );
  OR2_X1 U12983 ( .A1(n12831), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20107) );
  NOR2_X1 U12984 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14032) );
  NOR2_X2 U12985 ( .A1(n20262), .A2(n20516), .ZN(n20218) );
  OR2_X1 U12986 ( .A1(n20223), .A2(n20222), .ZN(n20576) );
  OAI211_X1 U12987 ( .C1(n20230), .C2(n20229), .A(n20228), .B(n20465), .ZN(
        n20252) );
  OAI21_X1 U12988 ( .B1(n20310), .B2(n20295), .A(n20605), .ZN(n20313) );
  AND2_X1 U12989 ( .A1(n20370), .A2(n20321), .ZN(n20364) );
  AND2_X1 U12990 ( .A1(n20370), .A2(n20596), .ZN(n20394) );
  INV_X1 U12991 ( .A(n20404), .ZN(n20425) );
  INV_X1 U12992 ( .A(n20516), .ZN(n20398) );
  NOR2_X2 U12993 ( .A1(n20493), .A2(n20576), .ZN(n20481) );
  INV_X1 U12994 ( .A(n20369), .ZN(n20486) );
  INV_X1 U12995 ( .A(n21072), .ZN(n20564) );
  OR2_X1 U12996 ( .A1(n20223), .A2(n20138), .ZN(n20516) );
  AND2_X1 U12997 ( .A1(n20160), .A2(n20187), .ZN(n20667) );
  AND2_X1 U12998 ( .A1(n20176), .A2(n20187), .ZN(n20685) );
  AND2_X1 U12999 ( .A1(n20188), .A2(n20187), .ZN(n20697) );
  INV_X1 U13000 ( .A(n19030), .ZN(n19061) );
  INV_X1 U13001 ( .A(n19072), .ZN(n19043) );
  AND2_X1 U13002 ( .A1(n19875), .A2(n12902), .ZN(n19030) );
  AND2_X1 U13003 ( .A1(n19152), .A2(n12912), .ZN(n19042) );
  OR2_X1 U13004 ( .A1(n13761), .A2(n13803), .ZN(n13802) );
  OR2_X1 U13005 ( .A1(n11566), .A2(n11565), .ZN(n13633) );
  XNOR2_X1 U13006 ( .A(n14233), .B(n14234), .ZN(n14972) );
  INV_X1 U13007 ( .A(n19150), .ZN(n19143) );
  AND2_X1 U13008 ( .A1(n13650), .A2(n10206), .ZN(n18964) );
  INV_X1 U13009 ( .A(n19177), .ZN(n16200) );
  INV_X1 U13010 ( .A(n16204), .ZN(n19169) );
  INV_X1 U13011 ( .A(n19196), .ZN(n16281) );
  AND2_X1 U13012 ( .A1(n13543), .A2(n19884), .ZN(n19651) );
  AND2_X1 U13013 ( .A1(n16315), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16352) );
  OAI21_X1 U13014 ( .B1(n19206), .B2(n19242), .A(n19651), .ZN(n19245) );
  AND2_X1 U13015 ( .A1(n19251), .A2(n19248), .ZN(n19368) );
  INV_X1 U13016 ( .A(n19337), .ZN(n19329) );
  AND2_X1 U13017 ( .A1(n19368), .A2(n19826), .ZN(n19364) );
  AND2_X1 U13018 ( .A1(n19251), .A2(n19857), .ZN(n19399) );
  AOI22_X1 U13019 ( .A1(n19475), .A2(n19474), .B1(n19473), .B2(n19872), .ZN(
        n19491) );
  NOR2_X1 U13020 ( .A1(n19282), .A2(n19848), .ZN(n19463) );
  NOR2_X1 U13021 ( .A1(n19496), .A2(n19567), .ZN(n19552) );
  NOR2_X1 U13022 ( .A1(n19282), .A2(n19281), .ZN(n19826) );
  NOR2_X2 U13023 ( .A1(n19567), .A2(n19566), .ZN(n19622) );
  AND2_X1 U13024 ( .A1(n13578), .A2(n13577), .ZN(n19639) );
  INV_X1 U13025 ( .A(n19691), .ZN(n19678) );
  OAI22_X1 U13026 ( .A1(n19239), .A2(n19238), .B1(n19237), .B2(n19236), .ZN(
        n19730) );
  INV_X1 U13027 ( .A(n19880), .ZN(n19876) );
  NOR2_X1 U13028 ( .A1(n17392), .A2(n18210), .ZN(n10540) );
  NOR2_X1 U13029 ( .A1(n18682), .A2(n16508), .ZN(n18648) );
  INV_X1 U13030 ( .A(n16855), .ZN(n16874) );
  NOR2_X1 U13031 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16658), .ZN(n16639) );
  NOR2_X1 U13032 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16680), .ZN(n16662) );
  NOR2_X1 U13033 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16703), .ZN(n16684) );
  NOR2_X1 U13034 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16746), .ZN(n16730) );
  NOR2_X1 U13035 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16764), .ZN(n16757) );
  NOR2_X1 U13036 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16821), .ZN(n16804) );
  INV_X1 U13037 ( .A(n16870), .ZN(n16807) );
  NOR2_X2 U13038 ( .A1(n18706), .A2(n16512), .ZN(n16855) );
  NAND2_X1 U13039 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17080), .ZN(n17051) );
  INV_X1 U13040 ( .A(n18240), .ZN(n17218) );
  NOR2_X1 U13041 ( .A1(n17417), .A2(n17308), .ZN(n17304) );
  INV_X2 U13042 ( .A(n9800), .ZN(n17181) );
  NOR2_X1 U13043 ( .A1(n17450), .A2(n17447), .ZN(n17444) );
  INV_X1 U13044 ( .A(n17426), .ZN(n17449) );
  NOR2_X1 U13045 ( .A1(n17505), .A2(n17622), .ZN(n17574) );
  NAND2_X1 U13046 ( .A1(n10556), .A2(n18056), .ZN(n17581) );
  INV_X1 U13047 ( .A(n17839), .ZN(n17849) );
  INV_X1 U13048 ( .A(n10347), .ZN(n17854) );
  INV_X1 U13049 ( .A(n17706), .ZN(n18051) );
  NOR3_X1 U13050 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n16513), .ZN(n18496) );
  NOR2_X1 U13051 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18810), .ZN(
        n18835) );
  NAND2_X1 U13052 ( .A1(n18554), .A2(n18496), .ZN(n18356) );
  INV_X1 U13053 ( .A(n18355), .ZN(n18348) );
  INV_X1 U13054 ( .A(n18377), .ZN(n18370) );
  INV_X1 U13055 ( .A(n18554), .ZN(n18472) );
  INV_X1 U13056 ( .A(n18586), .ZN(n18572) );
  INV_X1 U13057 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18729) );
  NAND2_X1 U13058 ( .A1(n14351), .A2(n12836), .ZN(n12956) );
  AND2_X1 U13059 ( .A1(n12956), .A2(n12932), .ZN(n20798) );
  INV_X1 U13060 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21079) );
  INV_X1 U13061 ( .A(n19949), .ZN(n15751) );
  INV_X1 U13062 ( .A(n19991), .ZN(n19988) );
  NAND2_X2 U13063 ( .A1(n12608), .A2(n12607), .ZN(n20012) );
  OR2_X1 U13064 ( .A1(n13892), .A2(n13891), .ZN(n15817) );
  INV_X1 U13065 ( .A(n15770), .ZN(n20014) );
  INV_X2 U13066 ( .A(n15771), .ZN(n20016) );
  NAND2_X1 U13067 ( .A1(n20051), .A2(n20800), .ZN(n20044) );
  NOR2_X1 U13068 ( .A1(n12956), .A2(n12955), .ZN(n13212) );
  NAND2_X1 U13069 ( .A1(n19900), .A2(n12825), .ZN(n15784) );
  OAI21_X1 U13070 ( .B1(n13892), .B2(n13863), .A(n9780), .ZN(n14743) );
  INV_X1 U13071 ( .A(n15820), .ZN(n20085) );
  INV_X1 U13072 ( .A(n20128), .ZN(n15913) );
  OR2_X1 U13073 ( .A1(n20262), .A2(n20576), .ZN(n20250) );
  AOI22_X1 U13074 ( .A1(n20227), .A2(n20229), .B1(n10220), .B2(n20459), .ZN(
        n20255) );
  NAND2_X1 U13075 ( .A1(n20370), .A2(n20398), .ZN(n20341) );
  AOI22_X1 U13076 ( .A1(n20347), .A2(n20344), .B1(n10220), .B2(n20523), .ZN(
        n20368) );
  NAND2_X1 U13077 ( .A1(n20370), .A2(n20486), .ZN(n20404) );
  NAND2_X1 U13078 ( .A1(n20487), .A2(n20398), .ZN(n20453) );
  AOI22_X1 U13079 ( .A1(n20463), .A2(n20460), .B1(n20459), .B2(n20458), .ZN(
        n20485) );
  NAND2_X1 U13080 ( .A1(n20487), .A2(n20486), .ZN(n21072) );
  AOI22_X1 U13081 ( .A1(n20530), .A2(n20527), .B1(n20523), .B2(n20522), .ZN(
        n21075) );
  OR2_X1 U13082 ( .A1(n20651), .A2(n20516), .ZN(n21071) );
  NAND2_X1 U13083 ( .A1(n20597), .A2(n20596), .ZN(n20705) );
  INV_X1 U13084 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20707) );
  INV_X1 U13085 ( .A(n20786), .ZN(n20783) );
  OR2_X1 U13086 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n19893), .ZN(n20794) );
  INV_X1 U13087 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19746) );
  INV_X1 U13088 ( .A(n19042), .ZN(n19063) );
  AND2_X2 U13089 ( .A1(n13019), .A2(n19737), .ZN(n14992) );
  OR2_X1 U13090 ( .A1(n13807), .A2(n15029), .ZN(n15043) );
  AND2_X1 U13091 ( .A1(n13039), .A2(n19737), .ZN(n19103) );
  NAND2_X1 U13092 ( .A1(n19103), .A2(n10699), .ZN(n19107) );
  INV_X1 U13093 ( .A(n19147), .ZN(n19877) );
  INV_X1 U13094 ( .A(n19148), .ZN(n19146) );
  OR2_X1 U13095 ( .A1(n13156), .A2(n10757), .ZN(n13294) );
  INV_X1 U13096 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16146) );
  INV_X1 U13097 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16170) );
  INV_X1 U13098 ( .A(n19175), .ZN(n19161) );
  INV_X1 U13099 ( .A(n19171), .ZN(n16158) );
  NAND2_X1 U13100 ( .A1(n11704), .A2(n11703), .ZN(n19196) );
  NAND2_X1 U13101 ( .A1(n11704), .A2(n11242), .ZN(n16305) );
  INV_X1 U13102 ( .A(n19192), .ZN(n16266) );
  INV_X1 U13103 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20834) );
  NAND2_X1 U13104 ( .A1(n19463), .A2(n19399), .ZN(n19256) );
  NAND2_X1 U13105 ( .A1(n19463), .A2(n19368), .ZN(n19308) );
  INV_X1 U13106 ( .A(n19364), .ZN(n19342) );
  NAND2_X1 U13107 ( .A1(n19399), .A2(n19369), .ZN(n19398) );
  INV_X1 U13108 ( .A(n19412), .ZN(n19433) );
  OR2_X1 U13109 ( .A1(n19438), .A2(n19434), .ZN(n19495) );
  INV_X1 U13110 ( .A(n19552), .ZN(n19532) );
  NAND2_X1 U13111 ( .A1(n19527), .A2(n19826), .ZN(n19587) );
  NAND2_X1 U13112 ( .A1(n19527), .A2(n19369), .ZN(n19643) );
  NAND2_X1 U13113 ( .A1(n13580), .A2(n19369), .ZN(n19691) );
  INV_X1 U13114 ( .A(n19610), .ZN(n19711) );
  NAND2_X1 U13115 ( .A1(n13580), .A2(n13552), .ZN(n19735) );
  INV_X1 U13116 ( .A(n19824), .ZN(n19744) );
  CLKBUF_X1 U13117 ( .A(n19815), .Z(n19812) );
  INV_X1 U13118 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16513) );
  INV_X1 U13119 ( .A(n16882), .ZN(n16873) );
  INV_X1 U13120 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17693) );
  NOR2_X1 U13121 ( .A1(n16896), .A2(n16895), .ZN(n16923) );
  NOR3_X1 U13122 ( .A1(n17414), .A2(n17416), .A3(n17309), .ZN(n17302) );
  AND2_X1 U13123 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17339), .ZN(n17342) );
  NAND2_X1 U13124 ( .A1(n17447), .A2(n17392), .ZN(n17419) );
  INV_X1 U13125 ( .A(n17447), .ZN(n17452) );
  AOI211_X1 U13126 ( .C1(n18864), .C2(n18855), .A(n17454), .B(n17455), .ZN(
        n17474) );
  INV_X1 U13127 ( .A(n17498), .ZN(n17490) );
  NAND2_X1 U13128 ( .A1(n17474), .A2(n18855), .ZN(n17495) );
  INV_X1 U13129 ( .A(n17708), .ZN(n17704) );
  INV_X1 U13130 ( .A(n17766), .ZN(n17741) );
  NAND2_X1 U13131 ( .A1(n12719), .A2(n18855), .ZN(n17860) );
  NAND2_X1 U13132 ( .A1(n18210), .A2(n12719), .ZN(n17861) );
  INV_X1 U13133 ( .A(n18163), .ZN(n18185) );
  INV_X1 U13134 ( .A(n18164), .ZN(n18169) );
  INV_X1 U13135 ( .A(n18184), .ZN(n18177) );
  INV_X1 U13136 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18696) );
  INV_X1 U13137 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18655) );
  INV_X1 U13138 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18230) );
  INV_X1 U13139 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18268) );
  INV_X1 U13140 ( .A(n16861), .ZN(n18721) );
  INV_X1 U13141 ( .A(n18807), .ZN(n18724) );
  INV_X1 U13142 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18734) );
  INV_X1 U13143 ( .A(n16449), .ZN(n16445) );
  OAI21_X1 U13144 ( .B1(n14629), .B2(n14561), .A(n12706), .ZN(P1_U2842) );
  NAND2_X1 U13145 ( .A1(n12723), .A2(n10219), .ZN(P3_U2799) );
  INV_X1 U13146 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16898) );
  NOR2_X2 U13147 ( .A1(n10245), .A2(n18685), .ZN(n10309) );
  AOI22_X1 U13148 ( .A1(n17177), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10240) );
  OAI21_X1 U13149 ( .B1(n17170), .B2(n16898), .A(n10240), .ZN(n10255) );
  INV_X4 U13150 ( .A(n9796), .ZN(n17159) );
  INV_X4 U13151 ( .A(n10464), .ZN(n17173) );
  AOI22_X1 U13152 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10253) );
  INV_X1 U13153 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16899) );
  INV_X1 U13154 ( .A(n10241), .ZN(n10242) );
  OR2_X2 U13155 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10242), .ZN(
        n10275) );
  AOI22_X1 U13156 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17038), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10243) );
  OAI21_X1 U13157 ( .B1(n10221), .B2(n16899), .A(n10243), .ZN(n10251) );
  NOR3_X1 U13158 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n21016), .ZN(n10244) );
  NAND2_X1 U13159 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10244), .ZN(
        n10301) );
  INV_X1 U13160 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18469) );
  INV_X2 U13161 ( .A(n9798), .ZN(n17185) );
  AOI22_X1 U13162 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U13163 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10248) );
  OAI211_X1 U13164 ( .C1(n17143), .C2(n18469), .A(n10249), .B(n10248), .ZN(
        n10250) );
  AOI211_X1 U13165 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n10251), .B(n10250), .ZN(n10252) );
  OAI211_X1 U13166 ( .C1(n10298), .C2(n20968), .A(n10253), .B(n10252), .ZN(
        n10254) );
  AOI211_X4 U13167 ( .C1(n17181), .C2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n10255), .B(n10254), .ZN(n17358) );
  AOI22_X1 U13168 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10256) );
  OAI21_X1 U13169 ( .B1(n17118), .B2(n18230), .A(n10256), .ZN(n10266) );
  INV_X2 U13170 ( .A(n10221), .ZN(n17138) );
  AOI22_X1 U13171 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10264) );
  INV_X1 U13172 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10257) );
  INV_X1 U13173 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18281) );
  OAI22_X1 U13174 ( .A1(n9800), .A2(n10257), .B1(n10268), .B2(n18281), .ZN(
        n10262) );
  AOI22_X1 U13175 ( .A1(n9733), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10395), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U13176 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10259) );
  INV_X2 U13177 ( .A(n10301), .ZN(n17191) );
  AOI22_X1 U13178 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17031), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10258) );
  NAND3_X1 U13179 ( .A1(n10260), .A2(n10259), .A3(n10258), .ZN(n10261) );
  AOI211_X1 U13180 ( .C1(n9727), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n10262), .B(n10261), .ZN(n10263) );
  OAI211_X1 U13181 ( .C1(n10298), .C2(n20858), .A(n10264), .B(n10263), .ZN(
        n10265) );
  OAI22_X1 U13182 ( .A1(n17118), .A2(n18222), .B1(n10298), .B2(n20882), .ZN(
        n10273) );
  AOI22_X1 U13183 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U13184 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10395), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10270) );
  AOI22_X1 U13185 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10269) );
  NAND3_X1 U13186 ( .A1(n10271), .A2(n10270), .A3(n10269), .ZN(n10272) );
  AOI211_X1 U13187 ( .C1(n10309), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n10273), .B(n10272), .ZN(n10282) );
  INV_X1 U13188 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U13189 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10274) );
  OAI21_X1 U13190 ( .B1(n17170), .B2(n17119), .A(n10274), .ZN(n10280) );
  AOI22_X1 U13191 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17031), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10278) );
  INV_X1 U13192 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17117) );
  NOR2_X1 U13193 ( .A1(n10464), .A2(n17117), .ZN(n10276) );
  NAND2_X1 U13194 ( .A1(n10278), .A2(n10277), .ZN(n10279) );
  AOI22_X1 U13195 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10286) );
  INV_X1 U13196 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10283) );
  AOI21_X1 U13197 ( .B1(n17191), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n10284), .ZN(n10285) );
  NAND2_X1 U13198 ( .A1(n10286), .A2(n10285), .ZN(n10296) );
  INV_X1 U13199 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U13200 ( .A1(n10334), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9733), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10289) );
  AOI22_X1 U13201 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10288) );
  OAI211_X1 U13202 ( .C1(n17188), .C2(n17151), .A(n10289), .B(n10288), .ZN(
        n10295) );
  AOI22_X1 U13203 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U13204 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10395), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10292) );
  AOI22_X1 U13205 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10309), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10291) );
  NAND2_X1 U13206 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10290) );
  NAND4_X1 U13207 ( .A1(n10293), .A2(n10292), .A3(n10291), .A4(n10290), .ZN(
        n10294) );
  INV_X1 U13208 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U13209 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n9795), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n10395), .ZN(n10297) );
  OAI21_X1 U13210 ( .B1(n10298), .B2(n17169), .A(n10297), .ZN(n10299) );
  AOI22_X1 U13211 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17185), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10306) );
  AOI22_X1 U13212 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10334), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10300) );
  INV_X1 U13213 ( .A(n10300), .ZN(n10304) );
  INV_X1 U13214 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n20876) );
  AOI22_X1 U13215 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17104), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17156), .ZN(n10308) );
  AOI22_X1 U13216 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n16998), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n9733), .ZN(n10310) );
  AOI22_X1 U13217 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13218 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10313) );
  AOI22_X1 U13219 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10312) );
  OAI211_X1 U13220 ( .C1(n17188), .C2(n17101), .A(n10313), .B(n10312), .ZN(
        n10319) );
  AOI22_X1 U13221 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13222 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9733), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U13223 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U13224 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10314) );
  NAND4_X1 U13225 ( .A1(n10317), .A2(n10316), .A3(n10315), .A4(n10314), .ZN(
        n10318) );
  AOI211_X1 U13226 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n10319), .B(n10318), .ZN(n10320) );
  NAND2_X1 U13227 ( .A1(n10359), .A2(n10522), .ZN(n10333) );
  INV_X1 U13228 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U13229 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10331) );
  INV_X1 U13230 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U13231 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13232 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10322) );
  OAI211_X1 U13233 ( .C1(n17188), .C2(n17070), .A(n10323), .B(n10322), .ZN(
        n10329) );
  AOI22_X1 U13234 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13235 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13236 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9733), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10325) );
  NAND2_X1 U13237 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10324) );
  NAND4_X1 U13238 ( .A1(n10327), .A2(n10326), .A3(n10325), .A4(n10324), .ZN(
        n10328) );
  AOI211_X1 U13239 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n10329), .B(n10328), .ZN(n10330) );
  NAND2_X4 U13240 ( .A1(n16391), .A2(n16394), .ZN(n17679) );
  INV_X1 U13241 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18820) );
  AOI22_X1 U13242 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17765), .B1(
        n17679), .B2(n18820), .ZN(n10393) );
  NOR2_X1 U13243 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18820), .ZN(
        n10570) );
  INV_X1 U13244 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16387) );
  INV_X1 U13245 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17896) );
  XOR2_X1 U13246 ( .A(n17362), .B(n10332), .Z(n10362) );
  NAND2_X1 U13247 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10362), .ZN(
        n10363) );
  INV_X1 U13248 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21107) );
  XOR2_X1 U13249 ( .A(n17366), .B(n10333), .Z(n17799) );
  NAND2_X1 U13250 ( .A1(n10350), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10349) );
  INV_X1 U13251 ( .A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18450) );
  OAI22_X1 U13252 ( .A1(n17143), .A2(n18450), .B1(n10221), .B2(n17179), .ZN(
        n10339) );
  AOI22_X1 U13253 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13254 ( .A1(n10334), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9733), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13255 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17038), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10335) );
  NAND3_X1 U13256 ( .A1(n10337), .A2(n10336), .A3(n10335), .ZN(n10338) );
  AOI211_X1 U13257 ( .C1(n9727), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n10339), .B(n10338), .ZN(n10346) );
  AOI22_X1 U13258 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10309), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10342) );
  INV_X1 U13259 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n20856) );
  AOI21_X1 U13260 ( .B1(n17159), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n10340), .ZN(n10341) );
  INV_X1 U13261 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17194) );
  AOI22_X1 U13262 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10395), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10343) );
  OAI21_X1 U13263 ( .B1(n9794), .B2(n17194), .A(n10343), .ZN(n10344) );
  INV_X1 U13264 ( .A(n10344), .ZN(n10345) );
  NAND3_X1 U13265 ( .A1(n10346), .A2(n10224), .A3(n10345), .ZN(n10347) );
  INV_X1 U13266 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18838) );
  NOR2_X1 U13267 ( .A1(n17854), .A2(n18838), .ZN(n17853) );
  XNOR2_X1 U13268 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n10348), .ZN(
        n17845) );
  NAND2_X1 U13269 ( .A1(n17853), .A2(n17845), .ZN(n17844) );
  NAND2_X1 U13270 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10352), .ZN(
        n10353) );
  XOR2_X1 U13271 ( .A(n17373), .B(n10354), .Z(n10357) );
  INV_X1 U13272 ( .A(n10357), .ZN(n10355) );
  NAND2_X1 U13273 ( .A1(n10357), .A2(n10356), .ZN(n10358) );
  INV_X1 U13274 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18139) );
  XOR2_X1 U13275 ( .A(n10522), .B(n10359), .Z(n10360) );
  XNOR2_X1 U13276 ( .A(n18139), .B(n10360), .ZN(n17809) );
  NAND2_X1 U13277 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n10360), .ZN(
        n10361) );
  INV_X1 U13278 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18120) );
  XNOR2_X1 U13279 ( .A(n18120), .B(n10362), .ZN(n17785) );
  NAND2_X1 U13280 ( .A1(n10363), .A2(n17784), .ZN(n10366) );
  XNOR2_X1 U13281 ( .A(n10366), .B(n10365), .ZN(n17771) );
  NAND2_X1 U13282 ( .A1(n10367), .A2(n10366), .ZN(n10368) );
  NAND2_X1 U13283 ( .A1(n17770), .A2(n10368), .ZN(n10372) );
  NOR2_X1 U13284 ( .A1(n10372), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10371) );
  NAND2_X1 U13285 ( .A1(n9719), .A2(n17679), .ZN(n17743) );
  INV_X1 U13286 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17731) );
  INV_X1 U13287 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n20895) );
  NOR2_X2 U13288 ( .A1(n17662), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17680) );
  NOR2_X1 U13289 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10369) );
  INV_X1 U13290 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17967) );
  NAND2_X1 U13291 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18059) );
  INV_X1 U13292 ( .A(n18059), .ZN(n17724) );
  NAND2_X1 U13293 ( .A1(n17724), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17706) );
  NAND2_X1 U13294 ( .A1(n18051), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18016) );
  NOR2_X1 U13295 ( .A1(n20895), .A2(n18016), .ZN(n18017) );
  NAND2_X1 U13296 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18017), .ZN(
        n18002) );
  INV_X1 U13297 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18013) );
  NOR2_X1 U13298 ( .A1(n18002), .A2(n18013), .ZN(n10556) );
  INV_X1 U13299 ( .A(n9719), .ZN(n10373) );
  INV_X1 U13300 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17981) );
  NAND2_X1 U13301 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17972) );
  INV_X1 U13302 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17929) );
  NOR2_X1 U13303 ( .A1(n17972), .A2(n17929), .ZN(n17922) );
  INV_X1 U13304 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17961) );
  INV_X1 U13305 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17606) );
  NOR2_X1 U13306 ( .A1(n17961), .A2(n17606), .ZN(n17923) );
  NAND3_X1 U13307 ( .A1(n17922), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n17923), .ZN(n17931) );
  INV_X1 U13308 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17920) );
  NOR2_X1 U13309 ( .A1(n17931), .A2(n17920), .ZN(n17913) );
  INV_X1 U13310 ( .A(n17913), .ZN(n10375) );
  INV_X1 U13311 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20826) );
  NOR2_X1 U13312 ( .A1(n10375), .A2(n20826), .ZN(n17558) );
  NAND2_X1 U13313 ( .A1(n17629), .A2(n17961), .ZN(n10376) );
  INV_X1 U13314 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17934) );
  NAND2_X1 U13315 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17923), .ZN(
        n10379) );
  NOR2_X1 U13316 ( .A1(n10379), .A2(n17920), .ZN(n17932) );
  INV_X1 U13317 ( .A(n17972), .ZN(n17926) );
  NAND2_X1 U13318 ( .A1(n17926), .A2(n10380), .ZN(n17599) );
  NAND2_X1 U13319 ( .A1(n17570), .A2(n17599), .ZN(n17600) );
  NAND3_X1 U13320 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17932), .A3(
        n17600), .ZN(n17571) );
  OAI221_X2 U13321 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17679), 
        .C1(n17896), .C2(n17550), .A(n17549), .ZN(n17532) );
  NOR2_X1 U13322 ( .A1(n17550), .A2(n17679), .ZN(n10383) );
  NAND2_X1 U13323 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17864) );
  NAND3_X1 U13324 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17765), .A3(
        n17521), .ZN(n15548) );
  NOR2_X2 U13325 ( .A1(n16387), .A2(n15548), .ZN(n10388) );
  INV_X1 U13326 ( .A(n10388), .ZN(n10387) );
  INV_X1 U13327 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21105) );
  NOR2_X1 U13328 ( .A1(n17765), .A2(n10389), .ZN(n10390) );
  INV_X1 U13329 ( .A(n10390), .ZN(n10386) );
  NAND2_X1 U13330 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18820), .ZN(
        n10385) );
  OAI211_X1 U13331 ( .C1(n10570), .C2(n10387), .A(n10386), .B(n10385), .ZN(
        n10392) );
  NOR2_X2 U13332 ( .A1(n10389), .A2(n10388), .ZN(n15618) );
  INV_X1 U13333 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16364) );
  NOR2_X2 U13334 ( .A1(n15618), .A2(n16364), .ZN(n15617) );
  OAI21_X1 U13335 ( .B1(n10390), .B2(n15617), .A(n10393), .ZN(n10391) );
  OAI21_X1 U13336 ( .B1(n10393), .B2(n10392), .A(n10391), .ZN(n12709) );
  AOI22_X1 U13337 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n9722), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10394) );
  OAI21_X1 U13338 ( .B1(n20831), .B2(n10464), .A(n10394), .ZN(n10404) );
  INV_X1 U13339 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U13340 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10402) );
  INV_X1 U13341 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17161) );
  OAI22_X1 U13342 ( .A1(n10298), .A2(n17161), .B1(n20881), .B2(n17170), .ZN(
        n10400) );
  AOI22_X1 U13343 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U13344 ( .A1(n17104), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10397) );
  AOI22_X1 U13345 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17038), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10396) );
  NAND3_X1 U13346 ( .A1(n10398), .A2(n10397), .A3(n10396), .ZN(n10399) );
  AOI211_X1 U13347 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n10400), .B(n10399), .ZN(n10401) );
  OAI211_X1 U13348 ( .C1(n10275), .C2(n17025), .A(n10402), .B(n10401), .ZN(
        n10403) );
  AOI22_X1 U13349 ( .A1(n9733), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10414) );
  INV_X1 U13350 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U13351 ( .A1(n17177), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10406) );
  AOI22_X1 U13352 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10405) );
  OAI211_X1 U13353 ( .C1(n17143), .C2(n17137), .A(n10406), .B(n10405), .ZN(
        n10412) );
  AOI22_X1 U13354 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U13355 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U13356 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U13357 ( .A1(n17031), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10407) );
  NAND4_X1 U13358 ( .A1(n10410), .A2(n10409), .A3(n10408), .A4(n10407), .ZN(
        n10411) );
  NOR2_X1 U13359 ( .A1(n18210), .A2(n10537), .ZN(n10488) );
  INV_X1 U13360 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10425) );
  AOI22_X1 U13361 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17031), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10424) );
  INV_X1 U13362 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U13363 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10309), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10416) );
  AOI22_X1 U13364 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10415) );
  OAI211_X1 U13365 ( .C1(n17143), .C2(n16962), .A(n10416), .B(n10415), .ZN(
        n10422) );
  AOI22_X1 U13366 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10420) );
  AOI22_X1 U13367 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10419) );
  AOI22_X1 U13368 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10418) );
  NAND2_X1 U13369 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10417) );
  NAND4_X1 U13370 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n10417), .ZN(
        n10421) );
  AOI211_X1 U13371 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n10422), .B(n10421), .ZN(n10423) );
  NAND2_X1 U13372 ( .A1(n10488), .A2(n17231), .ZN(n10489) );
  INV_X1 U13373 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U13374 ( .A1(n17177), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10426) );
  OAI21_X1 U13375 ( .B1(n17170), .B2(n17042), .A(n10426), .ZN(n10432) );
  AOI22_X1 U13376 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10430) );
  INV_X1 U13377 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18208) );
  OAI22_X1 U13378 ( .A1(n10464), .A2(n18208), .B1(n17143), .B2(n17179), .ZN(
        n10429) );
  AOI22_X1 U13379 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13380 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10427) );
  OAI211_X1 U13381 ( .C1(n9796), .C2(n18268), .A(n10430), .B(n9813), .ZN(
        n10431) );
  NOR2_X1 U13382 ( .A1(n10537), .A2(n10540), .ZN(n10490) );
  AOI22_X1 U13383 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10309), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10433) );
  OAI21_X1 U13384 ( .B1(n17118), .B2(n17101), .A(n10433), .ZN(n10442) );
  AOI22_X1 U13385 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10440) );
  INV_X1 U13386 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n20909) );
  INV_X1 U13387 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16985) );
  OAI22_X1 U13388 ( .A1(n10275), .A2(n20909), .B1(n17170), .B2(n16985), .ZN(
        n10438) );
  AOI22_X1 U13389 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13390 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10435) );
  AOI22_X1 U13391 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17031), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10434) );
  NAND3_X1 U13392 ( .A1(n10436), .A2(n10435), .A3(n10434), .ZN(n10437) );
  AOI211_X1 U13393 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n10438), .B(n10437), .ZN(n10439) );
  OAI211_X1 U13394 ( .C1(n9794), .C2(n20841), .A(n10440), .B(n10439), .ZN(
        n10441) );
  AOI211_X2 U13395 ( .C1(n17155), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n10442), .B(n10441), .ZN(n18224) );
  INV_X1 U13396 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16969) );
  OAI22_X1 U13397 ( .A1(n10464), .A2(n18230), .B1(n17170), .B2(n16969), .ZN(
        n10452) );
  AOI22_X1 U13398 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U13399 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10449) );
  INV_X1 U13400 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17087) );
  AOI22_X1 U13401 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10443) );
  OAI21_X1 U13402 ( .B1(n10298), .B2(n17087), .A(n10443), .ZN(n10447) );
  AOI22_X1 U13403 ( .A1(n16998), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13404 ( .A1(n17177), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10444) );
  OAI211_X1 U13405 ( .C1(n17188), .C2(n20858), .A(n10445), .B(n10444), .ZN(
        n10446) );
  AOI211_X1 U13406 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n10447), .B(n10446), .ZN(n10448) );
  NAND3_X1 U13407 ( .A1(n10450), .A2(n10449), .A3(n10448), .ZN(n10451) );
  NOR2_X1 U13408 ( .A1(n18227), .A2(n17231), .ZN(n15644) );
  INV_X1 U13409 ( .A(n15644), .ZN(n18669) );
  INV_X1 U13410 ( .A(n17231), .ZN(n18232) );
  INV_X1 U13411 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13945) );
  AOI22_X1 U13412 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10453) );
  OAI21_X1 U13413 ( .B1(n9800), .B2(n13945), .A(n10453), .ZN(n10462) );
  AOI22_X1 U13414 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10460) );
  INV_X1 U13415 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17062) );
  OAI22_X1 U13416 ( .A1(n17170), .A2(n17062), .B1(n17188), .B2(n20968), .ZN(
        n10458) );
  AOI22_X1 U13417 ( .A1(n17104), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10456) );
  AOI22_X1 U13418 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10455) );
  AOI22_X1 U13419 ( .A1(n9795), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10454) );
  NAND3_X1 U13420 ( .A1(n10456), .A2(n10455), .A3(n10454), .ZN(n10457) );
  AOI211_X1 U13421 ( .C1(n17182), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n10458), .B(n10457), .ZN(n10459) );
  OAI211_X1 U13422 ( .C1(n10464), .C2(n21001), .A(n10460), .B(n10459), .ZN(
        n10461) );
  AOI211_X4 U13423 ( .C1(n9722), .C2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A(
        n10462), .B(n10461), .ZN(n18240) );
  AOI22_X1 U13424 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n10309), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10463) );
  OAI21_X1 U13425 ( .B1(n10464), .B2(n18222), .A(n10463), .ZN(n10470) );
  INV_X1 U13426 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17120) );
  AOI22_X1 U13427 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10469) );
  AOI22_X1 U13428 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9795), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10465) );
  OAI21_X1 U13429 ( .B1(n10298), .B2(n17119), .A(n10465), .ZN(n10468) );
  AOI22_X1 U13430 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U13431 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10466) );
  INV_X1 U13432 ( .A(n10552), .ZN(n10471) );
  AOI211_X1 U13433 ( .C1(n13906), .C2(n18669), .A(n10538), .B(n10471), .ZN(
        n10472) );
  NAND2_X1 U13434 ( .A1(n10490), .A2(n10472), .ZN(n10498) );
  INV_X1 U13435 ( .A(n16392), .ZN(n18651) );
  OAI22_X1 U13436 ( .A1(n18834), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n18675), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10504) );
  NAND2_X1 U13437 ( .A1(n18674), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10485) );
  NOR2_X1 U13438 ( .A1(n10504), .A2(n10485), .ZN(n10473) );
  AOI21_X1 U13439 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18675), .A(
        n10473), .ZN(n10478) );
  AOI22_X1 U13440 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18197), .B2(n18826), .ZN(
        n10477) );
  NOR2_X1 U13441 ( .A1(n10478), .A2(n10477), .ZN(n10474) );
  AOI21_X1 U13442 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18197), .A(
        n10474), .ZN(n10475) );
  AOI22_X1 U13443 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18655), .B1(
        n10475), .B2(n18819), .ZN(n10480) );
  NOR2_X1 U13444 ( .A1(n10475), .A2(n18819), .ZN(n10479) );
  NAND2_X1 U13445 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18655), .ZN(
        n10476) );
  OAI22_X1 U13446 ( .A1(n10480), .A2(n18696), .B1(n10479), .B2(n10476), .ZN(
        n10483) );
  XNOR2_X1 U13447 ( .A(n10478), .B(n10477), .ZN(n10486) );
  XNOR2_X1 U13448 ( .A(n10504), .B(n10485), .ZN(n10482) );
  INV_X1 U13449 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20840) );
  OR2_X1 U13450 ( .A1(n10479), .A2(n18696), .ZN(n10481) );
  AOI22_X1 U13451 ( .A1(n20840), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n10481), .B2(n10480), .ZN(n10501) );
  INV_X1 U13452 ( .A(n10483), .ZN(n10484) );
  OAI211_X1 U13453 ( .C1(n18674), .C2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10485), .B(n10484), .ZN(n10503) );
  NOR2_X1 U13454 ( .A1(n10486), .A2(n10503), .ZN(n12708) );
  INV_X1 U13455 ( .A(n10537), .ZN(n18214) );
  NOR2_X2 U13456 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18729), .ZN(n18800) );
  OAI211_X1 U13457 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(P3_STATE_REG_1__SCAN_IN), .A(n18734), .B(n18794), .ZN(n18732) );
  OAI21_X1 U13458 ( .B1(n18214), .B2(n18855), .A(n18732), .ZN(n10487) );
  NAND2_X1 U13459 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18707) );
  OAI21_X1 U13460 ( .B1(n10488), .B2(n10487), .A(n18707), .ZN(n16491) );
  OAI22_X1 U13461 ( .A1(n12708), .A2(n10489), .B1(n10545), .B2(n16491), .ZN(
        n10500) );
  NAND2_X1 U13462 ( .A1(n17238), .A2(n17231), .ZN(n10496) );
  NOR2_X1 U13463 ( .A1(n10537), .A2(n10496), .ZN(n10505) );
  NOR2_X1 U13464 ( .A1(n10544), .A2(n10505), .ZN(n10495) );
  AOI22_X1 U13465 ( .A1(n18219), .A2(n10497), .B1(n18224), .B2(n15644), .ZN(
        n10494) );
  NAND2_X1 U13466 ( .A1(n17218), .A2(n10496), .ZN(n10492) );
  INV_X1 U13467 ( .A(n10490), .ZN(n10491) );
  AOI22_X1 U13468 ( .A1(n10492), .A2(n13906), .B1(n10491), .B2(n10496), .ZN(
        n10493) );
  OAI211_X1 U13469 ( .C1(n10495), .C2(n17392), .A(n10494), .B(n10493), .ZN(
        n10546) );
  INV_X1 U13470 ( .A(n18219), .ZN(n10548) );
  NAND2_X1 U13471 ( .A1(n10549), .A2(n10537), .ZN(n10539) );
  OAI21_X1 U13472 ( .B1(n10498), .B2(n10546), .A(n10539), .ZN(n10499) );
  NOR2_X1 U13473 ( .A1(n18855), .A2(n18204), .ZN(n10536) );
  OAI21_X1 U13474 ( .B1(n18240), .B2(n15644), .A(n10536), .ZN(n10543) );
  NAND2_X1 U13475 ( .A1(n10499), .A2(n10543), .ZN(n15536) );
  OAI211_X1 U13476 ( .C1(n10504), .C2(n10503), .A(n10502), .B(n10501), .ZN(
        n13909) );
  INV_X1 U13477 ( .A(n13909), .ZN(n18646) );
  OAI21_X1 U13478 ( .B1(n10505), .B2(n13906), .A(n18646), .ZN(n10506) );
  NOR2_X1 U13479 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18859), .ZN(n18718) );
  NAND2_X1 U13480 ( .A1(n18718), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18713) );
  NOR3_X4 U13481 ( .A1(n17358), .A2(n18651), .A3(n18185), .ZN(n18099) );
  NAND2_X1 U13482 ( .A1(n12709), .A2(n18099), .ZN(n10575) );
  NOR2_X1 U13483 ( .A1(n17854), .A2(n10350), .ZN(n10515) );
  NOR2_X1 U13484 ( .A1(n10515), .A2(n10508), .ZN(n10513) );
  NOR2_X1 U13485 ( .A1(n10513), .A2(n17373), .ZN(n10523) );
  NAND2_X1 U13486 ( .A1(n10523), .A2(n10522), .ZN(n10511) );
  NOR2_X1 U13487 ( .A1(n17366), .A2(n10511), .ZN(n10510) );
  NAND2_X1 U13488 ( .A1(n10510), .A2(n17362), .ZN(n10509) );
  NOR2_X1 U13489 ( .A1(n17358), .A2(n10509), .ZN(n10533) );
  XNOR2_X1 U13490 ( .A(n10509), .B(n16391), .ZN(n17777) );
  XOR2_X1 U13491 ( .A(n10510), .B(n17362), .Z(n10527) );
  XOR2_X1 U13492 ( .A(n10511), .B(n17366), .Z(n10512) );
  NAND2_X1 U13493 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n10512), .ZN(
        n10525) );
  XNOR2_X1 U13494 ( .A(n21107), .B(n10512), .ZN(n17796) );
  XOR2_X1 U13495 ( .A(n10513), .B(n17373), .Z(n10514) );
  NAND2_X1 U13496 ( .A1(n10514), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10520) );
  INV_X1 U13497 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18151) );
  XNOR2_X1 U13498 ( .A(n18151), .B(n10514), .ZN(n17821) );
  XOR2_X1 U13499 ( .A(n17379), .B(n10515), .Z(n10516) );
  NAND2_X1 U13500 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10516), .ZN(
        n10519) );
  XOR2_X1 U13501 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10516), .Z(
        n17834) );
  AOI21_X1 U13502 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10348), .A(
        n10347), .ZN(n10518) );
  NOR2_X1 U13503 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n10348), .ZN(
        n10517) );
  AOI221_X1 U13504 ( .B1(n10347), .B2(n10348), .C1(n10518), .C2(n18838), .A(
        n10517), .ZN(n17833) );
  NAND2_X1 U13505 ( .A1(n17834), .A2(n17833), .ZN(n17832) );
  NAND2_X1 U13506 ( .A1(n10519), .A2(n17832), .ZN(n17820) );
  NAND2_X1 U13507 ( .A1(n17821), .A2(n17820), .ZN(n17819) );
  NAND2_X1 U13508 ( .A1(n10520), .A2(n17819), .ZN(n10521) );
  NAND2_X1 U13509 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n10521), .ZN(
        n10524) );
  XOR2_X1 U13510 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n10521), .Z(
        n17812) );
  INV_X1 U13511 ( .A(n10522), .ZN(n17370) );
  XNOR2_X1 U13512 ( .A(n10523), .B(n17370), .ZN(n17811) );
  NAND2_X1 U13513 ( .A1(n17812), .A2(n17811), .ZN(n17810) );
  NAND2_X1 U13514 ( .A1(n10524), .A2(n17810), .ZN(n17795) );
  NAND2_X1 U13515 ( .A1(n17796), .A2(n17795), .ZN(n17794) );
  NAND2_X1 U13516 ( .A1(n10525), .A2(n17794), .ZN(n10526) );
  NAND2_X1 U13517 ( .A1(n10527), .A2(n10526), .ZN(n10528) );
  XOR2_X1 U13518 ( .A(n10527), .B(n10526), .Z(n17783) );
  NAND2_X1 U13519 ( .A1(n17783), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17782) );
  INV_X1 U13520 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18106) );
  NAND2_X1 U13521 ( .A1(n10533), .A2(n10529), .ZN(n10534) );
  INV_X1 U13522 ( .A(n10529), .ZN(n10532) );
  NAND2_X1 U13523 ( .A1(n17777), .A2(n17776), .ZN(n10531) );
  NAND2_X1 U13524 ( .A1(n10533), .A2(n10532), .ZN(n10530) );
  OAI211_X1 U13525 ( .C1(n10533), .C2(n10532), .A(n10531), .B(n10530), .ZN(
        n17756) );
  NAND2_X1 U13526 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17756), .ZN(
        n17755) );
  INV_X1 U13527 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17876) );
  INV_X1 U13528 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17904) );
  NOR2_X1 U13529 ( .A1(n20826), .A2(n17904), .ZN(n17883) );
  NAND2_X1 U13530 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17883), .ZN(
        n17538) );
  NOR2_X1 U13531 ( .A1(n17876), .A2(n17538), .ZN(n10563) );
  NAND2_X1 U13532 ( .A1(n17913), .A2(n10563), .ZN(n17862) );
  NAND2_X1 U13533 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16396) );
  NOR2_X1 U13534 ( .A1(n16396), .A2(n16387), .ZN(n15616) );
  NAND3_X1 U13535 ( .A1(n17506), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15616), .ZN(n10535) );
  XOR2_X1 U13536 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n10535), .Z(
        n12720) );
  OR2_X1 U13537 ( .A1(n10540), .A2(n10536), .ZN(n18871) );
  NOR2_X1 U13538 ( .A1(n18224), .A2(n17231), .ZN(n18662) );
  NAND3_X1 U13539 ( .A1(n10552), .A2(n10545), .A3(n18662), .ZN(n13908) );
  NAND2_X1 U13540 ( .A1(n18661), .A2(n10538), .ZN(n13907) );
  NAND2_X1 U13541 ( .A1(n10540), .A2(n16492), .ZN(n10550) );
  OAI21_X1 U13542 ( .B1(n10545), .B2(n10544), .A(n10543), .ZN(n10547) );
  NAND2_X1 U13543 ( .A1(n18855), .A2(n10550), .ZN(n15534) );
  NAND2_X1 U13544 ( .A1(n9766), .A2(n18163), .ZN(n18145) );
  NAND3_X1 U13545 ( .A1(n15616), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n18820), .ZN(n10560) );
  INV_X1 U13546 ( .A(n10560), .ZN(n10561) );
  NAND3_X1 U13547 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10555) );
  INV_X1 U13548 ( .A(n10555), .ZN(n10553) );
  AOI21_X1 U13549 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18158) );
  NAND3_X1 U13550 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10554) );
  NOR2_X1 U13551 ( .A1(n18158), .A2(n10554), .ZN(n18086) );
  NAND2_X1 U13552 ( .A1(n10553), .A2(n18086), .ZN(n18054) );
  NOR2_X1 U13553 ( .A1(n17974), .A2(n18054), .ZN(n17925) );
  NAND2_X1 U13554 ( .A1(n17913), .A2(n17925), .ZN(n10565) );
  INV_X1 U13555 ( .A(n10565), .ZN(n10558) );
  INV_X1 U13556 ( .A(n18673), .ZN(n18171) );
  INV_X1 U13557 ( .A(n10554), .ZN(n18090) );
  NAND3_X1 U13558 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18090), .ZN(n18084) );
  NOR2_X1 U13559 ( .A1(n18084), .A2(n10555), .ZN(n17921) );
  NAND2_X1 U13560 ( .A1(n10556), .A2(n17921), .ZN(n17968) );
  INV_X1 U13561 ( .A(n17968), .ZN(n17927) );
  NAND2_X1 U13562 ( .A1(n17913), .A2(n17927), .ZN(n17863) );
  AOI221_X1 U13563 ( .B1(n18670), .B2(n18171), .C1(n18838), .C2(n18171), .A(
        n17863), .ZN(n10557) );
  AOI21_X1 U13564 ( .B1(n18658), .B2(n10558), .A(n10557), .ZN(n17884) );
  INV_X1 U13565 ( .A(n10563), .ZN(n10566) );
  NOR2_X1 U13566 ( .A1(n17884), .A2(n10566), .ZN(n15551) );
  INV_X1 U13567 ( .A(n17862), .ZN(n16361) );
  NAND2_X1 U13568 ( .A1(n16361), .A2(n18000), .ZN(n16395) );
  INV_X1 U13569 ( .A(n16395), .ZN(n17867) );
  NAND2_X1 U13570 ( .A1(n15616), .A2(n17867), .ZN(n16362) );
  OAI21_X1 U13571 ( .B1(n16364), .B2(n16362), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10559) );
  OAI21_X1 U13572 ( .B1(n10560), .B2(n16395), .A(n10559), .ZN(n12718) );
  AOI22_X1 U13573 ( .A1(n10561), .A2(n15551), .B1(n18094), .B2(n12718), .ZN(
        n10562) );
  OAI22_X1 U13574 ( .A1(n12720), .A2(n18145), .B1(n10562), .B2(n18185), .ZN(
        n10573) );
  INV_X1 U13575 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n17857) );
  NAND2_X1 U13576 ( .A1(n17857), .A2(n18810), .ZN(n18829) );
  NOR2_X1 U13577 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18829), .ZN(n18874) );
  NAND2_X2 U13578 ( .A1(n18874), .A2(n18859), .ZN(n18179) );
  AOI221_X1 U13579 ( .B1(n17862), .B2(n18673), .C1(n17968), .C2(n18673), .A(
        n18164), .ZN(n10568) );
  OR2_X1 U13580 ( .A1(n18838), .A2(n17863), .ZN(n10564) );
  NAND2_X1 U13581 ( .A1(n10563), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16389) );
  INV_X1 U13582 ( .A(n18670), .ZN(n18015) );
  OAI21_X1 U13583 ( .B1(n10564), .B2(n16389), .A(n18015), .ZN(n10567) );
  NAND2_X1 U13584 ( .A1(n18658), .A2(n10565), .ZN(n17901) );
  NAND2_X1 U13585 ( .A1(n18658), .A2(n10566), .ZN(n17865) );
  NAND4_X1 U13586 ( .A1(n10568), .A2(n10567), .A3(n17901), .A4(n17865), .ZN(
        n15543) );
  INV_X1 U13587 ( .A(n15616), .ZN(n10569) );
  OAI221_X1 U13588 ( .B1(n15543), .B2(n18088), .C1(n15543), .C2(n10569), .A(
        n18179), .ZN(n15619) );
  NAND2_X1 U13589 ( .A1(n18088), .A2(n18163), .ZN(n18170) );
  INV_X1 U13590 ( .A(n18170), .ZN(n18132) );
  INV_X1 U13591 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n21051) );
  NOR2_X1 U13592 ( .A1(n21051), .A2(n18179), .ZN(n12717) );
  AOI21_X1 U13593 ( .B1(n10570), .B2(n18132), .A(n12717), .ZN(n10571) );
  OAI21_X1 U13594 ( .B1(n15619), .B2(n18820), .A(n10571), .ZN(n10572) );
  NOR2_X1 U13595 ( .A1(n10573), .A2(n10572), .ZN(n10574) );
  NAND2_X1 U13596 ( .A1(n10575), .A2(n10574), .ZN(P3_U2831) );
  INV_X1 U13597 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U13598 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__5__SCAN_IN), .B2(n10639), .ZN(n10579) );
  AOI22_X1 U13599 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14125), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10578) );
  AND2_X2 U13600 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10787) );
  AND2_X4 U13601 ( .A1(n10787), .A2(n15527), .ZN(n14166) );
  AND2_X2 U13602 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11191) );
  AOI22_X1 U13603 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10795), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10577) );
  AND2_X4 U13604 ( .A1(n10789), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10786) );
  AND2_X4 U13605 ( .A1(n10787), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10793) );
  AOI22_X1 U13606 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10793), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10576) );
  NAND4_X1 U13607 ( .A1(n10579), .A2(n10578), .A3(n10577), .A4(n10576), .ZN(
        n10580) );
  AOI22_X1 U13608 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10584) );
  AOI22_X1 U13609 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10583) );
  AOI22_X1 U13610 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10793), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10582) );
  AOI22_X1 U13611 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14303), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10581) );
  NAND4_X1 U13612 ( .A1(n10584), .A2(n10583), .A3(n10582), .A4(n10581), .ZN(
        n10585) );
  AOI22_X1 U13613 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10587) );
  AOI22_X1 U13614 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9718), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10586) );
  AND3_X1 U13615 ( .A1(n10587), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10586), .ZN(n10590) );
  AOI22_X1 U13616 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10589) );
  AOI22_X1 U13617 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14125), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10588) );
  NAND3_X1 U13618 ( .A1(n10590), .A2(n10589), .A3(n10588), .ZN(n10597) );
  AOI22_X1 U13619 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9718), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13620 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9760), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10591) );
  AND3_X1 U13621 ( .A1(n10592), .A2(n10614), .A3(n10591), .ZN(n10595) );
  AOI22_X1 U13622 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9763), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10594) );
  AOI22_X1 U13623 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10593) );
  NAND3_X1 U13624 ( .A1(n10595), .A2(n10594), .A3(n10593), .ZN(n10596) );
  INV_X2 U13625 ( .A(n14309), .ZN(n14303) );
  AOI22_X1 U13626 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9764), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10602) );
  AOI22_X1 U13627 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14166), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10599) );
  AOI22_X1 U13628 ( .A1(n9718), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10598) );
  AND2_X1 U13629 ( .A1(n10599), .A2(n10598), .ZN(n10601) );
  AOI22_X1 U13630 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10600) );
  NAND3_X1 U13631 ( .A1(n10602), .A2(n10601), .A3(n10600), .ZN(n10603) );
  AOI22_X1 U13632 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13633 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14303), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13634 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14166), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13635 ( .A1(n10793), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10604) );
  NAND4_X1 U13636 ( .A1(n10607), .A2(n10606), .A3(n10605), .A4(n10604), .ZN(
        n10608) );
  INV_X2 U13637 ( .A(n10609), .ZN(n10657) );
  AOI22_X1 U13638 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10663), .B1(
        n10639), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13639 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10795), .B1(
        n14166), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13640 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9718), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13641 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n10639), .ZN(n10618) );
  AOI22_X1 U13642 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14125), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13643 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9718), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13644 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9760), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13645 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9764), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10622) );
  AOI22_X1 U13646 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n10639), .ZN(n10621) );
  AOI22_X1 U13647 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10793), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13648 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10795), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13649 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10793), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13650 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10795), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10624) );
  AND3_X1 U13651 ( .A1(n10625), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10624), .ZN(n10628) );
  AOI22_X1 U13652 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__4__SCAN_IN), .B2(n10639), .ZN(n10627) );
  AOI22_X1 U13653 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14303), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10626) );
  NAND3_X1 U13654 ( .A1(n10628), .A2(n10627), .A3(n10626), .ZN(n10629) );
  NAND2_X1 U13655 ( .A1(n19224), .A2(n13814), .ZN(n10656) );
  AOI22_X1 U13656 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14303), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10635) );
  AOI22_X1 U13657 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10793), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10634) );
  NAND4_X1 U13658 ( .A1(n10636), .A2(n10635), .A3(n10634), .A4(n10633), .ZN(
        n10645) );
  NAND2_X1 U13659 ( .A1(n10795), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10638) );
  AOI22_X1 U13660 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9763), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U13661 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10793), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U13662 ( .A1(n10663), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n10639), .ZN(n10640) );
  NAND4_X1 U13663 ( .A1(n10643), .A2(n10642), .A3(n10641), .A4(n10640), .ZN(
        n10644) );
  AOI22_X1 U13664 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13665 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9764), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13666 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10793), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10647) );
  AOI22_X1 U13667 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10795), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10646) );
  NAND4_X1 U13668 ( .A1(n10649), .A2(n10648), .A3(n10647), .A4(n10646), .ZN(
        n10655) );
  AOI22_X1 U13669 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13670 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14125), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10652) );
  AOI22_X1 U13671 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10793), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13672 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10795), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10650) );
  NAND4_X1 U13673 ( .A1(n10653), .A2(n10652), .A3(n10651), .A4(n10650), .ZN(
        n10654) );
  NAND2_X1 U13674 ( .A1(n10689), .A2(n10672), .ZN(n11198) );
  NOR2_X2 U13675 ( .A1(n10656), .A2(n11198), .ZN(n10658) );
  NAND2_X1 U13676 ( .A1(n10658), .A2(n10675), .ZN(n11195) );
  AND2_X2 U13677 ( .A1(n10658), .A2(n10679), .ZN(n10706) );
  AOI22_X1 U13678 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9763), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13679 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10661) );
  AOI22_X1 U13680 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10793), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10660) );
  AOI22_X1 U13681 ( .A1(n14166), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10795), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10659) );
  NAND4_X1 U13682 ( .A1(n10662), .A2(n10661), .A3(n10660), .A4(n10659), .ZN(
        n10669) );
  AOI22_X1 U13683 ( .A1(n10801), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14303), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13684 ( .A1(n10639), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10663), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13685 ( .A1(n10786), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9760), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13686 ( .A1(n10793), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14166), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10664) );
  NAND4_X1 U13687 ( .A1(n10667), .A2(n10666), .A3(n10665), .A4(n10664), .ZN(
        n10668) );
  MUX2_X2 U13688 ( .A(n10669), .B(n10668), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19883) );
  MUX2_X1 U13689 ( .A(n10657), .B(n13814), .S(n9726), .Z(n10671) );
  NAND2_X1 U13690 ( .A1(n11419), .A2(n10711), .ZN(n10670) );
  NAND4_X1 U13691 ( .A1(n10671), .A2(n10689), .A3(n10680), .A4(n10670), .ZN(
        n10678) );
  INV_X1 U13692 ( .A(n13814), .ZN(n10673) );
  NAND3_X1 U13693 ( .A1(n10676), .A2(n10675), .A3(n10674), .ZN(n10686) );
  AND2_X1 U13694 ( .A1(n10686), .A2(n9730), .ZN(n10677) );
  NAND2_X1 U13695 ( .A1(n10678), .A2(n10677), .ZN(n11385) );
  NAND2_X1 U13696 ( .A1(n10721), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10685) );
  INV_X1 U13697 ( .A(n10679), .ZN(n10697) );
  NAND2_X1 U13698 ( .A1(n11199), .A2(n19224), .ZN(n10682) );
  NAND2_X1 U13699 ( .A1(n11206), .A2(n13814), .ZN(n11371) );
  INV_X2 U13700 ( .A(n10711), .ZN(n19218) );
  INV_X1 U13701 ( .A(n11383), .ZN(n10683) );
  INV_X1 U13702 ( .A(n11228), .ZN(n10712) );
  NAND2_X1 U13703 ( .A1(n10728), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10694) );
  NAND2_X1 U13704 ( .A1(n10706), .A2(n19883), .ZN(n12899) );
  INV_X1 U13705 ( .A(n10686), .ZN(n10687) );
  NAND2_X1 U13706 ( .A1(n10687), .A2(n9730), .ZN(n11197) );
  INV_X1 U13707 ( .A(n11646), .ZN(n10692) );
  INV_X1 U13708 ( .A(n11381), .ZN(n10691) );
  NOR2_X1 U13709 ( .A1(n10711), .A2(n11380), .ZN(n10690) );
  AND2_X1 U13710 ( .A1(n13814), .A2(n10657), .ZN(n13810) );
  NOR2_X1 U13711 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19873) );
  AOI22_X1 U13712 ( .A1(n10695), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19873), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10693) );
  NAND2_X1 U13713 ( .A1(n10695), .A2(n14257), .ZN(n10704) );
  NAND2_X2 U13714 ( .A1(n11381), .A2(n12907), .ZN(n11376) );
  NAND2_X2 U13715 ( .A1(n10704), .A2(n13319), .ZN(n11243) );
  INV_X1 U13716 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15510) );
  NOR2_X1 U13717 ( .A1(n12907), .A2(n11380), .ZN(n10705) );
  AOI22_X1 U13718 ( .A1(n11248), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10708) );
  OAI21_X2 U13719 ( .B1(n9752), .B2(n15510), .A(n10710), .ZN(n10726) );
  NOR2_X1 U13720 ( .A1(n10712), .A2(n10711), .ZN(n10713) );
  INV_X1 U13721 ( .A(n19873), .ZN(n10717) );
  OAI22_X1 U13722 ( .A1(n13319), .A2(n19884), .B1(n10717), .B2(n19861), .ZN(
        n10714) );
  INV_X1 U13723 ( .A(n10714), .ZN(n10715) );
  INV_X1 U13724 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16301) );
  INV_X1 U13725 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19060) );
  NAND2_X1 U13726 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10716) );
  OAI211_X1 U13727 ( .C1(n10742), .C2(n19060), .A(n10717), .B(n10716), .ZN(
        n10718) );
  AOI21_X1 U13728 ( .B1(n11272), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10718), .ZN(
        n10724) );
  NOR2_X1 U13729 ( .A1(n9745), .A2(n10719), .ZN(n10722) );
  OAI21_X1 U13730 ( .B1(n10722), .B2(n10721), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10723) );
  OAI211_X1 U13731 ( .C1(n9753), .C2(n16301), .A(n10724), .B(n10723), .ZN(
        n10750) );
  INV_X1 U13732 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n11189) );
  OAI21_X1 U13733 ( .B1(n19845), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11189), 
        .ZN(n10729) );
  INV_X1 U13734 ( .A(n9753), .ZN(n10730) );
  NAND2_X1 U13735 ( .A1(n11272), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10732) );
  AOI22_X1 U13736 ( .A1(n11248), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10731) );
  INV_X1 U13737 ( .A(n10735), .ZN(n10737) );
  NAND2_X1 U13738 ( .A1(n10737), .A2(n10736), .ZN(n10738) );
  AND2_X1 U13739 ( .A1(n19873), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10739) );
  INV_X1 U13740 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16297) );
  NAND2_X1 U13741 ( .A1(n11272), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13742 ( .A1(n11361), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10743) );
  INV_X1 U13743 ( .A(n13296), .ZN(n10747) );
  NAND2_X2 U13744 ( .A1(n10747), .A2(n15517), .ZN(n10772) );
  INV_X1 U13745 ( .A(n10749), .ZN(n10753) );
  OR2_X1 U13746 ( .A1(n10751), .A2(n10750), .ZN(n10752) );
  INV_X1 U13747 ( .A(n19170), .ZN(n13021) );
  INV_X1 U13748 ( .A(n10763), .ZN(n10771) );
  OR2_X2 U13749 ( .A1(n10772), .A2(n10771), .ZN(n19409) );
  NOR2_X2 U13750 ( .A1(n10772), .A2(n10760), .ZN(n19338) );
  INV_X1 U13751 ( .A(n10754), .ZN(n10767) );
  NAND2_X2 U13752 ( .A1(n13296), .A2(n15517), .ZN(n10768) );
  INV_X1 U13753 ( .A(n10756), .ZN(n10755) );
  NAND2_X1 U13754 ( .A1(n19170), .A2(n10756), .ZN(n10776) );
  NAND2_X2 U13755 ( .A1(n10747), .A2(n13678), .ZN(n10779) );
  NOR2_X2 U13756 ( .A1(n10779), .A2(n10760), .ZN(n19203) );
  AOI22_X1 U13757 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19203), .B1(
        n19590), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U13758 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19472), .B1(
        n19528), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10764) );
  INV_X1 U13759 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n19633) );
  OR2_X2 U13760 ( .A1(n10768), .A2(n10776), .ZN(n13574) );
  INV_X1 U13761 ( .A(n10768), .ZN(n10769) );
  NAND2_X2 U13762 ( .A1(n10763), .A2(n10769), .ZN(n19653) );
  INV_X1 U13763 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11515) );
  OAI22_X1 U13764 ( .A1(n19633), .A2(n13574), .B1(n19653), .B2(n11515), .ZN(
        n10770) );
  INV_X1 U13765 ( .A(n10770), .ZN(n10785) );
  INV_X1 U13766 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10774) );
  INV_X1 U13767 ( .A(n10780), .ZN(n10778) );
  OR2_X2 U13768 ( .A1(n10772), .A2(n10778), .ZN(n10951) );
  INV_X1 U13769 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10773) );
  OAI22_X1 U13770 ( .A1(n10774), .A2(n10941), .B1(n10951), .B2(n10773), .ZN(
        n10775) );
  INV_X1 U13771 ( .A(n10775), .ZN(n10784) );
  INV_X1 U13772 ( .A(n10776), .ZN(n10777) );
  INV_X1 U13773 ( .A(n10994), .ZN(n19502) );
  AOI22_X1 U13774 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19249), .B1(
        n19502), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13775 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19313), .B1(
        n19559), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10782) );
  OR2_X1 U13776 ( .A1(n9762), .A2(n13326), .ZN(n11530) );
  INV_X2 U13777 ( .A(n11530), .ZN(n14144) );
  AOI22_X1 U13778 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n14144), .B1(
        n14136), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10800) );
  OR2_X2 U13779 ( .A1(n14274), .A2(n13326), .ZN(n14099) );
  NAND2_X1 U13780 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10791) );
  NAND2_X1 U13781 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10790) );
  OAI211_X1 U13782 ( .C1(n14099), .C2(n19633), .A(n10791), .B(n10790), .ZN(
        n10792) );
  INV_X1 U13783 ( .A(n10792), .ZN(n10799) );
  INV_X2 U13784 ( .A(n14141), .ZN(n14096) );
  INV_X1 U13785 ( .A(n10793), .ZN(n10794) );
  INV_X4 U13786 ( .A(n10794), .ZN(n14302) );
  AND2_X2 U13787 ( .A1(n14302), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10884) );
  AOI22_X1 U13788 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10798) );
  AND2_X2 U13789 ( .A1(n10796), .A2(n13326), .ZN(n14145) );
  AND2_X1 U13790 ( .A1(n14166), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10965) );
  AOI22_X1 U13791 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14145), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10797) );
  NAND4_X1 U13792 ( .A1(n10800), .A2(n10799), .A3(n10798), .A4(n10797), .ZN(
        n10810) );
  AND2_X2 U13793 ( .A1(n9717), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14077) );
  AOI22_X1 U13794 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14150), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10808) );
  AND2_X2 U13795 ( .A1(n14315), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10833) );
  AOI22_X1 U13796 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10833), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10807) );
  AND2_X1 U13797 ( .A1(n10802), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10803) );
  AND2_X2 U13798 ( .A1(n14115), .A2(n10803), .ZN(n14154) );
  AND2_X1 U13799 ( .A1(n15505), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10804) );
  AOI22_X1 U13800 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10806) );
  AND2_X2 U13801 ( .A1(n9763), .A2(n13326), .ZN(n14152) );
  NAND2_X1 U13802 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n10805) );
  NAND4_X1 U13803 ( .A1(n10808), .A2(n10807), .A3(n10806), .A4(n10805), .ZN(
        n10809) );
  INV_X1 U13804 ( .A(n11430), .ZN(n10811) );
  INV_X1 U13805 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10814) );
  INV_X1 U13806 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10813) );
  OAI22_X1 U13807 ( .A1(n10946), .A2(n10814), .B1(n10941), .B2(n10813), .ZN(
        n10817) );
  INV_X1 U13808 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14168) );
  INV_X1 U13809 ( .A(n19249), .ZN(n10939) );
  INV_X1 U13810 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10815) );
  OAI22_X1 U13811 ( .A1(n14168), .A2(n10951), .B1(n10939), .B2(n10815), .ZN(
        n10816) );
  NOR2_X1 U13812 ( .A1(n10817), .A2(n10816), .ZN(n10832) );
  INV_X1 U13813 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10819) );
  NAND2_X1 U13814 ( .A1(n19338), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10818) );
  OAI211_X1 U13815 ( .C1(n10819), .C2(n10950), .A(n10818), .B(n10757), .ZN(
        n10822) );
  INV_X1 U13816 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11471) );
  INV_X1 U13817 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14175) );
  NOR2_X1 U13818 ( .A1(n10822), .A2(n10821), .ZN(n10831) );
  INV_X1 U13819 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13072) );
  INV_X1 U13820 ( .A(n19203), .ZN(n10954) );
  INV_X1 U13821 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11475) );
  OAI22_X1 U13822 ( .A1(n13072), .A2(n10954), .B1(n19653), .B2(n11475), .ZN(
        n10825) );
  INV_X1 U13823 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10846) );
  INV_X1 U13824 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10823) );
  OAI22_X1 U13825 ( .A1(n10846), .A2(n13574), .B1(n10994), .B2(n10823), .ZN(
        n10824) );
  NOR2_X1 U13826 ( .A1(n10825), .A2(n10824), .ZN(n10830) );
  INV_X1 U13827 ( .A(n10826), .ZN(n10827) );
  NOR2_X1 U13828 ( .A1(n10828), .A2(n10827), .ZN(n10829) );
  AOI22_X1 U13829 ( .A1(n14135), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14144), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10837) );
  AOI22_X1 U13830 ( .A1(n14145), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10833), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13831 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13832 ( .A1(n14136), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10834) );
  NAND4_X1 U13833 ( .A1(n10837), .A2(n10836), .A3(n10835), .A4(n10834), .ZN(
        n10843) );
  AOI22_X1 U13834 ( .A1(n14153), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14137), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13835 ( .A1(n14154), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14138), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13836 ( .A1(n10965), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13837 ( .A1(n10884), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10838) );
  NAND4_X1 U13838 ( .A1(n10841), .A2(n10840), .A3(n10839), .A4(n10838), .ZN(
        n10842) );
  NOR2_X1 U13839 ( .A1(n10843), .A2(n10842), .ZN(n11666) );
  OR2_X1 U13840 ( .A1(n11666), .A2(n10757), .ZN(n16304) );
  INV_X1 U13841 ( .A(n16304), .ZN(n10858) );
  AOI22_X1 U13842 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14096), .B1(
        n14136), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10851) );
  NAND2_X1 U13843 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10845) );
  NAND2_X1 U13844 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10844) );
  OAI211_X1 U13845 ( .C1(n14099), .C2(n10846), .A(n10845), .B(n10844), .ZN(
        n10847) );
  INV_X1 U13846 ( .A(n10847), .ZN(n10850) );
  AOI22_X1 U13847 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U13848 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14145), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10848) );
  NAND4_X1 U13849 ( .A1(n10851), .A2(n10850), .A3(n10849), .A4(n10848), .ZN(
        n10857) );
  AOI22_X1 U13850 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n14150), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10855) );
  AOI22_X1 U13851 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n14152), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10854) );
  AOI22_X1 U13852 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10853) );
  NAND2_X1 U13853 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10852) );
  NAND4_X1 U13854 ( .A1(n10855), .A2(n10854), .A3(n10853), .A4(n10852), .ZN(
        n10856) );
  NAND2_X1 U13855 ( .A1(n10858), .A2(n11665), .ZN(n11671) );
  AOI22_X1 U13856 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n14150), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13857 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n14152), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U13858 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10860) );
  NAND2_X1 U13859 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10859) );
  AOI22_X1 U13860 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14137), .B1(
        n14138), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10866) );
  NAND2_X1 U13861 ( .A1(n14135), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10865) );
  NAND2_X1 U13862 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10864) );
  NAND2_X1 U13863 ( .A1(n14136), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10863) );
  NAND4_X1 U13864 ( .A1(n10866), .A2(n10865), .A3(n10864), .A4(n10863), .ZN(
        n10871) );
  NAND2_X1 U13865 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10870) );
  NAND2_X1 U13866 ( .A1(n10884), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10869) );
  NAND2_X1 U13867 ( .A1(n14145), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10868) );
  NAND2_X1 U13868 ( .A1(n10965), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10867) );
  NAND2_X1 U13869 ( .A1(n11671), .A2(n11672), .ZN(n10872) );
  NAND2_X1 U13870 ( .A1(n10874), .A2(n10873), .ZN(n10875) );
  AOI22_X1 U13871 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n14150), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U13872 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n14152), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13873 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n14153), .B1(
        n14138), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10877) );
  NAND2_X1 U13874 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10876) );
  AOI22_X1 U13875 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14137), .B1(
        n14154), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10883) );
  NAND2_X1 U13876 ( .A1(n14135), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10882) );
  NAND2_X1 U13877 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10881) );
  NAND2_X1 U13878 ( .A1(n14136), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10880) );
  NAND4_X1 U13879 ( .A1(n10883), .A2(n10882), .A3(n10881), .A4(n10880), .ZN(
        n10890) );
  NAND2_X1 U13880 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10888) );
  NAND2_X1 U13881 ( .A1(n14145), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10887) );
  NAND2_X1 U13882 ( .A1(n14143), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10886) );
  NAND2_X1 U13883 ( .A1(n10884), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10885) );
  NAND4_X1 U13884 ( .A1(n10888), .A2(n10887), .A3(n10886), .A4(n10885), .ZN(
        n10889) );
  AND2_X4 U13885 ( .A1(n10892), .A2(n10891), .ZN(n14045) );
  MUX2_X1 U13886 ( .A(n10893), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11172) );
  NAND2_X1 U13887 ( .A1(n11172), .A2(n11184), .ZN(n10895) );
  NAND2_X1 U13888 ( .A1(n10893), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10894) );
  NAND2_X1 U13889 ( .A1(n10895), .A2(n10894), .ZN(n10900) );
  XNOR2_X1 U13890 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10899) );
  NAND2_X1 U13891 ( .A1(n10900), .A2(n10899), .ZN(n10897) );
  NAND2_X1 U13892 ( .A1(n19845), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10896) );
  NAND2_X1 U13893 ( .A1(n10897), .A2(n10896), .ZN(n10933) );
  MUX2_X1 U13894 ( .A(n13299), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10932) );
  INV_X1 U13895 ( .A(n10932), .ZN(n10898) );
  XNOR2_X1 U13896 ( .A(n10933), .B(n10898), .ZN(n11209) );
  MUX2_X1 U13897 ( .A(n11430), .B(n11209), .S(n12907), .Z(n11176) );
  INV_X1 U13898 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13662) );
  MUX2_X1 U13899 ( .A(n11176), .B(n13662), .S(n9755), .Z(n10904) );
  XNOR2_X1 U13900 ( .A(n10900), .B(n10899), .ZN(n11218) );
  INV_X1 U13901 ( .A(n11218), .ZN(n11188) );
  NAND2_X1 U13902 ( .A1(n12907), .A2(n11188), .ZN(n11221) );
  INV_X1 U13903 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10901) );
  NOR2_X1 U13904 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10902) );
  MUX2_X1 U13905 ( .A(n11665), .B(n10902), .S(n9755), .Z(n10907) );
  OAI21_X1 U13906 ( .B1(n10904), .B2(n10903), .A(n10985), .ZN(n13666) );
  INV_X1 U13907 ( .A(n11184), .ZN(n10906) );
  NAND2_X1 U13908 ( .A1(n10802), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10905) );
  AND2_X1 U13909 ( .A1(n10906), .A2(n10905), .ZN(n11213) );
  INV_X1 U13910 ( .A(n11213), .ZN(n11216) );
  MUX2_X1 U13911 ( .A(n11216), .B(n11666), .S(n10702), .Z(n11175) );
  INV_X1 U13912 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13020) );
  MUX2_X1 U13913 ( .A(n11175), .B(n13020), .S(n9755), .Z(n19068) );
  INV_X1 U13914 ( .A(n10907), .ZN(n10910) );
  NAND3_X1 U13915 ( .A1(n9755), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10908) );
  NAND2_X1 U13916 ( .A1(n10910), .A2(n10908), .ZN(n13693) );
  NOR2_X1 U13917 ( .A1(n10225), .A2(n13693), .ZN(n10909) );
  NAND2_X1 U13918 ( .A1(n10225), .A2(n13693), .ZN(n13007) );
  OAI21_X1 U13919 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10909), .A(
        n13007), .ZN(n13996) );
  XNOR2_X1 U13920 ( .A(n10911), .B(n10910), .ZN(n13674) );
  XNOR2_X1 U13921 ( .A(n13674), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13995) );
  OR2_X1 U13922 ( .A1(n13996), .A2(n13995), .ZN(n14003) );
  NAND2_X1 U13923 ( .A1(n13674), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10912) );
  NAND2_X1 U13924 ( .A1(n14003), .A2(n10912), .ZN(n13601) );
  NAND2_X1 U13925 ( .A1(n13600), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10913) );
  INV_X1 U13926 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10915) );
  INV_X1 U13927 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10914) );
  OAI22_X1 U13928 ( .A1(n10915), .A2(n14099), .B1(n11530), .B2(n10914), .ZN(
        n10916) );
  INV_X1 U13929 ( .A(n10916), .ZN(n10924) );
  AOI22_X1 U13930 ( .A1(n14136), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U13931 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10884), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10922) );
  INV_X1 U13932 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10919) );
  NAND2_X1 U13933 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10918) );
  NAND2_X1 U13934 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10917) );
  OAI211_X1 U13935 ( .C1(n14141), .C2(n10919), .A(n10918), .B(n10917), .ZN(
        n10920) );
  INV_X1 U13936 ( .A(n10920), .ZN(n10921) );
  NAND4_X1 U13937 ( .A1(n10924), .A2(n10923), .A3(n10922), .A4(n10921), .ZN(
        n10930) );
  AOI22_X1 U13938 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n14143), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U13939 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10833), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U13940 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10926) );
  NAND2_X1 U13941 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10925) );
  NAND4_X1 U13942 ( .A1(n10928), .A2(n10927), .A3(n10926), .A4(n10925), .ZN(
        n10929) );
  NOR2_X1 U13943 ( .A1(n13326), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10931) );
  AOI21_X1 U13944 ( .B1(n10933), .B2(n10932), .A(n10931), .ZN(n11179) );
  NOR2_X1 U13945 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20834), .ZN(
        n10934) );
  NAND2_X1 U13946 ( .A1(n11179), .A2(n10934), .ZN(n11183) );
  MUX2_X1 U13947 ( .A(n11435), .B(n11183), .S(n12907), .Z(n11210) );
  INV_X1 U13948 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13392) );
  MUX2_X1 U13949 ( .A(n11210), .B(n13392), .S(n9755), .Z(n10935) );
  XNOR2_X1 U13950 ( .A(n10985), .B(n10984), .ZN(n10936) );
  XNOR2_X1 U13951 ( .A(n10936), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19155) );
  NAND2_X1 U13952 ( .A1(n19157), .A2(n19155), .ZN(n10938) );
  INV_X1 U13953 ( .A(n10936), .ZN(n19040) );
  NAND2_X1 U13954 ( .A1(n19040), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10937) );
  INV_X1 U13955 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14078) );
  INV_X1 U13956 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10940) );
  OAI22_X1 U13957 ( .A1(n14078), .A2(n10939), .B1(n10994), .B2(n10940), .ZN(
        n10944) );
  INV_X1 U13958 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10942) );
  INV_X1 U13959 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11555) );
  OAI22_X1 U13960 ( .A1(n10942), .A2(n10941), .B1(n19653), .B2(n11555), .ZN(
        n10943) );
  NOR2_X1 U13961 ( .A1(n10944), .A2(n10943), .ZN(n10961) );
  INV_X1 U13962 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14088) );
  INV_X1 U13963 ( .A(n19528), .ZN(n11005) );
  INV_X1 U13964 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10945) );
  OAI22_X1 U13965 ( .A1(n14088), .A2(n19593), .B1(n11005), .B2(n10945), .ZN(
        n10949) );
  INV_X1 U13966 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10947) );
  INV_X1 U13967 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14266) );
  OAI22_X1 U13968 ( .A1(n10947), .A2(n10946), .B1(n11008), .B2(n14266), .ZN(
        n10948) );
  NOR2_X1 U13969 ( .A1(n10949), .A2(n10948), .ZN(n10960) );
  INV_X1 U13970 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14086) );
  INV_X1 U13971 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11551) );
  OAI22_X1 U13972 ( .A1(n14086), .A2(n10950), .B1(n10995), .B2(n11551), .ZN(
        n10953) );
  INV_X1 U13973 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14259) );
  INV_X1 U13974 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14081) );
  OAI22_X1 U13975 ( .A1(n14259), .A2(n10951), .B1(n13574), .B2(n14081), .ZN(
        n10952) );
  NOR2_X1 U13976 ( .A1(n10953), .A2(n10952), .ZN(n10959) );
  INV_X1 U13977 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14084) );
  INV_X1 U13978 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13452) );
  INV_X1 U13979 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10955) );
  OAI22_X1 U13980 ( .A1(n13452), .A2(n10954), .B1(n19469), .B2(n10955), .ZN(
        n10956) );
  NOR2_X1 U13981 ( .A1(n10957), .A2(n10956), .ZN(n10958) );
  NAND4_X1 U13982 ( .A1(n10961), .A2(n10960), .A3(n10959), .A4(n10958), .ZN(
        n10979) );
  AOI22_X1 U13983 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14136), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10969) );
  NAND2_X1 U13984 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10963) );
  NAND2_X1 U13985 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10962) );
  OAI211_X1 U13986 ( .C1(n14099), .C2(n14081), .A(n10963), .B(n10962), .ZN(
        n10964) );
  INV_X1 U13987 ( .A(n10964), .ZN(n10968) );
  AOI22_X1 U13988 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U13989 ( .A1(n14143), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10966) );
  NAND4_X1 U13990 ( .A1(n10969), .A2(n10968), .A3(n10967), .A4(n10966), .ZN(
        n10976) );
  AOI22_X1 U13991 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U13992 ( .A1(n10970), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10973) );
  AOI22_X1 U13993 ( .A1(n14154), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10972) );
  NAND2_X1 U13994 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10971) );
  NAND4_X1 U13995 ( .A1(n10974), .A2(n10973), .A3(n10972), .A4(n10971), .ZN(
        n10975) );
  INV_X1 U13996 ( .A(n11440), .ZN(n10977) );
  NAND2_X1 U13997 ( .A1(n10977), .A2(n14257), .ZN(n10978) );
  NAND2_X1 U13998 ( .A1(n10981), .A2(n10980), .ZN(n11664) );
  NAND3_X1 U13999 ( .A1(n11664), .A2(n11663), .A3(n14045), .ZN(n10990) );
  NOR2_X2 U14000 ( .A1(n10985), .A2(n10984), .ZN(n10987) );
  INV_X1 U14001 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13419) );
  MUX2_X1 U14002 ( .A(n11440), .B(n13419), .S(n9755), .Z(n10986) );
  INV_X1 U14003 ( .A(n11036), .ZN(n10989) );
  OR2_X1 U14004 ( .A1(n10987), .A2(n10986), .ZN(n10988) );
  NAND2_X1 U14005 ( .A1(n10989), .A2(n10988), .ZN(n19027) );
  NAND2_X1 U14006 ( .A1(n10990), .A2(n19027), .ZN(n10991) );
  INV_X1 U14007 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13781) );
  XNOR2_X1 U14008 ( .A(n10991), .B(n13781), .ZN(n13773) );
  NAND2_X1 U14009 ( .A1(n13772), .A2(n13773), .ZN(n10993) );
  INV_X1 U14010 ( .A(n10991), .ZN(n10992) );
  INV_X1 U14011 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14110) );
  INV_X1 U14012 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11018) );
  OAI22_X1 U14013 ( .A1(n14110), .A2(n10939), .B1(n10994), .B2(n11018), .ZN(
        n10998) );
  INV_X1 U14014 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10996) );
  INV_X1 U14015 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11574) );
  OAI22_X1 U14016 ( .A1(n10996), .A2(n10950), .B1(n10995), .B2(n11574), .ZN(
        n10997) );
  NOR2_X1 U14017 ( .A1(n10998), .A2(n10997), .ZN(n11015) );
  INV_X1 U14018 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10999) );
  INV_X1 U14019 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14286) );
  OAI22_X1 U14020 ( .A1(n10999), .A2(n10941), .B1(n10951), .B2(n14286), .ZN(
        n11001) );
  INV_X1 U14021 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14106) );
  INV_X1 U14022 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11569) );
  OAI22_X1 U14023 ( .A1(n14106), .A2(n13574), .B1(n19653), .B2(n11569), .ZN(
        n11000) );
  NOR2_X1 U14024 ( .A1(n11001), .A2(n11000), .ZN(n11014) );
  INV_X1 U14025 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11003) );
  INV_X1 U14026 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11002) );
  OAI22_X1 U14027 ( .A1(n11003), .A2(n10954), .B1(n19593), .B2(n11002), .ZN(
        n11007) );
  INV_X1 U14028 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14107) );
  INV_X1 U14029 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11004) );
  OAI22_X1 U14030 ( .A1(n14107), .A2(n11005), .B1(n19469), .B2(n11004), .ZN(
        n11006) );
  NOR2_X1 U14031 ( .A1(n11007), .A2(n11006), .ZN(n11013) );
  INV_X1 U14032 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11570) );
  INV_X1 U14033 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11009) );
  INV_X1 U14034 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14279) );
  OAI22_X1 U14035 ( .A1(n11009), .A2(n10946), .B1(n11008), .B2(n14279), .ZN(
        n11010) );
  NOR2_X1 U14036 ( .A1(n11011), .A2(n11010), .ZN(n11012) );
  NAND4_X1 U14037 ( .A1(n11015), .A2(n11014), .A3(n11013), .A4(n11012), .ZN(
        n11032) );
  AOI22_X1 U14038 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n14135), .B1(
        n14136), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11023) );
  NAND2_X1 U14039 ( .A1(n14154), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11017) );
  NAND2_X1 U14040 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11016) );
  OAI211_X1 U14041 ( .C1(n11530), .C2(n11018), .A(n11017), .B(n11016), .ZN(
        n11019) );
  INV_X1 U14042 ( .A(n11019), .ZN(n11022) );
  AOI22_X1 U14043 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U14044 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10884), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11020) );
  NAND4_X1 U14045 ( .A1(n11023), .A2(n11022), .A3(n11021), .A4(n11020), .ZN(
        n11029) );
  AOI22_X1 U14046 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n14145), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U14047 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n14155), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U14048 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14153), .B1(
        n14138), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11025) );
  NAND2_X1 U14049 ( .A1(n14152), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11024) );
  NAND4_X1 U14050 ( .A1(n11027), .A2(n11026), .A3(n11025), .A4(n11024), .ZN(
        n11028) );
  INV_X1 U14051 ( .A(n11443), .ZN(n11030) );
  NAND2_X1 U14052 ( .A1(n11030), .A2(n14257), .ZN(n11031) );
  INV_X1 U14053 ( .A(n11686), .ZN(n11033) );
  INV_X1 U14054 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13461) );
  MUX2_X1 U14055 ( .A(n11443), .B(n13461), .S(n9755), .Z(n11035) );
  OAI21_X1 U14056 ( .B1(n11036), .B2(n11035), .A(n11042), .ZN(n19015) );
  INV_X1 U14057 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15483) );
  NAND2_X1 U14058 ( .A1(n11038), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11039) );
  MUX2_X1 U14059 ( .A(n14045), .B(P2_EBX_REG_7__SCAN_IN), .S(n9755), .Z(n11041) );
  AND2_X1 U14060 ( .A1(n9755), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11040) );
  XNOR2_X1 U14061 ( .A(n11047), .B(n11040), .ZN(n19007) );
  INV_X1 U14062 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16285) );
  NOR2_X1 U14063 ( .A1(n14045), .A2(n16285), .ZN(n11699) );
  NAND2_X1 U14064 ( .A1(n19007), .A2(n11699), .ZN(n16186) );
  XNOR2_X1 U14065 ( .A(n11042), .B(n10052), .ZN(n13685) );
  NAND2_X1 U14066 ( .A1(n13685), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16188) );
  NAND2_X1 U14067 ( .A1(n19007), .A2(n11694), .ZN(n11043) );
  NAND2_X1 U14068 ( .A1(n11043), .A2(n16285), .ZN(n16187) );
  INV_X1 U14069 ( .A(n13685), .ZN(n11044) );
  INV_X1 U14070 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11696) );
  NAND2_X1 U14071 ( .A1(n11044), .A2(n11696), .ZN(n16190) );
  AND2_X1 U14072 ( .A1(n16187), .A2(n16190), .ZN(n11045) );
  INV_X1 U14073 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13491) );
  NAND2_X1 U14074 ( .A1(n11047), .A2(n13491), .ZN(n11048) );
  AND2_X1 U14075 ( .A1(n9755), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11049) );
  XNOR2_X1 U14076 ( .A(n11050), .B(n11049), .ZN(n18996) );
  NAND2_X1 U14077 ( .A1(n18996), .A2(n11694), .ZN(n11060) );
  INV_X1 U14078 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15470) );
  NAND2_X1 U14079 ( .A1(n9755), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11051) );
  INV_X1 U14080 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13495) );
  MUX2_X1 U14081 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n11051), .S(n11053), .Z(
        n11052) );
  NAND2_X1 U14082 ( .A1(n11052), .A2(n11145), .ZN(n18982) );
  OR2_X1 U14083 ( .A1(n18982), .A2(n14045), .ZN(n11061) );
  INV_X1 U14084 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16153) );
  NAND2_X1 U14085 ( .A1(n11061), .A2(n16153), .ZN(n15447) );
  NOR2_X2 U14086 ( .A1(n11053), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11055) );
  NAND2_X1 U14087 ( .A1(n9755), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11054) );
  OR2_X1 U14088 ( .A1(n11055), .A2(n11054), .ZN(n11057) );
  INV_X1 U14089 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13521) );
  INV_X1 U14090 ( .A(n11062), .ZN(n11056) );
  NAND2_X1 U14091 ( .A1(n11057), .A2(n11056), .ZN(n18970) );
  OR2_X1 U14092 ( .A1(n18970), .A2(n14045), .ZN(n11067) );
  INV_X1 U14093 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16152) );
  INV_X1 U14094 ( .A(n16162), .ZN(n11058) );
  NOR2_X1 U14095 ( .A1(n11060), .A2(n15470), .ZN(n15462) );
  NOR2_X1 U14096 ( .A1(n16153), .A2(n11061), .ZN(n15445) );
  NOR2_X1 U14097 ( .A1(n15462), .A2(n15445), .ZN(n16159) );
  NAND2_X1 U14098 ( .A1(n9755), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11063) );
  INV_X1 U14099 ( .A(n11063), .ZN(n11065) );
  NAND2_X1 U14100 ( .A1(n11065), .A2(n11064), .ZN(n11066) );
  NAND2_X1 U14101 ( .A1(n11089), .A2(n11066), .ZN(n18957) );
  INV_X1 U14102 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15425) );
  OR3_X1 U14103 ( .A1(n18957), .A2(n14045), .A3(n15425), .ZN(n15416) );
  OR2_X1 U14104 ( .A1(n11067), .A2(n16152), .ZN(n16161) );
  AND2_X1 U14105 ( .A1(n9755), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11087) );
  INV_X1 U14106 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n11294) );
  INV_X1 U14107 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13733) );
  NAND2_X1 U14108 ( .A1(n11294), .A2(n13733), .ZN(n11068) );
  INV_X1 U14109 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n15041) );
  INV_X1 U14110 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11069) );
  NAND2_X1 U14111 ( .A1(n15041), .A2(n11069), .ZN(n11070) );
  AND2_X1 U14112 ( .A1(n9755), .A2(n11070), .ZN(n11071) );
  NAND2_X1 U14113 ( .A1(n9755), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11105) );
  AND2_X1 U14114 ( .A1(n9755), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11102) );
  OR2_X2 U14115 ( .A1(n11104), .A2(n11102), .ZN(n11098) );
  OR2_X2 U14116 ( .A1(n11098), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11123) );
  NAND2_X1 U14117 ( .A1(n11123), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11072) );
  OAI21_X1 U14118 ( .B1(n11072), .B2(n11034), .A(n11145), .ZN(n11073) );
  INV_X1 U14119 ( .A(n11073), .ZN(n11074) );
  OAI21_X1 U14120 ( .B1(n11123), .B2(P2_EBX_REG_21__SCAN_IN), .A(n11074), .ZN(
        n14927) );
  OR2_X1 U14121 ( .A1(n14927), .A2(n14045), .ZN(n11075) );
  INV_X1 U14122 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15181) );
  NAND2_X1 U14123 ( .A1(n11075), .A2(n15181), .ZN(n15170) );
  INV_X1 U14124 ( .A(n11076), .ZN(n11106) );
  OR2_X1 U14125 ( .A1(n11092), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11094) );
  NAND3_X1 U14126 ( .A1(n11094), .A2(P2_EBX_REG_17__SCAN_IN), .A3(n9755), .ZN(
        n11077) );
  NAND2_X1 U14127 ( .A1(n11106), .A2(n11077), .ZN(n18925) );
  INV_X1 U14128 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11397) );
  OAI21_X1 U14129 ( .B1(n18925), .B2(n14045), .A(n11397), .ZN(n15176) );
  OR2_X1 U14130 ( .A1(n11083), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11084) );
  AND2_X1 U14131 ( .A1(n9755), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11078) );
  NAND2_X1 U14132 ( .A1(n11084), .A2(n11078), .ZN(n11079) );
  NAND2_X1 U14133 ( .A1(n11079), .A2(n11092), .ZN(n12910) );
  OR2_X1 U14134 ( .A1(n12910), .A2(n14045), .ZN(n11080) );
  INV_X1 U14135 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15237) );
  NAND2_X1 U14136 ( .A1(n11080), .A2(n15237), .ZN(n16119) );
  OR2_X1 U14137 ( .A1(n18957), .A2(n14045), .ZN(n11081) );
  NAND2_X1 U14138 ( .A1(n11081), .A2(n15425), .ZN(n15417) );
  AND2_X1 U14139 ( .A1(n16119), .A2(n15417), .ZN(n11091) );
  NAND2_X1 U14140 ( .A1(n11083), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11082) );
  MUX2_X1 U14141 ( .A(n11083), .B(n11082), .S(n9755), .Z(n11085) );
  NAND2_X1 U14142 ( .A1(n18949), .A2(n11694), .ZN(n11086) );
  INV_X1 U14143 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16251) );
  NAND2_X1 U14144 ( .A1(n11086), .A2(n16251), .ZN(n16131) );
  INV_X1 U14145 ( .A(n11087), .ZN(n11088) );
  XNOR2_X1 U14146 ( .A(n11089), .B(n11088), .ZN(n13715) );
  NAND2_X1 U14147 ( .A1(n13715), .A2(n11694), .ZN(n11090) );
  INV_X1 U14148 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15426) );
  NAND2_X1 U14149 ( .A1(n11090), .A2(n15426), .ZN(n15419) );
  AND4_X1 U14150 ( .A1(n15176), .A2(n11091), .A3(n16131), .A4(n15419), .ZN(
        n11101) );
  NAND3_X1 U14151 ( .A1(n11092), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n9755), .ZN(
        n11093) );
  AND3_X1 U14152 ( .A1(n11094), .A2(n11145), .A3(n11093), .ZN(n18937) );
  NAND2_X1 U14153 ( .A1(n18937), .A2(n11694), .ZN(n11095) );
  XNOR2_X1 U14154 ( .A(n11095), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15171) );
  AND2_X1 U14155 ( .A1(n9755), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11097) );
  INV_X1 U14156 ( .A(n11145), .ZN(n11096) );
  AOI21_X1 U14157 ( .B1(n11098), .B2(n11097), .A(n11096), .ZN(n11099) );
  AND2_X1 U14158 ( .A1(n11123), .A2(n11099), .ZN(n14944) );
  NAND2_X1 U14159 ( .A1(n14944), .A2(n11694), .ZN(n11100) );
  INV_X1 U14160 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15196) );
  NAND2_X1 U14161 ( .A1(n11100), .A2(n15196), .ZN(n15189) );
  NAND4_X1 U14162 ( .A1(n15170), .A2(n11101), .A3(n15171), .A4(n15189), .ZN(
        n11108) );
  INV_X1 U14163 ( .A(n11102), .ZN(n11103) );
  XNOR2_X1 U14164 ( .A(n11104), .B(n11103), .ZN(n18900) );
  NAND2_X1 U14165 ( .A1(n18900), .A2(n11694), .ZN(n11120) );
  INV_X1 U14166 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11308) );
  NAND2_X1 U14167 ( .A1(n11120), .A2(n11308), .ZN(n15203) );
  XNOR2_X1 U14168 ( .A(n11106), .B(n11105), .ZN(n18912) );
  NAND2_X1 U14169 ( .A1(n18912), .A2(n11694), .ZN(n11107) );
  INV_X1 U14170 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21055) );
  NAND2_X1 U14171 ( .A1(n11107), .A2(n21055), .ZN(n15215) );
  NAND2_X1 U14172 ( .A1(n15203), .A2(n15215), .ZN(n15190) );
  NOR2_X1 U14173 ( .A1(n11108), .A2(n15190), .ZN(n11109) );
  OR2_X1 U14174 ( .A1(n14045), .A2(n15181), .ZN(n11110) );
  OR2_X1 U14175 ( .A1(n14927), .A2(n11110), .ZN(n15169) );
  NOR2_X1 U14176 ( .A1(n14045), .A2(n16251), .ZN(n11111) );
  NAND2_X1 U14177 ( .A1(n18949), .A2(n11111), .ZN(n16130) );
  OR2_X1 U14178 ( .A1(n14045), .A2(n15237), .ZN(n11112) );
  OR2_X1 U14179 ( .A1(n12910), .A2(n11112), .ZN(n16118) );
  INV_X1 U14180 ( .A(n18925), .ZN(n11114) );
  NOR2_X1 U14181 ( .A1(n14045), .A2(n11397), .ZN(n11113) );
  NAND2_X1 U14182 ( .A1(n11114), .A2(n11113), .ZN(n15175) );
  NOR2_X1 U14183 ( .A1(n14045), .A2(n21055), .ZN(n11115) );
  NAND2_X1 U14184 ( .A1(n18912), .A2(n11115), .ZN(n15214) );
  INV_X1 U14185 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15236) );
  NOR2_X1 U14186 ( .A1(n14045), .A2(n15236), .ZN(n11116) );
  NAND2_X1 U14187 ( .A1(n18937), .A2(n11116), .ZN(n15172) );
  INV_X1 U14188 ( .A(n13715), .ZN(n11117) );
  OR3_X1 U14189 ( .A1(n11117), .A2(n14045), .A3(n15426), .ZN(n15418) );
  AND4_X1 U14190 ( .A1(n15175), .A2(n15214), .A3(n15172), .A4(n15418), .ZN(
        n11119) );
  NOR2_X1 U14191 ( .A1(n14045), .A2(n15196), .ZN(n11118) );
  NAND2_X1 U14192 ( .A1(n14944), .A2(n11118), .ZN(n15188) );
  NAND4_X1 U14193 ( .A1(n15169), .A2(n14025), .A3(n11119), .A4(n15188), .ZN(
        n11122) );
  INV_X1 U14194 ( .A(n11120), .ZN(n11121) );
  INV_X1 U14195 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15013) );
  AND2_X1 U14196 ( .A1(n9755), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11126) );
  INV_X1 U14197 ( .A(n11137), .ZN(n11131) );
  NAND2_X1 U14198 ( .A1(n11126), .A2(n11125), .ZN(n11127) );
  AND2_X1 U14199 ( .A1(n11131), .A2(n11127), .ZN(n15564) );
  NAND2_X1 U14200 ( .A1(n15564), .A2(n11694), .ZN(n11128) );
  INV_X1 U14201 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15165) );
  NAND2_X1 U14202 ( .A1(n11128), .A2(n15165), .ZN(n15158) );
  INV_X1 U14203 ( .A(n11128), .ZN(n11129) );
  NAND2_X1 U14204 ( .A1(n11129), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15159) );
  AND2_X1 U14205 ( .A1(n9755), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11130) );
  XNOR2_X1 U14206 ( .A(n11131), .B(n11130), .ZN(n11132) );
  INV_X1 U14207 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11325) );
  OAI21_X1 U14208 ( .B1(n11132), .B2(n14045), .A(n11325), .ZN(n11134) );
  INV_X1 U14209 ( .A(n11132), .ZN(n16064) );
  AND2_X1 U14210 ( .A1(n11694), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11133) );
  NAND2_X1 U14211 ( .A1(n16064), .A2(n11133), .ZN(n11135) );
  INV_X1 U14212 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n11136) );
  INV_X1 U14213 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11138) );
  INV_X1 U14214 ( .A(n11147), .ZN(n11142) );
  INV_X1 U14215 ( .A(n11139), .ZN(n11140) );
  NAND3_X1 U14216 ( .A1(n11140), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n9755), .ZN(
        n11141) );
  NAND3_X1 U14217 ( .A1(n11142), .A2(n11145), .A3(n11141), .ZN(n14920) );
  NOR2_X1 U14218 ( .A1(n14920), .A2(n14045), .ZN(n15152) );
  INV_X1 U14219 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14984) );
  NAND2_X1 U14220 ( .A1(n9755), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n11143) );
  INV_X1 U14221 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11340) );
  INV_X1 U14222 ( .A(n11153), .ZN(n11168) );
  OAI21_X1 U14223 ( .B1(n11149), .B2(n11143), .A(n11168), .ZN(n16041) );
  NOR2_X1 U14224 ( .A1(n16041), .A2(n14045), .ZN(n11144) );
  INV_X1 U14225 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15317) );
  OAI21_X1 U14226 ( .B1(n11144), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n11156), .ZN(n15139) );
  NAND2_X1 U14227 ( .A1(n9755), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11146) );
  OAI21_X1 U14228 ( .B1(n11147), .B2(n11146), .A(n11145), .ZN(n11148) );
  NOR2_X1 U14229 ( .A1(n11149), .A2(n11148), .ZN(n16057) );
  NAND2_X1 U14230 ( .A1(n16057), .A2(n11694), .ZN(n11154) );
  INV_X1 U14231 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15335) );
  NOR2_X1 U14232 ( .A1(n15139), .A2(n15323), .ZN(n11150) );
  NAND2_X1 U14233 ( .A1(n9755), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11152) );
  NAND2_X1 U14234 ( .A1(n9755), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11157) );
  XNOR2_X1 U14235 ( .A(n14044), .B(n11157), .ZN(n16019) );
  NAND2_X1 U14236 ( .A1(n16019), .A2(n11694), .ZN(n14048) );
  INV_X1 U14237 ( .A(n11154), .ZN(n11155) );
  NAND2_X1 U14238 ( .A1(n11155), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15322) );
  INV_X1 U14239 ( .A(n14044), .ZN(n11158) );
  NAND2_X1 U14240 ( .A1(n11158), .A2(n11157), .ZN(n11159) );
  AND2_X1 U14241 ( .A1(n9755), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11160) );
  XNOR2_X1 U14242 ( .A(n11159), .B(n11160), .ZN(n11165) );
  INV_X1 U14243 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11350) );
  OAI21_X1 U14244 ( .B1(n11165), .B2(n14045), .A(n11350), .ZN(n15118) );
  INV_X1 U14245 ( .A(n11159), .ZN(n11162) );
  INV_X1 U14246 ( .A(n11160), .ZN(n11161) );
  NAND2_X1 U14247 ( .A1(n11162), .A2(n11161), .ZN(n11166) );
  NAND2_X1 U14248 ( .A1(n9755), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11163) );
  XNOR2_X1 U14249 ( .A(n11166), .B(n11163), .ZN(n15996) );
  AOI21_X1 U14250 ( .B1(n15996), .B2(n11694), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15107) );
  INV_X1 U14251 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11659) );
  NOR2_X1 U14252 ( .A1(n14045), .A2(n11659), .ZN(n11164) );
  NAND2_X1 U14253 ( .A1(n15996), .A2(n11164), .ZN(n15108) );
  INV_X1 U14254 ( .A(n11165), .ZN(n16009) );
  NAND3_X1 U14255 ( .A1(n16009), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11694), .ZN(n15117) );
  OAI211_X1 U14256 ( .C1(n15106), .C2(n15107), .A(n15108), .B(n15117), .ZN(
        n11171) );
  NOR2_X1 U14257 ( .A1(n11166), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11167) );
  MUX2_X1 U14258 ( .A(n11168), .B(n11167), .S(n9755), .Z(n15991) );
  NAND2_X1 U14259 ( .A1(n15991), .A2(n11694), .ZN(n11169) );
  XOR2_X1 U14260 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11169), .Z(
        n11170) );
  XNOR2_X1 U14261 ( .A(n11171), .B(n11170), .ZN(n11708) );
  INV_X1 U14262 ( .A(n11172), .ZN(n11217) );
  INV_X1 U14263 ( .A(n11173), .ZN(n11174) );
  OAI21_X1 U14264 ( .B1(n11175), .B2(n11217), .A(n11174), .ZN(n11177) );
  NAND3_X1 U14265 ( .A1(n11177), .A2(n11176), .A3(n11210), .ZN(n11182) );
  NAND2_X1 U14266 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20834), .ZN(
        n11178) );
  NAND2_X1 U14267 ( .A1(n11179), .A2(n11178), .ZN(n11181) );
  NAND2_X1 U14268 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13036), .ZN(
        n11180) );
  INV_X1 U14269 ( .A(n11232), .ZN(n11186) );
  NAND2_X1 U14270 ( .A1(n11182), .A2(n11186), .ZN(n19866) );
  AND2_X1 U14271 ( .A1(n14257), .A2(n19883), .ZN(n19865) );
  INV_X1 U14272 ( .A(n19865), .ZN(n16348) );
  NAND2_X1 U14273 ( .A1(n11183), .A2(n11209), .ZN(n11227) );
  XNOR2_X1 U14274 ( .A(n11217), .B(n11184), .ZN(n11212) );
  NAND2_X1 U14275 ( .A1(n11188), .A2(n11212), .ZN(n11185) );
  OR2_X1 U14276 ( .A1(n11227), .A2(n11185), .ZN(n11187) );
  NAND2_X1 U14277 ( .A1(n11187), .A2(n11186), .ZN(n16313) );
  NAND2_X1 U14278 ( .A1(n11188), .A2(n11213), .ZN(n11190) );
  OAI21_X1 U14279 ( .B1(n11227), .B2(n11190), .A(n11189), .ZN(n11194) );
  NAND2_X1 U14280 ( .A1(n11191), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11192) );
  NAND2_X1 U14281 ( .A1(n11192), .A2(n13036), .ZN(n16321) );
  INV_X1 U14282 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12929) );
  OAI21_X1 U14283 ( .B1(n10970), .B2(n16321), .A(n12929), .ZN(n11193) );
  NAND2_X1 U14284 ( .A1(n11193), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19855) );
  OAI21_X1 U14285 ( .B1(n16313), .B2(n11194), .A(n19855), .ZN(n16344) );
  INV_X1 U14286 ( .A(n16344), .ZN(n19864) );
  OAI22_X1 U14287 ( .A1(n19866), .A2(n16348), .B1(n14257), .B2(n19864), .ZN(
        n11196) );
  INV_X1 U14288 ( .A(n11195), .ZN(n16320) );
  NAND2_X1 U14289 ( .A1(n11196), .A2(n16320), .ZN(n11707) );
  NAND2_X1 U14290 ( .A1(n13033), .A2(n11198), .ZN(n11201) );
  NAND2_X1 U14291 ( .A1(n11199), .A2(n13814), .ZN(n11200) );
  NAND2_X1 U14292 ( .A1(n11200), .A2(n19865), .ZN(n11372) );
  NAND2_X1 U14293 ( .A1(n11201), .A2(n11372), .ZN(n11370) );
  INV_X1 U14294 ( .A(n11370), .ZN(n11205) );
  AND2_X1 U14295 ( .A1(n9726), .A2(n14257), .ZN(n11368) );
  OAI21_X1 U14296 ( .B1(n11368), .B2(n19883), .A(n13814), .ZN(n11202) );
  NAND2_X1 U14297 ( .A1(n11202), .A2(n10689), .ZN(n11204) );
  INV_X1 U14298 ( .A(n16313), .ZN(n12898) );
  NAND2_X1 U14299 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19880) );
  INV_X1 U14300 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21048) );
  INV_X1 U14301 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19745) );
  NOR2_X1 U14302 ( .A1(n21048), .A2(n19745), .ZN(n19755) );
  NOR2_X1 U14303 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n19757) );
  OR3_X1 U14304 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19755), .A3(n19757), .ZN(
        n19881) );
  NOR2_X1 U14305 ( .A1(n19876), .A2(n19881), .ZN(n12927) );
  NAND3_X1 U14306 ( .A1(n10706), .A2(n12898), .A3(n12927), .ZN(n11203) );
  NAND4_X1 U14307 ( .A1(n11206), .A2(n11205), .A3(n11204), .A4(n11203), .ZN(
        n13028) );
  MUX2_X1 U14308 ( .A(n10706), .B(n11380), .S(n14257), .Z(n11207) );
  NOR2_X1 U14309 ( .A1(n16313), .A2(n19876), .ZN(n13026) );
  AND2_X1 U14310 ( .A1(n11207), .A2(n13026), .ZN(n11208) );
  NOR2_X1 U14311 ( .A1(n13028), .A2(n11208), .ZN(n11240) );
  NAND2_X1 U14312 ( .A1(n11210), .A2(n11209), .ZN(n11211) );
  NAND2_X1 U14313 ( .A1(n11211), .A2(n12907), .ZN(n11225) );
  OAI21_X1 U14314 ( .B1(n10757), .B2(n11213), .A(n11212), .ZN(n11214) );
  OAI21_X1 U14315 ( .B1(n10757), .B2(n11218), .A(n11214), .ZN(n11215) );
  NAND2_X1 U14316 ( .A1(n11215), .A2(n9730), .ZN(n11223) );
  OAI21_X1 U14317 ( .B1(n11217), .B2(n11216), .A(n10702), .ZN(n11222) );
  NAND2_X1 U14318 ( .A1(n19883), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11231) );
  NAND2_X1 U14319 ( .A1(n11231), .A2(n10757), .ZN(n11219) );
  NAND2_X1 U14320 ( .A1(n11219), .A2(n11218), .ZN(n11220) );
  AOI22_X1 U14321 ( .A1(n11223), .A2(n11222), .B1(n11221), .B2(n11220), .ZN(
        n11224) );
  AOI21_X1 U14322 ( .B1(n11225), .B2(n11224), .A(n11232), .ZN(n11226) );
  MUX2_X1 U14323 ( .A(n11226), .B(n13036), .S(n19884), .Z(n11230) );
  NAND2_X1 U14324 ( .A1(n11228), .A2(n11227), .ZN(n11229) );
  INV_X1 U14325 ( .A(n13025), .ZN(n11236) );
  AOI21_X1 U14326 ( .B1(n11234), .B2(n9730), .A(n19224), .ZN(n11235) );
  NAND2_X1 U14327 ( .A1(n11236), .A2(n11235), .ZN(n11239) );
  INV_X1 U14328 ( .A(n12927), .ZN(n13023) );
  NOR2_X1 U14329 ( .A1(n10689), .A2(n13023), .ZN(n11237) );
  NAND2_X1 U14330 ( .A1(n13025), .A2(n11237), .ZN(n11238) );
  NAND4_X1 U14331 ( .A1(n11707), .A2(n11240), .A3(n11239), .A4(n11238), .ZN(
        n11241) );
  AND2_X1 U14332 ( .A1(n11189), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16346) );
  NOR2_X1 U14333 ( .A1(n11195), .A2(n12907), .ZN(n11242) );
  NAND2_X1 U14334 ( .A1(n11708), .A2(n19187), .ZN(n11705) );
  AND2_X1 U14335 ( .A1(n11243), .A2(n11704), .ZN(n19192) );
  OR2_X1 U14336 ( .A1(n11355), .A2(n15237), .ZN(n11247) );
  NAND2_X1 U14337 ( .A1(n11362), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14338 ( .A1(n11361), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11244) );
  AND2_X1 U14339 ( .A1(n11245), .A2(n11244), .ZN(n11246) );
  NAND2_X1 U14340 ( .A1(n11247), .A2(n11246), .ZN(n12913) );
  OR2_X1 U14341 ( .A1(n11355), .A2(n15425), .ZN(n11252) );
  NAND2_X1 U14342 ( .A1(n11362), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14343 ( .A1(n11361), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11249) );
  AND2_X1 U14344 ( .A1(n11250), .A2(n11249), .ZN(n11251) );
  OR2_X1 U14345 ( .A1(n11355), .A2(n15470), .ZN(n11256) );
  NAND2_X1 U14346 ( .A1(n11362), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14347 ( .A1(n11361), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11253) );
  AND2_X1 U14348 ( .A1(n11254), .A2(n11253), .ZN(n11255) );
  NAND2_X1 U14349 ( .A1(n11256), .A2(n11255), .ZN(n13493) );
  OR2_X1 U14350 ( .A1(n11355), .A2(n15483), .ZN(n11260) );
  NAND2_X1 U14351 ( .A1(n11362), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14352 ( .A1(n11361), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11257) );
  AND2_X1 U14353 ( .A1(n11258), .A2(n11257), .ZN(n11259) );
  NAND2_X1 U14354 ( .A1(n11262), .A2(n11261), .ZN(n11267) );
  INV_X1 U14355 ( .A(n11263), .ZN(n11265) );
  NAND2_X1 U14356 ( .A1(n11265), .A2(n11264), .ZN(n11266) );
  INV_X1 U14357 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19190) );
  OR2_X1 U14358 ( .A1(n11355), .A2(n19190), .ZN(n11271) );
  NAND2_X1 U14359 ( .A1(n11362), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n11269) );
  AOI22_X1 U14360 ( .A1(n11361), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11268) );
  AND2_X1 U14361 ( .A1(n11269), .A2(n11268), .ZN(n11270) );
  OR2_X1 U14362 ( .A1(n11355), .A2(n13781), .ZN(n11274) );
  AOI22_X1 U14363 ( .A1(n11361), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11273) );
  OAI211_X1 U14364 ( .C1(n13419), .C2(n11341), .A(n11274), .B(n11273), .ZN(
        n13416) );
  OR2_X1 U14365 ( .A1(n11355), .A2(n11696), .ZN(n11278) );
  NAND2_X1 U14366 ( .A1(n11362), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11276) );
  AOI22_X1 U14367 ( .A1(n11361), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11275) );
  AND2_X1 U14368 ( .A1(n11276), .A2(n11275), .ZN(n11277) );
  NAND2_X1 U14369 ( .A1(n11278), .A2(n11277), .ZN(n13448) );
  AOI22_X1 U14370 ( .A1(n11361), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11279) );
  OAI21_X1 U14371 ( .B1(n11341), .B2(n13491), .A(n11279), .ZN(n11280) );
  AOI21_X1 U14372 ( .B1(n10730), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n11280), .ZN(n13488) );
  OR2_X1 U14373 ( .A1(n11355), .A2(n16153), .ZN(n11284) );
  NAND2_X1 U14374 ( .A1(n11362), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14375 ( .A1(n11361), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n11281) );
  AND2_X1 U14376 ( .A1(n11282), .A2(n11281), .ZN(n11283) );
  NAND2_X1 U14377 ( .A1(n11284), .A2(n11283), .ZN(n13532) );
  OR2_X1 U14378 ( .A1(n11355), .A2(n16152), .ZN(n11288) );
  NAND2_X1 U14379 ( .A1(n11362), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14380 ( .A1(n11361), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n11285) );
  AND2_X1 U14381 ( .A1(n11286), .A2(n11285), .ZN(n11287) );
  NAND2_X1 U14382 ( .A1(n11288), .A2(n11287), .ZN(n13520) );
  OR2_X1 U14383 ( .A1(n11355), .A2(n15426), .ZN(n11292) );
  NAND2_X1 U14384 ( .A1(n11362), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14385 ( .A1(n11361), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n11289) );
  AND2_X1 U14386 ( .A1(n11290), .A2(n11289), .ZN(n11291) );
  NAND2_X1 U14387 ( .A1(n11292), .A2(n11291), .ZN(n13559) );
  AOI22_X1 U14388 ( .A1(n11361), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n11293) );
  OAI21_X1 U14389 ( .B1(n11341), .B2(n11294), .A(n11293), .ZN(n11295) );
  AOI21_X1 U14390 ( .B1(n10730), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n11295), .ZN(n13640) );
  OR2_X1 U14391 ( .A1(n11355), .A2(n15236), .ZN(n11299) );
  NAND2_X1 U14392 ( .A1(n11362), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11297) );
  AOI22_X1 U14393 ( .A1(n11361), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11296) );
  AND2_X1 U14394 ( .A1(n11297), .A2(n11296), .ZN(n11298) );
  NAND2_X1 U14395 ( .A1(n11299), .A2(n11298), .ZN(n13763) );
  OR2_X1 U14396 ( .A1(n11355), .A2(n11397), .ZN(n11303) );
  NAND2_X1 U14397 ( .A1(n11362), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14398 ( .A1(n11361), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n11300) );
  AND2_X1 U14399 ( .A1(n11301), .A2(n11300), .ZN(n11302) );
  OR2_X1 U14400 ( .A1(n11355), .A2(n21055), .ZN(n11307) );
  NAND2_X1 U14401 ( .A1(n11362), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U14402 ( .A1(n11361), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n11304) );
  AND2_X1 U14403 ( .A1(n11305), .A2(n11304), .ZN(n11306) );
  NAND2_X1 U14404 ( .A1(n11307), .A2(n11306), .ZN(n15032) );
  OR2_X1 U14405 ( .A1(n11355), .A2(n11308), .ZN(n11312) );
  NAND2_X1 U14406 ( .A1(n11362), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14407 ( .A1(n11361), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11309) );
  AND2_X1 U14408 ( .A1(n11310), .A2(n11309), .ZN(n11311) );
  OR2_X1 U14409 ( .A1(n11355), .A2(n15196), .ZN(n11316) );
  NAND2_X1 U14410 ( .A1(n11362), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14411 ( .A1(n11361), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n11313) );
  AND2_X1 U14412 ( .A1(n11314), .A2(n11313), .ZN(n11315) );
  OR2_X1 U14413 ( .A1(n11355), .A2(n15181), .ZN(n11320) );
  NAND2_X1 U14414 ( .A1(n11362), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11318) );
  AOI22_X1 U14415 ( .A1(n11361), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n11317) );
  AND2_X1 U14416 ( .A1(n11318), .A2(n11317), .ZN(n11319) );
  OR2_X1 U14417 ( .A1(n11355), .A2(n15165), .ZN(n11324) );
  NAND2_X1 U14418 ( .A1(n11362), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11322) );
  AOI22_X1 U14419 ( .A1(n11361), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n11321) );
  AND2_X1 U14420 ( .A1(n11322), .A2(n11321), .ZN(n11323) );
  NAND2_X1 U14421 ( .A1(n11324), .A2(n11323), .ZN(n15002) );
  OR2_X1 U14422 ( .A1(n11355), .A2(n11325), .ZN(n11329) );
  NAND2_X1 U14423 ( .A1(n11362), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11327) );
  AOI22_X1 U14424 ( .A1(n11361), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n11326) );
  AND2_X1 U14425 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  INV_X1 U14426 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16210) );
  OR2_X1 U14427 ( .A1(n11355), .A2(n16210), .ZN(n11333) );
  NAND2_X1 U14428 ( .A1(n11362), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14429 ( .A1(n11361), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n11330) );
  AND2_X1 U14430 ( .A1(n11331), .A2(n11330), .ZN(n11332) );
  OR2_X1 U14431 ( .A1(n11355), .A2(n15335), .ZN(n11337) );
  NAND2_X1 U14432 ( .A1(n11362), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14433 ( .A1(n11361), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n11334) );
  AND2_X1 U14434 ( .A1(n11335), .A2(n11334), .ZN(n11336) );
  NAND2_X1 U14435 ( .A1(n11337), .A2(n11336), .ZN(n14980) );
  OR2_X1 U14436 ( .A1(n11355), .A2(n15317), .ZN(n11339) );
  AOI22_X1 U14437 ( .A1(n11361), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n11338) );
  OAI211_X1 U14438 ( .C1(n11341), .C2(n11340), .A(n11339), .B(n11338), .ZN(
        n14973) );
  INV_X1 U14439 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15301) );
  OR2_X1 U14440 ( .A1(n11355), .A2(n15301), .ZN(n11345) );
  NAND2_X1 U14441 ( .A1(n11362), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14442 ( .A1(n11361), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n11342) );
  AND2_X1 U14443 ( .A1(n11343), .A2(n11342), .ZN(n11344) );
  INV_X1 U14444 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15276) );
  OR2_X1 U14445 ( .A1(n11355), .A2(n15276), .ZN(n11349) );
  NAND2_X1 U14446 ( .A1(n11362), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14447 ( .A1(n11361), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n11346) );
  AND2_X1 U14448 ( .A1(n11347), .A2(n11346), .ZN(n11348) );
  NAND2_X1 U14449 ( .A1(n11349), .A2(n11348), .ZN(n14050) );
  NAND2_X1 U14450 ( .A1(n14051), .A2(n14050), .ZN(n14948) );
  OR2_X1 U14451 ( .A1(n11355), .A2(n11350), .ZN(n11354) );
  NAND2_X1 U14452 ( .A1(n11362), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14453 ( .A1(n11361), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11351) );
  AND2_X1 U14454 ( .A1(n11352), .A2(n11351), .ZN(n11353) );
  AND2_X1 U14455 ( .A1(n11354), .A2(n11353), .ZN(n14947) );
  OR2_X1 U14456 ( .A1(n11355), .A2(n11659), .ZN(n11359) );
  NAND2_X1 U14457 ( .A1(n11362), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14458 ( .A1(n11361), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11356) );
  AND2_X1 U14459 ( .A1(n11357), .A2(n11356), .ZN(n11358) );
  NAND2_X1 U14460 ( .A1(n11359), .A2(n11358), .ZN(n14331) );
  INV_X1 U14461 ( .A(n14331), .ZN(n11360) );
  AOI22_X1 U14462 ( .A1(n11361), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11364) );
  NAND2_X1 U14463 ( .A1(n11362), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n11363) );
  NAND2_X1 U14464 ( .A1(n11364), .A2(n11363), .ZN(n11365) );
  AOI21_X1 U14465 ( .B1(n10730), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n11365), .ZN(n11366) );
  INV_X1 U14466 ( .A(n11715), .ZN(n15993) );
  NAND3_X1 U14467 ( .A1(n10699), .A2(n11368), .A3(n13814), .ZN(n11369) );
  NAND2_X1 U14468 ( .A1(n11704), .A2(n16316), .ZN(n14013) );
  NAND2_X1 U14469 ( .A1(n9735), .A2(n10757), .ZN(n15496) );
  NAND2_X1 U14470 ( .A1(n15496), .A2(n11372), .ZN(n11379) );
  INV_X1 U14471 ( .A(n11373), .ZN(n11375) );
  NAND2_X1 U14472 ( .A1(n11375), .A2(n11374), .ZN(n11377) );
  AOI21_X1 U14473 ( .B1(n11377), .B2(n11376), .A(n11380), .ZN(n11378) );
  MUX2_X1 U14474 ( .A(n11379), .B(n11378), .S(n19218), .Z(n11388) );
  NOR2_X1 U14475 ( .A1(n11381), .A2(n11380), .ZN(n11382) );
  NAND2_X1 U14476 ( .A1(n11383), .A2(n11382), .ZN(n13037) );
  OAI22_X1 U14477 ( .A1(n11376), .A2(n19224), .B1(n9730), .B2(n10689), .ZN(
        n11384) );
  INV_X1 U14478 ( .A(n11384), .ZN(n11386) );
  NAND3_X1 U14479 ( .A1(n13037), .A2(n11386), .A3(n11385), .ZN(n11387) );
  NOR2_X1 U14480 ( .A1(n11388), .A2(n11387), .ZN(n15507) );
  NAND2_X1 U14481 ( .A1(n15507), .A2(n9827), .ZN(n11389) );
  NAND2_X1 U14482 ( .A1(n11704), .A2(n11389), .ZN(n13992) );
  NOR3_X1 U14483 ( .A1(n19190), .A2(n16297), .A3(n13781), .ZN(n15484) );
  NAND2_X1 U14484 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15484), .ZN(
        n11655) );
  INV_X1 U14485 ( .A(n11655), .ZN(n11390) );
  OR2_X1 U14486 ( .A1(n16309), .A2(n11390), .ZN(n11394) );
  INV_X1 U14487 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11670) );
  NAND2_X1 U14488 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13081) );
  NAND2_X1 U14489 ( .A1(n11670), .A2(n13081), .ZN(n13990) );
  NOR2_X1 U14490 ( .A1(n11670), .A2(n13081), .ZN(n11652) );
  INV_X1 U14491 ( .A(n11704), .ZN(n11391) );
  NOR2_X2 U14492 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19825) );
  AND2_X1 U14493 ( .A1(n19825), .A2(n11189), .ZN(n18878) );
  INV_X2 U14494 ( .A(n19029), .ZN(n19045) );
  NAND2_X1 U14495 ( .A1(n11391), .A2(n19045), .ZN(n13986) );
  OAI21_X1 U14496 ( .B1(n13992), .B2(n11652), .A(n13986), .ZN(n11392) );
  INV_X1 U14497 ( .A(n11392), .ZN(n11393) );
  OAI21_X1 U14498 ( .B1(n14013), .B2(n13990), .A(n11393), .ZN(n13780) );
  INV_X1 U14499 ( .A(n13780), .ZN(n16296) );
  NAND2_X1 U14500 ( .A1(n11394), .A2(n16296), .ZN(n15474) );
  NOR2_X1 U14501 ( .A1(n11696), .A2(n16285), .ZN(n16273) );
  NOR2_X1 U14502 ( .A1(n16309), .A2(n16273), .ZN(n11395) );
  NOR2_X1 U14503 ( .A1(n15474), .A2(n11395), .ZN(n15465) );
  NAND2_X1 U14504 ( .A1(n15465), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16206) );
  AND3_X1 U14505 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11396) );
  AND2_X1 U14506 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15422) );
  NAND2_X1 U14507 ( .A1(n11396), .A2(n15422), .ZN(n16250) );
  NOR2_X1 U14508 ( .A1(n16250), .A2(n16251), .ZN(n14019) );
  NAND2_X1 U14509 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15403) );
  NOR2_X1 U14510 ( .A1(n15403), .A2(n11397), .ZN(n11398) );
  NAND2_X1 U14511 ( .A1(n14019), .A2(n11398), .ZN(n15218) );
  NOR2_X1 U14512 ( .A1(n21055), .A2(n15218), .ZN(n15369) );
  NAND3_X1 U14513 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n15369), .ZN(n15340) );
  NAND2_X1 U14514 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16221) );
  NOR3_X1 U14515 ( .A1(n15181), .A2(n15340), .A3(n16221), .ZN(n11701) );
  INV_X1 U14516 ( .A(n11701), .ZN(n16208) );
  OR2_X1 U14517 ( .A1(n16206), .A2(n16208), .ZN(n11399) );
  NAND2_X1 U14518 ( .A1(n16309), .A2(n13986), .ZN(n16207) );
  NAND2_X1 U14519 ( .A1(n11399), .A2(n16207), .ZN(n15336) );
  AND2_X1 U14520 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11658) );
  INV_X1 U14521 ( .A(n11658), .ZN(n11400) );
  NAND2_X1 U14522 ( .A1(n16207), .A2(n11400), .ZN(n11401) );
  NAND3_X1 U14523 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15267) );
  NAND2_X1 U14524 ( .A1(n16207), .A2(n15267), .ZN(n11402) );
  NAND2_X1 U14525 ( .A1(n15302), .A2(n11402), .ZN(n15264) );
  NOR2_X1 U14526 ( .A1(n16309), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11403) );
  OAI21_X1 U14527 ( .B1(n15264), .B2(n11403), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11651) );
  NAND2_X1 U14528 ( .A1(n19029), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11714) );
  INV_X1 U14529 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19798) );
  AOI22_X1 U14530 ( .A1(n11637), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11405) );
  OAI21_X1 U14531 ( .B1(n11639), .B2(n19798), .A(n11405), .ZN(n15091) );
  NOR2_X1 U14532 ( .A1(n9755), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11406) );
  OR2_X1 U14533 ( .A1(n11666), .A2(n11588), .ZN(n11411) );
  NAND2_X1 U14534 ( .A1(n10699), .A2(n11635), .ZN(n11423) );
  INV_X1 U14535 ( .A(n11418), .ZN(n11408) );
  NOR2_X1 U14536 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19871), .ZN(
        n19858) );
  INV_X1 U14537 ( .A(n19858), .ZN(n11407) );
  NAND2_X1 U14538 ( .A1(n11408), .A2(n11407), .ZN(n11409) );
  AND2_X1 U14539 ( .A1(n11423), .A2(n11409), .ZN(n11410) );
  NAND2_X1 U14540 ( .A1(n11411), .A2(n11410), .ZN(n13041) );
  NOR2_X1 U14541 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(P2_EAX_REG_0__SCAN_IN), 
        .ZN(n11412) );
  OAI22_X1 U14542 ( .A1(n11418), .A2(n11412), .B1(n14257), .B2(n16301), .ZN(
        n11413) );
  INV_X1 U14543 ( .A(n11413), .ZN(n11414) );
  OAI21_X1 U14544 ( .B1(n11639), .B2(n19060), .A(n11414), .ZN(n13042) );
  INV_X1 U14545 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U14546 ( .A1(n11404), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11635), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11415) );
  OAI21_X1 U14547 ( .B1(n11639), .B2(n19763), .A(n11415), .ZN(n11422) );
  INV_X1 U14548 ( .A(n11422), .ZN(n11416) );
  AND2_X1 U14549 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n11417) );
  AOI21_X1 U14550 ( .B1(n11419), .B2(n11418), .A(n11417), .ZN(n11421) );
  NAND2_X1 U14551 ( .A1(n11608), .A2(n11665), .ZN(n11420) );
  NAND2_X1 U14552 ( .A1(n13084), .A2(n13083), .ZN(n13082) );
  NAND2_X1 U14553 ( .A1(n11608), .A2(n10039), .ZN(n11424) );
  OAI211_X1 U14554 ( .C1(n19871), .C2(n19845), .A(n11424), .B(n11423), .ZN(
        n11425) );
  AND3_X1 U14555 ( .A1(n13082), .A2(n11426), .A3(n11425), .ZN(n11427) );
  INV_X1 U14556 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20918) );
  AOI22_X1 U14557 ( .A1(n11637), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11635), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11428) );
  OAI21_X1 U14558 ( .B1(n11639), .B2(n20918), .A(n11428), .ZN(n13427) );
  NAND2_X1 U14559 ( .A1(n11632), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14560 ( .A1(n11635), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11433) );
  NAND2_X1 U14561 ( .A1(n11608), .A2(n11430), .ZN(n11432) );
  NAND2_X1 U14562 ( .A1(n11404), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11431) );
  NAND4_X1 U14563 ( .A1(n11434), .A2(n11433), .A3(n11432), .A4(n11431), .ZN(
        n13477) );
  NAND2_X1 U14564 ( .A1(n13476), .A2(n13477), .ZN(n13478) );
  INV_X1 U14565 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n11438) );
  NAND2_X1 U14566 ( .A1(n11608), .A2(n11435), .ZN(n11437) );
  AOI22_X1 U14567 ( .A1(n11404), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11635), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11436) );
  OAI211_X1 U14568 ( .C1(n11639), .C2(n11438), .A(n11437), .B(n11436), .ZN(
        n13565) );
  INV_X1 U14569 ( .A(n13565), .ZN(n11439) );
  AOI22_X1 U14570 ( .A1(n11632), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11608), 
        .B2(n11440), .ZN(n11442) );
  AOI22_X1 U14571 ( .A1(n11404), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11635), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U14572 ( .A1(n11442), .A2(n11441), .ZN(n13779) );
  NAND2_X1 U14573 ( .A1(n13566), .A2(n13779), .ZN(n13778) );
  NAND2_X1 U14574 ( .A1(n11608), .A2(n11443), .ZN(n11444) );
  INV_X1 U14575 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19769) );
  AOI22_X1 U14576 ( .A1(n11637), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11635), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11445) );
  OAI21_X1 U14577 ( .B1(n11639), .B2(n19769), .A(n11445), .ZN(n13108) );
  NAND2_X1 U14578 ( .A1(n13109), .A2(n13108), .ZN(n11447) );
  NAND2_X1 U14579 ( .A1(n11608), .A2(n11694), .ZN(n11446) );
  INV_X1 U14580 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19771) );
  AOI22_X1 U14581 ( .A1(n11637), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11635), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11448) );
  OAI21_X1 U14582 ( .B1(n11639), .B2(n19771), .A(n11448), .ZN(n13160) );
  INV_X1 U14583 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11468) );
  INV_X1 U14584 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11450) );
  INV_X1 U14585 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11449) );
  OAI22_X1 U14586 ( .A1(n14141), .A2(n11450), .B1(n14099), .B2(n11449), .ZN(
        n11451) );
  INV_X1 U14587 ( .A(n11451), .ZN(n11459) );
  AOI22_X1 U14588 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14589 ( .A1(n14143), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11457) );
  INV_X1 U14590 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11454) );
  NAND2_X1 U14591 ( .A1(n14154), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11453) );
  NAND2_X1 U14592 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11452) );
  OAI211_X1 U14593 ( .C1(n14089), .C2(n11454), .A(n11453), .B(n11452), .ZN(
        n11455) );
  INV_X1 U14594 ( .A(n11455), .ZN(n11456) );
  NAND4_X1 U14595 ( .A1(n11459), .A2(n11458), .A3(n11457), .A4(n11456), .ZN(
        n11465) );
  AOI22_X1 U14596 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14597 ( .A1(n10970), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14598 ( .A1(n14153), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14138), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11461) );
  NAND2_X1 U14599 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11460) );
  NAND4_X1 U14600 ( .A1(n11463), .A2(n11462), .A3(n11461), .A4(n11460), .ZN(
        n11464) );
  NAND2_X1 U14601 ( .A1(n11608), .A2(n13486), .ZN(n11467) );
  AOI22_X1 U14602 ( .A1(n11637), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11635), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11466) );
  OAI211_X1 U14603 ( .C1(n11639), .C2(n11468), .A(n11467), .B(n11466), .ZN(
        n16274) );
  INV_X1 U14604 ( .A(n16274), .ZN(n11469) );
  AOI22_X1 U14605 ( .A1(n11632), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n11404), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11488) );
  INV_X1 U14606 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11470) );
  OAI22_X1 U14607 ( .A1(n11471), .A2(n14141), .B1(n14089), .B2(n11470), .ZN(
        n11472) );
  INV_X1 U14608 ( .A(n11472), .ZN(n11480) );
  AOI22_X1 U14609 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U14610 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n14143), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11478) );
  NAND2_X1 U14611 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11474) );
  NAND2_X1 U14612 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11473) );
  OAI211_X1 U14613 ( .C1(n14099), .C2(n11475), .A(n11474), .B(n11473), .ZN(
        n11476) );
  INV_X1 U14614 ( .A(n11476), .ZN(n11477) );
  NAND4_X1 U14615 ( .A1(n11480), .A2(n11479), .A3(n11478), .A4(n11477), .ZN(
        n11486) );
  AOI22_X1 U14616 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n14077), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14617 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14152), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11483) );
  AOI22_X1 U14618 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11482) );
  NAND2_X1 U14619 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11481) );
  NAND4_X1 U14620 ( .A1(n11484), .A2(n11483), .A3(n11482), .A4(n11481), .ZN(
        n11485) );
  AOI22_X1 U14621 ( .A1(n11608), .A2(n13518), .B1(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n11635), .ZN(n11487) );
  NAND2_X1 U14622 ( .A1(n11488), .A2(n11487), .ZN(n13317) );
  INV_X1 U14623 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11508) );
  INV_X1 U14624 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11490) );
  INV_X1 U14625 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11489) );
  OAI22_X1 U14626 ( .A1(n11490), .A2(n14141), .B1(n14099), .B2(n11489), .ZN(
        n11491) );
  INV_X1 U14627 ( .A(n11491), .ZN(n11499) );
  AOI22_X1 U14628 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11498) );
  AOI22_X1 U14629 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10884), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11497) );
  INV_X1 U14630 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11494) );
  NAND2_X1 U14631 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11493) );
  NAND2_X1 U14632 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11492) );
  OAI211_X1 U14633 ( .C1(n14089), .C2(n11494), .A(n11493), .B(n11492), .ZN(
        n11495) );
  INV_X1 U14634 ( .A(n11495), .ZN(n11496) );
  NAND4_X1 U14635 ( .A1(n11499), .A2(n11498), .A3(n11497), .A4(n11496), .ZN(
        n11505) );
  AOI22_X1 U14636 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n14077), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14637 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14152), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14638 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11501) );
  NAND2_X1 U14639 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11500) );
  NAND4_X1 U14640 ( .A1(n11503), .A2(n11502), .A3(n11501), .A4(n11500), .ZN(
        n11504) );
  NAND2_X1 U14641 ( .A1(n11608), .A2(n13530), .ZN(n11507) );
  AOI22_X1 U14642 ( .A1(n11637), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11506) );
  OAI211_X1 U14643 ( .C1(n11639), .C2(n11508), .A(n11507), .B(n11506), .ZN(
        n11509) );
  INV_X1 U14644 ( .A(n11509), .ZN(n15450) );
  INV_X1 U14645 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11510) );
  OAI22_X1 U14646 ( .A1(n11511), .A2(n14141), .B1(n14089), .B2(n11510), .ZN(
        n11512) );
  INV_X1 U14647 ( .A(n11512), .ZN(n11520) );
  AOI22_X1 U14648 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14649 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n14143), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11518) );
  NAND2_X1 U14650 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11514) );
  NAND2_X1 U14651 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11513) );
  OAI211_X1 U14652 ( .C1(n14099), .C2(n11515), .A(n11514), .B(n11513), .ZN(
        n11516) );
  INV_X1 U14653 ( .A(n11516), .ZN(n11517) );
  NAND4_X1 U14654 ( .A1(n11520), .A2(n11519), .A3(n11518), .A4(n11517), .ZN(
        n11526) );
  AOI22_X1 U14655 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n14150), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11524) );
  AOI22_X1 U14656 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14152), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11523) );
  AOI22_X1 U14657 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11522) );
  NAND2_X1 U14658 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n11521) );
  NAND4_X1 U14659 ( .A1(n11524), .A2(n11523), .A3(n11522), .A4(n11521), .ZN(
        n11525) );
  AOI22_X1 U14660 ( .A1(n11632), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11608), 
        .B2(n13652), .ZN(n11528) );
  AOI22_X1 U14661 ( .A1(n11637), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11527) );
  NAND2_X1 U14662 ( .A1(n11528), .A2(n11527), .ZN(n13464) );
  INV_X1 U14663 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11549) );
  INV_X1 U14664 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11531) );
  INV_X1 U14665 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11529) );
  OAI22_X1 U14666 ( .A1(n11531), .A2(n14089), .B1(n11530), .B2(n11529), .ZN(
        n11532) );
  INV_X1 U14667 ( .A(n11532), .ZN(n11540) );
  AOI22_X1 U14668 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11539) );
  AOI22_X1 U14669 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10884), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11538) );
  INV_X1 U14670 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11535) );
  NAND2_X1 U14671 ( .A1(n14154), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11534) );
  NAND2_X1 U14672 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11533) );
  OAI211_X1 U14673 ( .C1(n14099), .C2(n11535), .A(n11534), .B(n11533), .ZN(
        n11536) );
  INV_X1 U14674 ( .A(n11536), .ZN(n11537) );
  NAND4_X1 U14675 ( .A1(n11540), .A2(n11539), .A3(n11538), .A4(n11537), .ZN(
        n11546) );
  AOI22_X1 U14676 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n14077), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U14677 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n14155), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11543) );
  AOI22_X1 U14678 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14153), .B1(
        n14138), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11542) );
  NAND2_X1 U14679 ( .A1(n10970), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11541) );
  NAND4_X1 U14680 ( .A1(n11544), .A2(n11543), .A3(n11542), .A4(n11541), .ZN(
        n11545) );
  NAND2_X1 U14681 ( .A1(n11608), .A2(n13651), .ZN(n11548) );
  AOI22_X1 U14682 ( .A1(n11637), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11547) );
  OAI211_X1 U14683 ( .C1(n11639), .C2(n11549), .A(n11548), .B(n11547), .ZN(
        n11550) );
  INV_X1 U14684 ( .A(n11550), .ZN(n13471) );
  NOR2_X2 U14685 ( .A1(n13472), .A2(n13471), .ZN(n13525) );
  OAI22_X1 U14686 ( .A1(n14141), .A2(n14084), .B1(n14089), .B2(n11551), .ZN(
        n11552) );
  INV_X1 U14687 ( .A(n11552), .ZN(n11560) );
  AOI22_X1 U14688 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14689 ( .A1(n14143), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U14690 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11554) );
  NAND2_X1 U14691 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11553) );
  OAI211_X1 U14692 ( .C1(n14099), .C2(n11555), .A(n11554), .B(n11553), .ZN(
        n11556) );
  INV_X1 U14693 ( .A(n11556), .ZN(n11557) );
  NAND4_X1 U14694 ( .A1(n11560), .A2(n11559), .A3(n11558), .A4(n11557), .ZN(
        n11566) );
  AOI22_X1 U14695 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14696 ( .A1(n10970), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14697 ( .A1(n14154), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11562) );
  NAND2_X1 U14698 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11561) );
  NAND4_X1 U14699 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .ZN(
        n11565) );
  AOI22_X1 U14700 ( .A1(n11632), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n11608), 
        .B2(n13633), .ZN(n11568) );
  AOI22_X1 U14701 ( .A1(n11637), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11567) );
  NAND2_X1 U14702 ( .A1(n11568), .A2(n11567), .ZN(n13524) );
  NAND2_X1 U14703 ( .A1(n13525), .A2(n13524), .ZN(n16248) );
  OAI22_X1 U14704 ( .A1(n11570), .A2(n14141), .B1(n14099), .B2(n11569), .ZN(
        n11571) );
  INV_X1 U14705 ( .A(n11571), .ZN(n11579) );
  AOI22_X1 U14706 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14707 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n14143), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11577) );
  NAND2_X1 U14708 ( .A1(n14154), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11573) );
  NAND2_X1 U14709 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11572) );
  OAI211_X1 U14710 ( .C1(n14089), .C2(n11574), .A(n11573), .B(n11572), .ZN(
        n11575) );
  INV_X1 U14711 ( .A(n11575), .ZN(n11576) );
  NAND4_X1 U14712 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n11585) );
  AOI22_X1 U14713 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n14077), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14714 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n14152), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14715 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14153), .B1(
        n14138), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U14716 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11580) );
  NAND4_X1 U14717 ( .A1(n11583), .A2(n11582), .A3(n11581), .A4(n11580), .ZN(
        n11584) );
  INV_X1 U14718 ( .A(n13636), .ZN(n11587) );
  AOI22_X1 U14719 ( .A1(n11637), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11586) );
  OAI21_X1 U14720 ( .B1(n11588), .B2(n11587), .A(n11586), .ZN(n11589) );
  AOI21_X1 U14721 ( .B1(n11632), .B2(P2_REIP_REG_14__SCAN_IN), .A(n11589), 
        .ZN(n16247) );
  NOR2_X4 U14722 ( .A1(n16248), .A2(n16247), .ZN(n16246) );
  AOI22_X1 U14723 ( .A1(n11632), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n11404), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n11610) );
  INV_X1 U14724 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11591) );
  INV_X1 U14725 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11590) );
  OAI22_X1 U14726 ( .A1(n11591), .A2(n14141), .B1(n14089), .B2(n11590), .ZN(
        n11592) );
  INV_X1 U14727 ( .A(n11592), .ZN(n11600) );
  AOI22_X1 U14728 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14729 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n14143), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11598) );
  INV_X1 U14730 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11595) );
  NAND2_X1 U14731 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11594) );
  NAND2_X1 U14732 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11593) );
  OAI211_X1 U14733 ( .C1(n14099), .C2(n11595), .A(n11594), .B(n11593), .ZN(
        n11596) );
  INV_X1 U14734 ( .A(n11596), .ZN(n11597) );
  NAND4_X1 U14735 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(
        n11606) );
  AOI22_X1 U14736 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n14077), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14737 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n14152), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14738 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11602) );
  INV_X1 U14739 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n20819) );
  OR2_X1 U14740 ( .A1(n14105), .A2(n20819), .ZN(n11601) );
  NAND4_X1 U14741 ( .A1(n11604), .A2(n11603), .A3(n11602), .A4(n11601), .ZN(
        n11605) );
  NOR2_X1 U14742 ( .A1(n11606), .A2(n11605), .ZN(n13805) );
  INV_X1 U14743 ( .A(n13805), .ZN(n11607) );
  AOI22_X1 U14744 ( .A1(n11608), .A2(n11607), .B1(n11635), .B2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11609) );
  NAND2_X1 U14745 ( .A1(n11610), .A2(n11609), .ZN(n12911) );
  INV_X1 U14746 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U14747 ( .A1(n11637), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11611) );
  OAI21_X1 U14748 ( .B1(n11639), .B2(n19785), .A(n11611), .ZN(n11612) );
  INV_X1 U14749 ( .A(n11612), .ZN(n14015) );
  INV_X1 U14750 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19787) );
  AOI22_X1 U14751 ( .A1(n11637), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11613) );
  OAI21_X1 U14752 ( .B1(n11639), .B2(n19787), .A(n11613), .ZN(n13808) );
  INV_X1 U14753 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19789) );
  AOI22_X1 U14754 ( .A1(n11637), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11614) );
  OAI21_X1 U14755 ( .B1(n11639), .B2(n19789), .A(n11614), .ZN(n11615) );
  INV_X1 U14756 ( .A(n11615), .ZN(n15388) );
  INV_X1 U14757 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19790) );
  AOI22_X1 U14758 ( .A1(n11637), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11616) );
  OAI21_X1 U14759 ( .B1(n11639), .B2(n19790), .A(n11616), .ZN(n13853) );
  INV_X1 U14760 ( .A(n13853), .ZN(n11617) );
  NOR2_X2 U14761 ( .A1(n15391), .A2(n11617), .ZN(n14932) );
  INV_X1 U14762 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19792) );
  AOI22_X1 U14763 ( .A1(n11637), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11618) );
  OAI21_X1 U14764 ( .B1(n11639), .B2(n19792), .A(n11618), .ZN(n14931) );
  AND2_X2 U14765 ( .A1(n14932), .A2(n14931), .ZN(n14934) );
  INV_X1 U14766 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19794) );
  INV_X1 U14767 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n12947) );
  OAI222_X1 U14768 ( .A1(n11639), .A2(n19794), .B1(n11620), .B2(n12947), .C1(
        n15181), .C2(n11619), .ZN(n14921) );
  NAND2_X1 U14769 ( .A1(n11632), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14770 ( .A1(n11637), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11621) );
  AND2_X1 U14771 ( .A1(n11622), .A2(n11621), .ZN(n15343) );
  NAND2_X1 U14772 ( .A1(n11632), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14773 ( .A1(n11637), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11623) );
  NAND2_X1 U14774 ( .A1(n11624), .A2(n11623), .ZN(n14911) );
  NAND2_X1 U14775 ( .A1(n11632), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11626) );
  AOI22_X1 U14776 ( .A1(n11637), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11625) );
  AND2_X1 U14777 ( .A1(n11626), .A2(n11625), .ZN(n15081) );
  OR2_X2 U14778 ( .A1(n15082), .A2(n15081), .ZN(n15084) );
  NAND2_X1 U14779 ( .A1(n11632), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U14780 ( .A1(n11637), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11627) );
  AND2_X1 U14781 ( .A1(n11628), .A2(n11627), .ZN(n15074) );
  INV_X1 U14782 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19807) );
  AOI22_X1 U14783 ( .A1(n11637), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11629) );
  OAI21_X1 U14784 ( .B1(n11639), .B2(n19807), .A(n11629), .ZN(n15065) );
  NAND2_X1 U14785 ( .A1(n11632), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U14786 ( .A1(n11637), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11630) );
  AND2_X1 U14787 ( .A1(n11631), .A2(n11630), .ZN(n15055) );
  NAND2_X1 U14788 ( .A1(n11632), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14789 ( .A1(n11637), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11633) );
  AND2_X1 U14790 ( .A1(n11634), .A2(n11633), .ZN(n15046) );
  INV_X1 U14791 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20975) );
  AOI22_X1 U14792 ( .A1(n11637), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11636) );
  OAI21_X1 U14793 ( .B1(n11639), .B2(n20975), .A(n11636), .ZN(n14325) );
  INV_X1 U14794 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19814) );
  AOI22_X1 U14795 ( .A1(n11637), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n11635), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11638) );
  OAI21_X1 U14796 ( .B1(n11639), .B2(n19814), .A(n11638), .ZN(n11640) );
  XNOR2_X1 U14797 ( .A(n9805), .B(n11640), .ZN(n15992) );
  NOR2_X1 U14798 ( .A1(n19241), .A2(n19224), .ZN(n11641) );
  AND2_X1 U14799 ( .A1(n11376), .A2(n11641), .ZN(n11642) );
  NAND2_X1 U14800 ( .A1(n11643), .A2(n11642), .ZN(n15495) );
  INV_X1 U14801 ( .A(n15495), .ZN(n11644) );
  AND2_X1 U14802 ( .A1(n11645), .A2(n11644), .ZN(n16314) );
  INV_X1 U14803 ( .A(n16314), .ZN(n11649) );
  NAND2_X1 U14804 ( .A1(n11647), .A2(n10757), .ZN(n11648) );
  NAND2_X1 U14805 ( .A1(n11649), .A2(n11648), .ZN(n11650) );
  INV_X1 U14806 ( .A(n11652), .ZN(n13989) );
  NAND2_X1 U14807 ( .A1(n14013), .A2(n13989), .ZN(n11653) );
  NAND2_X1 U14808 ( .A1(n11653), .A2(n13990), .ZN(n11654) );
  INV_X1 U14809 ( .A(n15340), .ZN(n15164) );
  NAND2_X1 U14810 ( .A1(n15471), .A2(n15164), .ZN(n15353) );
  INV_X1 U14811 ( .A(n16221), .ZN(n11656) );
  NAND2_X1 U14812 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n11656), .ZN(
        n11657) );
  NOR2_X1 U14813 ( .A1(n16224), .A2(n11657), .ZN(n15330) );
  NAND2_X1 U14814 ( .A1(n15330), .A2(n11658), .ZN(n15305) );
  NOR4_X1 U14815 ( .A1(n15305), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15267), .A4(n11659), .ZN(n11660) );
  NAND2_X1 U14816 ( .A1(n11663), .A2(n11664), .ZN(n11684) );
  NAND2_X1 U14817 ( .A1(n11691), .A2(n13775), .ZN(n11685) );
  NAND2_X1 U14818 ( .A1(n16304), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16303) );
  INV_X1 U14819 ( .A(n16303), .ZN(n11668) );
  XNOR2_X1 U14820 ( .A(n11666), .B(n11665), .ZN(n11667) );
  NAND2_X1 U14821 ( .A1(n11668), .A2(n11667), .ZN(n11669) );
  XOR2_X1 U14822 ( .A(n11668), .B(n11667), .Z(n13006) );
  NAND2_X1 U14823 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13006), .ZN(
        n13005) );
  NAND2_X1 U14824 ( .A1(n11669), .A2(n13005), .ZN(n11673) );
  XNOR2_X1 U14825 ( .A(n11670), .B(n11673), .ZN(n13988) );
  XNOR2_X1 U14826 ( .A(n11672), .B(n11671), .ZN(n13987) );
  NAND2_X1 U14827 ( .A1(n13988), .A2(n13987), .ZN(n11675) );
  NAND2_X1 U14828 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11673), .ZN(
        n11674) );
  NAND2_X1 U14829 ( .A1(n11675), .A2(n11674), .ZN(n11676) );
  XNOR2_X1 U14830 ( .A(n11676), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13598) );
  INV_X1 U14831 ( .A(n11676), .ZN(n11677) );
  OAI22_X1 U14832 ( .A1(n13599), .A2(n13598), .B1(n11677), .B2(n16297), .ZN(
        n19158) );
  XNOR2_X1 U14833 ( .A(n11678), .B(n11679), .ZN(n19159) );
  NAND2_X1 U14834 ( .A1(n19159), .A2(n19190), .ZN(n11680) );
  NAND2_X1 U14835 ( .A1(n19158), .A2(n11680), .ZN(n11683) );
  INV_X1 U14836 ( .A(n19159), .ZN(n11681) );
  NAND2_X1 U14837 ( .A1(n11681), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11682) );
  NAND2_X1 U14838 ( .A1(n11683), .A2(n11682), .ZN(n13776) );
  NAND2_X1 U14839 ( .A1(n11684), .A2(n13781), .ZN(n13774) );
  NAND2_X1 U14840 ( .A1(n13776), .A2(n13774), .ZN(n11690) );
  MUX2_X1 U14841 ( .A(n11691), .B(n11685), .S(n11690), .Z(n11689) );
  INV_X1 U14842 ( .A(n13775), .ZN(n11687) );
  NAND2_X1 U14843 ( .A1(n11687), .A2(n11686), .ZN(n11688) );
  NAND2_X1 U14844 ( .A1(n11689), .A2(n11688), .ZN(n15257) );
  NAND2_X1 U14845 ( .A1(n15257), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15256) );
  NAND2_X1 U14846 ( .A1(n11690), .A2(n13775), .ZN(n11692) );
  NAND2_X1 U14847 ( .A1(n11692), .A2(n11691), .ZN(n11693) );
  XNOR2_X1 U14848 ( .A(n11661), .B(n11694), .ZN(n11695) );
  INV_X1 U14849 ( .A(n11695), .ZN(n11697) );
  NAND2_X1 U14850 ( .A1(n11697), .A2(n11696), .ZN(n15242) );
  NOR2_X1 U14851 ( .A1(n11661), .A2(n14045), .ZN(n11698) );
  XNOR2_X1 U14852 ( .A(n11698), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16185) );
  INV_X1 U14853 ( .A(n11661), .ZN(n11700) );
  NOR2_X2 U14854 ( .A1(n16109), .A2(n16210), .ZN(n15327) );
  XOR2_X1 U14855 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11702), .Z(
        n11717) );
  NOR2_X1 U14856 ( .A1(n11195), .A2(n16348), .ZN(n11703) );
  NAND2_X1 U14857 ( .A1(n19883), .A2(n19737), .ZN(n11706) );
  NOR2_X2 U14858 ( .A1(n12928), .A2(n14257), .ZN(n19175) );
  NAND2_X1 U14859 ( .A1(n11708), .A2(n19175), .ZN(n11719) );
  NOR2_X1 U14860 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19827) );
  OR2_X1 U14861 ( .A1(n19825), .A2(n19827), .ZN(n19846) );
  NAND2_X1 U14862 ( .A1(n19846), .A2(n19884), .ZN(n11709) );
  INV_X1 U14863 ( .A(n16345), .ZN(n11711) );
  INV_X1 U14864 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19882) );
  NAND2_X1 U14865 ( .A1(n19882), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11710) );
  NAND2_X1 U14866 ( .A1(n11711), .A2(n11710), .ZN(n19168) );
  INV_X1 U14867 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16114) );
  INV_X1 U14868 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15182) );
  INV_X1 U14869 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16128) );
  INV_X1 U14870 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18924) );
  INV_X1 U14871 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16097) );
  INV_X1 U14872 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15133) );
  INV_X1 U14873 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14053) );
  INV_X1 U14874 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15123) );
  NOR2_X1 U14875 ( .A1(n11189), .A2(n19882), .ZN(n19847) );
  NAND2_X1 U14876 ( .A1(n19169), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11713) );
  INV_X1 U14877 ( .A(n12928), .ZN(n11716) );
  NAND2_X1 U14878 ( .A1(n11716), .A2(n14257), .ZN(n19177) );
  NAND2_X1 U14879 ( .A1(n11719), .A2(n11718), .ZN(P2_U2983) );
  NOR2_X4 U14880 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11952), .ZN(
        n11729) );
  NOR2_X4 U14881 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13361) );
  AOI22_X1 U14882 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11917), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11722) );
  AND2_X2 U14883 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13344) );
  AND3_X4 U14884 ( .A1(n13344), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n14035), .ZN(n11910) );
  NOR2_X2 U14885 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14886 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9720), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11721) );
  AND2_X2 U14887 ( .A1(n11723), .A2(n13361), .ZN(n11901) );
  AOI22_X1 U14888 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14889 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11725) );
  AND2_X4 U14890 ( .A1(n11853), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11731) );
  AND2_X4 U14891 ( .A1(n11732), .A2(n11731), .ZN(n11965) );
  AND2_X4 U14892 ( .A1(n13345), .A2(n11731), .ZN(n11959) );
  AOI22_X1 U14893 ( .A1(n11965), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14894 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12015), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11735) );
  AND2_X2 U14895 ( .A1(n13361), .A2(n13346), .ZN(n12016) );
  AOI22_X1 U14896 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11734) );
  AND2_X4 U14897 ( .A1(n11731), .A2(n13346), .ZN(n12010) );
  AOI22_X1 U14898 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11898), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11733) );
  INV_X1 U14899 ( .A(n11841), .ZN(n11845) );
  AOI22_X1 U14900 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11739) );
  AOI22_X1 U14901 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11738) );
  AOI22_X1 U14902 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11737) );
  AOI22_X1 U14903 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14904 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14905 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14906 ( .A1(n11965), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14907 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11917), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11740) );
  NAND2_X2 U14908 ( .A1(n9801), .A2(n10238), .ZN(n20176) );
  NAND2_X1 U14909 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11747) );
  NAND2_X1 U14910 ( .A1(n11965), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11746) );
  NAND2_X1 U14911 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11745) );
  NAND2_X1 U14912 ( .A1(n12016), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11744) );
  NAND2_X1 U14913 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11751) );
  NAND2_X1 U14914 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11750) );
  NAND2_X1 U14915 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11749) );
  NAND2_X1 U14916 ( .A1(n11917), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11748) );
  NAND2_X1 U14917 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11755) );
  NAND2_X1 U14918 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11754) );
  NAND2_X1 U14919 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11753) );
  NAND2_X1 U14920 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11752) );
  NAND2_X1 U14921 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11759) );
  NAND2_X1 U14922 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11758) );
  NAND2_X1 U14923 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11757) );
  NAND2_X1 U14924 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11756) );
  NAND3_X1 U14926 ( .A1(n11845), .A2(n11849), .A3(n20171), .ZN(n11783) );
  AOI22_X1 U14927 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11769) );
  NAND2_X1 U14928 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11765) );
  NAND2_X1 U14929 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11764) );
  AOI22_X1 U14930 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11767) );
  AOI22_X1 U14931 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U14932 ( .A1(n11965), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11772) );
  AOI22_X1 U14933 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U14934 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11917), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11770) );
  AOI22_X1 U14935 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11965), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11777) );
  AOI22_X1 U14936 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U14937 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14938 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U14939 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U14940 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14941 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11917), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11778) );
  NAND2_X1 U14942 ( .A1(n11978), .A2(n20165), .ZN(n11782) );
  NOR2_X2 U14943 ( .A1(n11783), .A2(n11782), .ZN(n12962) );
  AOI22_X1 U14944 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11965), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14945 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9758), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14946 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14947 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11819), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11784) );
  NAND4_X1 U14948 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11793) );
  AOI22_X1 U14949 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U14950 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U14951 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U14952 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11917), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11788) );
  NAND4_X1 U14953 ( .A1(n11791), .A2(n11790), .A3(n11789), .A4(n11788), .ZN(
        n11792) );
  NAND2_X1 U14954 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11797) );
  NAND2_X1 U14955 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11796) );
  NAND2_X1 U14956 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11795) );
  NAND2_X1 U14957 ( .A1(n11917), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11794) );
  NAND2_X1 U14958 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11801) );
  NAND2_X1 U14959 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11800) );
  NAND2_X1 U14960 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11799) );
  NAND2_X1 U14961 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11798) );
  NAND2_X1 U14962 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11805) );
  NAND2_X1 U14963 ( .A1(n11965), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11804) );
  NAND2_X1 U14964 ( .A1(n11819), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11803) );
  NAND2_X1 U14965 ( .A1(n12016), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11802) );
  NAND2_X1 U14966 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11809) );
  NAND2_X1 U14967 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11808) );
  NAND2_X1 U14968 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11807) );
  NAND2_X1 U14969 ( .A1(n9757), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11806) );
  NAND2_X1 U14971 ( .A1(n11965), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11818) );
  NAND2_X1 U14972 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11817) );
  NAND2_X1 U14973 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11816) );
  NAND2_X1 U14974 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11815) );
  NAND2_X1 U14975 ( .A1(n11898), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11823) );
  NAND2_X1 U14976 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11822) );
  NAND2_X1 U14977 ( .A1(n11916), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11821) );
  NAND2_X1 U14978 ( .A1(n11876), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11827) );
  NAND2_X1 U14979 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11826) );
  NAND2_X1 U14980 ( .A1(n11901), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11825) );
  NAND2_X1 U14981 ( .A1(n12016), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11824) );
  NAND2_X1 U14982 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11830) );
  NAND2_X1 U14983 ( .A1(n11917), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11829) );
  NAND2_X1 U14984 ( .A1(n11960), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11828) );
  NAND3_X1 U14985 ( .A1(n11830), .A2(n11829), .A3(n11828), .ZN(n11831) );
  INV_X2 U14986 ( .A(n20171), .ZN(n13136) );
  NAND2_X1 U14987 ( .A1(n13136), .A2(n20188), .ZN(n12254) );
  NAND2_X1 U14988 ( .A1(n12254), .A2(n12863), .ZN(n11836) );
  NAND2_X1 U14989 ( .A1(n12733), .A2(n20181), .ZN(n11835) );
  NAND2_X1 U14990 ( .A1(n11836), .A2(n11835), .ZN(n11842) );
  INV_X1 U14991 ( .A(n11842), .ZN(n11837) );
  NAND2_X1 U14992 ( .A1(n11837), .A2(n9772), .ZN(n12930) );
  OR2_X2 U14993 ( .A1(n12930), .A2(n20155), .ZN(n12591) );
  AND2_X1 U14994 ( .A1(n20144), .A2(n20165), .ZN(n12726) );
  NAND2_X1 U14995 ( .A1(n12726), .A2(n12595), .ZN(n11843) );
  OR2_X1 U14996 ( .A1(n11845), .A2(n20144), .ZN(n11866) );
  OAI211_X1 U14997 ( .C1(n12551), .C2(n12619), .A(n13141), .B(n11866), .ZN(
        n12589) );
  INV_X1 U14998 ( .A(n11846), .ZN(n11865) );
  NAND2_X1 U14999 ( .A1(n20144), .A2(n20155), .ZN(n14474) );
  NAND2_X1 U15000 ( .A1(n11865), .A2(n14474), .ZN(n11847) );
  OR2_X2 U15001 ( .A1(n20155), .A2(n20144), .ZN(n20803) );
  NAND2_X1 U15002 ( .A1(n11848), .A2(n20803), .ZN(n12597) );
  NAND2_X1 U15003 ( .A1(n11848), .A2(n20171), .ZN(n11851) );
  NAND2_X1 U15004 ( .A1(n11849), .A2(n20181), .ZN(n12602) );
  AND2_X1 U15005 ( .A1(n12602), .A2(n20188), .ZN(n11850) );
  INV_X1 U15006 ( .A(n12816), .ZN(n11870) );
  NAND2_X1 U15007 ( .A1(n14032), .A2(n20708), .ZN(n12831) );
  NAND2_X1 U15008 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11949) );
  OAI21_X1 U15009 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11949), .ZN(n20457) );
  NAND2_X1 U15010 ( .A1(n20707), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15568) );
  NAND2_X1 U15011 ( .A1(n15568), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11944) );
  OAI21_X1 U15012 ( .B1(n12831), .B2(n20457), .A(n11944), .ZN(n11854) );
  INV_X1 U15013 ( .A(n11854), .ZN(n11855) );
  INV_X1 U15014 ( .A(n20257), .ZN(n11874) );
  INV_X1 U15015 ( .A(n15568), .ZN(n11858) );
  MUX2_X1 U15016 ( .A(n11858), .B(n12831), .S(n20568), .Z(n11859) );
  OAI21_X2 U15017 ( .B1(n11951), .B2(n14035), .A(n11859), .ZN(n11890) );
  NAND2_X1 U15018 ( .A1(n11849), .A2(n20188), .ZN(n14564) );
  NAND2_X1 U15019 ( .A1(n14564), .A2(n12863), .ZN(n13113) );
  NAND3_X1 U15020 ( .A1(n13113), .A2(n20165), .A3(n12602), .ZN(n11860) );
  NAND2_X1 U15021 ( .A1(n11860), .A2(n12619), .ZN(n11863) );
  INV_X1 U15022 ( .A(n11861), .ZN(n11862) );
  NAND2_X1 U15023 ( .A1(n11863), .A2(n11862), .ZN(n11864) );
  AND2_X1 U15024 ( .A1(n20144), .A2(n12606), .ZN(n14350) );
  INV_X1 U15025 ( .A(n14350), .ZN(n14472) );
  NAND2_X1 U15026 ( .A1(n11864), .A2(n14472), .ZN(n11869) );
  OR2_X1 U15027 ( .A1(n11865), .A2(n20181), .ZN(n11867) );
  NAND2_X1 U15028 ( .A1(n14032), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19897) );
  INV_X1 U15029 ( .A(n19897), .ZN(n11868) );
  NAND4_X1 U15030 ( .A1(n11869), .A2(n13142), .A3(n11868), .A4(n14474), .ZN(
        n11872) );
  INV_X1 U15031 ( .A(n11875), .ZN(n11873) );
  AOI22_X1 U15032 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12515), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U15033 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U15034 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U15035 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11877) );
  NAND4_X1 U15036 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(
        n11886) );
  AOI22_X1 U15037 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U15038 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U15039 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U15040 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11881) );
  NAND4_X1 U15041 ( .A1(n11884), .A2(n11883), .A3(n11882), .A4(n11881), .ZN(
        n11885) );
  BUF_X1 U15042 ( .A(n11891), .Z(n12498) );
  BUF_X1 U15043 ( .A(n11959), .Z(n11892) );
  AOI22_X1 U15044 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U15045 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11896) );
  BUF_X1 U15046 ( .A(n11910), .Z(n12493) );
  AOI22_X1 U15047 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U15048 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11894) );
  NAND4_X1 U15049 ( .A1(n11897), .A2(n11896), .A3(n11895), .A4(n11894), .ZN(
        n11909) );
  AOI22_X1 U15050 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11898), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U15051 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U15052 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U15053 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11904) );
  NAND4_X1 U15054 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11908) );
  NOR2_X1 U15055 ( .A1(n12009), .A2(n12780), .ZN(n11934) );
  AOI22_X1 U15056 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U15057 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U15058 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U15059 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11912) );
  NAND4_X1 U15060 ( .A1(n11915), .A2(n11914), .A3(n11913), .A4(n11912), .ZN(
        n11923) );
  AOI22_X1 U15061 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11921) );
  AOI22_X1 U15062 ( .A1(n11958), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U15063 ( .A1(n11893), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U15064 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11918) );
  NAND4_X1 U15065 ( .A1(n11921), .A2(n11920), .A3(n11919), .A4(n11918), .ZN(
        n11922) );
  MUX2_X1 U15066 ( .A(n11934), .B(n12787), .S(n12727), .Z(n11924) );
  INV_X1 U15067 ( .A(n11924), .ZN(n11925) );
  NOR2_X1 U15068 ( .A1(n20144), .A2(n20708), .ZN(n11926) );
  INV_X1 U15069 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11927) );
  OR2_X1 U15070 ( .A1(n12568), .A2(n11927), .ZN(n11931) );
  NAND2_X1 U15071 ( .A1(n20144), .A2(n12730), .ZN(n11929) );
  NAND2_X1 U15072 ( .A1(n20171), .A2(n12780), .ZN(n11928) );
  INV_X1 U15073 ( .A(n12787), .ZN(n11932) );
  NAND2_X1 U15074 ( .A1(n20144), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12008) );
  INV_X1 U15075 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11933) );
  OR2_X1 U15076 ( .A1(n12568), .A2(n11933), .ZN(n11936) );
  INV_X1 U15077 ( .A(n11934), .ZN(n11935) );
  OAI211_X1 U15078 ( .C1(n11937), .C2(n12008), .A(n11936), .B(n11935), .ZN(
        n11985) );
  INV_X1 U15079 ( .A(n12734), .ZN(n11940) );
  NAND2_X1 U15080 ( .A1(n11987), .A2(n11942), .ZN(n11976) );
  INV_X1 U15081 ( .A(n11943), .ZN(n11946) );
  NAND2_X1 U15082 ( .A1(n11944), .A2(n11853), .ZN(n11945) );
  NAND2_X1 U15083 ( .A1(n11946), .A2(n11945), .ZN(n11947) );
  INV_X1 U15084 ( .A(n11949), .ZN(n11948) );
  NAND2_X1 U15085 ( .A1(n11948), .A2(n12539), .ZN(n20489) );
  NAND2_X1 U15086 ( .A1(n11949), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11950) );
  OR2_X1 U15087 ( .A1(n11951), .A2(n11952), .ZN(n11954) );
  NAND2_X1 U15088 ( .A1(n15568), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11953) );
  AOI22_X1 U15089 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U15090 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15091 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15092 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11961) );
  NAND4_X1 U15093 ( .A1(n11964), .A2(n11963), .A3(n11962), .A4(n11961), .ZN(
        n11971) );
  INV_X1 U15094 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n21080) );
  AOI22_X1 U15095 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11969) );
  AOI22_X1 U15096 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U15097 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U15098 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11966) );
  NAND4_X1 U15099 ( .A1(n11969), .A2(n11968), .A3(n11967), .A4(n11966), .ZN(
        n11970) );
  INV_X1 U15100 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11972) );
  OAI22_X1 U15101 ( .A1(n12568), .A2(n11972), .B1(n12741), .B2(n12008), .ZN(
        n11973) );
  XNOR2_X1 U15102 ( .A(n11974), .B(n11973), .ZN(n11975) );
  NAND2_X1 U15103 ( .A1(n11975), .A2(n11976), .ZN(n11977) );
  INV_X1 U15104 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11979) );
  XNOR2_X1 U15105 ( .A(n11979), .B(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n19983) );
  NAND2_X1 U15106 ( .A1(n11980), .A2(n21079), .ZN(n12055) );
  NAND2_X1 U15107 ( .A1(n11980), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12273) );
  OAI21_X1 U15108 ( .B1(n19983), .B2(n12055), .A(n12273), .ZN(n11981) );
  AOI21_X1 U15109 ( .B1(n12534), .B2(P1_EAX_REG_2__SCAN_IN), .A(n11981), .ZN(
        n11983) );
  AND2_X1 U15110 ( .A1(n13120), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11996) );
  NAND2_X1 U15111 ( .A1(n11996), .A2(n9746), .ZN(n11982) );
  NAND2_X1 U15112 ( .A1(n12820), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12004) );
  NAND2_X1 U15113 ( .A1(n11984), .A2(n12004), .ZN(n13337) );
  INV_X1 U15114 ( .A(n11985), .ZN(n11986) );
  NAND2_X1 U15115 ( .A1(n20223), .A2(n12231), .ZN(n11992) );
  AOI22_X1 U15116 ( .A1(n12075), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n11980), .ZN(n11990) );
  NAND2_X1 U15117 ( .A1(n11996), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11989) );
  AND2_X1 U15118 ( .A1(n11990), .A2(n11989), .ZN(n11991) );
  NAND2_X1 U15119 ( .A1(n11992), .A2(n11991), .ZN(n13111) );
  NAND2_X1 U15120 ( .A1(n20222), .A2(n11978), .ZN(n11994) );
  NAND2_X1 U15121 ( .A1(n11994), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13092) );
  INV_X1 U15122 ( .A(n11996), .ZN(n12059) );
  NAND2_X1 U15123 ( .A1(n12075), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11998) );
  NAND2_X1 U15124 ( .A1(n11980), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11997) );
  OAI211_X1 U15125 ( .C1(n12059), .C2(n14035), .A(n11998), .B(n11997), .ZN(
        n11999) );
  AOI21_X1 U15126 ( .B1(n20256), .B2(n12231), .A(n11999), .ZN(n12000) );
  OR2_X1 U15127 ( .A1(n13092), .A2(n12000), .ZN(n13093) );
  INV_X1 U15128 ( .A(n12000), .ZN(n13094) );
  OR2_X1 U15129 ( .A1(n13094), .A2(n12055), .ZN(n12001) );
  NAND2_X1 U15130 ( .A1(n13093), .A2(n12001), .ZN(n13110) );
  NAND2_X1 U15131 ( .A1(n13111), .A2(n13110), .ZN(n13336) );
  NOR3_X1 U15132 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12539), .A3(
        n20524), .ZN(n20377) );
  NAND2_X1 U15133 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20377), .ZN(
        n20371) );
  NAND3_X1 U15134 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20647) );
  NOR2_X1 U15135 ( .A1(n20568), .A2(n20647), .ZN(n20696) );
  AOI21_X1 U15136 ( .B1(n20371), .B2(n20488), .A(n20696), .ZN(n20400) );
  INV_X1 U15137 ( .A(n12831), .ZN(n12005) );
  AOI22_X1 U15138 ( .A1(n20400), .A2(n12005), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15568), .ZN(n12006) );
  AOI22_X1 U15139 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15140 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12013) );
  INV_X1 U15141 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n20827) );
  AOI22_X1 U15142 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11960), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12012) );
  AOI22_X1 U15143 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12011) );
  NAND4_X1 U15144 ( .A1(n12014), .A2(n12013), .A3(n12012), .A4(n12011), .ZN(
        n12022) );
  AOI22_X1 U15145 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U15146 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15147 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15148 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12017) );
  NAND4_X1 U15149 ( .A1(n12020), .A2(n12019), .A3(n12018), .A4(n12017), .ZN(
        n12021) );
  AOI22_X1 U15150 ( .A1(n12582), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12585), .B2(n12755), .ZN(n12023) );
  INV_X1 U15151 ( .A(n13373), .ZN(n12024) );
  NAND2_X1 U15152 ( .A1(n12025), .A2(n12024), .ZN(n12026) );
  INV_X1 U15153 ( .A(n20137), .ZN(n12027) );
  INV_X1 U15154 ( .A(n12029), .ZN(n12031) );
  INV_X1 U15155 ( .A(n12054), .ZN(n12030) );
  OAI21_X1 U15156 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12031), .A(
        n12030), .ZN(n14477) );
  AOI22_X1 U15157 ( .A1(n13611), .A2(n14477), .B1(n12820), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12033) );
  NAND2_X1 U15158 ( .A1(n12534), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12032) );
  OAI211_X1 U15159 ( .C1(n12059), .C2(n12543), .A(n12033), .B(n12032), .ZN(
        n12034) );
  INV_X1 U15160 ( .A(n12034), .ZN(n12035) );
  NAND2_X1 U15161 ( .A1(n12036), .A2(n12035), .ZN(n13404) );
  INV_X1 U15162 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15163 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12498), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U15164 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11903), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U15165 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11892), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U15166 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12520), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12038) );
  NAND4_X1 U15167 ( .A1(n12041), .A2(n12040), .A3(n12039), .A4(n12038), .ZN(
        n12047) );
  AOI22_X1 U15168 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15169 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11911), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15170 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U15171 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12042) );
  NAND4_X1 U15172 ( .A1(n12045), .A2(n12044), .A3(n12043), .A4(n12042), .ZN(
        n12046) );
  NAND2_X1 U15173 ( .A1(n12585), .A2(n12756), .ZN(n12048) );
  INV_X1 U15174 ( .A(n12052), .ZN(n12050) );
  NAND2_X1 U15175 ( .A1(n9895), .A2(n12052), .ZN(n12053) );
  NAND2_X1 U15176 ( .A1(n12082), .A2(n12053), .ZN(n12749) );
  OAI21_X1 U15177 ( .B1(n12054), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n12076), .ZN(n20084) );
  INV_X1 U15178 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12056) );
  AOI21_X1 U15179 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n12056), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12057) );
  AOI21_X1 U15180 ( .B1(n12534), .B2(P1_EAX_REG_4__SCAN_IN), .A(n12057), .ZN(
        n12058) );
  OAI21_X1 U15181 ( .B1(n12975), .B2(n12059), .A(n12058), .ZN(n12060) );
  OAI21_X1 U15182 ( .B1(n20084), .B2(n12055), .A(n12060), .ZN(n12061) );
  OAI21_X1 U15183 ( .B1(n12749), .B2(n12220), .A(n12061), .ZN(n13439) );
  INV_X1 U15184 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12062) );
  OR2_X1 U15185 ( .A1(n12568), .A2(n12062), .ZN(n12074) );
  AOI22_X1 U15186 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15187 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15188 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15189 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12063) );
  NAND4_X1 U15190 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12072) );
  AOI22_X1 U15191 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15192 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15193 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12068) );
  INV_X1 U15194 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n20944) );
  AOI22_X1 U15195 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12067) );
  NAND4_X1 U15196 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12071) );
  NAND2_X1 U15197 ( .A1(n12585), .A2(n12768), .ZN(n12073) );
  NAND2_X1 U15198 ( .A1(n12074), .A2(n12073), .ZN(n12083) );
  XNOR2_X1 U15199 ( .A(n12082), .B(n12083), .ZN(n12754) );
  INV_X1 U15200 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12080) );
  NAND2_X1 U15201 ( .A1(n12076), .A2(n19956), .ZN(n12078) );
  NAND2_X1 U15202 ( .A1(n12078), .A2(n12097), .ZN(n19962) );
  AOI22_X1 U15203 ( .A1(n19962), .A2(n13611), .B1(n12820), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12079) );
  OAI21_X1 U15204 ( .B1(n11988), .B2(n12080), .A(n12079), .ZN(n12081) );
  INV_X1 U15205 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12084) );
  OR2_X1 U15206 ( .A1(n12568), .A2(n12084), .ZN(n12096) );
  AOI22_X1 U15207 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U15208 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15209 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15210 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12085) );
  NAND4_X1 U15211 ( .A1(n12088), .A2(n12087), .A3(n12086), .A4(n12085), .ZN(
        n12094) );
  AOI22_X1 U15212 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15213 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15214 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U15215 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12089) );
  NAND4_X1 U15216 ( .A1(n12092), .A2(n12091), .A3(n12090), .A4(n12089), .ZN(
        n12093) );
  NAND2_X1 U15217 ( .A1(n12585), .A2(n12778), .ZN(n12095) );
  NAND2_X1 U15218 ( .A1(n12106), .A2(n12105), .ZN(n12766) );
  NAND2_X1 U15219 ( .A1(n12766), .A2(n12231), .ZN(n12104) );
  INV_X1 U15220 ( .A(n12097), .ZN(n12099) );
  INV_X1 U15221 ( .A(n12110), .ZN(n12098) );
  OAI21_X1 U15222 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12099), .A(
        n12098), .ZN(n19953) );
  NAND2_X1 U15223 ( .A1(n19953), .A2(n13611), .ZN(n12100) );
  OAI21_X1 U15224 ( .B1(n12101), .B2(n12273), .A(n12100), .ZN(n12102) );
  AOI21_X1 U15225 ( .B1(n12534), .B2(P1_EAX_REG_6__SCAN_IN), .A(n12102), .ZN(
        n12103) );
  NAND2_X1 U15226 ( .A1(n13499), .A2(n13498), .ZN(n13504) );
  INV_X1 U15227 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12108) );
  NAND2_X1 U15228 ( .A1(n12585), .A2(n12780), .ZN(n12107) );
  OAI21_X1 U15229 ( .B1(n12568), .B2(n12108), .A(n12107), .ZN(n12109) );
  INV_X1 U15230 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12112) );
  OAI21_X1 U15231 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12110), .A(
        n12126), .ZN(n19939) );
  AOI22_X1 U15232 ( .A1(n13611), .A2(n19939), .B1(n12820), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12111) );
  OAI21_X1 U15233 ( .B1(n11988), .B2(n12112), .A(n12111), .ZN(n12113) );
  AOI21_X1 U15234 ( .B1(n12776), .B2(n12231), .A(n12113), .ZN(n13503) );
  AOI22_X1 U15235 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15236 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15237 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15238 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12116) );
  NAND4_X1 U15239 ( .A1(n12119), .A2(n12118), .A3(n12117), .A4(n12116), .ZN(
        n12125) );
  AOI22_X1 U15240 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12522), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15241 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12122) );
  AOI22_X1 U15242 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15243 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12120) );
  NAND4_X1 U15244 ( .A1(n12123), .A2(n12122), .A3(n12121), .A4(n12120), .ZN(
        n12124) );
  OAI21_X1 U15245 ( .B1(n12125), .B2(n12124), .A(n12231), .ZN(n12129) );
  XNOR2_X1 U15246 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12131), .ZN(
        n13741) );
  AOI22_X1 U15247 ( .A1(n13611), .A2(n13741), .B1(n12820), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12128) );
  NAND2_X1 U15248 ( .A1(n12534), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12127) );
  XNOR2_X1 U15249 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12156), .ZN(
        n19916) );
  INV_X1 U15250 ( .A(n19916), .ZN(n13769) );
  AOI22_X1 U15251 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12522), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15252 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15253 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15254 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11960), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12132) );
  NAND4_X1 U15255 ( .A1(n12135), .A2(n12134), .A3(n12133), .A4(n12132), .ZN(
        n12141) );
  AOI22_X1 U15256 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15257 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12138) );
  AOI22_X1 U15258 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12137) );
  AOI22_X1 U15259 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12136) );
  NAND4_X1 U15260 ( .A1(n12139), .A2(n12138), .A3(n12137), .A4(n12136), .ZN(
        n12140) );
  OAI21_X1 U15261 ( .B1(n12141), .B2(n12140), .A(n12231), .ZN(n12144) );
  NAND2_X1 U15262 ( .A1(n12534), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12143) );
  NAND2_X1 U15263 ( .A1(n12820), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12142) );
  NAND3_X1 U15264 ( .A1(n12144), .A2(n12143), .A3(n12142), .ZN(n12145) );
  AOI21_X1 U15265 ( .B1(n13769), .B2(n13611), .A(n12145), .ZN(n13719) );
  AOI22_X1 U15266 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15267 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12522), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15268 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15269 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12146) );
  NAND4_X1 U15270 ( .A1(n12149), .A2(n12148), .A3(n12147), .A4(n12146), .ZN(
        n12155) );
  AOI22_X1 U15271 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15272 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15273 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15274 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12150) );
  NAND4_X1 U15275 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n12154) );
  NOR2_X1 U15276 ( .A1(n12155), .A2(n12154), .ZN(n12159) );
  XNOR2_X1 U15277 ( .A(n12160), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14751) );
  NAND2_X1 U15278 ( .A1(n14751), .A2(n13611), .ZN(n12158) );
  AOI22_X1 U15279 ( .A1(n12534), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12820), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12157) );
  OAI211_X1 U15280 ( .C1(n12159), .C2(n12220), .A(n12158), .B(n12157), .ZN(
        n13645) );
  INV_X1 U15281 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12163) );
  OAI21_X1 U15282 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12161), .A(
        n12191), .ZN(n15830) );
  NAND2_X1 U15283 ( .A1(n15830), .A2(n13611), .ZN(n12162) );
  OAI21_X1 U15284 ( .B1(n12163), .B2(n12273), .A(n12162), .ZN(n12164) );
  AOI21_X1 U15285 ( .B1(n12534), .B2(P1_EAX_REG_11__SCAN_IN), .A(n12164), .ZN(
        n13860) );
  INV_X1 U15286 ( .A(n13860), .ZN(n12165) );
  AOI22_X1 U15287 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15288 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15289 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11960), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15290 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12166) );
  NAND4_X1 U15291 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n12175) );
  AOI22_X1 U15292 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15293 ( .A1(n11893), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15294 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15295 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12170) );
  NAND4_X1 U15296 ( .A1(n12173), .A2(n12172), .A3(n12171), .A4(n12170), .ZN(
        n12174) );
  OR2_X1 U15297 ( .A1(n12175), .A2(n12174), .ZN(n12176) );
  NAND2_X1 U15298 ( .A1(n12231), .A2(n12176), .ZN(n15753) );
  XOR2_X1 U15299 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12217), .Z(
        n14740) );
  AOI22_X1 U15300 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15301 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15302 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15303 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12178) );
  NAND4_X1 U15304 ( .A1(n12181), .A2(n12180), .A3(n12179), .A4(n12178), .ZN(
        n12187) );
  AOI22_X1 U15305 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12522), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15306 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15307 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15308 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12182) );
  NAND4_X1 U15309 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        n12186) );
  OR2_X1 U15310 ( .A1(n12187), .A2(n12186), .ZN(n12188) );
  AOI22_X1 U15311 ( .A1(n12231), .A2(n12188), .B1(n12820), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12190) );
  NAND2_X1 U15312 ( .A1(n12534), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12189) );
  OAI211_X1 U15313 ( .C1(n14740), .C2(n12055), .A(n12190), .B(n12189), .ZN(
        n13863) );
  AOI21_X1 U15314 ( .B1(n21034), .B2(n12191), .A(n12217), .ZN(n15819) );
  OR2_X1 U15315 ( .A1(n15819), .A2(n12055), .ZN(n12206) );
  AOI22_X1 U15316 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11911), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15317 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11903), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15318 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9757), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15319 ( .A1(n11893), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12192) );
  NAND4_X1 U15320 ( .A1(n12195), .A2(n12194), .A3(n12193), .A4(n12192), .ZN(
        n12201) );
  AOI22_X1 U15321 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12522), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15322 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15323 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11902), .B1(
        n12515), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15324 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12498), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12196) );
  NAND4_X1 U15325 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12196), .ZN(
        n12200) );
  OAI21_X1 U15326 ( .B1(n12201), .B2(n12200), .A(n12231), .ZN(n12204) );
  NAND2_X1 U15327 ( .A1(n12534), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12203) );
  NAND2_X1 U15328 ( .A1(n12820), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12202) );
  AND3_X1 U15329 ( .A1(n12204), .A2(n12203), .A3(n12202), .ZN(n12205) );
  NAND2_X1 U15330 ( .A1(n12206), .A2(n12205), .ZN(n13889) );
  AOI22_X1 U15331 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15332 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15333 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15334 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12207) );
  NAND4_X1 U15335 ( .A1(n12210), .A2(n12209), .A3(n12208), .A4(n12207), .ZN(
        n12216) );
  AOI22_X1 U15336 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15337 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15338 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15339 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12211) );
  NAND4_X1 U15340 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n12215) );
  NOR2_X1 U15341 ( .A1(n12216), .A2(n12215), .ZN(n12221) );
  XNOR2_X1 U15342 ( .A(n12222), .B(n15730), .ZN(n15734) );
  NAND2_X1 U15343 ( .A1(n15734), .A2(n13611), .ZN(n12219) );
  AOI22_X1 U15344 ( .A1(n12534), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n12820), 
        .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12218) );
  OAI211_X1 U15345 ( .C1(n12221), .C2(n12220), .A(n12219), .B(n12218), .ZN(
        n13881) );
  XNOR2_X1 U15346 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12241), .ZN(
        n15809) );
  INV_X1 U15347 ( .A(n15809), .ZN(n12238) );
  AOI22_X1 U15348 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15349 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15350 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15351 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12223) );
  NAND4_X1 U15352 ( .A1(n12226), .A2(n12225), .A3(n12224), .A4(n12223), .ZN(
        n12233) );
  AOI22_X1 U15353 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12515), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15354 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15355 ( .A1(n11893), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15356 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12227) );
  NAND4_X1 U15357 ( .A1(n12230), .A2(n12229), .A3(n12228), .A4(n12227), .ZN(
        n12232) );
  OAI21_X1 U15358 ( .B1(n12233), .B2(n12232), .A(n12231), .ZN(n12236) );
  NAND2_X1 U15359 ( .A1(n12534), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12235) );
  NAND2_X1 U15360 ( .A1(n12820), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12234) );
  NAND3_X1 U15361 ( .A1(n12236), .A2(n12235), .A3(n12234), .ZN(n12237) );
  AOI21_X1 U15362 ( .B1(n12238), .B2(n13611), .A(n12237), .ZN(n13900) );
  INV_X1 U15363 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12242) );
  XNOR2_X1 U15364 ( .A(n12261), .B(n12242), .ZN(n14712) );
  NAND2_X1 U15365 ( .A1(n14712), .A2(n13611), .ZN(n12260) );
  AOI22_X1 U15366 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15367 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15368 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12493), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15369 ( .A1(n11893), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12244) );
  NAND4_X1 U15370 ( .A1(n12247), .A2(n12246), .A3(n12245), .A4(n12244), .ZN(
        n12256) );
  AOI22_X1 U15371 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15372 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12515), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15373 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12251) );
  AOI21_X1 U15374 ( .B1(n9756), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A(n13611), .ZN(n12249) );
  NAND2_X1 U15375 ( .A1(n12521), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12248) );
  AND2_X1 U15376 ( .A1(n12249), .A2(n12248), .ZN(n12250) );
  NAND4_X1 U15377 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12255) );
  NAND2_X1 U15378 ( .A1(n12509), .A2(n12055), .ZN(n12357) );
  OAI21_X1 U15379 ( .B1(n12256), .B2(n12255), .A(n12357), .ZN(n12258) );
  AOI22_X1 U15380 ( .A1(n12534), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11980), .ZN(n12257) );
  NAND2_X1 U15381 ( .A1(n12258), .A2(n12257), .ZN(n12259) );
  NAND2_X1 U15382 ( .A1(n12260), .A2(n12259), .ZN(n14452) );
  AOI21_X1 U15383 ( .B1(n20990), .B2(n12262), .A(n12306), .ZN(n15798) );
  OR2_X1 U15384 ( .A1(n15798), .A2(n12055), .ZN(n12277) );
  INV_X1 U15385 ( .A(n12509), .ZN(n12531) );
  AOI22_X1 U15386 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15387 ( .A1(n11965), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15388 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12264) );
  AOI22_X1 U15389 ( .A1(n11893), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12263) );
  NAND4_X1 U15390 ( .A1(n12266), .A2(n12265), .A3(n12264), .A4(n12263), .ZN(
        n12272) );
  AOI22_X1 U15391 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12522), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15392 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15393 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15394 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12267) );
  NAND4_X1 U15395 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n12271) );
  OR2_X1 U15396 ( .A1(n12272), .A2(n12271), .ZN(n12275) );
  INV_X1 U15397 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14610) );
  OAI22_X1 U15398 ( .A1(n11988), .A2(n14610), .B1(n12273), .B2(n20990), .ZN(
        n12274) );
  AOI21_X1 U15399 ( .B1(n12531), .B2(n12275), .A(n12274), .ZN(n12276) );
  NAND2_X1 U15400 ( .A1(n12277), .A2(n12276), .ZN(n14437) );
  AND2_X2 U15401 ( .A1(n14438), .A2(n14437), .ZN(n14547) );
  INV_X1 U15402 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15709) );
  XNOR2_X1 U15403 ( .A(n12306), .B(n15709), .ZN(n15711) );
  AOI22_X1 U15404 ( .A1(n12075), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11980), .ZN(n12291) );
  AOI22_X1 U15405 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12522), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15406 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15407 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15408 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12278) );
  NAND4_X1 U15409 ( .A1(n12281), .A2(n12280), .A3(n12279), .A4(n12278), .ZN(
        n12289) );
  AOI22_X1 U15410 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12287) );
  AOI21_X1 U15411 ( .B1(n12493), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n13611), .ZN(n12283) );
  NAND2_X1 U15412 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12282) );
  AND2_X1 U15413 ( .A1(n12283), .A2(n12282), .ZN(n12286) );
  AOI22_X1 U15414 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15415 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12284) );
  NAND4_X1 U15416 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12284), .ZN(
        n12288) );
  OAI21_X1 U15417 ( .B1(n12289), .B2(n12288), .A(n12357), .ZN(n12290) );
  AOI22_X1 U15418 ( .A1(n15711), .A2(n13611), .B1(n12291), .B2(n12290), .ZN(
        n14546) );
  AOI22_X1 U15419 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15420 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15421 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15422 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12292) );
  NAND4_X1 U15423 ( .A1(n12295), .A2(n12294), .A3(n12293), .A4(n12292), .ZN(
        n12301) );
  AOI22_X1 U15424 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15425 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15426 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15427 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12296) );
  NAND4_X1 U15428 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12300) );
  NOR2_X1 U15429 ( .A1(n12301), .A2(n12300), .ZN(n12305) );
  NAND2_X1 U15430 ( .A1(n11980), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12302) );
  NAND2_X1 U15431 ( .A1(n12055), .A2(n12302), .ZN(n12303) );
  AOI21_X1 U15432 ( .B1(n12534), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12303), .ZN(
        n12304) );
  OAI21_X1 U15433 ( .B1(n12509), .B2(n12305), .A(n12304), .ZN(n12309) );
  OAI21_X1 U15434 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12307), .A(
        n12340), .ZN(n15791) );
  OR2_X1 U15435 ( .A1(n12055), .A2(n15791), .ZN(n12308) );
  NAND2_X1 U15436 ( .A1(n12309), .A2(n12308), .ZN(n14542) );
  AOI22_X1 U15437 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n11903), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15438 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12515), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15439 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12311) );
  AOI22_X1 U15440 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12310) );
  NAND4_X1 U15441 ( .A1(n12313), .A2(n12312), .A3(n12311), .A4(n12310), .ZN(
        n12321) );
  AOI22_X1 U15442 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12522), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U15443 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12318) );
  AOI22_X1 U15444 ( .A1(n11911), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12317) );
  NAND2_X1 U15445 ( .A1(n12521), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12315) );
  NAND2_X1 U15446 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12314) );
  AND3_X1 U15447 ( .A1(n12315), .A2(n12314), .A3(n12055), .ZN(n12316) );
  NAND4_X1 U15448 ( .A1(n12319), .A2(n12318), .A3(n12317), .A4(n12316), .ZN(
        n12320) );
  OAI21_X1 U15449 ( .B1(n12321), .B2(n12320), .A(n12357), .ZN(n12323) );
  AOI22_X1 U15450 ( .A1(n12075), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11980), .ZN(n12322) );
  NAND2_X1 U15451 ( .A1(n12323), .A2(n12322), .ZN(n12325) );
  XNOR2_X1 U15452 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12340), .ZN(
        n14427) );
  NAND2_X1 U15453 ( .A1(n13611), .A2(n14427), .ZN(n12324) );
  AOI22_X1 U15454 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12522), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15455 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12515), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15456 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11965), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15457 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12326) );
  NAND4_X1 U15458 ( .A1(n12329), .A2(n12328), .A3(n12327), .A4(n12326), .ZN(
        n12335) );
  AOI22_X1 U15459 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15460 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U15461 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15462 ( .A1(n11893), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12330) );
  NAND4_X1 U15463 ( .A1(n12333), .A2(n12332), .A3(n12331), .A4(n12330), .ZN(
        n12334) );
  NOR2_X1 U15464 ( .A1(n12335), .A2(n12334), .ZN(n12339) );
  NAND2_X1 U15465 ( .A1(n11980), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12336) );
  NAND2_X1 U15466 ( .A1(n12055), .A2(n12336), .ZN(n12337) );
  AOI21_X1 U15467 ( .B1(n12534), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12337), .ZN(
        n12338) );
  OAI21_X1 U15468 ( .B1(n12509), .B2(n12339), .A(n12338), .ZN(n12343) );
  INV_X1 U15469 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14428) );
  OAI21_X1 U15470 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12341), .A(
        n12362), .ZN(n15780) );
  OR2_X1 U15471 ( .A1(n12055), .A2(n15780), .ZN(n12342) );
  NAND2_X1 U15472 ( .A1(n12343), .A2(n12342), .ZN(n14531) );
  AOI22_X1 U15473 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12349) );
  AOI22_X1 U15474 ( .A1(n11893), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12348) );
  NAND2_X1 U15475 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12345) );
  NAND2_X1 U15476 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n12344) );
  AND3_X1 U15477 ( .A1(n12345), .A2(n12344), .A3(n12055), .ZN(n12347) );
  AOI22_X1 U15478 ( .A1(n11959), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12346) );
  NAND4_X1 U15479 ( .A1(n12349), .A2(n12348), .A3(n12347), .A4(n12346), .ZN(
        n12355) );
  AOI22_X1 U15480 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11965), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15481 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15482 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15483 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12350) );
  NAND4_X1 U15484 ( .A1(n12353), .A2(n12352), .A3(n12351), .A4(n12350), .ZN(
        n12354) );
  OR2_X1 U15485 ( .A1(n12355), .A2(n12354), .ZN(n12356) );
  NAND2_X1 U15486 ( .A1(n12357), .A2(n12356), .ZN(n12360) );
  AOI22_X1 U15487 ( .A1(n12075), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n11980), .ZN(n12359) );
  XNOR2_X1 U15488 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n12362), .ZN(
        n15681) );
  INV_X1 U15489 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12361) );
  OR2_X1 U15490 ( .A1(n12363), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12364) );
  NAND2_X1 U15491 ( .A1(n12364), .A2(n12424), .ZN(n15777) );
  AOI22_X1 U15492 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U15493 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15494 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15495 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12365) );
  NAND4_X1 U15496 ( .A1(n12368), .A2(n12367), .A3(n12366), .A4(n12365), .ZN(
        n12374) );
  AOI22_X1 U15497 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15498 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15499 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15500 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12369) );
  NAND4_X1 U15501 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12373) );
  NOR2_X1 U15502 ( .A1(n12374), .A2(n12373), .ZN(n12389) );
  AOI22_X1 U15503 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U15504 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12377) );
  AOI22_X1 U15505 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12493), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15506 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12375) );
  NAND4_X1 U15507 ( .A1(n12378), .A2(n12377), .A3(n12376), .A4(n12375), .ZN(
        n12384) );
  AOI22_X1 U15508 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15509 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15510 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15511 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12379) );
  NAND4_X1 U15512 ( .A1(n12382), .A2(n12381), .A3(n12380), .A4(n12379), .ZN(
        n12383) );
  NOR2_X1 U15513 ( .A1(n12384), .A2(n12383), .ZN(n12390) );
  XNOR2_X1 U15514 ( .A(n12389), .B(n12390), .ZN(n12385) );
  NOR2_X1 U15515 ( .A1(n12509), .A2(n12385), .ZN(n12388) );
  INV_X1 U15516 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14593) );
  NAND2_X1 U15517 ( .A1(n11980), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12386) );
  OAI211_X1 U15518 ( .C1(n11988), .C2(n14593), .A(n12055), .B(n12386), .ZN(
        n12387) );
  OAI22_X1 U15519 ( .A1(n15777), .A2(n12055), .B1(n12388), .B2(n12387), .ZN(
        n14516) );
  NOR2_X2 U15520 ( .A1(n14513), .A2(n14516), .ZN(n14412) );
  NOR2_X1 U15521 ( .A1(n12390), .A2(n12389), .ZN(n12419) );
  AOI22_X1 U15522 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15523 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11892), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15524 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12392) );
  AOI22_X1 U15525 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12391) );
  NAND4_X1 U15526 ( .A1(n12394), .A2(n12393), .A3(n12392), .A4(n12391), .ZN(
        n12400) );
  AOI22_X1 U15527 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15528 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15529 ( .A1(n11902), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12396) );
  INV_X1 U15530 ( .A(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n21088) );
  AOI22_X1 U15531 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12395) );
  NAND4_X1 U15532 ( .A1(n12398), .A2(n12397), .A3(n12396), .A4(n12395), .ZN(
        n12399) );
  OR2_X1 U15533 ( .A1(n12400), .A2(n12399), .ZN(n12418) );
  XNOR2_X1 U15534 ( .A(n12419), .B(n12418), .ZN(n12404) );
  NAND2_X1 U15535 ( .A1(n11980), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12401) );
  NAND2_X1 U15536 ( .A1(n12055), .A2(n12401), .ZN(n12402) );
  AOI21_X1 U15537 ( .B1(n12534), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12402), .ZN(
        n12403) );
  OAI21_X1 U15538 ( .B1(n12404), .B2(n12509), .A(n12403), .ZN(n12406) );
  XNOR2_X1 U15539 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n12424), .ZN(
        n14416) );
  NAND2_X1 U15540 ( .A1(n13611), .A2(n14416), .ZN(n12405) );
  NAND2_X1 U15541 ( .A1(n12406), .A2(n12405), .ZN(n14414) );
  AOI22_X1 U15542 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15543 ( .A1(n11893), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15544 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U15545 ( .A1(n11892), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12408) );
  NAND4_X1 U15546 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12417) );
  AOI22_X1 U15547 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15548 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11902), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15549 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15550 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12412) );
  NAND4_X1 U15551 ( .A1(n12415), .A2(n12414), .A3(n12413), .A4(n12412), .ZN(
        n12416) );
  NOR2_X1 U15552 ( .A1(n12417), .A2(n12416), .ZN(n12433) );
  NAND2_X1 U15553 ( .A1(n12419), .A2(n12418), .ZN(n12432) );
  XNOR2_X1 U15554 ( .A(n12433), .B(n12432), .ZN(n12423) );
  NAND2_X1 U15555 ( .A1(n11980), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12420) );
  NAND2_X1 U15556 ( .A1(n12055), .A2(n12420), .ZN(n12421) );
  AOI21_X1 U15557 ( .B1(n12534), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12421), .ZN(
        n12422) );
  OAI21_X1 U15558 ( .B1(n12423), .B2(n12509), .A(n12422), .ZN(n12431) );
  INV_X1 U15559 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12428) );
  INV_X1 U15560 ( .A(n12426), .ZN(n12427) );
  NAND2_X1 U15561 ( .A1(n12428), .A2(n12427), .ZN(n12429) );
  NAND2_X1 U15562 ( .A1(n12451), .A2(n12429), .ZN(n15672) );
  NOR2_X1 U15563 ( .A1(n12433), .A2(n12432), .ZN(n12467) );
  AOI22_X1 U15564 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15565 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12436) );
  AOI22_X1 U15566 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15567 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12434) );
  NAND4_X1 U15568 ( .A1(n12437), .A2(n12436), .A3(n12435), .A4(n12434), .ZN(
        n12443) );
  AOI22_X1 U15569 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U15570 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U15571 ( .A1(n11965), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15572 ( .A1(n11903), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12438) );
  NAND4_X1 U15573 ( .A1(n12441), .A2(n12440), .A3(n12439), .A4(n12438), .ZN(
        n12442) );
  OR2_X1 U15574 ( .A1(n12443), .A2(n12442), .ZN(n12466) );
  INV_X1 U15575 ( .A(n12466), .ZN(n12444) );
  XNOR2_X1 U15576 ( .A(n12467), .B(n12444), .ZN(n12445) );
  NAND2_X1 U15577 ( .A1(n12445), .A2(n12531), .ZN(n12450) );
  NAND2_X1 U15578 ( .A1(n11980), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12446) );
  NAND2_X1 U15579 ( .A1(n12055), .A2(n12446), .ZN(n12447) );
  AOI21_X1 U15580 ( .B1(n12534), .B2(P1_EAX_REG_26__SCAN_IN), .A(n12447), .ZN(
        n12449) );
  XNOR2_X1 U15581 ( .A(n12451), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15655) );
  INV_X1 U15582 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15650) );
  INV_X1 U15583 ( .A(n12452), .ZN(n12454) );
  INV_X1 U15584 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12453) );
  NAND2_X1 U15585 ( .A1(n12454), .A2(n12453), .ZN(n12455) );
  NAND2_X1 U15586 ( .A1(n12488), .A2(n12455), .ZN(n14657) );
  AOI22_X1 U15587 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12522), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U15588 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11959), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15589 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12457) );
  AOI22_X1 U15590 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12015), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12456) );
  NAND4_X1 U15591 ( .A1(n12459), .A2(n12458), .A3(n12457), .A4(n12456), .ZN(
        n12465) );
  AOI22_X1 U15592 ( .A1(n11900), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12498), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15593 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12515), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15594 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11965), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12461) );
  AOI22_X1 U15595 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12460) );
  NAND4_X1 U15596 ( .A1(n12463), .A2(n12462), .A3(n12461), .A4(n12460), .ZN(
        n12464) );
  NOR2_X1 U15597 ( .A1(n12465), .A2(n12464), .ZN(n12483) );
  NAND2_X1 U15598 ( .A1(n12467), .A2(n12466), .ZN(n12482) );
  XNOR2_X1 U15599 ( .A(n12483), .B(n12482), .ZN(n12470) );
  AOI21_X1 U15600 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n11980), .A(
        n13611), .ZN(n12469) );
  NAND2_X1 U15601 ( .A1(n12075), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12468) );
  OAI211_X1 U15602 ( .C1(n12470), .C2(n12509), .A(n12469), .B(n12468), .ZN(
        n12471) );
  AOI22_X1 U15603 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11899), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15604 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U15605 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15606 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12472) );
  NAND4_X1 U15607 ( .A1(n12475), .A2(n12474), .A3(n12473), .A4(n12472), .ZN(
        n12481) );
  AOI22_X1 U15608 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11893), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U15609 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11911), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15610 ( .A1(n11965), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12243), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15611 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12476) );
  NAND4_X1 U15612 ( .A1(n12479), .A2(n12478), .A3(n12477), .A4(n12476), .ZN(
        n12480) );
  OR2_X1 U15613 ( .A1(n12481), .A2(n12480), .ZN(n12505) );
  NOR2_X1 U15614 ( .A1(n12483), .A2(n12482), .ZN(n12506) );
  XOR2_X1 U15615 ( .A(n12505), .B(n12506), .Z(n12484) );
  NAND2_X1 U15616 ( .A1(n12484), .A2(n12531), .ZN(n12487) );
  INV_X1 U15617 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14639) );
  AOI21_X1 U15618 ( .B1(n14639), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12485) );
  AOI21_X1 U15619 ( .B1(n12534), .B2(P1_EAX_REG_28__SCAN_IN), .A(n12485), .ZN(
        n12486) );
  XNOR2_X1 U15620 ( .A(n12488), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14641) );
  AOI22_X1 U15621 ( .A1(n12487), .A2(n12486), .B1(n13611), .B2(n14641), .ZN(
        n14389) );
  INV_X1 U15622 ( .A(n12488), .ZN(n12489) );
  INV_X1 U15623 ( .A(n12490), .ZN(n12491) );
  INV_X1 U15624 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14381) );
  NAND2_X1 U15625 ( .A1(n12491), .A2(n14381), .ZN(n12492) );
  NAND2_X1 U15626 ( .A1(n12829), .A2(n12492), .ZN(n14634) );
  AOI22_X1 U15627 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12497) );
  AOI22_X1 U15628 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U15629 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12495) );
  AOI22_X1 U15630 ( .A1(n12493), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12494) );
  NAND4_X1 U15631 ( .A1(n12497), .A2(n12496), .A3(n12495), .A4(n12494), .ZN(
        n12504) );
  AOI22_X1 U15632 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12522), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12502) );
  AOI22_X1 U15633 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11965), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12501) );
  AOI22_X1 U15634 ( .A1(n12498), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12500) );
  AOI22_X1 U15635 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12499) );
  NAND4_X1 U15636 ( .A1(n12502), .A2(n12501), .A3(n12500), .A4(n12499), .ZN(
        n12503) );
  NOR2_X1 U15637 ( .A1(n12504), .A2(n12503), .ZN(n12513) );
  NAND2_X1 U15638 ( .A1(n12506), .A2(n12505), .ZN(n12512) );
  XNOR2_X1 U15639 ( .A(n12513), .B(n12512), .ZN(n12510) );
  AOI21_X1 U15640 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n11980), .A(
        n13611), .ZN(n12508) );
  NAND2_X1 U15641 ( .A1(n12075), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12507) );
  OAI211_X1 U15642 ( .C1(n12510), .C2(n12509), .A(n12508), .B(n12507), .ZN(
        n12511) );
  NOR2_X2 U15643 ( .A1(n14376), .A2(n14378), .ZN(n12819) );
  NOR2_X1 U15644 ( .A1(n12513), .A2(n12512), .ZN(n12530) );
  AOI22_X1 U15645 ( .A1(n11899), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12519) );
  AOI22_X1 U15646 ( .A1(n11891), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11959), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U15647 ( .A1(n12015), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11965), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U15648 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11916), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12516) );
  NAND4_X1 U15649 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12528) );
  AOI22_X1 U15650 ( .A1(n12520), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11901), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12526) );
  AOI22_X1 U15651 ( .A1(n12243), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12521), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U15652 ( .A1(n11910), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9756), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U15653 ( .A1(n12522), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13351), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12523) );
  NAND4_X1 U15654 ( .A1(n12526), .A2(n12525), .A3(n12524), .A4(n12523), .ZN(
        n12527) );
  NOR2_X1 U15655 ( .A1(n12528), .A2(n12527), .ZN(n12529) );
  XNOR2_X1 U15656 ( .A(n12530), .B(n12529), .ZN(n12532) );
  NAND2_X1 U15657 ( .A1(n12532), .A2(n12531), .ZN(n12536) );
  INV_X1 U15658 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14623) );
  NOR2_X1 U15659 ( .A1(n14623), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12533) );
  AOI211_X1 U15660 ( .C1(n12534), .C2(P1_EAX_REG_30__SCAN_IN), .A(n12533), .B(
        n13611), .ZN(n12535) );
  XNOR2_X1 U15661 ( .A(n12829), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14625) );
  AOI22_X1 U15662 ( .A1(n12536), .A2(n12535), .B1(n14625), .B2(n13611), .ZN(
        n12818) );
  NAND2_X1 U15663 ( .A1(n11853), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12537) );
  NAND2_X1 U15664 ( .A1(n12538), .A2(n12537), .ZN(n12554) );
  MUX2_X1 U15665 ( .A(n12539), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n11952), .Z(n12563) );
  XNOR2_X1 U15666 ( .A(n12543), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12574) );
  AOI222_X1 U15667 ( .A1(n12544), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n12544), .B2(n12975), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n12975), .ZN(n12842) );
  NOR2_X1 U15668 ( .A1(n20176), .A2(n20708), .ZN(n12546) );
  AOI21_X1 U15669 ( .B1(n12585), .B2(n20155), .A(n12546), .ZN(n12559) );
  NAND2_X1 U15670 ( .A1(n12559), .A2(n20155), .ZN(n12580) );
  INV_X1 U15671 ( .A(n12585), .ZN(n12547) );
  OAI21_X1 U15672 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20568), .A(
        n12555), .ZN(n12549) );
  NOR2_X1 U15673 ( .A1(n12547), .A2(n12549), .ZN(n12553) );
  OR2_X1 U15674 ( .A1(n20176), .A2(n20144), .ZN(n12548) );
  NAND2_X1 U15675 ( .A1(n12548), .A2(n12606), .ZN(n12576) );
  INV_X1 U15676 ( .A(n12549), .ZN(n12550) );
  OAI211_X1 U15677 ( .C1(n12551), .C2(n20144), .A(n12576), .B(n12550), .ZN(
        n12552) );
  OAI21_X1 U15678 ( .B1(n12553), .B2(n12586), .A(n12552), .ZN(n12561) );
  INV_X1 U15679 ( .A(n12554), .ZN(n12558) );
  INV_X1 U15680 ( .A(n12555), .ZN(n12557) );
  OAI21_X1 U15681 ( .B1(n12558), .B2(n12557), .A(n12556), .ZN(n12839) );
  OAI211_X1 U15682 ( .C1(n12561), .C2(n12559), .A(n12839), .B(n12580), .ZN(
        n12571) );
  INV_X1 U15683 ( .A(n12559), .ZN(n12560) );
  NOR2_X1 U15684 ( .A1(n12839), .A2(n12560), .ZN(n12562) );
  NAND2_X1 U15685 ( .A1(n12562), .A2(n12561), .ZN(n12570) );
  NAND2_X1 U15686 ( .A1(n12564), .A2(n12563), .ZN(n12566) );
  NAND2_X1 U15687 ( .A1(n12566), .A2(n12565), .ZN(n12838) );
  INV_X1 U15688 ( .A(n12838), .ZN(n12567) );
  NAND2_X1 U15689 ( .A1(n12585), .A2(n12567), .ZN(n12575) );
  OAI211_X1 U15690 ( .C1(n12568), .C2(n12567), .A(n12576), .B(n12575), .ZN(
        n12569) );
  AOI21_X1 U15691 ( .B1(n12574), .B2(n12573), .A(n12572), .ZN(n12837) );
  INV_X1 U15692 ( .A(n12786), .ZN(n12740) );
  OAI22_X1 U15693 ( .A1(n12837), .A2(n12740), .B1(n12576), .B2(n12575), .ZN(
        n12577) );
  OAI22_X1 U15694 ( .A1(n12578), .A2(n12577), .B1(n12582), .B2(n12837), .ZN(
        n12579) );
  OAI21_X1 U15695 ( .B1(n12841), .B2(n12580), .A(n12579), .ZN(n12581) );
  OAI21_X1 U15696 ( .B1(n12582), .B2(n12841), .A(n12581), .ZN(n12583) );
  OAI21_X1 U15697 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n12975), .A(n12583), 
        .ZN(n12584) );
  AOI21_X1 U15698 ( .B1(n12585), .B2(n12842), .A(n12584), .ZN(n12588) );
  AND2_X1 U15699 ( .A1(n12842), .A2(n12586), .ZN(n12587) );
  INV_X1 U15700 ( .A(n13145), .ZN(n12600) );
  NOR2_X1 U15701 ( .A1(n12817), .A2(n14474), .ZN(n13139) );
  NOR2_X1 U15702 ( .A1(n13139), .A2(n12589), .ZN(n12590) );
  AND2_X1 U15703 ( .A1(n12590), .A2(n20176), .ZN(n12599) );
  AND2_X1 U15704 ( .A1(n11978), .A2(n20171), .ZN(n12592) );
  OAI21_X1 U15705 ( .B1(n12817), .B2(n12592), .A(n20188), .ZN(n12594) );
  NAND2_X1 U15706 ( .A1(n12594), .A2(n12593), .ZN(n12596) );
  NAND2_X1 U15707 ( .A1(n12596), .A2(n12595), .ZN(n12598) );
  NAND2_X1 U15708 ( .A1(n12598), .A2(n12597), .ZN(n13143) );
  NAND4_X1 U15709 ( .A1(n12600), .A2(n12599), .A3(n12591), .A4(n13143), .ZN(
        n14882) );
  NAND2_X1 U15710 ( .A1(n12593), .A2(n9740), .ZN(n12601) );
  NOR2_X1 U15711 ( .A1(n14351), .A2(n14343), .ZN(n12959) );
  OR2_X1 U15712 ( .A1(n15568), .A2(n20708), .ZN(n19894) );
  NAND2_X1 U15713 ( .A1(n12959), .A2(n13129), .ZN(n12608) );
  INV_X1 U15714 ( .A(n12602), .ZN(n12605) );
  INV_X1 U15715 ( .A(n20188), .ZN(n14345) );
  AND3_X1 U15716 ( .A1(n14345), .A2(n20171), .A3(n13129), .ZN(n12604) );
  AND3_X1 U15717 ( .A1(n12605), .A2(n12604), .A3(n12603), .ZN(n12846) );
  INV_X1 U15718 ( .A(n12610), .ZN(n13162) );
  NAND2_X1 U15719 ( .A1(n12846), .A2(n13162), .ZN(n12607) );
  NAND2_X2 U15720 ( .A1(n20012), .A2(n20188), .ZN(n14561) );
  NOR2_X4 U15721 ( .A1(n12610), .A2(n12619), .ZN(n12695) );
  INV_X1 U15722 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n14483) );
  NAND2_X1 U15723 ( .A1(n12695), .A2(n14483), .ZN(n12613) );
  INV_X1 U15724 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20135) );
  NAND2_X1 U15725 ( .A1(n13141), .A2(n20135), .ZN(n12611) );
  OAI211_X1 U15726 ( .C1(n12610), .C2(P1_EBX_REG_1__SCAN_IN), .A(n12611), .B(
        n12619), .ZN(n12612) );
  NAND2_X1 U15727 ( .A1(n13141), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12615) );
  INV_X1 U15728 ( .A(n12609), .ZN(n12688) );
  INV_X1 U15729 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13100) );
  NAND2_X1 U15730 ( .A1(n12688), .A2(n13100), .ZN(n12614) );
  NAND2_X1 U15731 ( .A1(n12615), .A2(n12614), .ZN(n13097) );
  INV_X1 U15732 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13341) );
  NAND2_X1 U15733 ( .A1(n12695), .A2(n13341), .ZN(n12618) );
  INV_X1 U15734 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20120) );
  NAND2_X1 U15735 ( .A1(n13141), .A2(n20120), .ZN(n12616) );
  OAI211_X1 U15736 ( .C1(n12610), .C2(P1_EBX_REG_2__SCAN_IN), .A(n12616), .B(
        n12619), .ZN(n12617) );
  AND2_X1 U15737 ( .A1(n12618), .A2(n12617), .ZN(n13338) );
  MUX2_X1 U15738 ( .A(n12692), .B(n12609), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12621) );
  NOR2_X1 U15739 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12620) );
  NOR2_X1 U15740 ( .A1(n12621), .A2(n12620), .ZN(n13405) );
  NAND2_X1 U15741 ( .A1(n13406), .A2(n13405), .ZN(n13444) );
  MUX2_X1 U15742 ( .A(n12695), .B(n12670), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12623) );
  INV_X1 U15743 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20092) );
  OAI21_X1 U15744 ( .B1(n13162), .B2(n20092), .A(n12673), .ZN(n12622) );
  NOR2_X1 U15745 ( .A1(n12623), .A2(n12622), .ZN(n13445) );
  INV_X1 U15746 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20011) );
  NAND2_X1 U15747 ( .A1(n12692), .A2(n20011), .ZN(n12626) );
  NAND2_X1 U15748 ( .A1(n12688), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12624) );
  OAI211_X1 U15749 ( .C1(n12610), .C2(P1_EBX_REG_5__SCAN_IN), .A(n13141), .B(
        n12624), .ZN(n12625) );
  MUX2_X1 U15750 ( .A(n12695), .B(n12670), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12629) );
  NAND2_X1 U15751 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12610), .ZN(
        n12627) );
  NAND2_X1 U15752 ( .A1(n12673), .A2(n12627), .ZN(n12628) );
  NOR2_X1 U15753 ( .A1(n12629), .A2(n12628), .ZN(n13500) );
  INV_X1 U15754 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13510) );
  NAND2_X1 U15755 ( .A1(n12692), .A2(n13510), .ZN(n12632) );
  NAND2_X1 U15756 ( .A1(n12688), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12630) );
  OAI211_X1 U15757 ( .C1(n12610), .C2(P1_EBX_REG_7__SCAN_IN), .A(n13141), .B(
        n12630), .ZN(n12631) );
  NAND2_X1 U15758 ( .A1(n13508), .A2(n13507), .ZN(n13506) );
  MUX2_X1 U15759 ( .A(n12695), .B(n12670), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12635) );
  NAND2_X1 U15760 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n12610), .ZN(
        n12633) );
  NAND2_X1 U15761 ( .A1(n12673), .A2(n12633), .ZN(n12634) );
  NOR2_X1 U15762 ( .A1(n12635), .A2(n12634), .ZN(n13621) );
  INV_X1 U15763 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20005) );
  NAND2_X1 U15764 ( .A1(n12692), .A2(n20005), .ZN(n12638) );
  NAND2_X1 U15765 ( .A1(n12688), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12636) );
  OAI211_X1 U15766 ( .C1(n12610), .C2(P1_EBX_REG_9__SCAN_IN), .A(n13141), .B(
        n12636), .ZN(n12637) );
  NAND2_X1 U15767 ( .A1(n12638), .A2(n12637), .ZN(n15934) );
  INV_X1 U15768 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13729) );
  NAND2_X1 U15769 ( .A1(n12695), .A2(n13729), .ZN(n12641) );
  INV_X1 U15770 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14747) );
  NAND2_X1 U15771 ( .A1(n13141), .A2(n14747), .ZN(n12639) );
  OAI211_X1 U15772 ( .C1(n12610), .C2(P1_EBX_REG_10__SCAN_IN), .A(n12639), .B(
        n12688), .ZN(n12640) );
  MUX2_X1 U15773 ( .A(n12692), .B(n12609), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12643) );
  NOR2_X1 U15774 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12642) );
  NOR2_X1 U15775 ( .A1(n12643), .A2(n12642), .ZN(n15757) );
  MUX2_X1 U15776 ( .A(n12695), .B(n12670), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12644) );
  INV_X1 U15777 ( .A(n12644), .ZN(n12647) );
  NAND2_X1 U15778 ( .A1(n12610), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12645) );
  AND2_X1 U15779 ( .A1(n12673), .A2(n12645), .ZN(n12646) );
  NAND2_X1 U15780 ( .A1(n12647), .A2(n12646), .ZN(n13886) );
  MUX2_X1 U15781 ( .A(n12692), .B(n12609), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12648) );
  INV_X1 U15782 ( .A(n12648), .ZN(n12650) );
  INV_X1 U15783 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15899) );
  NAND2_X1 U15784 ( .A1(n13096), .A2(n15899), .ZN(n12649) );
  NAND2_X1 U15785 ( .A1(n12650), .A2(n12649), .ZN(n13875) );
  MUX2_X1 U15786 ( .A(n12695), .B(n12670), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12653) );
  NAND2_X1 U15787 ( .A1(n12610), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12651) );
  NAND2_X1 U15788 ( .A1(n12673), .A2(n12651), .ZN(n12652) );
  NOR2_X1 U15789 ( .A1(n12653), .A2(n12652), .ZN(n13894) );
  MUX2_X1 U15790 ( .A(n12692), .B(n12609), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12655) );
  NOR2_X1 U15791 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12654) );
  NOR2_X1 U15792 ( .A1(n12655), .A2(n12654), .ZN(n14558) );
  MUX2_X1 U15793 ( .A(n12695), .B(n12670), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n12658) );
  NAND2_X1 U15794 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n12610), .ZN(
        n12656) );
  NAND2_X1 U15795 ( .A1(n12673), .A2(n12656), .ZN(n12657) );
  NOR2_X1 U15796 ( .A1(n12658), .A2(n12657), .ZN(n14456) );
  MUX2_X1 U15797 ( .A(n12692), .B(n12609), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12659) );
  INV_X1 U15798 ( .A(n12659), .ZN(n12661) );
  NAND2_X1 U15799 ( .A1(n13096), .A2(n12801), .ZN(n12660) );
  NAND2_X1 U15800 ( .A1(n12661), .A2(n12660), .ZN(n14442) );
  INV_X1 U15801 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15714) );
  NAND2_X1 U15802 ( .A1(n12695), .A2(n15714), .ZN(n12665) );
  INV_X1 U15803 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12662) );
  NAND2_X1 U15804 ( .A1(n13141), .A2(n12662), .ZN(n12663) );
  OAI211_X1 U15805 ( .C1(n12610), .C2(P1_EBX_REG_18__SCAN_IN), .A(n12663), .B(
        n12688), .ZN(n12664) );
  MUX2_X1 U15806 ( .A(n12692), .B(n12609), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12667) );
  NOR2_X1 U15807 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12666) );
  NOR2_X1 U15808 ( .A1(n12667), .A2(n12666), .ZN(n14539) );
  AND2_X2 U15809 ( .A1(n14552), .A2(n14539), .ZN(n14541) );
  MUX2_X1 U15810 ( .A(n12692), .B(n12609), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12669) );
  NOR2_X1 U15811 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12668) );
  NOR2_X1 U15812 ( .A1(n12669), .A2(n12668), .ZN(n14533) );
  MUX2_X1 U15813 ( .A(n12695), .B(n12670), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12671) );
  INV_X1 U15814 ( .A(n12671), .ZN(n12675) );
  NAND2_X1 U15815 ( .A1(n12610), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12672) );
  AND2_X1 U15816 ( .A1(n12673), .A2(n12672), .ZN(n12674) );
  NAND2_X1 U15817 ( .A1(n12675), .A2(n12674), .ZN(n14534) );
  AND2_X1 U15818 ( .A1(n14533), .A2(n14534), .ZN(n12676) );
  NAND2_X1 U15819 ( .A1(n12695), .A2(n15683), .ZN(n12679) );
  INV_X1 U15820 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14687) );
  NAND2_X1 U15821 ( .A1(n13141), .A2(n14687), .ZN(n12677) );
  OAI211_X1 U15822 ( .C1(n12610), .C2(P1_EBX_REG_22__SCAN_IN), .A(n12677), .B(
        n12688), .ZN(n12678) );
  NAND2_X1 U15823 ( .A1(n12679), .A2(n12678), .ZN(n14526) );
  MUX2_X1 U15824 ( .A(n12692), .B(n12609), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12680) );
  INV_X1 U15825 ( .A(n12680), .ZN(n12682) );
  INV_X1 U15826 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15864) );
  NAND2_X1 U15827 ( .A1(n13096), .A2(n15864), .ZN(n12681) );
  NAND2_X1 U15828 ( .A1(n12682), .A2(n12681), .ZN(n14517) );
  MUX2_X1 U15829 ( .A(n12692), .B(n12609), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12684) );
  NOR2_X1 U15830 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12683) );
  NOR2_X1 U15831 ( .A1(n12684), .A2(n12683), .ZN(n14505) );
  INV_X1 U15832 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14415) );
  NAND2_X1 U15833 ( .A1(n12695), .A2(n14415), .ZN(n12687) );
  INV_X1 U15834 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15851) );
  NAND2_X1 U15835 ( .A1(n13141), .A2(n15851), .ZN(n12685) );
  OAI211_X1 U15836 ( .C1(n12610), .C2(P1_EBX_REG_24__SCAN_IN), .A(n12685), .B(
        n12688), .ZN(n12686) );
  NAND2_X1 U15837 ( .A1(n12687), .A2(n12686), .ZN(n14506) );
  INV_X1 U15838 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15651) );
  NAND2_X1 U15839 ( .A1(n12695), .A2(n15651), .ZN(n12691) );
  INV_X1 U15840 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14824) );
  NAND2_X1 U15841 ( .A1(n13141), .A2(n14824), .ZN(n12689) );
  OAI211_X1 U15842 ( .C1(n12610), .C2(P1_EBX_REG_26__SCAN_IN), .A(n12689), .B(
        n12688), .ZN(n12690) );
  NAND2_X1 U15843 ( .A1(n12691), .A2(n12690), .ZN(n14500) );
  AND2_X2 U15844 ( .A1(n14508), .A2(n14500), .ZN(n14502) );
  MUX2_X1 U15845 ( .A(n12692), .B(n12609), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12694) );
  NOR2_X1 U15846 ( .A1(n14354), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12693) );
  NOR2_X1 U15847 ( .A1(n12694), .A2(n12693), .ZN(n14401) );
  INV_X1 U15848 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14493) );
  NAND2_X1 U15849 ( .A1(n12695), .A2(n14493), .ZN(n12699) );
  INV_X1 U15850 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12696) );
  NAND2_X1 U15851 ( .A1(n13141), .A2(n12696), .ZN(n12697) );
  OAI211_X1 U15852 ( .C1(n12610), .C2(P1_EBX_REG_28__SCAN_IN), .A(n12697), .B(
        n12688), .ZN(n12698) );
  AND2_X1 U15853 ( .A1(n12699), .A2(n12698), .ZN(n14391) );
  INV_X1 U15854 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n12700) );
  NAND2_X1 U15855 ( .A1(n13162), .A2(n12700), .ZN(n12701) );
  OAI21_X1 U15856 ( .B1(n14354), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n12701), .ZN(n12702) );
  MUX2_X1 U15857 ( .A(n12702), .B(n12701), .S(n12609), .Z(n14380) );
  OAI22_X1 U15858 ( .A1(n14379), .A2(n12688), .B1(n12702), .B2(n14393), .ZN(
        n12704) );
  AOI22_X1 U15859 ( .A1(n14354), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12610), .ZN(n14353) );
  INV_X1 U15860 ( .A(n14353), .ZN(n12703) );
  XNOR2_X1 U15861 ( .A(n12704), .B(n12703), .ZN(n14780) );
  INV_X1 U15862 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14370) );
  OAI21_X1 U15863 ( .B1(n14780), .B2(n20001), .A(n10229), .ZN(n12705) );
  INV_X1 U15864 ( .A(n12705), .ZN(n12706) );
  NOR2_X1 U15865 ( .A1(n12708), .A2(n12707), .ZN(n18650) );
  NAND2_X1 U15866 ( .A1(n12709), .A2(n17766), .ZN(n12723) );
  NAND2_X1 U15867 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18189) );
  NAND2_X1 U15868 ( .A1(n18810), .A2(n18189), .ZN(n18861) );
  NAND2_X1 U15869 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17822) );
  NAND3_X1 U15870 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17718) );
  NAND2_X1 U15871 ( .A1(n16753), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16647) );
  NAND2_X1 U15872 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17655) );
  INV_X1 U15873 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17635) );
  INV_X1 U15874 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16654) );
  NAND2_X1 U15875 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17586) );
  NAND2_X1 U15876 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17545) );
  NAND2_X1 U15877 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17533), .ZN(
        n17513) );
  NAND2_X1 U15878 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17514) );
  NAND2_X1 U15879 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n12713), .ZN(
        n12714) );
  INV_X1 U15880 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17848) );
  NAND2_X1 U15881 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16374), .ZN(
        n12711) );
  INV_X1 U15882 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18856) );
  NOR2_X1 U15883 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18856), .ZN(n17689) );
  NAND2_X1 U15884 ( .A1(n17857), .A2(n18856), .ZN(n18858) );
  AOI21_X1 U15885 ( .B1(n18189), .B2(n18858), .A(n18835), .ZN(n18201) );
  INV_X2 U15886 ( .A(n18356), .ZN(n18241) );
  OR2_X1 U15887 ( .A1(n12714), .A2(n17691), .ZN(n16367) );
  INV_X1 U15888 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16534) );
  XOR2_X1 U15889 ( .A(n16534), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12715) );
  NOR2_X1 U15890 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17607), .ZN(
        n16376) );
  INV_X1 U15891 ( .A(n12713), .ZN(n16379) );
  NOR2_X1 U15892 ( .A1(n16379), .A2(n17848), .ZN(n16514) );
  INV_X1 U15893 ( .A(n17689), .ZN(n17856) );
  NAND2_X1 U15894 ( .A1(n18241), .A2(n12714), .ZN(n16380) );
  OAI211_X1 U15895 ( .C1(n16514), .C2(n17856), .A(n16380), .B(n17855), .ZN(
        n16385) );
  NOR2_X1 U15896 ( .A1(n16376), .A2(n16385), .ZN(n16366) );
  OAI22_X1 U15897 ( .A1(n16367), .A2(n12715), .B1(n16366), .B2(n16534), .ZN(
        n12716) );
  AOI211_X1 U15898 ( .C1(n17708), .C2(n16525), .A(n12717), .B(n12716), .ZN(
        n12722) );
  NAND2_X1 U15899 ( .A1(n12718), .A2(n17767), .ZN(n12721) );
  NAND2_X1 U15900 ( .A1(n12731), .A2(n12730), .ZN(n12742) );
  XNOR2_X1 U15901 ( .A(n12742), .B(n12741), .ZN(n12724) );
  AOI21_X1 U15902 ( .B1(n12724), .B2(n13117), .A(n12726), .ZN(n12725) );
  AOI21_X1 U15903 ( .B1(n13117), .B2(n12727), .A(n12726), .ZN(n12728) );
  OAI211_X1 U15904 ( .C1(n12731), .C2(n12730), .A(n13117), .B(n12742), .ZN(
        n12732) );
  OAI211_X1 U15905 ( .C1(n12734), .C2(n12606), .A(n12733), .B(n12732), .ZN(
        n12735) );
  XNOR2_X1 U15906 ( .A(n13103), .B(n12735), .ZN(n13313) );
  NAND2_X1 U15907 ( .A1(n13313), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13314) );
  INV_X1 U15908 ( .A(n13103), .ZN(n12736) );
  NAND2_X1 U15909 ( .A1(n12736), .A2(n12735), .ZN(n12737) );
  XNOR2_X1 U15910 ( .A(n12738), .B(n20120), .ZN(n13396) );
  NAND2_X1 U15911 ( .A1(n13395), .A2(n13396), .ZN(n13394) );
  NAND2_X1 U15912 ( .A1(n12738), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12739) );
  NAND2_X2 U15913 ( .A1(n13394), .A2(n12739), .ZN(n12747) );
  INV_X1 U15914 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20101) );
  OR2_X1 U15915 ( .A1(n20137), .A2(n12740), .ZN(n12746) );
  NAND2_X1 U15916 ( .A1(n12742), .A2(n12741), .ZN(n12758) );
  INV_X1 U15917 ( .A(n12755), .ZN(n12743) );
  XNOR2_X1 U15918 ( .A(n12758), .B(n12743), .ZN(n12744) );
  NAND2_X1 U15919 ( .A1(n12744), .A2(n13117), .ZN(n12745) );
  NAND2_X1 U15920 ( .A1(n12746), .A2(n12745), .ZN(n13410) );
  NAND2_X1 U15921 ( .A1(n12747), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12748) );
  INV_X1 U15923 ( .A(n12749), .ZN(n12753) );
  NAND2_X1 U15924 ( .A1(n12758), .A2(n12755), .ZN(n12750) );
  XNOR2_X1 U15925 ( .A(n12750), .B(n12756), .ZN(n12751) );
  AND2_X1 U15926 ( .A1(n12751), .A2(n13117), .ZN(n12752) );
  AOI21_X1 U15927 ( .B1(n12753), .B2(n12786), .A(n12752), .ZN(n20077) );
  NAND2_X1 U15928 ( .A1(n12754), .A2(n12786), .ZN(n12761) );
  AND2_X1 U15929 ( .A1(n12756), .A2(n12755), .ZN(n12757) );
  NAND2_X1 U15930 ( .A1(n12758), .A2(n12757), .ZN(n12767) );
  XNOR2_X1 U15931 ( .A(n12767), .B(n12768), .ZN(n12759) );
  NAND2_X1 U15932 ( .A1(n12759), .A2(n13117), .ZN(n12760) );
  NAND2_X1 U15933 ( .A1(n12761), .A2(n12760), .ZN(n12764) );
  XNOR2_X1 U15934 ( .A(n12764), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15846) );
  NAND2_X1 U15935 ( .A1(n12763), .A2(n12762), .ZN(n15843) );
  NAND2_X1 U15936 ( .A1(n12764), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12765) );
  NAND3_X1 U15937 ( .A1(n12789), .A2(n12766), .A3(n12786), .ZN(n12772) );
  INV_X1 U15938 ( .A(n12767), .ZN(n12769) );
  NAND2_X1 U15939 ( .A1(n12769), .A2(n12768), .ZN(n12777) );
  XNOR2_X1 U15940 ( .A(n12777), .B(n12778), .ZN(n12770) );
  NAND2_X1 U15941 ( .A1(n12770), .A2(n13117), .ZN(n12771) );
  INV_X1 U15942 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15837) );
  NAND2_X1 U15943 ( .A1(n15838), .A2(n15837), .ZN(n12773) );
  INV_X1 U15944 ( .A(n15838), .ZN(n12774) );
  NAND2_X1 U15945 ( .A1(n12774), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12775) );
  NAND2_X1 U15946 ( .A1(n12776), .A2(n12786), .ZN(n12783) );
  INV_X1 U15947 ( .A(n12777), .ZN(n12779) );
  NAND2_X1 U15948 ( .A1(n12779), .A2(n12778), .ZN(n12791) );
  XNOR2_X1 U15949 ( .A(n12791), .B(n12780), .ZN(n12781) );
  NAND2_X1 U15950 ( .A1(n12781), .A2(n13117), .ZN(n12782) );
  NAND2_X1 U15951 ( .A1(n12783), .A2(n12782), .ZN(n12784) );
  OR2_X1 U15952 ( .A1(n12784), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15833) );
  NAND2_X1 U15953 ( .A1(n12784), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15832) );
  AND2_X1 U15954 ( .A1(n12787), .A2(n12786), .ZN(n12788) );
  INV_X1 U15955 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13736) );
  NAND2_X1 U15956 ( .A1(n13737), .A2(n13736), .ZN(n12792) );
  INV_X1 U15957 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15943) );
  NAND2_X1 U15958 ( .A1(n9738), .A2(n15943), .ZN(n12794) );
  NAND2_X1 U15959 ( .A1(n9738), .A2(n15899), .ZN(n12795) );
  NAND2_X1 U15960 ( .A1(n14719), .A2(n12795), .ZN(n14737) );
  INV_X1 U15961 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14734) );
  NAND2_X1 U15962 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12796) );
  NAND2_X1 U15963 ( .A1(n9738), .A2(n12796), .ZN(n14728) );
  NAND2_X1 U15964 ( .A1(n14735), .A2(n14728), .ZN(n12797) );
  NOR2_X1 U15965 ( .A1(n14737), .A2(n12797), .ZN(n14721) );
  NAND2_X1 U15966 ( .A1(n9738), .A2(n14856), .ZN(n12798) );
  NAND2_X1 U15967 ( .A1(n14721), .A2(n12798), .ZN(n14707) );
  NAND2_X1 U15968 ( .A1(n15794), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12799) );
  NAND2_X1 U15969 ( .A1(n14719), .A2(n12799), .ZN(n15805) );
  INV_X1 U15970 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14855) );
  NAND2_X1 U15971 ( .A1(n9738), .A2(n14855), .ZN(n15802) );
  OAI21_X1 U15972 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n15794), .ZN(n12800) );
  INV_X1 U15973 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12801) );
  NAND2_X1 U15974 ( .A1(n9738), .A2(n12801), .ZN(n12802) );
  NOR2_X1 U15975 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14730) );
  NAND2_X1 U15976 ( .A1(n14730), .A2(n14734), .ZN(n12803) );
  NAND2_X1 U15977 ( .A1(n15794), .A2(n12803), .ZN(n14718) );
  NOR2_X1 U15978 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15638) );
  INV_X1 U15979 ( .A(n15638), .ZN(n15607) );
  XNOR2_X1 U15980 ( .A(n9738), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14701) );
  AND2_X1 U15981 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15629) );
  INV_X1 U15982 ( .A(n15629), .ZN(n12805) );
  INV_X1 U15983 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12804) );
  INV_X1 U15984 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14820) );
  NAND3_X1 U15985 ( .A1(n15864), .A2(n15851), .A3(n14820), .ZN(n14644) );
  AND2_X1 U15986 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14821) );
  AND2_X1 U15987 ( .A1(n14821), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14822) );
  INV_X1 U15988 ( .A(n14822), .ZN(n14643) );
  INV_X1 U15989 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14795) );
  NAND3_X1 U15990 ( .A1(n14630), .A2(n15794), .A3(n14795), .ZN(n12810) );
  AND2_X1 U15991 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14796) );
  INV_X1 U15992 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14783) );
  XNOR2_X1 U15993 ( .A(n12812), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14778) );
  NOR2_X1 U15994 ( .A1(n12813), .A2(n20160), .ZN(n12815) );
  NAND2_X1 U15995 ( .A1(n14879), .A2(n20144), .ZN(n12814) );
  AND2_X1 U15996 ( .A1(n12965), .A2(n12817), .ZN(n13131) );
  NAND2_X1 U15997 ( .A1(n12819), .A2(n12818), .ZN(n12823) );
  AOI22_X1 U15998 ( .A1(n12075), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12820), .ZN(n12821) );
  INV_X1 U15999 ( .A(n12821), .ZN(n12822) );
  XNOR2_X2 U16000 ( .A(n12823), .B(n12822), .ZN(n14357) );
  NOR2_X1 U16001 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20654) );
  NOR2_X1 U16002 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20707), .ZN(n15605) );
  AND2_X1 U16003 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n15605), .ZN(n12824) );
  NAND2_X1 U16004 ( .A1(n14357), .A2(n14666), .ZN(n12835) );
  NAND2_X1 U16005 ( .A1(n20644), .A2(n12831), .ZN(n20796) );
  NAND2_X1 U16006 ( .A1(n20796), .A2(n20708), .ZN(n12825) );
  NAND2_X1 U16007 ( .A1(n20708), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12827) );
  NAND2_X1 U16008 ( .A1(n21079), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12826) );
  AND2_X1 U16009 ( .A1(n12827), .A2(n12826), .ZN(n13101) );
  INV_X1 U16010 ( .A(n13101), .ZN(n12828) );
  INV_X1 U16011 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14362) );
  INV_X1 U16012 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20776) );
  NOR2_X1 U16013 ( .A1(n20107), .A2(n20776), .ZN(n14774) );
  AOI21_X1 U16014 ( .B1(n20076), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14774), .ZN(n12832) );
  OAI21_X1 U16015 ( .B1(n20085), .B2(n13616), .A(n12832), .ZN(n12833) );
  INV_X1 U16016 ( .A(n12833), .ZN(n12834) );
  OAI211_X1 U16017 ( .C1(n14778), .C2(n19900), .A(n12835), .B(n12834), .ZN(
        P1_U2968) );
  NOR2_X1 U16018 ( .A1(n14348), .A2(n19894), .ZN(n12836) );
  NAND2_X1 U16019 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n15977) );
  NAND2_X1 U16020 ( .A1(n20155), .A2(n15977), .ZN(n12849) );
  AND2_X1 U16021 ( .A1(n12965), .A2(n14350), .ZN(n13059) );
  NAND2_X1 U16022 ( .A1(n14351), .A2(n13059), .ZN(n12845) );
  INV_X1 U16023 ( .A(n12591), .ZN(n13362) );
  INV_X1 U16024 ( .A(n12837), .ZN(n12840) );
  NOR3_X1 U16025 ( .A1(n12840), .A2(n12839), .A3(n12838), .ZN(n12843) );
  OAI21_X1 U16026 ( .B1(n12843), .B2(n12842), .A(n12841), .ZN(n14338) );
  AND2_X1 U16027 ( .A1(n15977), .A2(n14338), .ZN(n13121) );
  NAND2_X1 U16028 ( .A1(n13362), .A2(n13121), .ZN(n12844) );
  NAND2_X1 U16029 ( .A1(n12845), .A2(n12844), .ZN(n12960) );
  NAND2_X1 U16030 ( .A1(n12960), .A2(n13129), .ZN(n12848) );
  NAND2_X1 U16031 ( .A1(n12846), .A2(n14350), .ZN(n12847) );
  AND2_X1 U16032 ( .A1(n20015), .A2(n14345), .ZN(n12850) );
  NAND2_X1 U16033 ( .A1(n14357), .A2(n12850), .ZN(n12869) );
  NOR4_X1 U16034 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12854) );
  NOR4_X1 U16035 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_15__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n12853) );
  NOR4_X1 U16036 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12852) );
  NOR4_X1 U16037 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12851) );
  AND4_X1 U16038 ( .A1(n12854), .A2(n12853), .A3(n12852), .A4(n12851), .ZN(
        n12859) );
  NOR4_X1 U16039 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_14__SCAN_IN), .ZN(n12857) );
  NOR4_X1 U16040 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12856) );
  NOR4_X1 U16041 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12855) );
  INV_X1 U16042 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20725) );
  AND4_X1 U16043 ( .A1(n12857), .A2(n12856), .A3(n12855), .A4(n20725), .ZN(
        n12858) );
  NAND2_X1 U16044 ( .A1(n12859), .A2(n12858), .ZN(n12860) );
  AND2_X2 U16045 ( .A1(n12860), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20143)
         );
  INV_X1 U16046 ( .A(n20143), .ZN(n12861) );
  NOR2_X1 U16047 ( .A1(n9740), .A2(n12861), .ZN(n12862) );
  NAND2_X1 U16048 ( .A1(n20015), .A2(n12862), .ZN(n14612) );
  INV_X1 U16049 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19239) );
  NOR2_X1 U16050 ( .A1(n14612), .A2(n19239), .ZN(n12867) );
  NOR3_X1 U16051 ( .A1(n15768), .A2(n20143), .A3(n9740), .ZN(n12864) );
  AOI22_X1 U16052 ( .A1(n14619), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15768), .ZN(n12865) );
  INV_X1 U16053 ( .A(n12865), .ZN(n12866) );
  NOR2_X1 U16054 ( .A1(n12867), .A2(n12866), .ZN(n12868) );
  NAND2_X1 U16055 ( .A1(n12869), .A2(n12868), .ZN(P1_U2873) );
  INV_X1 U16056 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19863) );
  NOR2_X1 U16057 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(n19863), .ZN(n12871) );
  NOR4_X1 U16058 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12870) );
  INV_X1 U16059 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20987) );
  NAND4_X1 U16060 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(n12871), .A3(n12870), .A4(
        n20987), .ZN(n12883) );
  NOR2_X1 U16061 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12883), .ZN(n16473)
         );
  INV_X1 U16062 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20913) );
  INV_X1 U16063 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20962) );
  AND4_X1 U16064 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(P1_W_R_N_REG_SCAN_IN), .A3(
        n20913), .A4(n20962), .ZN(n12873) );
  NOR4_X1 U16065 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_BE_N_REG_3__SCAN_IN), .A4(P1_D_C_N_REG_SCAN_IN), .ZN(n12872) );
  NAND3_X1 U16066 ( .A1(n20143), .A2(n12873), .A3(n12872), .ZN(U214) );
  NOR4_X1 U16067 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n12877) );
  NOR4_X1 U16068 ( .A1(P2_ADDRESS_REG_21__SCAN_IN), .A2(
        P2_ADDRESS_REG_20__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_18__SCAN_IN), .ZN(n12876) );
  NOR4_X1 U16069 ( .A1(P2_ADDRESS_REG_8__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n12875) );
  NOR4_X1 U16070 ( .A1(P2_ADDRESS_REG_12__SCAN_IN), .A2(
        P2_ADDRESS_REG_11__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_9__SCAN_IN), .ZN(n12874) );
  NAND4_X1 U16071 ( .A1(n12877), .A2(n12876), .A3(n12875), .A4(n12874), .ZN(
        n12882) );
  NOR2_X1 U16072 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .ZN(n21092) );
  NOR3_X1 U16073 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_2__SCAN_IN), .A3(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n12880) );
  NOR4_X1 U16074 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_23__SCAN_IN), .A4(
        P2_ADDRESS_REG_22__SCAN_IN), .ZN(n12879) );
  NOR4_X1 U16075 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12878) );
  NAND4_X1 U16076 ( .A1(n21092), .A2(n12880), .A3(n12879), .A4(n12878), .ZN(
        n12881) );
  NOR2_X1 U16077 ( .A1(n13811), .A2(n12883), .ZN(n16408) );
  NAND2_X1 U16078 ( .A1(n16408), .A2(U214), .ZN(U212) );
  AOI21_X1 U16079 ( .B1(n16128), .B2(n12895), .A(n14901), .ZN(n16115) );
  AOI21_X1 U16080 ( .B1(n16146), .B2(n12893), .A(n9834), .ZN(n16138) );
  AOI21_X1 U16081 ( .B1(n16170), .B2(n12891), .A(n12894), .ZN(n18974) );
  AOI21_X1 U16082 ( .B1(n21003), .B2(n12889), .A(n12892), .ZN(n18994) );
  AOI21_X1 U16083 ( .B1(n15248), .B2(n12887), .A(n12890), .ZN(n15249) );
  AOI21_X1 U16084 ( .B1(n16205), .B2(n12885), .A(n12888), .ZN(n19034) );
  AOI21_X1 U16085 ( .B1(n13661), .B2(n12884), .A(n12886), .ZN(n13659) );
  OAI22_X1 U16086 ( .A1(n19884), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19078) );
  INV_X1 U16087 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13695) );
  OAI22_X1 U16088 ( .A1(n19884), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n13695), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13702) );
  AND2_X1 U16089 ( .A1(n19078), .A2(n13702), .ZN(n13670) );
  OAI21_X1 U16090 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n12884), .ZN(n13672) );
  NAND2_X1 U16091 ( .A1(n13670), .A2(n13672), .ZN(n13657) );
  NOR2_X1 U16092 ( .A1(n13659), .A2(n13657), .ZN(n19051) );
  OAI21_X1 U16093 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n12886), .A(
        n12885), .ZN(n19166) );
  NAND2_X1 U16094 ( .A1(n19051), .A2(n19166), .ZN(n19031) );
  NOR2_X1 U16095 ( .A1(n19034), .A2(n19031), .ZN(n19018) );
  OAI21_X1 U16096 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n12888), .A(
        n12887), .ZN(n19019) );
  NAND2_X1 U16097 ( .A1(n19018), .A2(n19019), .ZN(n13683) );
  NOR2_X1 U16098 ( .A1(n15249), .A2(n13683), .ZN(n19004) );
  OAI21_X1 U16099 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n12890), .A(
        n12889), .ZN(n19005) );
  NAND2_X1 U16100 ( .A1(n19004), .A2(n19005), .ZN(n18993) );
  NOR2_X1 U16101 ( .A1(n18994), .A2(n18993), .ZN(n18986) );
  OAI21_X1 U16102 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n12892), .A(
        n12891), .ZN(n18987) );
  NAND2_X1 U16103 ( .A1(n18986), .A2(n18987), .ZN(n18972) );
  NOR2_X1 U16104 ( .A1(n18974), .A2(n18972), .ZN(n18961) );
  OAI21_X1 U16105 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n12894), .A(
        n12893), .ZN(n18962) );
  NAND2_X1 U16106 ( .A1(n18961), .A2(n18962), .ZN(n13708) );
  NOR2_X1 U16107 ( .A1(n16138), .A2(n13708), .ZN(n13709) );
  OAI21_X1 U16108 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n9834), .A(
        n12895), .ZN(n18947) );
  NAND2_X1 U16109 ( .A1(n13709), .A2(n18947), .ZN(n12897) );
  NOR2_X1 U16110 ( .A1(n16115), .A2(n12897), .ZN(n18934) );
  NOR3_X1 U16111 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15640) );
  NAND2_X1 U16112 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15640), .ZN(n19741) );
  NAND2_X1 U16113 ( .A1(n19036), .A2(n19032), .ZN(n19077) );
  AOI211_X1 U16114 ( .C1(n16115), .C2(n12897), .A(n18934), .B(n19077), .ZN(
        n12921) );
  INV_X1 U16115 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19783) );
  NAND2_X1 U16116 ( .A1(n12898), .A2(n19737), .ZN(n12900) );
  OR2_X1 U16117 ( .A1(n13033), .A2(n12900), .ZN(n19049) );
  NAND2_X1 U16118 ( .A1(n19872), .A2(n11189), .ZN(n15639) );
  NOR3_X1 U16119 ( .A1(n19884), .A2(n19871), .A3(n15639), .ZN(n16342) );
  OR2_X1 U16120 ( .A1(n19029), .A2(n16342), .ZN(n12901) );
  NOR2_X1 U16121 ( .A1(n19036), .A2(n12901), .ZN(n12902) );
  INV_X2 U16122 ( .A(n13294), .ZN(n19152) );
  NAND2_X1 U16123 ( .A1(n19882), .A2(n12927), .ZN(n16349) );
  AND2_X1 U16124 ( .A1(n19152), .A2(n16349), .ZN(n15988) );
  INV_X1 U16125 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n12903) );
  NAND2_X1 U16126 ( .A1(n19882), .A2(n19880), .ZN(n12915) );
  NAND2_X1 U16127 ( .A1(n12903), .A2(n12915), .ZN(n12904) );
  NOR2_X1 U16128 ( .A1(n13156), .A2(n12904), .ZN(n12905) );
  OR2_X2 U16129 ( .A1(n15988), .A2(n12905), .ZN(n19065) );
  AOI22_X1 U16130 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19043), .B1(
        P2_EBX_REG_15__SCAN_IN), .B2(n19065), .ZN(n12906) );
  OAI211_X1 U16131 ( .C1(n19783), .C2(n19061), .A(n12906), .B(n19045), .ZN(
        n12920) );
  NOR2_X1 U16132 ( .A1(n19875), .A2(n12907), .ZN(n12917) );
  AND2_X1 U16133 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n12915), .ZN(n12908) );
  NAND2_X1 U16134 ( .A1(n12917), .A2(n12908), .ZN(n19067) );
  NAND2_X1 U16135 ( .A1(n19052), .A2(n19036), .ZN(n19071) );
  INV_X1 U16136 ( .A(n16115), .ZN(n12909) );
  OAI22_X1 U16137 ( .A1(n12910), .A2(n19067), .B1(n19071), .B2(n12909), .ZN(
        n12919) );
  OAI21_X1 U16138 ( .B1(n16246), .B2(n12911), .A(n14016), .ZN(n16236) );
  INV_X1 U16139 ( .A(n16349), .ZN(n12912) );
  NOR2_X1 U16140 ( .A1(n12913), .A2(n13638), .ZN(n12914) );
  NOR2_X1 U16141 ( .A1(n13764), .A2(n12914), .ZN(n16241) );
  INV_X1 U16142 ( .A(n16241), .ZN(n13732) );
  INV_X1 U16143 ( .A(n12915), .ZN(n12916) );
  NAND2_X1 U16144 ( .A1(n12917), .A2(n12916), .ZN(n19047) );
  OAI22_X1 U16145 ( .A1(n16236), .A2(n19063), .B1(n13732), .B2(n19047), .ZN(
        n12918) );
  OR4_X1 U16146 ( .A1(n12921), .A2(n12920), .A3(n12919), .A4(n12918), .ZN(
        P2_U2840) );
  INV_X1 U16147 ( .A(n19049), .ZN(n19074) );
  INV_X1 U16148 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12923) );
  INV_X1 U16149 ( .A(n18878), .ZN(n12922) );
  OAI211_X1 U16150 ( .C1(n19074), .C2(n12923), .A(n12922), .B(n13156), .ZN(
        P2_U2814) );
  INV_X1 U16151 ( .A(n11376), .ZN(n12925) );
  OAI21_X1 U16152 ( .B1(n18878), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19875), 
        .ZN(n12924) );
  OAI21_X1 U16153 ( .B1(n12925), .B2(n19875), .A(n12924), .ZN(P2_U3612) );
  NOR2_X1 U16154 ( .A1(n12925), .A2(n19876), .ZN(n12926) );
  NOR4_X1 U16155 ( .A1(n10692), .A2(n12927), .A3(n12926), .A4(n16313), .ZN(
        n16323) );
  INV_X1 U16156 ( .A(n19737), .ZN(n16357) );
  NOR2_X1 U16157 ( .A1(n16323), .A2(n16357), .ZN(n19869) );
  OAI21_X1 U16158 ( .B1(n12929), .B2(n19869), .A(n12928), .ZN(P2_U2819) );
  INV_X1 U16159 ( .A(n12930), .ZN(n14340) );
  AND2_X1 U16160 ( .A1(n14338), .A2(n14340), .ZN(n14349) );
  NAND2_X1 U16161 ( .A1(n14349), .A2(n13129), .ZN(n12932) );
  AND2_X1 U16162 ( .A1(n20654), .A2(n20707), .ZN(n13627) );
  AOI21_X1 U16163 ( .B1(n12932), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13627), 
        .ZN(n12931) );
  NAND2_X1 U16164 ( .A1(n12956), .A2(n12931), .ZN(P1_U2801) );
  NOR2_X1 U16165 ( .A1(n14350), .A2(n12609), .ZN(n12934) );
  OAI21_X1 U16166 ( .B1(n13627), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n20798), 
        .ZN(n12933) );
  OAI21_X1 U16167 ( .B1(n20798), .B2(n12934), .A(n12933), .ZN(P1_U3487) );
  NOR2_X1 U16168 ( .A1(n13033), .A2(n16357), .ZN(n12935) );
  NAND2_X1 U16169 ( .A1(n13025), .A2(n12935), .ZN(n12936) );
  NAND2_X1 U16170 ( .A1(n19148), .A2(n12937), .ZN(n19115) );
  INV_X1 U16171 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15085) );
  NAND2_X1 U16172 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n13540) );
  NOR2_X1 U16173 ( .A1(n13540), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19147) );
  INV_X1 U16174 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n12938) );
  INV_X1 U16175 ( .A(n19877), .ZN(n19144) );
  INV_X1 U16176 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n21025) );
  OAI222_X1 U16177 ( .A1(n19115), .A2(n15085), .B1(n19877), .B2(n12938), .C1(
        n19150), .C2(n21025), .ZN(P2_U2926) );
  INV_X1 U16178 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n16480) );
  INV_X1 U16179 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13238) );
  INV_X1 U16180 ( .A(P2_UWORD_REG_14__SCAN_IN), .ZN(n20814) );
  OAI222_X1 U16181 ( .A1(n19150), .A2(n16480), .B1(n19115), .B2(n13238), .C1(
        n20814), .C2(n19877), .ZN(P2_U2921) );
  INV_X1 U16182 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U16183 ( .A1(n19144), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12939) );
  OAI21_X1 U16184 ( .B1(n12940), .B2(n19115), .A(n12939), .ZN(P2_U2934) );
  INV_X1 U16185 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U16186 ( .A1(n19147), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12941) );
  OAI21_X1 U16187 ( .B1(n12942), .B2(n19115), .A(n12941), .ZN(P2_U2928) );
  INV_X1 U16188 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15068) );
  AOI22_X1 U16189 ( .A1(n19144), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12943) );
  OAI21_X1 U16190 ( .B1(n15068), .B2(n19115), .A(n12943), .ZN(P2_U2924) );
  INV_X1 U16191 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15049) );
  AOI22_X1 U16192 ( .A1(n19144), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12944) );
  OAI21_X1 U16193 ( .B1(n15049), .B2(n19115), .A(n12944), .ZN(P2_U2922) );
  INV_X1 U16194 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n20848) );
  AOI22_X1 U16195 ( .A1(n19147), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12945) );
  OAI21_X1 U16196 ( .B1(n20848), .B2(n19115), .A(n12945), .ZN(P2_U2931) );
  AOI22_X1 U16197 ( .A1(n19147), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12946) );
  OAI21_X1 U16198 ( .B1(n12947), .B2(n19115), .A(n12946), .ZN(P2_U2930) );
  INV_X1 U16199 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U16200 ( .A1(n19147), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12948) );
  OAI21_X1 U16201 ( .B1(n15058), .B2(n19115), .A(n12948), .ZN(P2_U2923) );
  INV_X1 U16202 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n12950) );
  AOI22_X1 U16203 ( .A1(n19147), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12949) );
  OAI21_X1 U16204 ( .B1(n12950), .B2(n19115), .A(n12949), .ZN(P2_U2932) );
  INV_X1 U16205 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12952) );
  AOI22_X1 U16206 ( .A1(n19144), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12951) );
  OAI21_X1 U16207 ( .B1(n12952), .B2(n19115), .A(n12951), .ZN(P2_U2933) );
  INV_X1 U16208 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13295) );
  AOI22_X1 U16209 ( .A1(n19147), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12953) );
  OAI21_X1 U16210 ( .B1(n13295), .B2(n19115), .A(n12953), .ZN(P2_U2925) );
  INV_X1 U16211 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13291) );
  AOI22_X1 U16212 ( .A1(n19147), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12954) );
  OAI21_X1 U16213 ( .B1(n13291), .B2(n19115), .A(n12954), .ZN(P2_U2927) );
  INV_X1 U16214 ( .A(n15977), .ZN(n20799) );
  AND2_X1 U16215 ( .A1(n20803), .A2(n20799), .ZN(n12955) );
  NAND2_X1 U16216 ( .A1(n13212), .A2(n12606), .ZN(n13174) );
  INV_X1 U16217 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n20022) );
  NAND2_X1 U16218 ( .A1(n13212), .A2(n20155), .ZN(n13051) );
  INV_X1 U16219 ( .A(DATAI_15_), .ZN(n12958) );
  INV_X1 U16220 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12957) );
  MUX2_X1 U16221 ( .A(n12958), .B(n12957), .S(n20143), .Z(n13901) );
  INV_X1 U16222 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20023) );
  OAI222_X1 U16223 ( .A1(n13174), .A2(n20022), .B1(n13051), .B2(n13901), .C1(
        n13212), .C2(n20023), .ZN(P1_U2967) );
  INV_X1 U16224 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20532) );
  INV_X1 U16225 ( .A(n12959), .ZN(n12971) );
  INV_X1 U16226 ( .A(n12960), .ZN(n12970) );
  NOR2_X1 U16227 ( .A1(n12930), .A2(n12606), .ZN(n14031) );
  INV_X1 U16228 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12961) );
  NAND2_X1 U16229 ( .A1(n10231), .A2(n12961), .ZN(n15624) );
  INV_X1 U16230 ( .A(n15624), .ZN(n12976) );
  NAND2_X1 U16231 ( .A1(n14031), .A2(n12976), .ZN(n12978) );
  AND2_X1 U16232 ( .A1(n12610), .A2(n15624), .ZN(n12963) );
  NAND2_X1 U16233 ( .A1(n12962), .A2(n20188), .ZN(n13135) );
  OR2_X1 U16234 ( .A1(n12963), .A2(n13135), .ZN(n12964) );
  AOI21_X1 U16235 ( .B1(n12978), .B2(n12964), .A(n20799), .ZN(n12968) );
  AOI21_X1 U16236 ( .B1(n12965), .B2(n13143), .A(n14340), .ZN(n13125) );
  NOR2_X1 U16237 ( .A1(n14474), .A2(n20160), .ZN(n12966) );
  OR2_X1 U16238 ( .A1(n13125), .A2(n12966), .ZN(n12967) );
  AOI21_X1 U16239 ( .B1(n14351), .B2(n12968), .A(n12967), .ZN(n12969) );
  NAND3_X1 U16240 ( .A1(n12971), .A2(n12970), .A3(n12969), .ZN(n15584) );
  NAND2_X1 U16241 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15981) );
  NOR2_X1 U16242 ( .A1(n20708), .A2(n15981), .ZN(n13368) );
  AOI22_X1 U16243 ( .A1(n15584), .A2(n13129), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n13368), .ZN(n12974) );
  OAI21_X1 U16244 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20532), .A(n12974), 
        .ZN(n14894) );
  INV_X1 U16245 ( .A(n20288), .ZN(n20519) );
  XNOR2_X1 U16246 ( .A(n12972), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19963) );
  NAND3_X1 U16247 ( .A1(n19963), .A2(n14032), .A3(n13362), .ZN(n12973) );
  OAI22_X1 U16248 ( .A1(n14894), .A2(n12975), .B1(n12974), .B2(n12973), .ZN(
        P1_U3468) );
  INV_X1 U16249 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12983) );
  NAND2_X1 U16250 ( .A1(n13117), .A2(n12976), .ZN(n12977) );
  NOR2_X1 U16251 ( .A1(n13135), .A2(n12977), .ZN(n15570) );
  INV_X1 U16252 ( .A(n15570), .ZN(n12979) );
  AOI21_X1 U16253 ( .B1(n12979), .B2(n12978), .A(n19894), .ZN(n12980) );
  INV_X1 U16254 ( .A(n20051), .ZN(n12981) );
  NAND2_X1 U16255 ( .A1(n12981), .A2(n12593), .ZN(n20018) );
  OR2_X1 U16256 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15981), .ZN(n20800) );
  AOI22_X1 U16257 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12982) );
  OAI21_X1 U16258 ( .B1(n12983), .B2(n20018), .A(n12982), .ZN(P1_U2911) );
  INV_X1 U16259 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U16260 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12984) );
  OAI21_X1 U16261 ( .B1(n12985), .B2(n20018), .A(n12984), .ZN(P1_U2920) );
  AOI22_X1 U16262 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12986) );
  OAI21_X1 U16263 ( .B1(n14593), .B2(n20018), .A(n12986), .ZN(P1_U2913) );
  INV_X1 U16264 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U16265 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12987) );
  OAI21_X1 U16266 ( .B1(n12988), .B2(n20018), .A(n12987), .ZN(P1_U2914) );
  INV_X1 U16267 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12990) );
  AOI22_X1 U16268 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12989) );
  OAI21_X1 U16269 ( .B1(n12990), .B2(n20018), .A(n12989), .ZN(P1_U2906) );
  INV_X1 U16270 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n21018) );
  AOI22_X1 U16271 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12991) );
  OAI21_X1 U16272 ( .B1(n21018), .B2(n20018), .A(n12991), .ZN(P1_U2907) );
  INV_X1 U16273 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U16274 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12992) );
  OAI21_X1 U16275 ( .B1(n12993), .B2(n20018), .A(n12992), .ZN(P1_U2908) );
  INV_X1 U16276 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12995) );
  AOI22_X1 U16277 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12994) );
  OAI21_X1 U16278 ( .B1(n12995), .B2(n20018), .A(n12994), .ZN(P1_U2909) );
  AOI22_X1 U16279 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12996) );
  OAI21_X1 U16280 ( .B1(n14610), .B2(n20018), .A(n12996), .ZN(P1_U2919) );
  INV_X1 U16281 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U16282 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12997) );
  OAI21_X1 U16283 ( .B1(n12998), .B2(n20018), .A(n12997), .ZN(P1_U2916) );
  INV_X1 U16284 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13000) );
  AOI22_X1 U16285 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12999) );
  OAI21_X1 U16286 ( .B1(n13000), .B2(n20018), .A(n12999), .ZN(P1_U2915) );
  INV_X1 U16287 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U16288 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13001) );
  OAI21_X1 U16289 ( .B1(n13002), .B2(n20018), .A(n13001), .ZN(P1_U2918) );
  INV_X1 U16290 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13004) );
  AOI22_X1 U16291 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13003) );
  OAI21_X1 U16292 ( .B1(n13004), .B2(n20018), .A(n13003), .ZN(P1_U2917) );
  MUX2_X1 U16293 ( .A(n16198), .B(n19169), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13011) );
  OAI21_X1 U16294 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13006), .A(
        n13005), .ZN(n13087) );
  OAI21_X1 U16295 ( .B1(n13693), .B2(n10225), .A(n13007), .ZN(n13008) );
  XNOR2_X1 U16296 ( .A(n13008), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13090) );
  NAND2_X1 U16297 ( .A1(n13090), .A2(n19175), .ZN(n13009) );
  NAND2_X1 U16298 ( .A1(n19029), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13080) );
  OAI211_X1 U16299 ( .C1(n13087), .C2(n19177), .A(n13009), .B(n13080), .ZN(
        n13010) );
  AOI211_X1 U16300 ( .C1(n19171), .C2(n13078), .A(n13011), .B(n13010), .ZN(
        n13012) );
  INV_X1 U16301 ( .A(n13012), .ZN(P2_U3013) );
  NAND2_X1 U16302 ( .A1(n10657), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U16303 ( .A1(n13301), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19825), .B2(n19861), .ZN(n13014) );
  AOI21_X1 U16304 ( .B1(n10757), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13016) );
  AND2_X1 U16305 ( .A1(n13017), .A2(n13016), .ZN(n13018) );
  INV_X1 U16306 ( .A(n16315), .ZN(n16317) );
  NAND2_X1 U16307 ( .A1(n16317), .A2(n16314), .ZN(n13029) );
  NAND2_X1 U16308 ( .A1(n13029), .A2(n9827), .ZN(n13019) );
  MUX2_X1 U16309 ( .A(n13021), .B(n13020), .S(n15040), .Z(n13022) );
  OAI21_X1 U16310 ( .B1(n19857), .B2(n15026), .A(n13022), .ZN(P2_U2887) );
  NOR2_X1 U16311 ( .A1(n19884), .A2(n13540), .ZN(n16359) );
  NOR2_X1 U16312 ( .A1(n13033), .A2(n13023), .ZN(n13024) );
  NAND2_X1 U16313 ( .A1(n13025), .A2(n13024), .ZN(n13031) );
  AND3_X1 U16314 ( .A1(n11647), .A2(n13026), .A3(n11376), .ZN(n13027) );
  AOI21_X1 U16315 ( .B1(n16315), .B2(n16316), .A(n13027), .ZN(n13038) );
  INV_X1 U16316 ( .A(n13028), .ZN(n13030) );
  AND4_X1 U16317 ( .A1(n13031), .A2(n13038), .A3(n13030), .A4(n13029), .ZN(
        n16331) );
  OAI22_X1 U16318 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19871), .B1(n16331), 
        .B2(n16357), .ZN(n13032) );
  AOI21_X1 U16319 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16359), .A(n13032), .ZN(
        n15526) );
  INV_X1 U16320 ( .A(n15526), .ZN(n13035) );
  NOR2_X1 U16321 ( .A1(n13033), .A2(n10757), .ZN(n16322) );
  NAND4_X1 U16322 ( .A1(n13035), .A2(n16322), .A3(n16321), .A4(n19827), .ZN(
        n13034) );
  OAI21_X1 U16323 ( .B1(n13036), .B2(n13035), .A(n13034), .ZN(P2_U3595) );
  NAND2_X1 U16324 ( .A1(n13038), .A2(n13037), .ZN(n13039) );
  INV_X1 U16325 ( .A(n19107), .ZN(n16079) );
  NAND2_X1 U16326 ( .A1(n19103), .A2(n19241), .ZN(n16092) );
  AOI21_X1 U16327 ( .B1(n19857), .B2(n16079), .A(n19087), .ZN(n13050) );
  INV_X1 U16328 ( .A(n13040), .ZN(n13046) );
  INV_X1 U16329 ( .A(n13041), .ZN(n13044) );
  INV_X1 U16330 ( .A(n13042), .ZN(n13043) );
  NAND2_X1 U16331 ( .A1(n13044), .A2(n13043), .ZN(n13045) );
  NAND2_X1 U16332 ( .A1(n13046), .A2(n13045), .ZN(n19062) );
  NOR2_X1 U16333 ( .A1(n10699), .A2(n19241), .ZN(n13047) );
  NAND2_X1 U16334 ( .A1(n19103), .A2(n13047), .ZN(n13593) );
  INV_X1 U16335 ( .A(n13593), .ZN(n19106) );
  OAI22_X1 U16336 ( .A1(n13811), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13812), .ZN(n13585) );
  INV_X1 U16337 ( .A(n13585), .ZN(n19081) );
  AOI22_X1 U16338 ( .A1(n19106), .A2(n19081), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19104), .ZN(n13049) );
  NAND3_X1 U16339 ( .A1(n19248), .A2(n16079), .A3(n19062), .ZN(n13048) );
  OAI211_X1 U16340 ( .C1(n13050), .C2(n19062), .A(n13049), .B(n13048), .ZN(
        P2_U2919) );
  INV_X1 U16341 ( .A(DATAI_13_), .ZN(n13053) );
  NAND2_X1 U16342 ( .A1(n20143), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13052) );
  OAI21_X1 U16343 ( .B1(n20143), .B2(n13053), .A(n13052), .ZN(n14567) );
  NAND2_X1 U16344 ( .A1(n20060), .A2(n14567), .ZN(n20070) );
  INV_X2 U16345 ( .A(n13212), .ZN(n20072) );
  NAND2_X1 U16346 ( .A1(n20072), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13054) );
  OAI211_X1 U16347 ( .C1(n13174), .C2(n21018), .A(n20070), .B(n13054), .ZN(
        P1_U2950) );
  INV_X1 U16348 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20036) );
  NAND2_X1 U16349 ( .A1(n20072), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13057) );
  INV_X1 U16350 ( .A(DATAI_8_), .ZN(n13056) );
  NAND2_X1 U16351 ( .A1(n20143), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13055) );
  OAI21_X1 U16352 ( .B1(n20143), .B2(n13056), .A(n13055), .ZN(n14589) );
  NAND2_X1 U16353 ( .A1(n20060), .A2(n14589), .ZN(n13211) );
  OAI211_X1 U16354 ( .C1(n13174), .C2(n20036), .A(n13057), .B(n13211), .ZN(
        P1_U2960) );
  INV_X1 U16355 ( .A(n14894), .ZN(n13070) );
  INV_X1 U16356 ( .A(n20520), .ZN(n20140) );
  INV_X1 U16357 ( .A(n13059), .ZN(n14337) );
  NAND2_X1 U16358 ( .A1(n14343), .A2(n14337), .ZN(n13349) );
  XNOR2_X1 U16359 ( .A(n14884), .B(n9746), .ZN(n13065) );
  NAND2_X1 U16360 ( .A1(n13349), .A2(n13065), .ZN(n13063) );
  XNOR2_X1 U16361 ( .A(n11952), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13061) );
  NOR2_X1 U16362 ( .A1(n14879), .A2(n13065), .ZN(n13060) );
  AOI22_X1 U16363 ( .A1(n14031), .A2(n13061), .B1(n13353), .B2(n13060), .ZN(
        n13062) );
  NAND2_X1 U16364 ( .A1(n13063), .A2(n13062), .ZN(n13064) );
  AOI21_X1 U16365 ( .B1(n20140), .B2(n14882), .A(n13064), .ZN(n15579) );
  INV_X1 U16366 ( .A(n15579), .ZN(n13067) );
  INV_X1 U16367 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20110) );
  NOR2_X1 U16368 ( .A1(n20707), .A2(n20110), .ZN(n14886) );
  INV_X1 U16369 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20879) );
  AOI22_X1 U16370 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n20135), .B2(n20879), .ZN(
        n14883) );
  INV_X1 U16371 ( .A(n13065), .ZN(n13066) );
  AOI222_X1 U16372 ( .A1(n13067), .A2(n14032), .B1(n14886), .B2(n14883), .C1(
        n13066), .C2(n15602), .ZN(n13069) );
  NAND2_X1 U16373 ( .A1(n13070), .A2(n9746), .ZN(n13068) );
  OAI21_X1 U16374 ( .B1(n13070), .B2(n13069), .A(n13068), .ZN(P1_U3472) );
  NAND2_X1 U16375 ( .A1(n13301), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13073) );
  NAND2_X1 U16376 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19558) );
  NAND2_X1 U16377 ( .A1(n10893), .A2(n19861), .ZN(n19464) );
  AND2_X1 U16378 ( .A1(n19558), .A2(n19464), .ZN(n19402) );
  NAND2_X1 U16379 ( .A1(n19402), .A2(n19825), .ZN(n19530) );
  NAND2_X1 U16380 ( .A1(n13073), .A2(n19530), .ZN(n13074) );
  INV_X1 U16381 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13694) );
  INV_X1 U16382 ( .A(n13078), .ZN(n15508) );
  MUX2_X1 U16383 ( .A(n13694), .B(n15508), .S(n14992), .Z(n13079) );
  OAI21_X1 U16384 ( .B1(n19281), .B2(n15026), .A(n13079), .ZN(P2_U2886) );
  OAI21_X1 U16385 ( .B1(n13986), .B2(n15510), .A(n13080), .ZN(n13089) );
  INV_X1 U16386 ( .A(n16309), .ZN(n15365) );
  OAI211_X1 U16387 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15365), .B(n13081), .ZN(n13086) );
  OAI21_X1 U16388 ( .B1(n13084), .B2(n13083), .A(n13082), .ZN(n19852) );
  NAND2_X1 U16389 ( .A1(n19186), .A2(n19852), .ZN(n13085) );
  OAI211_X1 U16390 ( .C1(n13087), .C2(n19196), .A(n13086), .B(n13085), .ZN(
        n13088) );
  AOI211_X1 U16391 ( .C1(n19187), .C2(n13090), .A(n13089), .B(n13088), .ZN(
        n13091) );
  OAI21_X1 U16392 ( .B1(n15508), .B2(n16266), .A(n13091), .ZN(P2_U3045) );
  INV_X1 U16393 ( .A(n13092), .ZN(n13095) );
  OAI21_X1 U16394 ( .B1(n13095), .B2(n13094), .A(n13093), .ZN(n20017) );
  NAND2_X1 U16395 ( .A1(n13096), .A2(n20110), .ZN(n13098) );
  AND2_X1 U16396 ( .A1(n13098), .A2(n13097), .ZN(n19990) );
  INV_X1 U16397 ( .A(n19990), .ZN(n13099) );
  OAI222_X1 U16398 ( .A1(n20017), .A2(n14561), .B1(n20012), .B2(n13100), .C1(
        n13099), .C2(n20001), .ZN(P1_U2872) );
  NAND2_X1 U16399 ( .A1(n13101), .A2(n15784), .ZN(n13106) );
  INV_X1 U16400 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13102) );
  NOR2_X1 U16401 ( .A1(n20107), .A2(n13102), .ZN(n13148) );
  OAI21_X1 U16402 ( .B1(n13104), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13103), .ZN(n13155) );
  NOR2_X1 U16403 ( .A1(n19900), .A2(n13155), .ZN(n13105) );
  AOI211_X1 U16404 ( .C1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13106), .A(
        n13148), .B(n13105), .ZN(n13107) );
  OAI21_X1 U16405 ( .B1(n20142), .B2(n20017), .A(n13107), .ZN(P1_U2999) );
  OAI22_X1 U16406 ( .A1(n13811), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13812), .ZN(n19231) );
  XNOR2_X1 U16407 ( .A(n13109), .B(n13108), .ZN(n19025) );
  INV_X1 U16408 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19135) );
  OAI222_X1 U16409 ( .A1(n13593), .A2(n19231), .B1(n19025), .B2(n19113), .C1(
        n19135), .C2(n19103), .ZN(P2_U2913) );
  OAI21_X1 U16410 ( .B1(n13111), .B2(n13110), .A(n13336), .ZN(n14484) );
  INV_X1 U16411 ( .A(n13113), .ZN(n13112) );
  AND2_X1 U16412 ( .A1(n20015), .A2(n13113), .ZN(n15770) );
  INV_X1 U16413 ( .A(DATAI_1_), .ZN(n13115) );
  NAND2_X1 U16414 ( .A1(n20143), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13114) );
  OAI21_X1 U16415 ( .B1(n20143), .B2(n13115), .A(n13114), .ZN(n20154) );
  INV_X1 U16416 ( .A(n20154), .ZN(n13116) );
  INV_X1 U16417 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20048) );
  OAI222_X1 U16418 ( .A1(n14484), .A2(n20016), .B1(n20014), .B2(n13116), .C1(
        n20015), .C2(n20048), .ZN(P1_U2903) );
  OR2_X1 U16419 ( .A1(n13135), .A2(n20799), .ZN(n13118) );
  AOI22_X1 U16420 ( .A1(n13118), .A2(n12593), .B1(n13117), .B2(n15624), .ZN(
        n13119) );
  OAI21_X1 U16421 ( .B1(n13120), .B2(n13119), .A(n14351), .ZN(n13124) );
  NAND2_X1 U16422 ( .A1(n20155), .A2(n15624), .ZN(n13122) );
  NAND2_X1 U16423 ( .A1(n13122), .A2(n13121), .ZN(n13123) );
  MUX2_X1 U16424 ( .A(n13124), .B(n13123), .S(n20160), .Z(n13128) );
  NOR2_X1 U16425 ( .A1(n14879), .A2(n12606), .ZN(n13126) );
  AOI21_X1 U16426 ( .B1(n14342), .B2(n13126), .A(n13125), .ZN(n13127) );
  NAND2_X1 U16427 ( .A1(n13128), .A2(n13127), .ZN(n13130) );
  INV_X1 U16428 ( .A(n13131), .ZN(n14336) );
  INV_X1 U16429 ( .A(n13137), .ZN(n13132) );
  NAND2_X1 U16430 ( .A1(n13132), .A2(n13136), .ZN(n13133) );
  AND4_X1 U16431 ( .A1(n14337), .A2(n14336), .A3(n9779), .A4(n13133), .ZN(
        n13134) );
  NOR2_X2 U16432 ( .A1(n13150), .A2(n13134), .ZN(n20128) );
  OAI22_X1 U16433 ( .A1(n13137), .A2(n13136), .B1(n20803), .B2(n13135), .ZN(
        n13138) );
  INV_X1 U16434 ( .A(n13139), .ZN(n13140) );
  NAND4_X1 U16435 ( .A1(n13143), .A2(n13142), .A3(n13141), .A4(n13140), .ZN(
        n13144) );
  OR2_X1 U16436 ( .A1(n13145), .A2(n13144), .ZN(n13146) );
  NAND2_X1 U16437 ( .A1(n13149), .A2(n13146), .ZN(n15626) );
  NAND2_X1 U16438 ( .A1(n15626), .A2(n20114), .ZN(n14760) );
  NAND2_X1 U16439 ( .A1(n20110), .A2(n14760), .ZN(n20133) );
  INV_X1 U16440 ( .A(n20133), .ZN(n13147) );
  AOI211_X1 U16441 ( .C1(n20126), .C2(n19990), .A(n13148), .B(n13147), .ZN(
        n13154) );
  INV_X1 U16442 ( .A(n15893), .ZN(n13152) );
  NAND2_X1 U16443 ( .A1(n13150), .A2(n20107), .ZN(n20134) );
  INV_X1 U16444 ( .A(n20134), .ZN(n13151) );
  OAI21_X1 U16445 ( .B1(n13152), .B2(n13151), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13153) );
  OAI211_X1 U16446 ( .C1(n15913), .C2(n13155), .A(n13154), .B(n13153), .ZN(
        P1_U3031) );
  NOR3_X4 U16447 ( .A1(n13156), .A2(n14257), .A3(n19876), .ZN(n13287) );
  INV_X1 U16448 ( .A(n13287), .ZN(n13159) );
  AOI22_X1 U16449 ( .A1(n13812), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13550), .ZN(n13592) );
  INV_X1 U16450 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19120) );
  INV_X1 U16451 ( .A(n13156), .ZN(n13158) );
  NAND2_X1 U16452 ( .A1(n10757), .A2(n19876), .ZN(n13157) );
  NAND2_X2 U16453 ( .A1(n13158), .A2(n13157), .ZN(n19151) );
  INV_X1 U16454 ( .A(n19151), .ZN(n13286) );
  INV_X1 U16455 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n19119) );
  OAI222_X1 U16456 ( .A1(n13159), .A2(n13592), .B1(n13294), .B2(n19120), .C1(
        n13286), .C2(n19119), .ZN(P2_U2982) );
  AOI22_X1 U16457 ( .A1(n13812), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13550), .ZN(n19243) );
  XNOR2_X1 U16458 ( .A(n13161), .B(n13160), .ZN(n15477) );
  INV_X1 U16459 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19133) );
  OAI222_X1 U16460 ( .A1(n13593), .A2(n19243), .B1(n15477), .B2(n19113), .C1(
        n19133), .C2(n19103), .ZN(P2_U2912) );
  OR2_X1 U16461 ( .A1(n13163), .A2(n13162), .ZN(n13164) );
  NAND2_X1 U16462 ( .A1(n13165), .A2(n13164), .ZN(n20125) );
  INV_X1 U16463 ( .A(n20125), .ZN(n14485) );
  OAI22_X1 U16464 ( .A1(n20001), .A2(n14485), .B1(n14483), .B2(n20012), .ZN(
        n13166) );
  INV_X1 U16465 ( .A(n13166), .ZN(n13167) );
  OAI21_X1 U16466 ( .B1(n14561), .B2(n14484), .A(n13167), .ZN(P1_U2871) );
  AOI22_X1 U16467 ( .A1(n20073), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20072), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13170) );
  INV_X1 U16468 ( .A(DATAI_2_), .ZN(n13169) );
  NAND2_X1 U16469 ( .A1(n20143), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13168) );
  OAI21_X1 U16470 ( .B1(n20143), .B2(n13169), .A(n13168), .ZN(n20159) );
  NAND2_X1 U16471 ( .A1(n20060), .A2(n20159), .ZN(n13178) );
  NAND2_X1 U16472 ( .A1(n13170), .A2(n13178), .ZN(P1_U2954) );
  AOI22_X1 U16473 ( .A1(n20073), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20072), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13173) );
  INV_X1 U16474 ( .A(DATAI_5_), .ZN(n13172) );
  NAND2_X1 U16475 ( .A1(n20143), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13171) );
  OAI21_X1 U16476 ( .B1(n20143), .B2(n13172), .A(n13171), .ZN(n20175) );
  NAND2_X1 U16477 ( .A1(n20060), .A2(n20175), .ZN(n13197) );
  NAND2_X1 U16478 ( .A1(n13173), .A2(n13197), .ZN(P1_U2942) );
  INV_X2 U16479 ( .A(n13174), .ZN(n20073) );
  AOI22_X1 U16480 ( .A1(n20073), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20072), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13177) );
  INV_X1 U16481 ( .A(DATAI_3_), .ZN(n13176) );
  NAND2_X1 U16482 ( .A1(n20143), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13175) );
  OAI21_X1 U16483 ( .B1(n20143), .B2(n13176), .A(n13175), .ZN(n20164) );
  NAND2_X1 U16484 ( .A1(n20060), .A2(n20164), .ZN(n13189) );
  NAND2_X1 U16485 ( .A1(n13177), .A2(n13189), .ZN(P1_U2940) );
  AOI22_X1 U16486 ( .A1(n20073), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20072), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13179) );
  NAND2_X1 U16487 ( .A1(n13179), .A2(n13178), .ZN(P1_U2939) );
  AOI22_X1 U16488 ( .A1(n20073), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20072), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13182) );
  INV_X1 U16489 ( .A(DATAI_7_), .ZN(n13181) );
  NAND2_X1 U16490 ( .A1(n20143), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13180) );
  OAI21_X1 U16491 ( .B1(n20143), .B2(n13181), .A(n13180), .ZN(n20186) );
  NAND2_X1 U16492 ( .A1(n20060), .A2(n20186), .ZN(n13193) );
  NAND2_X1 U16493 ( .A1(n13182), .A2(n13193), .ZN(P1_U2944) );
  AOI22_X1 U16494 ( .A1(n20073), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20072), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13185) );
  INV_X1 U16495 ( .A(DATAI_6_), .ZN(n13184) );
  NAND2_X1 U16496 ( .A1(n20143), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13183) );
  OAI21_X1 U16497 ( .B1(n20143), .B2(n13184), .A(n13183), .ZN(n20180) );
  NAND2_X1 U16498 ( .A1(n20060), .A2(n20180), .ZN(n13191) );
  NAND2_X1 U16499 ( .A1(n13185), .A2(n13191), .ZN(P1_U2943) );
  AOI22_X1 U16500 ( .A1(n20073), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20072), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13188) );
  INV_X1 U16501 ( .A(DATAI_4_), .ZN(n13187) );
  NAND2_X1 U16502 ( .A1(n20143), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13186) );
  OAI21_X1 U16503 ( .B1(n20143), .B2(n13187), .A(n13186), .ZN(n20169) );
  NAND2_X1 U16504 ( .A1(n20060), .A2(n20169), .ZN(n13195) );
  NAND2_X1 U16505 ( .A1(n13188), .A2(n13195), .ZN(P1_U2941) );
  AOI22_X1 U16506 ( .A1(n20073), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20072), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13190) );
  NAND2_X1 U16507 ( .A1(n13190), .A2(n13189), .ZN(P1_U2955) );
  AOI22_X1 U16508 ( .A1(n20073), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20072), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13192) );
  NAND2_X1 U16509 ( .A1(n13192), .A2(n13191), .ZN(P1_U2958) );
  AOI22_X1 U16510 ( .A1(n20073), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20072), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13194) );
  NAND2_X1 U16511 ( .A1(n13194), .A2(n13193), .ZN(P1_U2959) );
  AOI22_X1 U16512 ( .A1(n20073), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20072), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13196) );
  NAND2_X1 U16513 ( .A1(n13196), .A2(n13195), .ZN(P1_U2956) );
  AOI22_X1 U16514 ( .A1(n20073), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20072), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13198) );
  NAND2_X1 U16515 ( .A1(n13198), .A2(n13197), .ZN(P1_U2957) );
  AOI22_X1 U16516 ( .A1(n20073), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20072), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13201) );
  INV_X1 U16517 ( .A(DATAI_0_), .ZN(n13200) );
  NAND2_X1 U16518 ( .A1(n20143), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13199) );
  OAI21_X1 U16519 ( .B1(n20143), .B2(n13200), .A(n13199), .ZN(n20141) );
  NAND2_X1 U16520 ( .A1(n20060), .A2(n20141), .ZN(n13205) );
  NAND2_X1 U16521 ( .A1(n13201), .A2(n13205), .ZN(P1_U2952) );
  AOI22_X1 U16522 ( .A1(n20073), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20072), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13202) );
  NAND2_X1 U16523 ( .A1(n20060), .A2(n20154), .ZN(n13203) );
  NAND2_X1 U16524 ( .A1(n13202), .A2(n13203), .ZN(P1_U2953) );
  AOI22_X1 U16525 ( .A1(n20073), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20072), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13204) );
  NAND2_X1 U16526 ( .A1(n13204), .A2(n13203), .ZN(P1_U2938) );
  AOI22_X1 U16527 ( .A1(n20073), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20072), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13206) );
  NAND2_X1 U16528 ( .A1(n13206), .A2(n13205), .ZN(P1_U2937) );
  INV_X1 U16529 ( .A(P1_UWORD_REG_10__SCAN_IN), .ZN(n20976) );
  INV_X1 U16530 ( .A(DATAI_10_), .ZN(n13208) );
  NAND2_X1 U16531 ( .A1(n20143), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13207) );
  OAI21_X1 U16532 ( .B1(n20143), .B2(n13208), .A(n13207), .ZN(n14580) );
  NAND2_X1 U16533 ( .A1(n20060), .A2(n14580), .ZN(n20064) );
  NAND2_X1 U16534 ( .A1(n20073), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n13209) );
  OAI211_X1 U16535 ( .C1(n13212), .C2(n20976), .A(n20064), .B(n13209), .ZN(
        P1_U2947) );
  INV_X1 U16536 ( .A(P1_UWORD_REG_8__SCAN_IN), .ZN(n21024) );
  NAND2_X1 U16537 ( .A1(n20073), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n13210) );
  OAI211_X1 U16538 ( .C1(n13212), .C2(n21024), .A(n13211), .B(n13210), .ZN(
        P1_U2945) );
  NAND2_X1 U16539 ( .A1(n15517), .A2(n16345), .ZN(n13216) );
  NAND2_X1 U16540 ( .A1(n19558), .A2(n19845), .ZN(n13214) );
  NAND2_X1 U16541 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19644) );
  INV_X1 U16542 ( .A(n19644), .ZN(n13213) );
  AND2_X1 U16543 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13213), .ZN(
        n13297) );
  INV_X1 U16544 ( .A(n13297), .ZN(n13298) );
  AND2_X1 U16545 ( .A1(n13214), .A2(n13298), .ZN(n19339) );
  AOI22_X1 U16546 ( .A1(n13301), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19825), .B2(n19339), .ZN(n13215) );
  INV_X1 U16547 ( .A(n13220), .ZN(n15500) );
  NAND2_X1 U16548 ( .A1(n15500), .A2(n13221), .ZN(n13222) );
  NAND2_X1 U16549 ( .A1(n13223), .A2(n13222), .ZN(n13225) );
  NAND2_X1 U16550 ( .A1(n13226), .A2(n13225), .ZN(n13227) );
  MUX2_X1 U16551 ( .A(n15517), .B(P2_EBX_REG_2__SCAN_IN), .S(n15040), .Z(
        n13228) );
  AOI21_X1 U16552 ( .B1(n19282), .B2(n15007), .A(n13228), .ZN(n13229) );
  INV_X1 U16553 ( .A(n13229), .ZN(P2_U2885) );
  NOR2_X1 U16554 ( .A1(n19857), .A2(n19062), .ZN(n13232) );
  INV_X1 U16555 ( .A(n19852), .ZN(n13230) );
  NAND2_X1 U16556 ( .A1(n19281), .A2(n13230), .ZN(n13424) );
  OAI21_X1 U16557 ( .B1(n19281), .B2(n13230), .A(n13424), .ZN(n13231) );
  NOR2_X1 U16558 ( .A1(n13231), .A2(n13232), .ZN(n13426) );
  AOI21_X1 U16559 ( .B1(n13232), .B2(n13231), .A(n13426), .ZN(n13236) );
  AOI22_X1 U16560 ( .A1(n13812), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13550), .ZN(n13549) );
  INV_X1 U16561 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n13233) );
  OAI22_X1 U16562 ( .A1(n13593), .A2(n13549), .B1(n19103), .B2(n13233), .ZN(
        n13234) );
  AOI21_X1 U16563 ( .B1(n19087), .B2(n19852), .A(n13234), .ZN(n13235) );
  OAI21_X1 U16564 ( .B1(n13236), .B2(n19107), .A(n13235), .ZN(P2_U2918) );
  MUX2_X1 U16565 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n13550), .Z(n19093) );
  NAND2_X1 U16566 ( .A1(n13287), .A2(n19093), .ZN(n19153) );
  NAND2_X1 U16567 ( .A1(n19151), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13237) );
  OAI211_X1 U16568 ( .C1(n13238), .C2(n13294), .A(n19153), .B(n13237), .ZN(
        P2_U2966) );
  AOI22_X1 U16569 ( .A1(P2_EAX_REG_16__SCAN_IN), .A2(n19152), .B1(n19151), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13239) );
  NAND2_X1 U16570 ( .A1(n13287), .A2(n19081), .ZN(n13259) );
  NAND2_X1 U16571 ( .A1(n13239), .A2(n13259), .ZN(P2_U2952) );
  AOI22_X1 U16572 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n19152), .B1(n19151), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13243) );
  INV_X1 U16573 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13240) );
  OR2_X1 U16574 ( .A1(n13550), .A2(n13240), .ZN(n13242) );
  NAND2_X1 U16575 ( .A1(n13550), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13241) );
  NAND2_X1 U16576 ( .A1(n13242), .A2(n13241), .ZN(n15087) );
  NAND2_X1 U16577 ( .A1(n13287), .A2(n15087), .ZN(n13255) );
  NAND2_X1 U16578 ( .A1(n13243), .A2(n13255), .ZN(P2_U2961) );
  AOI22_X1 U16579 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n19152), .B1(n19151), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13247) );
  INV_X1 U16580 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13244) );
  OR2_X1 U16581 ( .A1(n13811), .A2(n13244), .ZN(n13246) );
  NAND2_X1 U16582 ( .A1(n13550), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13245) );
  NAND2_X1 U16583 ( .A1(n13246), .A2(n13245), .ZN(n15051) );
  NAND2_X1 U16584 ( .A1(n13287), .A2(n15051), .ZN(n13277) );
  NAND2_X1 U16585 ( .A1(n13247), .A2(n13277), .ZN(P2_U2965) );
  AOI22_X1 U16586 ( .A1(n19152), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n19151), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13248) );
  INV_X1 U16587 ( .A(n19243), .ZN(n15094) );
  NAND2_X1 U16588 ( .A1(n13287), .A2(n15094), .ZN(n13261) );
  NAND2_X1 U16589 ( .A1(n13248), .A2(n13261), .ZN(P2_U2959) );
  AOI22_X1 U16590 ( .A1(P2_EAX_REG_22__SCAN_IN), .A2(n19152), .B1(n19151), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13249) );
  INV_X1 U16591 ( .A(n19231), .ZN(n16077) );
  NAND2_X1 U16592 ( .A1(n13287), .A2(n16077), .ZN(n13263) );
  NAND2_X1 U16593 ( .A1(n13249), .A2(n13263), .ZN(P2_U2958) );
  AOI22_X1 U16594 ( .A1(n19152), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n19151), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13250) );
  AOI22_X1 U16595 ( .A1(n13812), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13550), .ZN(n13579) );
  INV_X1 U16596 ( .A(n13579), .ZN(n19105) );
  NAND2_X1 U16597 ( .A1(n13287), .A2(n19105), .ZN(n13265) );
  NAND2_X1 U16598 ( .A1(n13250), .A2(n13265), .ZN(P2_U2957) );
  AOI22_X1 U16599 ( .A1(P2_EAX_REG_20__SCAN_IN), .A2(n19152), .B1(n19151), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13251) );
  OAI22_X1 U16600 ( .A1(n13811), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13812), .ZN(n19225) );
  INV_X1 U16601 ( .A(n19225), .ZN(n16084) );
  NAND2_X1 U16602 ( .A1(n13287), .A2(n16084), .ZN(n13267) );
  NAND2_X1 U16603 ( .A1(n13251), .A2(n13267), .ZN(P2_U2956) );
  AOI22_X1 U16604 ( .A1(n19152), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n19151), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13252) );
  AOI22_X1 U16605 ( .A1(n13812), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13811), .ZN(n19219) );
  INV_X1 U16606 ( .A(n19219), .ZN(n13854) );
  NAND2_X1 U16607 ( .A1(n13287), .A2(n13854), .ZN(n13269) );
  NAND2_X1 U16608 ( .A1(n13252), .A2(n13269), .ZN(P2_U2955) );
  AOI22_X1 U16609 ( .A1(P2_EAX_REG_18__SCAN_IN), .A2(n19152), .B1(n19151), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13253) );
  INV_X1 U16610 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16446) );
  INV_X1 U16611 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18213) );
  AOI22_X1 U16612 ( .A1(n13812), .A2(n16446), .B1(n18213), .B2(n13811), .ZN(
        n19214) );
  NAND2_X1 U16613 ( .A1(n13287), .A2(n19214), .ZN(n13271) );
  NAND2_X1 U16614 ( .A1(n13253), .A2(n13271), .ZN(P2_U2954) );
  AOI22_X1 U16615 ( .A1(n19152), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n19151), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13254) );
  INV_X1 U16616 ( .A(n13549), .ZN(n13816) );
  NAND2_X1 U16617 ( .A1(n13287), .A2(n13816), .ZN(n13257) );
  NAND2_X1 U16618 ( .A1(n13254), .A2(n13257), .ZN(P2_U2953) );
  AOI22_X1 U16619 ( .A1(n19152), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n19151), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13256) );
  NAND2_X1 U16620 ( .A1(n13256), .A2(n13255), .ZN(P2_U2976) );
  AOI22_X1 U16621 ( .A1(n19152), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n19151), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13258) );
  NAND2_X1 U16622 ( .A1(n13258), .A2(n13257), .ZN(P2_U2968) );
  AOI22_X1 U16623 ( .A1(n19152), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n19151), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13260) );
  NAND2_X1 U16624 ( .A1(n13260), .A2(n13259), .ZN(P2_U2967) );
  AOI22_X1 U16625 ( .A1(n19152), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n19151), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13262) );
  NAND2_X1 U16626 ( .A1(n13262), .A2(n13261), .ZN(P2_U2974) );
  AOI22_X1 U16627 ( .A1(n19152), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n19151), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13264) );
  NAND2_X1 U16628 ( .A1(n13264), .A2(n13263), .ZN(P2_U2973) );
  AOI22_X1 U16629 ( .A1(n19152), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n19151), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13266) );
  NAND2_X1 U16630 ( .A1(n13266), .A2(n13265), .ZN(P2_U2972) );
  AOI22_X1 U16631 ( .A1(n19152), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n19151), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13268) );
  NAND2_X1 U16632 ( .A1(n13268), .A2(n13267), .ZN(P2_U2971) );
  AOI22_X1 U16633 ( .A1(n19152), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n19151), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13270) );
  NAND2_X1 U16634 ( .A1(n13270), .A2(n13269), .ZN(P2_U2970) );
  AOI22_X1 U16635 ( .A1(n19152), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n19151), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13272) );
  NAND2_X1 U16636 ( .A1(n13272), .A2(n13271), .ZN(P2_U2969) );
  AOI22_X1 U16637 ( .A1(n19152), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n19151), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13276) );
  INV_X1 U16638 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13273) );
  OR2_X1 U16639 ( .A1(n13550), .A2(n13273), .ZN(n13275) );
  NAND2_X1 U16640 ( .A1(n13550), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13274) );
  NAND2_X1 U16641 ( .A1(n13275), .A2(n13274), .ZN(n15070) );
  NAND2_X1 U16642 ( .A1(n13287), .A2(n15070), .ZN(n13283) );
  NAND2_X1 U16643 ( .A1(n13276), .A2(n13283), .ZN(P2_U2978) );
  AOI22_X1 U16644 ( .A1(n19152), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n19151), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13278) );
  NAND2_X1 U16645 ( .A1(n13278), .A2(n13277), .ZN(P2_U2980) );
  AOI22_X1 U16646 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(n19152), .B1(n19151), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13280) );
  AOI22_X1 U16647 ( .A1(n13812), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n13550), .ZN(n15059) );
  INV_X1 U16648 ( .A(n15059), .ZN(n13279) );
  NAND2_X1 U16649 ( .A1(n13287), .A2(n13279), .ZN(n13281) );
  NAND2_X1 U16650 ( .A1(n13280), .A2(n13281), .ZN(P2_U2964) );
  AOI22_X1 U16651 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19152), .B1(n19151), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13282) );
  NAND2_X1 U16652 ( .A1(n13282), .A2(n13281), .ZN(P2_U2979) );
  AOI22_X1 U16653 ( .A1(P2_EAX_REG_27__SCAN_IN), .A2(n19152), .B1(n19151), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13284) );
  NAND2_X1 U16654 ( .A1(n13284), .A2(n13283), .ZN(P2_U2963) );
  INV_X1 U16655 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n20820) );
  MUX2_X1 U16656 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n13550), .Z(n19096) );
  NAND2_X1 U16657 ( .A1(n13287), .A2(n19096), .ZN(n13293) );
  NAND2_X1 U16658 ( .A1(n19152), .A2(P2_EAX_REG_10__SCAN_IN), .ZN(n13285) );
  OAI211_X1 U16659 ( .C1(n13286), .C2(n20820), .A(n13293), .B(n13285), .ZN(
        P2_U2977) );
  INV_X1 U16660 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20860) );
  INV_X1 U16661 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16438) );
  INV_X1 U16662 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U16663 ( .A1(n13812), .A2(n16438), .B1(n17482), .B2(n13811), .ZN(
        n19099) );
  NAND2_X1 U16664 ( .A1(n13287), .A2(n19099), .ZN(n13290) );
  NAND2_X1 U16665 ( .A1(n19151), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13288) );
  OAI211_X1 U16666 ( .C1(n20860), .C2(n13294), .A(n13290), .B(n13288), .ZN(
        P2_U2975) );
  NAND2_X1 U16667 ( .A1(n19151), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13289) );
  OAI211_X1 U16668 ( .C1(n13291), .C2(n13294), .A(n13290), .B(n13289), .ZN(
        P2_U2960) );
  NAND2_X1 U16669 ( .A1(n19151), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13292) );
  OAI211_X1 U16670 ( .C1(n13295), .C2(n13294), .A(n13293), .B(n13292), .ZN(
        P2_U2962) );
  NAND2_X1 U16671 ( .A1(n13297), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19205) );
  NAND2_X1 U16672 ( .A1(n13299), .A2(n13298), .ZN(n13300) );
  AND3_X1 U16673 ( .A1(n19205), .A2(n19825), .A3(n13300), .ZN(n19588) );
  AOI21_X1 U16674 ( .B1(n13301), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19588), .ZN(n13302) );
  NAND2_X1 U16675 ( .A1(n13381), .A2(n13304), .ZN(n13385) );
  NAND2_X1 U16676 ( .A1(n15040), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13311) );
  NAND2_X1 U16677 ( .A1(n13296), .A2(n14992), .ZN(n13310) );
  OAI211_X1 U16678 ( .C1(n19251), .C2(n15026), .A(n13311), .B(n13310), .ZN(
        P2_U2884) );
  NOR2_X1 U16679 ( .A1(n20107), .A2(n20788), .ZN(n20124) );
  NOR2_X1 U16680 ( .A1(n20085), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13312) );
  AOI211_X1 U16681 ( .C1(n20076), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n20124), .B(n13312), .ZN(n13316) );
  OR2_X1 U16682 ( .A1(n13313), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20127) );
  NAND3_X1 U16683 ( .A1(n20127), .A2(n13314), .A3(n20081), .ZN(n13315) );
  OAI211_X1 U16684 ( .C1(n20142), .C2(n14484), .A(n13316), .B(n13315), .ZN(
        P1_U2998) );
  INV_X1 U16685 ( .A(n15087), .ZN(n13318) );
  INV_X1 U16686 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19130) );
  OAI21_X1 U16687 ( .B1(n16275), .B2(n13317), .A(n15451), .ZN(n18999) );
  OAI222_X1 U16688 ( .A1(n13593), .A2(n13318), .B1(n19103), .B2(n19130), .C1(
        n19113), .C2(n18999), .ZN(P2_U2910) );
  INV_X1 U16689 ( .A(n19251), .ZN(n19830) );
  INV_X1 U16690 ( .A(n15507), .ZN(n15516) );
  INV_X1 U16691 ( .A(n11191), .ZN(n13323) );
  NAND2_X1 U16692 ( .A1(n9741), .A2(n13323), .ZN(n13322) );
  NAND2_X1 U16693 ( .A1(n9827), .A2(n13319), .ZN(n15518) );
  NAND2_X1 U16694 ( .A1(n15518), .A2(n10794), .ZN(n13321) );
  INV_X1 U16695 ( .A(n10788), .ZN(n13320) );
  NAND2_X1 U16696 ( .A1(n13320), .A2(n15527), .ZN(n15515) );
  NAND3_X1 U16697 ( .A1(n13322), .A2(n13321), .A3(n15515), .ZN(n13328) );
  NOR2_X1 U16698 ( .A1(n16314), .A2(n16316), .ZN(n15523) );
  INV_X1 U16699 ( .A(n15515), .ZN(n13325) );
  INV_X1 U16700 ( .A(n10695), .ZN(n13324) );
  OAI22_X1 U16701 ( .A1(n15523), .A2(n13325), .B1(n13324), .B2(n13323), .ZN(
        n13327) );
  MUX2_X1 U16702 ( .A(n13328), .B(n13327), .S(n13326), .Z(n13329) );
  INV_X1 U16703 ( .A(n13329), .ZN(n13330) );
  INV_X1 U16704 ( .A(n14150), .ZN(n14108) );
  NAND2_X1 U16705 ( .A1(n13330), .A2(n14108), .ZN(n13331) );
  AOI21_X1 U16706 ( .B1(n13296), .B2(n15516), .A(n13331), .ZN(n16332) );
  INV_X1 U16707 ( .A(n16332), .ZN(n16310) );
  AOI22_X1 U16708 ( .A1(n19830), .A2(n16352), .B1(n19827), .B2(n16310), .ZN(
        n13333) );
  NAND2_X1 U16709 ( .A1(n15526), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13332) );
  OAI21_X1 U16710 ( .B1(n13333), .B2(n15526), .A(n13332), .ZN(P2_U3596) );
  INV_X1 U16711 ( .A(n13334), .ZN(n13335) );
  AOI21_X1 U16712 ( .B1(n13337), .B2(n13336), .A(n13335), .ZN(n13401) );
  INV_X1 U16713 ( .A(n14561), .ZN(n20008) );
  AND2_X1 U16714 ( .A1(n13339), .A2(n13338), .ZN(n13340) );
  OR2_X1 U16715 ( .A1(n13406), .A2(n13340), .ZN(n20108) );
  OAI22_X1 U16716 ( .A1(n20001), .A2(n20108), .B1(n13341), .B2(n20012), .ZN(
        n13342) );
  AOI21_X1 U16717 ( .B1(n13401), .B2(n20008), .A(n13342), .ZN(n13343) );
  INV_X1 U16718 ( .A(n13343), .ZN(P1_U2870) );
  AOI21_X1 U16719 ( .B1(n15584), .B2(n20707), .A(n13346), .ZN(n13360) );
  INV_X1 U16720 ( .A(n14031), .ZN(n14878) );
  XNOR2_X1 U16721 ( .A(n13344), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13356) );
  MUX2_X1 U16722 ( .A(n13345), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n14884), .Z(n13347) );
  NOR2_X1 U16723 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  NAND2_X1 U16724 ( .A1(n13349), .A2(n13348), .ZN(n13355) );
  AOI21_X1 U16725 ( .B1(n14884), .B2(n9746), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13350) );
  NOR2_X1 U16726 ( .A1(n13351), .A2(n13350), .ZN(n14890) );
  NAND3_X1 U16727 ( .A1(n13353), .A2(n13352), .A3(n14890), .ZN(n13354) );
  OAI211_X1 U16728 ( .C1(n14878), .C2(n13356), .A(n13355), .B(n13354), .ZN(
        n13357) );
  AOI21_X1 U16729 ( .B1(n20399), .B2(n14882), .A(n13357), .ZN(n15582) );
  OAI21_X1 U16730 ( .B1(n15582), .B2(n15579), .A(n15584), .ZN(n13358) );
  INV_X1 U16731 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19901) );
  AND2_X1 U16732 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n19901), .ZN(n13365) );
  AOI21_X1 U16733 ( .B1(n13358), .B2(n20707), .A(n13365), .ZN(n13359) );
  OR2_X1 U16734 ( .A1(n13360), .A2(n13359), .ZN(n15587) );
  NAND2_X1 U16735 ( .A1(n19963), .A2(n13362), .ZN(n13363) );
  NAND2_X1 U16736 ( .A1(n15584), .A2(n13363), .ZN(n13364) );
  OAI211_X1 U16737 ( .C1(n15584), .C2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13364), .B(n20707), .ZN(n13367) );
  NAND2_X1 U16738 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13365), .ZN(
        n13366) );
  AND2_X1 U16739 ( .A1(n13367), .A2(n13366), .ZN(n15588) );
  OAI21_X1 U16740 ( .B1(n15587), .B2(n13361), .A(n15588), .ZN(n14873) );
  OR2_X1 U16741 ( .A1(n14873), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n13369) );
  NAND2_X1 U16742 ( .A1(n13369), .A2(n13368), .ZN(n13370) );
  NOR2_X1 U16743 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20801) );
  INV_X1 U16744 ( .A(n20801), .ZN(n15976) );
  AND2_X1 U16745 ( .A1(n13370), .A2(n20294), .ZN(n20136) );
  INV_X1 U16746 ( .A(n20136), .ZN(n14036) );
  NAND2_X1 U16747 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20532), .ZN(n14874) );
  NAND2_X1 U16748 ( .A1(n14036), .A2(n14874), .ZN(n14063) );
  INV_X1 U16749 ( .A(n20399), .ZN(n13377) );
  NOR2_X1 U16750 ( .A1(n20136), .A2(n20644), .ZN(n14060) );
  INV_X1 U16751 ( .A(n14060), .ZN(n14038) );
  NAND2_X1 U16752 ( .A1(n20223), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20650) );
  INV_X1 U16753 ( .A(n20650), .ZN(n20259) );
  NAND2_X1 U16754 ( .A1(n20370), .A2(n20259), .ZN(n20375) );
  NAND2_X1 U16755 ( .A1(n20375), .A2(n20493), .ZN(n13375) );
  OR2_X1 U16756 ( .A1(n20223), .A2(n21079), .ZN(n20431) );
  NOR2_X1 U16757 ( .A1(n20651), .A2(n20431), .ZN(n20571) );
  AOI211_X1 U16758 ( .C1(n12027), .C2(n21079), .A(n13375), .B(n20571), .ZN(
        n13376) );
  OAI222_X1 U16759 ( .A1(n14036), .A2(n20488), .B1(n14063), .B2(n13377), .C1(
        n14038), .C2(n13376), .ZN(P1_U3475) );
  INV_X1 U16760 ( .A(n13401), .ZN(n19980) );
  INV_X1 U16761 ( .A(n20159), .ZN(n13378) );
  INV_X1 U16762 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20046) );
  OAI222_X1 U16763 ( .A1(n19980), .A2(n20016), .B1(n20014), .B2(n13378), .C1(
        n20015), .C2(n20046), .ZN(P1_U2902) );
  NAND2_X1 U16764 ( .A1(n10657), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13379) );
  INV_X1 U16765 ( .A(n13383), .ZN(n13384) );
  NAND2_X1 U16766 ( .A1(n13385), .A2(n13384), .ZN(n13386) );
  OR2_X1 U16767 ( .A1(n13387), .A2(n13386), .ZN(n13388) );
  NAND2_X1 U16768 ( .A1(n13447), .A2(n13388), .ZN(n19108) );
  NAND2_X1 U16769 ( .A1(n13390), .A2(n13389), .ZN(n13391) );
  AND2_X1 U16770 ( .A1(n13391), .A2(n9858), .ZN(n19193) );
  INV_X1 U16771 ( .A(n19193), .ZN(n19048) );
  MUX2_X1 U16772 ( .A(n13392), .B(n19048), .S(n14992), .Z(n13393) );
  OAI21_X1 U16773 ( .B1(n19108), .B2(n15026), .A(n13393), .ZN(P2_U2883) );
  OAI21_X1 U16774 ( .B1(n13396), .B2(n13395), .A(n13394), .ZN(n20106) );
  INV_X1 U16775 ( .A(n19983), .ZN(n13399) );
  AOI22_X1 U16776 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13398) );
  OAI21_X1 U16777 ( .B1(n20085), .B2(n13399), .A(n13398), .ZN(n13400) );
  AOI21_X1 U16778 ( .B1(n13401), .B2(n14666), .A(n13400), .ZN(n13402) );
  OAI21_X1 U16779 ( .B1(n19900), .B2(n20106), .A(n13402), .ZN(P1_U2997) );
  XOR2_X1 U16780 ( .A(n13403), .B(n13404), .Z(n13414) );
  INV_X1 U16781 ( .A(n13414), .ZN(n14482) );
  OR2_X1 U16782 ( .A1(n13406), .A2(n13405), .ZN(n13407) );
  AND2_X1 U16783 ( .A1(n13444), .A2(n13407), .ZN(n20095) );
  INV_X1 U16784 ( .A(n20012), .ZN(n14520) );
  AOI22_X1 U16785 ( .A1(n20007), .A2(n20095), .B1(n14520), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13408) );
  OAI21_X1 U16786 ( .B1(n14482), .B2(n14561), .A(n13408), .ZN(P1_U2869) );
  OAI21_X1 U16787 ( .B1(n9748), .B2(n13410), .A(n13409), .ZN(n20096) );
  NAND2_X1 U16788 ( .A1(n13397), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n20093) );
  NAND2_X1 U16789 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13412) );
  OAI211_X1 U16790 ( .C1(n20085), .C2(n14477), .A(n20093), .B(n13412), .ZN(
        n13413) );
  AOI21_X1 U16791 ( .B1(n13414), .B2(n14666), .A(n13413), .ZN(n13415) );
  OAI21_X1 U16792 ( .B1(n20096), .B2(n19900), .A(n13415), .ZN(P1_U2996) );
  XOR2_X1 U16793 ( .A(n13447), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13422)
         );
  INV_X1 U16794 ( .A(n13416), .ZN(n13417) );
  NAND2_X1 U16795 ( .A1(n13417), .A2(n9858), .ZN(n13418) );
  AND2_X1 U16796 ( .A1(n13418), .A2(n13455), .ZN(n19035) );
  NOR2_X1 U16797 ( .A1(n14992), .A2(n13419), .ZN(n13420) );
  AOI21_X1 U16798 ( .B1(n19035), .B2(n14992), .A(n13420), .ZN(n13421) );
  OAI21_X1 U16799 ( .B1(n13422), .B2(n15026), .A(n13421), .ZN(P2_U2882) );
  INV_X1 U16800 ( .A(n20164), .ZN(n13423) );
  INV_X1 U16801 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20888) );
  OAI222_X1 U16802 ( .A1(n14482), .A2(n20016), .B1(n20014), .B2(n13423), .C1(
        n20015), .C2(n20888), .ZN(P1_U2901) );
  INV_X1 U16803 ( .A(n13424), .ZN(n13425) );
  NOR2_X1 U16804 ( .A1(n13426), .A2(n13425), .ZN(n13434) );
  INV_X1 U16805 ( .A(n19282), .ZN(n19841) );
  NAND2_X1 U16806 ( .A1(n13428), .A2(n13427), .ZN(n13431) );
  INV_X1 U16807 ( .A(n13429), .ZN(n13430) );
  NAND2_X1 U16808 ( .A1(n13431), .A2(n13430), .ZN(n19843) );
  INV_X1 U16809 ( .A(n19843), .ZN(n13432) );
  NAND2_X1 U16810 ( .A1(n19841), .A2(n13432), .ZN(n13473) );
  OAI21_X1 U16811 ( .B1(n19841), .B2(n13432), .A(n13473), .ZN(n13433) );
  NOR2_X1 U16812 ( .A1(n13434), .A2(n13433), .ZN(n13475) );
  AOI21_X1 U16813 ( .B1(n13434), .B2(n13433), .A(n13475), .ZN(n13437) );
  AOI22_X1 U16814 ( .A1(n19106), .A2(n19214), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19104), .ZN(n13436) );
  NAND2_X1 U16815 ( .A1(n19843), .A2(n19087), .ZN(n13435) );
  OAI211_X1 U16816 ( .C1(n13437), .C2(n19107), .A(n13436), .B(n13435), .ZN(
        P2_U2917) );
  INV_X1 U16817 ( .A(n13438), .ZN(n13441) );
  INV_X1 U16818 ( .A(n13439), .ZN(n13440) );
  NAND2_X1 U16819 ( .A1(n13441), .A2(n13440), .ZN(n13442) );
  AND2_X1 U16820 ( .A1(n13442), .A2(n13468), .ZN(n20080) );
  INV_X1 U16821 ( .A(n20080), .ZN(n13463) );
  AOI21_X1 U16822 ( .B1(n13445), .B2(n13444), .A(n13443), .ZN(n20088) );
  AOI22_X1 U16823 ( .A1(n20007), .A2(n20088), .B1(n14520), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13446) );
  OAI21_X1 U16824 ( .B1(n13463), .B2(n14561), .A(n13446), .ZN(P1_U2868) );
  XNOR2_X1 U16825 ( .A(n13485), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13451) );
  INV_X1 U16826 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13449) );
  OAI21_X1 U16827 ( .B1(n13448), .B2(n13457), .A(n13487), .ZN(n15476) );
  MUX2_X1 U16828 ( .A(n13449), .B(n15476), .S(n14992), .Z(n13450) );
  OAI21_X1 U16829 ( .B1(n13451), .B2(n15026), .A(n13450), .ZN(P2_U2880) );
  NOR2_X1 U16830 ( .A1(n13447), .A2(n13452), .ZN(n13454) );
  INV_X1 U16831 ( .A(n13485), .ZN(n13453) );
  OAI211_X1 U16832 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13454), .A(
        n13453), .B(n15007), .ZN(n13460) );
  NAND2_X1 U16833 ( .A1(n13456), .A2(n13455), .ZN(n13458) );
  NAND2_X1 U16834 ( .A1(n13458), .A2(n10195), .ZN(n15259) );
  INV_X1 U16835 ( .A(n15259), .ZN(n19021) );
  NAND2_X1 U16836 ( .A1(n19021), .A2(n14992), .ZN(n13459) );
  OAI211_X1 U16837 ( .C1(n14992), .C2(n13461), .A(n13460), .B(n13459), .ZN(
        P2_U2881) );
  INV_X1 U16838 ( .A(n20169), .ZN(n13462) );
  INV_X1 U16839 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20042) );
  OAI222_X1 U16840 ( .A1(n20016), .A2(n13463), .B1(n20014), .B2(n13462), .C1(
        n20015), .C2(n20042), .ZN(P1_U2900) );
  INV_X1 U16841 ( .A(n15070), .ZN(n13466) );
  INV_X1 U16842 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19127) );
  OAI21_X1 U16843 ( .B1(n13465), .B2(n13464), .A(n13472), .ZN(n18980) );
  OAI222_X1 U16844 ( .A1(n13593), .A2(n13466), .B1(n19103), .B2(n19127), .C1(
        n18980), .C2(n19113), .ZN(P2_U2908) );
  AND2_X1 U16845 ( .A1(n13468), .A2(n13467), .ZN(n13469) );
  OR2_X1 U16846 ( .A1(n13469), .A2(n13499), .ZN(n15847) );
  INV_X1 U16847 ( .A(n20175), .ZN(n13470) );
  OAI222_X1 U16848 ( .A1(n15847), .A2(n20016), .B1(n20014), .B2(n13470), .C1(
        n20015), .C2(n12080), .ZN(P1_U2899) );
  XNOR2_X1 U16849 ( .A(n13472), .B(n13471), .ZN(n18968) );
  INV_X1 U16850 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19125) );
  OAI222_X1 U16851 ( .A1(n13593), .A2(n15059), .B1(n18968), .B2(n19113), .C1(
        n19125), .C2(n19103), .ZN(P2_U2907) );
  INV_X1 U16852 ( .A(n13473), .ZN(n13474) );
  NOR2_X1 U16853 ( .A1(n13475), .A2(n13474), .ZN(n13481) );
  OR2_X1 U16854 ( .A1(n13477), .A2(n13476), .ZN(n13479) );
  NAND2_X1 U16855 ( .A1(n13479), .A2(n13478), .ZN(n16288) );
  XNOR2_X1 U16856 ( .A(n19251), .B(n16288), .ZN(n13480) );
  NOR2_X1 U16857 ( .A1(n13481), .A2(n13480), .ZN(n13563) );
  AOI21_X1 U16858 ( .B1(n13481), .B2(n13480), .A(n13563), .ZN(n13484) );
  INV_X1 U16859 ( .A(n16288), .ZN(n19832) );
  AOI22_X1 U16860 ( .A1(n19087), .A2(n19832), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19104), .ZN(n13483) );
  NAND2_X1 U16861 ( .A1(n19106), .A2(n13854), .ZN(n13482) );
  OAI211_X1 U16862 ( .C1(n13484), .C2(n19107), .A(n13483), .B(n13482), .ZN(
        P2_U2916) );
  OAI211_X1 U16863 ( .C1(n10235), .C2(n13486), .A(n15007), .B(n13528), .ZN(
        n13490) );
  AOI21_X1 U16864 ( .B1(n13488), .B2(n13487), .A(n13492), .ZN(n19010) );
  NAND2_X1 U16865 ( .A1(n19010), .A2(n14992), .ZN(n13489) );
  OAI211_X1 U16866 ( .C1(n14992), .C2(n13491), .A(n13490), .B(n13489), .ZN(
        P2_U2879) );
  INV_X1 U16867 ( .A(n13518), .ZN(n13527) );
  XNOR2_X1 U16868 ( .A(n13528), .B(n13527), .ZN(n13497) );
  NOR2_X1 U16869 ( .A1(n13493), .A2(n13492), .ZN(n13494) );
  NOR2_X1 U16870 ( .A1(n13533), .A2(n13494), .ZN(n16181) );
  INV_X1 U16871 ( .A(n16181), .ZN(n18998) );
  MUX2_X1 U16872 ( .A(n13495), .B(n18998), .S(n14992), .Z(n13496) );
  OAI21_X1 U16873 ( .B1(n13497), .B2(n15026), .A(n13496), .ZN(P2_U2878) );
  XOR2_X1 U16874 ( .A(n13499), .B(n13498), .Z(n19950) );
  INV_X1 U16875 ( .A(n19950), .ZN(n13515) );
  XOR2_X1 U16876 ( .A(n13500), .B(n15967), .Z(n19941) );
  AOI22_X1 U16877 ( .A1(n20007), .A2(n19941), .B1(n14520), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n13501) );
  OAI21_X1 U16878 ( .B1(n13515), .B2(n14561), .A(n13501), .ZN(P1_U2866) );
  NAND2_X1 U16879 ( .A1(n13504), .A2(n13503), .ZN(n13505) );
  AND2_X1 U16880 ( .A1(n13502), .A2(n13505), .ZN(n19937) );
  OR2_X1 U16881 ( .A1(n13508), .A2(n13507), .ZN(n13509) );
  AND2_X1 U16882 ( .A1(n13506), .A2(n13509), .ZN(n19929) );
  INV_X1 U16883 ( .A(n19929), .ZN(n13511) );
  OAI22_X1 U16884 ( .A1(n20001), .A2(n13511), .B1(n13510), .B2(n20012), .ZN(
        n13512) );
  AOI21_X1 U16885 ( .B1(n19937), .B2(n20008), .A(n13512), .ZN(n13513) );
  INV_X1 U16886 ( .A(n13513), .ZN(P1_U2865) );
  INV_X1 U16887 ( .A(n20180), .ZN(n13514) );
  INV_X1 U16888 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20039) );
  OAI222_X1 U16889 ( .A1(n20016), .A2(n13515), .B1(n20014), .B2(n13514), .C1(
        n20015), .C2(n20039), .ZN(P1_U2898) );
  INV_X1 U16890 ( .A(n19937), .ZN(n13517) );
  INV_X1 U16891 ( .A(n20186), .ZN(n13516) );
  OAI222_X1 U16892 ( .A1(n13517), .A2(n20016), .B1(n20014), .B2(n13516), .C1(
        n20015), .C2(n12112), .ZN(P1_U2897) );
  NAND2_X1 U16893 ( .A1(n13518), .A2(n13530), .ZN(n13519) );
  XNOR2_X1 U16894 ( .A(n13558), .B(n13652), .ZN(n13523) );
  OAI21_X1 U16895 ( .B1(n13535), .B2(n13520), .A(n13647), .ZN(n18975) );
  MUX2_X1 U16896 ( .A(n13521), .B(n18975), .S(n14992), .Z(n13522) );
  OAI21_X1 U16897 ( .B1(n13523), .B2(n15026), .A(n13522), .ZN(P2_U2876) );
  INV_X1 U16898 ( .A(n15051), .ZN(n13526) );
  XOR2_X1 U16899 ( .A(n13525), .B(n13524), .Z(n15429) );
  INV_X1 U16900 ( .A(n15429), .ZN(n13718) );
  INV_X1 U16901 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19123) );
  OAI222_X1 U16902 ( .A1(n13593), .A2(n13526), .B1(n13718), .B2(n19113), .C1(
        n19123), .C2(n19103), .ZN(P2_U2906) );
  INV_X1 U16903 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13538) );
  NOR2_X1 U16904 ( .A1(n13528), .A2(n13527), .ZN(n13531) );
  INV_X1 U16905 ( .A(n13558), .ZN(n13529) );
  OAI211_X1 U16906 ( .C1(n13531), .C2(n13530), .A(n13529), .B(n15007), .ZN(
        n13537) );
  NOR2_X1 U16907 ( .A1(n13533), .A2(n13532), .ZN(n13534) );
  NOR2_X1 U16908 ( .A1(n13535), .A2(n13534), .ZN(n18989) );
  NAND2_X1 U16909 ( .A1(n18989), .A2(n14992), .ZN(n13536) );
  OAI211_X1 U16910 ( .C1(n14992), .C2(n13538), .A(n13537), .B(n13536), .ZN(
        P2_U2877) );
  NOR2_X1 U16911 ( .A1(n19251), .A2(n19882), .ZN(n19561) );
  NAND2_X1 U16912 ( .A1(n19561), .A2(n13552), .ZN(n13545) );
  OR2_X1 U16913 ( .A1(n13299), .A2(n19644), .ZN(n13546) );
  INV_X1 U16914 ( .A(n19205), .ZN(n19727) );
  NAND2_X1 U16915 ( .A1(n15639), .A2(n13540), .ZN(n13541) );
  OAI211_X1 U16916 ( .C1(n19727), .C2(n19871), .A(n13548), .B(n19651), .ZN(
        n13544) );
  AOI21_X1 U16917 ( .B1(n13545), .B2(n13546), .A(n13544), .ZN(n19695) );
  OAI21_X1 U16918 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n13546), .A(n19872), 
        .ZN(n13547) );
  AND2_X1 U16919 ( .A1(n13548), .A2(n13547), .ZN(n19729) );
  NOR2_X2 U16920 ( .A1(n13549), .A2(n19498), .ZN(n19664) );
  INV_X1 U16921 ( .A(n19240), .ZN(n13586) );
  INV_X1 U16922 ( .A(n19662), .ZN(n13554) );
  AOI22_X1 U16923 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19235), .ZN(n19605) );
  INV_X1 U16924 ( .A(n19605), .ZN(n19663) );
  AOI22_X1 U16925 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19235), .ZN(n19667) );
  AOI22_X1 U16926 ( .A1(n19721), .A2(n19663), .B1(n19731), .B2(n19602), .ZN(
        n13553) );
  OAI21_X1 U16927 ( .B1(n13554), .B2(n19205), .A(n13553), .ZN(n13555) );
  AOI21_X1 U16928 ( .B1(n19729), .B2(n19664), .A(n13555), .ZN(n13556) );
  OAI21_X1 U16929 ( .B1(n19695), .B2(n14175), .A(n13556), .ZN(P2_U3169) );
  AND2_X1 U16930 ( .A1(n13652), .A2(n13651), .ZN(n13557) );
  XNOR2_X1 U16931 ( .A(n13635), .B(n13633), .ZN(n13562) );
  INV_X1 U16932 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13560) );
  OAI21_X1 U16933 ( .B1(n13559), .B2(n13649), .A(n13639), .ZN(n16140) );
  MUX2_X1 U16934 ( .A(n13560), .B(n16140), .S(n14992), .Z(n13561) );
  OAI21_X1 U16935 ( .B1(n13562), .B2(n15026), .A(n13561), .ZN(P2_U2874) );
  AOI21_X1 U16936 ( .B1(n16288), .B2(n19251), .A(n13563), .ZN(n13569) );
  INV_X1 U16937 ( .A(n13478), .ZN(n13564) );
  OR2_X1 U16938 ( .A1(n13565), .A2(n13564), .ZN(n13568) );
  INV_X1 U16939 ( .A(n13566), .ZN(n13567) );
  AND2_X1 U16940 ( .A1(n13568), .A2(n13567), .ZN(n19185) );
  NOR2_X1 U16941 ( .A1(n13569), .A2(n19185), .ZN(n19109) );
  XOR2_X1 U16942 ( .A(n19108), .B(n19109), .Z(n13570) );
  NAND2_X1 U16943 ( .A1(n13570), .A2(n16079), .ZN(n13572) );
  AOI22_X1 U16944 ( .A1(n19087), .A2(n19185), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19104), .ZN(n13571) );
  OAI211_X1 U16945 ( .C1(n19225), .C2(n13593), .A(n13572), .B(n13571), .ZN(
        P2_U2915) );
  NAND2_X1 U16946 ( .A1(n19561), .A2(n19369), .ZN(n13576) );
  NAND3_X1 U16947 ( .A1(n10893), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19589) );
  NOR2_X1 U16948 ( .A1(n19861), .A2(n19589), .ZN(n19648) );
  INV_X1 U16949 ( .A(n19648), .ZN(n13588) );
  AND2_X1 U16950 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13588), .ZN(n13573) );
  NAND2_X1 U16951 ( .A1(n13574), .A2(n13573), .ZN(n13578) );
  OAI211_X1 U16952 ( .C1(n19871), .C2(n19648), .A(n13578), .B(n19651), .ZN(
        n13575) );
  AOI21_X1 U16953 ( .B1(n13576), .B2(n19589), .A(n13575), .ZN(n19634) );
  OAI21_X1 U16954 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19589), .A(n19872), 
        .ZN(n13577) );
  NOR2_X2 U16955 ( .A1(n13579), .A2(n19498), .ZN(n19713) );
  NOR2_X2 U16956 ( .A1(n9755), .A2(n19240), .ZN(n19712) );
  INV_X1 U16957 ( .A(n19712), .ZN(n13582) );
  INV_X1 U16958 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n17248) );
  INV_X1 U16959 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20924) );
  OAI22_X2 U16960 ( .A1(n17248), .A2(n19236), .B1(n20924), .B2(n19238), .ZN(
        n19679) );
  AOI22_X1 U16961 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19235), .ZN(n19682) );
  INV_X1 U16962 ( .A(n19682), .ZN(n19714) );
  AOI22_X1 U16963 ( .A1(n19630), .A2(n19679), .B1(n19678), .B2(n19714), .ZN(
        n13581) );
  OAI21_X1 U16964 ( .B1(n13582), .B2(n13588), .A(n13581), .ZN(n13583) );
  AOI21_X1 U16965 ( .B1(n19639), .B2(n19713), .A(n13583), .ZN(n13584) );
  OAI21_X1 U16966 ( .B1(n19634), .B2(n14081), .A(n13584), .ZN(P2_U3157) );
  INV_X1 U16967 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13591) );
  NOR2_X2 U16968 ( .A1(n13585), .A2(n19498), .ZN(n19658) );
  AND2_X1 U16969 ( .A1(n19883), .A2(n13586), .ZN(n19645) );
  INV_X1 U16970 ( .A(n19645), .ZN(n13595) );
  AOI22_X1 U16971 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19235), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19234), .ZN(n19661) );
  AOI22_X1 U16972 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19235), .ZN(n19601) );
  INV_X1 U16973 ( .A(n19601), .ZN(n19646) );
  AOI22_X1 U16974 ( .A1(n19630), .A2(n19598), .B1(n19678), .B2(n19646), .ZN(
        n13587) );
  OAI21_X1 U16975 ( .B1(n13595), .B2(n13588), .A(n13587), .ZN(n13589) );
  AOI21_X1 U16976 ( .B1(n19639), .B2(n19658), .A(n13589), .ZN(n13590) );
  OAI21_X1 U16977 ( .B1(n19634), .B2(n13591), .A(n13590), .ZN(P2_U3152) );
  OAI222_X1 U16978 ( .A1(n13593), .A2(n13592), .B1(n19103), .B2(n19120), .C1(
        n19113), .C2(n16236), .ZN(P2_U2904) );
  INV_X1 U16979 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13749) );
  AOI22_X1 U16980 ( .A1(n19731), .A2(n19598), .B1(n19721), .B2(n19646), .ZN(
        n13594) );
  OAI21_X1 U16981 ( .B1(n13595), .B2(n19205), .A(n13594), .ZN(n13596) );
  AOI21_X1 U16982 ( .B1(n19729), .B2(n19658), .A(n13596), .ZN(n13597) );
  OAI21_X1 U16983 ( .B1(n19695), .B2(n13749), .A(n13597), .ZN(P2_U3168) );
  XNOR2_X1 U16984 ( .A(n13599), .B(n13598), .ZN(n16292) );
  XNOR2_X1 U16985 ( .A(n13601), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13602) );
  XNOR2_X1 U16986 ( .A(n13600), .B(n13602), .ZN(n16294) );
  NAND2_X1 U16987 ( .A1(n16294), .A2(n19175), .ZN(n13606) );
  NAND2_X1 U16988 ( .A1(n16198), .A2(n13659), .ZN(n13603) );
  NAND2_X1 U16989 ( .A1(n19029), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16287) );
  OAI211_X1 U16990 ( .C1(n13661), .C2(n16204), .A(n13603), .B(n16287), .ZN(
        n13604) );
  AOI21_X1 U16991 ( .B1(n13296), .B2(n19171), .A(n13604), .ZN(n13605) );
  OAI211_X1 U16992 ( .C1(n16292), .C2(n19177), .A(n13606), .B(n13605), .ZN(
        P2_U3011) );
  INV_X1 U16993 ( .A(n13607), .ZN(n13608) );
  AOI21_X1 U16994 ( .B1(n13609), .B2(n13502), .A(n13608), .ZN(n13743) );
  INV_X1 U16995 ( .A(n13743), .ZN(n13706) );
  AOI22_X1 U16996 ( .A1(n15770), .A2(n14589), .B1(n15768), .B2(
        P1_EAX_REG_8__SCAN_IN), .ZN(n13610) );
  OAI21_X1 U16997 ( .B1(n13706), .B2(n20016), .A(n13610), .ZN(P1_U2896) );
  NAND2_X1 U16998 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20801), .ZN(n15598) );
  NAND2_X1 U16999 ( .A1(n13611), .A2(n15605), .ZN(n13612) );
  OAI211_X1 U17000 ( .C1(n15598), .C2(n20708), .A(n20107), .B(n13612), .ZN(
        n13613) );
  INV_X1 U17001 ( .A(n13613), .ZN(n13614) );
  NOR2_X1 U17002 ( .A1(n13616), .A2(n20707), .ZN(n13617) );
  NAND2_X1 U17003 ( .A1(n13743), .A2(n19949), .ZN(n13632) );
  INV_X1 U17004 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20737) );
  NAND3_X1 U17005 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n14467) );
  NOR2_X1 U17006 ( .A1(n20737), .A2(n14467), .ZN(n13865) );
  INV_X1 U17007 ( .A(n14417), .ZN(n19974) );
  INV_X1 U17008 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20728) );
  NAND2_X1 U17009 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n19984) );
  NOR2_X1 U17010 ( .A1(n20728), .A2(n19984), .ZN(n19965) );
  NAND2_X1 U17011 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n19965), .ZN(n13866) );
  NOR2_X1 U17012 ( .A1(n19974), .A2(n13866), .ZN(n13869) );
  OR2_X1 U17013 ( .A1(n14475), .A2(n20144), .ZN(n13620) );
  AND2_X1 U17014 ( .A1(n15977), .A2(n21079), .ZN(n15569) );
  INV_X1 U17015 ( .A(n15569), .ZN(n13618) );
  AOI21_X1 U17016 ( .B1(n12606), .B2(n15624), .A(n13618), .ZN(n13624) );
  NAND2_X1 U17017 ( .A1(n15662), .A2(n14417), .ZN(n19989) );
  AOI21_X1 U17018 ( .B1(n13865), .B2(n13869), .A(n15647), .ZN(n19922) );
  OR2_X1 U17019 ( .A1(n15662), .A2(n13866), .ZN(n19959) );
  NOR2_X1 U17020 ( .A1(n14467), .A2(n19959), .ZN(n13630) );
  AND2_X1 U17021 ( .A1(n20155), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13623) );
  NAND2_X1 U17022 ( .A1(n13623), .A2(n13618), .ZN(n13619) );
  NOR2_X2 U17023 ( .A1(n13620), .A2(n13619), .ZN(n19991) );
  NAND2_X1 U17024 ( .A1(n13506), .A2(n13621), .ZN(n13622) );
  NAND2_X1 U17025 ( .A1(n15935), .A2(n13622), .ZN(n15950) );
  NOR2_X1 U17026 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  AOI22_X1 U17027 ( .A1(n19994), .A2(P1_EBX_REG_8__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19975), .ZN(n13628) );
  NAND2_X1 U17028 ( .A1(n14417), .A2(n13627), .ZN(n19954) );
  OAI211_X1 U17029 ( .C1(n19988), .C2(n15950), .A(n13628), .B(n19954), .ZN(
        n13629) );
  AOI221_X1 U17030 ( .B1(n19922), .B2(P1_REIP_REG_8__SCAN_IN), .C1(n13630), 
        .C2(n20737), .A(n13629), .ZN(n13631) );
  OAI211_X1 U17031 ( .C1(n13741), .C2(n19992), .A(n13632), .B(n13631), .ZN(
        P1_U2832) );
  AND2_X1 U17032 ( .A1(n13635), .A2(n13633), .ZN(n13637) );
  AND2_X1 U17033 ( .A1(n13633), .A2(n13636), .ZN(n13634) );
  INV_X1 U17034 ( .A(n9838), .ZN(n13746) );
  OAI211_X1 U17035 ( .C1(n13637), .C2(n13636), .A(n15007), .B(n13746), .ZN(
        n13642) );
  AOI21_X1 U17036 ( .B1(n13640), .B2(n13639), .A(n13638), .ZN(n18953) );
  NAND2_X1 U17037 ( .A1(n18953), .A2(n14992), .ZN(n13641) );
  OAI211_X1 U17038 ( .C1(n14992), .C2(n11294), .A(n13642), .B(n13641), .ZN(
        P2_U2873) );
  OAI21_X1 U17039 ( .B1(n13721), .B2(n13645), .A(n13644), .ZN(n13726) );
  AOI22_X1 U17040 ( .A1(n15770), .A2(n14580), .B1(n15768), .B2(
        P1_EAX_REG_10__SCAN_IN), .ZN(n13646) );
  OAI21_X1 U17041 ( .B1(n13726), .B2(n20016), .A(n13646), .ZN(P1_U2894) );
  NAND2_X1 U17042 ( .A1(n13648), .A2(n13647), .ZN(n13650) );
  INV_X1 U17043 ( .A(n18964), .ZN(n13656) );
  AOI21_X1 U17044 ( .B1(n13558), .B2(n13652), .A(n13651), .ZN(n13653) );
  OR3_X1 U17045 ( .A1(n13635), .A2(n13653), .A3(n15026), .ZN(n13655) );
  NAND2_X1 U17046 ( .A1(n15040), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13654) );
  OAI211_X1 U17047 ( .C1(n13656), .C2(n15040), .A(n13655), .B(n13654), .ZN(
        P2_U2875) );
  NAND2_X1 U17048 ( .A1(n19032), .A2(n13657), .ZN(n13658) );
  XNOR2_X1 U17049 ( .A(n13659), .B(n13658), .ZN(n13660) );
  NAND2_X1 U17050 ( .A1(n13660), .A2(n19036), .ZN(n13669) );
  INV_X1 U17051 ( .A(n19065), .ZN(n19014) );
  OAI22_X1 U17052 ( .A1(n19014), .A2(n13662), .B1(n13661), .B2(n19072), .ZN(
        n13664) );
  INV_X1 U17053 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19766) );
  NOR2_X1 U17054 ( .A1(n19061), .A2(n19766), .ZN(n13663) );
  AOI211_X1 U17055 ( .C1(n19832), .C2(n19042), .A(n13664), .B(n13663), .ZN(
        n13665) );
  OAI21_X1 U17056 ( .B1(n13666), .B2(n19067), .A(n13665), .ZN(n13667) );
  AOI21_X1 U17057 ( .B1(n13296), .B2(n19070), .A(n13667), .ZN(n13668) );
  OAI211_X1 U17058 ( .C1(n19251), .C2(n19049), .A(n13669), .B(n13668), .ZN(
        P2_U2852) );
  INV_X1 U17059 ( .A(n13672), .ZN(n14006) );
  NOR2_X1 U17060 ( .A1(n19052), .A2(n13670), .ZN(n13701) );
  INV_X1 U17061 ( .A(n13701), .ZN(n13671) );
  AOI221_X1 U17062 ( .B1(n14006), .B2(n13701), .C1(n13672), .C2(n13671), .A(
        n19741), .ZN(n13673) );
  INV_X1 U17063 ( .A(n13673), .ZN(n13682) );
  INV_X1 U17064 ( .A(n13674), .ZN(n13677) );
  AOI22_X1 U17065 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n19043), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(n19065), .ZN(n13676) );
  NAND2_X1 U17066 ( .A1(n19030), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13675) );
  OAI211_X1 U17067 ( .C1(n19067), .C2(n13677), .A(n13676), .B(n13675), .ZN(
        n13680) );
  NOR2_X1 U17068 ( .A1(n13678), .A2(n19047), .ZN(n13679) );
  AOI211_X1 U17069 ( .C1(n19042), .C2(n19843), .A(n13680), .B(n13679), .ZN(
        n13681) );
  OAI211_X1 U17070 ( .C1(n19841), .C2(n19049), .A(n13682), .B(n13681), .ZN(
        P2_U2853) );
  NAND2_X1 U17071 ( .A1(n19032), .A2(n13683), .ZN(n13684) );
  XNOR2_X1 U17072 ( .A(n15249), .B(n13684), .ZN(n13691) );
  NOR2_X1 U17073 ( .A1(n15477), .A2(n19063), .ZN(n13690) );
  AOI22_X1 U17074 ( .A1(n13685), .A2(n19041), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19043), .ZN(n13686) );
  OAI211_X1 U17075 ( .C1(n19771), .C2(n19061), .A(n13686), .B(n19045), .ZN(
        n13687) );
  AOI21_X1 U17076 ( .B1(P2_EBX_REG_7__SCAN_IN), .B2(n19065), .A(n13687), .ZN(
        n13688) );
  OAI21_X1 U17077 ( .B1(n15476), .B2(n19047), .A(n13688), .ZN(n13689) );
  AOI211_X1 U17078 ( .C1(n13691), .C2(n19036), .A(n13690), .B(n13689), .ZN(
        n13692) );
  INV_X1 U17079 ( .A(n13692), .ZN(P2_U2848) );
  INV_X1 U17080 ( .A(n13693), .ZN(n13698) );
  OAI22_X1 U17081 ( .A1(n19014), .A2(n13694), .B1(n19763), .B2(n19061), .ZN(
        n13697) );
  NOR2_X1 U17082 ( .A1(n19072), .A2(n13695), .ZN(n13696) );
  AOI211_X1 U17083 ( .C1(n19041), .C2(n13698), .A(n13697), .B(n13696), .ZN(
        n13700) );
  NAND2_X1 U17084 ( .A1(n19852), .A2(n19042), .ZN(n13699) );
  OAI211_X1 U17085 ( .C1(n15508), .C2(n19047), .A(n13700), .B(n13699), .ZN(
        n13704) );
  OAI21_X1 U17086 ( .B1(n19078), .B2(n13702), .A(n13701), .ZN(n15509) );
  OAI22_X1 U17087 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19071), .B1(
        n15509), .B2(n19741), .ZN(n13703) );
  AOI211_X1 U17088 ( .C1(n19074), .C2(n19848), .A(n13704), .B(n13703), .ZN(
        n13705) );
  INV_X1 U17089 ( .A(n13705), .ZN(P2_U2854) );
  INV_X1 U17090 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13707) );
  OAI222_X1 U17091 ( .A1(n15950), .A2(n20001), .B1(n20012), .B2(n13707), .C1(
        n14561), .C2(n13706), .ZN(P1_U2864) );
  INV_X1 U17092 ( .A(n13708), .ZN(n13710) );
  INV_X1 U17093 ( .A(n16138), .ZN(n13711) );
  NOR2_X1 U17094 ( .A1(n19052), .A2(n13709), .ZN(n18948) );
  OAI211_X1 U17095 ( .C1(n13710), .C2(n13711), .A(n19036), .B(n18948), .ZN(
        n13717) );
  OAI22_X1 U17096 ( .A1(n16140), .A2(n19047), .B1(n13711), .B2(n19071), .ZN(
        n13714) );
  INV_X1 U17097 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19779) );
  AOI22_X1 U17098 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19043), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19065), .ZN(n13712) );
  OAI211_X1 U17099 ( .C1(n19779), .C2(n19061), .A(n13712), .B(n19045), .ZN(
        n13713) );
  AOI211_X1 U17100 ( .C1(n19041), .C2(n13715), .A(n13714), .B(n13713), .ZN(
        n13716) );
  OAI211_X1 U17101 ( .C1(n13718), .C2(n19063), .A(n13717), .B(n13716), .ZN(
        P2_U2842) );
  AND2_X1 U17102 ( .A1(n13607), .A2(n13719), .ZN(n13720) );
  NOR2_X1 U17103 ( .A1(n13721), .A2(n13720), .ZN(n20003) );
  INV_X1 U17104 ( .A(n20003), .ZN(n13725) );
  INV_X1 U17105 ( .A(DATAI_9_), .ZN(n13723) );
  NAND2_X1 U17106 ( .A1(n20143), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13722) );
  OAI21_X1 U17107 ( .B1(n20143), .B2(n13723), .A(n13722), .ZN(n20053) );
  AOI22_X1 U17108 ( .A1(n15770), .A2(n20053), .B1(n15768), .B2(
        P1_EAX_REG_9__SCAN_IN), .ZN(n13724) );
  OAI21_X1 U17109 ( .B1(n13725), .B2(n20016), .A(n13724), .ZN(P1_U2895) );
  INV_X1 U17110 ( .A(n13726), .ZN(n14753) );
  AND2_X1 U17111 ( .A1(n15937), .A2(n13727), .ZN(n13728) );
  OR2_X1 U17112 ( .A1(n13728), .A2(n15758), .ZN(n15927) );
  OAI22_X1 U17113 ( .A1(n20001), .A2(n15927), .B1(n13729), .B2(n20012), .ZN(
        n13730) );
  AOI21_X1 U17114 ( .B1(n14753), .B2(n20008), .A(n13730), .ZN(n13731) );
  INV_X1 U17115 ( .A(n13731), .ZN(P1_U2862) );
  XNOR2_X1 U17116 ( .A(n13746), .B(n13805), .ZN(n13735) );
  MUX2_X1 U17117 ( .A(n13733), .B(n13732), .S(n14992), .Z(n13734) );
  OAI21_X1 U17118 ( .B1(n13735), .B2(n15026), .A(n13734), .ZN(P2_U2872) );
  XNOR2_X1 U17119 ( .A(n13737), .B(n13736), .ZN(n13738) );
  XNOR2_X1 U17120 ( .A(n13739), .B(n13738), .ZN(n15954) );
  INV_X1 U17121 ( .A(n15954), .ZN(n13745) );
  AOI22_X1 U17122 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13740) );
  OAI21_X1 U17123 ( .B1(n20085), .B2(n13741), .A(n13740), .ZN(n13742) );
  AOI21_X1 U17124 ( .B1(n13743), .B2(n14666), .A(n13742), .ZN(n13744) );
  OAI21_X1 U17125 ( .B1(n13745), .B2(n19900), .A(n13744), .ZN(P1_U2991) );
  OR2_X1 U17126 ( .A1(n13746), .A2(n13805), .ZN(n13761) );
  AOI22_X1 U17127 ( .A1(n14096), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14136), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13754) );
  NAND2_X1 U17128 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13748) );
  NAND2_X1 U17129 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13747) );
  OAI211_X1 U17130 ( .C1(n14099), .C2(n13749), .A(n13748), .B(n13747), .ZN(
        n13750) );
  INV_X1 U17131 ( .A(n13750), .ZN(n13753) );
  AOI22_X1 U17132 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13752) );
  AOI22_X1 U17133 ( .A1(n14143), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13751) );
  NAND4_X1 U17134 ( .A1(n13754), .A2(n13753), .A3(n13752), .A4(n13751), .ZN(
        n13760) );
  AOI22_X1 U17135 ( .A1(n14150), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14077), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13758) );
  AOI22_X1 U17136 ( .A1(n10970), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13757) );
  AOI22_X1 U17137 ( .A1(n14154), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13756) );
  NAND2_X1 U17138 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13755) );
  NAND4_X1 U17139 ( .A1(n13758), .A2(n13757), .A3(n13756), .A4(n13755), .ZN(
        n13759) );
  NOR2_X1 U17140 ( .A1(n13760), .A2(n13759), .ZN(n13803) );
  NAND2_X1 U17141 ( .A1(n13761), .A2(n13803), .ZN(n13762) );
  NAND2_X1 U17142 ( .A1(n13802), .A2(n13762), .ZN(n19085) );
  OAI21_X1 U17143 ( .B1(n13764), .B2(n13763), .A(n15037), .ZN(n18942) );
  MUX2_X1 U17144 ( .A(n18942), .B(n11069), .S(n15040), .Z(n13765) );
  OAI21_X1 U17145 ( .B1(n19085), .B2(n15026), .A(n13765), .ZN(P2_U2871) );
  XNOR2_X1 U17146 ( .A(n9738), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13767) );
  XNOR2_X1 U17147 ( .A(n13766), .B(n13767), .ZN(n15932) );
  AOI22_X1 U17148 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n13768) );
  OAI21_X1 U17149 ( .B1(n20085), .B2(n13769), .A(n13768), .ZN(n13770) );
  AOI21_X1 U17150 ( .B1(n20003), .B2(n14666), .A(n13770), .ZN(n13771) );
  OAI21_X1 U17151 ( .B1(n15932), .B2(n19900), .A(n13771), .ZN(P1_U2990) );
  XOR2_X1 U17152 ( .A(n13773), .B(n13772), .Z(n16199) );
  INV_X1 U17153 ( .A(n16199), .ZN(n13788) );
  NAND2_X1 U17154 ( .A1(n13775), .A2(n13774), .ZN(n13777) );
  XNOR2_X1 U17155 ( .A(n13777), .B(n13776), .ZN(n16201) );
  OR2_X1 U17156 ( .A1(n16297), .A2(n16298), .ZN(n19201) );
  AOI221_X1 U17157 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n19190), .C2(n13781), .A(
        n19201), .ZN(n13786) );
  OAI21_X1 U17158 ( .B1(n13566), .B2(n13779), .A(n13778), .ZN(n19112) );
  INV_X1 U17159 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13782) );
  OAI21_X1 U17160 ( .B1(n16297), .B2(n13780), .A(n16207), .ZN(n19189) );
  OAI22_X1 U17161 ( .A1(n19045), .A2(n13782), .B1(n19189), .B2(n13781), .ZN(
        n13783) );
  AOI21_X1 U17162 ( .B1(n19192), .B2(n19035), .A(n13783), .ZN(n13784) );
  OAI21_X1 U17163 ( .B1(n19112), .B2(n16289), .A(n13784), .ZN(n13785) );
  AOI211_X1 U17164 ( .C1(n16201), .C2(n16281), .A(n13786), .B(n13785), .ZN(
        n13787) );
  OAI21_X1 U17165 ( .B1(n13788), .B2(n16305), .A(n13787), .ZN(P2_U3041) );
  AOI22_X1 U17166 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n14096), .B1(
        n14136), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13795) );
  NAND2_X1 U17167 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13790) );
  NAND2_X1 U17168 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13789) );
  OAI211_X1 U17169 ( .C1(n14099), .C2(n14175), .A(n13790), .B(n13789), .ZN(
        n13791) );
  INV_X1 U17170 ( .A(n13791), .ZN(n13794) );
  AOI22_X1 U17171 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13793) );
  AOI22_X1 U17172 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n14143), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13792) );
  NAND4_X1 U17173 ( .A1(n13795), .A2(n13794), .A3(n13793), .A4(n13792), .ZN(
        n13801) );
  AOI22_X1 U17174 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n14077), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13799) );
  AOI22_X1 U17175 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10970), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13798) );
  AOI22_X1 U17176 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13797) );
  NAND2_X1 U17177 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13796) );
  NAND4_X1 U17178 ( .A1(n13799), .A2(n13798), .A3(n13797), .A4(n13796), .ZN(
        n13800) );
  NOR2_X1 U17179 ( .A1(n13801), .A2(n13800), .ZN(n13804) );
  AND2_X1 U17180 ( .A1(n13802), .A2(n13804), .ZN(n13807) );
  OR2_X1 U17181 ( .A1(n13804), .A2(n13803), .ZN(n13806) );
  NOR2_X1 U17182 ( .A1(n13806), .A2(n13805), .ZN(n13835) );
  AND2_X1 U17183 ( .A1(n9838), .A2(n13835), .ZN(n15029) );
  OR2_X1 U17184 ( .A1(n14018), .A2(n13808), .ZN(n13809) );
  AND2_X1 U17185 ( .A1(n15389), .A2(n13809), .ZN(n18930) );
  AND2_X1 U17186 ( .A1(n19103), .A2(n13810), .ZN(n13813) );
  NAND2_X1 U17187 ( .A1(n19084), .A2(BUF2_REG_17__SCAN_IN), .ZN(n13819) );
  NAND2_X1 U17188 ( .A1(n19083), .A2(BUF1_REG_17__SCAN_IN), .ZN(n13818) );
  AND2_X1 U17189 ( .A1(n13814), .A2(n9755), .ZN(n13815) );
  AOI22_X1 U17190 ( .A1(n19082), .A2(n13816), .B1(n19104), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n13817) );
  NAND3_X1 U17191 ( .A1(n13819), .A2(n13818), .A3(n13817), .ZN(n13820) );
  AOI21_X1 U17192 ( .B1(n18930), .B2(n19087), .A(n13820), .ZN(n13821) );
  OAI21_X1 U17193 ( .B1(n19107), .B2(n15043), .A(n13821), .ZN(P2_U2902) );
  AOI22_X1 U17194 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n14096), .B1(
        n14136), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13828) );
  INV_X1 U17195 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14199) );
  NAND2_X1 U17196 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13823) );
  NAND2_X1 U17197 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n13822) );
  OAI211_X1 U17198 ( .C1(n14099), .C2(n14199), .A(n13823), .B(n13822), .ZN(
        n13824) );
  INV_X1 U17199 ( .A(n13824), .ZN(n13827) );
  AOI22_X1 U17200 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13826) );
  AOI22_X1 U17201 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n14143), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13825) );
  NAND4_X1 U17202 ( .A1(n13828), .A2(n13827), .A3(n13826), .A4(n13825), .ZN(
        n13834) );
  AOI22_X1 U17203 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n14077), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13832) );
  AOI22_X1 U17204 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10970), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13831) );
  AOI22_X1 U17205 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13830) );
  NAND2_X1 U17206 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13829) );
  NAND4_X1 U17207 ( .A1(n13832), .A2(n13831), .A3(n13830), .A4(n13829), .ZN(
        n13833) );
  OR2_X1 U17208 ( .A1(n13834), .A2(n13833), .ZN(n15028) );
  AND2_X1 U17209 ( .A1(n15028), .A2(n13835), .ZN(n13849) );
  NAND2_X1 U17210 ( .A1(n13849), .A2(n9838), .ZN(n15031) );
  INV_X1 U17211 ( .A(n15031), .ZN(n13852) );
  AOI22_X1 U17212 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14096), .B1(
        n14136), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13842) );
  INV_X1 U17213 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14222) );
  NAND2_X1 U17214 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n13837) );
  NAND2_X1 U17215 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n13836) );
  OAI211_X1 U17216 ( .C1(n14099), .C2(n14222), .A(n13837), .B(n13836), .ZN(
        n13838) );
  INV_X1 U17217 ( .A(n13838), .ZN(n13841) );
  AOI22_X1 U17218 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13840) );
  AOI22_X1 U17219 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n14143), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13839) );
  NAND4_X1 U17220 ( .A1(n13842), .A2(n13841), .A3(n13840), .A4(n13839), .ZN(
        n13848) );
  AOI22_X1 U17221 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n14077), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U17222 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n14152), .B1(
        n10970), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13845) );
  AOI22_X1 U17223 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13844) );
  NAND2_X1 U17224 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13843) );
  NAND4_X1 U17225 ( .A1(n13846), .A2(n13845), .A3(n13844), .A4(n13843), .ZN(
        n13847) );
  OR2_X1 U17226 ( .A1(n13848), .A2(n13847), .ZN(n13851) );
  OAI21_X1 U17227 ( .B1(n13852), .B2(n13851), .A(n15016), .ZN(n15027) );
  XNOR2_X1 U17228 ( .A(n15391), .B(n13853), .ZN(n18905) );
  NAND2_X1 U17229 ( .A1(n19084), .A2(BUF2_REG_19__SCAN_IN), .ZN(n13857) );
  NAND2_X1 U17230 ( .A1(n19083), .A2(BUF1_REG_19__SCAN_IN), .ZN(n13856) );
  AOI22_X1 U17231 ( .A1(n19082), .A2(n13854), .B1(n19104), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n13855) );
  NAND3_X1 U17232 ( .A1(n13857), .A2(n13856), .A3(n13855), .ZN(n13858) );
  AOI21_X1 U17233 ( .B1(n18905), .B2(n19087), .A(n13858), .ZN(n13859) );
  OAI21_X1 U17234 ( .B1(n19107), .B2(n15027), .A(n13859), .ZN(P2_U2900) );
  NAND2_X1 U17235 ( .A1(n13644), .A2(n13860), .ZN(n13861) );
  NAND2_X1 U17236 ( .A1(n13862), .A2(n13861), .ZN(n15752) );
  OAI21_X1 U17237 ( .B1(n15752), .B2(n15753), .A(n13862), .ZN(n13890) );
  AOI22_X1 U17238 ( .A1(n15770), .A2(n14567), .B1(n15768), .B2(
        P1_EAX_REG_13__SCAN_IN), .ZN(n13864) );
  OAI21_X1 U17239 ( .B1(n14743), .B2(n20016), .A(n13864), .ZN(P1_U2891) );
  INV_X1 U17240 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20744) );
  INV_X1 U17241 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20741) );
  NAND3_X1 U17242 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(n13865), .ZN(n13868) );
  NOR2_X1 U17243 ( .A1(n13866), .A2(n13868), .ZN(n15755) );
  NAND3_X1 U17244 ( .A1(n19985), .A2(n15755), .A3(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n15747) );
  NOR2_X1 U17245 ( .A1(n20741), .A2(n15747), .ZN(n15729) );
  INV_X1 U17246 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14738) );
  INV_X1 U17247 ( .A(n19954), .ZN(n19964) );
  AOI21_X1 U17248 ( .B1(n14740), .B2(n19982), .A(n19964), .ZN(n13867) );
  OAI21_X1 U17249 ( .B1(n14738), .B2(n19993), .A(n13867), .ZN(n13878) );
  NAND2_X1 U17250 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n13873) );
  INV_X1 U17251 ( .A(n13868), .ZN(n13872) );
  INV_X1 U17252 ( .A(n13869), .ZN(n13870) );
  AND2_X1 U17253 ( .A1(n19989), .A2(n13870), .ZN(n19970) );
  INV_X1 U17254 ( .A(n19970), .ZN(n13871) );
  OAI21_X1 U17255 ( .B1(n15647), .B2(n13872), .A(n13871), .ZN(n15761) );
  AOI21_X1 U17256 ( .B1(n13873), .B2(n19989), .A(n15761), .ZN(n15746) );
  INV_X1 U17257 ( .A(n13895), .ZN(n13874) );
  AOI21_X1 U17258 ( .B1(n13875), .B2(n13888), .A(n13874), .ZN(n15895) );
  AOI22_X1 U17259 ( .A1(n19991), .A2(n15895), .B1(n19994), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n13876) );
  OAI21_X1 U17260 ( .B1(n15746), .B2(n20744), .A(n13876), .ZN(n13877) );
  AOI211_X1 U17261 ( .C1(n20744), .C2(n15729), .A(n13878), .B(n13877), .ZN(
        n13879) );
  OAI21_X1 U17262 ( .B1(n14743), .B2(n15751), .A(n13879), .ZN(P1_U2827) );
  AOI22_X1 U17263 ( .A1(n15895), .A2(n20007), .B1(n14520), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n13880) );
  OAI21_X1 U17264 ( .B1(n14743), .B2(n14561), .A(n13880), .ZN(P1_U2859) );
  AOI21_X1 U17265 ( .B1(n10124), .B2(n9780), .A(n12240), .ZN(n15736) );
  INV_X1 U17266 ( .A(n15736), .ZN(n13897) );
  INV_X1 U17267 ( .A(DATAI_14_), .ZN(n13884) );
  NAND2_X1 U17268 ( .A1(n20143), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13883) );
  OAI21_X1 U17269 ( .B1(n20143), .B2(n13884), .A(n13883), .ZN(n20059) );
  AOI22_X1 U17270 ( .A1(n15770), .A2(n20059), .B1(n15768), .B2(
        P1_EAX_REG_14__SCAN_IN), .ZN(n13885) );
  OAI21_X1 U17271 ( .B1(n13897), .B2(n20016), .A(n13885), .ZN(P1_U2890) );
  OR2_X1 U17272 ( .A1(n15760), .A2(n13886), .ZN(n13887) );
  NAND2_X1 U17273 ( .A1(n13888), .A2(n13887), .ZN(n15908) );
  INV_X1 U17274 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n13893) );
  NOR2_X1 U17275 ( .A1(n13890), .A2(n13889), .ZN(n13891) );
  OAI222_X1 U17276 ( .A1(n15908), .A2(n20001), .B1(n20012), .B2(n13893), .C1(
        n14561), .C2(n15817), .ZN(P1_U2860) );
  AND2_X1 U17277 ( .A1(n13895), .A2(n13894), .ZN(n13896) );
  OR2_X1 U17278 ( .A1(n13896), .A2(n9839), .ZN(n15731) );
  INV_X1 U17279 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n13898) );
  OAI222_X1 U17280 ( .A1(n15731), .A2(n20001), .B1(n20012), .B2(n13898), .C1(
        n14561), .C2(n13897), .ZN(P1_U2858) );
  INV_X1 U17281 ( .A(n14451), .ZN(n13899) );
  AOI21_X1 U17282 ( .B1(n13900), .B2(n13882), .A(n13899), .ZN(n15810) );
  INV_X1 U17283 ( .A(n15810), .ZN(n14562) );
  OAI222_X1 U17284 ( .A1(n14562), .A2(n20016), .B1(n20014), .B2(n13901), .C1(
        n20015), .C2(n20022), .ZN(P1_U2889) );
  OAI211_X1 U17285 ( .C1(n18819), .C2(n18666), .A(n10298), .B(n18655), .ZN(
        n18190) );
  NOR2_X1 U17286 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18190), .ZN(n13902) );
  NAND3_X1 U17287 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18808)
         );
  OAI21_X1 U17288 ( .B1(n13902), .B2(n18808), .A(n18472), .ZN(n18196) );
  INV_X1 U17289 ( .A(n18196), .ZN(n13903) );
  INV_X1 U17290 ( .A(n17822), .ZN(n17687) );
  NOR2_X1 U17291 ( .A1(n17687), .A2(n18861), .ZN(n15531) );
  AOI21_X1 U17292 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15531), .ZN(n15532) );
  NOR2_X1 U17293 ( .A1(n13903), .A2(n15532), .ZN(n13905) );
  OAI21_X1 U17294 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n18810), .A(
        n18196), .ZN(n15530) );
  OR2_X1 U17295 ( .A1(n18496), .A2(n15530), .ZN(n13904) );
  MUX2_X1 U17296 ( .A(n13905), .B(n13904), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AND2_X1 U17297 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16930) );
  NAND2_X1 U17298 ( .A1(n18240), .A2(n17230), .ZN(n17224) );
  INV_X2 U17299 ( .A(n17227), .ZN(n17222) );
  INV_X1 U17300 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16888) );
  INV_X1 U17301 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16940) );
  INV_X1 U17302 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n13911) );
  INV_X1 U17303 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16995) );
  INV_X1 U17304 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16661) );
  INV_X1 U17305 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16681) );
  INV_X1 U17306 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n21047) );
  INV_X1 U17307 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17083) );
  INV_X1 U17308 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16822) );
  INV_X1 U17309 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16847) );
  NAND3_X1 U17310 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17215) );
  NOR2_X1 U17311 ( .A1(n16847), .A2(n17215), .ZN(n17205) );
  AND2_X1 U17312 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_9__SCAN_IN), 
        .ZN(n17116) );
  NAND4_X1 U17313 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(P3_EBX_REG_7__SCAN_IN), .A4(n17116), .ZN(n17081) );
  NAND2_X1 U17314 ( .A1(n18240), .A2(n17010), .ZN(n16994) );
  NAND2_X1 U17315 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n9828), .ZN(n16936) );
  NAND2_X1 U17316 ( .A1(n17222), .A2(n16936), .ZN(n16934) );
  OAI21_X1 U17317 ( .B1(n16930), .B2(n17224), .A(n16934), .ZN(n16928) );
  OAI22_X1 U17318 ( .A1(n10298), .A2(n17117), .B1(n17170), .B2(n18222), .ZN(
        n13921) );
  AOI22_X1 U17319 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10309), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13919) );
  AOI22_X1 U17320 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13918) );
  INV_X1 U17321 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18276) );
  AOI22_X1 U17322 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13912) );
  OAI21_X1 U17323 ( .B1(n17188), .B2(n18276), .A(n13912), .ZN(n13916) );
  AOI22_X1 U17324 ( .A1(n17104), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13914) );
  AOI22_X1 U17325 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13913) );
  OAI211_X1 U17326 ( .C1(n17143), .C2(n17119), .A(n13914), .B(n13913), .ZN(
        n13915) );
  AOI211_X1 U17327 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n13916), .B(n13915), .ZN(n13917) );
  NAND3_X1 U17328 ( .A1(n13919), .A2(n13918), .A3(n13917), .ZN(n13920) );
  AOI211_X1 U17329 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n13921), .B(n13920), .ZN(n16937) );
  AOI22_X1 U17330 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13922) );
  OAI21_X1 U17331 ( .B1(n20831), .B2(n17170), .A(n13922), .ZN(n13931) );
  AOI22_X1 U17332 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17182), .ZN(n13929) );
  AOI22_X1 U17333 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17139), .ZN(n13923) );
  OAI21_X1 U17334 ( .B1(n17025), .B2(n10268), .A(n13923), .ZN(n13927) );
  AOI22_X1 U17335 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n17177), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13925) );
  AOI22_X1 U17336 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17104), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13924) );
  OAI211_X1 U17337 ( .C1(n17161), .C2(n17143), .A(n13925), .B(n13924), .ZN(
        n13926) );
  AOI211_X1 U17338 ( .C1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(n17038), .A(
        n13927), .B(n13926), .ZN(n13928) );
  OAI211_X1 U17339 ( .C1(n20881), .C2(n10221), .A(n13929), .B(n13928), .ZN(
        n13930) );
  AOI211_X1 U17340 ( .C1(n17159), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n13931), .B(n13930), .ZN(n16946) );
  AOI22_X1 U17341 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13941) );
  AOI22_X1 U17342 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13933) );
  AOI22_X1 U17343 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10309), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13932) );
  OAI211_X1 U17344 ( .C1(n17188), .C2(n18268), .A(n13933), .B(n13932), .ZN(
        n13939) );
  AOI22_X1 U17345 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13937) );
  AOI22_X1 U17346 ( .A1(n9733), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13936) );
  AOI22_X1 U17347 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13935) );
  NAND2_X1 U17348 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13934) );
  NAND4_X1 U17349 ( .A1(n13937), .A2(n13936), .A3(n13935), .A4(n13934), .ZN(
        n13938) );
  AOI211_X1 U17350 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n13939), .B(n13938), .ZN(n13940) );
  OAI211_X1 U17351 ( .C1(n10275), .C2(n17179), .A(n13941), .B(n13940), .ZN(
        n16950) );
  AOI22_X1 U17352 ( .A1(n9733), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13952) );
  AOI22_X1 U17353 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13942) );
  OAI21_X1 U17354 ( .B1(n10234), .B2(n18469), .A(n13942), .ZN(n13950) );
  AOI22_X1 U17355 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13948) );
  AOI22_X1 U17356 ( .A1(n17177), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13944) );
  AOI22_X1 U17357 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13943) );
  OAI211_X1 U17358 ( .C1(n10268), .C2(n13945), .A(n13944), .B(n13943), .ZN(
        n13946) );
  AOI21_X1 U17359 ( .B1(n17038), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n13946), .ZN(n13947) );
  OAI211_X1 U17360 ( .C1(n17143), .C2(n17062), .A(n13948), .B(n13947), .ZN(
        n13949) );
  AOI211_X1 U17361 ( .C1(n17173), .C2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n13950), .B(n13949), .ZN(n13951) );
  OAI211_X1 U17362 ( .C1(n10298), .C2(n21001), .A(n13952), .B(n13951), .ZN(
        n16951) );
  NAND2_X1 U17363 ( .A1(n16950), .A2(n16951), .ZN(n16949) );
  NOR2_X1 U17364 ( .A1(n16946), .A2(n16949), .ZN(n16943) );
  AOI22_X1 U17365 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17038), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13962) );
  AOI22_X1 U17366 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U17367 ( .A1(n9733), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17104), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13953) );
  OAI211_X1 U17368 ( .C1(n17143), .C2(n20961), .A(n13954), .B(n13953), .ZN(
        n13960) );
  AOI22_X1 U17369 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13958) );
  AOI22_X1 U17370 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10309), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13957) );
  AOI22_X1 U17371 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13956) );
  NAND2_X1 U17372 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13955) );
  NAND4_X1 U17373 ( .A1(n13958), .A2(n13957), .A3(n13956), .A4(n13955), .ZN(
        n13959) );
  AOI211_X1 U17374 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n13960), .B(n13959), .ZN(n13961) );
  OAI211_X1 U17375 ( .C1(n10275), .C2(n17137), .A(n13962), .B(n13961), .ZN(
        n16942) );
  NAND2_X1 U17376 ( .A1(n16943), .A2(n16942), .ZN(n16941) );
  NOR2_X1 U17377 ( .A1(n16937), .A2(n16941), .ZN(n17256) );
  INV_X1 U17378 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17103) );
  AOI22_X1 U17379 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13972) );
  AOI22_X1 U17380 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13964) );
  AOI22_X1 U17381 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10309), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13963) );
  OAI211_X1 U17382 ( .C1(n10268), .C2(n20909), .A(n13964), .B(n13963), .ZN(
        n13970) );
  AOI22_X1 U17383 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9733), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13968) );
  AOI22_X1 U17384 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13967) );
  AOI22_X1 U17385 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13966) );
  NAND2_X1 U17386 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13965) );
  NAND4_X1 U17387 ( .A1(n13968), .A2(n13967), .A3(n13966), .A4(n13965), .ZN(
        n13969) );
  AOI211_X1 U17388 ( .C1(n17038), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n13970), .B(n13969), .ZN(n13971) );
  OAI211_X1 U17389 ( .C1(n10234), .C2(n17103), .A(n13972), .B(n13971), .ZN(
        n17255) );
  NAND2_X1 U17390 ( .A1(n17256), .A2(n17255), .ZN(n17254) );
  AOI22_X1 U17391 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13982) );
  INV_X1 U17392 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n21035) );
  AOI22_X1 U17393 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13973) );
  OAI21_X1 U17394 ( .B1(n9800), .B2(n21035), .A(n13973), .ZN(n13980) );
  AOI22_X1 U17395 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13978) );
  AOI22_X1 U17396 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10309), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13975) );
  AOI22_X1 U17397 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9733), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13974) );
  OAI211_X1 U17398 ( .C1(n17188), .C2(n18281), .A(n13975), .B(n13974), .ZN(
        n13976) );
  AOI21_X1 U17399 ( .B1(n17183), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n13976), .ZN(n13977) );
  OAI211_X1 U17400 ( .C1(n17143), .C2(n17087), .A(n13978), .B(n13977), .ZN(
        n13979) );
  AOI211_X1 U17401 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n13980), .B(n13979), .ZN(n13981) );
  OAI211_X1 U17402 ( .C1(n10221), .C2(n16969), .A(n13982), .B(n13981), .ZN(
        n16925) );
  XNOR2_X1 U17403 ( .A(n17254), .B(n16925), .ZN(n17249) );
  AOI22_X1 U17404 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16928), .B1(n17227), 
        .B2(n17249), .ZN(n13985) );
  INV_X1 U17405 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n13983) );
  INV_X1 U17406 ( .A(n16936), .ZN(n16939) );
  NAND3_X1 U17407 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n13983), .A3(n16939), 
        .ZN(n13984) );
  NAND2_X1 U17408 ( .A1(n13985), .A2(n13984), .ZN(P3_U2675) );
  INV_X1 U17409 ( .A(n13986), .ZN(n16300) );
  AOI22_X1 U17410 ( .A1(n16300), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n19186), .B2(n19843), .ZN(n14000) );
  XOR2_X1 U17411 ( .A(n13988), .B(n13987), .Z(n14005) );
  INV_X1 U17412 ( .A(n14013), .ZN(n13991) );
  NAND2_X1 U17413 ( .A1(n13990), .A2(n13989), .ZN(n13993) );
  AOI22_X1 U17414 ( .A1(n16281), .A2(n14005), .B1(n13991), .B2(n13993), .ZN(
        n13999) );
  INV_X1 U17415 ( .A(n13992), .ZN(n14014) );
  INV_X1 U17416 ( .A(n13993), .ZN(n13994) );
  AND2_X1 U17417 ( .A1(n19029), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14004) );
  AOI21_X1 U17418 ( .B1(n14014), .B2(n13994), .A(n14004), .ZN(n13998) );
  NAND2_X1 U17419 ( .A1(n13996), .A2(n13995), .ZN(n14002) );
  NAND3_X1 U17420 ( .A1(n14003), .A2(n19187), .A3(n14002), .ZN(n13997) );
  AND4_X1 U17421 ( .A1(n14000), .A2(n13999), .A3(n13998), .A4(n13997), .ZN(
        n14001) );
  OAI21_X1 U17422 ( .B1(n13678), .B2(n16266), .A(n14001), .ZN(P2_U3044) );
  NAND3_X1 U17423 ( .A1(n14003), .A2(n19175), .A3(n14002), .ZN(n14010) );
  AOI21_X1 U17424 ( .B1(n16200), .B2(n14005), .A(n14004), .ZN(n14009) );
  NAND2_X1 U17425 ( .A1(n19169), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14008) );
  NAND2_X1 U17426 ( .A1(n16198), .A2(n14006), .ZN(n14007) );
  AND4_X1 U17427 ( .A1(n14010), .A2(n14009), .A3(n14008), .A4(n14007), .ZN(
        n14011) );
  OAI21_X1 U17428 ( .B1(n13678), .B2(n16158), .A(n14011), .ZN(P2_U3012) );
  OR2_X1 U17429 ( .A1(n16309), .A2(n14019), .ZN(n14012) );
  NAND2_X1 U17430 ( .A1(n15465), .A2(n14012), .ZN(n16240) );
  INV_X1 U17431 ( .A(n15422), .ZN(n16261) );
  NOR2_X2 U17432 ( .A1(n16154), .A2(n16261), .ZN(n16156) );
  NAND2_X1 U17433 ( .A1(n16156), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15436) );
  OR2_X2 U17434 ( .A1(n15436), .A2(n15426), .ZN(n16129) );
  AND2_X1 U17435 ( .A1(n14016), .A2(n14015), .ZN(n14017) );
  NOR2_X1 U17436 ( .A1(n14018), .A2(n14017), .ZN(n19088) );
  OAI22_X1 U17437 ( .A1(n16266), .A2(n18942), .B1(n19785), .B2(n19045), .ZN(
        n14022) );
  INV_X1 U17438 ( .A(n15471), .ZN(n16249) );
  INV_X1 U17439 ( .A(n14019), .ZN(n14020) );
  NOR2_X1 U17440 ( .A1(n16249), .A2(n14020), .ZN(n16235) );
  AOI21_X1 U17441 ( .B1(n10168), .B2(n16281), .A(n16235), .ZN(n15404) );
  NOR3_X1 U17442 ( .A1(n15404), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15237), .ZN(n14021) );
  AOI211_X1 U17443 ( .C1(n19186), .C2(n19088), .A(n14022), .B(n14021), .ZN(
        n14028) );
  INV_X1 U17444 ( .A(n15417), .ZN(n15433) );
  NAND2_X1 U17445 ( .A1(n16161), .A2(n16159), .ZN(n15413) );
  NAND2_X1 U17446 ( .A1(n15418), .A2(n15416), .ZN(n14023) );
  NOR2_X1 U17447 ( .A1(n15413), .A2(n14023), .ZN(n14024) );
  INV_X1 U17448 ( .A(n14025), .ZN(n14026) );
  XNOR2_X1 U17449 ( .A(n15174), .B(n15171), .ZN(n15231) );
  NAND2_X1 U17450 ( .A1(n15231), .A2(n19187), .ZN(n14027) );
  OAI211_X1 U17451 ( .C1(n15402), .C2(n15236), .A(n14028), .B(n14027), .ZN(
        P2_U3030) );
  NOR2_X1 U17452 ( .A1(n14879), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14029) );
  AOI21_X1 U17453 ( .B1(n20256), .B2(n14882), .A(n14029), .ZN(n15573) );
  INV_X1 U17454 ( .A(n14032), .ZN(n14893) );
  AOI22_X1 U17455 ( .A1(n14035), .A2(n15602), .B1(n20110), .B2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n14030) );
  OAI21_X1 U17456 ( .B1(n15573), .B2(n14893), .A(n14030), .ZN(n14033) );
  AND2_X1 U17457 ( .A1(n14031), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15571) );
  AOI22_X1 U17458 ( .A1(n14894), .A2(n14033), .B1(n14032), .B2(n15571), .ZN(
        n14034) );
  OAI21_X1 U17459 ( .B1(n14035), .B2(n14894), .A(n14034), .ZN(P1_U3474) );
  XNOR2_X1 U17460 ( .A(n13372), .B(n20650), .ZN(n14037) );
  OAI222_X1 U17461 ( .A1(n14038), .A2(n14037), .B1(n14036), .B2(n12539), .C1(
        n20520), .C2(n14063), .ZN(P1_U3476) );
  XNOR2_X1 U17462 ( .A(n15136), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15294) );
  NAND3_X1 U17463 ( .A1(n9755), .A2(P2_EBX_REG_27__SCAN_IN), .A3(n14041), .ZN(
        n14043) );
  NAND2_X1 U17464 ( .A1(n14044), .A2(n14043), .ZN(n16032) );
  NOR2_X1 U17465 ( .A1(n16032), .A2(n14045), .ZN(n14047) );
  XNOR2_X1 U17466 ( .A(n14048), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14049) );
  NAND2_X1 U17467 ( .A1(n15285), .A2(n19175), .ZN(n14058) );
  OR2_X1 U17468 ( .A1(n14051), .A2(n14050), .ZN(n14052) );
  NAND2_X1 U17469 ( .A1(n14948), .A2(n14052), .ZN(n15288) );
  INV_X1 U17470 ( .A(n15288), .ZN(n16021) );
  NAND2_X1 U17471 ( .A1(n19029), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n15287) );
  OAI21_X1 U17472 ( .B1(n16204), .B2(n14053), .A(n15287), .ZN(n14056) );
  NAND2_X1 U17473 ( .A1(n15131), .A2(n14053), .ZN(n14054) );
  NAND2_X1 U17474 ( .A1(n15122), .A2(n14054), .ZN(n16024) );
  NOR2_X1 U17475 ( .A1(n16024), .A2(n19167), .ZN(n14055) );
  AOI211_X1 U17476 ( .C1(n16021), .C2(n19171), .A(n14056), .B(n14055), .ZN(
        n14057) );
  OAI211_X1 U17477 ( .C1(n19177), .C2(n15294), .A(n14058), .B(n14057), .ZN(
        P2_U2986) );
  OAI211_X1 U17478 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20223), .A(n14060), 
        .B(n20650), .ZN(n14062) );
  NAND2_X1 U17479 ( .A1(n20136), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14061) );
  OAI211_X1 U17480 ( .C1(n14063), .C2(n20521), .A(n14062), .B(n14061), .ZN(
        P1_U3477) );
  AOI22_X1 U17481 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14096), .B1(
        n14136), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14070) );
  INV_X1 U17482 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14245) );
  NAND2_X1 U17483 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14065) );
  NAND2_X1 U17484 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14064) );
  OAI211_X1 U17485 ( .C1(n14099), .C2(n14245), .A(n14065), .B(n14064), .ZN(
        n14066) );
  INV_X1 U17486 ( .A(n14066), .ZN(n14069) );
  AOI22_X1 U17487 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10884), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14068) );
  AOI22_X1 U17488 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n14143), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14067) );
  NAND4_X1 U17489 ( .A1(n14070), .A2(n14069), .A3(n14068), .A4(n14067), .ZN(
        n14076) );
  AOI22_X1 U17490 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n14077), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14074) );
  AOI22_X1 U17491 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10970), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14073) );
  AOI22_X1 U17492 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14072) );
  NAND2_X1 U17493 ( .A1(n10833), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n14071) );
  NAND4_X1 U17494 ( .A1(n14074), .A2(n14073), .A3(n14072), .A4(n14071), .ZN(
        n14075) );
  NOR2_X1 U17495 ( .A1(n14076), .A2(n14075), .ZN(n15015) );
  INV_X1 U17496 ( .A(n14077), .ZN(n14109) );
  NOR2_X1 U17497 ( .A1(n14109), .A2(n14078), .ZN(n14083) );
  AOI22_X1 U17498 ( .A1(n10970), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14080) );
  AOI22_X1 U17499 ( .A1(n14154), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14079) );
  OAI211_X1 U17500 ( .C1(n14105), .C2(n14081), .A(n14080), .B(n14079), .ZN(
        n14082) );
  AOI211_X1 U17501 ( .C1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .C2(n14150), .A(
        n14083), .B(n14082), .ZN(n14095) );
  INV_X1 U17502 ( .A(n14138), .ZN(n14087) );
  INV_X1 U17503 ( .A(n14137), .ZN(n14085) );
  OAI22_X1 U17504 ( .A1(n14087), .A2(n14086), .B1(n14085), .B2(n14084), .ZN(
        n14091) );
  OAI22_X1 U17505 ( .A1(n14141), .A2(n14259), .B1(n14089), .B2(n14088), .ZN(
        n14090) );
  AOI211_X1 U17506 ( .C1(n14135), .C2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n14091), .B(n14090), .ZN(n14094) );
  AOI22_X1 U17507 ( .A1(n10884), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14144), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14093) );
  AOI22_X1 U17508 ( .A1(n14143), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14092) );
  NAND4_X1 U17509 ( .A1(n14095), .A2(n14094), .A3(n14093), .A4(n14092), .ZN(
        n15012) );
  AOI22_X1 U17510 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n14096), .B1(
        n14136), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14098) );
  AOI22_X1 U17511 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n14137), .B1(
        n14138), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14097) );
  OAI211_X1 U17512 ( .C1(n14279), .C2(n14099), .A(n14098), .B(n14097), .ZN(
        n14114) );
  AOI22_X1 U17513 ( .A1(n10884), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n14144), .ZN(n14101) );
  AOI22_X1 U17514 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n14143), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14100) );
  NAND2_X1 U17515 ( .A1(n14101), .A2(n14100), .ZN(n14113) );
  AOI22_X1 U17516 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10970), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14104) );
  AOI22_X1 U17517 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14103) );
  OAI211_X1 U17518 ( .C1(n14106), .C2(n14105), .A(n14104), .B(n14103), .ZN(
        n14112) );
  OAI22_X1 U17519 ( .A1(n14110), .A2(n14109), .B1(n14108), .B2(n14107), .ZN(
        n14111) );
  NOR4_X1 U17520 ( .A1(n14114), .A2(n14113), .A3(n14112), .A4(n14111), .ZN(
        n15006) );
  NOR2_X2 U17521 ( .A1(n15004), .A2(n15006), .ZN(n15005) );
  AOI22_X1 U17522 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14125), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14123) );
  AOI22_X1 U17523 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14166), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14122) );
  INV_X1 U17524 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14119) );
  NAND2_X1 U17525 ( .A1(n14315), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n14118) );
  INV_X1 U17526 ( .A(n14115), .ZN(n14117) );
  NAND2_X1 U17527 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14116) );
  NAND2_X1 U17528 ( .A1(n14117), .A2(n14116), .ZN(n14307) );
  OAI211_X1 U17529 ( .C1(n14165), .C2(n14119), .A(n14118), .B(n14307), .ZN(
        n14120) );
  INV_X1 U17530 ( .A(n14120), .ZN(n14121) );
  NAND4_X1 U17531 ( .A1(n14124), .A2(n14123), .A3(n14122), .A4(n14121), .ZN(
        n14134) );
  AOI22_X1 U17532 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14132) );
  AOI22_X1 U17533 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14166), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14130) );
  INV_X1 U17534 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14127) );
  NAND2_X1 U17535 ( .A1(n14303), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n14126) );
  OAI211_X1 U17536 ( .C1(n14165), .C2(n14127), .A(n14126), .B(n14277), .ZN(
        n14128) );
  INV_X1 U17537 ( .A(n14128), .ZN(n14129) );
  NAND4_X1 U17538 ( .A1(n14132), .A2(n14131), .A3(n14130), .A4(n14129), .ZN(
        n14133) );
  AND2_X1 U17539 ( .A1(n14134), .A2(n14133), .ZN(n14185) );
  NAND2_X1 U17540 ( .A1(n10757), .A2(n14185), .ZN(n14162) );
  AOI22_X1 U17541 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n14136), .B1(
        n14135), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14149) );
  INV_X1 U17542 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U17543 ( .A1(n14137), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n14140) );
  NAND2_X1 U17544 ( .A1(n14138), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n14139) );
  OAI211_X1 U17545 ( .C1(n14141), .C2(n14310), .A(n14140), .B(n14139), .ZN(
        n14142) );
  INV_X1 U17546 ( .A(n14142), .ZN(n14148) );
  AOI22_X1 U17547 ( .A1(n14144), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14143), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14147) );
  AOI22_X1 U17548 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14077), .B1(
        n14145), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14146) );
  NAND4_X1 U17549 ( .A1(n14149), .A2(n14148), .A3(n14147), .A4(n14146), .ZN(
        n14161) );
  AOI22_X1 U17550 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10884), .B1(
        n14150), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14159) );
  AOI22_X1 U17551 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10970), .B1(
        n14152), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14158) );
  AOI22_X1 U17552 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n14154), .B1(
        n14153), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14157) );
  NAND2_X1 U17553 ( .A1(n14155), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n14156) );
  NAND4_X1 U17554 ( .A1(n14159), .A2(n14158), .A3(n14157), .A4(n14156), .ZN(
        n14160) );
  OR2_X1 U17555 ( .A1(n14161), .A2(n14160), .ZN(n14164) );
  XNOR2_X1 U17556 ( .A(n14162), .B(n14164), .ZN(n14188) );
  XNOR2_X1 U17557 ( .A(n15005), .B(n14188), .ZN(n14999) );
  NAND2_X1 U17558 ( .A1(n14257), .A2(n14185), .ZN(n14998) );
  NAND2_X1 U17559 ( .A1(n14164), .A2(n14185), .ZN(n14190) );
  INV_X1 U17560 ( .A(n14274), .ZN(n14316) );
  AOI22_X1 U17561 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14173) );
  AOI22_X1 U17562 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10796), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14171) );
  INV_X1 U17563 ( .A(n14166), .ZN(n14311) );
  NAND2_X1 U17564 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n14167) );
  OAI211_X1 U17565 ( .C1(n14311), .C2(n14168), .A(n14167), .B(n14307), .ZN(
        n14169) );
  INV_X1 U17566 ( .A(n14169), .ZN(n14170) );
  NAND4_X1 U17567 ( .A1(n14173), .A2(n14172), .A3(n14171), .A4(n14170), .ZN(
        n14182) );
  AOI22_X1 U17568 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14180) );
  AOI22_X1 U17569 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10796), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14178) );
  NAND2_X1 U17570 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n14174) );
  OAI211_X1 U17571 ( .C1(n14311), .C2(n14175), .A(n14174), .B(n14277), .ZN(
        n14176) );
  INV_X1 U17572 ( .A(n14176), .ZN(n14177) );
  NAND4_X1 U17573 ( .A1(n14180), .A2(n14179), .A3(n14178), .A4(n14177), .ZN(
        n14181) );
  NAND2_X1 U17574 ( .A1(n14182), .A2(n14181), .ZN(n14189) );
  XOR2_X1 U17575 ( .A(n14190), .B(n14189), .Z(n14183) );
  NAND2_X1 U17576 ( .A1(n14183), .A2(n14207), .ZN(n14986) );
  INV_X1 U17577 ( .A(n14189), .ZN(n14184) );
  NAND2_X1 U17578 ( .A1(n14257), .A2(n14184), .ZN(n14988) );
  INV_X1 U17579 ( .A(n14185), .ZN(n14186) );
  NOR2_X1 U17580 ( .A1(n14988), .A2(n14186), .ZN(n14187) );
  NOR2_X1 U17581 ( .A1(n14190), .A2(n14189), .ZN(n14208) );
  AOI22_X1 U17582 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14197) );
  AOI22_X1 U17583 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9717), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14195) );
  INV_X1 U17584 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14192) );
  NAND2_X1 U17585 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n14191) );
  OAI211_X1 U17586 ( .C1(n14311), .C2(n14192), .A(n14191), .B(n14307), .ZN(
        n14193) );
  INV_X1 U17587 ( .A(n14193), .ZN(n14194) );
  NAND4_X1 U17588 ( .A1(n14197), .A2(n14196), .A3(n14195), .A4(n14194), .ZN(
        n14206) );
  AOI22_X1 U17589 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14204) );
  AOI22_X1 U17590 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10796), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14202) );
  NAND2_X1 U17591 ( .A1(n14303), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n14198) );
  OAI211_X1 U17592 ( .C1(n14311), .C2(n14199), .A(n14198), .B(n14277), .ZN(
        n14200) );
  INV_X1 U17593 ( .A(n14200), .ZN(n14201) );
  NAND4_X1 U17594 ( .A1(n14204), .A2(n14203), .A3(n14202), .A4(n14201), .ZN(
        n14205) );
  AND2_X1 U17595 ( .A1(n14206), .A2(n14205), .ZN(n14210) );
  NAND2_X1 U17596 ( .A1(n14208), .A2(n14210), .ZN(n14230) );
  OAI211_X1 U17597 ( .C1(n14208), .C2(n14210), .A(n14207), .B(n14230), .ZN(
        n14212) );
  INV_X1 U17598 ( .A(n14212), .ZN(n14209) );
  INV_X1 U17599 ( .A(n14210), .ZN(n14211) );
  NOR2_X1 U17600 ( .A1(n10757), .A2(n14211), .ZN(n14978) );
  NAND2_X1 U17601 ( .A1(n14979), .A2(n14978), .ZN(n14977) );
  AOI22_X1 U17602 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14220) );
  AOI22_X1 U17603 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9717), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14218) );
  NAND2_X1 U17604 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n14215) );
  OAI211_X1 U17605 ( .C1(n14311), .C2(n10773), .A(n14215), .B(n14307), .ZN(
        n14216) );
  INV_X1 U17606 ( .A(n14216), .ZN(n14217) );
  NAND4_X1 U17607 ( .A1(n14220), .A2(n14219), .A3(n14218), .A4(n14217), .ZN(
        n14229) );
  AOI22_X1 U17608 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14227) );
  AOI22_X1 U17609 ( .A1(n10038), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14315), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14226) );
  AOI22_X1 U17610 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10796), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14225) );
  NAND2_X1 U17611 ( .A1(n14125), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n14221) );
  OAI211_X1 U17612 ( .C1(n14311), .C2(n14222), .A(n14221), .B(n14277), .ZN(
        n14223) );
  INV_X1 U17613 ( .A(n14223), .ZN(n14224) );
  NAND4_X1 U17614 ( .A1(n14227), .A2(n14226), .A3(n14225), .A4(n14224), .ZN(
        n14228) );
  NAND2_X1 U17615 ( .A1(n14229), .A2(n14228), .ZN(n14232) );
  AOI21_X1 U17616 ( .B1(n14230), .B2(n14232), .A(n13071), .ZN(n14231) );
  OR2_X1 U17617 ( .A1(n14230), .A2(n14232), .ZN(n14253) );
  NAND2_X1 U17618 ( .A1(n14231), .A2(n14253), .ZN(n14234) );
  NOR2_X1 U17619 ( .A1(n10757), .A2(n14232), .ZN(n14971) );
  NAND2_X1 U17620 ( .A1(n14972), .A2(n14971), .ZN(n14970) );
  INV_X1 U17621 ( .A(n14233), .ZN(n14235) );
  AOI22_X1 U17622 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14243) );
  AOI22_X1 U17623 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9717), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14241) );
  INV_X1 U17624 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14238) );
  NAND2_X1 U17625 ( .A1(n9764), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n14237) );
  OAI211_X1 U17626 ( .C1(n14311), .C2(n14238), .A(n14237), .B(n14307), .ZN(
        n14239) );
  INV_X1 U17627 ( .A(n14239), .ZN(n14240) );
  NAND4_X1 U17628 ( .A1(n14243), .A2(n14242), .A3(n14241), .A4(n14240), .ZN(
        n14252) );
  AOI22_X1 U17629 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14250) );
  AOI22_X1 U17630 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10796), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14248) );
  NAND2_X1 U17631 ( .A1(n14303), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n14244) );
  OAI211_X1 U17632 ( .C1(n14311), .C2(n14245), .A(n14244), .B(n14277), .ZN(
        n14246) );
  INV_X1 U17633 ( .A(n14246), .ZN(n14247) );
  NAND4_X1 U17634 ( .A1(n14250), .A2(n14249), .A3(n14248), .A4(n14247), .ZN(
        n14251) );
  NAND2_X1 U17635 ( .A1(n14252), .A2(n14251), .ZN(n14255) );
  NOR2_X1 U17636 ( .A1(n14253), .A2(n14255), .ZN(n14294) );
  AOI211_X1 U17637 ( .C1(n14255), .C2(n14253), .A(n13071), .B(n14294), .ZN(
        n14254) );
  INV_X1 U17638 ( .A(n14255), .ZN(n14256) );
  NAND2_X1 U17639 ( .A1(n14257), .A2(n14256), .ZN(n14963) );
  AOI22_X1 U17640 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14264) );
  AOI22_X1 U17641 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9717), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14262) );
  NAND2_X1 U17642 ( .A1(n14303), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n14258) );
  OAI211_X1 U17643 ( .C1(n14311), .C2(n14259), .A(n14258), .B(n14307), .ZN(
        n14260) );
  INV_X1 U17644 ( .A(n14260), .ZN(n14261) );
  NAND4_X1 U17645 ( .A1(n14264), .A2(n14263), .A3(n14262), .A4(n14261), .ZN(
        n14273) );
  AOI22_X1 U17646 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14271) );
  AOI22_X1 U17647 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10796), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14269) );
  NAND2_X1 U17648 ( .A1(n14125), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n14265) );
  OAI211_X1 U17649 ( .C1(n14311), .C2(n14266), .A(n14265), .B(n14277), .ZN(
        n14267) );
  INV_X1 U17650 ( .A(n14267), .ZN(n14268) );
  NAND4_X1 U17651 ( .A1(n14271), .A2(n14270), .A3(n14269), .A4(n14268), .ZN(
        n14272) );
  AND2_X1 U17652 ( .A1(n14273), .A2(n14272), .ZN(n14958) );
  OAI22_X1 U17653 ( .A1(n11002), .A2(n9762), .B1(n14274), .B2(n11004), .ZN(
        n14276) );
  INV_X1 U17654 ( .A(n14276), .ZN(n14284) );
  AOI22_X1 U17655 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9717), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14282) );
  NAND2_X1 U17656 ( .A1(n9763), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n14278) );
  OAI211_X1 U17657 ( .C1(n14311), .C2(n14279), .A(n14278), .B(n14277), .ZN(
        n14280) );
  INV_X1 U17658 ( .A(n14280), .ZN(n14281) );
  NAND4_X1 U17659 ( .A1(n14284), .A2(n14283), .A3(n14282), .A4(n14281), .ZN(
        n14293) );
  AOI22_X1 U17660 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14236), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14291) );
  AOI22_X1 U17661 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10796), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14289) );
  NAND2_X1 U17662 ( .A1(n14303), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n14285) );
  OAI211_X1 U17663 ( .C1(n14311), .C2(n14286), .A(n14285), .B(n14307), .ZN(
        n14287) );
  INV_X1 U17664 ( .A(n14287), .ZN(n14288) );
  NAND4_X1 U17665 ( .A1(n14291), .A2(n14290), .A3(n14289), .A4(n14288), .ZN(
        n14292) );
  AND2_X1 U17666 ( .A1(n14293), .A2(n14292), .ZN(n14297) );
  INV_X1 U17667 ( .A(n14294), .ZN(n14956) );
  NAND2_X1 U17668 ( .A1(n10757), .A2(n14958), .ZN(n14295) );
  NOR2_X1 U17669 ( .A1(n14956), .A2(n14295), .ZN(n14296) );
  NAND2_X1 U17670 ( .A1(n14296), .A2(n14297), .ZN(n14298) );
  OAI21_X1 U17671 ( .B1(n14297), .B2(n14296), .A(n14298), .ZN(n14952) );
  NOR2_X1 U17672 ( .A1(n14953), .A2(n14952), .ZN(n14951) );
  INV_X1 U17673 ( .A(n14298), .ZN(n14299) );
  NOR2_X1 U17674 ( .A1(n14951), .A2(n14299), .ZN(n14324) );
  AOI22_X1 U17675 ( .A1(n14236), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14315), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14300) );
  NAND2_X1 U17676 ( .A1(n14301), .A2(n14300), .ZN(n14322) );
  INV_X1 U17677 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14306) );
  AOI22_X1 U17678 ( .A1(n14302), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10796), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14305) );
  AOI21_X1 U17679 ( .B1(n14125), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n14307), .ZN(n14304) );
  OAI211_X1 U17680 ( .C1(n14311), .C2(n14306), .A(n14305), .B(n14304), .ZN(
        n14321) );
  INV_X1 U17681 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14308) );
  OAI21_X1 U17682 ( .B1(n14309), .B2(n14308), .A(n14307), .ZN(n14314) );
  INV_X1 U17683 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14312) );
  OAI22_X1 U17684 ( .A1(n10794), .A2(n14312), .B1(n14311), .B2(n14310), .ZN(
        n14313) );
  AOI211_X1 U17685 ( .C1(n9717), .C2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n14314), .B(n14313), .ZN(n14319) );
  AOI22_X1 U17686 ( .A1(n14316), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14315), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14318) );
  NAND3_X1 U17687 ( .A1(n14319), .A2(n14318), .A3(n14317), .ZN(n14320) );
  OAI21_X1 U17688 ( .B1(n14322), .B2(n14321), .A(n14320), .ZN(n14323) );
  XNOR2_X1 U17689 ( .A(n14324), .B(n14323), .ZN(n14334) );
  INV_X1 U17690 ( .A(n15048), .ZN(n14326) );
  NAND2_X1 U17691 ( .A1(n14326), .A2(n10177), .ZN(n14327) );
  NAND2_X1 U17692 ( .A1(n9805), .A2(n14327), .ZN(n15997) );
  OAI22_X1 U17693 ( .A1(n15997), .A2(n16092), .B1(n19103), .B2(n13238), .ZN(
        n14328) );
  AOI21_X1 U17694 ( .B1(n19082), .B2(n19093), .A(n14328), .ZN(n14330) );
  AOI22_X1 U17695 ( .A1(n19083), .A2(BUF1_REG_30__SCAN_IN), .B1(n19084), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n14329) );
  OAI211_X1 U17696 ( .C1(n14334), .C2(n19107), .A(n14330), .B(n14329), .ZN(
        P2_U2889) );
  NAND2_X1 U17697 ( .A1(n15999), .A2(n14992), .ZN(n14333) );
  NAND2_X1 U17698 ( .A1(n15040), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14332) );
  OAI211_X1 U17699 ( .C1(n14334), .C2(n15026), .A(n14333), .B(n14332), .ZN(
        P2_U2857) );
  NAND2_X1 U17700 ( .A1(n12962), .A2(n12593), .ZN(n14335) );
  NAND3_X1 U17701 ( .A1(n14337), .A2(n14336), .A3(n14335), .ZN(n14341) );
  INV_X1 U17702 ( .A(n14338), .ZN(n14339) );
  AOI22_X1 U17703 ( .A1(n14342), .A2(n14341), .B1(n14340), .B2(n14339), .ZN(
        n14347) );
  INV_X1 U17704 ( .A(n14343), .ZN(n14344) );
  NAND2_X1 U17705 ( .A1(n14351), .A2(n14344), .ZN(n14346) );
  AOI21_X1 U17706 ( .B1(n14347), .B2(n14346), .A(n14345), .ZN(n15592) );
  OAI22_X1 U17707 ( .A1(n14351), .A2(n14350), .B1(n11839), .B2(n14349), .ZN(
        n19895) );
  NAND3_X1 U17708 ( .A1(n14472), .A2(n15624), .A3(n12610), .ZN(n14352) );
  AND2_X1 U17709 ( .A1(n14352), .A2(n15977), .ZN(n20802) );
  NOR2_X1 U17710 ( .A1(n19895), .A2(n20802), .ZN(n15594) );
  NOR2_X1 U17711 ( .A1(n15594), .A2(n19894), .ZN(n19902) );
  MUX2_X1 U17712 ( .A(P1_MORE_REG_SCAN_IN), .B(n15592), .S(n19902), .Z(
        P1_U3484) );
  AOI22_X1 U17713 ( .A1(n14354), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n12610), .ZN(n14355) );
  NAND2_X1 U17714 ( .A1(n14357), .A2(n19949), .ZN(n14367) );
  NAND2_X1 U17715 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n14363) );
  INV_X1 U17716 ( .A(n14363), .ZN(n14361) );
  INV_X1 U17717 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20764) );
  NAND4_X1 U17718 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_14__SCAN_IN), .A4(P1_REIP_REG_13__SCAN_IN), .ZN(n14431) );
  INV_X1 U17719 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20749) );
  NAND2_X1 U17720 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14454) );
  NOR2_X1 U17721 ( .A1(n20749), .A2(n14454), .ZN(n14441) );
  NAND4_X1 U17722 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n14441), .A3(
        P1_REIP_REG_19__SCAN_IN), .A4(P1_REIP_REG_18__SCAN_IN), .ZN(n15680) );
  NAND4_X1 U17723 ( .A1(n15755), .A2(P1_REIP_REG_23__SCAN_IN), .A3(
        P1_REIP_REG_22__SCAN_IN), .A4(P1_REIP_REG_21__SCAN_IN), .ZN(n14358) );
  NOR3_X1 U17724 ( .A1(n14431), .A2(n15680), .A3(n14358), .ZN(n14419) );
  NAND2_X1 U17725 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14419), .ZN(n15661) );
  NOR2_X1 U17726 ( .A1(n20764), .A2(n15661), .ZN(n15648) );
  NAND2_X1 U17727 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n15648), .ZN(n14405) );
  INV_X1 U17728 ( .A(n14405), .ZN(n14359) );
  AND2_X1 U17729 ( .A1(n14417), .A2(n14359), .ZN(n15646) );
  NAND3_X1 U17730 ( .A1(n15646), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14360) );
  NAND2_X1 U17731 ( .A1(n19989), .A2(n14360), .ZN(n14394) );
  OAI21_X1 U17732 ( .B1(n15647), .B2(n14361), .A(n14394), .ZN(n14374) );
  INV_X1 U17733 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14491) );
  OAI22_X1 U17734 ( .A1(n19946), .A2(n14491), .B1(n14362), .B2(n19993), .ZN(
        n14365) );
  INV_X1 U17735 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20766) );
  NOR3_X1 U17736 ( .A1(n15662), .A2(n14405), .A3(n20766), .ZN(n14396) );
  NAND2_X1 U17737 ( .A1(n14396), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14382) );
  NOR3_X1 U17738 ( .A1(n14382), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14363), 
        .ZN(n14364) );
  AOI211_X1 U17739 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14374), .A(n14365), 
        .B(n14364), .ZN(n14366) );
  OAI211_X1 U17740 ( .C1(n14756), .C2(n19988), .A(n14367), .B(n14366), .ZN(
        P1_U2809) );
  INV_X1 U17741 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20772) );
  INV_X1 U17742 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14368) );
  OAI21_X1 U17743 ( .B1(n14382), .B2(n20772), .A(n14368), .ZN(n14373) );
  AOI22_X1 U17744 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19975), .B1(
        n19982), .B2(n14625), .ZN(n14369) );
  OAI21_X1 U17745 ( .B1(n19946), .B2(n14370), .A(n14369), .ZN(n14372) );
  NOR2_X1 U17746 ( .A1(n14780), .A2(n19988), .ZN(n14371) );
  OAI21_X1 U17747 ( .B1(n14629), .B2(n15751), .A(n14375), .ZN(P1_U2810) );
  AOI21_X1 U17748 ( .B1(n14378), .B2(n14376), .A(n14377), .ZN(n14636) );
  INV_X1 U17749 ( .A(n14636), .ZN(n14570) );
  AOI21_X1 U17750 ( .B1(n14380), .B2(n14393), .A(n14379), .ZN(n14790) );
  OAI22_X1 U17751 ( .A1(n14381), .A2(n19993), .B1(n19992), .B2(n14634), .ZN(
        n14384) );
  NOR2_X1 U17752 ( .A1(n14382), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14383) );
  AOI211_X1 U17753 ( .C1(P1_EBX_REG_29__SCAN_IN), .C2(n19994), .A(n14384), .B(
        n14383), .ZN(n14385) );
  OAI21_X1 U17754 ( .B1(n20772), .B2(n14394), .A(n14385), .ZN(n14386) );
  AOI21_X1 U17755 ( .B1(n14790), .B2(n19991), .A(n14386), .ZN(n14387) );
  OAI21_X1 U17756 ( .B1(n14570), .B2(n15751), .A(n14387), .ZN(P1_U2811) );
  NAND2_X1 U17757 ( .A1(n14390), .A2(n14391), .ZN(n14392) );
  INV_X1 U17758 ( .A(n14394), .ZN(n14395) );
  OAI21_X1 U17759 ( .B1(n14396), .B2(P1_REIP_REG_28__SCAN_IN), .A(n14395), 
        .ZN(n14398) );
  AOI22_X1 U17760 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19975), .B1(
        n19982), .B2(n14641), .ZN(n14397) );
  OAI211_X1 U17761 ( .C1(n19946), .C2(n14493), .A(n14398), .B(n14397), .ZN(
        n14399) );
  AOI21_X1 U17762 ( .B1(n14805), .B2(n19991), .A(n14399), .ZN(n14400) );
  OAI21_X1 U17763 ( .B1(n14651), .B2(n15751), .A(n14400), .ZN(P1_U2812) );
  OR2_X1 U17764 ( .A1(n14502), .A2(n14401), .ZN(n14402) );
  NAND2_X1 U17765 ( .A1(n14390), .A2(n14402), .ZN(n14813) );
  AOI21_X1 U17766 ( .B1(n14404), .B2(n14403), .A(n14388), .ZN(n14659) );
  NAND2_X1 U17767 ( .A1(n14659), .A2(n19949), .ZN(n14411) );
  NOR3_X1 U17768 ( .A1(n15647), .A2(n15646), .A3(n20766), .ZN(n14409) );
  NOR3_X1 U17769 ( .A1(n15662), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14405), 
        .ZN(n14408) );
  INV_X1 U17770 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14496) );
  NOR2_X1 U17771 ( .A1(n19946), .A2(n14496), .ZN(n14407) );
  OAI22_X1 U17772 ( .A1(n12453), .A2(n19993), .B1(n19992), .B2(n14657), .ZN(
        n14406) );
  NOR4_X1 U17773 ( .A1(n14409), .A2(n14408), .A3(n14407), .A4(n14406), .ZN(
        n14410) );
  OAI211_X1 U17774 ( .C1(n19988), .C2(n14813), .A(n14411), .B(n14410), .ZN(
        P1_U2813) );
  INV_X1 U17775 ( .A(n14412), .ZN(n14514) );
  AOI21_X1 U17776 ( .B1(n14414), .B2(n14514), .A(n14413), .ZN(n14682) );
  INV_X1 U17777 ( .A(n14682), .ZN(n14592) );
  XNOR2_X1 U17778 ( .A(n14519), .B(n14506), .ZN(n15853) );
  NOR2_X1 U17779 ( .A1(n19946), .A2(n14415), .ZN(n14423) );
  INV_X1 U17780 ( .A(n14416), .ZN(n14680) );
  NOR2_X1 U17781 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15662), .ZN(n14418) );
  OAI21_X1 U17782 ( .B1(n14419), .B2(n15662), .A(n14417), .ZN(n15673) );
  AOI22_X1 U17783 ( .A1(n14419), .A2(n14418), .B1(P1_REIP_REG_24__SCAN_IN), 
        .B2(n15673), .ZN(n14421) );
  NAND2_X1 U17784 ( .A1(n19975), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14420) );
  OAI211_X1 U17785 ( .C1(n19992), .C2(n14680), .A(n14421), .B(n14420), .ZN(
        n14422) );
  AOI211_X1 U17786 ( .C1(n15853), .C2(n19991), .A(n14423), .B(n14422), .ZN(
        n14424) );
  OAI21_X1 U17787 ( .B1(n14592), .B2(n15751), .A(n14424), .ZN(P1_U2816) );
  OAI21_X1 U17788 ( .B1(n14425), .B2(n10233), .A(n14426), .ZN(n14699) );
  XNOR2_X1 U17789 ( .A(n14541), .B(n14534), .ZN(n14538) );
  INV_X1 U17790 ( .A(n14538), .ZN(n15632) );
  INV_X1 U17791 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14537) );
  NOR2_X1 U17792 ( .A1(n19946), .A2(n14537), .ZN(n14430) );
  INV_X1 U17793 ( .A(n14427), .ZN(n14695) );
  OAI22_X1 U17794 ( .A1(n14695), .A2(n19992), .B1(n19993), .B2(n14428), .ZN(
        n14429) );
  AOI211_X1 U17795 ( .C1(n15632), .C2(n19991), .A(n14430), .B(n14429), .ZN(
        n14436) );
  AOI21_X1 U17796 ( .B1(n14431), .B2(n19989), .A(n15761), .ZN(n15740) );
  INV_X1 U17797 ( .A(n15740), .ZN(n15721) );
  AOI21_X1 U17798 ( .B1(n15680), .B2(n19989), .A(n15721), .ZN(n14432) );
  INV_X1 U17799 ( .A(n14432), .ZN(n15691) );
  NAND2_X1 U17800 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14433) );
  NAND3_X1 U17801 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(n15729), .ZN(n15728) );
  INV_X1 U17802 ( .A(n15728), .ZN(n14455) );
  NAND2_X1 U17803 ( .A1(n14441), .A2(n14455), .ZN(n15703) );
  INV_X1 U17804 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20754) );
  OAI21_X1 U17805 ( .B1(n14433), .B2(n15703), .A(n20754), .ZN(n14434) );
  NAND2_X1 U17806 ( .A1(n15691), .A2(n14434), .ZN(n14435) );
  OAI211_X1 U17807 ( .C1(n14699), .C2(n15751), .A(n14436), .B(n14435), .ZN(
        P1_U2820) );
  INV_X1 U17808 ( .A(n14437), .ZN(n14440) );
  INV_X1 U17809 ( .A(n14438), .ZN(n14439) );
  AOI21_X1 U17810 ( .B1(n14440), .B2(n14439), .A(n14547), .ZN(n15799) );
  INV_X1 U17811 ( .A(n15799), .ZN(n14616) );
  OAI21_X1 U17812 ( .B1(n14441), .B2(n15647), .A(n15740), .ZN(n15718) );
  OAI21_X1 U17813 ( .B1(n14454), .B2(n15728), .A(n20749), .ZN(n14449) );
  INV_X1 U17814 ( .A(n14458), .ZN(n14444) );
  INV_X1 U17815 ( .A(n14442), .ZN(n14443) );
  OAI21_X1 U17816 ( .B1(n14444), .B2(n14443), .A(n14551), .ZN(n15876) );
  NAND2_X1 U17817 ( .A1(n19982), .A2(n15798), .ZN(n14445) );
  OAI211_X1 U17818 ( .C1(n19993), .C2(n20990), .A(n19954), .B(n14445), .ZN(
        n14446) );
  AOI21_X1 U17819 ( .B1(n19994), .B2(P1_EBX_REG_17__SCAN_IN), .A(n14446), .ZN(
        n14447) );
  OAI21_X1 U17820 ( .B1(n15876), .B2(n19988), .A(n14447), .ZN(n14448) );
  AOI21_X1 U17821 ( .B1(n15718), .B2(n14449), .A(n14448), .ZN(n14450) );
  OAI21_X1 U17822 ( .B1(n14616), .B2(n15751), .A(n14450), .ZN(P1_U2823) );
  AOI21_X1 U17823 ( .B1(n14452), .B2(n14451), .A(n14438), .ZN(n14716) );
  INV_X1 U17824 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20748) );
  AOI22_X1 U17825 ( .A1(n19994), .A2(P1_EBX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19975), .ZN(n14453) );
  OAI211_X1 U17826 ( .C1(n15740), .C2(n20748), .A(n14453), .B(n19954), .ZN(
        n14463) );
  OAI211_X1 U17827 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n14455), .B(n14454), .ZN(n14461) );
  NAND2_X1 U17828 ( .A1(n14560), .A2(n14456), .ZN(n14457) );
  NAND2_X1 U17829 ( .A1(n14458), .A2(n14457), .ZN(n14860) );
  NOR2_X1 U17830 ( .A1(n19988), .A2(n14860), .ZN(n14459) );
  AOI21_X1 U17831 ( .B1(n19982), .B2(n14712), .A(n14459), .ZN(n14460) );
  NAND2_X1 U17832 ( .A1(n14461), .A2(n14460), .ZN(n14462) );
  AOI211_X1 U17833 ( .C1(n14716), .C2(n19949), .A(n14463), .B(n14462), .ZN(
        n14464) );
  INV_X1 U17834 ( .A(n14464), .ZN(P1_U2824) );
  AOI21_X1 U17835 ( .B1(n19975), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19964), .ZN(n14466) );
  AOI22_X1 U17836 ( .A1(n15761), .A2(P1_REIP_REG_10__SCAN_IN), .B1(n19994), 
        .B2(P1_EBX_REG_10__SCAN_IN), .ZN(n14465) );
  OAI211_X1 U17837 ( .C1(n19988), .C2(n15927), .A(n14466), .B(n14465), .ZN(
        n14470) );
  NOR3_X1 U17838 ( .A1(n20737), .A2(n14467), .A3(n19959), .ZN(n19921) );
  INV_X1 U17839 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21000) );
  NAND3_X1 U17840 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19921), .A3(n21000), 
        .ZN(n14468) );
  OAI21_X1 U17841 ( .B1(n14751), .B2(n19992), .A(n14468), .ZN(n14469) );
  AOI211_X1 U17842 ( .C1(n14753), .C2(n19949), .A(n14470), .B(n14469), .ZN(
        n14471) );
  INV_X1 U17843 ( .A(n14471), .ZN(P1_U2830) );
  OR2_X1 U17844 ( .A1(n14475), .A2(n14472), .ZN(n14473) );
  NOR2_X1 U17845 ( .A1(n14475), .A2(n14474), .ZN(n19995) );
  AOI22_X1 U17846 ( .A1(n19975), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n19974), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n14476) );
  OAI21_X1 U17847 ( .B1(n19992), .B2(n14477), .A(n14476), .ZN(n14479) );
  AOI211_X1 U17848 ( .C1(n19984), .C2(n20728), .A(n19965), .B(n15662), .ZN(
        n14478) );
  AOI211_X1 U17849 ( .C1(n19995), .C2(n20399), .A(n14479), .B(n14478), .ZN(
        n14481) );
  AOI22_X1 U17850 ( .A1(n19994), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n19991), .B2(
        n20095), .ZN(n14480) );
  OAI211_X1 U17851 ( .C1(n19999), .C2(n14482), .A(n14481), .B(n14480), .ZN(
        P1_U2837) );
  OAI22_X1 U17852 ( .A1(n19999), .A2(n14484), .B1(n19946), .B2(n14483), .ZN(
        n14490) );
  OAI22_X1 U17853 ( .A1(n19988), .A2(n14485), .B1(P1_REIP_REG_1__SCAN_IN), 
        .B2(n15662), .ZN(n14489) );
  INV_X1 U17854 ( .A(n20521), .ZN(n20598) );
  NAND2_X1 U17855 ( .A1(n19995), .A2(n20598), .ZN(n14487) );
  AOI22_X1 U17856 ( .A1(n19975), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n19974), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14486) );
  OAI211_X1 U17857 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19992), .A(
        n14487), .B(n14486), .ZN(n14488) );
  OR3_X1 U17858 ( .A1(n14490), .A2(n14489), .A3(n14488), .ZN(P1_U2839) );
  OAI22_X1 U17859 ( .A1(n14756), .A2(n20001), .B1(n14491), .B2(n20012), .ZN(
        P1_U2841) );
  AOI22_X1 U17860 ( .A1(n14790), .A2(n20007), .B1(n14520), .B2(
        P1_EBX_REG_29__SCAN_IN), .ZN(n14492) );
  OAI21_X1 U17861 ( .B1(n14570), .B2(n14561), .A(n14492), .ZN(P1_U2843) );
  NOR2_X1 U17862 ( .A1(n20012), .A2(n14493), .ZN(n14494) );
  AOI21_X1 U17863 ( .B1(n14805), .B2(n20007), .A(n14494), .ZN(n14495) );
  OAI21_X1 U17864 ( .B1(n14651), .B2(n14561), .A(n14495), .ZN(P1_U2844) );
  INV_X1 U17865 ( .A(n14659), .ZN(n14579) );
  OAI222_X1 U17866 ( .A1(n14496), .A2(n20012), .B1(n20001), .B2(n14813), .C1(
        n14579), .C2(n14561), .ZN(P1_U2845) );
  OR2_X1 U17867 ( .A1(n14497), .A2(n14498), .ZN(n14499) );
  INV_X1 U17868 ( .A(n15656), .ZN(n14583) );
  NOR2_X1 U17869 ( .A1(n14508), .A2(n14500), .ZN(n14501) );
  OR2_X1 U17870 ( .A1(n14502), .A2(n14501), .ZN(n15659) );
  OAI22_X1 U17871 ( .A1(n15659), .A2(n20001), .B1(n15651), .B2(n20012), .ZN(
        n14503) );
  INV_X1 U17872 ( .A(n14503), .ZN(n14504) );
  OAI21_X1 U17873 ( .B1(n14583), .B2(n14561), .A(n14504), .ZN(P1_U2846) );
  INV_X1 U17874 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15663) );
  INV_X1 U17875 ( .A(n14519), .ZN(n14507) );
  AOI21_X1 U17876 ( .B1(n14507), .B2(n14506), .A(n14505), .ZN(n14509) );
  OR2_X1 U17877 ( .A1(n14509), .A2(n14508), .ZN(n15667) );
  NOR2_X1 U17878 ( .A1(n14413), .A2(n14510), .ZN(n14511) );
  OR2_X1 U17879 ( .A1(n14497), .A2(n14511), .ZN(n15668) );
  OAI222_X1 U17880 ( .A1(n15663), .A2(n20012), .B1(n20001), .B2(n15667), .C1(
        n15668), .C2(n14561), .ZN(P1_U2847) );
  AOI22_X1 U17881 ( .A1(n15853), .A2(n20007), .B1(n14520), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n14512) );
  OAI21_X1 U17882 ( .B1(n14592), .B2(n14561), .A(n14512), .ZN(P1_U2848) );
  INV_X1 U17883 ( .A(n14514), .ZN(n14515) );
  AOI21_X1 U17884 ( .B1(n14516), .B2(n14513), .A(n14515), .ZN(n15774) );
  INV_X1 U17885 ( .A(n15774), .ZN(n14598) );
  NAND2_X1 U17886 ( .A1(n14528), .A2(n14517), .ZN(n14518) );
  AND2_X1 U17887 ( .A1(n14519), .A2(n14518), .ZN(n15860) );
  AOI22_X1 U17888 ( .A1(n15860), .A2(n20007), .B1(n14520), .B2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n14521) );
  OAI21_X1 U17889 ( .B1(n14598), .B2(n14561), .A(n14521), .ZN(P1_U2849) );
  OAI21_X1 U17890 ( .B1(n14523), .B2(n14524), .A(n14513), .ZN(n15687) );
  OR2_X1 U17891 ( .A1(n14525), .A2(n14526), .ZN(n14527) );
  NAND2_X1 U17892 ( .A1(n14528), .A2(n14527), .ZN(n15690) );
  OAI22_X1 U17893 ( .A1(n15690), .A2(n20001), .B1(n15683), .B2(n20012), .ZN(
        n14529) );
  INV_X1 U17894 ( .A(n14529), .ZN(n14530) );
  OAI21_X1 U17895 ( .B1(n15687), .B2(n14561), .A(n14530), .ZN(P1_U2850) );
  INV_X1 U17896 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14536) );
  AND2_X1 U17897 ( .A1(n14426), .A2(n14531), .ZN(n14532) );
  OR2_X1 U17898 ( .A1(n14532), .A2(n14523), .ZN(n15778) );
  AOI21_X1 U17899 ( .B1(n14541), .B2(n14534), .A(n14533), .ZN(n14535) );
  OR2_X1 U17900 ( .A1(n14525), .A2(n14535), .ZN(n15693) );
  OAI222_X1 U17901 ( .A1(n14536), .A2(n20012), .B1(n14561), .B2(n15778), .C1(
        n15693), .C2(n20001), .ZN(P1_U2851) );
  OAI222_X1 U17902 ( .A1(n14699), .A2(n14561), .B1(n20001), .B2(n14538), .C1(
        n20012), .C2(n14537), .ZN(P1_U2852) );
  INV_X1 U17903 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14545) );
  NOR2_X1 U17904 ( .A1(n14552), .A2(n14539), .ZN(n14540) );
  OR2_X1 U17905 ( .A1(n14541), .A2(n14540), .ZN(n15867) );
  NAND2_X1 U17906 ( .A1(n14549), .A2(n14542), .ZN(n14543) );
  AND2_X1 U17907 ( .A1(n14544), .A2(n14543), .ZN(n15788) );
  INV_X1 U17908 ( .A(n15788), .ZN(n14607) );
  OAI222_X1 U17909 ( .A1(n14545), .A2(n20012), .B1(n20001), .B2(n15867), .C1(
        n14607), .C2(n14561), .ZN(P1_U2853) );
  OR2_X1 U17910 ( .A1(n14547), .A2(n14546), .ZN(n14548) );
  NAND2_X1 U17911 ( .A1(n14549), .A2(n14548), .ZN(n15715) );
  AND2_X1 U17912 ( .A1(n14551), .A2(n14550), .ZN(n14553) );
  OR2_X1 U17913 ( .A1(n14553), .A2(n14552), .ZN(n15720) );
  OAI22_X1 U17914 ( .A1(n15720), .A2(n20001), .B1(n15714), .B2(n20012), .ZN(
        n14554) );
  INV_X1 U17915 ( .A(n14554), .ZN(n14555) );
  OAI21_X1 U17916 ( .B1(n15715), .B2(n14561), .A(n14555), .ZN(P1_U2854) );
  INV_X1 U17917 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14556) );
  OAI222_X1 U17918 ( .A1(n15876), .A2(n20001), .B1(n14556), .B2(n20012), .C1(
        n14561), .C2(n14616), .ZN(P1_U2855) );
  INV_X1 U17919 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n14557) );
  INV_X1 U17920 ( .A(n14716), .ZN(n14622) );
  OAI222_X1 U17921 ( .A1(n14860), .A2(n20001), .B1(n20012), .B2(n14557), .C1(
        n14561), .C2(n14622), .ZN(P1_U2856) );
  OR2_X1 U17922 ( .A1(n9839), .A2(n14558), .ZN(n14559) );
  NAND2_X1 U17923 ( .A1(n14560), .A2(n14559), .ZN(n15884) );
  INV_X1 U17924 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14563) );
  OAI222_X1 U17925 ( .A1(n15884), .A2(n20001), .B1(n14563), .B2(n20012), .C1(
        n14562), .C2(n14561), .ZN(P1_U2857) );
  AOI22_X1 U17926 ( .A1(n14617), .A2(BUF1_REG_30__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n14566) );
  NOR2_X2 U17927 ( .A1(n15768), .A2(n14564), .ZN(n14618) );
  AOI22_X1 U17928 ( .A1(n14619), .A2(DATAI_30_), .B1(n14618), .B2(n20059), 
        .ZN(n14565) );
  OAI211_X1 U17929 ( .C1(n14629), .C2(n20016), .A(n14566), .B(n14565), .ZN(
        P1_U2874) );
  AOI22_X1 U17930 ( .A1(n14617), .A2(BUF1_REG_29__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n14569) );
  AOI22_X1 U17931 ( .A1(n14619), .A2(DATAI_29_), .B1(n14618), .B2(n14567), 
        .ZN(n14568) );
  OAI211_X1 U17932 ( .C1(n14570), .C2(n20016), .A(n14569), .B(n14568), .ZN(
        P1_U2875) );
  AOI22_X1 U17933 ( .A1(n14617), .A2(BUF1_REG_28__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n14574) );
  INV_X1 U17934 ( .A(DATAI_12_), .ZN(n14572) );
  NAND2_X1 U17935 ( .A1(n20143), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14571) );
  OAI21_X1 U17936 ( .B1(n20143), .B2(n14572), .A(n14571), .ZN(n20057) );
  AOI22_X1 U17937 ( .A1(n14619), .A2(DATAI_28_), .B1(n14618), .B2(n20057), 
        .ZN(n14573) );
  OAI211_X1 U17938 ( .C1(n14651), .C2(n20016), .A(n14574), .B(n14573), .ZN(
        P1_U2876) );
  AOI22_X1 U17939 ( .A1(n14617), .A2(BUF1_REG_27__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n14578) );
  INV_X1 U17940 ( .A(DATAI_11_), .ZN(n14576) );
  NAND2_X1 U17941 ( .A1(n20143), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14575) );
  OAI21_X1 U17942 ( .B1(n20143), .B2(n14576), .A(n14575), .ZN(n20055) );
  AOI22_X1 U17943 ( .A1(n14619), .A2(DATAI_27_), .B1(n14618), .B2(n20055), 
        .ZN(n14577) );
  OAI211_X1 U17944 ( .C1(n14579), .C2(n20016), .A(n14578), .B(n14577), .ZN(
        P1_U2877) );
  AOI22_X1 U17945 ( .A1(n14617), .A2(BUF1_REG_26__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_26__SCAN_IN), .ZN(n14582) );
  AOI22_X1 U17946 ( .A1(n14619), .A2(DATAI_26_), .B1(n14618), .B2(n14580), 
        .ZN(n14581) );
  OAI211_X1 U17947 ( .C1(n14583), .C2(n20016), .A(n14582), .B(n14581), .ZN(
        P1_U2878) );
  AOI22_X1 U17948 ( .A1(n14617), .A2(BUF1_REG_25__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n14585) );
  AOI22_X1 U17949 ( .A1(n14619), .A2(DATAI_25_), .B1(n14618), .B2(n20053), 
        .ZN(n14584) );
  OAI211_X1 U17950 ( .C1(n15668), .C2(n20016), .A(n14585), .B(n14584), .ZN(
        P1_U2879) );
  INV_X1 U17951 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n14587) );
  INV_X1 U17952 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14586) );
  OAI22_X1 U17953 ( .A1(n14612), .A2(n14587), .B1(n14586), .B2(n20015), .ZN(
        n14588) );
  INV_X1 U17954 ( .A(n14588), .ZN(n14591) );
  AOI22_X1 U17955 ( .A1(n14619), .A2(DATAI_24_), .B1(n14618), .B2(n14589), 
        .ZN(n14590) );
  OAI211_X1 U17956 ( .C1(n14592), .C2(n20016), .A(n14591), .B(n14590), .ZN(
        P1_U2880) );
  INV_X1 U17957 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n14594) );
  OAI22_X1 U17958 ( .A1(n14612), .A2(n14594), .B1(n14593), .B2(n20015), .ZN(
        n14595) );
  INV_X1 U17959 ( .A(n14595), .ZN(n14597) );
  AOI22_X1 U17960 ( .A1(n14619), .A2(DATAI_23_), .B1(n14618), .B2(n20186), 
        .ZN(n14596) );
  OAI211_X1 U17961 ( .C1(n14598), .C2(n20016), .A(n14597), .B(n14596), .ZN(
        P1_U2881) );
  AOI22_X1 U17962 ( .A1(n14617), .A2(BUF1_REG_22__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n14600) );
  AOI22_X1 U17963 ( .A1(n14619), .A2(DATAI_22_), .B1(n14618), .B2(n20180), 
        .ZN(n14599) );
  OAI211_X1 U17964 ( .C1(n15687), .C2(n20016), .A(n14600), .B(n14599), .ZN(
        P1_U2882) );
  AOI22_X1 U17965 ( .A1(n14617), .A2(BUF1_REG_21__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_21__SCAN_IN), .ZN(n14602) );
  AOI22_X1 U17966 ( .A1(n14619), .A2(DATAI_21_), .B1(n14618), .B2(n20175), 
        .ZN(n14601) );
  OAI211_X1 U17967 ( .C1(n15778), .C2(n20016), .A(n14602), .B(n14601), .ZN(
        P1_U2883) );
  AOI22_X1 U17968 ( .A1(n14617), .A2(BUF1_REG_20__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_20__SCAN_IN), .ZN(n14604) );
  AOI22_X1 U17969 ( .A1(n14619), .A2(DATAI_20_), .B1(n14618), .B2(n20169), 
        .ZN(n14603) );
  OAI211_X1 U17970 ( .C1(n14699), .C2(n20016), .A(n14604), .B(n14603), .ZN(
        P1_U2884) );
  AOI22_X1 U17971 ( .A1(n14617), .A2(BUF1_REG_19__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_19__SCAN_IN), .ZN(n14606) );
  AOI22_X1 U17972 ( .A1(n14619), .A2(DATAI_19_), .B1(n14618), .B2(n20164), 
        .ZN(n14605) );
  OAI211_X1 U17973 ( .C1(n14607), .C2(n20016), .A(n14606), .B(n14605), .ZN(
        P1_U2885) );
  AOI22_X1 U17974 ( .A1(n14617), .A2(BUF1_REG_18__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n14609) );
  AOI22_X1 U17975 ( .A1(n14619), .A2(DATAI_18_), .B1(n14618), .B2(n20159), 
        .ZN(n14608) );
  OAI211_X1 U17976 ( .C1(n15715), .C2(n20016), .A(n14609), .B(n14608), .ZN(
        P1_U2886) );
  INV_X1 U17977 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14611) );
  OAI22_X1 U17978 ( .A1(n14612), .A2(n14611), .B1(n14610), .B2(n20015), .ZN(
        n14613) );
  INV_X1 U17979 ( .A(n14613), .ZN(n14615) );
  AOI22_X1 U17980 ( .A1(n14619), .A2(DATAI_17_), .B1(n14618), .B2(n20154), 
        .ZN(n14614) );
  OAI211_X1 U17981 ( .C1(n14616), .C2(n20016), .A(n14615), .B(n14614), .ZN(
        P1_U2887) );
  AOI22_X1 U17982 ( .A1(n14617), .A2(BUF1_REG_16__SCAN_IN), .B1(n15768), .B2(
        P1_EAX_REG_16__SCAN_IN), .ZN(n14621) );
  AOI22_X1 U17983 ( .A1(n14619), .A2(DATAI_16_), .B1(n14618), .B2(n20141), 
        .ZN(n14620) );
  OAI211_X1 U17984 ( .C1(n14622), .C2(n20016), .A(n14621), .B(n14620), .ZN(
        P1_U2888) );
  NAND2_X1 U17985 ( .A1(n13397), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14781) );
  OAI21_X1 U17986 ( .B1(n15784), .B2(n14623), .A(n14781), .ZN(n14624) );
  AOI21_X1 U17987 ( .B1(n14625), .B2(n15820), .A(n14624), .ZN(n14628) );
  NAND2_X1 U17988 ( .A1(n14779), .A2(n20081), .ZN(n14627) );
  OAI211_X1 U17989 ( .C1(n14629), .C2(n20142), .A(n14628), .B(n14627), .ZN(
        P1_U2969) );
  MUX2_X1 U17990 ( .A(n14631), .B(n14630), .S(n15794), .Z(n14632) );
  XNOR2_X1 U17991 ( .A(n14632), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14799) );
  NOR2_X1 U17992 ( .A1(n20107), .A2(n20772), .ZN(n14793) );
  AOI21_X1 U17993 ( .B1(n20076), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14793), .ZN(n14633) );
  OAI21_X1 U17994 ( .B1(n20085), .B2(n14634), .A(n14633), .ZN(n14635) );
  AOI21_X1 U17995 ( .B1(n14636), .B2(n14666), .A(n14635), .ZN(n14637) );
  OAI21_X1 U17996 ( .B1(n19900), .B2(n14799), .A(n14637), .ZN(P1_U2970) );
  INV_X1 U17997 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14638) );
  NOR2_X1 U17998 ( .A1(n20107), .A2(n14638), .ZN(n14803) );
  NOR2_X1 U17999 ( .A1(n15784), .A2(n14639), .ZN(n14640) );
  AOI211_X1 U18000 ( .C1(n15820), .C2(n14641), .A(n14803), .B(n14640), .ZN(
        n14650) );
  NAND2_X1 U18001 ( .A1(n9738), .A2(n14643), .ZN(n14661) );
  NAND2_X1 U18002 ( .A1(n14642), .A2(n14661), .ZN(n14647) );
  OAI21_X1 U18003 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14644), .A(
        n14647), .ZN(n14646) );
  INV_X1 U18004 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14816) );
  MUX2_X1 U18005 ( .A(n14816), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n9738), .Z(n14645) );
  OAI211_X1 U18006 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14647), .A(
        n14646), .B(n14645), .ZN(n14648) );
  XNOR2_X1 U18007 ( .A(n14648), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14800) );
  NAND2_X1 U18008 ( .A1(n14800), .A2(n20081), .ZN(n14649) );
  OAI211_X1 U18009 ( .C1(n14651), .C2(n20142), .A(n14650), .B(n14649), .ZN(
        P1_U2971) );
  INV_X1 U18010 ( .A(n14652), .ZN(n14654) );
  MUX2_X1 U18011 ( .A(n14654), .B(n14653), .S(n15794), .Z(n14655) );
  NOR2_X1 U18012 ( .A1(n20107), .A2(n20766), .ZN(n14810) );
  AOI21_X1 U18013 ( .B1(n20076), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14810), .ZN(n14656) );
  OAI21_X1 U18014 ( .B1(n20085), .B2(n14657), .A(n14656), .ZN(n14658) );
  AOI21_X1 U18015 ( .B1(n14659), .B2(n14666), .A(n14658), .ZN(n14660) );
  OAI21_X1 U18016 ( .B1(n19900), .B2(n14814), .A(n14660), .ZN(P1_U2972) );
  OAI211_X1 U18017 ( .C1(n15794), .C2(n14642), .A(n14662), .B(n14661), .ZN(
        n14663) );
  XNOR2_X1 U18018 ( .A(n14663), .B(n14824), .ZN(n14830) );
  NAND2_X1 U18019 ( .A1(n15820), .A2(n15655), .ZN(n14664) );
  NAND2_X1 U18020 ( .A1(n13397), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14818) );
  OAI211_X1 U18021 ( .C1(n15784), .C2(n15650), .A(n14664), .B(n14818), .ZN(
        n14665) );
  AOI21_X1 U18022 ( .B1(n15656), .B2(n14666), .A(n14665), .ZN(n14667) );
  OAI21_X1 U18023 ( .B1(n19900), .B2(n14830), .A(n14667), .ZN(P1_U2973) );
  NOR2_X1 U18024 ( .A1(n20107), .A2(n20764), .ZN(n14833) );
  NOR2_X1 U18025 ( .A1(n20085), .A2(n15672), .ZN(n14668) );
  AOI211_X1 U18026 ( .C1(n20076), .C2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14833), .B(n14668), .ZN(n14674) );
  NOR3_X1 U18027 ( .A1(n14642), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14671) );
  NAND2_X1 U18028 ( .A1(n14669), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14677) );
  NOR2_X1 U18029 ( .A1(n14677), .A2(n15851), .ZN(n14670) );
  MUX2_X1 U18030 ( .A(n14671), .B(n14670), .S(n9738), .Z(n14672) );
  XNOR2_X1 U18031 ( .A(n14672), .B(n14820), .ZN(n14831) );
  NAND2_X1 U18032 ( .A1(n14831), .A2(n20081), .ZN(n14673) );
  OAI211_X1 U18033 ( .C1(n15668), .C2(n20142), .A(n14674), .B(n14673), .ZN(
        P1_U2974) );
  INV_X1 U18034 ( .A(n14642), .ZN(n14675) );
  NAND2_X1 U18035 ( .A1(n14675), .A2(n14677), .ZN(n14676) );
  MUX2_X1 U18036 ( .A(n14677), .B(n14676), .S(n15794), .Z(n14678) );
  XNOR2_X1 U18037 ( .A(n14678), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15854) );
  INV_X1 U18038 ( .A(n15854), .ZN(n14684) );
  AOI22_X1 U18039 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n14679) );
  OAI21_X1 U18040 ( .B1(n20085), .B2(n14680), .A(n14679), .ZN(n14681) );
  AOI21_X1 U18041 ( .B1(n14682), .B2(n14666), .A(n14681), .ZN(n14683) );
  OAI21_X1 U18042 ( .B1(n19900), .B2(n14684), .A(n14683), .ZN(P1_U2975) );
  NAND2_X1 U18043 ( .A1(n14686), .A2(n14685), .ZN(n14688) );
  XNOR2_X1 U18044 ( .A(n14688), .B(n14687), .ZN(n14846) );
  NAND2_X1 U18045 ( .A1(n13397), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n14840) );
  OAI21_X1 U18046 ( .B1(n15784), .B2(n12361), .A(n14840), .ZN(n14690) );
  NOR2_X1 U18047 ( .A1(n15687), .A2(n20142), .ZN(n14689) );
  AOI211_X1 U18048 ( .C1(n15820), .C2(n15681), .A(n14690), .B(n14689), .ZN(
        n14691) );
  OAI21_X1 U18049 ( .B1(n19900), .B2(n14846), .A(n14691), .ZN(P1_U2977) );
  NOR2_X1 U18050 ( .A1(n9738), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15786) );
  NAND2_X1 U18051 ( .A1(n10110), .A2(n15786), .ZN(n15606) );
  INV_X1 U18052 ( .A(n14692), .ZN(n14693) );
  NAND3_X1 U18053 ( .A1(n14693), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n9738), .ZN(n15609) );
  OAI21_X1 U18054 ( .B1(n15606), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15609), .ZN(n14694) );
  INV_X1 U18055 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15608) );
  XNOR2_X1 U18056 ( .A(n14694), .B(n15608), .ZN(n15633) );
  NAND2_X1 U18057 ( .A1(n15633), .A2(n20081), .ZN(n14698) );
  NOR2_X1 U18058 ( .A1(n20107), .A2(n20754), .ZN(n15634) );
  NOR2_X1 U18059 ( .A1(n20085), .A2(n14695), .ZN(n14696) );
  AOI211_X1 U18060 ( .C1(n20076), .C2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15634), .B(n14696), .ZN(n14697) );
  OAI211_X1 U18061 ( .C1(n20142), .C2(n14699), .A(n14698), .B(n14697), .ZN(
        P1_U2979) );
  NAND2_X1 U18062 ( .A1(n13397), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14849) );
  OAI21_X1 U18063 ( .B1(n15784), .B2(n15709), .A(n14849), .ZN(n14700) );
  AOI21_X1 U18064 ( .B1(n15711), .B2(n15820), .A(n14700), .ZN(n14704) );
  OR2_X1 U18065 ( .A1(n14702), .A2(n14701), .ZN(n14847) );
  NAND3_X1 U18066 ( .A1(n14847), .A2(n14692), .A3(n20081), .ZN(n14703) );
  OAI211_X1 U18067 ( .C1(n15715), .C2(n20142), .A(n14704), .B(n14703), .ZN(
        P1_U2981) );
  OAI21_X1 U18068 ( .B1(n14706), .B2(n14707), .A(n14718), .ZN(n15806) );
  INV_X1 U18069 ( .A(n14708), .ZN(n14709) );
  OAI21_X1 U18070 ( .B1(n15806), .B2(n14709), .A(n15802), .ZN(n14710) );
  XOR2_X1 U18071 ( .A(n14711), .B(n14710), .Z(n14864) );
  INV_X1 U18072 ( .A(n14712), .ZN(n14714) );
  AOI22_X1 U18073 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14713) );
  OAI21_X1 U18074 ( .B1(n20085), .B2(n14714), .A(n14713), .ZN(n14715) );
  AOI21_X1 U18075 ( .B1(n14716), .B2(n14666), .A(n14715), .ZN(n14717) );
  OAI21_X1 U18076 ( .B1(n14864), .B2(n19900), .A(n14717), .ZN(P1_U2983) );
  NAND2_X1 U18077 ( .A1(n14706), .A2(n14718), .ZN(n14722) );
  INV_X1 U18078 ( .A(n14719), .ZN(n14720) );
  AOI21_X1 U18079 ( .B1(n14722), .B2(n14721), .A(n14720), .ZN(n14724) );
  INV_X1 U18080 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14856) );
  MUX2_X1 U18081 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n14856), .S(
        n9738), .Z(n14723) );
  XNOR2_X1 U18082 ( .A(n14724), .B(n14723), .ZN(n14872) );
  NAND2_X1 U18083 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14725) );
  NAND2_X1 U18084 ( .A1(n13397), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n14866) );
  OAI211_X1 U18085 ( .C1(n20085), .C2(n15734), .A(n14725), .B(n14866), .ZN(
        n14726) );
  AOI21_X1 U18086 ( .B1(n15736), .B2(n14666), .A(n14726), .ZN(n14727) );
  OAI21_X1 U18087 ( .B1(n14872), .B2(n19900), .A(n14727), .ZN(P1_U2985) );
  INV_X1 U18088 ( .A(n14728), .ZN(n14729) );
  OR2_X1 U18089 ( .A1(n14706), .A2(n14729), .ZN(n14733) );
  INV_X1 U18090 ( .A(n14730), .ZN(n14731) );
  NAND2_X1 U18091 ( .A1(n15794), .A2(n14731), .ZN(n14732) );
  NAND2_X1 U18092 ( .A1(n14733), .A2(n14732), .ZN(n15816) );
  OAI21_X1 U18093 ( .B1(n9738), .B2(n14734), .A(n14735), .ZN(n15815) );
  NAND2_X1 U18094 ( .A1(n15813), .A2(n14735), .ZN(n14736) );
  XOR2_X1 U18095 ( .A(n14737), .B(n14736), .Z(n15896) );
  NAND2_X1 U18096 ( .A1(n15896), .A2(n20081), .ZN(n14742) );
  OAI22_X1 U18097 ( .A1(n15784), .A2(n14738), .B1(n20107), .B2(n20744), .ZN(
        n14739) );
  AOI21_X1 U18098 ( .B1(n15820), .B2(n14740), .A(n14739), .ZN(n14741) );
  OAI211_X1 U18099 ( .C1(n20142), .C2(n14743), .A(n14742), .B(n14741), .ZN(
        P1_U2986) );
  NAND2_X1 U18100 ( .A1(n14744), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14746) );
  XNOR2_X1 U18101 ( .A(n14706), .B(n14747), .ZN(n14745) );
  MUX2_X1 U18102 ( .A(n14746), .B(n14745), .S(n9738), .Z(n14749) );
  INV_X1 U18103 ( .A(n14744), .ZN(n14748) );
  NAND3_X1 U18104 ( .A1(n14748), .A2(n15794), .A3(n14747), .ZN(n15824) );
  NAND2_X1 U18105 ( .A1(n14749), .A2(n15824), .ZN(n15930) );
  INV_X1 U18106 ( .A(n15930), .ZN(n14755) );
  AOI22_X1 U18107 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n14750) );
  OAI21_X1 U18108 ( .B1(n20085), .B2(n14751), .A(n14750), .ZN(n14752) );
  AOI21_X1 U18109 ( .B1(n14753), .B2(n14666), .A(n14752), .ZN(n14754) );
  OAI21_X1 U18110 ( .B1(n14755), .B2(n19900), .A(n14754), .ZN(P1_U2989) );
  NOR2_X1 U18111 ( .A1(n14756), .A2(n20109), .ZN(n14776) );
  INV_X1 U18112 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15972) );
  NAND2_X1 U18113 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20089) );
  NOR2_X1 U18114 ( .A1(n15972), .A2(n20089), .ZN(n15906) );
  INV_X1 U18115 ( .A(n15906), .ZN(n14757) );
  AOI21_X1 U18116 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20111) );
  OR2_X1 U18117 ( .A1(n14757), .A2(n20111), .ZN(n15902) );
  INV_X1 U18118 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15959) );
  NOR3_X1 U18119 ( .A1(n13736), .A2(n15959), .A3(n15837), .ZN(n15926) );
  NAND3_X1 U18120 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n15926), .ZN(n15907) );
  NOR2_X1 U18121 ( .A1(n15902), .A2(n15907), .ZN(n15918) );
  NAND3_X1 U18122 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n15918), .ZN(n14762) );
  NOR2_X1 U18123 ( .A1(n20114), .A2(n14762), .ZN(n15627) );
  NAND2_X1 U18124 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14758) );
  INV_X1 U18125 ( .A(n15907), .ZN(n15901) );
  NOR3_X1 U18126 ( .A1(n20120), .A2(n20135), .A3(n14757), .ZN(n15923) );
  NAND2_X1 U18127 ( .A1(n15901), .A2(n15923), .ZN(n15905) );
  NOR2_X1 U18128 ( .A1(n14758), .A2(n15905), .ZN(n15890) );
  NAND2_X1 U18129 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15890), .ZN(
        n14763) );
  NAND2_X1 U18130 ( .A1(n15893), .A2(n15626), .ZN(n15947) );
  NAND2_X1 U18131 ( .A1(n20110), .A2(n15893), .ZN(n20122) );
  NAND2_X1 U18132 ( .A1(n15947), .A2(n20122), .ZN(n20103) );
  NOR2_X1 U18133 ( .A1(n14763), .A2(n20103), .ZN(n15852) );
  NAND3_X1 U18134 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15874) );
  NOR2_X1 U18135 ( .A1(n12801), .A2(n15874), .ZN(n14851) );
  NAND2_X1 U18136 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14851), .ZN(
        n14765) );
  NOR2_X1 U18137 ( .A1(n15875), .A2(n14765), .ZN(n15866) );
  NAND2_X1 U18138 ( .A1(n15866), .A2(n15629), .ZN(n14838) );
  NAND2_X1 U18139 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14844) );
  NAND2_X1 U18140 ( .A1(n14822), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14759) );
  NOR2_X1 U18141 ( .A1(n14819), .A2(n14759), .ZN(n14817) );
  NAND3_X1 U18142 ( .A1(n14817), .A2(n14796), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14784) );
  NOR3_X1 U18143 ( .A1(n14784), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14783), .ZN(n14775) );
  INV_X1 U18144 ( .A(n14760), .ZN(n14761) );
  NAND2_X1 U18145 ( .A1(n20086), .A2(n15864), .ZN(n14767) );
  OAI21_X1 U18146 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15626), .A(
        n20134), .ZN(n20104) );
  NOR2_X1 U18147 ( .A1(n20123), .A2(n20104), .ZN(n14766) );
  NOR2_X1 U18148 ( .A1(n15899), .A2(n14762), .ZN(n14869) );
  AOI21_X1 U18149 ( .B1(n15947), .B2(n14763), .A(n20104), .ZN(n14764) );
  OAI21_X1 U18150 ( .B1(n14869), .B2(n20114), .A(n14764), .ZN(n14865) );
  INV_X1 U18151 ( .A(n14766), .ZN(n15924) );
  OAI21_X1 U18152 ( .B1(n14865), .B2(n14765), .A(n15924), .ZN(n15872) );
  OAI21_X1 U18153 ( .B1(n15629), .B2(n14766), .A(n15872), .ZN(n15613) );
  AOI21_X1 U18154 ( .B1(n20123), .B2(n14844), .A(n15613), .ZN(n15865) );
  NAND2_X1 U18155 ( .A1(n14767), .A2(n15865), .ZN(n15850) );
  INV_X1 U18156 ( .A(n15850), .ZN(n14770) );
  INV_X1 U18157 ( .A(n14821), .ZN(n14768) );
  NAND2_X1 U18158 ( .A1(n15947), .A2(n14768), .ZN(n14769) );
  OAI211_X1 U18159 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n20114), .A(
        n14770), .B(n14769), .ZN(n14834) );
  NOR2_X1 U18160 ( .A1(n14834), .A2(n14824), .ZN(n14825) );
  INV_X1 U18161 ( .A(n14796), .ZN(n14804) );
  NOR2_X1 U18162 ( .A1(n14804), .A2(n14820), .ZN(n14771) );
  NOR2_X1 U18163 ( .A1(n14834), .A2(n20123), .ZN(n14772) );
  AOI21_X1 U18164 ( .B1(n14825), .B2(n14771), .A(n14772), .ZN(n14794) );
  AOI211_X1 U18165 ( .C1(n14795), .C2(n20123), .A(n14783), .B(n14794), .ZN(
        n14782) );
  NOR3_X1 U18166 ( .A1(n14782), .A2(n14772), .A3(n20879), .ZN(n14773) );
  NOR4_X1 U18167 ( .A1(n14776), .A2(n14775), .A3(n14774), .A4(n14773), .ZN(
        n14777) );
  OAI21_X1 U18168 ( .B1(n14778), .B2(n15913), .A(n14777), .ZN(P1_U3000) );
  INV_X1 U18169 ( .A(n14779), .ZN(n14789) );
  INV_X1 U18170 ( .A(n14780), .ZN(n14787) );
  INV_X1 U18171 ( .A(n14781), .ZN(n14786) );
  AOI21_X1 U18172 ( .B1(n14784), .B2(n14783), .A(n14782), .ZN(n14785) );
  AOI211_X1 U18173 ( .C1(n14787), .C2(n20126), .A(n14786), .B(n14785), .ZN(
        n14788) );
  OAI21_X1 U18174 ( .B1(n14789), .B2(n15913), .A(n14788), .ZN(P1_U3001) );
  INV_X1 U18175 ( .A(n14790), .ZN(n14791) );
  NOR2_X1 U18176 ( .A1(n14791), .A2(n20109), .ZN(n14792) );
  AOI211_X1 U18177 ( .C1(n14794), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14793), .B(n14792), .ZN(n14798) );
  NAND3_X1 U18178 ( .A1(n14817), .A2(n14796), .A3(n14795), .ZN(n14797) );
  OAI211_X1 U18179 ( .C1(n14799), .C2(n15913), .A(n14798), .B(n14797), .ZN(
        P1_U3002) );
  NAND2_X1 U18180 ( .A1(n14800), .A2(n20128), .ZN(n14809) );
  AND2_X1 U18181 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14801) );
  NOR2_X1 U18182 ( .A1(n14857), .A2(n14801), .ZN(n14802) );
  OR2_X1 U18183 ( .A1(n14834), .A2(n14802), .ZN(n14811) );
  AOI21_X1 U18184 ( .B1(n14811), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14803), .ZN(n14808) );
  NAND3_X1 U18185 ( .A1(n14817), .A2(n9872), .A3(n14804), .ZN(n14807) );
  NAND2_X1 U18186 ( .A1(n14805), .A2(n20126), .ZN(n14806) );
  NAND4_X1 U18187 ( .A1(n14809), .A2(n14808), .A3(n14807), .A4(n14806), .ZN(
        P1_U3003) );
  AOI21_X1 U18188 ( .B1(n14811), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14810), .ZN(n14812) );
  OAI21_X1 U18189 ( .B1(n14813), .B2(n20109), .A(n14812), .ZN(n14815) );
  INV_X1 U18190 ( .A(n15659), .ZN(n14828) );
  INV_X1 U18191 ( .A(n14818), .ZN(n14827) );
  NAND3_X1 U18192 ( .A1(n15859), .A2(n14821), .A3(n14820), .ZN(n14835) );
  NAND2_X1 U18193 ( .A1(n14822), .A2(n15859), .ZN(n14823) );
  AOI22_X1 U18194 ( .A1(n14825), .A2(n14835), .B1(n14824), .B2(n14823), .ZN(
        n14826) );
  AOI211_X1 U18195 ( .C1(n20126), .C2(n14828), .A(n14827), .B(n14826), .ZN(
        n14829) );
  OAI21_X1 U18196 ( .B1(n14830), .B2(n15913), .A(n14829), .ZN(P1_U3005) );
  INV_X1 U18197 ( .A(n14831), .ZN(n14837) );
  NOR2_X1 U18198 ( .A1(n15667), .A2(n20109), .ZN(n14832) );
  AOI211_X1 U18199 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n14834), .A(
        n14833), .B(n14832), .ZN(n14836) );
  OAI211_X1 U18200 ( .C1(n14837), .C2(n15913), .A(n14836), .B(n14835), .ZN(
        P1_U3006) );
  INV_X1 U18201 ( .A(n14838), .ZN(n15611) );
  OAI21_X1 U18202 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15611), .ZN(n14839) );
  INV_X1 U18203 ( .A(n14839), .ZN(n14843) );
  NAND2_X1 U18204 ( .A1(n15613), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14841) );
  OAI211_X1 U18205 ( .C1(n20109), .C2(n15690), .A(n14841), .B(n14840), .ZN(
        n14842) );
  AOI21_X1 U18206 ( .B1(n14844), .B2(n14843), .A(n14842), .ZN(n14845) );
  OAI21_X1 U18207 ( .B1(n14846), .B2(n15913), .A(n14845), .ZN(P1_U3009) );
  NAND3_X1 U18208 ( .A1(n14847), .A2(n14692), .A3(n20128), .ZN(n14854) );
  NOR2_X1 U18209 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15875), .ZN(
        n14852) );
  INV_X1 U18210 ( .A(n14865), .ZN(n15900) );
  OAI21_X1 U18211 ( .B1(n14857), .B2(n14851), .A(n15900), .ZN(n15878) );
  NAND2_X1 U18212 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15878), .ZN(
        n14848) );
  OAI211_X1 U18213 ( .C1(n15720), .C2(n20109), .A(n14849), .B(n14848), .ZN(
        n14850) );
  AOI21_X1 U18214 ( .B1(n14852), .B2(n14851), .A(n14850), .ZN(n14853) );
  NAND2_X1 U18215 ( .A1(n14854), .A2(n14853), .ZN(P1_U3013) );
  NOR4_X1 U18216 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15875), .A3(
        n14856), .A4(n14855), .ZN(n14862) );
  NOR3_X1 U18217 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15875), .A3(
        n14856), .ZN(n15886) );
  OAI21_X1 U18218 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14857), .A(
        n15900), .ZN(n15883) );
  OAI21_X1 U18219 ( .B1(n15886), .B2(n15883), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14859) );
  OR2_X1 U18220 ( .A1(n20107), .A2(n20748), .ZN(n14858) );
  OAI211_X1 U18221 ( .C1(n20109), .C2(n14860), .A(n14859), .B(n14858), .ZN(
        n14861) );
  NOR2_X1 U18222 ( .A1(n14862), .A2(n14861), .ZN(n14863) );
  OAI21_X1 U18223 ( .B1(n14864), .B2(n15913), .A(n14863), .ZN(P1_U3015) );
  NOR3_X1 U18224 ( .A1(n20120), .A2(n20135), .A3(n20103), .ZN(n15944) );
  NOR2_X1 U18225 ( .A1(n20086), .A2(n15944), .ZN(n15915) );
  NOR2_X1 U18226 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15915), .ZN(
        n14870) );
  NAND2_X1 U18227 ( .A1(n14865), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14867) );
  OAI211_X1 U18228 ( .C1(n20109), .C2(n15731), .A(n14867), .B(n14866), .ZN(
        n14868) );
  AOI21_X1 U18229 ( .B1(n14870), .B2(n14869), .A(n14868), .ZN(n14871) );
  OAI21_X1 U18230 ( .B1(n14872), .B2(n15913), .A(n14871), .ZN(P1_U3017) );
  NOR2_X1 U18231 ( .A1(n14873), .A2(n15981), .ZN(n15601) );
  INV_X1 U18232 ( .A(n15601), .ZN(n14876) );
  NAND2_X1 U18233 ( .A1(n20256), .A2(n14874), .ZN(n14875) );
  OAI211_X1 U18234 ( .C1(n20644), .C2(n20222), .A(n14876), .B(n14875), .ZN(
        n14877) );
  MUX2_X1 U18235 ( .A(n14877), .B(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .S(
        n20136), .Z(P1_U3478) );
  NOR2_X1 U18236 ( .A1(n14878), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14881) );
  NOR3_X1 U18237 ( .A1(n14879), .A2(n14884), .A3(n13361), .ZN(n14880) );
  AOI211_X1 U18238 ( .C1(n20598), .C2(n14882), .A(n14881), .B(n14880), .ZN(
        n15575) );
  INV_X1 U18239 ( .A(n14883), .ZN(n14887) );
  INV_X1 U18240 ( .A(n15602), .ZN(n14891) );
  NOR3_X1 U18241 ( .A1(n13361), .A2(n14884), .A3(n14891), .ZN(n14885) );
  AOI21_X1 U18242 ( .B1(n14887), .B2(n14886), .A(n14885), .ZN(n14888) );
  OAI21_X1 U18243 ( .B1(n15575), .B2(n14893), .A(n14888), .ZN(n14889) );
  MUX2_X1 U18244 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14889), .S(
        n14894), .Z(P1_U3473) );
  INV_X1 U18245 ( .A(n14890), .ZN(n14892) );
  OAI22_X1 U18246 ( .A1(n15582), .A2(n14893), .B1(n14892), .B2(n14891), .ZN(
        n14895) );
  MUX2_X1 U18247 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14895), .S(
        n14894), .Z(P1_U3469) );
  OAI21_X1 U18248 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n14896), .A(
        n15986), .ZN(n15153) );
  AOI21_X1 U18249 ( .B1(n16114), .B2(n14907), .A(n14896), .ZN(n16105) );
  INV_X1 U18250 ( .A(n16105), .ZN(n16068) );
  NAND2_X1 U18251 ( .A1(n15182), .A2(n14905), .ZN(n14898) );
  INV_X1 U18252 ( .A(n9831), .ZN(n14897) );
  AND2_X1 U18253 ( .A1(n14898), .A2(n14897), .ZN(n15184) );
  NOR2_X1 U18254 ( .A1(n14902), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14899) );
  NOR2_X1 U18255 ( .A1(n14906), .A2(n14899), .ZN(n18899) );
  AOI21_X1 U18256 ( .B1(n18924), .B2(n14900), .A(n14904), .ZN(n18923) );
  OAI21_X1 U18257 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n14901), .A(
        n14900), .ZN(n18935) );
  NAND2_X1 U18258 ( .A1(n18934), .A2(n18935), .ZN(n18921) );
  NOR2_X1 U18259 ( .A1(n18923), .A2(n18921), .ZN(n18909) );
  INV_X1 U18260 ( .A(n14902), .ZN(n14903) );
  OAI21_X1 U18261 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n14904), .A(
        n14903), .ZN(n18910) );
  NAND2_X1 U18262 ( .A1(n18909), .A2(n18910), .ZN(n18897) );
  NOR2_X1 U18263 ( .A1(n18899), .A2(n18897), .ZN(n14936) );
  OAI21_X1 U18264 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n14906), .A(
        n14905), .ZN(n15198) );
  OAI21_X1 U18265 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n9831), .A(
        n14907), .ZN(n15559) );
  NAND2_X1 U18266 ( .A1(n15560), .A2(n15559), .ZN(n15558) );
  NAND2_X1 U18267 ( .A1(n19032), .A2(n15558), .ZN(n16067) );
  NAND2_X1 U18268 ( .A1(n16068), .A2(n16067), .ZN(n16066) );
  NAND2_X1 U18269 ( .A1(n19032), .A2(n16066), .ZN(n14908) );
  NAND2_X1 U18270 ( .A1(n15153), .A2(n14908), .ZN(n15987) );
  OAI211_X1 U18271 ( .C1(n15153), .C2(n14908), .A(n19036), .B(n15987), .ZN(
        n14919) );
  AND2_X1 U18272 ( .A1(n14996), .A2(n14909), .ZN(n14910) );
  OR2_X1 U18273 ( .A1(n14910), .A2(n14981), .ZN(n15154) );
  OR2_X1 U18274 ( .A1(n15093), .A2(n14911), .ZN(n14912) );
  AND2_X1 U18275 ( .A1(n15082), .A2(n14912), .ZN(n16215) );
  INV_X1 U18276 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19800) );
  OAI22_X1 U18277 ( .A1(n19014), .A2(n11138), .B1(n19800), .B2(n19061), .ZN(
        n14915) );
  INV_X1 U18278 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14913) );
  NOR2_X1 U18279 ( .A1(n19072), .A2(n14913), .ZN(n14914) );
  AOI211_X1 U18280 ( .C1(n19042), .C2(n16215), .A(n14915), .B(n14914), .ZN(
        n14916) );
  OAI21_X1 U18281 ( .B1(n15154), .B2(n19047), .A(n14916), .ZN(n14917) );
  INV_X1 U18282 ( .A(n14917), .ZN(n14918) );
  OAI211_X1 U18283 ( .C1(n14920), .C2(n19067), .A(n14919), .B(n14918), .ZN(
        P2_U2831) );
  OAI21_X1 U18284 ( .B1(n14934), .B2(n14921), .A(n15342), .ZN(n15358) );
  OAI22_X1 U18285 ( .A1(n15182), .A2(n19072), .B1(n19794), .B2(n19061), .ZN(
        n14924) );
  INV_X1 U18286 ( .A(n14935), .ZN(n14922) );
  AOI221_X1 U18287 ( .B1(n15184), .B2(n14935), .C1(n10064), .C2(n14922), .A(
        n19741), .ZN(n14923) );
  AOI211_X1 U18288 ( .C1(P2_EBX_REG_21__SCAN_IN), .C2(n19065), .A(n14924), .B(
        n14923), .ZN(n14930) );
  AND2_X1 U18289 ( .A1(n14942), .A2(n14925), .ZN(n14926) );
  OR2_X1 U18290 ( .A1(n14926), .A2(n15003), .ZN(n15357) );
  OAI22_X1 U18291 ( .A1(n14927), .A2(n19067), .B1(n15357), .B2(n19047), .ZN(
        n14928) );
  INV_X1 U18292 ( .A(n14928), .ZN(n14929) );
  OAI211_X1 U18293 ( .C1(n15358), .C2(n19063), .A(n14930), .B(n14929), .ZN(
        P2_U2834) );
  NOR2_X1 U18294 ( .A1(n14932), .A2(n14931), .ZN(n14933) );
  OR2_X1 U18295 ( .A1(n14934), .A2(n14933), .ZN(n16086) );
  AOI22_X1 U18296 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(n19030), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n19065), .ZN(n14938) );
  OAI211_X1 U18297 ( .C1(n14936), .C2(n15198), .A(n19036), .B(n14935), .ZN(
        n14937) );
  OAI211_X1 U18298 ( .C1(n15198), .C2(n19071), .A(n14938), .B(n14937), .ZN(
        n14939) );
  AOI21_X1 U18299 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19043), .A(
        n14939), .ZN(n14946) );
  NAND2_X1 U18300 ( .A1(n15023), .A2(n14940), .ZN(n14941) );
  NAND2_X1 U18301 ( .A1(n14942), .A2(n14941), .ZN(n15368) );
  NOR2_X1 U18302 ( .A1(n15368), .A2(n19047), .ZN(n14943) );
  AOI21_X1 U18303 ( .B1(n14944), .B2(n19041), .A(n14943), .ZN(n14945) );
  OAI211_X1 U18304 ( .C1(n16086), .C2(n19063), .A(n14946), .B(n14945), .ZN(
        P2_U2835) );
  MUX2_X1 U18305 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n15993), .S(n14992), .Z(
        P2_U2856) );
  NAND2_X1 U18306 ( .A1(n14948), .A2(n14947), .ZN(n14949) );
  NAND2_X1 U18307 ( .A1(n14950), .A2(n14949), .ZN(n16012) );
  INV_X1 U18308 ( .A(n14951), .ZN(n15045) );
  NAND2_X1 U18309 ( .A1(n14953), .A2(n14952), .ZN(n15044) );
  NAND3_X1 U18310 ( .A1(n15045), .A2(n15007), .A3(n15044), .ZN(n14955) );
  NAND2_X1 U18311 ( .A1(n15040), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14954) );
  OAI211_X1 U18312 ( .C1(n15040), .C2(n16012), .A(n14955), .B(n14954), .ZN(
        P2_U2858) );
  NAND2_X1 U18313 ( .A1(n14957), .A2(n14956), .ZN(n14959) );
  XNOR2_X1 U18314 ( .A(n14959), .B(n14958), .ZN(n15064) );
  NOR2_X1 U18315 ( .A1(n15288), .A2(n15040), .ZN(n14960) );
  AOI21_X1 U18316 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15040), .A(n14960), .ZN(
        n14961) );
  OAI21_X1 U18317 ( .B1(n15064), .B2(n15026), .A(n14961), .ZN(P2_U2859) );
  AOI21_X1 U18318 ( .B1(n14964), .B2(n14963), .A(n14962), .ZN(n14965) );
  INV_X1 U18319 ( .A(n14965), .ZN(n15073) );
  XNOR2_X1 U18320 ( .A(n14966), .B(n14967), .ZN(n15296) );
  NOR2_X1 U18321 ( .A1(n15296), .A2(n15040), .ZN(n14968) );
  AOI21_X1 U18322 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n15040), .A(n14968), .ZN(
        n14969) );
  OAI21_X1 U18323 ( .B1(n15073), .B2(n15026), .A(n14969), .ZN(P2_U2860) );
  OAI21_X1 U18324 ( .B1(n14972), .B2(n14971), .A(n14970), .ZN(n15080) );
  OR2_X1 U18325 ( .A1(n14983), .A2(n14973), .ZN(n14974) );
  NAND2_X1 U18326 ( .A1(n14966), .A2(n14974), .ZN(n16045) );
  NOR2_X1 U18327 ( .A1(n16045), .A2(n15040), .ZN(n14975) );
  AOI21_X1 U18328 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n15040), .A(n14975), .ZN(
        n14976) );
  OAI21_X1 U18329 ( .B1(n15080), .B2(n15026), .A(n14976), .ZN(P2_U2861) );
  OAI21_X1 U18330 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n15090) );
  NOR2_X1 U18331 ( .A1(n14981), .A2(n14980), .ZN(n14982) );
  OR2_X1 U18332 ( .A1(n14983), .A2(n14982), .ZN(n16104) );
  MUX2_X1 U18333 ( .A(n16104), .B(n14984), .S(n15040), .Z(n14985) );
  OAI21_X1 U18334 ( .B1(n15090), .B2(n15026), .A(n14985), .ZN(P2_U2862) );
  AOI21_X1 U18335 ( .B1(n14987), .B2(n14986), .A(n9809), .ZN(n14989) );
  XNOR2_X1 U18336 ( .A(n14989), .B(n14988), .ZN(n16073) );
  NAND2_X1 U18337 ( .A1(n16073), .A2(n15007), .ZN(n14991) );
  INV_X1 U18338 ( .A(n15154), .ZN(n16216) );
  NAND2_X1 U18339 ( .A1(n16216), .A2(n14992), .ZN(n14990) );
  OAI211_X1 U18340 ( .C1(n14992), .C2(n11138), .A(n14991), .B(n14990), .ZN(
        P2_U2863) );
  NAND2_X1 U18341 ( .A1(n14993), .A2(n14994), .ZN(n14995) );
  NAND2_X1 U18342 ( .A1(n14996), .A2(n14995), .ZN(n16229) );
  AOI21_X1 U18343 ( .B1(n14999), .B2(n14998), .A(n14997), .ZN(n15098) );
  NAND2_X1 U18344 ( .A1(n15098), .A2(n15007), .ZN(n15001) );
  NAND2_X1 U18345 ( .A1(n15040), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15000) );
  OAI211_X1 U18346 ( .C1(n16229), .C2(n15040), .A(n15001), .B(n15000), .ZN(
        P2_U2864) );
  OAI21_X1 U18347 ( .B1(n15003), .B2(n15002), .A(n14993), .ZN(n15556) );
  AOI21_X1 U18348 ( .B1(n15006), .B2(n15011), .A(n15005), .ZN(n16080) );
  NAND2_X1 U18349 ( .A1(n16080), .A2(n15007), .ZN(n15009) );
  NAND2_X1 U18350 ( .A1(n15040), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n15008) );
  OAI211_X1 U18351 ( .C1(n15556), .C2(n15040), .A(n15009), .B(n15008), .ZN(
        P2_U2865) );
  OAI21_X1 U18352 ( .B1(n15010), .B2(n15012), .A(n15011), .ZN(n15105) );
  MUX2_X1 U18353 ( .A(n15357), .B(n15013), .S(n15040), .Z(n15014) );
  OAI21_X1 U18354 ( .B1(n15105), .B2(n15026), .A(n15014), .ZN(P2_U2866) );
  NAND2_X1 U18355 ( .A1(n15016), .A2(n15015), .ZN(n15017) );
  NAND2_X1 U18356 ( .A1(n10159), .A2(n15017), .ZN(n16085) );
  INV_X1 U18357 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n15018) );
  MUX2_X1 U18358 ( .A(n15368), .B(n15018), .S(n15040), .Z(n15019) );
  OAI21_X1 U18359 ( .B1(n16085), .B2(n15026), .A(n15019), .ZN(P2_U2867) );
  NAND2_X1 U18360 ( .A1(n15020), .A2(n15021), .ZN(n15022) );
  NAND2_X1 U18361 ( .A1(n15023), .A2(n15022), .ZN(n18903) );
  NOR2_X1 U18362 ( .A1(n18903), .A2(n15040), .ZN(n15024) );
  AOI21_X1 U18363 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15040), .A(n15024), .ZN(
        n15025) );
  OAI21_X1 U18364 ( .B1(n15027), .B2(n15026), .A(n15025), .ZN(P2_U2868) );
  OR2_X1 U18365 ( .A1(n15029), .A2(n15028), .ZN(n15030) );
  NAND2_X1 U18366 ( .A1(n15031), .A2(n15030), .ZN(n16091) );
  OR2_X1 U18367 ( .A1(n15038), .A2(n15032), .ZN(n15033) );
  NAND2_X1 U18368 ( .A1(n15020), .A2(n15033), .ZN(n18915) );
  INV_X1 U18369 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n15034) );
  MUX2_X1 U18370 ( .A(n18915), .B(n15034), .S(n15040), .Z(n15035) );
  OAI21_X1 U18371 ( .B1(n16091), .B2(n15026), .A(n15035), .ZN(P2_U2869) );
  AND2_X1 U18372 ( .A1(n15037), .A2(n15036), .ZN(n15039) );
  OR2_X1 U18373 ( .A1(n15039), .A2(n15038), .ZN(n18928) );
  MUX2_X1 U18374 ( .A(n18928), .B(n15041), .S(n15040), .Z(n15042) );
  OAI21_X1 U18375 ( .B1(n15043), .B2(n15026), .A(n15042), .ZN(P2_U2870) );
  NAND3_X1 U18376 ( .A1(n15045), .A2(n16079), .A3(n15044), .ZN(n15054) );
  AND2_X1 U18377 ( .A1(n15057), .A2(n15046), .ZN(n15047) );
  OAI22_X1 U18378 ( .A1(n16092), .A2(n15274), .B1(n19103), .B2(n15049), .ZN(
        n15050) );
  AOI21_X1 U18379 ( .B1(n19082), .B2(n15051), .A(n15050), .ZN(n15053) );
  AOI22_X1 U18380 ( .A1(n19083), .A2(BUF1_REG_29__SCAN_IN), .B1(n19084), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15052) );
  NAND3_X1 U18381 ( .A1(n15054), .A2(n15053), .A3(n15052), .ZN(P2_U2890) );
  NAND2_X1 U18382 ( .A1(n15067), .A2(n15055), .ZN(n15056) );
  INV_X1 U18383 ( .A(n19082), .ZN(n15060) );
  OAI22_X1 U18384 ( .A1(n15060), .A2(n15059), .B1(n19103), .B2(n15058), .ZN(
        n15061) );
  AOI21_X1 U18385 ( .B1(n19087), .B2(n16020), .A(n15061), .ZN(n15063) );
  AOI22_X1 U18386 ( .A1(n19083), .A2(BUF1_REG_28__SCAN_IN), .B1(n19084), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15062) );
  OAI211_X1 U18387 ( .C1(n15064), .C2(n19107), .A(n15063), .B(n15062), .ZN(
        P2_U2891) );
  OR2_X1 U18388 ( .A1(n15076), .A2(n15065), .ZN(n15066) );
  NAND2_X1 U18389 ( .A1(n15067), .A2(n15066), .ZN(n16040) );
  OAI22_X1 U18390 ( .A1(n16092), .A2(n16040), .B1(n19103), .B2(n15068), .ZN(
        n15069) );
  AOI21_X1 U18391 ( .B1(n19082), .B2(n15070), .A(n15069), .ZN(n15072) );
  AOI22_X1 U18392 ( .A1(n19083), .A2(BUF1_REG_27__SCAN_IN), .B1(n19084), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n15071) );
  OAI211_X1 U18393 ( .C1(n15073), .C2(n19107), .A(n15072), .B(n15071), .ZN(
        P2_U2892) );
  AND2_X1 U18394 ( .A1(n15084), .A2(n15074), .ZN(n15075) );
  NOR2_X1 U18395 ( .A1(n15076), .A2(n15075), .ZN(n15314) );
  INV_X1 U18396 ( .A(n15314), .ZN(n16044) );
  OAI22_X1 U18397 ( .A1(n16092), .A2(n16044), .B1(n19103), .B2(n13295), .ZN(
        n15077) );
  AOI21_X1 U18398 ( .B1(n19082), .B2(n19096), .A(n15077), .ZN(n15079) );
  AOI22_X1 U18399 ( .A1(n19083), .A2(BUF1_REG_26__SCAN_IN), .B1(n19084), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15078) );
  OAI211_X1 U18400 ( .C1(n15080), .C2(n19107), .A(n15079), .B(n15078), .ZN(
        P2_U2893) );
  NAND2_X1 U18401 ( .A1(n15082), .A2(n15081), .ZN(n15083) );
  NAND2_X1 U18402 ( .A1(n15084), .A2(n15083), .ZN(n16063) );
  OAI22_X1 U18403 ( .A1(n16092), .A2(n16063), .B1(n19103), .B2(n15085), .ZN(
        n15086) );
  AOI21_X1 U18404 ( .B1(n19082), .B2(n15087), .A(n15086), .ZN(n15089) );
  AOI22_X1 U18405 ( .A1(n19083), .A2(BUF1_REG_25__SCAN_IN), .B1(n19084), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n15088) );
  OAI211_X1 U18406 ( .C1(n15090), .C2(n19107), .A(n15089), .B(n15088), .ZN(
        P2_U2894) );
  NOR2_X1 U18407 ( .A1(n15091), .A2(n9830), .ZN(n15092) );
  OR2_X1 U18408 ( .A1(n15093), .A2(n15092), .ZN(n16222) );
  AOI22_X1 U18409 ( .A1(n19083), .A2(BUF1_REG_23__SCAN_IN), .B1(n19084), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n15096) );
  AOI22_X1 U18410 ( .A1(n19082), .A2(n15094), .B1(n19104), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n15095) );
  OAI211_X1 U18411 ( .C1(n16092), .C2(n16222), .A(n15096), .B(n15095), .ZN(
        n15097) );
  AOI21_X1 U18412 ( .B1(n15098), .B2(n16079), .A(n15097), .ZN(n15099) );
  INV_X1 U18413 ( .A(n15099), .ZN(P2_U2896) );
  NAND2_X1 U18414 ( .A1(n19083), .A2(BUF1_REG_21__SCAN_IN), .ZN(n15101) );
  AOI22_X1 U18415 ( .A1(n19082), .A2(n19105), .B1(n19104), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15100) );
  NAND2_X1 U18416 ( .A1(n15101), .A2(n15100), .ZN(n15103) );
  NOR2_X1 U18417 ( .A1(n15358), .A2(n16092), .ZN(n15102) );
  AOI211_X1 U18418 ( .C1(n19084), .C2(BUF2_REG_21__SCAN_IN), .A(n15103), .B(
        n15102), .ZN(n15104) );
  OAI21_X1 U18419 ( .B1(n19107), .B2(n15105), .A(n15104), .ZN(P2_U2898) );
  XNOR2_X1 U18420 ( .A(n15126), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15272) );
  NAND2_X1 U18421 ( .A1(n15106), .A2(n15117), .ZN(n15111) );
  INV_X1 U18422 ( .A(n15107), .ZN(n15109) );
  NAND2_X1 U18423 ( .A1(n15109), .A2(n15108), .ZN(n15110) );
  NAND2_X1 U18424 ( .A1(n15263), .A2(n19175), .ZN(n15116) );
  INV_X1 U18425 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15112) );
  NAND2_X1 U18426 ( .A1(n19029), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15265) );
  OAI21_X1 U18427 ( .B1(n16204), .B2(n15112), .A(n15265), .ZN(n15114) );
  XNOR2_X1 U18428 ( .A(n15121), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16002) );
  NOR2_X1 U18429 ( .A1(n16002), .A2(n19167), .ZN(n15113) );
  AOI211_X1 U18430 ( .C1(n19171), .C2(n15999), .A(n15114), .B(n15113), .ZN(
        n15115) );
  OAI211_X1 U18431 ( .C1(n19177), .C2(n15272), .A(n15116), .B(n15115), .ZN(
        P2_U2984) );
  NAND2_X1 U18432 ( .A1(n15118), .A2(n15117), .ZN(n15120) );
  XOR2_X1 U18433 ( .A(n15120), .B(n15119), .Z(n15284) );
  AOI21_X1 U18434 ( .B1(n15123), .B2(n15122), .A(n15121), .ZN(n15983) );
  NAND2_X1 U18435 ( .A1(n19029), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15273) );
  OAI21_X1 U18436 ( .B1(n16204), .B2(n15123), .A(n15273), .ZN(n15125) );
  NOR2_X1 U18437 ( .A1(n16012), .A2(n16158), .ZN(n15124) );
  AOI211_X1 U18438 ( .C1(n15983), .C2(n16198), .A(n15125), .B(n15124), .ZN(
        n15129) );
  AOI21_X1 U18439 ( .B1(n15136), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U18440 ( .A1(n15127), .A2(n15126), .ZN(n15282) );
  NAND2_X1 U18441 ( .A1(n15282), .A2(n16200), .ZN(n15128) );
  OAI211_X1 U18442 ( .C1(n15284), .C2(n19161), .A(n15129), .B(n15128), .ZN(
        P2_U2985) );
  XNOR2_X1 U18443 ( .A(n15130), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15310) );
  INV_X1 U18444 ( .A(n15131), .ZN(n15132) );
  AOI21_X1 U18445 ( .B1(n15133), .B2(n15144), .A(n15132), .ZN(n15984) );
  NAND2_X1 U18446 ( .A1(n19029), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15297) );
  OAI21_X1 U18447 ( .B1(n16204), .B2(n15133), .A(n15297), .ZN(n15135) );
  NOR2_X1 U18448 ( .A1(n15296), .A2(n16158), .ZN(n15134) );
  AOI211_X1 U18449 ( .C1(n16198), .C2(n15984), .A(n15135), .B(n15134), .ZN(
        n15138) );
  INV_X1 U18450 ( .A(n15136), .ZN(n15308) );
  NAND2_X1 U18451 ( .A1(n15142), .A2(n15301), .ZN(n15295) );
  NAND3_X1 U18452 ( .A1(n15308), .A2(n16200), .A3(n15295), .ZN(n15137) );
  OAI211_X1 U18453 ( .C1(n15310), .C2(n19161), .A(n15138), .B(n15137), .ZN(
        P2_U2987) );
  AOI21_X1 U18454 ( .B1(n15326), .B2(n15322), .A(n15323), .ZN(n15140) );
  MUX2_X1 U18455 ( .A(n15322), .B(n15140), .S(n15139), .Z(n15141) );
  NAND2_X1 U18456 ( .A1(n14039), .A2(n15141), .ZN(n15321) );
  INV_X1 U18457 ( .A(n15142), .ZN(n15143) );
  AOI21_X1 U18458 ( .B1(n15317), .B2(n15329), .A(n15143), .ZN(n15319) );
  OAI21_X1 U18459 ( .B1(n15985), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15144), .ZN(n16049) );
  AND2_X1 U18460 ( .A1(n19029), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15313) );
  NOR2_X1 U18461 ( .A1(n16045), .A2(n16158), .ZN(n15145) );
  AOI211_X1 U18462 ( .C1(n19169), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15313), .B(n15145), .ZN(n15146) );
  OAI21_X1 U18463 ( .B1(n19167), .B2(n16049), .A(n15146), .ZN(n15147) );
  AOI21_X1 U18464 ( .B1(n15319), .B2(n16200), .A(n15147), .ZN(n15148) );
  OAI21_X1 U18465 ( .B1(n15321), .B2(n19161), .A(n15148), .ZN(P2_U2988) );
  NAND2_X1 U18466 ( .A1(n15150), .A2(n15149), .ZN(n15151) );
  XOR2_X1 U18467 ( .A(n15152), .B(n15151), .Z(n16220) );
  AOI21_X1 U18468 ( .B1(n16210), .B2(n16109), .A(n15327), .ZN(n16217) );
  OAI22_X1 U18469 ( .A1(n19800), .A2(n19045), .B1(n19167), .B2(n15153), .ZN(
        n15156) );
  OAI22_X1 U18470 ( .A1(n15154), .A2(n16158), .B1(n14913), .B2(n16204), .ZN(
        n15155) );
  AOI211_X1 U18471 ( .C1(n16217), .C2(n16200), .A(n15156), .B(n15155), .ZN(
        n15157) );
  OAI21_X1 U18472 ( .B1(n16220), .B2(n19161), .A(n15157), .ZN(P2_U2990) );
  NAND2_X1 U18473 ( .A1(n15159), .A2(n15158), .ZN(n15161) );
  XOR2_X1 U18474 ( .A(n15161), .B(n15160), .Z(n15352) );
  NOR2_X1 U18475 ( .A1(n15556), .A2(n16158), .ZN(n15163) );
  INV_X1 U18476 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19796) );
  OAI22_X1 U18477 ( .A1(n19796), .A2(n19045), .B1(n19167), .B2(n15559), .ZN(
        n15162) );
  AOI211_X1 U18478 ( .C1(n19169), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15163), .B(n15162), .ZN(n15168) );
  NAND2_X1 U18479 ( .A1(n15464), .A2(n15164), .ZN(n15194) );
  NOR2_X1 U18480 ( .A1(n15194), .A2(n15181), .ZN(n15180) );
  INV_X1 U18481 ( .A(n15180), .ZN(n15166) );
  NOR2_X1 U18482 ( .A1(n15166), .A2(n15165), .ZN(n16110) );
  INV_X1 U18483 ( .A(n16110), .ZN(n15349) );
  NAND2_X1 U18484 ( .A1(n15166), .A2(n15165), .ZN(n15348) );
  NAND3_X1 U18485 ( .A1(n15349), .A2(n16200), .A3(n15348), .ZN(n15167) );
  OAI211_X1 U18486 ( .C1(n15352), .C2(n19161), .A(n15168), .B(n15167), .ZN(
        P2_U2992) );
  INV_X1 U18487 ( .A(n15171), .ZN(n15173) );
  NAND2_X1 U18488 ( .A1(n15176), .A2(n15175), .ZN(n15225) );
  INV_X1 U18489 ( .A(n15190), .ZN(n15177) );
  NAND2_X1 U18490 ( .A1(n15177), .A2(n15189), .ZN(n15178) );
  AOI21_X1 U18491 ( .B1(n15181), .B2(n15194), .A(n15180), .ZN(n15361) );
  NAND2_X1 U18492 ( .A1(n19029), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15355) );
  OAI21_X1 U18493 ( .B1(n16204), .B2(n15182), .A(n15355), .ZN(n15183) );
  AOI21_X1 U18494 ( .B1(n16198), .B2(n15184), .A(n15183), .ZN(n15185) );
  OAI21_X1 U18495 ( .B1(n15357), .B2(n16158), .A(n15185), .ZN(n15186) );
  AOI21_X1 U18496 ( .B1(n15361), .B2(n16200), .A(n15186), .ZN(n15187) );
  OAI21_X1 U18497 ( .B1(n15363), .B2(n19161), .A(n15187), .ZN(P2_U2993) );
  NAND2_X1 U18498 ( .A1(n15189), .A2(n15188), .ZN(n15193) );
  XOR2_X1 U18499 ( .A(n15193), .B(n15192), .Z(n15377) );
  AND2_X1 U18500 ( .A1(n15464), .A2(n15369), .ZN(n15219) );
  NAND2_X1 U18501 ( .A1(n15219), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15207) );
  INV_X1 U18502 ( .A(n15194), .ZN(n15195) );
  AOI21_X1 U18503 ( .B1(n15207), .B2(n15196), .A(n15195), .ZN(n15375) );
  NOR2_X1 U18504 ( .A1(n15368), .A2(n16158), .ZN(n15200) );
  NAND2_X1 U18505 ( .A1(n19029), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15367) );
  NAND2_X1 U18506 ( .A1(n19169), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15197) );
  OAI211_X1 U18507 ( .C1(n19167), .C2(n15198), .A(n15367), .B(n15197), .ZN(
        n15199) );
  AOI211_X1 U18508 ( .C1(n15375), .C2(n16200), .A(n15200), .B(n15199), .ZN(
        n15201) );
  OAI21_X1 U18509 ( .B1(n15377), .B2(n19161), .A(n15201), .ZN(P2_U2994) );
  NAND2_X1 U18510 ( .A1(n9728), .A2(n15203), .ZN(n15206) );
  NAND2_X1 U18511 ( .A1(n15204), .A2(n15215), .ZN(n15205) );
  XOR2_X1 U18512 ( .A(n15206), .B(n15205), .Z(n15378) );
  OAI21_X1 U18513 ( .B1(n15219), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15207), .ZN(n15387) );
  INV_X1 U18514 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15208) );
  NAND2_X1 U18515 ( .A1(n19029), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15379) );
  OAI21_X1 U18516 ( .B1(n16204), .B2(n15208), .A(n15379), .ZN(n15209) );
  AOI21_X1 U18517 ( .B1(n18899), .B2(n16198), .A(n15209), .ZN(n15211) );
  OR2_X1 U18518 ( .A1(n18903), .A2(n16158), .ZN(n15210) );
  OAI211_X1 U18519 ( .C1(n15387), .C2(n19177), .A(n15211), .B(n15210), .ZN(
        n15212) );
  AOI21_X1 U18520 ( .B1(n15378), .B2(n19175), .A(n15212), .ZN(n15213) );
  INV_X1 U18521 ( .A(n15213), .ZN(P2_U2995) );
  NAND2_X1 U18522 ( .A1(n15215), .A2(n15214), .ZN(n15216) );
  XNOR2_X1 U18523 ( .A(n15217), .B(n15216), .ZN(n15401) );
  INV_X1 U18524 ( .A(n15218), .ZN(n15395) );
  NAND2_X1 U18525 ( .A1(n15464), .A2(n15395), .ZN(n15228) );
  AOI21_X1 U18526 ( .B1(n21055), .B2(n15228), .A(n15219), .ZN(n15399) );
  AND2_X1 U18527 ( .A1(n19029), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15393) );
  NOR2_X1 U18528 ( .A1(n18910), .A2(n19167), .ZN(n15220) );
  AOI211_X1 U18529 ( .C1(n19169), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15393), .B(n15220), .ZN(n15221) );
  OAI21_X1 U18530 ( .B1(n16158), .B2(n18915), .A(n15221), .ZN(n15222) );
  AOI21_X1 U18531 ( .B1(n15399), .B2(n16200), .A(n15222), .ZN(n15223) );
  OAI21_X1 U18532 ( .B1(n15401), .B2(n19161), .A(n15223), .ZN(P2_U2996) );
  XOR2_X1 U18533 ( .A(n15225), .B(n15224), .Z(n15411) );
  AOI22_X1 U18534 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19169), .B1(
        n16198), .B2(n18923), .ZN(n15226) );
  NAND2_X1 U18535 ( .A1(n19029), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15405) );
  OAI211_X1 U18536 ( .C1(n16158), .C2(n18928), .A(n15226), .B(n15405), .ZN(
        n15227) );
  INV_X1 U18537 ( .A(n15227), .ZN(n15230) );
  OAI211_X1 U18538 ( .C1(n15235), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16200), .B(n15228), .ZN(n15229) );
  OAI211_X1 U18539 ( .C1(n15411), .C2(n19161), .A(n15230), .B(n15229), .ZN(
        P2_U2997) );
  INV_X1 U18540 ( .A(n15231), .ZN(n15241) );
  INV_X1 U18541 ( .A(n18942), .ZN(n15234) );
  NOR2_X1 U18542 ( .A1(n19785), .A2(n19045), .ZN(n15233) );
  INV_X1 U18543 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18938) );
  OAI22_X1 U18544 ( .A1(n18938), .A2(n16204), .B1(n19167), .B2(n18935), .ZN(
        n15232) );
  AOI211_X1 U18545 ( .C1(n15234), .C2(n19171), .A(n15233), .B(n15232), .ZN(
        n15240) );
  OAI21_X1 U18546 ( .B1(n16122), .B2(n15237), .A(n15236), .ZN(n15238) );
  NAND3_X1 U18547 ( .A1(n10166), .A2(n16200), .A3(n15238), .ZN(n15239) );
  OAI211_X1 U18548 ( .C1(n15241), .C2(n19161), .A(n15240), .B(n15239), .ZN(
        P2_U2998) );
  INV_X1 U18549 ( .A(n15242), .ZN(n15244) );
  NOR2_X1 U18550 ( .A1(n15244), .A2(n15243), .ZN(n15245) );
  XNOR2_X1 U18551 ( .A(n15246), .B(n15245), .ZN(n15482) );
  NAND2_X1 U18552 ( .A1(n16188), .A2(n16190), .ZN(n15247) );
  XNOR2_X1 U18553 ( .A(n16191), .B(n15247), .ZN(n15480) );
  OAI22_X1 U18554 ( .A1(n15248), .A2(n16204), .B1(n19771), .B2(n19045), .ZN(
        n15252) );
  INV_X1 U18555 ( .A(n15249), .ZN(n15250) );
  OAI22_X1 U18556 ( .A1(n19167), .A2(n15250), .B1(n16158), .B2(n15476), .ZN(
        n15251) );
  AOI211_X1 U18557 ( .C1(n15480), .C2(n19175), .A(n15252), .B(n15251), .ZN(
        n15253) );
  OAI21_X1 U18558 ( .B1(n15482), .B2(n19177), .A(n15253), .ZN(P2_U3007) );
  XNOR2_X1 U18559 ( .A(n15254), .B(n15255), .ZN(n15494) );
  OAI21_X1 U18560 ( .B1(n15257), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15256), .ZN(n15258) );
  INV_X1 U18561 ( .A(n15258), .ZN(n15492) );
  OAI22_X1 U18562 ( .A1(n19769), .A2(n19045), .B1(n19167), .B2(n19019), .ZN(
        n15261) );
  OAI22_X1 U18563 ( .A1(n16158), .A2(n15259), .B1(n16204), .B2(n10069), .ZN(
        n15260) );
  AOI211_X1 U18564 ( .C1(n15492), .C2(n16200), .A(n15261), .B(n15260), .ZN(
        n15262) );
  OAI21_X1 U18565 ( .B1(n19161), .B2(n15494), .A(n15262), .ZN(P2_U3008) );
  NAND2_X1 U18566 ( .A1(n15263), .A2(n19187), .ZN(n15271) );
  NAND2_X1 U18567 ( .A1(n15264), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15266) );
  OAI211_X1 U18568 ( .C1(n16289), .C2(n15997), .A(n15266), .B(n15265), .ZN(
        n15269) );
  NOR3_X1 U18569 ( .A1(n15305), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n15267), .ZN(n15268) );
  AOI211_X1 U18570 ( .C1(n19192), .C2(n15999), .A(n15269), .B(n15268), .ZN(
        n15270) );
  OAI211_X1 U18571 ( .C1(n15272), .C2(n19196), .A(n15271), .B(n15270), .ZN(
        P2_U3016) );
  OAI21_X1 U18572 ( .B1(n16289), .B2(n15274), .A(n15273), .ZN(n15275) );
  INV_X1 U18573 ( .A(n15275), .ZN(n15277) );
  INV_X1 U18574 ( .A(n15278), .ZN(n15280) );
  NOR3_X1 U18575 ( .A1(n15305), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15301), .ZN(n15289) );
  OAI21_X1 U18576 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16309), .A(
        n15302), .ZN(n15291) );
  OAI21_X1 U18577 ( .B1(n15289), .B2(n15291), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15279) );
  NAND2_X1 U18578 ( .A1(n15280), .A2(n15279), .ZN(n15281) );
  AOI21_X1 U18579 ( .B1(n15282), .B2(n16281), .A(n15281), .ZN(n15283) );
  OAI21_X1 U18580 ( .B1(n15284), .B2(n16305), .A(n15283), .ZN(P2_U3017) );
  NAND2_X1 U18581 ( .A1(n15285), .A2(n19187), .ZN(n15293) );
  NAND2_X1 U18582 ( .A1(n19186), .A2(n16020), .ZN(n15286) );
  OAI211_X1 U18583 ( .C1(n15288), .C2(n16266), .A(n15287), .B(n15286), .ZN(
        n15290) );
  AOI211_X1 U18584 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15291), .A(
        n15290), .B(n15289), .ZN(n15292) );
  OAI211_X1 U18585 ( .C1(n15294), .C2(n19196), .A(n15293), .B(n15292), .ZN(
        P2_U3018) );
  AND2_X1 U18586 ( .A1(n15295), .A2(n16281), .ZN(n15307) );
  INV_X1 U18587 ( .A(n15296), .ZN(n16034) );
  INV_X1 U18588 ( .A(n16040), .ZN(n15299) );
  INV_X1 U18589 ( .A(n15297), .ZN(n15298) );
  AOI21_X1 U18590 ( .B1(n19186), .B2(n15299), .A(n15298), .ZN(n15300) );
  OAI21_X1 U18591 ( .B1(n15302), .B2(n15301), .A(n15300), .ZN(n15303) );
  AOI21_X1 U18592 ( .B1(n16034), .B2(n19192), .A(n15303), .ZN(n15304) );
  OAI21_X1 U18593 ( .B1(n15305), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15304), .ZN(n15306) );
  AOI21_X1 U18594 ( .B1(n15308), .B2(n15307), .A(n15306), .ZN(n15309) );
  OAI21_X1 U18595 ( .B1(n15310), .B2(n16305), .A(n15309), .ZN(P2_U3019) );
  XNOR2_X1 U18596 ( .A(n15317), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15311) );
  NAND2_X1 U18597 ( .A1(n15330), .A2(n15311), .ZN(n15316) );
  NOR2_X1 U18598 ( .A1(n16045), .A2(n16266), .ZN(n15312) );
  AOI211_X1 U18599 ( .C1(n19186), .C2(n15314), .A(n15313), .B(n15312), .ZN(
        n15315) );
  OAI211_X1 U18600 ( .C1(n15336), .C2(n15317), .A(n15316), .B(n15315), .ZN(
        n15318) );
  AOI21_X1 U18601 ( .B1(n15319), .B2(n16281), .A(n15318), .ZN(n15320) );
  OAI21_X1 U18602 ( .B1(n15321), .B2(n16305), .A(n15320), .ZN(P2_U3020) );
  INV_X1 U18603 ( .A(n15322), .ZN(n15324) );
  NOR2_X1 U18604 ( .A1(n15324), .A2(n15323), .ZN(n15325) );
  XNOR2_X1 U18605 ( .A(n15326), .B(n15325), .ZN(n16101) );
  INV_X1 U18606 ( .A(n16101), .ZN(n15339) );
  OR2_X1 U18607 ( .A1(n15327), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15328) );
  AND2_X1 U18608 ( .A1(n15329), .A2(n15328), .ZN(n16100) );
  NAND2_X1 U18609 ( .A1(n15330), .A2(n15335), .ZN(n15334) );
  INV_X1 U18610 ( .A(n16104), .ZN(n15332) );
  INV_X1 U18611 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19802) );
  OAI22_X1 U18612 ( .A1(n16289), .A2(n16063), .B1(n19802), .B2(n19045), .ZN(
        n15331) );
  AOI21_X1 U18613 ( .B1(n15332), .B2(n19192), .A(n15331), .ZN(n15333) );
  OAI211_X1 U18614 ( .C1(n15336), .C2(n15335), .A(n15334), .B(n15333), .ZN(
        n15337) );
  AOI21_X1 U18615 ( .B1(n16100), .B2(n16281), .A(n15337), .ZN(n15338) );
  OAI21_X1 U18616 ( .B1(n15339), .B2(n16305), .A(n15338), .ZN(P2_U3021) );
  NAND2_X1 U18617 ( .A1(n15365), .A2(n15340), .ZN(n15341) );
  OAI211_X1 U18618 ( .C1(n15353), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15465), .B(n15341), .ZN(n16227) );
  NAND2_X1 U18619 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19029), .ZN(n15345) );
  AOI21_X1 U18620 ( .B1(n15343), .B2(n15342), .A(n9830), .ZN(n16078) );
  NAND2_X1 U18621 ( .A1(n19186), .A2(n16078), .ZN(n15344) );
  OAI211_X1 U18622 ( .C1(n15556), .C2(n16266), .A(n15345), .B(n15344), .ZN(
        n15347) );
  NOR2_X1 U18623 ( .A1(n16224), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15346) );
  AOI211_X1 U18624 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n16227), .A(
        n15347), .B(n15346), .ZN(n15351) );
  NAND3_X1 U18625 ( .A1(n15349), .A2(n16281), .A3(n15348), .ZN(n15350) );
  OAI211_X1 U18626 ( .C1(n15352), .C2(n16305), .A(n15351), .B(n15350), .ZN(
        P2_U3024) );
  INV_X1 U18627 ( .A(n15353), .ZN(n15354) );
  OAI21_X1 U18628 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n15354), .A(
        n16227), .ZN(n15356) );
  OAI211_X1 U18629 ( .C1(n15357), .C2(n16266), .A(n15356), .B(n15355), .ZN(
        n15360) );
  NOR2_X1 U18630 ( .A1(n15358), .A2(n16289), .ZN(n15359) );
  AOI211_X1 U18631 ( .C1(n15361), .C2(n16281), .A(n15360), .B(n15359), .ZN(
        n15362) );
  OAI21_X1 U18632 ( .B1(n15363), .B2(n16305), .A(n15362), .ZN(P2_U3025) );
  INV_X1 U18633 ( .A(n15369), .ZN(n15364) );
  NAND2_X1 U18634 ( .A1(n15365), .A2(n15364), .ZN(n15366) );
  NAND2_X1 U18635 ( .A1(n15465), .A2(n15366), .ZN(n15381) );
  OAI21_X1 U18636 ( .B1(n15368), .B2(n16266), .A(n15367), .ZN(n15372) );
  NAND2_X1 U18637 ( .A1(n15369), .A2(n15471), .ZN(n15383) );
  XNOR2_X1 U18638 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15370) );
  NOR2_X1 U18639 ( .A1(n15383), .A2(n15370), .ZN(n15371) );
  AOI211_X1 U18640 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15381), .A(
        n15372), .B(n15371), .ZN(n15373) );
  OAI21_X1 U18641 ( .B1(n16086), .B2(n16289), .A(n15373), .ZN(n15374) );
  AOI21_X1 U18642 ( .B1(n15375), .B2(n16281), .A(n15374), .ZN(n15376) );
  OAI21_X1 U18643 ( .B1(n15377), .B2(n16305), .A(n15376), .ZN(P2_U3026) );
  NAND2_X1 U18644 ( .A1(n15378), .A2(n19187), .ZN(n15386) );
  OAI21_X1 U18645 ( .B1(n18903), .B2(n16266), .A(n15379), .ZN(n15380) );
  AOI21_X1 U18646 ( .B1(n15381), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15380), .ZN(n15382) );
  OAI21_X1 U18647 ( .B1(n15383), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15382), .ZN(n15384) );
  AOI21_X1 U18648 ( .B1(n18905), .B2(n19186), .A(n15384), .ZN(n15385) );
  OAI211_X1 U18649 ( .C1(n15387), .C2(n19196), .A(n15386), .B(n15385), .ZN(
        P2_U3027) );
  NAND2_X1 U18650 ( .A1(n15389), .A2(n15388), .ZN(n15390) );
  NAND2_X1 U18651 ( .A1(n15391), .A2(n15390), .ZN(n18916) );
  OAI21_X1 U18652 ( .B1(n16309), .B2(n15395), .A(n15465), .ZN(n15394) );
  NOR2_X1 U18653 ( .A1(n18915), .A2(n16266), .ZN(n15392) );
  AOI211_X1 U18654 ( .C1(n15394), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15393), .B(n15392), .ZN(n15397) );
  NAND3_X1 U18655 ( .A1(n15471), .A2(n15395), .A3(n21055), .ZN(n15396) );
  OAI211_X1 U18656 ( .C1(n18916), .C2(n16289), .A(n15397), .B(n15396), .ZN(
        n15398) );
  AOI21_X1 U18657 ( .B1(n15399), .B2(n16281), .A(n15398), .ZN(n15400) );
  OAI21_X1 U18658 ( .B1(n15401), .B2(n16305), .A(n15400), .ZN(P2_U3028) );
  OAI21_X1 U18659 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16309), .A(
        n15402), .ZN(n15409) );
  NOR3_X1 U18660 ( .A1(n15404), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15403), .ZN(n15408) );
  NAND2_X1 U18661 ( .A1(n18930), .A2(n19186), .ZN(n15406) );
  OAI211_X1 U18662 ( .C1(n16266), .C2(n18928), .A(n15406), .B(n15405), .ZN(
        n15407) );
  AOI211_X1 U18663 ( .C1(n15409), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15408), .B(n15407), .ZN(n15410) );
  OAI21_X1 U18664 ( .B1(n15411), .B2(n16305), .A(n15410), .ZN(P2_U3029) );
  NAND2_X1 U18665 ( .A1(n15436), .A2(n15426), .ZN(n15412) );
  NAND2_X1 U18666 ( .A1(n16129), .A2(n15412), .ZN(n16141) );
  INV_X1 U18667 ( .A(n15413), .ZN(n15414) );
  NAND2_X1 U18668 ( .A1(n15415), .A2(n15414), .ZN(n15435) );
  INV_X1 U18669 ( .A(n15416), .ZN(n15432) );
  OAI21_X1 U18670 ( .B1(n15435), .B2(n15432), .A(n15417), .ZN(n15421) );
  AND2_X1 U18671 ( .A1(n15419), .A2(n15418), .ZN(n15420) );
  XNOR2_X1 U18672 ( .A(n15421), .B(n15420), .ZN(n16139) );
  NAND2_X1 U18673 ( .A1(n16139), .A2(n19187), .ZN(n15431) );
  OAI22_X1 U18674 ( .A1(n16266), .A2(n16140), .B1(n19779), .B2(n19045), .ZN(
        n15428) );
  NOR2_X1 U18675 ( .A1(n15470), .A2(n16249), .ZN(n16260) );
  NAND2_X1 U18676 ( .A1(n15422), .A2(n16260), .ZN(n15424) );
  NOR2_X1 U18677 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15424), .ZN(
        n15438) );
  NOR2_X1 U18678 ( .A1(n15470), .A2(n16261), .ZN(n15423) );
  OAI21_X1 U18679 ( .B1(n15423), .B2(n16309), .A(n15465), .ZN(n15439) );
  NOR2_X1 U18680 ( .A1(n15438), .A2(n15439), .ZN(n16253) );
  OR2_X1 U18681 ( .A1(n15424), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16252) );
  OAI22_X1 U18682 ( .A1(n16253), .A2(n15426), .B1(n15425), .B2(n16252), .ZN(
        n15427) );
  AOI211_X1 U18683 ( .C1(n19186), .C2(n15429), .A(n15428), .B(n15427), .ZN(
        n15430) );
  OAI211_X1 U18684 ( .C1(n16141), .C2(n19196), .A(n15431), .B(n15430), .ZN(
        P2_U3033) );
  NOR2_X1 U18685 ( .A1(n15433), .A2(n15432), .ZN(n15434) );
  XNOR2_X1 U18686 ( .A(n15435), .B(n15434), .ZN(n16148) );
  OAI21_X1 U18687 ( .B1(n16156), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15436), .ZN(n16147) );
  INV_X1 U18688 ( .A(n16147), .ZN(n15443) );
  NOR2_X1 U18689 ( .A1(n11549), .A2(n19045), .ZN(n15437) );
  AOI211_X1 U18690 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15439), .A(
        n15438), .B(n15437), .ZN(n15441) );
  NAND2_X1 U18691 ( .A1(n19192), .A2(n18964), .ZN(n15440) );
  OAI211_X1 U18692 ( .C1(n16289), .C2(n18968), .A(n15441), .B(n15440), .ZN(
        n15442) );
  AOI21_X1 U18693 ( .B1(n15443), .B2(n16281), .A(n15442), .ZN(n15444) );
  OAI21_X1 U18694 ( .B1(n16148), .B2(n16305), .A(n15444), .ZN(P2_U3034) );
  XNOR2_X1 U18695 ( .A(n16154), .B(n16153), .ZN(n16171) );
  NOR2_X1 U18696 ( .A1(n15458), .A2(n15462), .ZN(n15449) );
  INV_X1 U18697 ( .A(n15445), .ZN(n15446) );
  NAND2_X1 U18698 ( .A1(n15447), .A2(n15446), .ZN(n15448) );
  XNOR2_X1 U18699 ( .A(n15449), .B(n15448), .ZN(n16172) );
  INV_X1 U18700 ( .A(n16172), .ZN(n15456) );
  XNOR2_X1 U18701 ( .A(n15451), .B(n15450), .ZN(n19098) );
  OAI21_X1 U18702 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16309), .A(
        n15465), .ZN(n16265) );
  NOR2_X1 U18703 ( .A1(n11508), .A2(n19045), .ZN(n15452) );
  AOI221_X1 U18704 ( .B1(n16260), .B2(n16153), .C1(n16265), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n15452), .ZN(n15454) );
  NAND2_X1 U18705 ( .A1(n18989), .A2(n19192), .ZN(n15453) );
  OAI211_X1 U18706 ( .C1(n16289), .C2(n19098), .A(n15454), .B(n15453), .ZN(
        n15455) );
  AOI21_X1 U18707 ( .B1(n15456), .B2(n19187), .A(n15455), .ZN(n15457) );
  OAI21_X1 U18708 ( .B1(n19196), .B2(n16171), .A(n15457), .ZN(P2_U3036) );
  INV_X1 U18709 ( .A(n15458), .ZN(n15463) );
  OAI21_X1 U18710 ( .B1(n15460), .B2(n15462), .A(n15459), .ZN(n15461) );
  OAI21_X1 U18711 ( .B1(n15463), .B2(n15462), .A(n15461), .ZN(n16176) );
  INV_X1 U18712 ( .A(n16154), .ZN(n16177) );
  NOR2_X1 U18713 ( .A1(n15464), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16178) );
  OR3_X1 U18714 ( .A1(n16177), .A2(n16178), .A3(n19196), .ZN(n15473) );
  INV_X1 U18715 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19773) );
  NOR2_X1 U18716 ( .A1(n19773), .A2(n19045), .ZN(n15467) );
  NOR2_X1 U18717 ( .A1(n15465), .A2(n15470), .ZN(n15466) );
  AOI211_X1 U18718 ( .C1(n16181), .C2(n19192), .A(n15467), .B(n15466), .ZN(
        n15468) );
  OAI21_X1 U18719 ( .B1(n18999), .B2(n16289), .A(n15468), .ZN(n15469) );
  AOI21_X1 U18720 ( .B1(n15471), .B2(n15470), .A(n15469), .ZN(n15472) );
  OAI211_X1 U18721 ( .C1(n16176), .C2(n16305), .A(n15473), .B(n15472), .ZN(
        P2_U3037) );
  INV_X1 U18722 ( .A(n15474), .ZN(n16286) );
  NAND2_X1 U18723 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19029), .ZN(n15475) );
  OAI221_X1 U18724 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16272), .C1(
        n11696), .C2(n16286), .A(n15475), .ZN(n15479) );
  OAI22_X1 U18725 ( .A1(n15477), .A2(n16289), .B1(n16266), .B2(n15476), .ZN(
        n15478) );
  AOI211_X1 U18726 ( .C1(n15480), .C2(n19187), .A(n15479), .B(n15478), .ZN(
        n15481) );
  OAI21_X1 U18727 ( .B1(n15482), .B2(n19196), .A(n15481), .ZN(P2_U3039) );
  NOR2_X1 U18728 ( .A1(n19025), .A2(n16289), .ZN(n15491) );
  NAND2_X1 U18729 ( .A1(n15484), .A2(n15483), .ZN(n15489) );
  OAI21_X1 U18730 ( .B1(n16309), .B2(n15484), .A(n16296), .ZN(n15485) );
  NAND2_X1 U18731 ( .A1(n15485), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15488) );
  NOR2_X1 U18732 ( .A1(n19769), .A2(n19045), .ZN(n15486) );
  AOI21_X1 U18733 ( .B1(n19192), .B2(n19021), .A(n15486), .ZN(n15487) );
  OAI211_X1 U18734 ( .C1(n15489), .C2(n16298), .A(n15488), .B(n15487), .ZN(
        n15490) );
  AOI211_X1 U18735 ( .C1(n15492), .C2(n16281), .A(n15491), .B(n15490), .ZN(
        n15493) );
  OAI21_X1 U18736 ( .B1(n16305), .B2(n15494), .A(n15493), .ZN(P2_U3040) );
  NAND2_X1 U18737 ( .A1(n15496), .A2(n15495), .ZN(n15504) );
  MUX2_X1 U18738 ( .A(n15504), .B(n9741), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15497) );
  AOI21_X1 U18739 ( .B1(n19170), .B2(n15516), .A(n15497), .ZN(n15498) );
  INV_X1 U18740 ( .A(n15498), .ZN(n16327) );
  INV_X1 U18741 ( .A(n19078), .ZN(n15499) );
  AOI22_X1 U18742 ( .A1(n19052), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n15499), .B2(n19032), .ZN(n15511) );
  AOI222_X1 U18743 ( .A1(n16327), .A2(n19827), .B1(n15500), .B2(n16352), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15511), .ZN(n15502) );
  NAND2_X1 U18744 ( .A1(n15526), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15501) );
  OAI21_X1 U18745 ( .B1(n15502), .B2(n15526), .A(n15501), .ZN(P2_U3601) );
  NOR2_X1 U18746 ( .A1(n10789), .A2(n10788), .ZN(n15503) );
  AOI22_X1 U18747 ( .A1(n9741), .A2(n15505), .B1(n15504), .B2(n15503), .ZN(
        n15506) );
  OAI21_X1 U18748 ( .B1(n15508), .B2(n15507), .A(n15506), .ZN(n16328) );
  OAI21_X1 U18749 ( .B1(n19032), .B2(n15510), .A(n15509), .ZN(n15525) );
  INV_X1 U18750 ( .A(n15525), .ZN(n15512) );
  NOR2_X1 U18751 ( .A1(n15511), .A2(n11189), .ZN(n15524) );
  AOI222_X1 U18752 ( .A1(n16328), .A2(n19827), .B1(n19848), .B2(n16352), .C1(
        n15512), .C2(n15524), .ZN(n15514) );
  NAND2_X1 U18753 ( .A1(n15526), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15513) );
  OAI21_X1 U18754 ( .B1(n15514), .B2(n15526), .A(n15513), .ZN(P2_U3600) );
  AND2_X1 U18755 ( .A1(n10794), .A2(n15515), .ZN(n15522) );
  NAND2_X1 U18756 ( .A1(n15517), .A2(n15516), .ZN(n15521) );
  AOI22_X1 U18757 ( .A1(n15519), .A2(n9741), .B1(n15518), .B2(n15522), .ZN(
        n15520) );
  OAI211_X1 U18758 ( .C1(n15523), .C2(n15522), .A(n15521), .B(n15520), .ZN(
        n16312) );
  AOI222_X1 U18759 ( .A1(n16312), .A2(n19827), .B1(n19282), .B2(n16352), .C1(
        n15525), .C2(n15524), .ZN(n15528) );
  MUX2_X1 U18760 ( .A(n15528), .B(n15527), .S(n15526), .Z(n15529) );
  INV_X1 U18761 ( .A(n15529), .ZN(P2_U3599) );
  NAND2_X1 U18762 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18378) );
  AOI221_X1 U18763 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18378), .C1(n15531), 
        .C2(n18378), .A(n15530), .ZN(n18195) );
  NOR2_X1 U18764 ( .A1(n15532), .A2(n18675), .ZN(n15533) );
  OAI21_X1 U18765 ( .B1(n15533), .B2(n18496), .A(n18196), .ZN(n18193) );
  AOI22_X1 U18766 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18195), .B1(
        n18193), .B2(n18197), .ZN(P3_U2865) );
  NOR2_X1 U18767 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18810), .ZN(n18203) );
  NAND2_X1 U18768 ( .A1(n18649), .A2(n18707), .ZN(n15539) );
  INV_X1 U18769 ( .A(n18732), .ZN(n18854) );
  NAND3_X1 U18770 ( .A1(n18854), .A2(n16508), .A3(n15534), .ZN(n17390) );
  NOR3_X1 U18771 ( .A1(n15537), .A2(n15643), .A3(n15536), .ZN(n15538) );
  OAI21_X1 U18772 ( .B1(n15539), .B2(n17390), .A(n15538), .ZN(n18689) );
  INV_X1 U18773 ( .A(n18689), .ZN(n18690) );
  INV_X1 U18774 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18191) );
  OAI22_X1 U18775 ( .A1(n18690), .A2(n18713), .B1(n18191), .B2(n18808), .ZN(
        n15540) );
  INV_X1 U18776 ( .A(n18829), .ZN(n18837) );
  INV_X1 U18777 ( .A(n18666), .ZN(n18659) );
  AOI21_X1 U18778 ( .B1(n18659), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15541) );
  NOR2_X1 U18779 ( .A1(n15541), .A2(n16507), .ZN(n18702) );
  NAND3_X1 U18780 ( .A1(n18839), .A2(n18837), .A3(n18702), .ZN(n15542) );
  OAI21_X1 U18781 ( .B1(n18839), .B2(n18655), .A(n15542), .ZN(P3_U3284) );
  INV_X1 U18782 ( .A(n18088), .ZN(n17993) );
  INV_X1 U18783 ( .A(n18068), .ZN(n18018) );
  AOI21_X1 U18784 ( .B1(n18018), .B2(n10076), .A(n15543), .ZN(n16398) );
  OAI21_X1 U18785 ( .B1(n17993), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16398), .ZN(n15546) );
  NOR2_X1 U18786 ( .A1(n18651), .A2(n18185), .ZN(n18184) );
  NOR2_X1 U18787 ( .A1(n16391), .A2(n18177), .ZN(n15544) );
  INV_X1 U18788 ( .A(n18145), .ZN(n18182) );
  NAND2_X1 U18789 ( .A1(n17506), .A2(n15616), .ZN(n16363) );
  AOI22_X1 U18790 ( .A1(n15544), .A2(n16362), .B1(n18182), .B2(n16363), .ZN(
        n15620) );
  INV_X1 U18791 ( .A(n15620), .ZN(n15545) );
  AOI21_X1 U18792 ( .B1(n18179), .B2(n15546), .A(n15545), .ZN(n15555) );
  NAND2_X1 U18793 ( .A1(n15548), .A2(n15547), .ZN(n15549) );
  INV_X1 U18794 ( .A(n16383), .ZN(n15553) );
  INV_X1 U18795 ( .A(n17506), .ZN(n17869) );
  OAI22_X1 U18796 ( .A1(n9765), .A2(n17869), .B1(n16395), .B2(n18023), .ZN(
        n15550) );
  OAI21_X1 U18797 ( .B1(n15551), .B2(n15550), .A(n18163), .ZN(n15623) );
  NOR3_X1 U18798 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16396), .A3(
        n15623), .ZN(n15552) );
  AOI21_X1 U18799 ( .B1(n18099), .B2(n15553), .A(n15552), .ZN(n15554) );
  NAND2_X1 U18800 ( .A1(n9732), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16378) );
  OAI211_X1 U18801 ( .C1(n15555), .C2(n16387), .A(n15554), .B(n16378), .ZN(
        P3_U2833) );
  INV_X1 U18802 ( .A(n15556), .ZN(n15557) );
  AOI22_X1 U18803 ( .A1(n15557), .A2(n19070), .B1(n16078), .B2(n19042), .ZN(
        n15566) );
  AOI22_X1 U18804 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19043), .B1(
        P2_EBX_REG_22__SCAN_IN), .B2(n19065), .ZN(n15562) );
  OAI211_X1 U18805 ( .C1(n15560), .C2(n15559), .A(n19036), .B(n15558), .ZN(
        n15561) );
  OAI211_X1 U18806 ( .C1(n19061), .C2(n19796), .A(n15562), .B(n15561), .ZN(
        n15563) );
  AOI21_X1 U18807 ( .B1(n19041), .B2(n15564), .A(n15563), .ZN(n15565) );
  NAND2_X1 U18808 ( .A1(n15566), .A2(n15565), .ZN(P2_U2833) );
  NAND3_X1 U18809 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20799), .A3(n20708), 
        .ZN(n15567) );
  AOI22_X1 U18810 ( .A1(n15570), .A2(n15569), .B1(n15568), .B2(n15567), .ZN(
        n15975) );
  NOR2_X1 U18811 ( .A1(n15571), .A2(n20568), .ZN(n15572) );
  AND2_X1 U18812 ( .A1(n15573), .A2(n15572), .ZN(n15574) );
  NAND2_X1 U18813 ( .A1(n15574), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n15578) );
  INV_X1 U18814 ( .A(n15584), .ZN(n15576) );
  OAI22_X1 U18815 ( .A1(n15576), .A2(n15575), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n15574), .ZN(n15577) );
  NAND2_X1 U18816 ( .A1(n15578), .A2(n15577), .ZN(n15581) );
  NAND2_X1 U18817 ( .A1(n15584), .A2(n13067), .ZN(n15580) );
  AOI222_X1 U18818 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15581), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15580), .C1(n15581), 
        .C2(n15580), .ZN(n15586) );
  INV_X1 U18819 ( .A(n15582), .ZN(n15583) );
  AND2_X1 U18820 ( .A1(n15584), .A2(n15583), .ZN(n15585) );
  AOI222_X1 U18821 ( .A1(n15586), .A2(n20488), .B1(n15586), .B2(n15585), .C1(
        n20488), .C2(n15585), .ZN(n15589) );
  OAI211_X1 U18822 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15589), .A(
        n15588), .B(n15587), .ZN(n15591) );
  NOR2_X1 U18823 ( .A1(n15591), .A2(n15590), .ZN(n15596) );
  OR2_X1 U18824 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n15593) );
  AOI21_X1 U18825 ( .B1(n15594), .B2(n15593), .A(n15592), .ZN(n15595) );
  AOI21_X1 U18826 ( .B1(n15596), .B2(n15595), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n15597) );
  INV_X1 U18827 ( .A(n15597), .ZN(n15599) );
  AOI21_X1 U18828 ( .B1(n15599), .B2(n15975), .A(n20708), .ZN(n15982) );
  INV_X1 U18829 ( .A(n15982), .ZN(n15980) );
  OAI221_X1 U18830 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15977), .C1(n11980), 
        .C2(n15599), .A(n15598), .ZN(n15600) );
  NOR3_X1 U18831 ( .A1(n15601), .A2(n15980), .A3(n15600), .ZN(n15604) );
  AND3_X1 U18832 ( .A1(n20708), .A2(n20801), .A3(n15602), .ZN(n15603) );
  AOI211_X1 U18833 ( .C1(n15975), .C2(n15605), .A(n15604), .B(n15603), .ZN(
        P1_U3161) );
  OAI22_X1 U18834 ( .A1(n15609), .A2(n15608), .B1(n15607), .B2(n15606), .ZN(
        n15610) );
  XNOR2_X1 U18835 ( .A(n15610), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15779) );
  AOI22_X1 U18836 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n13397), .B1(n15611), 
        .B2(n12804), .ZN(n15615) );
  INV_X1 U18837 ( .A(n15693), .ZN(n15612) );
  AOI22_X1 U18838 ( .A1(n15613), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n15612), .B2(n20126), .ZN(n15614) );
  OAI211_X1 U18839 ( .C1(n15779), .C2(n15913), .A(n15615), .B(n15614), .ZN(
        P1_U3010) );
  NAND2_X1 U18840 ( .A1(n15616), .A2(n16364), .ZN(n16373) );
  AOI21_X1 U18841 ( .B1(n15618), .B2(n16364), .A(n15617), .ZN(n16370) );
  AOI21_X1 U18842 ( .B1(n15620), .B2(n15619), .A(n16364), .ZN(n15621) );
  AOI21_X1 U18843 ( .B1(n18099), .B2(n16370), .A(n15621), .ZN(n15622) );
  NAND2_X1 U18844 ( .A1(n9732), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16365) );
  OAI211_X1 U18845 ( .C1(n16373), .C2(n15623), .A(n15622), .B(n16365), .ZN(
        P3_U2832) );
  INV_X1 U18846 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20877) );
  INV_X1 U18847 ( .A(HOLD), .ZN(n20717) );
  NOR2_X1 U18848 ( .A1(n20877), .A2(n20717), .ZN(n20713) );
  AOI22_X1 U18849 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15625) );
  NAND2_X1 U18850 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20799), .ZN(n20716) );
  OAI211_X1 U18851 ( .C1(n20713), .C2(n15625), .A(n15624), .B(n20716), .ZN(
        P1_U3195) );
  INV_X1 U18852 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16482) );
  NOR2_X1 U18853 ( .A1(n20044), .A2(n16482), .ZN(P1_U2905) );
  INV_X1 U18854 ( .A(n15872), .ZN(n15631) );
  NOR2_X1 U18855 ( .A1(n20110), .A2(n15626), .ZN(n15628) );
  AOI21_X1 U18856 ( .B1(n15890), .B2(n15628), .A(n15627), .ZN(n15891) );
  AOI21_X1 U18857 ( .B1(n15891), .B2(n15893), .A(n15629), .ZN(n15630) );
  OAI22_X1 U18858 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15866), .B1(
        n15631), .B2(n15630), .ZN(n15637) );
  AOI22_X1 U18859 ( .A1(n15633), .A2(n20128), .B1(n20126), .B2(n15632), .ZN(
        n15636) );
  INV_X1 U18860 ( .A(n15634), .ZN(n15635) );
  OAI211_X1 U18861 ( .C1(n15638), .C2(n15637), .A(n15636), .B(n15635), .ZN(
        P1_U3011) );
  INV_X1 U18862 ( .A(n15639), .ZN(n19878) );
  NOR3_X1 U18863 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19884), .A3(n19880), 
        .ZN(n16343) );
  NOR4_X1 U18864 ( .A1(n15640), .A2(n19878), .A3(n16343), .A4(n16359), .ZN(
        P2_U3178) );
  AOI221_X1 U18865 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16359), .C1(n19864), .C2(
        n16359), .A(n19651), .ZN(n19854) );
  INV_X1 U18866 ( .A(n19854), .ZN(n19862) );
  NOR2_X1 U18867 ( .A1(n20834), .A2(n19862), .ZN(P2_U3047) );
  NOR3_X1 U18868 ( .A1(n15641), .A2(n17392), .A3(n18855), .ZN(n15642) );
  NAND2_X1 U18869 ( .A1(n18240), .A2(n17233), .ZN(n17376) );
  INV_X1 U18870 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17453) );
  AOI22_X1 U18871 ( .A1(n17384), .A2(BUF2_REG_0__SCAN_IN), .B1(n17344), .B2(
        n10347), .ZN(n15645) );
  OAI221_X1 U18872 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17376), .C1(n17453), 
        .C2(n17233), .A(n15645), .ZN(P3_U2735) );
  NOR2_X1 U18873 ( .A1(n15647), .A2(n15646), .ZN(n15654) );
  INV_X1 U18874 ( .A(n15648), .ZN(n15649) );
  NOR3_X1 U18875 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n15662), .A3(n15649), 
        .ZN(n15653) );
  OAI22_X1 U18876 ( .A1(n19946), .A2(n15651), .B1(n19993), .B2(n15650), .ZN(
        n15652) );
  AOI211_X1 U18877 ( .C1(n15654), .C2(P1_REIP_REG_26__SCAN_IN), .A(n15653), 
        .B(n15652), .ZN(n15658) );
  AOI22_X1 U18878 ( .A1(n15656), .A2(n19949), .B1(n15655), .B2(n19982), .ZN(
        n15657) );
  OAI211_X1 U18879 ( .C1(n15659), .C2(n19988), .A(n15658), .B(n15657), .ZN(
        P1_U2814) );
  INV_X1 U18880 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20762) );
  AOI21_X1 U18881 ( .B1(n19985), .B2(n20762), .A(n15673), .ZN(n15660) );
  NOR2_X1 U18882 ( .A1(n15660), .A2(n20764), .ZN(n15666) );
  NOR3_X1 U18883 ( .A1(n15662), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n15661), 
        .ZN(n15665) );
  OAI22_X1 U18884 ( .A1(n19946), .A2(n15663), .B1(n12428), .B2(n19993), .ZN(
        n15664) );
  NOR3_X1 U18885 ( .A1(n15666), .A2(n15665), .A3(n15664), .ZN(n15671) );
  OAI22_X1 U18886 ( .A1(n15668), .A2(n15751), .B1(n15667), .B2(n19988), .ZN(
        n15669) );
  INV_X1 U18887 ( .A(n15669), .ZN(n15670) );
  OAI211_X1 U18888 ( .C1(n15672), .C2(n19992), .A(n15671), .B(n15670), .ZN(
        P1_U2815) );
  INV_X1 U18889 ( .A(n15673), .ZN(n15679) );
  INV_X1 U18890 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20757) );
  NOR3_X1 U18891 ( .A1(n15680), .A2(n20757), .A3(n15728), .ZN(n15685) );
  AOI21_X1 U18892 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15685), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15678) );
  INV_X1 U18893 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15674) );
  OAI22_X1 U18894 ( .A1(n15674), .A2(n19993), .B1(n19992), .B2(n15777), .ZN(
        n15675) );
  AOI21_X1 U18895 ( .B1(n19994), .B2(P1_EBX_REG_23__SCAN_IN), .A(n15675), .ZN(
        n15677) );
  AOI22_X1 U18896 ( .A1(n15774), .A2(n19949), .B1(n15860), .B2(n19991), .ZN(
        n15676) );
  OAI211_X1 U18897 ( .C1(n15679), .C2(n15678), .A(n15677), .B(n15676), .ZN(
        P1_U2817) );
  NOR3_X1 U18898 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15680), .A3(n15728), 
        .ZN(n15695) );
  INV_X1 U18899 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20759) );
  INV_X1 U18900 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15683) );
  AOI22_X1 U18901 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19975), .B1(
        n19982), .B2(n15681), .ZN(n15682) );
  OAI21_X1 U18902 ( .B1(n19946), .B2(n15683), .A(n15682), .ZN(n15684) );
  AOI21_X1 U18903 ( .B1(n15685), .B2(n20759), .A(n15684), .ZN(n15686) );
  OAI21_X1 U18904 ( .B1(n15687), .B2(n15751), .A(n15686), .ZN(n15688) );
  AOI221_X1 U18905 ( .B1(n15695), .B2(P1_REIP_REG_22__SCAN_IN), .C1(n15691), 
        .C2(P1_REIP_REG_22__SCAN_IN), .A(n15688), .ZN(n15689) );
  OAI21_X1 U18906 ( .B1(n19988), .B2(n15690), .A(n15689), .ZN(P1_U2818) );
  AOI22_X1 U18907 ( .A1(n19994), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n19975), .ZN(n15699) );
  INV_X1 U18908 ( .A(n15780), .ZN(n15692) );
  AOI22_X1 U18909 ( .A1(n15692), .A2(n19982), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n15691), .ZN(n15698) );
  OAI22_X1 U18910 ( .A1(n15778), .A2(n15751), .B1(n19988), .B2(n15693), .ZN(
        n15694) );
  INV_X1 U18911 ( .A(n15694), .ZN(n15697) );
  INV_X1 U18912 ( .A(n15695), .ZN(n15696) );
  NAND4_X1 U18913 ( .A1(n15699), .A2(n15698), .A3(n15697), .A4(n15696), .ZN(
        P1_U2819) );
  INV_X1 U18914 ( .A(n15791), .ZN(n15700) );
  AOI22_X1 U18915 ( .A1(n19994), .A2(P1_EBX_REG_19__SCAN_IN), .B1(n15700), 
        .B2(n19982), .ZN(n15707) );
  INV_X1 U18916 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20752) );
  NOR3_X1 U18917 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n20752), .A3(n15703), 
        .ZN(n15701) );
  AOI211_X1 U18918 ( .C1(n19975), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15701), .B(n19964), .ZN(n15706) );
  NOR2_X1 U18919 ( .A1(n15867), .A2(n19988), .ZN(n15702) );
  AOI21_X1 U18920 ( .B1(n15788), .B2(n19949), .A(n15702), .ZN(n15705) );
  NOR2_X1 U18921 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15703), .ZN(n15708) );
  OAI21_X1 U18922 ( .B1(n15708), .B2(n15718), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15704) );
  NAND4_X1 U18923 ( .A1(n15707), .A2(n15706), .A3(n15705), .A4(n15704), .ZN(
        P1_U2821) );
  INV_X1 U18924 ( .A(n15708), .ZN(n15713) );
  OAI21_X1 U18925 ( .B1(n19993), .B2(n15709), .A(n19954), .ZN(n15710) );
  AOI21_X1 U18926 ( .B1(n15711), .B2(n19982), .A(n15710), .ZN(n15712) );
  OAI211_X1 U18927 ( .C1(n15714), .C2(n19946), .A(n15713), .B(n15712), .ZN(
        n15717) );
  NOR2_X1 U18928 ( .A1(n15715), .A2(n15751), .ZN(n15716) );
  AOI211_X1 U18929 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15718), .A(n15717), 
        .B(n15716), .ZN(n15719) );
  OAI21_X1 U18930 ( .B1(n19988), .B2(n15720), .A(n15719), .ZN(P1_U2822) );
  AOI22_X1 U18931 ( .A1(n15809), .A2(n19982), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n15721), .ZN(n15727) );
  OAI21_X1 U18932 ( .B1(n19993), .B2(n15722), .A(n19954), .ZN(n15723) );
  AOI21_X1 U18933 ( .B1(n19994), .B2(P1_EBX_REG_15__SCAN_IN), .A(n15723), .ZN(
        n15724) );
  OAI21_X1 U18934 ( .B1(n19988), .B2(n15884), .A(n15724), .ZN(n15725) );
  AOI21_X1 U18935 ( .B1(n15810), .B2(n19949), .A(n15725), .ZN(n15726) );
  OAI211_X1 U18936 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15728), .A(n15727), 
        .B(n15726), .ZN(P1_U2825) );
  AOI21_X1 U18937 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n15729), .A(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15739) );
  OAI21_X1 U18938 ( .B1(n19993), .B2(n15730), .A(n19954), .ZN(n15733) );
  NOR2_X1 U18939 ( .A1(n19988), .A2(n15731), .ZN(n15732) );
  AOI211_X1 U18940 ( .C1(n19994), .C2(P1_EBX_REG_14__SCAN_IN), .A(n15733), .B(
        n15732), .ZN(n15738) );
  INV_X1 U18941 ( .A(n15734), .ZN(n15735) );
  AOI22_X1 U18942 ( .A1(n15736), .A2(n19949), .B1(n19982), .B2(n15735), .ZN(
        n15737) );
  OAI211_X1 U18943 ( .C1(n15740), .C2(n15739), .A(n15738), .B(n15737), .ZN(
        P1_U2826) );
  INV_X1 U18944 ( .A(n15908), .ZN(n15741) );
  NAND2_X1 U18945 ( .A1(n19991), .A2(n15741), .ZN(n15744) );
  NAND2_X1 U18946 ( .A1(n19975), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15742) );
  AND2_X1 U18947 ( .A1(n15742), .A2(n19954), .ZN(n15743) );
  OAI211_X1 U18948 ( .C1(n19946), .C2(n13893), .A(n15744), .B(n15743), .ZN(
        n15745) );
  INV_X1 U18949 ( .A(n15745), .ZN(n15750) );
  AOI21_X1 U18950 ( .B1(n20741), .B2(n15747), .A(n15746), .ZN(n15748) );
  AOI21_X1 U18951 ( .B1(n19982), .B2(n15819), .A(n15748), .ZN(n15749) );
  OAI211_X1 U18952 ( .C1(n15751), .C2(n15817), .A(n15750), .B(n15749), .ZN(
        P1_U2828) );
  XOR2_X1 U18953 ( .A(n15753), .B(n15752), .Z(n15827) );
  INV_X1 U18954 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15767) );
  INV_X1 U18955 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15754) );
  NAND3_X1 U18956 ( .A1(n19985), .A2(n15755), .A3(n15754), .ZN(n15756) );
  OAI21_X1 U18957 ( .B1(n15767), .B2(n19946), .A(n15756), .ZN(n15764) );
  NOR2_X1 U18958 ( .A1(n15758), .A2(n15757), .ZN(n15759) );
  AOI22_X1 U18959 ( .A1(n19991), .A2(n9826), .B1(P1_REIP_REG_11__SCAN_IN), 
        .B2(n15761), .ZN(n15762) );
  OAI211_X1 U18960 ( .C1(n19993), .C2(n12163), .A(n15762), .B(n19954), .ZN(
        n15763) );
  AOI211_X1 U18961 ( .C1(n19949), .C2(n15827), .A(n15764), .B(n15763), .ZN(
        n15765) );
  OAI21_X1 U18962 ( .B1(n15830), .B2(n19992), .A(n15765), .ZN(P1_U2829) );
  AOI22_X1 U18963 ( .A1(n15827), .A2(n20008), .B1(n20007), .B2(n9826), .ZN(
        n15766) );
  OAI21_X1 U18964 ( .B1(n20012), .B2(n15767), .A(n15766), .ZN(P1_U2861) );
  AOI22_X1 U18965 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(n15768), .B1(n15770), 
        .B2(n20057), .ZN(n15769) );
  OAI21_X1 U18966 ( .B1(n20016), .B2(n15817), .A(n15769), .ZN(P1_U2892) );
  INV_X1 U18967 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20896) );
  AOI22_X1 U18968 ( .A1(n15771), .A2(n15827), .B1(n15770), .B2(n20055), .ZN(
        n15772) );
  OAI21_X1 U18969 ( .B1(n20015), .B2(n20896), .A(n15772), .ZN(P1_U2893) );
  AOI22_X1 U18970 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n15776) );
  XNOR2_X1 U18971 ( .A(n9738), .B(n15864), .ZN(n15773) );
  XNOR2_X1 U18972 ( .A(n14642), .B(n15773), .ZN(n15861) );
  AOI22_X1 U18973 ( .A1(n15774), .A2(n14666), .B1(n20081), .B2(n15861), .ZN(
        n15775) );
  OAI211_X1 U18974 ( .C1(n20085), .C2(n15777), .A(n15776), .B(n15775), .ZN(
        P1_U2976) );
  INV_X1 U18975 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15785) );
  OAI222_X1 U18976 ( .A1(n20085), .A2(n15780), .B1(n19900), .B2(n15779), .C1(
        n20142), .C2(n15778), .ZN(n15781) );
  INV_X1 U18977 ( .A(n15781), .ZN(n15783) );
  NAND2_X1 U18978 ( .A1(n13397), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15782) );
  OAI211_X1 U18979 ( .C1(n15785), .C2(n15784), .A(n15783), .B(n15782), .ZN(
        P1_U2978) );
  AOI22_X1 U18980 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15790) );
  MUX2_X1 U18981 ( .A(n9738), .B(n15786), .S(n14692), .Z(n15787) );
  XOR2_X1 U18982 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n15787), .Z(
        n15869) );
  AOI22_X1 U18983 ( .A1(n15869), .A2(n20081), .B1(n14666), .B2(n15788), .ZN(
        n15789) );
  OAI211_X1 U18984 ( .C1(n20085), .C2(n15791), .A(n15790), .B(n15789), .ZN(
        P1_U2980) );
  AOI21_X1 U18985 ( .B1(n14706), .B2(n15793), .A(n15792), .ZN(n15796) );
  NOR2_X1 U18986 ( .A1(n15796), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15795) );
  MUX2_X1 U18987 ( .A(n15796), .B(n15795), .S(n15794), .Z(n15797) );
  XNOR2_X1 U18988 ( .A(n15797), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15882) );
  AOI22_X1 U18989 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15801) );
  AOI22_X1 U18990 ( .A1(n15799), .A2(n14666), .B1(n15820), .B2(n15798), .ZN(
        n15800) );
  OAI211_X1 U18991 ( .C1(n19900), .C2(n15882), .A(n15801), .B(n15800), .ZN(
        P1_U2982) );
  INV_X1 U18992 ( .A(n15802), .ZN(n15803) );
  NOR2_X1 U18993 ( .A1(n15804), .A2(n15803), .ZN(n15808) );
  NOR2_X1 U18994 ( .A1(n15806), .A2(n15805), .ZN(n15807) );
  XOR2_X1 U18995 ( .A(n15808), .B(n15807), .Z(n15889) );
  AOI22_X1 U18996 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15812) );
  AOI22_X1 U18997 ( .A1(n15810), .A2(n14666), .B1(n15809), .B2(n15820), .ZN(
        n15811) );
  OAI211_X1 U18998 ( .C1(n15889), .C2(n19900), .A(n15812), .B(n15811), .ZN(
        P1_U2984) );
  INV_X1 U18999 ( .A(n15813), .ZN(n15814) );
  AOI21_X1 U19000 ( .B1(n15816), .B2(n15815), .A(n15814), .ZN(n15914) );
  AOI22_X1 U19001 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15822) );
  INV_X1 U19002 ( .A(n15817), .ZN(n15818) );
  AOI22_X1 U19003 ( .A1(n15820), .A2(n15819), .B1(n14666), .B2(n15818), .ZN(
        n15821) );
  OAI211_X1 U19004 ( .C1(n15914), .C2(n19900), .A(n15822), .B(n15821), .ZN(
        P1_U2987) );
  AOI22_X1 U19005 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15829) );
  NAND2_X1 U19006 ( .A1(n9738), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15825) );
  OAI21_X1 U19007 ( .B1(n14706), .B2(n15825), .A(n15824), .ZN(n15826) );
  INV_X1 U19008 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15921) );
  XNOR2_X1 U19009 ( .A(n15826), .B(n15921), .ZN(n15916) );
  AOI22_X1 U19010 ( .A1(n20081), .A2(n15916), .B1(n14666), .B2(n15827), .ZN(
        n15828) );
  OAI211_X1 U19011 ( .C1(n20085), .C2(n15830), .A(n15829), .B(n15828), .ZN(
        P1_U2988) );
  AOI22_X1 U19012 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15836) );
  NAND2_X1 U19013 ( .A1(n15833), .A2(n15832), .ZN(n15834) );
  XNOR2_X1 U19014 ( .A(n15831), .B(n15834), .ZN(n15956) );
  AOI22_X1 U19015 ( .A1(n15956), .A2(n20081), .B1(n14666), .B2(n19937), .ZN(
        n15835) );
  OAI211_X1 U19016 ( .C1(n20085), .C2(n19939), .A(n15836), .B(n15835), .ZN(
        P1_U2992) );
  AOI22_X1 U19017 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15842) );
  XNOR2_X1 U19018 ( .A(n15838), .B(n15837), .ZN(n15839) );
  XNOR2_X1 U19019 ( .A(n15840), .B(n15839), .ZN(n15962) );
  AOI22_X1 U19020 ( .A1(n15962), .A2(n20081), .B1(n14666), .B2(n19950), .ZN(
        n15841) );
  OAI211_X1 U19021 ( .C1(n20085), .C2(n19953), .A(n15842), .B(n15841), .ZN(
        P1_U2993) );
  AOI22_X1 U19022 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15849) );
  INV_X1 U19023 ( .A(n15843), .ZN(n15844) );
  AOI21_X1 U19024 ( .B1(n15846), .B2(n15845), .A(n15844), .ZN(n15969) );
  INV_X1 U19025 ( .A(n15847), .ZN(n20009) );
  AOI22_X1 U19026 ( .A1(n15969), .A2(n20081), .B1(n14666), .B2(n20009), .ZN(
        n15848) );
  OAI211_X1 U19027 ( .C1(n20085), .C2(n19962), .A(n15849), .B(n15848), .ZN(
        P1_U2994) );
  AOI21_X1 U19028 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15859), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15858) );
  AOI211_X1 U19029 ( .C1(n15852), .C2(n15864), .A(n15851), .B(n15850), .ZN(
        n15857) );
  AOI22_X1 U19030 ( .A1(n15854), .A2(n20128), .B1(n20126), .B2(n15853), .ZN(
        n15856) );
  NAND2_X1 U19031 ( .A1(n13397), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15855) );
  OAI211_X1 U19032 ( .C1(n15858), .C2(n15857), .A(n15856), .B(n15855), .ZN(
        P1_U3007) );
  AOI22_X1 U19033 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n13397), .B1(n15859), 
        .B2(n15864), .ZN(n15863) );
  AOI22_X1 U19034 ( .A1(n15861), .A2(n20128), .B1(n20126), .B2(n15860), .ZN(
        n15862) );
  OAI211_X1 U19035 ( .C1(n15865), .C2(n15864), .A(n15863), .B(n15862), .ZN(
        P1_U3008) );
  INV_X1 U19036 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15873) );
  AOI22_X1 U19037 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n13397), .B1(n15866), 
        .B2(n15873), .ZN(n15871) );
  INV_X1 U19038 ( .A(n15867), .ZN(n15868) );
  AOI22_X1 U19039 ( .A1(n15869), .A2(n20128), .B1(n20126), .B2(n15868), .ZN(
        n15870) );
  OAI211_X1 U19040 ( .C1(n15873), .C2(n15872), .A(n15871), .B(n15870), .ZN(
        P1_U3012) );
  OAI21_X1 U19041 ( .B1(n15875), .B2(n15874), .A(n12801), .ZN(n15879) );
  INV_X1 U19042 ( .A(n15876), .ZN(n15877) );
  AOI22_X1 U19043 ( .A1(n15879), .A2(n15878), .B1(n20126), .B2(n15877), .ZN(
        n15881) );
  NAND2_X1 U19044 ( .A1(n13397), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15880) );
  OAI211_X1 U19045 ( .C1(n15882), .C2(n15913), .A(n15881), .B(n15880), .ZN(
        P1_U3014) );
  AOI22_X1 U19046 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15883), .B1(
        n13397), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15888) );
  NOR2_X1 U19047 ( .A1(n15884), .A2(n20109), .ZN(n15885) );
  NOR2_X1 U19048 ( .A1(n15886), .A2(n15885), .ZN(n15887) );
  OAI211_X1 U19049 ( .C1(n15889), .C2(n15913), .A(n15888), .B(n15887), .ZN(
        P1_U3016) );
  INV_X1 U19050 ( .A(n15890), .ZN(n15892) );
  OAI21_X1 U19051 ( .B1(n15893), .B2(n15892), .A(n15891), .ZN(n15894) );
  AOI22_X1 U19052 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n13397), .B1(n15899), 
        .B2(n15894), .ZN(n15898) );
  AOI22_X1 U19053 ( .A1(n15896), .A2(n20128), .B1(n20126), .B2(n15895), .ZN(
        n15897) );
  OAI211_X1 U19054 ( .C1(n15900), .C2(n15899), .A(n15898), .B(n15897), .ZN(
        P1_U3018) );
  AOI21_X1 U19055 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15901), .A(
        n20114), .ZN(n15904) );
  AOI21_X1 U19056 ( .B1(n15902), .B2(n20086), .A(n20104), .ZN(n15903) );
  INV_X1 U19057 ( .A(n15903), .ZN(n15946) );
  AOI211_X1 U19058 ( .C1(n15947), .C2(n15905), .A(n15904), .B(n15946), .ZN(
        n15922) );
  OAI21_X1 U19059 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n20103), .A(
        n15922), .ZN(n15911) );
  NAND2_X1 U19060 ( .A1(n15906), .A2(n20098), .ZN(n15965) );
  NOR4_X1 U19061 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15921), .A3(
        n15907), .A4(n15965), .ZN(n15910) );
  OAI22_X1 U19062 ( .A1(n20109), .A2(n15908), .B1(n20741), .B2(n20107), .ZN(
        n15909) );
  AOI211_X1 U19063 ( .C1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15911), .A(
        n15910), .B(n15909), .ZN(n15912) );
  OAI21_X1 U19064 ( .B1(n15914), .B2(n15913), .A(n15912), .ZN(P1_U3019) );
  AOI22_X1 U19065 ( .A1(n20126), .A2(n9826), .B1(n13397), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15920) );
  NOR2_X1 U19066 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15915), .ZN(
        n15917) );
  AOI22_X1 U19067 ( .A1(n15918), .A2(n15917), .B1(n20128), .B2(n15916), .ZN(
        n15919) );
  OAI211_X1 U19068 ( .C1(n15922), .C2(n15921), .A(n15920), .B(n15919), .ZN(
        P1_U3020) );
  INV_X1 U19069 ( .A(n15947), .ZN(n15945) );
  OAI21_X1 U19070 ( .B1(n15945), .B2(n15923), .A(n15926), .ZN(n15925) );
  OAI21_X1 U19071 ( .B1(n15946), .B2(n15925), .A(n15924), .ZN(n15942) );
  INV_X1 U19072 ( .A(n15965), .ZN(n15951) );
  NAND2_X1 U19073 ( .A1(n15926), .A2(n15951), .ZN(n15933) );
  AOI221_X1 U19074 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14747), .C2(n15943), .A(
        n15933), .ZN(n15929) );
  OAI22_X1 U19075 ( .A1(n20109), .A2(n15927), .B1(n21000), .B2(n20107), .ZN(
        n15928) );
  AOI211_X1 U19076 ( .C1(n15930), .C2(n20128), .A(n15929), .B(n15928), .ZN(
        n15931) );
  OAI21_X1 U19077 ( .B1(n14747), .B2(n15942), .A(n15931), .ZN(P1_U3021) );
  INV_X1 U19078 ( .A(n15932), .ZN(n15940) );
  NOR2_X1 U19079 ( .A1(n15933), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15939) );
  NAND2_X1 U19080 ( .A1(n15935), .A2(n15934), .ZN(n15936) );
  NAND2_X1 U19081 ( .A1(n15937), .A2(n15936), .ZN(n20000) );
  INV_X1 U19082 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20946) );
  OAI22_X1 U19083 ( .A1(n20109), .A2(n20000), .B1(n20946), .B2(n20107), .ZN(
        n15938) );
  AOI211_X1 U19084 ( .C1(n15940), .C2(n20128), .A(n15939), .B(n15938), .ZN(
        n15941) );
  OAI21_X1 U19085 ( .B1(n15943), .B2(n15942), .A(n15941), .ZN(P1_U3022) );
  INV_X1 U19086 ( .A(n15944), .ZN(n15949) );
  NOR2_X1 U19087 ( .A1(n20089), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15968) );
  INV_X1 U19088 ( .A(n15968), .ZN(n15948) );
  AOI21_X1 U19089 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n15945), .ZN(n20105) );
  AOI211_X1 U19090 ( .C1(n20089), .C2(n15947), .A(n20105), .B(n15946), .ZN(
        n15973) );
  OAI21_X1 U19091 ( .B1(n15949), .B2(n15948), .A(n15973), .ZN(n15961) );
  AOI21_X1 U19092 ( .B1(n15837), .B2(n20123), .A(n15961), .ZN(n15958) );
  OAI22_X1 U19093 ( .A1(n20109), .A2(n15950), .B1(n20737), .B2(n20107), .ZN(
        n15953) );
  NAND2_X1 U19094 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15951), .ZN(
        n15960) );
  AOI221_X1 U19095 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n13736), .C2(n15959), .A(
        n15960), .ZN(n15952) );
  AOI211_X1 U19096 ( .C1(n15954), .C2(n20128), .A(n15953), .B(n15952), .ZN(
        n15955) );
  OAI21_X1 U19097 ( .B1(n15958), .B2(n13736), .A(n15955), .ZN(P1_U3023) );
  AOI222_X1 U19098 ( .A1(n15956), .A2(n20128), .B1(n20126), .B2(n19929), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(n13397), .ZN(n15957) );
  OAI221_X1 U19099 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15960), .C1(
        n15959), .C2(n15958), .A(n15957), .ZN(P1_U3024) );
  AOI22_X1 U19100 ( .A1(n20126), .A2(n19941), .B1(n13397), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n15964) );
  AOI22_X1 U19101 ( .A1(n15962), .A2(n20128), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15961), .ZN(n15963) );
  OAI211_X1 U19102 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15965), .A(
        n15964), .B(n15963), .ZN(P1_U3025) );
  AND2_X1 U19103 ( .A1(n15967), .A2(n15966), .ZN(n20006) );
  AOI22_X1 U19104 ( .A1(n20126), .A2(n20006), .B1(n13397), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n15971) );
  AOI22_X1 U19105 ( .A1(n15969), .A2(n20128), .B1(n20098), .B2(n15968), .ZN(
        n15970) );
  OAI211_X1 U19106 ( .C1(n15973), .C2(n15972), .A(n15971), .B(n15970), .ZN(
        P1_U3026) );
  NOR2_X1 U19107 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20799), .ZN(n15974) );
  OAI221_X1 U19108 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n20708), .C2(n15974), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20709) );
  AOI21_X1 U19109 ( .B1(n20709), .B2(n15981), .A(n15975), .ZN(n15979) );
  AOI21_X1 U19110 ( .B1(n20532), .B2(n15977), .A(n15976), .ZN(n15978) );
  AOI211_X1 U19111 ( .C1(n20707), .C2(n15980), .A(n15979), .B(n15978), .ZN(
        P1_U3162) );
  OAI22_X1 U19112 ( .A1(n15982), .A2(n20532), .B1(n20708), .B2(n15981), .ZN(
        P1_U3466) );
  INV_X1 U19113 ( .A(n15983), .ZN(n16016) );
  INV_X1 U19114 ( .A(n15984), .ZN(n16037) );
  AOI21_X1 U19115 ( .B1(n16097), .B2(n15986), .A(n15985), .ZN(n16099) );
  INV_X1 U19116 ( .A(n16099), .ZN(n16060) );
  NAND2_X1 U19117 ( .A1(n19032), .A2(n15987), .ZN(n16059) );
  NAND2_X1 U19118 ( .A1(n16060), .A2(n16059), .ZN(n16058) );
  NAND2_X1 U19119 ( .A1(n19032), .A2(n16058), .ZN(n16048) );
  NAND2_X1 U19120 ( .A1(n16049), .A2(n16048), .ZN(n16047) );
  NAND2_X1 U19121 ( .A1(n19032), .A2(n16047), .ZN(n16036) );
  NAND2_X1 U19122 ( .A1(n16037), .A2(n16036), .ZN(n16035) );
  NAND2_X1 U19123 ( .A1(n19032), .A2(n16035), .ZN(n16023) );
  NAND2_X1 U19124 ( .A1(n16024), .A2(n16023), .ZN(n16022) );
  NAND2_X1 U19125 ( .A1(n19032), .A2(n16022), .ZN(n16015) );
  NAND2_X1 U19126 ( .A1(n16016), .A2(n16015), .ZN(n16014) );
  NAND2_X1 U19127 ( .A1(n19032), .A2(n16014), .ZN(n16001) );
  NAND2_X1 U19128 ( .A1(n16002), .A2(n16001), .ZN(n16000) );
  AOI22_X1 U19129 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n19043), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n15988), .ZN(n15989) );
  OAI21_X1 U19130 ( .B1(n19814), .B2(n19061), .A(n15989), .ZN(n15990) );
  AOI21_X1 U19131 ( .B1(n15991), .B2(n19041), .A(n15990), .ZN(n15995) );
  AOI22_X1 U19132 ( .A1(n15993), .A2(n19070), .B1(n19042), .B2(n15992), .ZN(
        n15994) );
  OAI211_X1 U19133 ( .C1(n19077), .C2(n16000), .A(n15995), .B(n15994), .ZN(
        P2_U2824) );
  AOI22_X1 U19134 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19065), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19030), .ZN(n16006) );
  AOI22_X1 U19135 ( .A1(n15996), .A2(n19041), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19043), .ZN(n16005) );
  NOR2_X1 U19136 ( .A1(n15997), .A2(n19063), .ZN(n15998) );
  AOI21_X1 U19137 ( .B1(n15999), .B2(n19070), .A(n15998), .ZN(n16004) );
  OAI211_X1 U19138 ( .C1(n16002), .C2(n16001), .A(n19036), .B(n16000), .ZN(
        n16003) );
  NAND4_X1 U19139 ( .A1(n16006), .A2(n16005), .A3(n16004), .A4(n16003), .ZN(
        P2_U2825) );
  AOI22_X1 U19140 ( .A1(n19065), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19030), .ZN(n16007) );
  INV_X1 U19141 ( .A(n16007), .ZN(n16008) );
  AOI21_X1 U19142 ( .B1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19043), .A(
        n16008), .ZN(n16011) );
  NAND2_X1 U19143 ( .A1(n16009), .A2(n19041), .ZN(n16010) );
  OAI211_X1 U19144 ( .C1(n16012), .C2(n19047), .A(n16011), .B(n16010), .ZN(
        n16013) );
  INV_X1 U19145 ( .A(n16013), .ZN(n16018) );
  OAI211_X1 U19146 ( .C1(n16016), .C2(n16015), .A(n19036), .B(n16014), .ZN(
        n16017) );
  OAI211_X1 U19147 ( .C1(n19063), .C2(n15274), .A(n16018), .B(n16017), .ZN(
        P2_U2826) );
  AOI22_X1 U19148 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n19030), .B1(
        P2_EBX_REG_28__SCAN_IN), .B2(n19065), .ZN(n16028) );
  AOI22_X1 U19149 ( .A1(n16019), .A2(n19041), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19043), .ZN(n16027) );
  AOI22_X1 U19150 ( .A1(n16021), .A2(n19070), .B1(n16020), .B2(n19042), .ZN(
        n16026) );
  OAI211_X1 U19151 ( .C1(n16024), .C2(n16023), .A(n19036), .B(n16022), .ZN(
        n16025) );
  NAND4_X1 U19152 ( .A1(n16028), .A2(n16027), .A3(n16026), .A4(n16025), .ZN(
        P2_U2827) );
  INV_X1 U19153 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n16029) );
  OAI22_X1 U19154 ( .A1(n19014), .A2(n16029), .B1(n19807), .B2(n19061), .ZN(
        n16030) );
  AOI21_X1 U19155 ( .B1(n19043), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16030), .ZN(n16031) );
  OAI21_X1 U19156 ( .B1(n16032), .B2(n19067), .A(n16031), .ZN(n16033) );
  AOI21_X1 U19157 ( .B1(n16034), .B2(n19070), .A(n16033), .ZN(n16039) );
  OAI211_X1 U19158 ( .C1(n16037), .C2(n16036), .A(n19036), .B(n16035), .ZN(
        n16038) );
  OAI211_X1 U19159 ( .C1(n19063), .C2(n16040), .A(n16039), .B(n16038), .ZN(
        P2_U2828) );
  AOI22_X1 U19160 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19030), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19065), .ZN(n16053) );
  OR2_X1 U19161 ( .A1(n16041), .A2(n19067), .ZN(n16043) );
  NAND2_X1 U19162 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19043), .ZN(
        n16042) );
  AND2_X1 U19163 ( .A1(n16043), .A2(n16042), .ZN(n16052) );
  OAI22_X1 U19164 ( .A1(n16045), .A2(n19047), .B1(n16044), .B2(n19063), .ZN(
        n16046) );
  INV_X1 U19165 ( .A(n16046), .ZN(n16051) );
  OAI211_X1 U19166 ( .C1(n16049), .C2(n16048), .A(n19036), .B(n16047), .ZN(
        n16050) );
  NAND4_X1 U19167 ( .A1(n16053), .A2(n16052), .A3(n16051), .A4(n16050), .ZN(
        P2_U2829) );
  AOI22_X1 U19168 ( .A1(n19065), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19030), .ZN(n16055) );
  NAND2_X1 U19169 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19043), .ZN(
        n16054) );
  OAI211_X1 U19170 ( .C1(n16104), .C2(n19047), .A(n16055), .B(n16054), .ZN(
        n16056) );
  AOI21_X1 U19171 ( .B1(n16057), .B2(n19041), .A(n16056), .ZN(n16062) );
  OAI211_X1 U19172 ( .C1(n16060), .C2(n16059), .A(n19036), .B(n16058), .ZN(
        n16061) );
  OAI211_X1 U19173 ( .C1(n19063), .C2(n16063), .A(n16062), .B(n16061), .ZN(
        P2_U2830) );
  AOI22_X1 U19174 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19030), .B1(
        P2_EBX_REG_23__SCAN_IN), .B2(n19065), .ZN(n16072) );
  AOI22_X1 U19175 ( .A1(n16064), .A2(n19041), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19043), .ZN(n16071) );
  OAI22_X1 U19176 ( .A1(n16229), .A2(n19047), .B1(n16222), .B2(n19063), .ZN(
        n16065) );
  INV_X1 U19177 ( .A(n16065), .ZN(n16070) );
  OAI211_X1 U19178 ( .C1(n16068), .C2(n16067), .A(n19036), .B(n16066), .ZN(
        n16069) );
  NAND4_X1 U19179 ( .A1(n16072), .A2(n16071), .A3(n16070), .A4(n16069), .ZN(
        P2_U2832) );
  AOI22_X1 U19180 ( .A1(n19082), .A2(n19099), .B1(n19104), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16076) );
  AOI22_X1 U19181 ( .A1(n19084), .A2(BUF2_REG_24__SCAN_IN), .B1(n19083), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n16075) );
  AOI22_X1 U19182 ( .A1(n16073), .A2(n16079), .B1(n19087), .B2(n16215), .ZN(
        n16074) );
  NAND3_X1 U19183 ( .A1(n16076), .A2(n16075), .A3(n16074), .ZN(P2_U2895) );
  AOI22_X1 U19184 ( .A1(n19082), .A2(n16077), .B1(n19104), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16083) );
  AOI22_X1 U19185 ( .A1(n19084), .A2(BUF2_REG_22__SCAN_IN), .B1(n19083), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n16082) );
  AOI22_X1 U19186 ( .A1(n16080), .A2(n16079), .B1(n19087), .B2(n16078), .ZN(
        n16081) );
  NAND3_X1 U19187 ( .A1(n16083), .A2(n16082), .A3(n16081), .ZN(P2_U2897) );
  AOI22_X1 U19188 ( .A1(n19082), .A2(n16084), .B1(n19104), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16090) );
  AOI22_X1 U19189 ( .A1(n19084), .A2(BUF2_REG_20__SCAN_IN), .B1(n19083), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16089) );
  OAI22_X1 U19190 ( .A1(n16086), .A2(n16092), .B1(n19107), .B2(n16085), .ZN(
        n16087) );
  INV_X1 U19191 ( .A(n16087), .ZN(n16088) );
  NAND3_X1 U19192 ( .A1(n16090), .A2(n16089), .A3(n16088), .ZN(P2_U2899) );
  AOI22_X1 U19193 ( .A1(n19082), .A2(n19214), .B1(n19104), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16096) );
  AOI22_X1 U19194 ( .A1(n19084), .A2(BUF2_REG_18__SCAN_IN), .B1(n19083), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16095) );
  OAI22_X1 U19195 ( .A1(n18916), .A2(n16092), .B1(n19107), .B2(n16091), .ZN(
        n16093) );
  INV_X1 U19196 ( .A(n16093), .ZN(n16094) );
  NAND3_X1 U19197 ( .A1(n16096), .A2(n16095), .A3(n16094), .ZN(P2_U2901) );
  OAI22_X1 U19198 ( .A1(n16097), .A2(n16204), .B1(n19802), .B2(n19045), .ZN(
        n16098) );
  AOI21_X1 U19199 ( .B1(n16198), .B2(n16099), .A(n16098), .ZN(n16103) );
  AOI22_X1 U19200 ( .A1(n16101), .A2(n19175), .B1(n16200), .B2(n16100), .ZN(
        n16102) );
  OAI211_X1 U19201 ( .C1(n16158), .C2(n16104), .A(n16103), .B(n16102), .ZN(
        P2_U2989) );
  AOI22_X1 U19202 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19029), .B1(n16198), 
        .B2(n16105), .ZN(n16113) );
  OAI21_X1 U19203 ( .B1(n16108), .B2(n16107), .A(n16106), .ZN(n16228) );
  OAI21_X1 U19204 ( .B1(n16110), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16109), .ZN(n16234) );
  OAI222_X1 U19205 ( .A1(n16229), .A2(n16158), .B1(n16228), .B2(n19161), .C1(
        n16234), .C2(n19177), .ZN(n16111) );
  INV_X1 U19206 ( .A(n16111), .ZN(n16112) );
  OAI211_X1 U19207 ( .C1(n16114), .C2(n16204), .A(n16113), .B(n16112), .ZN(
        P2_U2991) );
  AOI22_X1 U19208 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19029), .B1(n16198), 
        .B2(n16115), .ZN(n16127) );
  INV_X1 U19209 ( .A(n16130), .ZN(n16116) );
  OR2_X1 U19210 ( .A1(n16117), .A2(n16116), .ZN(n16121) );
  AND2_X1 U19211 ( .A1(n16119), .A2(n16118), .ZN(n16120) );
  XNOR2_X1 U19212 ( .A(n16121), .B(n16120), .ZN(n16245) );
  NAND2_X1 U19213 ( .A1(n19171), .A2(n16241), .ZN(n16124) );
  XNOR2_X1 U19214 ( .A(n16122), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16242) );
  NAND2_X1 U19215 ( .A1(n16242), .A2(n16200), .ZN(n16123) );
  OAI211_X1 U19216 ( .C1(n16245), .C2(n19161), .A(n16124), .B(n16123), .ZN(
        n16125) );
  INV_X1 U19217 ( .A(n16125), .ZN(n16126) );
  OAI211_X1 U19218 ( .C1(n16128), .C2(n16204), .A(n16127), .B(n16126), .ZN(
        P2_U2999) );
  AOI22_X1 U19219 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19169), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19029), .ZN(n16137) );
  AOI21_X1 U19220 ( .B1(n16251), .B2(n16129), .A(n10168), .ZN(n16257) );
  NAND2_X1 U19221 ( .A1(n16131), .A2(n16130), .ZN(n16132) );
  XNOR2_X1 U19222 ( .A(n16133), .B(n16132), .ZN(n16256) );
  AOI22_X1 U19223 ( .A1(n16257), .A2(n16200), .B1(n19175), .B2(n16256), .ZN(
        n16134) );
  INV_X1 U19224 ( .A(n16134), .ZN(n16135) );
  AOI21_X1 U19225 ( .B1(n19171), .B2(n18953), .A(n16135), .ZN(n16136) );
  OAI211_X1 U19226 ( .C1(n19167), .C2(n18947), .A(n16137), .B(n16136), .ZN(
        P2_U3000) );
  AOI22_X1 U19227 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19029), .B1(n16198), 
        .B2(n16138), .ZN(n16145) );
  AND2_X1 U19228 ( .A1(n16139), .A2(n19175), .ZN(n16143) );
  OAI22_X1 U19229 ( .A1(n16141), .A2(n19177), .B1(n16158), .B2(n16140), .ZN(
        n16142) );
  NOR2_X1 U19230 ( .A1(n16143), .A2(n16142), .ZN(n16144) );
  OAI211_X1 U19231 ( .C1(n16146), .C2(n16204), .A(n16145), .B(n16144), .ZN(
        P2_U3001) );
  AOI22_X1 U19232 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19169), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19029), .ZN(n16151) );
  OAI22_X1 U19233 ( .A1(n16148), .A2(n19161), .B1(n16147), .B2(n19177), .ZN(
        n16149) );
  AOI21_X1 U19234 ( .B1(n19171), .B2(n18964), .A(n16149), .ZN(n16150) );
  OAI211_X1 U19235 ( .C1(n19167), .C2(n18962), .A(n16151), .B(n16150), .ZN(
        P2_U3002) );
  AOI22_X1 U19236 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19029), .B1(n16198), 
        .B2(n18974), .ZN(n16169) );
  OAI21_X1 U19237 ( .B1(n16154), .B2(n16153), .A(n16152), .ZN(n16155) );
  INV_X1 U19238 ( .A(n16155), .ZN(n16157) );
  OR2_X1 U19239 ( .A1(n16157), .A2(n16156), .ZN(n16267) );
  OAI22_X1 U19240 ( .A1(n16267), .A2(n19177), .B1(n16158), .B2(n18975), .ZN(
        n16167) );
  NAND2_X1 U19241 ( .A1(n16160), .A2(n16159), .ZN(n16165) );
  INV_X1 U19242 ( .A(n16161), .ZN(n16163) );
  NOR2_X1 U19243 ( .A1(n16163), .A2(n16162), .ZN(n16164) );
  XNOR2_X1 U19244 ( .A(n16165), .B(n16164), .ZN(n16271) );
  NOR2_X1 U19245 ( .A1(n16271), .A2(n19161), .ZN(n16166) );
  NOR2_X1 U19246 ( .A1(n16167), .A2(n16166), .ZN(n16168) );
  OAI211_X1 U19247 ( .C1(n16170), .C2(n16204), .A(n16169), .B(n16168), .ZN(
        P2_U3003) );
  AOI22_X1 U19248 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19029), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19169), .ZN(n16175) );
  OAI22_X1 U19249 ( .A1(n16172), .A2(n19161), .B1(n16171), .B2(n19177), .ZN(
        n16173) );
  AOI21_X1 U19250 ( .B1(n19171), .B2(n18989), .A(n16173), .ZN(n16174) );
  OAI211_X1 U19251 ( .C1(n19167), .C2(n18987), .A(n16175), .B(n16174), .ZN(
        P2_U3004) );
  AOI22_X1 U19252 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19029), .B1(n16198), 
        .B2(n18994), .ZN(n16183) );
  NOR2_X1 U19253 ( .A1(n16176), .A2(n19161), .ZN(n16180) );
  NOR3_X1 U19254 ( .A1(n16178), .A2(n16177), .A3(n19177), .ZN(n16179) );
  AOI211_X1 U19255 ( .C1(n19171), .C2(n16181), .A(n16180), .B(n16179), .ZN(
        n16182) );
  OAI211_X1 U19256 ( .C1(n21003), .C2(n16204), .A(n16183), .B(n16182), .ZN(
        P2_U3005) );
  AOI22_X1 U19257 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19169), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19029), .ZN(n16197) );
  XOR2_X1 U19258 ( .A(n16185), .B(n16184), .Z(n16280) );
  NAND2_X1 U19259 ( .A1(n16187), .A2(n16186), .ZN(n16193) );
  INV_X1 U19260 ( .A(n16188), .ZN(n16189) );
  AOI21_X1 U19261 ( .B1(n16191), .B2(n16190), .A(n16189), .ZN(n16192) );
  XOR2_X1 U19262 ( .A(n16193), .B(n16192), .Z(n16282) );
  AOI22_X1 U19263 ( .A1(n16280), .A2(n16200), .B1(n16282), .B2(n19175), .ZN(
        n16194) );
  INV_X1 U19264 ( .A(n16194), .ZN(n16195) );
  AOI21_X1 U19265 ( .B1(n19171), .B2(n19010), .A(n16195), .ZN(n16196) );
  OAI211_X1 U19266 ( .C1(n19167), .C2(n19005), .A(n16197), .B(n16196), .ZN(
        P2_U3006) );
  AOI22_X1 U19267 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19029), .B1(n16198), 
        .B2(n19034), .ZN(n16203) );
  AOI222_X1 U19268 ( .A1(n16201), .A2(n16200), .B1(n19171), .B2(n19035), .C1(
        n19175), .C2(n16199), .ZN(n16202) );
  OAI211_X1 U19269 ( .C1(n16205), .C2(n16204), .A(n16203), .B(n16202), .ZN(
        P2_U3009) );
  NAND2_X1 U19270 ( .A1(n19029), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16213) );
  AOI21_X1 U19271 ( .B1(n16208), .B2(n16207), .A(n16206), .ZN(n16209) );
  AOI221_X1 U19272 ( .B1(n16221), .B2(n16210), .C1(n16224), .C2(n16210), .A(
        n16209), .ZN(n16211) );
  INV_X1 U19273 ( .A(n16211), .ZN(n16212) );
  NAND2_X1 U19274 ( .A1(n16213), .A2(n16212), .ZN(n16214) );
  AOI21_X1 U19275 ( .B1(n19186), .B2(n16215), .A(n16214), .ZN(n16219) );
  AOI22_X1 U19276 ( .A1(n16217), .A2(n16281), .B1(n19192), .B2(n16216), .ZN(
        n16218) );
  OAI211_X1 U19277 ( .C1(n16305), .C2(n16220), .A(n16219), .B(n16218), .ZN(
        P2_U3022) );
  NOR2_X1 U19278 ( .A1(n19798), .A2(n19045), .ZN(n16226) );
  OAI21_X1 U19279 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n16221), .ZN(n16223) );
  OAI22_X1 U19280 ( .A1(n16224), .A2(n16223), .B1(n16289), .B2(n16222), .ZN(
        n16225) );
  AOI211_X1 U19281 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n16227), .A(
        n16226), .B(n16225), .ZN(n16233) );
  INV_X1 U19282 ( .A(n16228), .ZN(n16231) );
  INV_X1 U19283 ( .A(n16229), .ZN(n16230) );
  AOI22_X1 U19284 ( .A1(n16231), .A2(n19187), .B1(n19192), .B2(n16230), .ZN(
        n16232) );
  OAI211_X1 U19285 ( .C1(n19196), .C2(n16234), .A(n16233), .B(n16232), .ZN(
        P2_U3023) );
  NOR2_X1 U19286 ( .A1(n19783), .A2(n19045), .ZN(n16239) );
  INV_X1 U19287 ( .A(n16235), .ZN(n16237) );
  OAI22_X1 U19288 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16237), .B1(
        n16236), .B2(n16289), .ZN(n16238) );
  AOI211_X1 U19289 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16240), .A(
        n16239), .B(n16238), .ZN(n16244) );
  AOI22_X1 U19290 ( .A1(n16242), .A2(n16281), .B1(n19192), .B2(n16241), .ZN(
        n16243) );
  OAI211_X1 U19291 ( .C1(n16245), .C2(n16305), .A(n16244), .B(n16243), .ZN(
        P2_U3031) );
  INV_X1 U19292 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19781) );
  AOI21_X1 U19293 ( .B1(n16248), .B2(n16247), .A(n16246), .ZN(n19092) );
  NOR3_X1 U19294 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16250), .A3(
        n16249), .ZN(n16255) );
  AOI21_X1 U19295 ( .B1(n16253), .B2(n16252), .A(n16251), .ZN(n16254) );
  AOI211_X1 U19296 ( .C1(n19186), .C2(n19092), .A(n16255), .B(n16254), .ZN(
        n16259) );
  AOI222_X1 U19297 ( .A1(n16257), .A2(n16281), .B1(n19187), .B2(n16256), .C1(
        n19192), .C2(n18953), .ZN(n16258) );
  OAI211_X1 U19298 ( .C1(n19781), .C2(n19045), .A(n16259), .B(n16258), .ZN(
        P2_U3032) );
  NAND2_X1 U19299 ( .A1(n19029), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n16263) );
  OAI211_X1 U19300 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n16261), .B(n16260), .ZN(
        n16262) );
  OAI211_X1 U19301 ( .C1(n18980), .C2(n16289), .A(n16263), .B(n16262), .ZN(
        n16264) );
  AOI21_X1 U19302 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16265), .A(
        n16264), .ZN(n16270) );
  OAI22_X1 U19303 ( .A1(n16267), .A2(n19196), .B1(n16266), .B2(n18975), .ZN(
        n16268) );
  INV_X1 U19304 ( .A(n16268), .ZN(n16269) );
  OAI211_X1 U19305 ( .C1(n16271), .C2(n16305), .A(n16270), .B(n16269), .ZN(
        P2_U3035) );
  AOI211_X1 U19306 ( .C1(n11696), .C2(n16285), .A(n16273), .B(n16272), .ZN(
        n16279) );
  OR2_X1 U19307 ( .A1(n16274), .A2(n9865), .ZN(n16276) );
  AND2_X1 U19308 ( .A1(n16276), .A2(n10174), .ZN(n19100) );
  NAND2_X1 U19309 ( .A1(n19186), .A2(n19100), .ZN(n16277) );
  OAI21_X1 U19310 ( .B1(n11468), .B2(n19045), .A(n16277), .ZN(n16278) );
  NOR2_X1 U19311 ( .A1(n16279), .A2(n16278), .ZN(n16284) );
  AOI222_X1 U19312 ( .A1(n16282), .A2(n19187), .B1(n19192), .B2(n19010), .C1(
        n16281), .C2(n16280), .ZN(n16283) );
  OAI211_X1 U19313 ( .C1(n16286), .C2(n16285), .A(n16284), .B(n16283), .ZN(
        P2_U3038) );
  OAI21_X1 U19314 ( .B1(n16289), .B2(n16288), .A(n16287), .ZN(n16290) );
  AOI21_X1 U19315 ( .B1(n13296), .B2(n19192), .A(n16290), .ZN(n16291) );
  OAI21_X1 U19316 ( .B1(n16292), .B2(n19196), .A(n16291), .ZN(n16293) );
  AOI21_X1 U19317 ( .B1(n19187), .B2(n16294), .A(n16293), .ZN(n16295) );
  OAI221_X1 U19318 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16298), .C1(
        n16297), .C2(n16296), .A(n16295), .ZN(P2_U3043) );
  INV_X1 U19319 ( .A(n19062), .ZN(n16299) );
  AOI22_X1 U19320 ( .A1(n16300), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19186), .B2(n16299), .ZN(n16308) );
  AND2_X1 U19321 ( .A1(n19029), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19172) );
  NAND2_X1 U19322 ( .A1(n19068), .A2(n16301), .ZN(n16302) );
  NAND2_X1 U19323 ( .A1(n10225), .A2(n16302), .ZN(n19173) );
  OAI21_X1 U19324 ( .B1(n16304), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n16303), .ZN(n19176) );
  OAI22_X1 U19325 ( .A1(n16305), .A2(n19173), .B1(n19196), .B2(n19176), .ZN(
        n16306) );
  AOI211_X1 U19326 ( .C1(n19192), .C2(n19170), .A(n19172), .B(n16306), .ZN(
        n16307) );
  OAI211_X1 U19327 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16309), .A(
        n16308), .B(n16307), .ZN(P2_U3046) );
  INV_X1 U19328 ( .A(n16331), .ZN(n16311) );
  MUX2_X1 U19329 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16310), .S(
        n16311), .Z(n16341) );
  MUX2_X1 U19330 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16312), .S(
        n16311), .Z(n16340) );
  NAND2_X1 U19331 ( .A1(n16331), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n16326) );
  AOI22_X1 U19332 ( .A1(n16315), .A2(n16314), .B1(n11647), .B2(n16313), .ZN(
        n16319) );
  NAND2_X1 U19333 ( .A1(n16317), .A2(n16316), .ZN(n16318) );
  AND2_X1 U19334 ( .A1(n16319), .A2(n16318), .ZN(n19867) );
  AOI22_X1 U19335 ( .A1(n16322), .A2(n16321), .B1(n16320), .B2(n19883), .ZN(
        n16325) );
  OAI21_X1 U19336 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n16323), .ZN(n16324) );
  NAND4_X1 U19337 ( .A1(n16326), .A2(n19867), .A3(n16325), .A4(n16324), .ZN(
        n16339) );
  AND2_X1 U19338 ( .A1(n16340), .A2(n13299), .ZN(n16335) );
  NAND2_X1 U19339 ( .A1(n10893), .A2(n16328), .ZN(n16330) );
  OAI22_X1 U19340 ( .A1(n10893), .A2(n16328), .B1(n16327), .B2(n19861), .ZN(
        n16329) );
  NAND2_X1 U19341 ( .A1(n16330), .A2(n16329), .ZN(n16334) );
  AOI21_X1 U19342 ( .B1(n16332), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16331), .ZN(n16333) );
  OAI211_X1 U19343 ( .C1(n16335), .C2(n19845), .A(n16334), .B(n16333), .ZN(
        n16337) );
  AOI22_X1 U19344 ( .A1(n16341), .A2(n13299), .B1(n16335), .B2(n19845), .ZN(
        n16336) );
  AOI21_X1 U19345 ( .B1(n16337), .B2(n16336), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16338) );
  AOI211_X1 U19346 ( .C1(n16341), .C2(n16340), .A(n16339), .B(n16338), .ZN(
        n16358) );
  AOI211_X1 U19347 ( .C1(n16359), .C2(n16344), .A(n16343), .B(n16342), .ZN(
        n16356) );
  AOI21_X1 U19348 ( .B1(n16358), .B2(n16346), .A(n16345), .ZN(n16351) );
  NOR3_X1 U19349 ( .A1(n16347), .A2(n16349), .A3(n16348), .ZN(n16350) );
  AOI21_X1 U19350 ( .B1(n19878), .B2(n16352), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16354) );
  NAND2_X1 U19351 ( .A1(n19743), .A2(n19876), .ZN(n16353) );
  AOI22_X1 U19352 ( .A1(n19743), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16354), 
        .B2(n16353), .ZN(n16355) );
  OAI211_X1 U19353 ( .C1(n16358), .C2(n16357), .A(n16356), .B(n16355), .ZN(
        P2_U3176) );
  AOI221_X1 U19354 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19884), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n19743), .A(n16359), .ZN(n16360) );
  INV_X1 U19355 ( .A(n16360), .ZN(P2_U3593) );
  AOI22_X1 U19356 ( .A1(n17847), .A2(n18056), .B1(n17767), .B2(n17726), .ZN(
        n17754) );
  NAND2_X1 U19357 ( .A1(n16361), .A2(n17637), .ZN(n17529) );
  XOR2_X1 U19358 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n16374), .Z(
        n16537) );
  NAND2_X1 U19359 ( .A1(n17767), .A2(n16362), .ZN(n16388) );
  NAND2_X1 U19360 ( .A1(n17847), .A2(n16363), .ZN(n16381) );
  AOI21_X1 U19361 ( .B1(n16388), .B2(n16381), .A(n16364), .ZN(n16369) );
  INV_X1 U19362 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16538) );
  OAI221_X1 U19363 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16367), .C1(
        n16538), .C2(n16366), .A(n16365), .ZN(n16368) );
  AOI211_X1 U19364 ( .C1(n17708), .C2(n16537), .A(n16369), .B(n16368), .ZN(
        n16372) );
  NAND2_X1 U19365 ( .A1(n17766), .A2(n16370), .ZN(n16371) );
  OAI211_X1 U19366 ( .C1(n17529), .C2(n16373), .A(n16372), .B(n16371), .ZN(
        P3_U2800) );
  OR2_X1 U19367 ( .A1(n16396), .A2(n16395), .ZN(n16386) );
  INV_X1 U19368 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16548) );
  INV_X1 U19369 ( .A(n16514), .ZN(n16375) );
  AOI21_X1 U19370 ( .B1(n16548), .B2(n16375), .A(n16374), .ZN(n16547) );
  OAI21_X1 U19371 ( .B1(n16376), .B2(n17708), .A(n16547), .ZN(n16377) );
  OAI211_X1 U19372 ( .C1(n16380), .C2(n16379), .A(n16378), .B(n16377), .ZN(
        n16384) );
  NOR2_X1 U19373 ( .A1(n17869), .A2(n16396), .ZN(n16399) );
  NOR2_X1 U19374 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16399), .ZN(
        n16382) );
  INV_X1 U19375 ( .A(n17932), .ZN(n17505) );
  AOI22_X1 U19376 ( .A1(n9766), .A2(n18056), .B1(n17726), .B2(n18094), .ZN(
        n17973) );
  INV_X1 U19377 ( .A(n18054), .ZN(n17990) );
  OAI21_X1 U19378 ( .B1(n18670), .B2(n18838), .A(n18171), .ZN(n18089) );
  AOI22_X1 U19379 ( .A1(n18658), .A2(n17990), .B1(n17921), .B2(n18089), .ZN(
        n18020) );
  AOI21_X1 U19380 ( .B1(n17973), .B2(n18020), .A(n17974), .ZN(n17912) );
  NAND3_X1 U19381 ( .A1(n17922), .A2(n18163), .A3(n17912), .ZN(n17960) );
  NOR2_X1 U19382 ( .A1(n17505), .A2(n17960), .ZN(n17908) );
  NOR2_X1 U19383 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n16389), .ZN(
        n17512) );
  AOI22_X1 U19384 ( .A1(n9732), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n17908), 
        .B2(n17512), .ZN(n16405) );
  AOI21_X1 U19385 ( .B1(n17765), .B2(n16390), .A(n17522), .ZN(n17509) );
  AOI22_X1 U19386 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17679), .B1(
        n17765), .B2(n21105), .ZN(n17508) );
  NOR2_X1 U19387 ( .A1(n17509), .A2(n17508), .ZN(n17507) );
  NAND2_X1 U19388 ( .A1(n16392), .A2(n16391), .ZN(n16393) );
  AOI211_X1 U19389 ( .C1(n17521), .C2(n16394), .A(n17507), .B(n16393), .ZN(
        n16401) );
  OAI21_X1 U19390 ( .B1(n16396), .B2(n16395), .A(n18094), .ZN(n16397) );
  OAI211_X1 U19391 ( .C1(n16399), .C2(n9765), .A(n16398), .B(n16397), .ZN(
        n16400) );
  OAI211_X1 U19392 ( .C1(n16401), .C2(n16400), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18179), .ZN(n16404) );
  NAND4_X1 U19393 ( .A1(n17765), .A2(n17509), .A3(n18184), .A4(n21105), .ZN(
        n16403) );
  NAND3_X1 U19394 ( .A1(n18099), .A2(n17522), .A3(n17508), .ZN(n16402) );
  NAND4_X1 U19395 ( .A1(n16405), .A2(n16404), .A3(n16403), .A4(n16402), .ZN(
        P3_U2834) );
  INV_X1 U19396 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n20937) );
  NOR4_X1 U19397 ( .A1(P3_BE_N_REG_0__SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .A4(n20937), .ZN(n16407) );
  NOR4_X1 U19398 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16406) );
  NAND3_X1 U19399 ( .A1(n16407), .A2(n16406), .A3(U215), .ZN(U213) );
  INV_X1 U19400 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19114) );
  INV_X2 U19401 ( .A(U214), .ZN(n16450) );
  NOR2_X2 U19402 ( .A1(n16450), .A2(n16408), .ZN(n16449) );
  OAI222_X1 U19403 ( .A1(U212), .A2(n19114), .B1(n16445), .B2(n19239), .C1(
        U214), .C2(n16482), .ZN(U216) );
  INV_X1 U19404 ( .A(U212), .ZN(n16448) );
  AOI222_X1 U19405 ( .A1(n16450), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16449), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16448), .C2(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n16409) );
  INV_X1 U19406 ( .A(n16409), .ZN(U217) );
  AOI22_X1 U19407 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16450), .ZN(n16410) );
  OAI21_X1 U19408 ( .B1(n20924), .B2(n16445), .A(n16410), .ZN(U218) );
  INV_X1 U19409 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n19223) );
  AOI22_X1 U19410 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16450), .ZN(n16411) );
  OAI21_X1 U19411 ( .B1(n19223), .B2(n16445), .A(n16411), .ZN(U219) );
  INV_X1 U19412 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16413) );
  AOI22_X1 U19413 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16450), .ZN(n16412) );
  OAI21_X1 U19414 ( .B1(n16413), .B2(n16445), .A(n16412), .ZN(U220) );
  INV_X1 U19415 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16415) );
  AOI22_X1 U19416 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16450), .ZN(n16414) );
  OAI21_X1 U19417 ( .B1(n16415), .B2(n16445), .A(n16414), .ZN(U221) );
  INV_X1 U19418 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n16416) );
  INV_X1 U19419 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20912) );
  OAI222_X1 U19420 ( .A1(U214), .A2(n16416), .B1(n16445), .B2(n20912), .C1(
        U212), .C2(n21025), .ZN(U222) );
  AOI22_X1 U19421 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16450), .ZN(n16417) );
  OAI21_X1 U19422 ( .B1(n14587), .B2(n16445), .A(n16417), .ZN(U223) );
  AOI22_X1 U19423 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16450), .ZN(n16418) );
  OAI21_X1 U19424 ( .B1(n14594), .B2(n16445), .A(n16418), .ZN(U224) );
  INV_X1 U19425 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16420) );
  AOI22_X1 U19426 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16450), .ZN(n16419) );
  OAI21_X1 U19427 ( .B1(n16420), .B2(n16445), .A(n16419), .ZN(U225) );
  INV_X1 U19428 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16422) );
  AOI22_X1 U19429 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16450), .ZN(n16421) );
  OAI21_X1 U19430 ( .B1(n16422), .B2(n16445), .A(n16421), .ZN(U226) );
  INV_X1 U19431 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16424) );
  AOI22_X1 U19432 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16450), .ZN(n16423) );
  OAI21_X1 U19433 ( .B1(n16424), .B2(n16445), .A(n16423), .ZN(U227) );
  INV_X1 U19434 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20921) );
  AOI22_X1 U19435 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16450), .ZN(n16425) );
  OAI21_X1 U19436 ( .B1(n20921), .B2(n16445), .A(n16425), .ZN(U228) );
  INV_X1 U19437 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16427) );
  AOI22_X1 U19438 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16450), .ZN(n16426) );
  OAI21_X1 U19439 ( .B1(n16427), .B2(n16445), .A(n16426), .ZN(U229) );
  AOI22_X1 U19440 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16450), .ZN(n16428) );
  OAI21_X1 U19441 ( .B1(n14611), .B2(n16445), .A(n16428), .ZN(U230) );
  AOI222_X1 U19442 ( .A1(n16450), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n16449), 
        .B2(BUF1_REG_16__SCAN_IN), .C1(n16448), .C2(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n16429) );
  INV_X1 U19443 ( .A(n16429), .ZN(U231) );
  INV_X1 U19444 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n20953) );
  INV_X1 U19445 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n20941) );
  OAI222_X1 U19446 ( .A1(U214), .A2(n20953), .B1(n16445), .B2(n12957), .C1(
        U212), .C2(n20941), .ZN(U232) );
  INV_X1 U19447 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n20811) );
  AOI22_X1 U19448 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16450), .ZN(n16430) );
  OAI21_X1 U19449 ( .B1(n20811), .B2(U212), .A(n16430), .ZN(U233) );
  INV_X1 U19450 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n20919) );
  AOI22_X1 U19451 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16450), .ZN(n16431) );
  OAI21_X1 U19452 ( .B1(n20919), .B2(U212), .A(n16431), .ZN(U234) );
  INV_X1 U19453 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16462) );
  AOI22_X1 U19454 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16450), .ZN(n16432) );
  OAI21_X1 U19455 ( .B1(n16462), .B2(U212), .A(n16432), .ZN(U235) );
  INV_X1 U19456 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16461) );
  AOI22_X1 U19457 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16450), .ZN(n16433) );
  OAI21_X1 U19458 ( .B1(n16461), .B2(U212), .A(n16433), .ZN(U236) );
  INV_X1 U19459 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16435) );
  AOI22_X1 U19460 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16450), .ZN(n16434) );
  OAI21_X1 U19461 ( .B1(n16435), .B2(n16445), .A(n16434), .ZN(U237) );
  INV_X1 U19462 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16459) );
  AOI22_X1 U19463 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16450), .ZN(n16436) );
  OAI21_X1 U19464 ( .B1(n16459), .B2(U212), .A(n16436), .ZN(U238) );
  AOI22_X1 U19465 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16450), .ZN(n16437) );
  OAI21_X1 U19466 ( .B1(n16438), .B2(n16445), .A(n16437), .ZN(U239) );
  INV_X1 U19467 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16457) );
  AOI22_X1 U19468 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16450), .ZN(n16439) );
  OAI21_X1 U19469 ( .B1(n16457), .B2(U212), .A(n16439), .ZN(U240) );
  AOI222_X1 U19470 ( .A1(n16450), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n16449), 
        .B2(BUF1_REG_6__SCAN_IN), .C1(n16448), .C2(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n16440) );
  INV_X1 U19471 ( .A(n16440), .ZN(U241) );
  INV_X1 U19472 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16456) );
  AOI22_X1 U19473 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16450), .ZN(n16441) );
  OAI21_X1 U19474 ( .B1(n16456), .B2(U212), .A(n16441), .ZN(U242) );
  INV_X1 U19475 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16443) );
  AOI22_X1 U19476 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16450), .ZN(n16442) );
  OAI21_X1 U19477 ( .B1(n16443), .B2(n16445), .A(n16442), .ZN(U243) );
  INV_X1 U19478 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n20043) );
  INV_X1 U19479 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20902) );
  INV_X1 U19480 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16454) );
  OAI222_X1 U19481 ( .A1(U214), .A2(n20043), .B1(n16445), .B2(n20902), .C1(
        U212), .C2(n16454), .ZN(U244) );
  AOI22_X1 U19482 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16448), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16450), .ZN(n16444) );
  OAI21_X1 U19483 ( .B1(n16446), .B2(n16445), .A(n16444), .ZN(U245) );
  INV_X1 U19484 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16452) );
  AOI22_X1 U19485 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16449), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16450), .ZN(n16447) );
  OAI21_X1 U19486 ( .B1(n16452), .B2(U212), .A(n16447), .ZN(U246) );
  AOI222_X1 U19487 ( .A1(n16450), .A2(P1_DATAO_REG_0__SCAN_IN), .B1(n16449), 
        .B2(BUF1_REG_0__SCAN_IN), .C1(n16448), .C2(P2_DATAO_REG_0__SCAN_IN), 
        .ZN(n16451) );
  INV_X1 U19488 ( .A(n16451), .ZN(U247) );
  INV_X1 U19489 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n20958) );
  INV_X1 U19490 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18200) );
  AOI22_X1 U19491 ( .A1(n16481), .A2(n20958), .B1(n18200), .B2(U215), .ZN(U251) );
  INV_X1 U19492 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18209) );
  AOI22_X1 U19493 ( .A1(n16481), .A2(n16452), .B1(n18209), .B2(U215), .ZN(U252) );
  INV_X1 U19494 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16453) );
  AOI22_X1 U19495 ( .A1(n16481), .A2(n16453), .B1(n18213), .B2(U215), .ZN(U253) );
  INV_X1 U19496 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18218) );
  AOI22_X1 U19497 ( .A1(n16481), .A2(n16454), .B1(n18218), .B2(U215), .ZN(U254) );
  INV_X1 U19498 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16455) );
  INV_X1 U19499 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18223) );
  AOI22_X1 U19500 ( .A1(n16481), .A2(n16455), .B1(n18223), .B2(U215), .ZN(U255) );
  INV_X1 U19501 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n20847) );
  AOI22_X1 U19502 ( .A1(n16481), .A2(n16456), .B1(n20847), .B2(U215), .ZN(U256) );
  INV_X1 U19503 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n19134) );
  INV_X1 U19504 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18231) );
  AOI22_X1 U19505 ( .A1(n16473), .A2(n19134), .B1(n18231), .B2(U215), .ZN(U257) );
  INV_X1 U19506 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18237) );
  AOI22_X1 U19507 ( .A1(n16481), .A2(n16457), .B1(n18237), .B2(U215), .ZN(U258) );
  INV_X1 U19508 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16458) );
  AOI22_X1 U19509 ( .A1(n16473), .A2(n16458), .B1(n17482), .B2(U215), .ZN(U259) );
  INV_X1 U19510 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U19511 ( .A1(n16481), .A2(n16459), .B1(n17484), .B2(U215), .ZN(U260) );
  INV_X1 U19512 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16460) );
  INV_X1 U19513 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17486) );
  AOI22_X1 U19514 ( .A1(n16473), .A2(n16460), .B1(n17486), .B2(U215), .ZN(U261) );
  INV_X1 U19515 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17488) );
  AOI22_X1 U19516 ( .A1(n16481), .A2(n16461), .B1(n17488), .B2(U215), .ZN(U262) );
  INV_X1 U19517 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17491) );
  AOI22_X1 U19518 ( .A1(n16473), .A2(n16462), .B1(n17491), .B2(U215), .ZN(U263) );
  INV_X1 U19519 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n16463) );
  AOI22_X1 U19520 ( .A1(n16481), .A2(n20919), .B1(n16463), .B2(U215), .ZN(U264) );
  INV_X1 U19521 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U19522 ( .A1(n16473), .A2(n20811), .B1(n17496), .B2(U215), .ZN(U265) );
  INV_X1 U19523 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n16464) );
  AOI22_X1 U19524 ( .A1(n16481), .A2(n20941), .B1(n16464), .B2(U215), .ZN(U266) );
  INV_X1 U19525 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n21032) );
  INV_X1 U19526 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n16465) );
  AOI22_X1 U19527 ( .A1(n16473), .A2(n21032), .B1(n16465), .B2(U215), .ZN(U267) );
  OAI22_X1 U19528 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16481), .ZN(n16466) );
  INV_X1 U19529 ( .A(n16466), .ZN(U268) );
  OAI22_X1 U19530 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16481), .ZN(n16467) );
  INV_X1 U19531 ( .A(n16467), .ZN(U269) );
  OAI22_X1 U19532 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16473), .ZN(n16468) );
  INV_X1 U19533 ( .A(n16468), .ZN(U270) );
  OAI22_X1 U19534 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16481), .ZN(n16469) );
  INV_X1 U19535 ( .A(n16469), .ZN(U271) );
  OAI22_X1 U19536 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16473), .ZN(n16470) );
  INV_X1 U19537 ( .A(n16470), .ZN(U272) );
  INV_X1 U19538 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n16471) );
  INV_X1 U19539 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18233) );
  AOI22_X1 U19540 ( .A1(n16473), .A2(n16471), .B1(n18233), .B2(U215), .ZN(U273) );
  OAI22_X1 U19541 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16481), .ZN(n16472) );
  INV_X1 U19542 ( .A(n16472), .ZN(U274) );
  OAI22_X1 U19543 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16473), .ZN(n16474) );
  INV_X1 U19544 ( .A(n16474), .ZN(U275) );
  OAI22_X1 U19545 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16481), .ZN(n16475) );
  INV_X1 U19546 ( .A(n16475), .ZN(U276) );
  OAI22_X1 U19547 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16481), .ZN(n16476) );
  INV_X1 U19548 ( .A(n16476), .ZN(U277) );
  OAI22_X1 U19549 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16481), .ZN(n16477) );
  INV_X1 U19550 ( .A(n16477), .ZN(U278) );
  INV_X1 U19551 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16478) );
  INV_X1 U19552 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19222) );
  AOI22_X1 U19553 ( .A1(n16481), .A2(n16478), .B1(n19222), .B2(U215), .ZN(U279) );
  INV_X1 U19554 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n16479) );
  AOI22_X1 U19555 ( .A1(n16481), .A2(n16479), .B1(n17248), .B2(U215), .ZN(U280) );
  INV_X1 U19556 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n17239) );
  AOI22_X1 U19557 ( .A1(n16481), .A2(n16480), .B1(n17239), .B2(U215), .ZN(U281) );
  INV_X1 U19558 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19237) );
  AOI22_X1 U19559 ( .A1(n16481), .A2(n19114), .B1(n19237), .B2(U215), .ZN(U282) );
  INV_X1 U19560 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17391) );
  AOI222_X1 U19561 ( .A1(n19114), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16482), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n17391), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16483) );
  INV_X2 U19562 ( .A(n16485), .ZN(n16484) );
  INV_X1 U19563 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n21019) );
  INV_X1 U19564 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19775) );
  AOI22_X1 U19565 ( .A1(n16484), .A2(n21019), .B1(n19775), .B2(n16485), .ZN(
        U347) );
  INV_X1 U19566 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18752) );
  INV_X1 U19567 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19774) );
  AOI22_X1 U19568 ( .A1(n16484), .A2(n18752), .B1(n19774), .B2(n16485), .ZN(
        U348) );
  INV_X1 U19569 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n20954) );
  INV_X1 U19570 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20982) );
  AOI22_X1 U19571 ( .A1(n16484), .A2(n20954), .B1(n20982), .B2(n16485), .ZN(
        U349) );
  INV_X1 U19572 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20855) );
  INV_X1 U19573 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19772) );
  AOI22_X1 U19574 ( .A1(n16484), .A2(n20855), .B1(n19772), .B2(n16485), .ZN(
        U350) );
  INV_X1 U19575 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18749) );
  INV_X1 U19576 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19770) );
  AOI22_X1 U19577 ( .A1(n16484), .A2(n18749), .B1(n19770), .B2(n16485), .ZN(
        U351) );
  INV_X1 U19578 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18746) );
  INV_X1 U19579 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19768) );
  AOI22_X1 U19580 ( .A1(n16484), .A2(n18746), .B1(n19768), .B2(n16485), .ZN(
        U352) );
  INV_X1 U19581 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18745) );
  INV_X1 U19582 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19767) );
  AOI22_X1 U19583 ( .A1(n16484), .A2(n18745), .B1(n19767), .B2(n16485), .ZN(
        U353) );
  INV_X1 U19584 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18743) );
  INV_X1 U19585 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19765) );
  AOI22_X1 U19586 ( .A1(n16484), .A2(n18743), .B1(n19765), .B2(n16485), .ZN(
        U354) );
  INV_X1 U19587 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18792) );
  INV_X1 U19588 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20956) );
  AOI22_X1 U19589 ( .A1(n16484), .A2(n18792), .B1(n20956), .B2(n16485), .ZN(
        U355) );
  INV_X1 U19590 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18790) );
  INV_X1 U19591 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19811) );
  AOI22_X1 U19592 ( .A1(n16484), .A2(n18790), .B1(n19811), .B2(n16485), .ZN(
        U356) );
  INV_X1 U19593 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18787) );
  INV_X1 U19594 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19809) );
  AOI22_X1 U19595 ( .A1(n16484), .A2(n18787), .B1(n19809), .B2(n16485), .ZN(
        U357) );
  INV_X1 U19596 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18786) );
  INV_X1 U19597 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19806) );
  AOI22_X1 U19598 ( .A1(n16484), .A2(n18786), .B1(n19806), .B2(n16485), .ZN(
        U358) );
  INV_X1 U19599 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18784) );
  INV_X1 U19600 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n21007) );
  AOI22_X1 U19601 ( .A1(n16484), .A2(n18784), .B1(n21007), .B2(n16485), .ZN(
        U359) );
  INV_X1 U19602 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18782) );
  INV_X1 U19603 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19803) );
  AOI22_X1 U19604 ( .A1(n16484), .A2(n18782), .B1(n19803), .B2(n16485), .ZN(
        U360) );
  INV_X1 U19605 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18780) );
  INV_X1 U19606 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19801) );
  AOI22_X1 U19607 ( .A1(n16484), .A2(n18780), .B1(n19801), .B2(n16485), .ZN(
        U361) );
  INV_X1 U19608 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18777) );
  INV_X1 U19609 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19799) );
  AOI22_X1 U19610 ( .A1(n16484), .A2(n18777), .B1(n19799), .B2(n16485), .ZN(
        U362) );
  INV_X1 U19611 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18776) );
  INV_X1 U19612 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19797) );
  AOI22_X1 U19613 ( .A1(n16484), .A2(n18776), .B1(n19797), .B2(n16485), .ZN(
        U363) );
  INV_X1 U19614 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18773) );
  INV_X1 U19615 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19795) );
  AOI22_X1 U19616 ( .A1(n16484), .A2(n18773), .B1(n19795), .B2(n16485), .ZN(
        U364) );
  INV_X1 U19617 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18741) );
  INV_X1 U19618 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19764) );
  AOI22_X1 U19619 ( .A1(n16484), .A2(n18741), .B1(n19764), .B2(n16485), .ZN(
        U365) );
  INV_X1 U19620 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18772) );
  INV_X1 U19621 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19793) );
  AOI22_X1 U19622 ( .A1(n16484), .A2(n18772), .B1(n19793), .B2(n16485), .ZN(
        U366) );
  INV_X1 U19623 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18769) );
  INV_X1 U19624 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19791) );
  AOI22_X1 U19625 ( .A1(n16484), .A2(n18769), .B1(n19791), .B2(n16485), .ZN(
        U367) );
  INV_X1 U19626 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18768) );
  INV_X1 U19627 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20832) );
  AOI22_X1 U19628 ( .A1(n16484), .A2(n18768), .B1(n20832), .B2(n16485), .ZN(
        U368) );
  INV_X1 U19629 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18766) );
  INV_X1 U19630 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U19631 ( .A1(n16484), .A2(n18766), .B1(n19788), .B2(n16485), .ZN(
        U369) );
  INV_X1 U19632 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18764) );
  INV_X1 U19633 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19786) );
  AOI22_X1 U19634 ( .A1(n16484), .A2(n18764), .B1(n19786), .B2(n16485), .ZN(
        U370) );
  INV_X1 U19635 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20829) );
  INV_X1 U19636 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19784) );
  AOI22_X1 U19637 ( .A1(n16484), .A2(n20829), .B1(n19784), .B2(n16485), .ZN(
        U371) );
  INV_X1 U19638 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18760) );
  INV_X1 U19639 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19782) );
  AOI22_X1 U19640 ( .A1(n16484), .A2(n18760), .B1(n19782), .B2(n16485), .ZN(
        U372) );
  INV_X1 U19641 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18759) );
  INV_X1 U19642 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19780) );
  AOI22_X1 U19643 ( .A1(n16484), .A2(n18759), .B1(n19780), .B2(n16485), .ZN(
        U373) );
  INV_X1 U19644 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18757) );
  INV_X1 U19645 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19778) );
  AOI22_X1 U19646 ( .A1(n16484), .A2(n18757), .B1(n19778), .B2(n16485), .ZN(
        U374) );
  INV_X1 U19647 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18755) );
  INV_X1 U19648 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19777) );
  AOI22_X1 U19649 ( .A1(n16484), .A2(n18755), .B1(n19777), .B2(n16485), .ZN(
        U375) );
  INV_X1 U19650 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18739) );
  INV_X1 U19651 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20972) );
  AOI22_X1 U19652 ( .A1(n16484), .A2(n18739), .B1(n20972), .B2(n16485), .ZN(
        U376) );
  INV_X1 U19653 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16486) );
  NOR2_X1 U19654 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18734), .ZN(n18731) );
  OAI22_X1 U19655 ( .A1(n18729), .A2(n18731), .B1(n18734), .B2(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18804) );
  OAI21_X1 U19656 ( .B1(n18734), .B2(n16486), .A(n18804), .ZN(P3_U2633) );
  INV_X1 U19657 ( .A(n18874), .ZN(n16489) );
  INV_X1 U19658 ( .A(n16492), .ZN(n16487) );
  OAI21_X1 U19659 ( .B1(n16487), .B2(n17455), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16488) );
  OAI21_X1 U19660 ( .B1(n16489), .B2(n18859), .A(n16488), .ZN(P3_U2634) );
  INV_X1 U19661 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21050) );
  AOI21_X1 U19662 ( .B1(n18734), .B2(n21050), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16490) );
  AOI22_X1 U19663 ( .A1(n18869), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16490), 
        .B2(n18868), .ZN(P3_U2635) );
  INV_X1 U19664 ( .A(n18804), .ZN(n18807) );
  NOR2_X1 U19665 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n18725) );
  OAI21_X1 U19666 ( .B1(n18725), .B2(BS16), .A(n18807), .ZN(n18805) );
  OAI21_X1 U19667 ( .B1(n18807), .B2(n16513), .A(n18805), .ZN(P3_U2636) );
  AND3_X1 U19668 ( .A1(n18649), .A2(n16492), .A3(n16491), .ZN(n18652) );
  NOR2_X1 U19669 ( .A1(n18652), .A2(n18713), .ZN(n18852) );
  OAI21_X1 U19670 ( .B1(n18852), .B2(n18191), .A(n16493), .ZN(P3_U2637) );
  NOR4_X1 U19671 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16497) );
  NOR4_X1 U19672 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16496) );
  NOR4_X1 U19673 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16495) );
  NOR4_X1 U19674 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16494) );
  NAND4_X1 U19675 ( .A1(n16497), .A2(n16496), .A3(n16495), .A4(n16494), .ZN(
        n16503) );
  NOR4_X1 U19676 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16501) );
  AOI211_X1 U19677 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_16__SCAN_IN), .B(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16500) );
  NOR4_X1 U19678 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n16499) );
  NOR4_X1 U19679 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16498) );
  NAND4_X1 U19680 ( .A1(n16501), .A2(n16500), .A3(n16499), .A4(n16498), .ZN(
        n16502) );
  NOR2_X1 U19681 ( .A1(n16503), .A2(n16502), .ZN(n18846) );
  INV_X1 U19682 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18799) );
  NOR3_X1 U19683 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16505) );
  OAI21_X1 U19684 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16505), .A(n18846), .ZN(
        n16504) );
  OAI21_X1 U19685 ( .B1(n18846), .B2(n18799), .A(n16504), .ZN(P3_U2638) );
  INV_X1 U19686 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18842) );
  INV_X1 U19687 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18806) );
  AOI21_X1 U19688 ( .B1(n18842), .B2(n18806), .A(n16505), .ZN(n16506) );
  INV_X1 U19689 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18796) );
  INV_X1 U19690 ( .A(n18846), .ZN(n18849) );
  AOI22_X1 U19691 ( .A1(n18846), .A2(n16506), .B1(n18796), .B2(n18849), .ZN(
        P3_U2639) );
  INV_X1 U19692 ( .A(n16507), .ZN(n18682) );
  NAND3_X1 U19693 ( .A1(n18859), .A2(n18856), .A3(n16513), .ZN(n18723) );
  NOR2_X2 U19694 ( .A1(n17857), .A2(n18723), .ZN(n16861) );
  NOR2_X1 U19695 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18810), .ZN(n18548) );
  NAND2_X1 U19696 ( .A1(n18718), .A2(n18548), .ZN(n18711) );
  OAI211_X1 U19697 ( .C1(n18854), .C2(n18855), .A(n18707), .B(n16513), .ZN(
        n18706) );
  INV_X1 U19698 ( .A(n18706), .ZN(n16509) );
  AOI211_X4 U19699 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18855), .A(n16509), .B(
        n16512), .ZN(n16882) );
  INV_X1 U19700 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18793) );
  INV_X1 U19701 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18785) );
  INV_X1 U19702 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18783) );
  INV_X1 U19703 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18779) );
  INV_X1 U19704 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18771) );
  INV_X1 U19705 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18767) );
  INV_X1 U19706 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18754) );
  INV_X1 U19707 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20903) );
  INV_X1 U19708 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18744) );
  NAND3_X1 U19709 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16833) );
  NOR2_X1 U19710 ( .A1(n18744), .A2(n16833), .ZN(n16814) );
  NAND2_X1 U19711 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16814), .ZN(n16787) );
  NAND2_X1 U19712 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16778) );
  NOR3_X1 U19713 ( .A1(n20903), .A2(n16787), .A3(n16778), .ZN(n16739) );
  INV_X1 U19714 ( .A(n16739), .ZN(n16751) );
  INV_X1 U19715 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18753) );
  INV_X1 U19716 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18751) );
  NOR4_X1 U19717 ( .A1(n18754), .A2(n16751), .A3(n18753), .A4(n18751), .ZN(
        n16733) );
  AND2_X1 U19718 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16733), .ZN(n16710) );
  NAND3_X1 U19719 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16710), .ZN(n16711) );
  NAND2_X1 U19720 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16685) );
  NOR2_X1 U19721 ( .A1(n16711), .A2(n16685), .ZN(n16672) );
  NAND2_X1 U19722 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16672), .ZN(n16650) );
  NOR2_X1 U19723 ( .A1(n18767), .A2(n16650), .ZN(n16652) );
  NAND2_X1 U19724 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16652), .ZN(n16642) );
  NOR2_X1 U19725 ( .A1(n18771), .A2(n16642), .ZN(n16619) );
  INV_X1 U19726 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18778) );
  NAND2_X1 U19727 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n16625) );
  NOR2_X1 U19728 ( .A1(n18778), .A2(n16625), .ZN(n16592) );
  NAND2_X1 U19729 ( .A1(n16619), .A2(n16592), .ZN(n16609) );
  NOR2_X1 U19730 ( .A1(n18779), .A2(n16609), .ZN(n16593) );
  NAND2_X1 U19731 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16593), .ZN(n16587) );
  NOR2_X1 U19732 ( .A1(n18783), .A2(n16587), .ZN(n16526) );
  NAND2_X1 U19733 ( .A1(n16855), .A2(n16526), .ZN(n16570) );
  NOR2_X1 U19734 ( .A1(n18785), .A2(n16570), .ZN(n16557) );
  NAND3_X1 U19735 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(n16557), .ZN(n16528) );
  NOR3_X1 U19736 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18793), .A3(n16528), 
        .ZN(n16510) );
  AOI21_X1 U19737 ( .B1(n16882), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16510), .ZN(
        n16533) );
  NAND2_X1 U19738 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18855), .ZN(n16511) );
  AOI211_X4 U19739 ( .C1(n16513), .C2(n18707), .A(n16512), .B(n16511), .ZN(
        n16881) );
  NOR3_X1 U19740 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16851) );
  NAND2_X1 U19741 ( .A1(n16851), .A2(n16847), .ZN(n16846) );
  NOR2_X1 U19742 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16846), .ZN(n16826) );
  NAND2_X1 U19743 ( .A1(n16826), .A2(n16822), .ZN(n16821) );
  INV_X1 U19744 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17197) );
  NAND2_X1 U19745 ( .A1(n16804), .A2(n17197), .ZN(n16794) );
  INV_X1 U19746 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16766) );
  NAND2_X1 U19747 ( .A1(n16777), .A2(n16766), .ZN(n16764) );
  INV_X1 U19748 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16747) );
  NAND2_X1 U19749 ( .A1(n16757), .A2(n16747), .ZN(n16746) );
  NAND2_X1 U19750 ( .A1(n16730), .A2(n17083), .ZN(n16727) );
  NAND2_X1 U19751 ( .A1(n16709), .A2(n21047), .ZN(n16703) );
  NAND2_X1 U19752 ( .A1(n16684), .A2(n16681), .ZN(n16680) );
  NAND2_X1 U19753 ( .A1(n16662), .A2(n16661), .ZN(n16658) );
  INV_X1 U19754 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16981) );
  NAND2_X1 U19755 ( .A1(n16639), .A2(n16981), .ZN(n16633) );
  NOR2_X1 U19756 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16633), .ZN(n16620) );
  INV_X1 U19757 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16890) );
  NAND2_X1 U19758 ( .A1(n16620), .A2(n16890), .ZN(n16615) );
  NOR2_X1 U19759 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16615), .ZN(n16588) );
  NAND2_X1 U19760 ( .A1(n16588), .A2(n16888), .ZN(n16578) );
  NOR2_X1 U19761 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16578), .ZN(n16577) );
  INV_X1 U19762 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16935) );
  NAND2_X1 U19763 ( .A1(n16577), .A2(n16935), .ZN(n16573) );
  NOR2_X1 U19764 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16573), .ZN(n16558) );
  INV_X1 U19765 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16929) );
  NAND2_X1 U19766 ( .A1(n16558), .A2(n16929), .ZN(n16535) );
  NOR2_X1 U19767 ( .A1(n16880), .A2(n16535), .ZN(n16542) );
  INV_X1 U19768 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16896) );
  INV_X1 U19769 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16566) );
  INV_X1 U19770 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20973) );
  NAND2_X1 U19771 ( .A1(n9857), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17543) );
  NOR2_X1 U19772 ( .A1(n9994), .A2(n17543), .ZN(n16520) );
  INV_X1 U19773 ( .A(n16520), .ZN(n16519) );
  NOR2_X1 U19774 ( .A1(n17545), .A2(n16519), .ZN(n17502) );
  INV_X1 U19775 ( .A(n17502), .ZN(n16517) );
  NOR2_X1 U19776 ( .A1(n20973), .A2(n16517), .ZN(n16516) );
  NAND2_X1 U19777 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16516), .ZN(
        n16515) );
  AOI21_X1 U19778 ( .B1(n16566), .B2(n16515), .A(n16514), .ZN(n17504) );
  OAI21_X1 U19779 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16516), .A(
        n16515), .ZN(n17519) );
  INV_X1 U19780 ( .A(n17519), .ZN(n16569) );
  AOI21_X1 U19781 ( .B1(n20973), .B2(n16517), .A(n16516), .ZN(n17537) );
  INV_X1 U19782 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17556) );
  NOR2_X1 U19783 ( .A1(n17556), .A2(n16519), .ZN(n16518) );
  OAI21_X1 U19784 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16518), .A(
        n16517), .ZN(n17547) );
  INV_X1 U19785 ( .A(n17547), .ZN(n16591) );
  AOI22_X1 U19786 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16519), .B1(
        n16520), .B2(n17556), .ZN(n17564) );
  INV_X1 U19787 ( .A(n17564), .ZN(n16603) );
  AOI21_X1 U19788 ( .B1(n9994), .B2(n17543), .A(n16520), .ZN(n17565) );
  INV_X1 U19789 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17597) );
  OR2_X1 U19790 ( .A1(n17585), .A2(n17848), .ZN(n16523) );
  NOR2_X1 U19791 ( .A1(n17597), .A2(n16523), .ZN(n16521) );
  OAI21_X1 U19792 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16521), .A(
        n17543), .ZN(n16522) );
  INV_X1 U19793 ( .A(n16522), .ZN(n17584) );
  XNOR2_X1 U19794 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n16523), .ZN(
        n17593) );
  NAND3_X1 U19795 ( .A1(n17640), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16673) );
  NOR2_X1 U19796 ( .A1(n9860), .A2(n16673), .ZN(n17582) );
  OAI21_X1 U19797 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17582), .A(
        n16523), .ZN(n16524) );
  INV_X1 U19798 ( .A(n16524), .ZN(n17612) );
  NOR2_X1 U19799 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17848), .ZN(
        n16862) );
  NAND2_X1 U19800 ( .A1(n17640), .A2(n16862), .ZN(n16674) );
  NOR2_X1 U19801 ( .A1(n16637), .A2(n16841), .ZN(n16630) );
  NOR2_X1 U19802 ( .A1(n17593), .A2(n16630), .ZN(n16629) );
  NOR2_X1 U19803 ( .A1(n16629), .A2(n16841), .ZN(n16622) );
  NOR2_X1 U19804 ( .A1(n16621), .A2(n16841), .ZN(n16611) );
  NOR2_X1 U19805 ( .A1(n17565), .A2(n16611), .ZN(n16610) );
  NOR2_X1 U19806 ( .A1(n16610), .A2(n16841), .ZN(n16602) );
  NOR2_X1 U19807 ( .A1(n16601), .A2(n16841), .ZN(n16590) );
  NOR2_X1 U19808 ( .A1(n16591), .A2(n16590), .ZN(n16589) );
  NOR2_X1 U19809 ( .A1(n16589), .A2(n16841), .ZN(n16580) );
  NOR2_X1 U19810 ( .A1(n16579), .A2(n16841), .ZN(n16568) );
  NOR2_X1 U19811 ( .A1(n16569), .A2(n16568), .ZN(n16567) );
  NOR2_X1 U19812 ( .A1(n16567), .A2(n16841), .ZN(n16560) );
  NOR2_X1 U19813 ( .A1(n16559), .A2(n16841), .ZN(n16546) );
  NOR2_X1 U19814 ( .A1(n16545), .A2(n16841), .ZN(n16536) );
  NAND2_X1 U19815 ( .A1(n16525), .A2(n16861), .ZN(n16871) );
  NOR3_X1 U19816 ( .A1(n16537), .A2(n16536), .A3(n16871), .ZN(n16531) );
  NAND2_X1 U19817 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .ZN(n16527) );
  OR2_X1 U19818 ( .A1(n16874), .A2(n16526), .ZN(n16586) );
  NAND2_X1 U19819 ( .A1(n16884), .A2(n16586), .ZN(n16583) );
  AOI221_X1 U19820 ( .B1(n18785), .B2(n16855), .C1(n16527), .C2(n16855), .A(
        n16583), .ZN(n16556) );
  NOR2_X1 U19821 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16528), .ZN(n16540) );
  INV_X1 U19822 ( .A(n16540), .ZN(n16529) );
  AOI21_X1 U19823 ( .B1(n16556), .B2(n16529), .A(n21051), .ZN(n16530) );
  AOI211_X1 U19824 ( .C1(n16542), .C2(n16896), .A(n16531), .B(n16530), .ZN(
        n16532) );
  OAI211_X1 U19825 ( .C1(n16534), .C2(n16870), .A(n16533), .B(n16532), .ZN(
        P3_U2640) );
  NAND2_X1 U19826 ( .A1(n16881), .A2(n16535), .ZN(n16552) );
  XOR2_X1 U19827 ( .A(n16537), .B(n16536), .Z(n16541) );
  OAI22_X1 U19828 ( .A1(n16556), .A2(n18793), .B1(n16538), .B2(n16870), .ZN(
        n16539) );
  AOI211_X1 U19829 ( .C1(n16541), .C2(n16861), .A(n16540), .B(n16539), .ZN(
        n16544) );
  OAI21_X1 U19830 ( .B1(n16882), .B2(n16542), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16543) );
  OAI211_X1 U19831 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16552), .A(n16544), .B(
        n16543), .ZN(P3_U2641) );
  INV_X1 U19832 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18789) );
  AOI211_X1 U19833 ( .C1(n16547), .C2(n16546), .A(n16545), .B(n18721), .ZN(
        n16551) );
  NAND2_X1 U19834 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16557), .ZN(n16549) );
  OAI22_X1 U19835 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16549), .B1(n16548), 
        .B2(n16870), .ZN(n16550) );
  AOI211_X1 U19836 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16882), .A(n16551), .B(
        n16550), .ZN(n16555) );
  INV_X1 U19837 ( .A(n16552), .ZN(n16553) );
  OAI21_X1 U19838 ( .B1(n16558), .B2(n16929), .A(n16553), .ZN(n16554) );
  OAI211_X1 U19839 ( .C1(n16556), .C2(n18789), .A(n16555), .B(n16554), .ZN(
        P3_U2642) );
  INV_X1 U19840 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18788) );
  AOI22_X1 U19841 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16882), .B1(n16557), 
        .B2(n18788), .ZN(n16565) );
  INV_X1 U19842 ( .A(n16583), .ZN(n16576) );
  OAI21_X1 U19843 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16570), .A(n16576), 
        .ZN(n16563) );
  AOI211_X1 U19844 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16573), .A(n16558), .B(
        n16880), .ZN(n16562) );
  AOI211_X1 U19845 ( .C1(n17504), .C2(n16560), .A(n16559), .B(n18721), .ZN(
        n16561) );
  AOI211_X1 U19846 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16563), .A(n16562), 
        .B(n16561), .ZN(n16564) );
  OAI211_X1 U19847 ( .C1(n16566), .C2(n16870), .A(n16565), .B(n16564), .ZN(
        P3_U2643) );
  AOI211_X1 U19848 ( .C1(n16569), .C2(n16568), .A(n16567), .B(n18721), .ZN(
        n16572) );
  OAI22_X1 U19849 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16570), .B1(n16935), 
        .B2(n16873), .ZN(n16571) );
  AOI211_X1 U19850 ( .C1(n16807), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16572), .B(n16571), .ZN(n16575) );
  OAI211_X1 U19851 ( .C1(n16577), .C2(n16935), .A(n16881), .B(n16573), .ZN(
        n16574) );
  OAI211_X1 U19852 ( .C1(n16576), .C2(n18785), .A(n16575), .B(n16574), .ZN(
        P3_U2644) );
  AOI22_X1 U19853 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16807), .B1(
        n16882), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16585) );
  AOI211_X1 U19854 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16578), .A(n16577), .B(
        n16880), .ZN(n16582) );
  AOI211_X1 U19855 ( .C1(n17537), .C2(n16580), .A(n16579), .B(n18721), .ZN(
        n16581) );
  AOI211_X1 U19856 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16583), .A(n16582), 
        .B(n16581), .ZN(n16584) );
  OAI211_X1 U19857 ( .C1(n16587), .C2(n16586), .A(n16585), .B(n16584), .ZN(
        P3_U2645) );
  OR2_X1 U19858 ( .A1(n16880), .A2(n16588), .ZN(n16600) );
  AOI21_X1 U19859 ( .B1(n16881), .B2(n16588), .A(n16882), .ZN(n16599) );
  AOI211_X1 U19860 ( .C1(n16591), .C2(n16590), .A(n16589), .B(n18721), .ZN(
        n16597) );
  OAI221_X1 U19861 ( .B1(n16874), .B2(n16619), .C1(n16874), .C2(n16592), .A(
        n16884), .ZN(n16614) );
  AOI21_X1 U19862 ( .B1(n16855), .B2(n18779), .A(n16614), .ZN(n16595) );
  NAND2_X1 U19863 ( .A1(n16855), .A2(n16593), .ZN(n16594) );
  INV_X1 U19864 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18781) );
  AOI22_X1 U19865 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16595), .B1(n16594), 
        .B2(n18781), .ZN(n16596) );
  AOI211_X1 U19866 ( .C1(n16807), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16597), .B(n16596), .ZN(n16598) );
  OAI221_X1 U19867 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16600), .C1(n16888), 
        .C2(n16599), .A(n16598), .ZN(P3_U2646) );
  NAND2_X1 U19868 ( .A1(n16855), .A2(n18779), .ZN(n16608) );
  AOI22_X1 U19869 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16807), .B1(
        n16882), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16607) );
  AOI21_X1 U19870 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16615), .A(n16600), .ZN(
        n16605) );
  AOI211_X1 U19871 ( .C1(n16603), .C2(n16602), .A(n16601), .B(n18721), .ZN(
        n16604) );
  AOI211_X1 U19872 ( .C1(n16614), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16605), 
        .B(n16604), .ZN(n16606) );
  OAI211_X1 U19873 ( .C1(n16609), .C2(n16608), .A(n16607), .B(n16606), .ZN(
        P3_U2647) );
  NOR3_X1 U19874 ( .A1(n16874), .A2(n18771), .A3(n16642), .ZN(n16632) );
  NAND2_X1 U19875 ( .A1(n16632), .A2(n18778), .ZN(n16618) );
  AOI211_X1 U19876 ( .C1(n17565), .C2(n16611), .A(n16610), .B(n18721), .ZN(
        n16613) );
  OAI22_X1 U19877 ( .A1(n9994), .A2(n16870), .B1(n16873), .B2(n16890), .ZN(
        n16612) );
  AOI211_X1 U19878 ( .C1(n16614), .C2(P3_REIP_REG_23__SCAN_IN), .A(n16613), 
        .B(n16612), .ZN(n16617) );
  OAI211_X1 U19879 ( .C1(n16620), .C2(n16890), .A(n16881), .B(n16615), .ZN(
        n16616) );
  OAI211_X1 U19880 ( .C1(n16618), .C2(n16625), .A(n16617), .B(n16616), .ZN(
        P3_U2648) );
  AOI22_X1 U19881 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16807), .B1(
        n16882), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16628) );
  OAI21_X1 U19882 ( .B1(n16619), .B2(n16874), .A(n16884), .ZN(n16643) );
  AOI211_X1 U19883 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16633), .A(n16620), .B(
        n16880), .ZN(n16624) );
  AOI211_X1 U19884 ( .C1(n17584), .C2(n16622), .A(n16621), .B(n18721), .ZN(
        n16623) );
  AOI211_X1 U19885 ( .C1(n16643), .C2(P3_REIP_REG_22__SCAN_IN), .A(n16624), 
        .B(n16623), .ZN(n16627) );
  OAI211_X1 U19886 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(P3_REIP_REG_22__SCAN_IN), .A(n16632), .B(n16625), .ZN(n16626) );
  NAND3_X1 U19887 ( .A1(n16628), .A2(n16627), .A3(n16626), .ZN(P3_U2649) );
  AOI22_X1 U19888 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16807), .B1(
        n16882), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16636) );
  INV_X1 U19889 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18774) );
  AOI211_X1 U19890 ( .C1(n17593), .C2(n16630), .A(n16629), .B(n18721), .ZN(
        n16631) );
  AOI221_X1 U19891 ( .B1(n16643), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n16632), 
        .C2(n18774), .A(n16631), .ZN(n16635) );
  OAI211_X1 U19892 ( .C1(n16639), .C2(n16981), .A(n16881), .B(n16633), .ZN(
        n16634) );
  NAND3_X1 U19893 ( .A1(n16636), .A2(n16635), .A3(n16634), .ZN(P3_U2650) );
  AOI211_X1 U19894 ( .C1(n17612), .C2(n16638), .A(n16637), .B(n18721), .ZN(
        n16641) );
  AOI211_X1 U19895 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16658), .A(n16639), .B(
        n16880), .ZN(n16640) );
  AOI211_X1 U19896 ( .C1(n16807), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16641), .B(n16640), .ZN(n16646) );
  NOR2_X1 U19897 ( .A1(n16874), .A2(n16642), .ZN(n16644) );
  OAI21_X1 U19898 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n16644), .A(n16643), 
        .ZN(n16645) );
  OAI211_X1 U19899 ( .C1(n16995), .C2(n16873), .A(n16646), .B(n16645), .ZN(
        P3_U2651) );
  INV_X1 U19900 ( .A(n16673), .ZN(n17618) );
  NAND2_X1 U19901 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17618), .ZN(
        n16666) );
  AOI21_X1 U19902 ( .B1(n16654), .B2(n16666), .A(n17582), .ZN(n17619) );
  NAND2_X1 U19903 ( .A1(n17692), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16648) );
  NOR2_X1 U19904 ( .A1(n17746), .A2(n17848), .ZN(n16798) );
  INV_X1 U19905 ( .A(n16798), .ZN(n16789) );
  NOR2_X1 U19906 ( .A1(n16647), .A2(n16789), .ZN(n16706) );
  INV_X1 U19907 ( .A(n16706), .ZN(n17688) );
  NOR2_X1 U19908 ( .A1(n16648), .A2(n17688), .ZN(n17652) );
  NAND2_X1 U19909 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17652), .ZN(
        n16695) );
  OAI21_X1 U19910 ( .B1(n16695), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16525), .ZN(n16697) );
  INV_X1 U19911 ( .A(n16697), .ZN(n16692) );
  AOI21_X1 U19912 ( .B1(n16525), .B2(n16666), .A(n16692), .ZN(n16649) );
  XNOR2_X1 U19913 ( .A(n17619), .B(n16649), .ZN(n16657) );
  AOI21_X1 U19914 ( .B1(n16855), .B2(n16650), .A(n16868), .ZN(n16678) );
  NOR3_X1 U19915 ( .A1(n16874), .A2(n16650), .A3(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16665) );
  INV_X1 U19916 ( .A(n16665), .ZN(n16651) );
  INV_X1 U19917 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18770) );
  AOI21_X1 U19918 ( .B1(n16678), .B2(n16651), .A(n18770), .ZN(n16656) );
  NAND3_X1 U19919 ( .A1(n16855), .A2(n16652), .A3(n18770), .ZN(n16653) );
  OAI211_X1 U19920 ( .C1(n16654), .C2(n16870), .A(n18179), .B(n16653), .ZN(
        n16655) );
  AOI211_X1 U19921 ( .C1(n16861), .C2(n16657), .A(n16656), .B(n16655), .ZN(
        n16660) );
  OAI211_X1 U19922 ( .C1(n16662), .C2(n16661), .A(n16881), .B(n16658), .ZN(
        n16659) );
  OAI211_X1 U19923 ( .C1(n16661), .C2(n16873), .A(n16660), .B(n16659), .ZN(
        P3_U2652) );
  AOI211_X1 U19924 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16680), .A(n16662), .B(
        n16880), .ZN(n16664) );
  OAI22_X1 U19925 ( .A1(n17635), .A2(n16870), .B1(n16873), .B2(n9971), .ZN(
        n16663) );
  NOR4_X1 U19926 ( .A1(n9732), .A2(n16665), .A3(n16664), .A4(n16663), .ZN(
        n16671) );
  INV_X1 U19927 ( .A(n16667), .ZN(n16669) );
  OAI21_X1 U19928 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17618), .A(
        n16666), .ZN(n17632) );
  INV_X1 U19929 ( .A(n17632), .ZN(n16668) );
  OAI221_X1 U19930 ( .B1(n16669), .B2(n16668), .C1(n16667), .C2(n17632), .A(
        n16861), .ZN(n16670) );
  OAI211_X1 U19931 ( .C1(n16678), .C2(n18767), .A(n16671), .B(n16670), .ZN(
        P3_U2653) );
  AOI21_X1 U19932 ( .B1(n16855), .B2(n16672), .A(P3_REIP_REG_17__SCAN_IN), 
        .ZN(n16677) );
  AND2_X1 U19933 ( .A1(n17640), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16689) );
  OAI21_X1 U19934 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16689), .A(
        n16673), .ZN(n17641) );
  NAND2_X1 U19935 ( .A1(n16525), .A2(n16674), .ZN(n16675) );
  XNOR2_X1 U19936 ( .A(n17641), .B(n16675), .ZN(n16676) );
  OAI22_X1 U19937 ( .A1(n16678), .A2(n16677), .B1(n18721), .B2(n16676), .ZN(
        n16679) );
  AOI211_X1 U19938 ( .C1(n16882), .C2(P3_EBX_REG_17__SCAN_IN), .A(n9732), .B(
        n16679), .ZN(n16683) );
  OAI211_X1 U19939 ( .C1(n16684), .C2(n16681), .A(n16881), .B(n16680), .ZN(
        n16682) );
  OAI211_X1 U19940 ( .C1(n16870), .C2(n9996), .A(n16683), .B(n16682), .ZN(
        P3_U2654) );
  AOI21_X1 U19941 ( .B1(n16855), .B2(n16711), .A(n16868), .ZN(n16719) );
  INV_X1 U19942 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18763) );
  AOI211_X1 U19943 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16703), .A(n16684), .B(
        n16880), .ZN(n16688) );
  INV_X1 U19944 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16690) );
  NOR2_X1 U19945 ( .A1(n16874), .A2(n16711), .ZN(n16698) );
  OAI211_X1 U19946 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16698), .B(n16685), .ZN(n16686) );
  OAI211_X1 U19947 ( .C1(n16690), .C2(n16870), .A(n18179), .B(n16686), .ZN(
        n16687) );
  AOI211_X1 U19948 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16882), .A(n16688), .B(
        n16687), .ZN(n16694) );
  AOI21_X1 U19949 ( .B1(n16690), .B2(n16695), .A(n16689), .ZN(n17653) );
  INV_X1 U19950 ( .A(n17653), .ZN(n16691) );
  OAI221_X1 U19951 ( .B1(n17653), .B2(n16692), .C1(n16691), .C2(n16697), .A(
        n16861), .ZN(n16693) );
  OAI211_X1 U19952 ( .C1(n16719), .C2(n18763), .A(n16694), .B(n16693), .ZN(
        P3_U2655) );
  INV_X1 U19953 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17669) );
  OAI21_X1 U19954 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17652), .A(
        n16695), .ZN(n17666) );
  NAND2_X1 U19955 ( .A1(n16525), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16696) );
  NAND2_X1 U19956 ( .A1(n16861), .A2(n16696), .ZN(n16869) );
  AOI211_X1 U19957 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16525), .A(
        n17666), .B(n16869), .ZN(n16702) );
  INV_X1 U19958 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18762) );
  NOR2_X1 U19959 ( .A1(n18721), .A2(n16697), .ZN(n16699) );
  AOI22_X1 U19960 ( .A1(n16699), .A2(n17666), .B1(n16698), .B2(n18762), .ZN(
        n16700) );
  OAI211_X1 U19961 ( .C1(n18762), .C2(n16719), .A(n16700), .B(n18179), .ZN(
        n16701) );
  AOI211_X1 U19962 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16882), .A(n16702), .B(
        n16701), .ZN(n16705) );
  OAI211_X1 U19963 ( .C1(n16709), .C2(n21047), .A(n16881), .B(n16703), .ZN(
        n16704) );
  OAI211_X1 U19964 ( .C1(n16870), .C2(n17669), .A(n16705), .B(n16704), .ZN(
        P3_U2656) );
  INV_X1 U19965 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18761) );
  INV_X1 U19966 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16872) );
  AND3_X1 U19967 ( .A1(n16872), .A2(n17692), .A3(n16706), .ZN(n16712) );
  NOR2_X1 U19968 ( .A1(n16712), .A2(n16871), .ZN(n16726) );
  INV_X1 U19969 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16707) );
  NAND2_X1 U19970 ( .A1(n17692), .A2(n16706), .ZN(n16720) );
  AOI21_X1 U19971 ( .B1(n16707), .B2(n16720), .A(n17652), .ZN(n17685) );
  INV_X1 U19972 ( .A(n17685), .ZN(n16708) );
  AOI22_X1 U19973 ( .A1(n16882), .A2(P3_EBX_REG_14__SCAN_IN), .B1(n16726), 
        .B2(n16708), .ZN(n16718) );
  AOI211_X1 U19974 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16727), .A(n16709), .B(
        n16880), .ZN(n16716) );
  NAND2_X1 U19975 ( .A1(n16855), .A2(n16710), .ZN(n16723) );
  NAND2_X1 U19976 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16711), .ZN(n16714) );
  OAI211_X1 U19977 ( .C1(n16712), .C2(n16841), .A(n16861), .B(n17685), .ZN(
        n16713) );
  OAI211_X1 U19978 ( .C1(n16723), .C2(n16714), .A(n18179), .B(n16713), .ZN(
        n16715) );
  AOI211_X1 U19979 ( .C1(n16807), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16716), .B(n16715), .ZN(n16717) );
  OAI211_X1 U19980 ( .C1(n18761), .C2(n16719), .A(n16718), .B(n16717), .ZN(
        P3_U2657) );
  NOR2_X1 U19981 ( .A1(n20927), .A2(n17688), .ZN(n16734) );
  OAI21_X1 U19982 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16734), .A(
        n16720), .ZN(n17703) );
  AOI211_X1 U19983 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16525), .A(
        n17703), .B(n16869), .ZN(n16725) );
  INV_X1 U19984 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18758) );
  INV_X1 U19985 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18756) );
  OAI21_X1 U19986 ( .B1(n16733), .B2(n16874), .A(n16884), .ZN(n16745) );
  AOI21_X1 U19987 ( .B1(n16855), .B2(n18756), .A(n16745), .ZN(n16722) );
  AOI21_X1 U19988 ( .B1(n16882), .B2(P3_EBX_REG_13__SCAN_IN), .A(n9732), .ZN(
        n16721) );
  OAI221_X1 U19989 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n16723), .C1(n18758), 
        .C2(n16722), .A(n16721), .ZN(n16724) );
  AOI211_X1 U19990 ( .C1(n16726), .C2(n17703), .A(n16725), .B(n16724), .ZN(
        n16729) );
  OAI211_X1 U19991 ( .C1(n16730), .C2(n17083), .A(n16881), .B(n16727), .ZN(
        n16728) );
  OAI211_X1 U19992 ( .C1(n16870), .C2(n17693), .A(n16729), .B(n16728), .ZN(
        P3_U2658) );
  AOI22_X1 U19993 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16807), .B1(
        n16882), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16738) );
  NOR2_X1 U19994 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16874), .ZN(n16732) );
  AOI211_X1 U19995 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16746), .A(n16730), .B(
        n16880), .ZN(n16731) );
  AOI211_X1 U19996 ( .C1(n16733), .C2(n16732), .A(n9732), .B(n16731), .ZN(
        n16737) );
  AOI21_X1 U19997 ( .B1(n20927), .B2(n17688), .A(n16734), .ZN(n17707) );
  OAI21_X1 U19998 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17688), .A(
        n16525), .ZN(n16742) );
  XNOR2_X1 U19999 ( .A(n17707), .B(n16742), .ZN(n16735) );
  AOI22_X1 U20000 ( .A1(n16861), .A2(n16735), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16745), .ZN(n16736) );
  NAND3_X1 U20001 ( .A1(n16738), .A2(n16737), .A3(n16736), .ZN(P3_U2659) );
  AOI22_X1 U20002 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n16807), .B1(
        n16882), .B2(P3_EBX_REG_11__SCAN_IN), .ZN(n16750) );
  NAND2_X1 U20003 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16740) );
  NAND2_X1 U20004 ( .A1(n16855), .A2(n16739), .ZN(n16767) );
  OAI21_X1 U20005 ( .B1(n16740), .B2(n16767), .A(n18754), .ZN(n16744) );
  OAI221_X1 U20006 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16753), .C1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n16798), .A(n17688), .ZN(
        n17719) );
  NOR2_X1 U20007 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16789), .ZN(
        n16790) );
  AOI211_X1 U20008 ( .C1(n16753), .C2(n16790), .A(n16841), .B(n17719), .ZN(
        n16741) );
  AOI211_X1 U20009 ( .C1(n17719), .C2(n16742), .A(n16741), .B(n18721), .ZN(
        n16743) );
  AOI21_X1 U20010 ( .B1(n16745), .B2(n16744), .A(n16743), .ZN(n16749) );
  OAI211_X1 U20011 ( .C1(n16757), .C2(n16747), .A(n16881), .B(n16746), .ZN(
        n16748) );
  NAND4_X1 U20012 ( .A1(n16750), .A2(n16749), .A3(n18179), .A4(n16748), .ZN(
        P3_U2660) );
  AOI21_X1 U20013 ( .B1(n16855), .B2(n16751), .A(n16868), .ZN(n16779) );
  AOI221_X1 U20014 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .C1(n18753), .C2(n18751), .A(n16767), .ZN(n16752) );
  AOI211_X1 U20015 ( .C1(n16882), .C2(P3_EBX_REG_10__SCAN_IN), .A(n9732), .B(
        n16752), .ZN(n16761) );
  INV_X1 U20016 ( .A(n17746), .ZN(n17757) );
  NAND2_X1 U20017 ( .A1(n17757), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17759) );
  NOR2_X1 U20018 ( .A1(n17848), .A2(n17759), .ZN(n16788) );
  NAND2_X1 U20019 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16788), .ZN(
        n16775) );
  INV_X1 U20020 ( .A(n16775), .ZN(n16763) );
  NAND2_X1 U20021 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16763), .ZN(
        n16762) );
  OAI21_X1 U20022 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16762), .A(
        n16525), .ZN(n16770) );
  INV_X1 U20023 ( .A(n16762), .ZN(n16755) );
  NAND2_X1 U20024 ( .A1(n16753), .A2(n16798), .ZN(n16754) );
  OAI21_X1 U20025 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16755), .A(
        n16754), .ZN(n17733) );
  OAI21_X1 U20026 ( .B1(n16770), .B2(n17733), .A(n16861), .ZN(n16756) );
  AOI21_X1 U20027 ( .B1(n16770), .B2(n17733), .A(n16756), .ZN(n16759) );
  AOI211_X1 U20028 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16764), .A(n16757), .B(
        n16880), .ZN(n16758) );
  AOI211_X1 U20029 ( .C1(n16807), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16759), .B(n16758), .ZN(n16760) );
  OAI211_X1 U20030 ( .C1(n18753), .C2(n16779), .A(n16761), .B(n16760), .ZN(
        P3_U2661) );
  OAI21_X1 U20031 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16763), .A(
        n16762), .ZN(n17747) );
  NAND2_X1 U20032 ( .A1(n16861), .A2(n16841), .ZN(n16865) );
  OAI211_X1 U20033 ( .C1(n16777), .C2(n16766), .A(n16881), .B(n16764), .ZN(
        n16765) );
  OAI211_X1 U20034 ( .C1(n17747), .C2(n16865), .A(n18179), .B(n16765), .ZN(
        n16769) );
  OAI22_X1 U20035 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16767), .B1(n16873), 
        .B2(n16766), .ZN(n16768) );
  AOI211_X1 U20036 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n16807), .A(
        n16769), .B(n16768), .ZN(n16774) );
  NOR2_X1 U20037 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16775), .ZN(
        n16772) );
  INV_X1 U20038 ( .A(n16770), .ZN(n16771) );
  OAI211_X1 U20039 ( .C1(n16772), .C2(n17747), .A(n16771), .B(n16861), .ZN(
        n16773) );
  OAI211_X1 U20040 ( .C1(n16779), .C2(n18751), .A(n16774), .B(n16773), .ZN(
        P3_U2662) );
  OAI21_X1 U20041 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16788), .A(
        n16775), .ZN(n17761) );
  INV_X1 U20042 ( .A(n16862), .ZN(n16831) );
  OAI21_X1 U20043 ( .B1(n16831), .B2(n17759), .A(n16525), .ZN(n16776) );
  XNOR2_X1 U20044 ( .A(n17761), .B(n16776), .ZN(n16786) );
  AOI211_X1 U20045 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16794), .A(n16777), .B(
        n16880), .ZN(n16784) );
  INV_X1 U20046 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17760) );
  INV_X1 U20047 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20850) );
  OAI22_X1 U20048 ( .A1(n17760), .A2(n16870), .B1(n16873), .B2(n20850), .ZN(
        n16783) );
  NAND3_X1 U20049 ( .A1(n16855), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n16814), 
        .ZN(n16803) );
  NOR2_X1 U20050 ( .A1(n16778), .A2(n16803), .ZN(n16781) );
  INV_X1 U20051 ( .A(n16779), .ZN(n16780) );
  MUX2_X1 U20052 ( .A(n16781), .B(n16780), .S(P3_REIP_REG_8__SCAN_IN), .Z(
        n16782) );
  NOR4_X1 U20053 ( .A1(n9732), .A2(n16784), .A3(n16783), .A4(n16782), .ZN(
        n16785) );
  OAI21_X1 U20054 ( .B1(n18721), .B2(n16786), .A(n16785), .ZN(P3_U2663) );
  AOI22_X1 U20055 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16807), .B1(
        n16882), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n16797) );
  NOR2_X1 U20056 ( .A1(n16868), .A2(n16787), .ZN(n16819) );
  NOR2_X1 U20057 ( .A1(n16868), .A2(n16855), .ZN(n16813) );
  AOI21_X1 U20058 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16819), .A(n16813), .ZN(
        n16801) );
  INV_X1 U20059 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18748) );
  NOR2_X1 U20060 ( .A1(n18748), .A2(n16803), .ZN(n16793) );
  INV_X1 U20061 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18750) );
  INV_X1 U20062 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17773) );
  AOI21_X1 U20063 ( .B1(n17773), .B2(n16789), .A(n16788), .ZN(n17779) );
  NOR2_X1 U20064 ( .A1(n16790), .A2(n16841), .ZN(n16809) );
  OAI21_X1 U20065 ( .B1(n17779), .B2(n16809), .A(n16861), .ZN(n16791) );
  AOI21_X1 U20066 ( .B1(n17779), .B2(n16809), .A(n16791), .ZN(n16792) );
  AOI221_X1 U20067 ( .B1(n16801), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n16793), 
        .C2(n18750), .A(n16792), .ZN(n16796) );
  OAI211_X1 U20068 ( .C1(n16804), .C2(n17197), .A(n16881), .B(n16794), .ZN(
        n16795) );
  NAND4_X1 U20069 ( .A1(n16797), .A2(n16796), .A3(n18179), .A4(n16795), .ZN(
        P3_U2664) );
  INV_X1 U20070 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16799) );
  NAND2_X1 U20071 ( .A1(n17790), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16815) );
  AOI21_X1 U20072 ( .B1(n16799), .B2(n16815), .A(n16798), .ZN(n17791) );
  AOI21_X1 U20073 ( .B1(n16525), .B2(n16815), .A(n16869), .ZN(n16800) );
  AOI22_X1 U20074 ( .A1(n16882), .A2(P3_EBX_REG_6__SCAN_IN), .B1(n17791), .B2(
        n16800), .ZN(n16812) );
  INV_X1 U20075 ( .A(n16801), .ZN(n16802) );
  AOI21_X1 U20076 ( .B1(n18748), .B2(n16803), .A(n16802), .ZN(n16806) );
  AOI211_X1 U20077 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16821), .A(n16804), .B(
        n16880), .ZN(n16805) );
  AOI211_X1 U20078 ( .C1(n16807), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16806), .B(n16805), .ZN(n16811) );
  INV_X1 U20079 ( .A(n17791), .ZN(n16808) );
  NAND3_X1 U20080 ( .A1(n16861), .A2(n16809), .A3(n16808), .ZN(n16810) );
  NAND4_X1 U20081 ( .A1(n16812), .A2(n16811), .A3(n18179), .A4(n16810), .ZN(
        P3_U2665) );
  INV_X1 U20082 ( .A(n16813), .ZN(n16883) );
  AOI22_X1 U20083 ( .A1(n16855), .A2(n16814), .B1(P3_REIP_REG_5__SCAN_IN), 
        .B2(n16883), .ZN(n16818) );
  INV_X1 U20084 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16830) );
  NAND2_X1 U20085 ( .A1(n17815), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16839) );
  NOR2_X1 U20086 ( .A1(n16830), .A2(n16839), .ZN(n16825) );
  OAI21_X1 U20087 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16825), .A(
        n16815), .ZN(n17802) );
  INV_X1 U20088 ( .A(n16825), .ZN(n16816) );
  OAI21_X1 U20089 ( .B1(n16816), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16525), .ZN(n16832) );
  XNOR2_X1 U20090 ( .A(n17802), .B(n16832), .ZN(n16817) );
  OAI22_X1 U20091 ( .A1(n16819), .A2(n16818), .B1(n18721), .B2(n16817), .ZN(
        n16820) );
  AOI211_X1 U20092 ( .C1(n16882), .C2(P3_EBX_REG_5__SCAN_IN), .A(n9732), .B(
        n16820), .ZN(n16824) );
  OAI211_X1 U20093 ( .C1(n16826), .C2(n16822), .A(n16881), .B(n16821), .ZN(
        n16823) );
  OAI211_X1 U20094 ( .C1(n16870), .C2(n20943), .A(n16824), .B(n16823), .ZN(
        P3_U2666) );
  AOI21_X1 U20095 ( .B1(n16855), .B2(n16833), .A(n16868), .ZN(n16842) );
  INV_X1 U20096 ( .A(n16865), .ZN(n16829) );
  AOI21_X1 U20097 ( .B1(n16830), .B2(n16839), .A(n16825), .ZN(n17816) );
  AOI211_X1 U20098 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16846), .A(n16826), .B(
        n16880), .ZN(n16828) );
  INV_X1 U20099 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n20813) );
  OAI22_X1 U20100 ( .A1(n16830), .A2(n16870), .B1(n16873), .B2(n20813), .ZN(
        n16827) );
  AOI211_X1 U20101 ( .C1(n16829), .C2(n17816), .A(n16828), .B(n16827), .ZN(
        n16838) );
  NAND2_X1 U20102 ( .A1(n17815), .A2(n16830), .ZN(n17813) );
  OAI22_X1 U20103 ( .A1(n17816), .A2(n16832), .B1(n16831), .B2(n17813), .ZN(
        n16836) );
  NOR3_X1 U20104 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16874), .A3(n16833), .ZN(
        n16835) );
  NAND2_X1 U20105 ( .A1(n18204), .A2(n18873), .ZN(n16853) );
  OAI221_X1 U20106 ( .B1(n16853), .B2(n17118), .C1(n16853), .C2(n18655), .A(
        n18179), .ZN(n16834) );
  AOI211_X1 U20107 ( .C1(n16861), .C2(n16836), .A(n16835), .B(n16834), .ZN(
        n16837) );
  OAI211_X1 U20108 ( .C1(n18744), .C2(n16842), .A(n16838), .B(n16837), .ZN(
        P3_U2667) );
  NAND2_X1 U20109 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16850) );
  INV_X1 U20110 ( .A(n16839), .ZN(n16840) );
  AOI21_X1 U20111 ( .B1(n17826), .B2(n16850), .A(n16840), .ZN(n17830) );
  AOI21_X1 U20112 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n16862), .A(
        n16841), .ZN(n16860) );
  XOR2_X1 U20113 ( .A(n17830), .B(n16860), .Z(n16845) );
  INV_X1 U20114 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18742) );
  NAND2_X1 U20115 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16854) );
  AOI221_X1 U20116 ( .B1(n16874), .B2(n18742), .C1(n16854), .C2(n18742), .A(
        n16842), .ZN(n16844) );
  NOR2_X1 U20117 ( .A1(n21016), .A2(n18666), .ZN(n18664) );
  OAI21_X1 U20118 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18664), .A(
        n17118), .ZN(n18813) );
  OAI22_X1 U20119 ( .A1(n16873), .A2(n16847), .B1(n18813), .B2(n16853), .ZN(
        n16843) );
  AOI211_X1 U20120 ( .C1(n16845), .C2(n16861), .A(n16844), .B(n16843), .ZN(
        n16849) );
  OAI211_X1 U20121 ( .C1(n16851), .C2(n16847), .A(n16881), .B(n16846), .ZN(
        n16848) );
  OAI211_X1 U20122 ( .C1(n16870), .C2(n17826), .A(n16849), .B(n16848), .ZN(
        P3_U2668) );
  OAI21_X1 U20123 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16850), .ZN(n17838) );
  INV_X1 U20124 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17229) );
  INV_X1 U20125 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17223) );
  NAND2_X1 U20126 ( .A1(n17229), .A2(n17223), .ZN(n16852) );
  AOI211_X1 U20127 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16852), .A(n16851), .B(
        n16880), .ZN(n16859) );
  AOI21_X1 U20128 ( .B1(n18826), .B2(n18685), .A(n18664), .ZN(n18822) );
  INV_X1 U20129 ( .A(n16853), .ZN(n18875) );
  AOI22_X1 U20130 ( .A1(n16868), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18822), 
        .B2(n18875), .ZN(n16857) );
  OAI211_X1 U20131 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16855), .B(n16854), .ZN(n16856) );
  OAI211_X1 U20132 ( .C1(n16870), .C2(n17841), .A(n16857), .B(n16856), .ZN(
        n16858) );
  AOI211_X1 U20133 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16882), .A(n16859), .B(
        n16858), .ZN(n16864) );
  OAI211_X1 U20134 ( .C1(n16862), .C2(n17838), .A(n16861), .B(n16860), .ZN(
        n16863) );
  OAI211_X1 U20135 ( .C1(n16865), .C2(n17838), .A(n16864), .B(n16863), .ZN(
        P3_U2669) );
  NOR2_X1 U20136 ( .A1(n17229), .A2(n17223), .ZN(n17219) );
  AOI21_X1 U20137 ( .B1(n17229), .B2(n17223), .A(n17219), .ZN(n16866) );
  INV_X1 U20138 ( .A(n16866), .ZN(n17225) );
  AND2_X1 U20139 ( .A1(n16867), .A2(n18685), .ZN(n18832) );
  AOI22_X1 U20140 ( .A1(n16868), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18832), 
        .B2(n18875), .ZN(n16879) );
  INV_X1 U20141 ( .A(n16869), .ZN(n16877) );
  OAI21_X1 U20142 ( .B1(n16872), .B2(n16871), .A(n16870), .ZN(n16876) );
  OAI22_X1 U20143 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16874), .B1(n16873), 
        .B2(n17223), .ZN(n16875) );
  AOI221_X1 U20144 ( .B1(n16877), .B2(n17848), .C1(n16876), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16875), .ZN(n16878) );
  OAI211_X1 U20145 ( .C1(n16880), .C2(n17225), .A(n16879), .B(n16878), .ZN(
        P3_U2670) );
  NOR2_X1 U20146 ( .A1(n16882), .A2(n16881), .ZN(n16887) );
  AOI22_X1 U20147 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16883), .B1(n18875), 
        .B2(n21016), .ZN(n16886) );
  NAND3_X1 U20148 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18829), .A3(
        n16884), .ZN(n16885) );
  OAI211_X1 U20149 ( .C1(n16887), .C2(n17229), .A(n16886), .B(n16885), .ZN(
        P3_U2671) );
  NOR2_X1 U20150 ( .A1(n16888), .A2(n16940), .ZN(n16892) );
  NAND2_X1 U20151 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16930), .ZN(n16889) );
  NAND2_X1 U20152 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17010), .ZN(n16967) );
  NOR4_X1 U20153 ( .A1(n16929), .A2(n16890), .A3(n16889), .A4(n16967), .ZN(
        n16891) );
  NAND4_X1 U20154 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n16892), .A4(n16891), .ZN(n16895) );
  NAND2_X1 U20155 ( .A1(n17222), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16894) );
  NAND2_X1 U20156 ( .A1(n16923), .A2(n18240), .ZN(n16893) );
  OAI22_X1 U20157 ( .A1(n16923), .A2(n16894), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16893), .ZN(P3_U2672) );
  NAND2_X1 U20158 ( .A1(n16896), .A2(n16895), .ZN(n16897) );
  NAND2_X1 U20159 ( .A1(n16897), .A2(n17222), .ZN(n16922) );
  AOI22_X1 U20160 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9733), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16909) );
  AOI22_X1 U20161 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16908) );
  AOI22_X1 U20162 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17038), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16907) );
  OAI22_X1 U20163 ( .A1(n10275), .A2(n16899), .B1(n17143), .B2(n16898), .ZN(
        n16905) );
  AOI22_X1 U20164 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16903) );
  AOI22_X1 U20165 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16902) );
  AOI22_X1 U20166 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16901) );
  NAND2_X1 U20167 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n16900) );
  NAND4_X1 U20168 ( .A1(n16903), .A2(n16902), .A3(n16901), .A4(n16900), .ZN(
        n16904) );
  AOI211_X1 U20169 ( .C1(n17181), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n16905), .B(n16904), .ZN(n16906) );
  NAND4_X1 U20170 ( .A1(n16909), .A2(n16908), .A3(n16907), .A4(n16906), .ZN(
        n16921) );
  AOI22_X1 U20171 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16919) );
  AOI22_X1 U20172 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16918) );
  AOI22_X1 U20173 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17031), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16917) );
  OAI22_X1 U20174 ( .A1(n10298), .A2(n17068), .B1(n10267), .B2(n17070), .ZN(
        n16915) );
  AOI22_X1 U20175 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20176 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9733), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20177 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16911) );
  NAND2_X1 U20178 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n16910) );
  NAND4_X1 U20179 ( .A1(n16913), .A2(n16912), .A3(n16911), .A4(n16910), .ZN(
        n16914) );
  AOI211_X1 U20180 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n16915), .B(n16914), .ZN(n16916) );
  NAND4_X1 U20181 ( .A1(n16919), .A2(n16918), .A3(n16917), .A4(n16916), .ZN(
        n16926) );
  INV_X1 U20182 ( .A(n17254), .ZN(n16924) );
  NAND3_X1 U20183 ( .A1(n16926), .A2(n16924), .A3(n16925), .ZN(n16920) );
  XOR2_X1 U20184 ( .A(n16921), .B(n16920), .Z(n17240) );
  OAI22_X1 U20185 ( .A1(n16923), .A2(n16922), .B1(n17240), .B2(n17222), .ZN(
        P3_U2673) );
  NAND2_X1 U20186 ( .A1(n16925), .A2(n16924), .ZN(n16927) );
  XNOR2_X1 U20187 ( .A(n16927), .B(n16926), .ZN(n17244) );
  AOI22_X1 U20188 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16928), .B1(n17227), 
        .B2(n17244), .ZN(n16932) );
  NAND4_X1 U20189 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n9828), .A3(n16930), .A4(
        n16929), .ZN(n16931) );
  NAND2_X1 U20190 ( .A1(n16932), .A2(n16931), .ZN(P3_U2674) );
  OAI211_X1 U20191 ( .C1(n17256), .C2(n17255), .A(n17227), .B(n17254), .ZN(
        n16933) );
  OAI221_X1 U20192 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16936), .C1(n16935), 
        .C2(n16934), .A(n16933), .ZN(P3_U2676) );
  AOI21_X1 U20193 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17222), .A(n9828), .ZN(
        n16938) );
  XNOR2_X1 U20194 ( .A(n16937), .B(n16941), .ZN(n17265) );
  OAI22_X1 U20195 ( .A1(n16939), .A2(n16938), .B1(n17222), .B2(n17265), .ZN(
        P3_U2677) );
  NOR2_X1 U20196 ( .A1(n16940), .A2(n16945), .ZN(n16948) );
  AOI21_X1 U20197 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17222), .A(n16948), .ZN(
        n16944) );
  OAI21_X1 U20198 ( .B1(n16943), .B2(n16942), .A(n16941), .ZN(n17269) );
  OAI22_X1 U20199 ( .A1(n9828), .A2(n16944), .B1(n17222), .B2(n17269), .ZN(
        P3_U2678) );
  INV_X1 U20200 ( .A(n16945), .ZN(n16953) );
  AOI21_X1 U20201 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17222), .A(n16953), .ZN(
        n16947) );
  XNOR2_X1 U20202 ( .A(n16946), .B(n16949), .ZN(n17276) );
  OAI22_X1 U20203 ( .A1(n16948), .A2(n16947), .B1(n17222), .B2(n17276), .ZN(
        P3_U2679) );
  AOI21_X1 U20204 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17222), .A(n9842), .ZN(
        n16952) );
  OAI21_X1 U20205 ( .B1(n16951), .B2(n16950), .A(n16949), .ZN(n17279) );
  OAI22_X1 U20206 ( .A1(n16953), .A2(n16952), .B1(n17222), .B2(n17279), .ZN(
        P3_U2680) );
  AOI22_X1 U20207 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16954) );
  OAI21_X1 U20208 ( .B1(n17170), .B2(n17070), .A(n16954), .ZN(n16964) );
  AOI22_X1 U20209 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16961) );
  INV_X1 U20210 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18236) );
  AOI22_X1 U20211 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16955) );
  OAI21_X1 U20212 ( .B1(n10298), .B2(n18236), .A(n16955), .ZN(n16959) );
  AOI22_X1 U20213 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20214 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16956) );
  OAI211_X1 U20215 ( .C1(n17188), .C2(n17068), .A(n16957), .B(n16956), .ZN(
        n16958) );
  AOI211_X1 U20216 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n16959), .B(n16958), .ZN(n16960) );
  OAI211_X1 U20217 ( .C1(n9794), .C2(n16962), .A(n16961), .B(n16960), .ZN(
        n16963) );
  AOI211_X1 U20218 ( .C1(n17173), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n16964), .B(n16963), .ZN(n17284) );
  NAND3_X1 U20219 ( .A1(n16966), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17222), 
        .ZN(n16965) );
  OAI221_X1 U20220 ( .B1(n16966), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17222), 
        .C2(n17284), .A(n16965), .ZN(P3_U2681) );
  NAND2_X1 U20221 ( .A1(n17222), .A2(n16967), .ZN(n16996) );
  AOI22_X1 U20222 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16978) );
  AOI22_X1 U20223 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16968) );
  OAI21_X1 U20224 ( .B1(n17118), .B2(n18281), .A(n16968), .ZN(n16976) );
  OAI22_X1 U20225 ( .A1(n10275), .A2(n21035), .B1(n17143), .B2(n16969), .ZN(
        n16970) );
  AOI21_X1 U20226 ( .B1(n9733), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n16970), .ZN(n16974) );
  AOI22_X1 U20227 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20228 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20229 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17031), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16971) );
  NAND4_X1 U20230 ( .A1(n16974), .A2(n16973), .A3(n16972), .A4(n16971), .ZN(
        n16975) );
  AOI211_X1 U20231 ( .C1(n17181), .C2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n16976), .B(n16975), .ZN(n16977) );
  OAI211_X1 U20232 ( .C1(n10298), .C2(n18230), .A(n16978), .B(n16977), .ZN(
        n17288) );
  AOI22_X1 U20233 ( .A1(n17227), .A2(n17288), .B1(n16979), .B2(n16981), .ZN(
        n16980) );
  OAI21_X1 U20234 ( .B1(n16981), .B2(n16996), .A(n16980), .ZN(P3_U2682) );
  AOI22_X1 U20235 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16992) );
  AOI22_X1 U20236 ( .A1(n17177), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16982) );
  OAI21_X1 U20237 ( .B1(n17170), .B2(n17101), .A(n16982), .ZN(n16990) );
  INV_X1 U20238 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n20874) );
  AOI22_X1 U20239 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20240 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16984) );
  AOI22_X1 U20241 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16983) );
  OAI211_X1 U20242 ( .C1(n17143), .C2(n16985), .A(n16984), .B(n16983), .ZN(
        n16986) );
  AOI21_X1 U20243 ( .B1(n17031), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n16986), .ZN(n16987) );
  OAI211_X1 U20244 ( .C1(n10298), .C2(n20874), .A(n16988), .B(n16987), .ZN(
        n16989) );
  AOI211_X1 U20245 ( .C1(n17181), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n16990), .B(n16989), .ZN(n16991) );
  OAI211_X1 U20246 ( .C1(n9796), .C2(n20909), .A(n16992), .B(n16991), .ZN(
        n17293) );
  NAND2_X1 U20247 ( .A1(n17227), .A2(n17293), .ZN(n16993) );
  OAI221_X1 U20248 ( .B1(n16996), .B2(n16995), .C1(n16996), .C2(n16994), .A(
        n16993), .ZN(P3_U2683) );
  NAND2_X1 U20249 ( .A1(n17222), .A2(n16997), .ZN(n17021) );
  AOI22_X1 U20250 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20251 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17007) );
  OAI22_X1 U20252 ( .A1(n17118), .A2(n18276), .B1(n10298), .B2(n18222), .ZN(
        n17005) );
  AOI22_X1 U20253 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20254 ( .A1(n9733), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20255 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n16998), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16999) );
  OAI211_X1 U20256 ( .C1(n17188), .C2(n17117), .A(n17000), .B(n16999), .ZN(
        n17001) );
  AOI21_X1 U20257 ( .B1(n17183), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n17001), .ZN(n17002) );
  OAI211_X1 U20258 ( .C1(n17143), .C2(n17120), .A(n17003), .B(n17002), .ZN(
        n17004) );
  AOI211_X1 U20259 ( .C1(n17138), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n17005), .B(n17004), .ZN(n17006) );
  NAND3_X1 U20260 ( .A1(n17008), .A2(n17007), .A3(n17006), .ZN(n17298) );
  OAI22_X1 U20261 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17021), .B1(n17298), 
        .B2(n17222), .ZN(n17009) );
  AOI21_X1 U20262 ( .B1(n17010), .B2(n17222), .A(n17009), .ZN(P3_U2684) );
  AOI22_X1 U20263 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17011) );
  OAI21_X1 U20264 ( .B1(n17170), .B2(n17151), .A(n17011), .ZN(n17020) );
  AOI22_X1 U20265 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17018) );
  INV_X1 U20266 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18217) );
  INV_X1 U20267 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17142) );
  OAI22_X1 U20268 ( .A1(n10298), .A2(n18217), .B1(n10221), .B2(n17142), .ZN(
        n17016) );
  AOI22_X1 U20269 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20270 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20271 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17038), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17012) );
  NAND3_X1 U20272 ( .A1(n17014), .A2(n17013), .A3(n17012), .ZN(n17015) );
  AOI211_X1 U20273 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17016), .B(n17015), .ZN(n17017) );
  OAI211_X1 U20274 ( .C1(n17121), .C2(n20961), .A(n17018), .B(n17017), .ZN(
        n17019) );
  AOI211_X1 U20275 ( .C1(n17173), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17020), .B(n17019), .ZN(n17307) );
  NOR2_X1 U20276 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n9829), .ZN(n17022) );
  OAI22_X1 U20277 ( .A1(n17307), .A2(n17222), .B1(n17022), .B2(n17021), .ZN(
        P3_U2685) );
  INV_X1 U20278 ( .A(n17049), .ZN(n17023) );
  OAI21_X1 U20279 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n17023), .A(n17222), .ZN(
        n17036) );
  AOI22_X1 U20280 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17104), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17024) );
  OAI21_X1 U20281 ( .B1(n9796), .B2(n17025), .A(n17024), .ZN(n17035) );
  AOI22_X1 U20282 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n9733), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20283 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17185), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17183), .ZN(n17026) );
  OAI21_X1 U20284 ( .B1(n20831), .B2(n10298), .A(n17026), .ZN(n17030) );
  AOI22_X1 U20285 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17156), .ZN(n17028) );
  AOI22_X1 U20286 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17177), .ZN(n17027) );
  OAI211_X1 U20287 ( .C1(n20881), .C2(n17143), .A(n17028), .B(n17027), .ZN(
        n17029) );
  AOI211_X1 U20288 ( .C1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .C2(n17031), .A(
        n17030), .B(n17029), .ZN(n17032) );
  OAI211_X1 U20289 ( .C1(n20876), .C2(n10234), .A(n17033), .B(n17032), .ZN(
        n17034) );
  AOI211_X1 U20290 ( .C1(n17173), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n17035), .B(n17034), .ZN(n17313) );
  OAI22_X1 U20291 ( .A1(n9829), .A2(n17036), .B1(n17313), .B2(n17222), .ZN(
        P3_U2686) );
  AOI22_X1 U20292 ( .A1(n17139), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17037) );
  OAI21_X1 U20293 ( .B1(n10234), .B2(n18450), .A(n17037), .ZN(n17048) );
  AOI22_X1 U20294 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17046) );
  AOI22_X1 U20295 ( .A1(n17038), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17039) );
  OAI21_X1 U20296 ( .B1(n10275), .B2(n20856), .A(n17039), .ZN(n17044) );
  AOI22_X1 U20297 ( .A1(n9733), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20298 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17040) );
  OAI211_X1 U20299 ( .C1(n17143), .C2(n17042), .A(n17041), .B(n17040), .ZN(
        n17043) );
  AOI211_X1 U20300 ( .C1(n9795), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17044), .B(n17043), .ZN(n17045) );
  OAI211_X1 U20301 ( .C1(n17118), .C2(n18268), .A(n17046), .B(n17045), .ZN(
        n17047) );
  AOI211_X1 U20302 ( .C1(n17173), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n17048), .B(n17047), .ZN(n17320) );
  OAI21_X1 U20303 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17066), .A(n17049), .ZN(
        n17050) );
  AOI22_X1 U20304 ( .A1(n17227), .A2(n17320), .B1(n17050), .B2(n17222), .ZN(
        P3_U2687) );
  INV_X1 U20305 ( .A(n17051), .ZN(n17052) );
  OAI21_X1 U20306 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17052), .A(n17222), .ZN(
        n17065) );
  AOI22_X1 U20307 ( .A1(n17104), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17053) );
  OAI21_X1 U20308 ( .B1(n17170), .B2(n20968), .A(n17053), .ZN(n17064) );
  AOI22_X1 U20309 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17061) );
  INV_X1 U20310 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20311 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17054) );
  OAI21_X1 U20312 ( .B1(n10268), .B2(n17055), .A(n17054), .ZN(n17059) );
  AOI22_X1 U20313 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20314 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17056) );
  OAI211_X1 U20315 ( .C1(n17188), .C2(n21001), .A(n17057), .B(n17056), .ZN(
        n17058) );
  AOI211_X1 U20316 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n17059), .B(n17058), .ZN(n17060) );
  OAI211_X1 U20317 ( .C1(n17121), .C2(n17062), .A(n17061), .B(n17060), .ZN(
        n17063) );
  AOI211_X1 U20318 ( .C1(n17185), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n17064), .B(n17063), .ZN(n17324) );
  OAI22_X1 U20319 ( .A1(n17066), .A2(n17065), .B1(n17324), .B2(n17222), .ZN(
        P3_U2688) );
  AOI22_X1 U20320 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17067) );
  OAI21_X1 U20321 ( .B1(n17118), .B2(n17068), .A(n17067), .ZN(n17079) );
  INV_X1 U20322 ( .A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17077) );
  AOI22_X1 U20323 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17076) );
  AOI22_X1 U20324 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17069) );
  OAI21_X1 U20325 ( .B1(n10298), .B2(n17070), .A(n17069), .ZN(n17074) );
  AOI22_X1 U20326 ( .A1(n9733), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20327 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17071) );
  OAI211_X1 U20328 ( .C1(n17188), .C2(n18236), .A(n17072), .B(n17071), .ZN(
        n17073) );
  AOI211_X1 U20329 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17074), .B(n17073), .ZN(n17075) );
  OAI211_X1 U20330 ( .C1(n9796), .C2(n17077), .A(n17076), .B(n17075), .ZN(
        n17078) );
  AOI211_X1 U20331 ( .C1(n9722), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n17079), .B(n17078), .ZN(n17328) );
  NOR2_X1 U20332 ( .A1(n17227), .A2(n17080), .ZN(n17097) );
  NOR2_X1 U20333 ( .A1(n17218), .A2(n17204), .ZN(n17202) );
  INV_X1 U20334 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17082) );
  NOR4_X1 U20335 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17083), .A3(n17082), .A4(
        n17081), .ZN(n17084) );
  AOI22_X1 U20336 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17097), .B1(n17202), 
        .B2(n17084), .ZN(n17085) );
  OAI21_X1 U20337 ( .B1(n17328), .B2(n17222), .A(n17085), .ZN(P3_U2689) );
  AOI22_X1 U20338 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20339 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17086) );
  OAI21_X1 U20340 ( .B1(n9794), .B2(n21035), .A(n17086), .ZN(n17094) );
  OAI22_X1 U20341 ( .A1(n17188), .A2(n18230), .B1(n10267), .B2(n17087), .ZN(
        n17088) );
  AOI21_X1 U20342 ( .B1(n17182), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n17088), .ZN(n17092) );
  AOI22_X1 U20343 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17091) );
  AOI22_X1 U20344 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17090) );
  AOI22_X1 U20345 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17089) );
  NAND4_X1 U20346 ( .A1(n17092), .A2(n17091), .A3(n17090), .A4(n17089), .ZN(
        n17093) );
  AOI211_X1 U20347 ( .C1(n17155), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n17094), .B(n17093), .ZN(n17095) );
  OAI211_X1 U20348 ( .C1(n17170), .C2(n20858), .A(n17096), .B(n17095), .ZN(
        n17332) );
  INV_X1 U20349 ( .A(n17332), .ZN(n17100) );
  INV_X1 U20350 ( .A(n17114), .ZN(n17098) );
  OAI21_X1 U20351 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17098), .A(n17097), .ZN(
        n17099) );
  OAI21_X1 U20352 ( .B1(n17100), .B2(n17222), .A(n17099), .ZN(P3_U2690) );
  OAI22_X1 U20353 ( .A1(n9800), .A2(n20841), .B1(n10298), .B2(n17101), .ZN(
        n17113) );
  AOI22_X1 U20354 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20355 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20356 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9727), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17102) );
  OAI21_X1 U20357 ( .B1(n17143), .B2(n17103), .A(n17102), .ZN(n17108) );
  AOI22_X1 U20358 ( .A1(n17104), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17106) );
  AOI22_X1 U20359 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9733), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17105) );
  OAI211_X1 U20360 ( .C1(n17188), .C2(n20874), .A(n17106), .B(n17105), .ZN(
        n17107) );
  AOI211_X1 U20361 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n17108), .B(n17107), .ZN(n17109) );
  NAND3_X1 U20362 ( .A1(n17111), .A2(n17110), .A3(n17109), .ZN(n17112) );
  AOI211_X1 U20363 ( .C1(n10309), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n17113), .B(n17112), .ZN(n17336) );
  OAI21_X1 U20364 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17135), .A(n17114), .ZN(
        n17115) );
  AOI22_X1 U20365 ( .A1(n17227), .A2(n17336), .B1(n17115), .B2(n17222), .ZN(
        P3_U2691) );
  NOR3_X1 U20366 ( .A1(n20850), .A2(n17197), .A3(n17204), .ZN(n17174) );
  AND2_X1 U20367 ( .A1(n17116), .A2(n17174), .ZN(n17153) );
  OAI21_X1 U20368 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17153), .A(n17222), .ZN(
        n17134) );
  OAI22_X1 U20369 ( .A1(n17118), .A2(n17117), .B1(n17170), .B2(n20882), .ZN(
        n17133) );
  OAI22_X1 U20370 ( .A1(n17121), .A2(n17120), .B1(n10267), .B2(n17119), .ZN(
        n17132) );
  INV_X1 U20371 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20372 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17129) );
  INV_X1 U20373 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17123) );
  AOI22_X1 U20374 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17122) );
  OAI21_X1 U20375 ( .B1(n17143), .B2(n17123), .A(n17122), .ZN(n17127) );
  AOI22_X1 U20376 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17125) );
  AOI22_X1 U20377 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17124) );
  OAI211_X1 U20378 ( .C1(n17188), .C2(n18222), .A(n17125), .B(n17124), .ZN(
        n17126) );
  AOI211_X1 U20379 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17127), .B(n17126), .ZN(n17128) );
  OAI211_X1 U20380 ( .C1(n10275), .C2(n17130), .A(n17129), .B(n17128), .ZN(
        n17131) );
  NOR3_X1 U20381 ( .A1(n17133), .A2(n17132), .A3(n17131), .ZN(n17340) );
  OAI22_X1 U20382 ( .A1(n17135), .A2(n17134), .B1(n17340), .B2(n17222), .ZN(
        P3_U2692) );
  AOI22_X1 U20383 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20384 ( .A1(n9733), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17136) );
  OAI21_X1 U20385 ( .B1(n10234), .B2(n17137), .A(n17136), .ZN(n17148) );
  AOI22_X1 U20386 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U20387 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20388 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17140) );
  OAI211_X1 U20389 ( .C1(n17143), .C2(n17142), .A(n17141), .B(n17140), .ZN(
        n17144) );
  AOI21_X1 U20390 ( .B1(n17183), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n17144), .ZN(n17145) );
  OAI211_X1 U20391 ( .C1(n17188), .C2(n18217), .A(n17146), .B(n17145), .ZN(
        n17147) );
  AOI211_X1 U20392 ( .C1(n17173), .C2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n17148), .B(n17147), .ZN(n17149) );
  OAI211_X1 U20393 ( .C1(n10298), .C2(n17151), .A(n17150), .B(n17149), .ZN(
        n17343) );
  INV_X1 U20394 ( .A(n17343), .ZN(n17154) );
  AND2_X1 U20395 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17174), .ZN(n17176) );
  OAI21_X1 U20396 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17176), .A(n17222), .ZN(
        n17152) );
  OAI22_X1 U20397 ( .A1(n17154), .A2(n17222), .B1(n17153), .B2(n17152), .ZN(
        P3_U2693) );
  AOI22_X1 U20398 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17156), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17157) );
  OAI21_X1 U20399 ( .B1(n9800), .B2(n17158), .A(n17157), .ZN(n17172) );
  AOI22_X1 U20400 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17182), .ZN(n17168) );
  AOI22_X1 U20401 ( .A1(n9727), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17191), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17160) );
  OAI21_X1 U20402 ( .B1(n17161), .B2(n10267), .A(n17160), .ZN(n17166) );
  AOI22_X1 U20403 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17139), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20404 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17163) );
  OAI211_X1 U20405 ( .C1(n20831), .C2(n17188), .A(n17164), .B(n17163), .ZN(
        n17165) );
  AOI211_X1 U20406 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n17166), .B(n17165), .ZN(n17167) );
  OAI211_X1 U20407 ( .C1(n17170), .C2(n17169), .A(n17168), .B(n17167), .ZN(
        n17171) );
  AOI211_X1 U20408 ( .C1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(n17173), .A(
        n17172), .B(n17171), .ZN(n17349) );
  OAI21_X1 U20409 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17174), .A(n17222), .ZN(
        n17175) );
  OAI22_X1 U20410 ( .A1(n17349), .A2(n17222), .B1(n17176), .B2(n17175), .ZN(
        P3_U2694) );
  AOI22_X1 U20411 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17177), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17178) );
  OAI21_X1 U20412 ( .B1(n10234), .B2(n17179), .A(n17178), .ZN(n17196) );
  AOI22_X1 U20413 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17193) );
  AOI22_X1 U20414 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17182), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17184) );
  OAI21_X1 U20415 ( .B1(n10221), .B2(n18450), .A(n17184), .ZN(n17190) );
  AOI22_X1 U20416 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9733), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17187) );
  AOI22_X1 U20417 ( .A1(n17185), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17139), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17186) );
  OAI211_X1 U20418 ( .C1(n17188), .C2(n18208), .A(n17187), .B(n17186), .ZN(
        n17189) );
  AOI211_X1 U20419 ( .C1(n17191), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17190), .B(n17189), .ZN(n17192) );
  OAI211_X1 U20420 ( .C1(n10275), .C2(n17194), .A(n17193), .B(n17192), .ZN(
        n17195) );
  AOI211_X1 U20421 ( .C1(n17159), .C2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A(
        n17196), .B(n17195), .ZN(n17357) );
  NOR2_X1 U20422 ( .A1(n17197), .A2(n17204), .ZN(n17200) );
  NAND2_X1 U20423 ( .A1(n17200), .A2(P3_EBX_REG_8__SCAN_IN), .ZN(n17198) );
  OAI211_X1 U20424 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17200), .A(n17222), .B(
        n17198), .ZN(n17199) );
  OAI21_X1 U20425 ( .B1(n17357), .B2(n17222), .A(n17199), .ZN(P3_U2695) );
  INV_X1 U20426 ( .A(n17200), .ZN(n17201) );
  OAI211_X1 U20427 ( .C1(P3_EBX_REG_7__SCAN_IN), .C2(n17202), .A(n17201), .B(
        n17222), .ZN(n17203) );
  OAI21_X1 U20428 ( .B1(n17222), .B2(n21001), .A(n17203), .ZN(P3_U2696) );
  INV_X1 U20429 ( .A(n17204), .ZN(n17207) );
  INV_X1 U20430 ( .A(n17224), .ZN(n17226) );
  NAND2_X1 U20431 ( .A1(n17205), .A2(n17226), .ZN(n17212) );
  NOR2_X1 U20432 ( .A1(n20813), .A2(n17212), .ZN(n17214) );
  AOI22_X1 U20433 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17222), .B1(
        P3_EBX_REG_5__SCAN_IN), .B2(n17214), .ZN(n17206) );
  OAI22_X1 U20434 ( .A1(n17207), .A2(n17206), .B1(n18236), .B2(n17222), .ZN(
        P3_U2697) );
  INV_X1 U20435 ( .A(n17208), .ZN(n17209) );
  OAI21_X1 U20436 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17209), .A(n17222), .ZN(
        n17210) );
  OAI22_X1 U20437 ( .A1(n17211), .A2(n17210), .B1(n18230), .B2(n17222), .ZN(
        P3_U2698) );
  INV_X1 U20438 ( .A(n17212), .ZN(n17217) );
  AOI21_X1 U20439 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17222), .A(n17217), .ZN(
        n17213) );
  OAI22_X1 U20440 ( .A1(n17214), .A2(n17213), .B1(n20874), .B2(n17222), .ZN(
        P3_U2699) );
  NOR2_X1 U20441 ( .A1(n17215), .A2(n17224), .ZN(n17220) );
  AOI21_X1 U20442 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17222), .A(n17220), .ZN(
        n17216) );
  OAI22_X1 U20443 ( .A1(n17217), .A2(n17216), .B1(n18222), .B2(n17222), .ZN(
        P3_U2700) );
  AOI221_X1 U20444 ( .B1(n17219), .B2(n17230), .C1(n17218), .C2(n17230), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17221) );
  AOI211_X1 U20445 ( .C1(n17227), .C2(n18217), .A(n17221), .B(n17220), .ZN(
        P3_U2701) );
  OAI222_X1 U20446 ( .A1(n17225), .A2(n17224), .B1(n17223), .B2(n17230), .C1(
        n20831), .C2(n17222), .ZN(P3_U2702) );
  AOI22_X1 U20447 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17227), .B1(
        n17226), .B2(n17229), .ZN(n17228) );
  OAI21_X1 U20448 ( .B1(n17230), .B2(n17229), .A(n17228), .ZN(P3_U2703) );
  NAND2_X1 U20449 ( .A1(n17353), .A2(n17231), .ZN(n17283) );
  INV_X1 U20450 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17397) );
  INV_X1 U20451 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17400) );
  INV_X1 U20452 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17404) );
  INV_X1 U20453 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17406) );
  INV_X1 U20454 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17420) );
  INV_X1 U20455 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17423) );
  NAND2_X1 U20456 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17385) );
  INV_X1 U20457 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17439) );
  INV_X1 U20458 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17441) );
  NAND4_X1 U20459 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17232) );
  NOR4_X1 U20460 ( .A1(n17385), .A2(n17439), .A3(n17441), .A4(n17232), .ZN(
        n17325) );
  INV_X1 U20461 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17429) );
  INV_X1 U20462 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17431) );
  INV_X1 U20463 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17433) );
  NOR3_X1 U20464 ( .A1(n17429), .A2(n17431), .A3(n17433), .ZN(n17331) );
  NAND4_X1 U20465 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .A4(n17331), .ZN(n17326) );
  INV_X1 U20466 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17408) );
  INV_X1 U20467 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17410) );
  INV_X1 U20468 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17412) );
  INV_X1 U20469 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17417) );
  NOR4_X1 U20470 ( .A1(n17408), .A2(n17410), .A3(n17412), .A4(n17417), .ZN(
        n17234) );
  NAND4_X1 U20471 ( .A1(n17316), .A2(P3_EAX_REG_19__SCAN_IN), .A3(
        P3_EAX_REG_18__SCAN_IN), .A4(n17234), .ZN(n17278) );
  NAND2_X1 U20472 ( .A1(n18240), .A2(n17277), .ZN(n17270) );
  NAND2_X1 U20473 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17250), .ZN(n17245) );
  NOR2_X1 U20474 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17245), .ZN(n17236) );
  NAND2_X1 U20475 ( .A1(n17378), .A2(n17245), .ZN(n17243) );
  OAI21_X1 U20476 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17376), .A(n17243), .ZN(
        n17235) );
  AOI22_X1 U20477 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17236), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17235), .ZN(n17237) );
  OAI21_X1 U20478 ( .B1(n19237), .B2(n17283), .A(n17237), .ZN(P3_U2704) );
  INV_X1 U20479 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17394) );
  NOR2_X2 U20480 ( .A1(n17238), .A2(n17378), .ZN(n17315) );
  OAI22_X1 U20481 ( .A1(n17240), .A2(n17389), .B1(n17239), .B2(n17283), .ZN(
        n17241) );
  AOI21_X1 U20482 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17315), .A(n17241), .ZN(
        n17242) );
  OAI221_X1 U20483 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17245), .C1(n17394), 
        .C2(n17243), .A(n17242), .ZN(P3_U2705) );
  AOI22_X1 U20484 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17315), .B1(n17244), .B2(
        n17344), .ZN(n17247) );
  OAI211_X1 U20485 ( .C1(n17250), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17378), .B(
        n17245), .ZN(n17246) );
  OAI211_X1 U20486 ( .C1(n17283), .C2(n17248), .A(n17247), .B(n17246), .ZN(
        P3_U2706) );
  AOI22_X1 U20487 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17315), .B1(n17249), .B2(
        n17344), .ZN(n17253) );
  AOI211_X1 U20488 ( .C1(n17397), .C2(n17257), .A(n17250), .B(n17353), .ZN(
        n17251) );
  INV_X1 U20489 ( .A(n17251), .ZN(n17252) );
  OAI211_X1 U20490 ( .C1(n17283), .C2(n19222), .A(n17253), .B(n17252), .ZN(
        P3_U2707) );
  OAI21_X1 U20491 ( .B1(n17256), .B2(n17255), .A(n17254), .ZN(n17260) );
  AOI22_X1 U20492 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17315), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17314), .ZN(n17259) );
  OAI211_X1 U20493 ( .C1(n17261), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17378), .B(
        n17257), .ZN(n17258) );
  OAI211_X1 U20494 ( .C1(n17389), .C2(n17260), .A(n17259), .B(n17258), .ZN(
        P3_U2708) );
  AOI22_X1 U20495 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17315), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17314), .ZN(n17264) );
  AOI211_X1 U20496 ( .C1(n17400), .C2(n17266), .A(n17261), .B(n17353), .ZN(
        n17262) );
  INV_X1 U20497 ( .A(n17262), .ZN(n17263) );
  OAI211_X1 U20498 ( .C1(n17389), .C2(n17265), .A(n17264), .B(n17263), .ZN(
        P3_U2709) );
  AOI22_X1 U20499 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17315), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17314), .ZN(n17268) );
  OAI211_X1 U20500 ( .C1(n17271), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17378), .B(
        n17266), .ZN(n17267) );
  OAI211_X1 U20501 ( .C1(n17389), .C2(n17269), .A(n17268), .B(n17267), .ZN(
        P3_U2710) );
  AOI22_X1 U20502 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17315), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17314), .ZN(n17275) );
  OAI21_X1 U20503 ( .B1(n17404), .B2(n17353), .A(n17270), .ZN(n17273) );
  INV_X1 U20504 ( .A(n17271), .ZN(n17272) );
  NAND2_X1 U20505 ( .A1(n17273), .A2(n17272), .ZN(n17274) );
  OAI211_X1 U20506 ( .C1(n17276), .C2(n17389), .A(n17275), .B(n17274), .ZN(
        P3_U2711) );
  AOI211_X1 U20507 ( .C1(n17406), .C2(n17278), .A(n17353), .B(n17277), .ZN(
        n17281) );
  INV_X1 U20508 ( .A(n17315), .ZN(n17297) );
  OAI22_X1 U20509 ( .A1(n18237), .A2(n17297), .B1(n17389), .B2(n17279), .ZN(
        n17280) );
  AOI211_X1 U20510 ( .C1(n17314), .C2(BUF2_REG_23__SCAN_IN), .A(n17281), .B(
        n17280), .ZN(n17282) );
  INV_X1 U20511 ( .A(n17282), .ZN(P3_U2712) );
  INV_X1 U20512 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17414) );
  INV_X1 U20513 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17416) );
  NAND2_X1 U20514 ( .A1(n18240), .A2(n17316), .ZN(n17308) );
  NAND2_X1 U20515 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17302), .ZN(n17294) );
  NAND2_X1 U20516 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17290), .ZN(n17289) );
  NAND2_X1 U20517 ( .A1(n17289), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17287) );
  OAI22_X1 U20518 ( .A1(n17284), .A2(n17389), .B1(n18233), .B2(n17283), .ZN(
        n17285) );
  AOI21_X1 U20519 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17315), .A(n17285), .ZN(
        n17286) );
  OAI221_X1 U20520 ( .B1(n17289), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17287), 
        .C2(n17353), .A(n17286), .ZN(P3_U2713) );
  AOI22_X1 U20521 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n17314), .B1(n17344), .B2(
        n17288), .ZN(n17292) );
  OAI211_X1 U20522 ( .C1(n17290), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17378), .B(
        n17289), .ZN(n17291) );
  OAI211_X1 U20523 ( .C1(n17297), .C2(n20847), .A(n17292), .B(n17291), .ZN(
        P3_U2714) );
  AOI22_X1 U20524 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17314), .B1(n17344), .B2(
        n17293), .ZN(n17296) );
  OAI211_X1 U20525 ( .C1(n17302), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17378), .B(
        n17294), .ZN(n17295) );
  OAI211_X1 U20526 ( .C1(n17297), .C2(n18223), .A(n17296), .B(n17295), .ZN(
        P3_U2715) );
  AOI22_X1 U20527 ( .A1(n17304), .A2(P3_EAX_REG_18__SCAN_IN), .B1(
        P3_EAX_REG_19__SCAN_IN), .B2(n17378), .ZN(n17301) );
  AOI22_X1 U20528 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n17314), .B1(n17344), .B2(
        n17298), .ZN(n17300) );
  NAND2_X1 U20529 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17315), .ZN(n17299) );
  OAI211_X1 U20530 ( .C1(n17302), .C2(n17301), .A(n17300), .B(n17299), .ZN(
        P3_U2716) );
  AOI22_X1 U20531 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17315), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17314), .ZN(n17306) );
  NAND2_X1 U20532 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17304), .ZN(n17303) );
  OAI211_X1 U20533 ( .C1(n17304), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17378), .B(
        n17303), .ZN(n17305) );
  OAI211_X1 U20534 ( .C1(n17307), .C2(n17389), .A(n17306), .B(n17305), .ZN(
        P3_U2717) );
  AOI22_X1 U20535 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17315), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17314), .ZN(n17312) );
  OAI21_X1 U20536 ( .B1(n17417), .B2(n17353), .A(n17308), .ZN(n17310) );
  NAND2_X1 U20537 ( .A1(n17310), .A2(n17309), .ZN(n17311) );
  OAI211_X1 U20538 ( .C1(n17313), .C2(n17389), .A(n17312), .B(n17311), .ZN(
        P3_U2718) );
  AOI22_X1 U20539 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17315), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17314), .ZN(n17319) );
  AOI211_X1 U20540 ( .C1(n17420), .C2(n17321), .A(n17353), .B(n17316), .ZN(
        n17317) );
  INV_X1 U20541 ( .A(n17317), .ZN(n17318) );
  OAI211_X1 U20542 ( .C1(n17320), .C2(n17389), .A(n17319), .B(n17318), .ZN(
        P3_U2719) );
  OAI211_X1 U20543 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17330), .A(n17378), .B(
        n17321), .ZN(n17323) );
  NAND2_X1 U20544 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17384), .ZN(n17322) );
  OAI211_X1 U20545 ( .C1(n17324), .C2(n17389), .A(n17323), .B(n17322), .ZN(
        P3_U2720) );
  INV_X1 U20546 ( .A(n17376), .ZN(n17386) );
  INV_X1 U20547 ( .A(n17326), .ZN(n17327) );
  AOI22_X1 U20548 ( .A1(n17360), .A2(n17327), .B1(P3_EAX_REG_14__SCAN_IN), 
        .B2(n17378), .ZN(n17329) );
  OAI222_X1 U20549 ( .A1(n17382), .A2(n17496), .B1(n17330), .B2(n17329), .C1(
        n17389), .C2(n17328), .ZN(P3_U2721) );
  NAND2_X1 U20550 ( .A1(n17331), .A2(n17360), .ZN(n17345) );
  INV_X1 U20551 ( .A(n17345), .ZN(n17339) );
  NAND2_X1 U20552 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17342), .ZN(n17335) );
  NAND2_X1 U20553 ( .A1(n17335), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U20554 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17384), .B1(n17344), .B2(
        n17332), .ZN(n17333) );
  OAI221_X1 U20555 ( .B1(n17335), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17334), 
        .C2(n17353), .A(n17333), .ZN(P3_U2722) );
  INV_X1 U20556 ( .A(n17335), .ZN(n17338) );
  AOI21_X1 U20557 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17378), .A(n17342), .ZN(
        n17337) );
  OAI222_X1 U20558 ( .A1(n17382), .A2(n17491), .B1(n17338), .B2(n17337), .C1(
        n17389), .C2(n17336), .ZN(P3_U2723) );
  AOI21_X1 U20559 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17378), .A(n17339), .ZN(
        n17341) );
  OAI222_X1 U20560 ( .A1(n17382), .A2(n17488), .B1(n17342), .B2(n17341), .C1(
        n17389), .C2(n17340), .ZN(P3_U2724) );
  AOI22_X1 U20561 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17384), .B1(n17344), .B2(
        n17343), .ZN(n17347) );
  NAND2_X1 U20562 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17360), .ZN(n17348) );
  NOR2_X1 U20563 ( .A1(n17431), .A2(n17348), .ZN(n17351) );
  OAI211_X1 U20564 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17351), .A(n17378), .B(
        n17345), .ZN(n17346) );
  NAND2_X1 U20565 ( .A1(n17347), .A2(n17346), .ZN(P3_U2725) );
  INV_X1 U20566 ( .A(n17348), .ZN(n17352) );
  AOI21_X1 U20567 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17378), .A(n17352), .ZN(
        n17350) );
  OAI222_X1 U20568 ( .A1(n17382), .A2(n17484), .B1(n17351), .B2(n17350), .C1(
        n17389), .C2(n17349), .ZN(P3_U2726) );
  AOI211_X1 U20569 ( .C1(n17354), .C2(n17433), .A(n17353), .B(n17352), .ZN(
        n17355) );
  AOI21_X1 U20570 ( .B1(n17384), .B2(BUF2_REG_8__SCAN_IN), .A(n17355), .ZN(
        n17356) );
  OAI21_X1 U20571 ( .B1(n17357), .B2(n17389), .A(n17356), .ZN(P3_U2727) );
  INV_X1 U20572 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17437) );
  INV_X1 U20573 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17446) );
  NOR3_X1 U20574 ( .A1(n17385), .A2(n17446), .A3(n17376), .ZN(n17381) );
  NAND2_X1 U20575 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17381), .ZN(n17369) );
  NOR2_X1 U20576 ( .A1(n17441), .A2(n17369), .ZN(n17372) );
  NAND2_X1 U20577 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17372), .ZN(n17361) );
  NOR2_X1 U20578 ( .A1(n17437), .A2(n17361), .ZN(n17365) );
  AOI21_X1 U20579 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17378), .A(n17365), .ZN(
        n17359) );
  OAI222_X1 U20580 ( .A1(n18237), .A2(n17382), .B1(n17360), .B2(n17359), .C1(
        n17389), .C2(n17358), .ZN(P3_U2728) );
  INV_X1 U20581 ( .A(n17361), .ZN(n17368) );
  AOI21_X1 U20582 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17378), .A(n17368), .ZN(
        n17364) );
  INV_X1 U20583 ( .A(n17362), .ZN(n17363) );
  OAI222_X1 U20584 ( .A1(n18231), .A2(n17382), .B1(n17365), .B2(n17364), .C1(
        n17389), .C2(n17363), .ZN(P3_U2729) );
  AOI21_X1 U20585 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17378), .A(n17372), .ZN(
        n17367) );
  OAI222_X1 U20586 ( .A1(n20847), .A2(n17382), .B1(n17368), .B2(n17367), .C1(
        n17389), .C2(n17366), .ZN(P3_U2730) );
  INV_X1 U20587 ( .A(n17369), .ZN(n17375) );
  AOI21_X1 U20588 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17378), .A(n17375), .ZN(
        n17371) );
  OAI222_X1 U20589 ( .A1(n18223), .A2(n17382), .B1(n17372), .B2(n17371), .C1(
        n17389), .C2(n17370), .ZN(P3_U2731) );
  AOI21_X1 U20590 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17378), .A(n17381), .ZN(
        n17374) );
  OAI222_X1 U20591 ( .A1(n18218), .A2(n17382), .B1(n17375), .B2(n17374), .C1(
        n17389), .C2(n17373), .ZN(P3_U2732) );
  NOR2_X1 U20592 ( .A1(n17385), .A2(n17376), .ZN(n17377) );
  AOI21_X1 U20593 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17378), .A(n17377), .ZN(
        n17380) );
  OAI222_X1 U20594 ( .A1(n18213), .A2(n17382), .B1(n17381), .B2(n17380), .C1(
        n17389), .C2(n17379), .ZN(P3_U2733) );
  AOI22_X1 U20595 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17384), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n17383), .ZN(n17388) );
  OAI211_X1 U20596 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17386), .B(n17385), .ZN(n17387) );
  OAI211_X1 U20597 ( .C1(n10350), .C2(n17389), .A(n17388), .B(n17387), .ZN(
        P3_U2734) );
  OR2_X1 U20598 ( .A1(n17857), .A2(n17856), .ZN(n18863) );
  NOR2_X1 U20599 ( .A1(n17426), .A2(n17391), .ZN(P3_U2736) );
  INV_X2 U20600 ( .A(n18863), .ZN(n17450) );
  AOI22_X1 U20601 ( .A1(n17450), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17444), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17393) );
  OAI21_X1 U20602 ( .B1(n17394), .B2(n17419), .A(n17393), .ZN(P3_U2737) );
  INV_X1 U20603 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17470) );
  AOI22_X1 U20604 ( .A1(n17450), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17395) );
  OAI21_X1 U20605 ( .B1(n17470), .B2(n17419), .A(n17395), .ZN(P3_U2738) );
  AOI22_X1 U20606 ( .A1(P3_UWORD_REG_12__SCAN_IN), .A2(n17450), .B1(n17449), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17396) );
  OAI21_X1 U20607 ( .B1(n17397), .B2(n17419), .A(n17396), .ZN(P3_U2739) );
  INV_X1 U20608 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n20947) );
  INV_X1 U20609 ( .A(n17419), .ZN(n17401) );
  AOI22_X1 U20610 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17401), .B1(n17450), 
        .B2(P3_UWORD_REG_11__SCAN_IN), .ZN(n17398) );
  OAI21_X1 U20611 ( .B1(n20947), .B2(n17426), .A(n17398), .ZN(P3_U2740) );
  AOI22_X1 U20612 ( .A1(n17450), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17399) );
  OAI21_X1 U20613 ( .B1(n17400), .B2(n17419), .A(n17399), .ZN(P3_U2741) );
  INV_X1 U20614 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n20938) );
  AOI22_X1 U20615 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17401), .B1(n17450), 
        .B2(P3_UWORD_REG_9__SCAN_IN), .ZN(n17402) );
  OAI21_X1 U20616 ( .B1(n20938), .B2(n17426), .A(n17402), .ZN(P3_U2742) );
  AOI22_X1 U20617 ( .A1(n17450), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17403) );
  OAI21_X1 U20618 ( .B1(n17404), .B2(n17419), .A(n17403), .ZN(P3_U2743) );
  AOI22_X1 U20619 ( .A1(n17450), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17405) );
  OAI21_X1 U20620 ( .B1(n17406), .B2(n17419), .A(n17405), .ZN(P3_U2744) );
  AOI22_X1 U20621 ( .A1(n17450), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17407) );
  OAI21_X1 U20622 ( .B1(n17408), .B2(n17419), .A(n17407), .ZN(P3_U2745) );
  AOI22_X1 U20623 ( .A1(n17450), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20624 ( .B1(n17410), .B2(n17419), .A(n17409), .ZN(P3_U2746) );
  AOI22_X1 U20625 ( .A1(P3_DATAO_REG_20__SCAN_IN), .A2(n17449), .B1(n17450), 
        .B2(P3_UWORD_REG_4__SCAN_IN), .ZN(n17411) );
  OAI21_X1 U20626 ( .B1(n17412), .B2(n17419), .A(n17411), .ZN(P3_U2747) );
  AOI22_X1 U20627 ( .A1(n17450), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17413) );
  OAI21_X1 U20628 ( .B1(n17414), .B2(n17419), .A(n17413), .ZN(P3_U2748) );
  AOI22_X1 U20629 ( .A1(n17450), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17415) );
  OAI21_X1 U20630 ( .B1(n17416), .B2(n17419), .A(n17415), .ZN(P3_U2749) );
  INV_X1 U20631 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n21040) );
  INV_X1 U20632 ( .A(P3_UWORD_REG_1__SCAN_IN), .ZN(n21004) );
  OAI222_X1 U20633 ( .A1(n17419), .A2(n17417), .B1(n17426), .B2(n21040), .C1(
        n18863), .C2(n21004), .ZN(P3_U2750) );
  AOI22_X1 U20634 ( .A1(n17450), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17418) );
  OAI21_X1 U20635 ( .B1(n17420), .B2(n17419), .A(n17418), .ZN(P3_U2751) );
  INV_X1 U20636 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17501) );
  AOI22_X1 U20637 ( .A1(n17450), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17421) );
  OAI21_X1 U20638 ( .B1(n17501), .B2(n17452), .A(n17421), .ZN(P3_U2752) );
  AOI22_X1 U20639 ( .A1(n17450), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17422) );
  OAI21_X1 U20640 ( .B1(n17423), .B2(n17452), .A(n17422), .ZN(P3_U2753) );
  INV_X1 U20641 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17493) );
  AOI22_X1 U20642 ( .A1(n17450), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17424) );
  OAI21_X1 U20643 ( .B1(n17493), .B2(n17452), .A(n17424), .ZN(P3_U2754) );
  INV_X1 U20644 ( .A(P3_DATAO_REG_12__SCAN_IN), .ZN(n20892) );
  AOI22_X1 U20645 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17447), .B1(n17450), 
        .B2(P3_LWORD_REG_12__SCAN_IN), .ZN(n17425) );
  OAI21_X1 U20646 ( .B1(n20892), .B2(n17426), .A(n17425), .ZN(P3_U2755) );
  AOI222_X1 U20647 ( .A1(P3_LWORD_REG_11__SCAN_IN), .A2(n17450), .B1(n17449), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .C1(P3_EAX_REG_11__SCAN_IN), .C2(n17447), .ZN(n17427) );
  INV_X1 U20648 ( .A(n17427), .ZN(P3_U2756) );
  AOI22_X1 U20649 ( .A1(n17450), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17428) );
  OAI21_X1 U20650 ( .B1(n17429), .B2(n17452), .A(n17428), .ZN(P3_U2757) );
  AOI22_X1 U20651 ( .A1(n17450), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17430) );
  OAI21_X1 U20652 ( .B1(n17431), .B2(n17452), .A(n17430), .ZN(P3_U2758) );
  AOI22_X1 U20653 ( .A1(n17450), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17444), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17432) );
  OAI21_X1 U20654 ( .B1(n17433), .B2(n17452), .A(n17432), .ZN(P3_U2759) );
  INV_X1 U20655 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17435) );
  AOI22_X1 U20656 ( .A1(n17450), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17444), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17434) );
  OAI21_X1 U20657 ( .B1(n17435), .B2(n17452), .A(n17434), .ZN(P3_U2760) );
  AOI22_X1 U20658 ( .A1(n17450), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17444), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17436) );
  OAI21_X1 U20659 ( .B1(n17437), .B2(n17452), .A(n17436), .ZN(P3_U2761) );
  AOI22_X1 U20660 ( .A1(n17450), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17444), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17438) );
  OAI21_X1 U20661 ( .B1(n17439), .B2(n17452), .A(n17438), .ZN(P3_U2762) );
  AOI22_X1 U20662 ( .A1(n17450), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17444), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17440) );
  OAI21_X1 U20663 ( .B1(n17441), .B2(n17452), .A(n17440), .ZN(P3_U2763) );
  INV_X1 U20664 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U20665 ( .A1(n17450), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17444), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17442) );
  OAI21_X1 U20666 ( .B1(n17443), .B2(n17452), .A(n17442), .ZN(P3_U2764) );
  AOI22_X1 U20667 ( .A1(n17450), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17444), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17445) );
  OAI21_X1 U20668 ( .B1(n17446), .B2(n17452), .A(n17445), .ZN(P3_U2765) );
  INV_X1 U20669 ( .A(P3_LWORD_REG_1__SCAN_IN), .ZN(n20988) );
  AOI22_X1 U20670 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17447), .B1(n17449), .B2(
        P3_DATAO_REG_1__SCAN_IN), .ZN(n17448) );
  OAI21_X1 U20671 ( .B1(n20988), .B2(n18863), .A(n17448), .ZN(P3_U2766) );
  AOI22_X1 U20672 ( .A1(n17450), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17449), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17451) );
  OAI21_X1 U20673 ( .B1(n17453), .B2(n17452), .A(n17451), .ZN(P3_U2767) );
  INV_X1 U20674 ( .A(n18707), .ZN(n18864) );
  OR2_X1 U20675 ( .A1(n18855), .A2(n17454), .ZN(n18705) );
  INV_X2 U20676 ( .A(n17474), .ZN(n17497) );
  AOI22_X1 U20677 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17497), .ZN(n17456) );
  OAI21_X1 U20678 ( .B1(n18200), .B2(n17495), .A(n17456), .ZN(P3_U2768) );
  AOI22_X1 U20679 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17498), .B1(
        P3_EAX_REG_17__SCAN_IN), .B2(n9729), .ZN(n17457) );
  OAI21_X1 U20680 ( .B1(n17474), .B2(n21004), .A(n17457), .ZN(P3_U2769) );
  AOI22_X1 U20681 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17497), .ZN(n17458) );
  OAI21_X1 U20682 ( .B1(n18213), .B2(n17495), .A(n17458), .ZN(P3_U2770) );
  AOI22_X1 U20683 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17497), .ZN(n17459) );
  OAI21_X1 U20684 ( .B1(n18218), .B2(n17495), .A(n17459), .ZN(P3_U2771) );
  AOI22_X1 U20685 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17497), .ZN(n17460) );
  OAI21_X1 U20686 ( .B1(n18223), .B2(n17495), .A(n17460), .ZN(P3_U2772) );
  AOI22_X1 U20687 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17497), .ZN(n17461) );
  OAI21_X1 U20688 ( .B1(n20847), .B2(n17495), .A(n17461), .ZN(P3_U2773) );
  AOI22_X1 U20689 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17497), .ZN(n17462) );
  OAI21_X1 U20690 ( .B1(n18231), .B2(n17495), .A(n17462), .ZN(P3_U2774) );
  AOI22_X1 U20691 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17497), .ZN(n17463) );
  OAI21_X1 U20692 ( .B1(n18237), .B2(n17495), .A(n17463), .ZN(P3_U2775) );
  AOI22_X1 U20693 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17497), .ZN(n17464) );
  OAI21_X1 U20694 ( .B1(n17482), .B2(n17495), .A(n17464), .ZN(P3_U2776) );
  AOI22_X1 U20695 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17497), .ZN(n17465) );
  OAI21_X1 U20696 ( .B1(n17484), .B2(n17495), .A(n17465), .ZN(P3_U2777) );
  AOI22_X1 U20697 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17497), .ZN(n17466) );
  OAI21_X1 U20698 ( .B1(n17486), .B2(n17495), .A(n17466), .ZN(P3_U2778) );
  AOI22_X1 U20699 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17497), .ZN(n17467) );
  OAI21_X1 U20700 ( .B1(n17488), .B2(n17490), .A(n17467), .ZN(P3_U2779) );
  AOI22_X1 U20701 ( .A1(P3_UWORD_REG_12__SCAN_IN), .A2(n17497), .B1(
        P3_EAX_REG_28__SCAN_IN), .B2(n9729), .ZN(n17468) );
  OAI21_X1 U20702 ( .B1(n17491), .B2(n17490), .A(n17468), .ZN(P3_U2780) );
  AOI22_X1 U20703 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17498), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17497), .ZN(n17469) );
  OAI21_X1 U20704 ( .B1(n17470), .B2(n17500), .A(n17469), .ZN(P3_U2781) );
  AOI22_X1 U20705 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n9729), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17497), .ZN(n17471) );
  OAI21_X1 U20706 ( .B1(n17496), .B2(n17490), .A(n17471), .ZN(P3_U2782) );
  AOI22_X1 U20707 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17497), .ZN(n17472) );
  OAI21_X1 U20708 ( .B1(n18200), .B2(n17490), .A(n17472), .ZN(P3_U2783) );
  AOI22_X1 U20709 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17498), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n9729), .ZN(n17473) );
  OAI21_X1 U20710 ( .B1(n17474), .B2(n20988), .A(n17473), .ZN(P3_U2784) );
  AOI22_X1 U20711 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17497), .ZN(n17475) );
  OAI21_X1 U20712 ( .B1(n18213), .B2(n17490), .A(n17475), .ZN(P3_U2785) );
  AOI22_X1 U20713 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17497), .ZN(n17476) );
  OAI21_X1 U20714 ( .B1(n18218), .B2(n17490), .A(n17476), .ZN(P3_U2786) );
  AOI22_X1 U20715 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17497), .ZN(n17477) );
  OAI21_X1 U20716 ( .B1(n18223), .B2(n17490), .A(n17477), .ZN(P3_U2787) );
  AOI22_X1 U20717 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17497), .ZN(n17478) );
  OAI21_X1 U20718 ( .B1(n20847), .B2(n17490), .A(n17478), .ZN(P3_U2788) );
  AOI22_X1 U20719 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17497), .ZN(n17479) );
  OAI21_X1 U20720 ( .B1(n18231), .B2(n17490), .A(n17479), .ZN(P3_U2789) );
  AOI22_X1 U20721 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17497), .ZN(n17480) );
  OAI21_X1 U20722 ( .B1(n18237), .B2(n17490), .A(n17480), .ZN(P3_U2790) );
  AOI22_X1 U20723 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17497), .ZN(n17481) );
  OAI21_X1 U20724 ( .B1(n17482), .B2(n17490), .A(n17481), .ZN(P3_U2791) );
  AOI22_X1 U20725 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17497), .ZN(n17483) );
  OAI21_X1 U20726 ( .B1(n17484), .B2(n17490), .A(n17483), .ZN(P3_U2792) );
  AOI22_X1 U20727 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17497), .ZN(n17485) );
  OAI21_X1 U20728 ( .B1(n17486), .B2(n17490), .A(n17485), .ZN(P3_U2793) );
  AOI22_X1 U20729 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17497), .ZN(n17487) );
  OAI21_X1 U20730 ( .B1(n17488), .B2(n17490), .A(n17487), .ZN(P3_U2794) );
  AOI22_X1 U20731 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17497), .ZN(n17489) );
  OAI21_X1 U20732 ( .B1(n17491), .B2(n17490), .A(n17489), .ZN(P3_U2795) );
  AOI22_X1 U20733 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17498), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17497), .ZN(n17492) );
  OAI21_X1 U20734 ( .B1(n17493), .B2(n17500), .A(n17492), .ZN(P3_U2796) );
  AOI22_X1 U20735 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n9729), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17497), .ZN(n17494) );
  OAI21_X1 U20736 ( .B1(n17496), .B2(n17495), .A(n17494), .ZN(P3_U2797) );
  AOI22_X1 U20737 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17498), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17497), .ZN(n17499) );
  OAI21_X1 U20738 ( .B1(n17501), .B2(n17500), .A(n17499), .ZN(P3_U2798) );
  OAI21_X1 U20739 ( .B1(n17502), .B2(n17856), .A(n17855), .ZN(n17503) );
  AOI21_X1 U20740 ( .B1(n17687), .B2(n17513), .A(n17503), .ZN(n17535) );
  OAI21_X1 U20741 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17607), .A(
        n17535), .ZN(n17527) );
  AOI22_X1 U20742 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17527), .B1(
        n17708), .B2(n17504), .ZN(n17518) );
  NAND2_X1 U20743 ( .A1(n17922), .A2(n17637), .ZN(n17622) );
  NOR2_X1 U20744 ( .A1(n17847), .A2(n17767), .ZN(n17614) );
  INV_X1 U20745 ( .A(n17767), .ZN(n17725) );
  OAI22_X1 U20746 ( .A1(n17506), .A2(n17861), .B1(n17867), .B2(n17725), .ZN(
        n17539) );
  NOR2_X1 U20747 ( .A1(n10076), .A2(n17539), .ZN(n17530) );
  NOR3_X1 U20748 ( .A1(n17614), .A2(n17530), .A3(n21105), .ZN(n17511) );
  AOI211_X1 U20749 ( .C1(n17509), .C2(n17508), .A(n17507), .B(n17741), .ZN(
        n17510) );
  AOI211_X1 U20750 ( .C1(n17512), .C2(n17574), .A(n17511), .B(n17510), .ZN(
        n17517) );
  NAND2_X1 U20751 ( .A1(n9732), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17516) );
  NOR2_X1 U20752 ( .A1(n17691), .A2(n17513), .ZN(n17520) );
  OAI211_X1 U20753 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17520), .B(n17514), .ZN(n17515) );
  NAND4_X1 U20754 ( .A1(n17518), .A2(n17517), .A3(n17516), .A4(n17515), .ZN(
        P3_U2802) );
  OAI22_X1 U20755 ( .A1(n18179), .A2(n18785), .B1(n17704), .B2(n17519), .ZN(
        n17526) );
  INV_X1 U20756 ( .A(n17520), .ZN(n17524) );
  NOR2_X1 U20757 ( .A1(n17522), .A2(n17521), .ZN(n17523) );
  XNOR2_X1 U20758 ( .A(n17523), .B(n17679), .ZN(n17875) );
  OAI22_X1 U20759 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17524), .B1(
        n17875), .B2(n17741), .ZN(n17525) );
  AOI211_X1 U20760 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17527), .A(
        n17526), .B(n17525), .ZN(n17528) );
  OAI221_X1 U20761 ( .B1(n17530), .B2(n10076), .C1(n17530), .C2(n17529), .A(
        n17528), .ZN(P3_U2803) );
  AOI21_X1 U20762 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17532), .A(
        n17531), .ZN(n17882) );
  AOI21_X1 U20763 ( .B1(n18241), .B2(n17533), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17534) );
  OAI22_X1 U20764 ( .A1(n17535), .A2(n17534), .B1(n18179), .B2(n18783), .ZN(
        n17536) );
  AOI221_X1 U20765 ( .B1(n17708), .B2(n17537), .C1(n12712), .C2(n17537), .A(
        n17536), .ZN(n17541) );
  NOR2_X1 U20766 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17538), .ZN(
        n17879) );
  AOI22_X1 U20767 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17539), .B1(
        n17574), .B2(n17879), .ZN(n17540) );
  OAI211_X1 U20768 ( .C1(n17882), .C2(n17741), .A(n17541), .B(n17540), .ZN(
        P3_U2804) );
  NAND3_X1 U20769 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17558), .A3(
        n18000), .ZN(n17542) );
  XNOR2_X1 U20770 ( .A(n17542), .B(n17896), .ZN(n17887) );
  INV_X1 U20771 ( .A(n17855), .ZN(n17842) );
  AND2_X1 U20772 ( .A1(n17544), .A2(n18241), .ZN(n17569) );
  AOI211_X1 U20773 ( .C1(n17689), .C2(n17543), .A(n17842), .B(n17569), .ZN(
        n17567) );
  OAI21_X1 U20774 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17607), .A(
        n17567), .ZN(n17555) );
  NOR2_X1 U20775 ( .A1(n17691), .A2(n17544), .ZN(n17557) );
  OAI211_X1 U20776 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17557), .B(n17545), .ZN(n17546) );
  NAND2_X1 U20777 ( .A1(n9732), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17894) );
  OAI211_X1 U20778 ( .C1(n17704), .C2(n17547), .A(n17546), .B(n17894), .ZN(
        n17553) );
  NAND2_X1 U20779 ( .A1(n17999), .A2(n17558), .ZN(n17898) );
  NOR2_X1 U20780 ( .A1(n17904), .A2(n17898), .ZN(n17548) );
  XNOR2_X1 U20781 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17548), .ZN(
        n17890) );
  OAI21_X1 U20782 ( .B1(n17679), .B2(n17550), .A(n17549), .ZN(n17551) );
  XNOR2_X1 U20783 ( .A(n17551), .B(n17896), .ZN(n17889) );
  OAI22_X1 U20784 ( .A1(n17861), .A2(n17890), .B1(n17741), .B2(n17889), .ZN(
        n17552) );
  AOI211_X1 U20785 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17555), .A(
        n17553), .B(n17552), .ZN(n17554) );
  OAI21_X1 U20786 ( .B1(n17725), .B2(n17887), .A(n17554), .ZN(P3_U2805) );
  NOR2_X1 U20787 ( .A1(n18179), .A2(n18779), .ZN(n17907) );
  AOI221_X1 U20788 ( .B1(n17557), .B2(n17556), .C1(n17555), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17907), .ZN(n17563) );
  NOR2_X1 U20789 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n20826), .ZN(
        n17909) );
  NAND2_X1 U20790 ( .A1(n18000), .A2(n17558), .ZN(n17897) );
  AOI22_X1 U20791 ( .A1(n17847), .A2(n17898), .B1(n17767), .B2(n17897), .ZN(
        n17577) );
  AOI21_X1 U20792 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17560), .A(
        n17559), .ZN(n17911) );
  OAI22_X1 U20793 ( .A1(n17577), .A2(n17904), .B1(n17911), .B2(n17741), .ZN(
        n17561) );
  AOI21_X1 U20794 ( .B1(n17574), .B2(n17909), .A(n17561), .ZN(n17562) );
  OAI211_X1 U20795 ( .C1(n17704), .C2(n17564), .A(n17563), .B(n17562), .ZN(
        P3_U2806) );
  NOR2_X1 U20796 ( .A1(n18179), .A2(n18778), .ZN(n17914) );
  NOR2_X1 U20797 ( .A1(n17708), .A2(n12712), .ZN(n17839) );
  INV_X1 U20798 ( .A(n17565), .ZN(n17566) );
  OAI22_X1 U20799 ( .A1(n17567), .A2(n9994), .B1(n17839), .B2(n17566), .ZN(
        n17568) );
  AOI211_X1 U20800 ( .C1(n17569), .C2(n9857), .A(n17914), .B(n17568), .ZN(
        n17576) );
  AOI22_X1 U20801 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17679), .B1(
        n17571), .B2(n17579), .ZN(n17572) );
  NAND2_X1 U20802 ( .A1(n17570), .A2(n17572), .ZN(n17573) );
  XNOR2_X1 U20803 ( .A(n17573), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17915) );
  AOI22_X1 U20804 ( .A1(n17915), .A2(n17766), .B1(n17574), .B2(n20826), .ZN(
        n17575) );
  OAI211_X1 U20805 ( .C1(n17577), .C2(n20826), .A(n17576), .B(n17575), .ZN(
        P3_U2807) );
  INV_X1 U20806 ( .A(n17570), .ZN(n17578) );
  AOI221_X1 U20807 ( .B1(n9744), .B2(n17579), .C1(n17931), .C2(n17579), .A(
        n17578), .ZN(n17580) );
  XNOR2_X1 U20808 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17580), .ZN(
        n17940) );
  INV_X1 U20809 ( .A(n17931), .ZN(n17590) );
  NOR2_X1 U20810 ( .A1(n18000), .A2(n17725), .ZN(n17672) );
  AOI21_X1 U20811 ( .B1(n17847), .B2(n17581), .A(n17672), .ZN(n17660) );
  OAI21_X1 U20812 ( .B1(n17590), .B2(n17614), .A(n17660), .ZN(n17603) );
  INV_X1 U20813 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18775) );
  OAI21_X1 U20814 ( .B1(n17582), .B2(n17856), .A(n17855), .ZN(n17583) );
  AOI21_X1 U20815 ( .B1(n17687), .B2(n17585), .A(n17583), .ZN(n17610) );
  OAI21_X1 U20816 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17607), .A(
        n17610), .ZN(n17596) );
  AOI22_X1 U20817 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17596), .B1(
        n17708), .B2(n17584), .ZN(n17588) );
  NOR2_X1 U20818 ( .A1(n17691), .A2(n17585), .ZN(n17598) );
  OAI211_X1 U20819 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17598), .B(n17586), .ZN(n17587) );
  OAI211_X1 U20820 ( .C1(n18775), .C2(n18179), .A(n17588), .B(n17587), .ZN(
        n17589) );
  AOI21_X1 U20821 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17603), .A(
        n17589), .ZN(n17592) );
  NAND3_X1 U20822 ( .A1(n17590), .A2(n17637), .A3(n17920), .ZN(n17591) );
  OAI211_X1 U20823 ( .C1(n17741), .C2(n17940), .A(n17592), .B(n17591), .ZN(
        P3_U2808) );
  NAND2_X1 U20824 ( .A1(n17923), .A2(n17934), .ZN(n17947) );
  INV_X1 U20825 ( .A(n17593), .ZN(n17594) );
  OAI22_X1 U20826 ( .A1(n18179), .A2(n18774), .B1(n17704), .B2(n17594), .ZN(
        n17595) );
  AOI221_X1 U20827 ( .B1(n17598), .B2(n17597), .C1(n17596), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17595), .ZN(n17605) );
  NOR3_X1 U20828 ( .A1(n17929), .A2(n17679), .A3(n17599), .ZN(n17620) );
  INV_X1 U20829 ( .A(n17600), .ZN(n17631) );
  AOI22_X1 U20830 ( .A1(n17923), .A2(n17620), .B1(n17631), .B2(n17601), .ZN(
        n17602) );
  XNOR2_X1 U20831 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17602), .ZN(
        n17941) );
  AOI22_X1 U20832 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17603), .B1(
        n17766), .B2(n17941), .ZN(n17604) );
  OAI211_X1 U20833 ( .C1(n17622), .C2(n17947), .A(n17605), .B(n17604), .ZN(
        P3_U2809) );
  NAND2_X1 U20834 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17606), .ZN(
        n17959) );
  AOI21_X1 U20835 ( .B1(n17608), .B2(n18241), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17609) );
  OAI22_X1 U20836 ( .A1(n17610), .A2(n17609), .B1(n18179), .B2(n18771), .ZN(
        n17611) );
  AOI221_X1 U20837 ( .B1(n17708), .B2(n17612), .C1(n12712), .C2(n17612), .A(
        n17611), .ZN(n17617) );
  INV_X1 U20838 ( .A(n17922), .ZN(n17613) );
  NOR2_X1 U20839 ( .A1(n17613), .A2(n17961), .ZN(n17955) );
  OAI21_X1 U20840 ( .B1(n17614), .B2(n17955), .A(n17660), .ZN(n17624) );
  OAI221_X1 U20841 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17629), 
        .C1(n17961), .C2(n17620), .A(n17570), .ZN(n17615) );
  XNOR2_X1 U20842 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17615), .ZN(
        n17948) );
  AOI22_X1 U20843 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17624), .B1(
        n17766), .B2(n17948), .ZN(n17616) );
  OAI211_X1 U20844 ( .C1(n17622), .C2(n17959), .A(n17617), .B(n17616), .ZN(
        P3_U2810) );
  AOI21_X1 U20845 ( .B1(n17687), .B2(n17625), .A(n17842), .ZN(n17642) );
  OAI21_X1 U20846 ( .B1(n17618), .B2(n17856), .A(n17642), .ZN(n17634) );
  AOI22_X1 U20847 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17634), .B1(
        n17708), .B2(n17619), .ZN(n17628) );
  AOI21_X1 U20848 ( .B1(n17631), .B2(n17629), .A(n17620), .ZN(n17621) );
  XNOR2_X1 U20849 ( .A(n17621), .B(n17961), .ZN(n17966) );
  OAI22_X1 U20850 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17622), .B1(
        n17966), .B2(n17741), .ZN(n17623) );
  AOI21_X1 U20851 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17624), .A(
        n17623), .ZN(n17627) );
  NAND2_X1 U20852 ( .A1(n9732), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17964) );
  NOR2_X1 U20853 ( .A1(n17691), .A2(n17625), .ZN(n17636) );
  OAI211_X1 U20854 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17636), .B(n9860), .ZN(n17626)
         );
  NAND4_X1 U20855 ( .A1(n17628), .A2(n17627), .A3(n17964), .A4(n17626), .ZN(
        P3_U2811) );
  AOI21_X1 U20856 ( .B1(n17765), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17629), .ZN(n17630) );
  XNOR2_X1 U20857 ( .A(n17631), .B(n17630), .ZN(n17979) );
  OAI22_X1 U20858 ( .A1(n18179), .A2(n18767), .B1(n17704), .B2(n17632), .ZN(
        n17633) );
  AOI221_X1 U20859 ( .B1(n17636), .B2(n17635), .C1(n17634), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17633), .ZN(n17639) );
  INV_X1 U20860 ( .A(n17637), .ZN(n17661) );
  OAI21_X1 U20861 ( .B1(n17926), .B2(n17661), .A(n17660), .ZN(n17647) );
  NOR2_X1 U20862 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17972), .ZN(
        n17975) );
  AOI22_X1 U20863 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17647), .B1(
        n17637), .B2(n17975), .ZN(n17638) );
  OAI211_X1 U20864 ( .C1(n17741), .C2(n17979), .A(n17639), .B(n17638), .ZN(
        P3_U2812) );
  NAND2_X1 U20865 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17981), .ZN(
        n17987) );
  AOI21_X1 U20866 ( .B1(n17640), .B2(n18241), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17643) );
  OAI22_X1 U20867 ( .A1(n17643), .A2(n17642), .B1(n17839), .B2(n17641), .ZN(
        n17644) );
  AOI21_X1 U20868 ( .B1(n9732), .B2(P3_REIP_REG_17__SCAN_IN), .A(n17644), .ZN(
        n17649) );
  OAI21_X1 U20869 ( .B1(n17646), .B2(n17981), .A(n17645), .ZN(n17984) );
  AOI22_X1 U20870 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17647), .B1(
        n17766), .B2(n17984), .ZN(n17648) );
  OAI211_X1 U20871 ( .C1(n17661), .C2(n17987), .A(n17649), .B(n17648), .ZN(
        P3_U2813) );
  AOI21_X1 U20872 ( .B1(n17765), .B2(n9744), .A(n17650), .ZN(n17651) );
  XNOR2_X1 U20873 ( .A(n17651), .B(n17967), .ZN(n17994) );
  AOI21_X1 U20874 ( .B1(n17687), .B2(n17654), .A(n17842), .ZN(n17678) );
  OAI21_X1 U20875 ( .B1(n17652), .B2(n17856), .A(n17678), .ZN(n17668) );
  AOI22_X1 U20876 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17668), .B1(
        n17708), .B2(n17653), .ZN(n17657) );
  NAND2_X1 U20877 ( .A1(n9732), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17996) );
  NOR2_X1 U20878 ( .A1(n17691), .A2(n17654), .ZN(n17670) );
  OAI211_X1 U20879 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17670), .B(n17655), .ZN(n17656) );
  NAND3_X1 U20880 ( .A1(n17657), .A2(n17996), .A3(n17656), .ZN(n17658) );
  AOI21_X1 U20881 ( .B1(n17766), .B2(n17994), .A(n17658), .ZN(n17659) );
  OAI221_X1 U20882 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17661), 
        .C1(n17967), .C2(n17660), .A(n17659), .ZN(P3_U2814) );
  INV_X1 U20883 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18029) );
  INV_X1 U20884 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18043) );
  NAND3_X1 U20885 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n18051), .ZN(n17663) );
  OAI21_X1 U20886 ( .B1(n17696), .B2(n17663), .A(n17662), .ZN(n17664) );
  OAI221_X1 U20887 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18029), 
        .C1(n18043), .C2(n17765), .A(n17664), .ZN(n17665) );
  XNOR2_X1 U20888 ( .A(n18013), .B(n17665), .ZN(n18006) );
  OAI22_X1 U20889 ( .A1(n18179), .A2(n18762), .B1(n17704), .B2(n17666), .ZN(
        n17667) );
  AOI221_X1 U20890 ( .B1(n17670), .B2(n17669), .C1(n17668), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17667), .ZN(n17675) );
  NOR2_X1 U20891 ( .A1(n17999), .A2(n17861), .ZN(n17673) );
  NAND2_X1 U20892 ( .A1(n18017), .A2(n18056), .ZN(n17676) );
  OAI21_X1 U20893 ( .B1(n18029), .B2(n17676), .A(n18013), .ZN(n18009) );
  INV_X1 U20894 ( .A(n18002), .ZN(n17671) );
  NAND2_X1 U20895 ( .A1(n17671), .A2(n17726), .ZN(n17682) );
  NAND2_X1 U20896 ( .A1(n18013), .A2(n17682), .ZN(n18004) );
  AOI22_X1 U20897 ( .A1(n17673), .A2(n18009), .B1(n17672), .B2(n18004), .ZN(
        n17674) );
  OAI211_X1 U20898 ( .C1(n17741), .C2(n18006), .A(n17675), .B(n17674), .ZN(
        P3_U2815) );
  XOR2_X1 U20899 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17676), .Z(
        n18024) );
  NOR2_X1 U20900 ( .A1(n18356), .A2(n9869), .ZN(n17721) );
  AOI21_X1 U20901 ( .B1(n17692), .B2(n17721), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17677) );
  NAND2_X1 U20902 ( .A1(n9732), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n18031) );
  OAI21_X1 U20903 ( .B1(n17678), .B2(n17677), .A(n18031), .ZN(n17684) );
  NOR2_X1 U20904 ( .A1(n17679), .A2(n18053), .ZN(n17730) );
  AOI21_X1 U20905 ( .B1(n18017), .B2(n17730), .A(n17680), .ZN(n17681) );
  XOR2_X1 U20906 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17681), .Z(
        n18028) );
  OAI221_X1 U20907 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18017), 
        .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17726), .A(n17682), .ZN(
        n18022) );
  OAI22_X1 U20908 ( .A1(n18028), .A2(n17741), .B1(n17725), .B2(n18022), .ZN(
        n17683) );
  AOI211_X1 U20909 ( .C1(n17685), .C2(n17849), .A(n17684), .B(n17683), .ZN(
        n17686) );
  OAI21_X1 U20910 ( .B1(n17861), .B2(n18024), .A(n17686), .ZN(P3_U2816) );
  AOI22_X1 U20911 ( .A1(n17689), .A2(n17688), .B1(n17687), .B2(n9869), .ZN(
        n17690) );
  NAND2_X1 U20912 ( .A1(n17690), .A2(n17855), .ZN(n17709) );
  OR2_X1 U20913 ( .A1(n9869), .A2(n17691), .ZN(n17711) );
  AOI211_X1 U20914 ( .C1(n20927), .C2(n17693), .A(n17692), .B(n17711), .ZN(
        n17695) );
  NOR2_X1 U20915 ( .A1(n18179), .A2(n18758), .ZN(n17694) );
  AOI211_X1 U20916 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17709), .A(
        n17695), .B(n17694), .ZN(n17702) );
  OAI22_X1 U20917 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17765), .B1(
        n17696), .B2(n18016), .ZN(n17697) );
  OAI21_X1 U20918 ( .B1(n17765), .B2(n9833), .A(n17697), .ZN(n17698) );
  XNOR2_X1 U20919 ( .A(n17698), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18034) );
  INV_X1 U20920 ( .A(n18016), .ZN(n17699) );
  NAND2_X1 U20921 ( .A1(n17699), .A2(n20895), .ZN(n18042) );
  NAND2_X1 U20922 ( .A1(n17699), .A2(n18056), .ZN(n18036) );
  NAND2_X1 U20923 ( .A1(n17699), .A2(n17726), .ZN(n18035) );
  AOI22_X1 U20924 ( .A1(n17847), .A2(n18036), .B1(n17767), .B2(n18035), .ZN(
        n17715) );
  OAI22_X1 U20925 ( .A1(n17754), .A2(n18042), .B1(n17715), .B2(n20895), .ZN(
        n17700) );
  AOI21_X1 U20926 ( .B1(n17766), .B2(n18034), .A(n17700), .ZN(n17701) );
  OAI211_X1 U20927 ( .C1(n17704), .C2(n17703), .A(n17702), .B(n17701), .ZN(
        P3_U2817) );
  AOI21_X1 U20928 ( .B1(n18051), .B2(n17730), .A(n9833), .ZN(n17705) );
  XNOR2_X1 U20929 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n17705), .ZN(
        n18046) );
  NOR3_X1 U20930 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17754), .A3(
        n17706), .ZN(n17713) );
  AOI22_X1 U20931 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17709), .B1(
        n17708), .B2(n17707), .ZN(n17710) );
  NAND2_X1 U20932 ( .A1(n9732), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18047) );
  OAI211_X1 U20933 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n17711), .A(
        n17710), .B(n18047), .ZN(n17712) );
  AOI211_X1 U20934 ( .C1(n17766), .C2(n18046), .A(n17713), .B(n17712), .ZN(
        n17714) );
  OAI21_X1 U20935 ( .B1(n17715), .B2(n18043), .A(n17714), .ZN(P3_U2818) );
  OR2_X1 U20936 ( .A1(n18059), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18064) );
  INV_X1 U20937 ( .A(n17730), .ZN(n17744) );
  OAI21_X1 U20938 ( .B1(n18059), .B2(n17744), .A(n17716), .ZN(n17717) );
  XOR2_X1 U20939 ( .A(n17717), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18050) );
  NOR2_X1 U20940 ( .A1(n18179), .A2(n18754), .ZN(n17723) );
  NOR3_X1 U20941 ( .A1(n18356), .A2(n17746), .A3(n17718), .ZN(n17749) );
  AND2_X1 U20942 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17749), .ZN(
        n17735) );
  AOI21_X1 U20943 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17850), .A(
        n17735), .ZN(n17720) );
  OAI22_X1 U20944 ( .A1(n17721), .A2(n17720), .B1(n17839), .B2(n17719), .ZN(
        n17722) );
  AOI211_X1 U20945 ( .C1(n17766), .C2(n18050), .A(n17723), .B(n17722), .ZN(
        n17728) );
  NOR2_X1 U20946 ( .A1(n17724), .A2(n17754), .ZN(n17738) );
  OAI22_X1 U20947 ( .A1(n17726), .A2(n17725), .B1(n17861), .B2(n18056), .ZN(
        n17742) );
  OAI21_X1 U20948 ( .B1(n17738), .B2(n17742), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17727) );
  OAI211_X1 U20949 ( .C1(n17754), .C2(n18064), .A(n17728), .B(n17727), .ZN(
        P3_U2819) );
  AOI21_X1 U20950 ( .B1(n17730), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17729), .ZN(n17732) );
  XNOR2_X1 U20951 ( .A(n17732), .B(n17731), .ZN(n18073) );
  NOR2_X1 U20952 ( .A1(n18179), .A2(n18753), .ZN(n17737) );
  AOI21_X1 U20953 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17850), .A(
        n17749), .ZN(n17734) );
  OAI22_X1 U20954 ( .A1(n17735), .A2(n17734), .B1(n17839), .B2(n17733), .ZN(
        n17736) );
  AOI211_X1 U20955 ( .C1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n17742), .A(
        n17737), .B(n17736), .ZN(n17740) );
  OAI21_X1 U20956 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17738), .ZN(n17739) );
  OAI211_X1 U20957 ( .C1(n18073), .C2(n17741), .A(n17740), .B(n17739), .ZN(
        P3_U2820) );
  INV_X1 U20958 ( .A(n17742), .ZN(n17753) );
  NAND2_X1 U20959 ( .A1(n17744), .A2(n17743), .ZN(n17745) );
  XOR2_X1 U20960 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n17745), .Z(
        n18074) );
  NOR2_X1 U20961 ( .A1(n18179), .A2(n18751), .ZN(n17751) );
  NOR2_X1 U20962 ( .A1(n17773), .A2(n17760), .ZN(n17758) );
  NOR2_X1 U20963 ( .A1(n18356), .A2(n17746), .ZN(n17774) );
  AOI22_X1 U20964 ( .A1(n17758), .A2(n17774), .B1(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17850), .ZN(n17748) );
  OAI22_X1 U20965 ( .A1(n17749), .A2(n17748), .B1(n17839), .B2(n17747), .ZN(
        n17750) );
  AOI211_X1 U20966 ( .C1(n17766), .C2(n18074), .A(n17751), .B(n17750), .ZN(
        n17752) );
  OAI221_X1 U20967 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17754), .C1(
        n10082), .C2(n17753), .A(n17752), .ZN(P3_U2821) );
  OAI21_X1 U20968 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17756), .A(
        n17755), .ZN(n18095) );
  OAI21_X1 U20969 ( .B1(n17757), .B2(n17822), .A(n17855), .ZN(n17772) );
  AOI211_X1 U20970 ( .C1(n17760), .C2(n17759), .A(n17758), .B(n18356), .ZN(
        n17763) );
  NAND2_X1 U20971 ( .A1(n9732), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18100) );
  OAI21_X1 U20972 ( .B1(n17839), .B2(n17761), .A(n18100), .ZN(n17762) );
  AOI211_X1 U20973 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17772), .A(
        n17763), .B(n17762), .ZN(n17769) );
  OAI21_X1 U20974 ( .B1(n17765), .B2(n18093), .A(n17764), .ZN(n18098) );
  AOI22_X1 U20975 ( .A1(n17767), .A2(n18093), .B1(n17766), .B2(n18098), .ZN(
        n17768) );
  OAI211_X1 U20976 ( .C1(n17861), .C2(n18095), .A(n17769), .B(n17768), .ZN(
        P3_U2822) );
  OAI21_X1 U20977 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17771), .A(
        n17770), .ZN(n18111) );
  NOR2_X1 U20978 ( .A1(n18179), .A2(n18750), .ZN(n18108) );
  AOI221_X1 U20979 ( .B1(n17774), .B2(n17773), .C1(n17772), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18108), .ZN(n17781) );
  AOI21_X1 U20980 ( .B1(n17777), .B2(n17776), .A(n17775), .ZN(n17778) );
  XNOR2_X1 U20981 ( .A(n17778), .B(n18106), .ZN(n18109) );
  AOI22_X1 U20982 ( .A1(n17847), .A2(n18109), .B1(n17779), .B2(n17849), .ZN(
        n17780) );
  OAI211_X1 U20983 ( .C1(n17860), .C2(n18111), .A(n17781), .B(n17780), .ZN(
        P3_U2823) );
  OAI21_X1 U20984 ( .B1(n17783), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17782), .ZN(n18115) );
  NAND2_X1 U20985 ( .A1(n18241), .A2(n17790), .ZN(n17787) );
  OAI21_X1 U20986 ( .B1(n17786), .B2(n17785), .A(n17784), .ZN(n18114) );
  OAI22_X1 U20987 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17787), .B1(
        n17860), .B2(n18114), .ZN(n17788) );
  AOI21_X1 U20988 ( .B1(n9732), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17788), .ZN(
        n17793) );
  INV_X1 U20989 ( .A(n17850), .ZN(n17789) );
  AOI21_X1 U20990 ( .B1(n17790), .B2(n18241), .A(n17789), .ZN(n17805) );
  AOI22_X1 U20991 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17805), .B1(
        n17791), .B2(n17849), .ZN(n17792) );
  OAI211_X1 U20992 ( .C1(n17861), .C2(n18115), .A(n17793), .B(n17792), .ZN(
        P3_U2824) );
  OAI21_X1 U20993 ( .B1(n17796), .B2(n17795), .A(n17794), .ZN(n18127) );
  OAI21_X1 U20994 ( .B1(n17842), .B2(n17797), .A(n20943), .ZN(n17804) );
  OAI21_X1 U20995 ( .B1(n17800), .B2(n17799), .A(n17798), .ZN(n17801) );
  XNOR2_X1 U20996 ( .A(n17801), .B(n21107), .ZN(n18121) );
  OAI22_X1 U20997 ( .A1(n17839), .A2(n17802), .B1(n17860), .B2(n18121), .ZN(
        n17803) );
  AOI21_X1 U20998 ( .B1(n17805), .B2(n17804), .A(n17803), .ZN(n17806) );
  NAND2_X1 U20999 ( .A1(n9732), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18125) );
  OAI211_X1 U21000 ( .C1(n17861), .C2(n18127), .A(n17806), .B(n18125), .ZN(
        P3_U2825) );
  OAI21_X1 U21001 ( .B1(n17809), .B2(n17808), .A(n17807), .ZN(n18134) );
  OAI21_X1 U21002 ( .B1(n17812), .B2(n17811), .A(n17810), .ZN(n18133) );
  OAI22_X1 U21003 ( .A1(n17861), .A2(n18133), .B1(n18356), .B2(n17813), .ZN(
        n17814) );
  AOI21_X1 U21004 ( .B1(n9732), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17814), .ZN(
        n17818) );
  OAI21_X1 U21005 ( .B1(n17815), .B2(n17822), .A(n17855), .ZN(n17823) );
  AOI22_X1 U21006 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17823), .B1(
        n17816), .B2(n17849), .ZN(n17817) );
  OAI211_X1 U21007 ( .C1(n17860), .C2(n18134), .A(n17818), .B(n17817), .ZN(
        P3_U2826) );
  OAI21_X1 U21008 ( .B1(n17821), .B2(n17820), .A(n17819), .ZN(n18144) );
  NOR4_X1 U21009 ( .A1(n17842), .A2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        n17841), .A4(n17822), .ZN(n17829) );
  INV_X1 U21010 ( .A(n17823), .ZN(n17827) );
  OAI21_X1 U21011 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17825), .A(
        n17824), .ZN(n18143) );
  OAI22_X1 U21012 ( .A1(n17827), .A2(n17826), .B1(n17860), .B2(n18143), .ZN(
        n17828) );
  AOI211_X1 U21013 ( .C1(n17830), .C2(n17849), .A(n17829), .B(n17828), .ZN(
        n17831) );
  NAND2_X1 U21014 ( .A1(n9732), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18149) );
  OAI211_X1 U21015 ( .C1(n17861), .C2(n18144), .A(n17831), .B(n18149), .ZN(
        P3_U2827) );
  OAI21_X1 U21016 ( .B1(n17834), .B2(n17833), .A(n17832), .ZN(n18161) );
  OAI21_X1 U21017 ( .B1(n17837), .B2(n17836), .A(n17835), .ZN(n18167) );
  OAI22_X1 U21018 ( .A1(n17839), .A2(n17838), .B1(n17860), .B2(n18167), .ZN(
        n17840) );
  AOI221_X1 U21019 ( .B1(n17842), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18241), .C2(n17841), .A(n17840), .ZN(n17843) );
  NAND2_X1 U21020 ( .A1(n9732), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18165) );
  OAI211_X1 U21021 ( .C1(n17861), .C2(n18161), .A(n17843), .B(n18165), .ZN(
        P3_U2828) );
  OAI21_X1 U21022 ( .B1(n17845), .B2(n17853), .A(n17844), .ZN(n18178) );
  NAND2_X1 U21023 ( .A1(n18838), .A2(n17854), .ZN(n17846) );
  XNOR2_X1 U21024 ( .A(n17846), .B(n17845), .ZN(n18174) );
  AOI22_X1 U21025 ( .A1(n17847), .A2(n18174), .B1(n9732), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17852) );
  AOI22_X1 U21026 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17850), .B1(
        n17849), .B2(n17848), .ZN(n17851) );
  OAI211_X1 U21027 ( .C1(n17860), .C2(n18178), .A(n17852), .B(n17851), .ZN(
        P3_U2829) );
  AOI21_X1 U21028 ( .B1(n17854), .B2(n18838), .A(n17853), .ZN(n18183) );
  INV_X1 U21029 ( .A(n18183), .ZN(n18181) );
  NAND3_X1 U21030 ( .A1(n17857), .A2(n17856), .A3(n17855), .ZN(n17858) );
  AOI22_X1 U21031 ( .A1(n9732), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17858), .ZN(n17859) );
  OAI221_X1 U21032 ( .B1(n18183), .B2(n17861), .C1(n18181), .C2(n17860), .A(
        n17859), .ZN(P3_U2830) );
  INV_X1 U21033 ( .A(n17912), .ZN(n17919) );
  NOR2_X1 U21034 ( .A1(n17862), .A2(n17919), .ZN(n17871) );
  NOR2_X1 U21035 ( .A1(n18673), .A2(n18015), .ZN(n18153) );
  NOR2_X1 U21036 ( .A1(n18670), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18157) );
  NOR2_X1 U21037 ( .A1(n18157), .A2(n17863), .ZN(n17900) );
  OAI221_X1 U21038 ( .B1(n18153), .B2(n17883), .C1(n18153), .C2(n17900), .A(
        n17901), .ZN(n17885) );
  INV_X1 U21039 ( .A(n18153), .ZN(n18128) );
  NAND2_X1 U21040 ( .A1(n17864), .A2(n18128), .ZN(n17866) );
  OAI211_X1 U21041 ( .C1(n17867), .C2(n18023), .A(n17866), .B(n17865), .ZN(
        n17868) );
  AOI211_X1 U21042 ( .C1(n9766), .C2(n17869), .A(n17885), .B(n17868), .ZN(
        n17877) );
  INV_X1 U21043 ( .A(n17877), .ZN(n17870) );
  MUX2_X1 U21044 ( .A(n17871), .B(n17870), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17872) );
  AOI22_X1 U21045 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18164), .B1(
        n18163), .B2(n17872), .ZN(n17874) );
  NAND2_X1 U21046 ( .A1(n9732), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17873) );
  OAI211_X1 U21047 ( .C1(n17875), .C2(n18072), .A(n17874), .B(n17873), .ZN(
        P3_U2835) );
  AOI211_X1 U21048 ( .C1(n18163), .C2(n17877), .A(n9732), .B(n17876), .ZN(
        n17878) );
  AOI21_X1 U21049 ( .B1(n17879), .B2(n17908), .A(n17878), .ZN(n17881) );
  NAND2_X1 U21050 ( .A1(n9732), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17880) );
  OAI211_X1 U21051 ( .C1(n17882), .C2(n18072), .A(n17881), .B(n17880), .ZN(
        P3_U2836) );
  INV_X1 U21052 ( .A(n17883), .ZN(n17886) );
  NOR3_X1 U21053 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17884), .A3(
        n17886), .ZN(n17893) );
  AOI21_X1 U21054 ( .B1(n18658), .B2(n17886), .A(n17885), .ZN(n17888) );
  OAI22_X1 U21055 ( .A1(n17888), .A2(n17896), .B1(n18023), .B2(n17887), .ZN(
        n17892) );
  OAI22_X1 U21056 ( .A1(n18145), .A2(n17890), .B1(n18072), .B2(n17889), .ZN(
        n17891) );
  AOI221_X1 U21057 ( .B1(n17893), .B2(n18163), .C1(n17892), .C2(n18163), .A(
        n17891), .ZN(n17895) );
  OAI211_X1 U21058 ( .C1(n18169), .C2(n17896), .A(n17895), .B(n17894), .ZN(
        P3_U2837) );
  AOI22_X1 U21059 ( .A1(n9766), .A2(n17898), .B1(n18094), .B2(n17897), .ZN(
        n17899) );
  OAI211_X1 U21060 ( .C1(n18153), .C2(n17900), .A(n17899), .B(n18169), .ZN(
        n17903) );
  INV_X1 U21061 ( .A(n17903), .ZN(n17905) );
  NAND2_X1 U21062 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17901), .ZN(
        n17902) );
  OAI21_X1 U21063 ( .B1(n17903), .B2(n17902), .A(n18179), .ZN(n17918) );
  AOI211_X1 U21064 ( .C1(n17993), .C2(n17905), .A(n17904), .B(n17918), .ZN(
        n17906) );
  AOI211_X1 U21065 ( .C1(n17909), .C2(n17908), .A(n17907), .B(n17906), .ZN(
        n17910) );
  OAI21_X1 U21066 ( .B1(n17911), .B2(n18072), .A(n17910), .ZN(P3_U2838) );
  NAND3_X1 U21067 ( .A1(n17913), .A2(n17912), .A3(n18169), .ZN(n17917) );
  AOI21_X1 U21068 ( .B1(n17915), .B2(n18099), .A(n17914), .ZN(n17916) );
  OAI221_X1 U21069 ( .B1(n17918), .B2(n20826), .C1(n17918), .C2(n17917), .A(
        n17916), .ZN(P3_U2839) );
  AOI221_X1 U21070 ( .B1(n17931), .B2(n17920), .C1(n17919), .C2(n17920), .A(
        n18185), .ZN(n17937) );
  NAND2_X1 U21071 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17921), .ZN(
        n18052) );
  NOR2_X1 U21072 ( .A1(n17974), .A2(n18052), .ZN(n17988) );
  AOI21_X1 U21073 ( .B1(n17922), .B2(n17988), .A(n18670), .ZN(n17952) );
  INV_X1 U21074 ( .A(n17923), .ZN(n17924) );
  NOR2_X1 U21075 ( .A1(n17952), .A2(n17924), .ZN(n17943) );
  NAND2_X1 U21076 ( .A1(n9765), .A2(n18023), .ZN(n18058) );
  INV_X1 U21077 ( .A(n18658), .ZN(n18688) );
  AOI21_X1 U21078 ( .B1(n17926), .B2(n17925), .A(n18688), .ZN(n17971) );
  AOI21_X1 U21079 ( .B1(n17927), .B2(n17955), .A(n18171), .ZN(n17928) );
  AOI211_X1 U21080 ( .C1(n18658), .C2(n17929), .A(n17971), .B(n17928), .ZN(
        n17949) );
  OAI21_X1 U21081 ( .B1(n18171), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n17949), .ZN(n17930) );
  AOI21_X1 U21082 ( .B1(n17931), .B2(n18058), .A(n17930), .ZN(n17942) );
  AOI21_X1 U21083 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18688), .A(
        n17932), .ZN(n17933) );
  OAI22_X1 U21084 ( .A1(n17999), .A2(n9765), .B1(n18000), .B2(n18023), .ZN(
        n17951) );
  AOI211_X1 U21085 ( .C1(n17934), .C2(n18128), .A(n17933), .B(n17951), .ZN(
        n17935) );
  OAI211_X1 U21086 ( .C1(n18670), .C2(n17943), .A(n17942), .B(n17935), .ZN(
        n17936) );
  AOI22_X1 U21087 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18164), .B1(
        n17937), .B2(n17936), .ZN(n17939) );
  NAND2_X1 U21088 ( .A1(n9732), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17938) );
  OAI211_X1 U21089 ( .C1(n17940), .C2(n18072), .A(n17939), .B(n17938), .ZN(
        P3_U2840) );
  AOI22_X1 U21090 ( .A1(n9732), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18099), 
        .B2(n17941), .ZN(n17946) );
  NOR2_X1 U21091 ( .A1(n18658), .A2(n18015), .ZN(n18168) );
  OAI211_X1 U21092 ( .C1(n18168), .C2(n17943), .A(n17992), .B(n17942), .ZN(
        n17944) );
  NAND3_X1 U21093 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18179), .A3(
        n17944), .ZN(n17945) );
  OAI211_X1 U21094 ( .C1(n17947), .C2(n17960), .A(n17946), .B(n17945), .ZN(
        P3_U2841) );
  AOI22_X1 U21095 ( .A1(n9732), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18099), 
        .B2(n17948), .ZN(n17958) );
  INV_X1 U21096 ( .A(n17949), .ZN(n17950) );
  NOR4_X1 U21097 ( .A1(n18164), .A2(n17952), .A3(n17951), .A4(n17950), .ZN(
        n17954) );
  INV_X1 U21098 ( .A(n18058), .ZN(n17953) );
  AOI221_X1 U21099 ( .B1(n17955), .B2(n17954), .C1(n17953), .C2(n17954), .A(
        n9732), .ZN(n17963) );
  NOR3_X1 U21100 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18168), .A3(
        n18856), .ZN(n17956) );
  OAI21_X1 U21101 ( .B1(n17963), .B2(n17956), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17957) );
  OAI211_X1 U21102 ( .C1(n17959), .C2(n17960), .A(n17958), .B(n17957), .ZN(
        P3_U2842) );
  INV_X1 U21103 ( .A(n17960), .ZN(n17962) );
  AOI22_X1 U21104 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17963), .B1(
        n17962), .B2(n17961), .ZN(n17965) );
  OAI211_X1 U21105 ( .C1(n17966), .C2(n18072), .A(n17965), .B(n17964), .ZN(
        P3_U2843) );
  NOR3_X1 U21106 ( .A1(n18157), .A2(n17968), .A3(n17967), .ZN(n17969) );
  OAI21_X1 U21107 ( .B1(n18153), .B2(n17969), .A(n17992), .ZN(n17970) );
  AOI221_X1 U21108 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17982), 
        .C1(n18153), .C2(n17982), .A(n9732), .ZN(n17976) );
  NAND2_X1 U21109 ( .A1(n17973), .A2(n18020), .ZN(n18045) );
  NAND2_X1 U21110 ( .A1(n18163), .A2(n18045), .ZN(n18083) );
  NOR2_X1 U21111 ( .A1(n17974), .A2(n18083), .ZN(n17980) );
  AOI22_X1 U21112 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17976), .B1(
        n17975), .B2(n17980), .ZN(n17978) );
  NAND2_X1 U21113 ( .A1(n9732), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17977) );
  OAI211_X1 U21114 ( .C1(n17979), .C2(n18072), .A(n17978), .B(n17977), .ZN(
        P3_U2844) );
  INV_X1 U21115 ( .A(n17980), .ZN(n17998) );
  NOR3_X1 U21116 ( .A1(n9732), .A2(n17982), .A3(n17981), .ZN(n17983) );
  AOI21_X1 U21117 ( .B1(n18099), .B2(n17984), .A(n17983), .ZN(n17986) );
  NAND2_X1 U21118 ( .A1(n9732), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17985) );
  OAI211_X1 U21119 ( .C1(n17987), .C2(n17998), .A(n17986), .B(n17985), .ZN(
        P3_U2845) );
  AOI21_X1 U21120 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18670), .A(
        n17988), .ZN(n17991) );
  INV_X1 U21121 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18102) );
  NAND2_X1 U21122 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18091) );
  OAI21_X1 U21123 ( .B1(n18084), .B2(n18091), .A(n18673), .ZN(n17989) );
  INV_X1 U21124 ( .A(n17989), .ZN(n18080) );
  AOI21_X1 U21125 ( .B1(n18673), .B2(n18102), .A(n18080), .ZN(n18067) );
  OAI21_X1 U21126 ( .B1(n17990), .B2(n18688), .A(n18067), .ZN(n18014) );
  AOI211_X1 U21127 ( .C1(n18018), .C2(n18002), .A(n17991), .B(n18014), .ZN(
        n18001) );
  AOI221_X1 U21128 ( .B1(n17993), .B2(n17992), .C1(n18001), .C2(n17992), .A(
        n9732), .ZN(n17995) );
  AOI22_X1 U21129 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17995), .B1(
        n18099), .B2(n17994), .ZN(n17997) );
  OAI211_X1 U21130 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17998), .A(
        n17997), .B(n17996), .ZN(P3_U2846) );
  NOR2_X1 U21131 ( .A1(n17999), .A2(n18145), .ZN(n18010) );
  NOR2_X1 U21132 ( .A1(n18000), .A2(n18023), .ZN(n18005) );
  AOI221_X1 U21133 ( .B1(n18002), .B2(n18013), .C1(n18020), .C2(n18013), .A(
        n18001), .ZN(n18003) );
  AOI21_X1 U21134 ( .B1(n18005), .B2(n18004), .A(n18003), .ZN(n18007) );
  OAI22_X1 U21135 ( .A1(n18007), .A2(n18185), .B1(n18072), .B2(n18006), .ZN(
        n18008) );
  AOI21_X1 U21136 ( .B1(n18010), .B2(n18009), .A(n18008), .ZN(n18012) );
  NAND2_X1 U21137 ( .A1(n9732), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18011) );
  OAI211_X1 U21138 ( .C1(n18169), .C2(n18013), .A(n18012), .B(n18011), .ZN(
        P3_U2847) );
  AOI221_X1 U21139 ( .B1(n18016), .B2(n18015), .C1(n18052), .C2(n18015), .A(
        n18014), .ZN(n18038) );
  INV_X1 U21140 ( .A(n18017), .ZN(n18021) );
  NAND2_X1 U21141 ( .A1(n18018), .A2(n18021), .ZN(n18019) );
  OAI211_X1 U21142 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18168), .A(
        n18038), .B(n18019), .ZN(n18027) );
  NOR3_X1 U21143 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18021), .A3(
        n18020), .ZN(n18026) );
  OAI22_X1 U21144 ( .A1(n9765), .A2(n18024), .B1(n18023), .B2(n18022), .ZN(
        n18025) );
  AOI211_X1 U21145 ( .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18027), .A(
        n18026), .B(n18025), .ZN(n18033) );
  OAI22_X1 U21146 ( .A1(n18029), .A2(n18169), .B1(n18072), .B2(n18028), .ZN(
        n18030) );
  INV_X1 U21147 ( .A(n18030), .ZN(n18032) );
  OAI211_X1 U21148 ( .C1(n18033), .C2(n18185), .A(n18032), .B(n18031), .ZN(
        P3_U2848) );
  AOI22_X1 U21149 ( .A1(n9732), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18099), 
        .B2(n18034), .ZN(n18041) );
  AOI22_X1 U21150 ( .A1(n9766), .A2(n18036), .B1(n18094), .B2(n18035), .ZN(
        n18037) );
  OAI211_X1 U21151 ( .C1(n18068), .C2(n18051), .A(n18038), .B(n18037), .ZN(
        n18044) );
  OAI21_X1 U21152 ( .B1(n18068), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18163), .ZN(n18039) );
  OAI211_X1 U21153 ( .C1(n18044), .C2(n18039), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18179), .ZN(n18040) );
  OAI211_X1 U21154 ( .C1(n18083), .C2(n18042), .A(n18041), .B(n18040), .ZN(
        P3_U2849) );
  OAI222_X1 U21155 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18051), 
        .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18045), .C1(n18044), 
        .C2(n18043), .ZN(n18049) );
  AOI22_X1 U21156 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18164), .B1(
        n18099), .B2(n18046), .ZN(n18048) );
  OAI211_X1 U21157 ( .C1(n18185), .C2(n18049), .A(n18048), .B(n18047), .ZN(
        P3_U2850) );
  AOI22_X1 U21158 ( .A1(n9732), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18099), 
        .B2(n18050), .ZN(n18063) );
  NOR2_X1 U21159 ( .A1(n18068), .A2(n18051), .ZN(n18061) );
  INV_X1 U21160 ( .A(n18052), .ZN(n18078) );
  AOI21_X1 U21161 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18078), .A(
        n18670), .ZN(n18057) );
  AOI22_X1 U21162 ( .A1(n18658), .A2(n18054), .B1(n18094), .B2(n18053), .ZN(
        n18055) );
  OAI211_X1 U21163 ( .C1(n9765), .C2(n18056), .A(n18163), .B(n18055), .ZN(
        n18075) );
  AOI211_X1 U21164 ( .C1(n18059), .C2(n18058), .A(n18057), .B(n18075), .ZN(
        n18066) );
  OAI211_X1 U21165 ( .C1(n18670), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18067), .B(n18066), .ZN(n18060) );
  OAI211_X1 U21166 ( .C1(n18061), .C2(n18060), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18179), .ZN(n18062) );
  OAI211_X1 U21167 ( .C1(n18064), .C2(n18083), .A(n18063), .B(n18062), .ZN(
        P3_U2851) );
  NOR2_X1 U21168 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18083), .ZN(
        n18065) );
  AOI22_X1 U21169 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18065), .B1(
        n9732), .B2(P3_REIP_REG_10__SCAN_IN), .ZN(n18071) );
  OAI211_X1 U21170 ( .C1(n18068), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18067), .B(n18066), .ZN(n18069) );
  NAND3_X1 U21171 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18179), .A3(
        n18069), .ZN(n18070) );
  OAI211_X1 U21172 ( .C1(n18073), .C2(n18072), .A(n18071), .B(n18070), .ZN(
        P3_U2852) );
  AOI22_X1 U21173 ( .A1(n9732), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18099), .B2(
        n18074), .ZN(n18082) );
  NAND2_X1 U21174 ( .A1(n18673), .A2(n18102), .ZN(n18077) );
  INV_X1 U21175 ( .A(n18075), .ZN(n18076) );
  OAI211_X1 U21176 ( .C1(n18078), .C2(n18670), .A(n18077), .B(n18076), .ZN(
        n18079) );
  OAI211_X1 U21177 ( .C1(n18080), .C2(n18079), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n18179), .ZN(n18081) );
  OAI211_X1 U21178 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18083), .A(
        n18082), .B(n18081), .ZN(P3_U2853) );
  AOI21_X1 U21179 ( .B1(n18084), .B2(n18128), .A(n18157), .ZN(n18085) );
  OAI21_X1 U21180 ( .B1(n18086), .B2(n18688), .A(n18085), .ZN(n18112) );
  AOI211_X1 U21181 ( .C1(n18088), .C2(n18120), .A(n18106), .B(n18112), .ZN(
        n18087) );
  NOR2_X1 U21182 ( .A1(n18087), .A2(n18185), .ZN(n18104) );
  AOI21_X1 U21183 ( .B1(n18104), .B2(n18088), .A(n18164), .ZN(n18103) );
  NAND2_X1 U21184 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18129) );
  INV_X1 U21185 ( .A(n18089), .ZN(n18154) );
  OAI22_X1 U21186 ( .A1(n18158), .A2(n18688), .B1(n18129), .B2(n18154), .ZN(
        n18141) );
  NAND2_X1 U21187 ( .A1(n18090), .A2(n18141), .ZN(n18113) );
  NOR2_X1 U21188 ( .A1(n18091), .A2(n18113), .ZN(n18092) );
  AOI22_X1 U21189 ( .A1(n18094), .A2(n18093), .B1(n18092), .B2(n18102), .ZN(
        n18096) );
  OAI22_X1 U21190 ( .A1(n18096), .A2(n18185), .B1(n18145), .B2(n18095), .ZN(
        n18097) );
  AOI21_X1 U21191 ( .B1(n18099), .B2(n18098), .A(n18097), .ZN(n18101) );
  OAI211_X1 U21192 ( .C1(n18103), .C2(n18102), .A(n18101), .B(n18100), .ZN(
        P3_U2854) );
  AOI21_X1 U21193 ( .B1(n18164), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18104), .ZN(n18105) );
  AOI221_X1 U21194 ( .B1(n18120), .B2(n18106), .C1(n18113), .C2(n18106), .A(
        n18105), .ZN(n18107) );
  AOI211_X1 U21195 ( .C1(n18109), .C2(n18182), .A(n18108), .B(n18107), .ZN(
        n18110) );
  OAI21_X1 U21196 ( .B1(n18177), .B2(n18111), .A(n18110), .ZN(P3_U2855) );
  OAI21_X1 U21197 ( .B1(n18185), .B2(n18112), .A(n18179), .ZN(n18122) );
  NOR2_X1 U21198 ( .A1(n18113), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18117) );
  OAI22_X1 U21199 ( .A1(n18145), .A2(n18115), .B1(n18177), .B2(n18114), .ZN(
        n18116) );
  AOI21_X1 U21200 ( .B1(n18117), .B2(n18163), .A(n18116), .ZN(n18119) );
  NAND2_X1 U21201 ( .A1(n9732), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18118) );
  OAI211_X1 U21202 ( .C1(n18120), .C2(n18122), .A(n18119), .B(n18118), .ZN(
        P3_U2856) );
  NAND3_X1 U21203 ( .A1(n18163), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18141), .ZN(n18140) );
  NOR2_X1 U21204 ( .A1(n18140), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18124) );
  OAI22_X1 U21205 ( .A1(n21107), .A2(n18122), .B1(n18177), .B2(n18121), .ZN(
        n18123) );
  AOI21_X1 U21206 ( .B1(n18124), .B2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n18123), .ZN(n18126) );
  OAI211_X1 U21207 ( .C1(n18145), .C2(n18127), .A(n18126), .B(n18125), .ZN(
        P3_U2857) );
  AOI22_X1 U21208 ( .A1(n18658), .A2(n18158), .B1(n18129), .B2(n18128), .ZN(
        n18131) );
  INV_X1 U21209 ( .A(n18157), .ZN(n18130) );
  NAND3_X1 U21210 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18131), .A3(
        n18130), .ZN(n18147) );
  AOI21_X1 U21211 ( .B1(n18132), .B2(n18147), .A(n18164), .ZN(n18138) );
  INV_X1 U21212 ( .A(n18133), .ZN(n18136) );
  OAI22_X1 U21213 ( .A1(n18179), .A2(n18744), .B1(n18177), .B2(n18134), .ZN(
        n18135) );
  AOI21_X1 U21214 ( .B1(n18182), .B2(n18136), .A(n18135), .ZN(n18137) );
  OAI221_X1 U21215 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18140), .C1(
        n18139), .C2(n18138), .A(n18137), .ZN(P3_U2858) );
  INV_X1 U21216 ( .A(n18141), .ZN(n18142) );
  AOI21_X1 U21217 ( .B1(n18142), .B2(n18151), .A(n18185), .ZN(n18148) );
  OAI22_X1 U21218 ( .A1(n18145), .A2(n18144), .B1(n18177), .B2(n18143), .ZN(
        n18146) );
  AOI21_X1 U21219 ( .B1(n18148), .B2(n18147), .A(n18146), .ZN(n18150) );
  OAI211_X1 U21220 ( .C1(n18169), .C2(n18151), .A(n18150), .B(n18149), .ZN(
        P3_U2859) );
  NAND2_X1 U21221 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18152) );
  OAI22_X1 U21222 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18153), .B1(
        n18688), .B2(n18152), .ZN(n18156) );
  INV_X1 U21223 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18821) );
  NOR3_X1 U21224 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18821), .A3(
        n18154), .ZN(n18155) );
  AOI221_X1 U21225 ( .B1(n18157), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18156), .C2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n18155), .ZN(
        n18160) );
  NAND2_X1 U21226 ( .A1(n18658), .A2(n18158), .ZN(n18159) );
  OAI211_X1 U21227 ( .C1(n18161), .C2(n9765), .A(n18160), .B(n18159), .ZN(
        n18162) );
  AOI22_X1 U21228 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18164), .B1(
        n18163), .B2(n18162), .ZN(n18166) );
  OAI211_X1 U21229 ( .C1(n18167), .C2(n18177), .A(n18166), .B(n18165), .ZN(
        P3_U2860) );
  OR3_X1 U21230 ( .A1(n18185), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18168), .ZN(n18187) );
  AOI21_X1 U21231 ( .B1(n18169), .B2(n18187), .A(n18821), .ZN(n18173) );
  AOI211_X1 U21232 ( .C1(n18171), .C2(n18838), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18170), .ZN(n18172) );
  AOI211_X1 U21233 ( .C1(n18182), .C2(n18174), .A(n18173), .B(n18172), .ZN(
        n18176) );
  NAND2_X1 U21234 ( .A1(n9732), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18175) );
  OAI211_X1 U21235 ( .C1(n18178), .C2(n18177), .A(n18176), .B(n18175), .ZN(
        P3_U2861) );
  INV_X1 U21236 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18848) );
  NOR2_X1 U21237 ( .A1(n18179), .A2(n18848), .ZN(n18180) );
  AOI221_X1 U21238 ( .B1(n18184), .B2(n18183), .C1(n18182), .C2(n18181), .A(
        n18180), .ZN(n18188) );
  OAI211_X1 U21239 ( .C1(n18673), .C2(n18185), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18179), .ZN(n18186) );
  NAND3_X1 U21240 ( .A1(n18188), .A2(n18187), .A3(n18186), .ZN(P3_U2862) );
  AOI21_X1 U21241 ( .B1(n18191), .B2(n18190), .A(n18189), .ZN(n18708) );
  NOR2_X1 U21242 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18810), .ZN(
        n18473) );
  OAI21_X1 U21243 ( .B1(n18708), .B2(n18473), .A(n18196), .ZN(n18192) );
  OAI221_X1 U21244 ( .B1(n18674), .B2(n18861), .C1(n18674), .C2(n18196), .A(
        n18192), .ZN(P3_U2863) );
  NOR2_X1 U21245 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18696), .ZN(
        n18495) );
  NOR2_X1 U21246 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18197), .ZN(
        n18380) );
  NOR2_X1 U21247 ( .A1(n18495), .A2(n18380), .ZN(n18194) );
  OAI22_X1 U21248 ( .A1(n18195), .A2(n18696), .B1(n18194), .B2(n18193), .ZN(
        P3_U2866) );
  NOR2_X1 U21249 ( .A1(n20840), .A2(n18196), .ZN(P3_U2867) );
  NOR2_X1 U21250 ( .A1(n18197), .A2(n18696), .ZN(n18523) );
  INV_X1 U21251 ( .A(n18523), .ZN(n18521) );
  NOR2_X1 U21252 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18675), .ZN(
        n18445) );
  NOR2_X1 U21253 ( .A1(n18674), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18425) );
  NOR2_X1 U21254 ( .A1(n18445), .A2(n18425), .ZN(n18498) );
  OR2_X1 U21255 ( .A1(n18521), .A2(n18498), .ZN(n18550) );
  NOR2_X1 U21256 ( .A1(n18696), .A2(n18378), .ZN(n18590) );
  NAND2_X1 U21257 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18590), .ZN(
        n18289) );
  INV_X1 U21258 ( .A(n18289), .ZN(n18638) );
  NOR2_X1 U21259 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18678) );
  NOR2_X1 U21260 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18291) );
  NAND2_X1 U21261 ( .A1(n18678), .A2(n18291), .ZN(n18306) );
  INV_X1 U21262 ( .A(n18306), .ZN(n18309) );
  NOR2_X1 U21263 ( .A1(n18638), .A2(n18309), .ZN(n18264) );
  AOI211_X1 U21264 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18472), .B(n18264), .ZN(
        n18198) );
  INV_X1 U21265 ( .A(n18198), .ZN(n18199) );
  OAI21_X1 U21266 ( .B1(n18550), .B2(n18356), .A(n18199), .ZN(n18244) );
  NAND2_X1 U21267 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18241), .ZN(n18595) );
  INV_X1 U21268 ( .A(n18595), .ZN(n18549) );
  NAND2_X1 U21269 ( .A1(n18425), .A2(n18523), .ZN(n18632) );
  INV_X1 U21270 ( .A(n18632), .ZN(n18636) );
  NOR2_X2 U21271 ( .A1(n18472), .A2(n18200), .ZN(n18587) );
  NOR2_X1 U21272 ( .A1(n18548), .A2(n18264), .ZN(n18238) );
  AOI22_X1 U21273 ( .A1(n18549), .A2(n18636), .B1(n18587), .B2(n18238), .ZN(
        n18207) );
  INV_X1 U21274 ( .A(n18201), .ZN(n18202) );
  NAND2_X1 U21275 ( .A1(n18203), .A2(n18202), .ZN(n18239) );
  NOR2_X2 U21276 ( .A1(n18204), .A2(n18239), .ZN(n18592) );
  NAND2_X1 U21277 ( .A1(n18241), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18557) );
  INV_X1 U21278 ( .A(n18557), .ZN(n18588) );
  INV_X1 U21279 ( .A(n18445), .ZN(n18205) );
  AOI22_X1 U21280 ( .A1(n18592), .A2(n18309), .B1(n18588), .B2(n9716), .ZN(
        n18206) );
  OAI211_X1 U21281 ( .C1(n18208), .C2(n18244), .A(n18207), .B(n18206), .ZN(
        P3_U2868) );
  NAND2_X1 U21282 ( .A1(n18241), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18601) );
  INV_X1 U21283 ( .A(n18601), .ZN(n18527) );
  NOR2_X2 U21284 ( .A1(n18472), .A2(n18209), .ZN(n18597) );
  AOI22_X1 U21285 ( .A1(n18527), .A2(n9716), .B1(n18597), .B2(n18238), .ZN(
        n18212) );
  NOR2_X2 U21286 ( .A1(n18210), .A2(n18239), .ZN(n18598) );
  NAND2_X1 U21287 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18241), .ZN(n18530) );
  INV_X1 U21288 ( .A(n18530), .ZN(n18596) );
  AOI22_X1 U21289 ( .A1(n18598), .A2(n18309), .B1(n18596), .B2(n18636), .ZN(
        n18211) );
  OAI211_X1 U21290 ( .C1(n20831), .C2(n18244), .A(n18212), .B(n18211), .ZN(
        P3_U2869) );
  NAND2_X1 U21291 ( .A1(n18241), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18607) );
  INV_X1 U21292 ( .A(n18607), .ZN(n18560) );
  NOR2_X2 U21293 ( .A1(n18472), .A2(n18213), .ZN(n18603) );
  AOI22_X1 U21294 ( .A1(n18560), .A2(n9716), .B1(n18603), .B2(n18238), .ZN(
        n18216) );
  NOR2_X2 U21295 ( .A1(n18214), .A2(n18239), .ZN(n18604) );
  NAND2_X1 U21296 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18241), .ZN(n18563) );
  INV_X1 U21297 ( .A(n18563), .ZN(n18602) );
  AOI22_X1 U21298 ( .A1(n18604), .A2(n18309), .B1(n18602), .B2(n18636), .ZN(
        n18215) );
  OAI211_X1 U21299 ( .C1(n18217), .C2(n18244), .A(n18216), .B(n18215), .ZN(
        P3_U2870) );
  NOR2_X2 U21300 ( .A1(n18472), .A2(n18218), .ZN(n18609) );
  NAND2_X1 U21301 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18241), .ZN(n18567) );
  INV_X1 U21302 ( .A(n18567), .ZN(n18608) );
  AOI22_X1 U21303 ( .A1(n18609), .A2(n18238), .B1(n18608), .B2(n18636), .ZN(
        n18221) );
  NAND2_X1 U21304 ( .A1(n18241), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18613) );
  INV_X1 U21305 ( .A(n18613), .ZN(n18564) );
  NOR2_X2 U21306 ( .A1(n18219), .A2(n18239), .ZN(n18610) );
  AOI22_X1 U21307 ( .A1(n18564), .A2(n9716), .B1(n18610), .B2(n18309), .ZN(
        n18220) );
  OAI211_X1 U21308 ( .C1(n18222), .C2(n18244), .A(n18221), .B(n18220), .ZN(
        P3_U2871) );
  NOR2_X1 U21309 ( .A1(n19222), .A2(n18356), .ZN(n18615) );
  NOR2_X2 U21310 ( .A1(n18472), .A2(n18223), .ZN(n18614) );
  AOI22_X1 U21311 ( .A1(n18615), .A2(n18636), .B1(n18614), .B2(n18238), .ZN(
        n18226) );
  NAND2_X1 U21312 ( .A1(n18241), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18619) );
  INV_X1 U21313 ( .A(n18619), .ZN(n18568) );
  NOR2_X2 U21314 ( .A1(n18224), .A2(n18239), .ZN(n18616) );
  AOI22_X1 U21315 ( .A1(n18568), .A2(n9716), .B1(n18616), .B2(n18309), .ZN(
        n18225) );
  OAI211_X1 U21316 ( .C1(n20874), .C2(n18244), .A(n18226), .B(n18225), .ZN(
        P3_U2872) );
  NAND2_X1 U21317 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18241), .ZN(n18625) );
  INV_X1 U21318 ( .A(n18625), .ZN(n18573) );
  NOR2_X2 U21319 ( .A1(n18472), .A2(n20847), .ZN(n18620) );
  AOI22_X1 U21320 ( .A1(n18573), .A2(n18636), .B1(n18620), .B2(n18238), .ZN(
        n18229) );
  NOR2_X2 U21321 ( .A1(n18227), .A2(n18239), .ZN(n18622) );
  NAND2_X1 U21322 ( .A1(n18241), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18576) );
  INV_X1 U21323 ( .A(n18576), .ZN(n18621) );
  AOI22_X1 U21324 ( .A1(n18622), .A2(n18309), .B1(n18621), .B2(n9716), .ZN(
        n18228) );
  OAI211_X1 U21325 ( .C1(n18230), .C2(n18244), .A(n18229), .B(n18228), .ZN(
        P3_U2873) );
  NAND2_X1 U21326 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18241), .ZN(n18580) );
  INV_X1 U21327 ( .A(n18580), .ZN(n18628) );
  NOR2_X2 U21328 ( .A1(n18472), .A2(n18231), .ZN(n18626) );
  AOI22_X1 U21329 ( .A1(n18628), .A2(n18636), .B1(n18626), .B2(n18238), .ZN(
        n18235) );
  NOR2_X2 U21330 ( .A1(n18232), .A2(n18239), .ZN(n18629) );
  NOR2_X1 U21331 ( .A1(n18356), .A2(n18233), .ZN(n18577) );
  AOI22_X1 U21332 ( .A1(n18629), .A2(n18309), .B1(n18577), .B2(n9716), .ZN(
        n18234) );
  OAI211_X1 U21333 ( .C1(n18236), .C2(n18244), .A(n18235), .B(n18234), .ZN(
        P3_U2874) );
  NOR2_X1 U21334 ( .A1(n18356), .A2(n19237), .ZN(n18542) );
  NOR2_X2 U21335 ( .A1(n18472), .A2(n18237), .ZN(n18635) );
  AOI22_X1 U21336 ( .A1(n18542), .A2(n18636), .B1(n18635), .B2(n18238), .ZN(
        n18243) );
  NOR2_X2 U21337 ( .A1(n18240), .A2(n18239), .ZN(n18639) );
  NAND2_X1 U21338 ( .A1(n18241), .A2(BUF2_REG_23__SCAN_IN), .ZN(n18547) );
  INV_X1 U21339 ( .A(n18547), .ZN(n18637) );
  AOI22_X1 U21340 ( .A1(n18639), .A2(n18309), .B1(n18637), .B2(n9716), .ZN(
        n18242) );
  OAI211_X1 U21341 ( .C1(n21001), .C2(n18244), .A(n18243), .B(n18242), .ZN(
        P3_U2875) );
  INV_X1 U21342 ( .A(n18291), .ZN(n18290) );
  INV_X1 U21343 ( .A(n18548), .ZN(n18716) );
  NAND2_X1 U21344 ( .A1(n18675), .A2(n18716), .ZN(n18520) );
  NOR2_X1 U21345 ( .A1(n18290), .A2(n18520), .ZN(n18260) );
  AOI22_X1 U21346 ( .A1(n18549), .A2(n9716), .B1(n18587), .B2(n18260), .ZN(
        n18246) );
  NOR3_X1 U21347 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18473), .A3(
        n18472), .ZN(n18522) );
  AOI22_X1 U21348 ( .A1(n18241), .A2(n18590), .B1(n18291), .B2(n18522), .ZN(
        n18261) );
  NAND2_X1 U21349 ( .A1(n18425), .A2(n18291), .ZN(n18333) );
  INV_X1 U21350 ( .A(n18333), .ZN(n18324) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18261), .B1(
        n18592), .B2(n18324), .ZN(n18245) );
  OAI211_X1 U21352 ( .C1(n18557), .C2(n18289), .A(n18246), .B(n18245), .ZN(
        P3_U2876) );
  AOI22_X1 U21353 ( .A1(n18597), .A2(n18260), .B1(n18596), .B2(n9716), .ZN(
        n18248) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18261), .B1(
        n18598), .B2(n18324), .ZN(n18247) );
  OAI211_X1 U21355 ( .C1(n18601), .C2(n18289), .A(n18248), .B(n18247), .ZN(
        P3_U2877) );
  INV_X1 U21356 ( .A(n9716), .ZN(n18259) );
  AOI22_X1 U21357 ( .A1(n18560), .A2(n18638), .B1(n18603), .B2(n18260), .ZN(
        n18250) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18261), .B1(
        n18604), .B2(n18324), .ZN(n18249) );
  OAI211_X1 U21359 ( .C1(n18563), .C2(n18259), .A(n18250), .B(n18249), .ZN(
        P3_U2878) );
  AOI22_X1 U21360 ( .A1(n18609), .A2(n18260), .B1(n18608), .B2(n9716), .ZN(
        n18252) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18261), .B1(
        n18610), .B2(n18324), .ZN(n18251) );
  OAI211_X1 U21362 ( .C1(n18613), .C2(n18289), .A(n18252), .B(n18251), .ZN(
        P3_U2879) );
  INV_X1 U21363 ( .A(n18615), .ZN(n18571) );
  AOI22_X1 U21364 ( .A1(n18568), .A2(n18638), .B1(n18614), .B2(n18260), .ZN(
        n18254) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18261), .B1(
        n18616), .B2(n18324), .ZN(n18253) );
  OAI211_X1 U21366 ( .C1(n18571), .C2(n18259), .A(n18254), .B(n18253), .ZN(
        P3_U2880) );
  AOI22_X1 U21367 ( .A1(n18621), .A2(n18638), .B1(n18620), .B2(n18260), .ZN(
        n18256) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18261), .B1(
        n18622), .B2(n18324), .ZN(n18255) );
  OAI211_X1 U21369 ( .C1(n18625), .C2(n18259), .A(n18256), .B(n18255), .ZN(
        P3_U2881) );
  AOI22_X1 U21370 ( .A1(n18577), .A2(n18638), .B1(n18626), .B2(n18260), .ZN(
        n18258) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18261), .B1(
        n18629), .B2(n18324), .ZN(n18257) );
  OAI211_X1 U21372 ( .C1(n18580), .C2(n18259), .A(n18258), .B(n18257), .ZN(
        P3_U2882) );
  AOI22_X1 U21373 ( .A1(n18542), .A2(n9716), .B1(n18635), .B2(n18260), .ZN(
        n18263) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18261), .B1(
        n18639), .B2(n18324), .ZN(n18262) );
  OAI211_X1 U21375 ( .C1(n18547), .C2(n18289), .A(n18263), .B(n18262), .ZN(
        P3_U2883) );
  NAND2_X1 U21376 ( .A1(n18445), .A2(n18291), .ZN(n18355) );
  INV_X1 U21377 ( .A(n18496), .ZN(n18551) );
  NOR2_X1 U21378 ( .A1(n18324), .A2(n18348), .ZN(n18312) );
  OAI21_X1 U21379 ( .B1(n18551), .B2(n18264), .A(n18312), .ZN(n18265) );
  OAI211_X1 U21380 ( .C1(n18810), .C2(n18348), .A(n18265), .B(n18554), .ZN(
        n18286) );
  INV_X1 U21381 ( .A(n18286), .ZN(n18282) );
  NOR2_X1 U21382 ( .A1(n18548), .A2(n18312), .ZN(n18285) );
  AOI22_X1 U21383 ( .A1(n18549), .A2(n18638), .B1(n18587), .B2(n18285), .ZN(
        n18267) );
  AOI22_X1 U21384 ( .A1(n18592), .A2(n18348), .B1(n18588), .B2(n18309), .ZN(
        n18266) );
  OAI211_X1 U21385 ( .C1(n18282), .C2(n18268), .A(n18267), .B(n18266), .ZN(
        P3_U2884) );
  INV_X1 U21386 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18271) );
  AOI22_X1 U21387 ( .A1(n18527), .A2(n18309), .B1(n18597), .B2(n18285), .ZN(
        n18270) );
  AOI22_X1 U21388 ( .A1(n18598), .A2(n18348), .B1(n18596), .B2(n18638), .ZN(
        n18269) );
  OAI211_X1 U21389 ( .C1(n18282), .C2(n18271), .A(n18270), .B(n18269), .ZN(
        P3_U2885) );
  AOI22_X1 U21390 ( .A1(n18603), .A2(n18285), .B1(n18602), .B2(n18638), .ZN(
        n18273) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18286), .B1(
        n18604), .B2(n18348), .ZN(n18272) );
  OAI211_X1 U21392 ( .C1(n18607), .C2(n18306), .A(n18273), .B(n18272), .ZN(
        P3_U2886) );
  AOI22_X1 U21393 ( .A1(n18609), .A2(n18285), .B1(n18608), .B2(n18638), .ZN(
        n18275) );
  AOI22_X1 U21394 ( .A1(n18564), .A2(n18309), .B1(n18610), .B2(n18348), .ZN(
        n18274) );
  OAI211_X1 U21395 ( .C1(n18282), .C2(n18276), .A(n18275), .B(n18274), .ZN(
        P3_U2887) );
  AOI22_X1 U21396 ( .A1(n18568), .A2(n18309), .B1(n18614), .B2(n18285), .ZN(
        n18278) );
  AOI22_X1 U21397 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18286), .B1(
        n18616), .B2(n18348), .ZN(n18277) );
  OAI211_X1 U21398 ( .C1(n18571), .C2(n18289), .A(n18278), .B(n18277), .ZN(
        P3_U2888) );
  AOI22_X1 U21399 ( .A1(n18621), .A2(n18309), .B1(n18620), .B2(n18285), .ZN(
        n18280) );
  AOI22_X1 U21400 ( .A1(n18573), .A2(n18638), .B1(n18622), .B2(n18348), .ZN(
        n18279) );
  OAI211_X1 U21401 ( .C1(n18282), .C2(n18281), .A(n18280), .B(n18279), .ZN(
        P3_U2889) );
  INV_X1 U21402 ( .A(n18577), .ZN(n18633) );
  AOI22_X1 U21403 ( .A1(n18628), .A2(n18638), .B1(n18626), .B2(n18285), .ZN(
        n18284) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18286), .B1(
        n18629), .B2(n18348), .ZN(n18283) );
  OAI211_X1 U21405 ( .C1(n18633), .C2(n18306), .A(n18284), .B(n18283), .ZN(
        P3_U2890) );
  INV_X1 U21406 ( .A(n18542), .ZN(n18644) );
  AOI22_X1 U21407 ( .A1(n18637), .A2(n18309), .B1(n18635), .B2(n18285), .ZN(
        n18288) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18286), .B1(
        n18639), .B2(n18348), .ZN(n18287) );
  OAI211_X1 U21409 ( .C1(n18644), .C2(n18289), .A(n18288), .B(n18287), .ZN(
        P3_U2891) );
  NOR2_X1 U21410 ( .A1(n18675), .A2(n18290), .ZN(n18335) );
  AND2_X1 U21411 ( .A1(n18716), .A2(n18335), .ZN(n18307) );
  AOI22_X1 U21412 ( .A1(n18549), .A2(n18309), .B1(n18587), .B2(n18307), .ZN(
        n18293) );
  NAND2_X1 U21413 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18335), .ZN(
        n18377) );
  AOI21_X1 U21414 ( .B1(n18675), .B2(n18551), .A(n18472), .ZN(n18379) );
  OAI211_X1 U21415 ( .C1(n18370), .C2(n18810), .A(n18291), .B(n18379), .ZN(
        n18308) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18308), .B1(
        n18592), .B2(n18370), .ZN(n18292) );
  OAI211_X1 U21417 ( .C1(n18557), .C2(n18333), .A(n18293), .B(n18292), .ZN(
        P3_U2892) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18308), .B1(
        n18597), .B2(n18307), .ZN(n18295) );
  AOI22_X1 U21419 ( .A1(n18598), .A2(n18370), .B1(n18596), .B2(n18309), .ZN(
        n18294) );
  OAI211_X1 U21420 ( .C1(n18601), .C2(n18333), .A(n18295), .B(n18294), .ZN(
        P3_U2893) );
  AOI22_X1 U21421 ( .A1(n18560), .A2(n18324), .B1(n18603), .B2(n18307), .ZN(
        n18297) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18308), .B1(
        n18604), .B2(n18370), .ZN(n18296) );
  OAI211_X1 U21423 ( .C1(n18563), .C2(n18306), .A(n18297), .B(n18296), .ZN(
        P3_U2894) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18308), .B1(
        n18609), .B2(n18307), .ZN(n18299) );
  AOI22_X1 U21425 ( .A1(n18610), .A2(n18370), .B1(n18608), .B2(n18309), .ZN(
        n18298) );
  OAI211_X1 U21426 ( .C1(n18613), .C2(n18333), .A(n18299), .B(n18298), .ZN(
        P3_U2895) );
  AOI22_X1 U21427 ( .A1(n18568), .A2(n18324), .B1(n18614), .B2(n18307), .ZN(
        n18301) );
  AOI22_X1 U21428 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18308), .B1(
        n18616), .B2(n18370), .ZN(n18300) );
  OAI211_X1 U21429 ( .C1(n18571), .C2(n18306), .A(n18301), .B(n18300), .ZN(
        P3_U2896) );
  AOI22_X1 U21430 ( .A1(n18621), .A2(n18324), .B1(n18620), .B2(n18307), .ZN(
        n18303) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18308), .B1(
        n18622), .B2(n18370), .ZN(n18302) );
  OAI211_X1 U21432 ( .C1(n18625), .C2(n18306), .A(n18303), .B(n18302), .ZN(
        P3_U2897) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18308), .B1(
        n18626), .B2(n18307), .ZN(n18305) );
  AOI22_X1 U21434 ( .A1(n18629), .A2(n18370), .B1(n18577), .B2(n18324), .ZN(
        n18304) );
  OAI211_X1 U21435 ( .C1(n18580), .C2(n18306), .A(n18305), .B(n18304), .ZN(
        P3_U2898) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18308), .B1(
        n18635), .B2(n18307), .ZN(n18311) );
  AOI22_X1 U21437 ( .A1(n18542), .A2(n18309), .B1(n18639), .B2(n18370), .ZN(
        n18310) );
  OAI211_X1 U21438 ( .C1(n18547), .C2(n18333), .A(n18311), .B(n18310), .ZN(
        P3_U2899) );
  NAND2_X1 U21439 ( .A1(n18678), .A2(n18380), .ZN(n18400) );
  AOI21_X1 U21440 ( .B1(n18377), .B2(n18400), .A(n18548), .ZN(n18329) );
  AOI22_X1 U21441 ( .A1(n18549), .A2(n18324), .B1(n18587), .B2(n18329), .ZN(
        n18315) );
  INV_X1 U21442 ( .A(n18400), .ZN(n18383) );
  AOI221_X1 U21443 ( .B1(n18312), .B2(n18377), .C1(n18551), .C2(n18377), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18313) );
  OAI21_X1 U21444 ( .B1(n18383), .B2(n18313), .A(n18554), .ZN(n18330) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18330), .B1(
        n18592), .B2(n18383), .ZN(n18314) );
  OAI211_X1 U21446 ( .C1(n18557), .C2(n18355), .A(n18315), .B(n18314), .ZN(
        P3_U2900) );
  AOI22_X1 U21447 ( .A1(n18527), .A2(n18348), .B1(n18597), .B2(n18329), .ZN(
        n18317) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18330), .B1(
        n18598), .B2(n18383), .ZN(n18316) );
  OAI211_X1 U21449 ( .C1(n18530), .C2(n18333), .A(n18317), .B(n18316), .ZN(
        P3_U2901) );
  AOI22_X1 U21450 ( .A1(n18603), .A2(n18329), .B1(n18602), .B2(n18324), .ZN(
        n18319) );
  AOI22_X1 U21451 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18330), .B1(
        n18604), .B2(n18383), .ZN(n18318) );
  OAI211_X1 U21452 ( .C1(n18607), .C2(n18355), .A(n18319), .B(n18318), .ZN(
        P3_U2902) );
  AOI22_X1 U21453 ( .A1(n18609), .A2(n18329), .B1(n18608), .B2(n18324), .ZN(
        n18321) );
  AOI22_X1 U21454 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18330), .B1(
        n18610), .B2(n18383), .ZN(n18320) );
  OAI211_X1 U21455 ( .C1(n18613), .C2(n18355), .A(n18321), .B(n18320), .ZN(
        P3_U2903) );
  AOI22_X1 U21456 ( .A1(n18615), .A2(n18324), .B1(n18614), .B2(n18329), .ZN(
        n18323) );
  AOI22_X1 U21457 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18330), .B1(
        n18616), .B2(n18383), .ZN(n18322) );
  OAI211_X1 U21458 ( .C1(n18619), .C2(n18355), .A(n18323), .B(n18322), .ZN(
        P3_U2904) );
  AOI22_X1 U21459 ( .A1(n18573), .A2(n18324), .B1(n18620), .B2(n18329), .ZN(
        n18326) );
  AOI22_X1 U21460 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18330), .B1(
        n18622), .B2(n18383), .ZN(n18325) );
  OAI211_X1 U21461 ( .C1(n18576), .C2(n18355), .A(n18326), .B(n18325), .ZN(
        P3_U2905) );
  AOI22_X1 U21462 ( .A1(n18577), .A2(n18348), .B1(n18626), .B2(n18329), .ZN(
        n18328) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18330), .B1(
        n18629), .B2(n18383), .ZN(n18327) );
  OAI211_X1 U21464 ( .C1(n18580), .C2(n18333), .A(n18328), .B(n18327), .ZN(
        P3_U2906) );
  AOI22_X1 U21465 ( .A1(n18637), .A2(n18348), .B1(n18635), .B2(n18329), .ZN(
        n18332) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18330), .B1(
        n18639), .B2(n18383), .ZN(n18331) );
  OAI211_X1 U21467 ( .C1(n18644), .C2(n18333), .A(n18332), .B(n18331), .ZN(
        P3_U2907) );
  INV_X1 U21468 ( .A(n18380), .ZN(n18334) );
  NOR2_X1 U21469 ( .A1(n18334), .A2(n18520), .ZN(n18351) );
  AOI22_X1 U21470 ( .A1(n18549), .A2(n18348), .B1(n18587), .B2(n18351), .ZN(
        n18337) );
  AOI22_X1 U21471 ( .A1(n18241), .A2(n18335), .B1(n18380), .B2(n18522), .ZN(
        n18352) );
  NAND2_X1 U21472 ( .A1(n18380), .A2(n18425), .ZN(n18414) );
  INV_X1 U21473 ( .A(n18414), .ZN(n18420) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18352), .B1(
        n18592), .B2(n18420), .ZN(n18336) );
  OAI211_X1 U21475 ( .C1(n18557), .C2(n18377), .A(n18337), .B(n18336), .ZN(
        P3_U2908) );
  AOI22_X1 U21476 ( .A1(n18597), .A2(n18351), .B1(n18596), .B2(n18348), .ZN(
        n18339) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18352), .B1(
        n18598), .B2(n18420), .ZN(n18338) );
  OAI211_X1 U21478 ( .C1(n18601), .C2(n18377), .A(n18339), .B(n18338), .ZN(
        P3_U2909) );
  AOI22_X1 U21479 ( .A1(n18560), .A2(n18370), .B1(n18603), .B2(n18351), .ZN(
        n18341) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18352), .B1(
        n18604), .B2(n18420), .ZN(n18340) );
  OAI211_X1 U21481 ( .C1(n18563), .C2(n18355), .A(n18341), .B(n18340), .ZN(
        P3_U2910) );
  AOI22_X1 U21482 ( .A1(n18609), .A2(n18351), .B1(n18608), .B2(n18348), .ZN(
        n18343) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18352), .B1(
        n18610), .B2(n18420), .ZN(n18342) );
  OAI211_X1 U21484 ( .C1(n18613), .C2(n18377), .A(n18343), .B(n18342), .ZN(
        P3_U2911) );
  AOI22_X1 U21485 ( .A1(n18615), .A2(n18348), .B1(n18614), .B2(n18351), .ZN(
        n18345) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18352), .B1(
        n18616), .B2(n18420), .ZN(n18344) );
  OAI211_X1 U21487 ( .C1(n18619), .C2(n18377), .A(n18345), .B(n18344), .ZN(
        P3_U2912) );
  AOI22_X1 U21488 ( .A1(n18621), .A2(n18370), .B1(n18620), .B2(n18351), .ZN(
        n18347) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18352), .B1(
        n18622), .B2(n18420), .ZN(n18346) );
  OAI211_X1 U21490 ( .C1(n18625), .C2(n18355), .A(n18347), .B(n18346), .ZN(
        P3_U2913) );
  AOI22_X1 U21491 ( .A1(n18628), .A2(n18348), .B1(n18626), .B2(n18351), .ZN(
        n18350) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18352), .B1(
        n18629), .B2(n18420), .ZN(n18349) );
  OAI211_X1 U21493 ( .C1(n18633), .C2(n18377), .A(n18350), .B(n18349), .ZN(
        P3_U2914) );
  AOI22_X1 U21494 ( .A1(n18637), .A2(n18370), .B1(n18635), .B2(n18351), .ZN(
        n18354) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18352), .B1(
        n18639), .B2(n18420), .ZN(n18353) );
  OAI211_X1 U21496 ( .C1(n18644), .C2(n18355), .A(n18354), .B(n18353), .ZN(
        P3_U2915) );
  NAND2_X1 U21497 ( .A1(n18380), .A2(n18445), .ZN(n18438) );
  AOI21_X1 U21498 ( .B1(n18414), .B2(n18438), .A(n18548), .ZN(n18373) );
  AOI22_X1 U21499 ( .A1(n18549), .A2(n18370), .B1(n18587), .B2(n18373), .ZN(
        n18359) );
  INV_X1 U21500 ( .A(n18438), .ZN(n18441) );
  AOI21_X1 U21501 ( .B1(n18414), .B2(n18438), .A(n18472), .ZN(n18401) );
  AOI21_X1 U21502 ( .B1(n18377), .B2(n18400), .A(n18356), .ZN(n18357) );
  OAI22_X1 U21503 ( .A1(n18441), .A2(n18810), .B1(n18401), .B2(n18357), .ZN(
        n18374) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18374), .B1(
        n18592), .B2(n18441), .ZN(n18358) );
  OAI211_X1 U21505 ( .C1(n18557), .C2(n18400), .A(n18359), .B(n18358), .ZN(
        P3_U2916) );
  AOI22_X1 U21506 ( .A1(n18597), .A2(n18373), .B1(n18596), .B2(n18370), .ZN(
        n18361) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18374), .B1(
        n18598), .B2(n18441), .ZN(n18360) );
  OAI211_X1 U21508 ( .C1(n18601), .C2(n18400), .A(n18361), .B(n18360), .ZN(
        P3_U2917) );
  AOI22_X1 U21509 ( .A1(n18603), .A2(n18373), .B1(n18602), .B2(n18370), .ZN(
        n18363) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18374), .B1(
        n18604), .B2(n18441), .ZN(n18362) );
  OAI211_X1 U21511 ( .C1(n18607), .C2(n18400), .A(n18363), .B(n18362), .ZN(
        P3_U2918) );
  AOI22_X1 U21512 ( .A1(n18564), .A2(n18383), .B1(n18609), .B2(n18373), .ZN(
        n18365) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18374), .B1(
        n18610), .B2(n18441), .ZN(n18364) );
  OAI211_X1 U21514 ( .C1(n18567), .C2(n18377), .A(n18365), .B(n18364), .ZN(
        P3_U2919) );
  AOI22_X1 U21515 ( .A1(n18615), .A2(n18370), .B1(n18614), .B2(n18373), .ZN(
        n18367) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18374), .B1(
        n18616), .B2(n18441), .ZN(n18366) );
  OAI211_X1 U21517 ( .C1(n18619), .C2(n18400), .A(n18367), .B(n18366), .ZN(
        P3_U2920) );
  AOI22_X1 U21518 ( .A1(n18573), .A2(n18370), .B1(n18620), .B2(n18373), .ZN(
        n18369) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18374), .B1(
        n18622), .B2(n18441), .ZN(n18368) );
  OAI211_X1 U21520 ( .C1(n18576), .C2(n18400), .A(n18369), .B(n18368), .ZN(
        P3_U2921) );
  AOI22_X1 U21521 ( .A1(n18628), .A2(n18370), .B1(n18626), .B2(n18373), .ZN(
        n18372) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18374), .B1(
        n18629), .B2(n18441), .ZN(n18371) );
  OAI211_X1 U21523 ( .C1(n18633), .C2(n18400), .A(n18372), .B(n18371), .ZN(
        P3_U2922) );
  AOI22_X1 U21524 ( .A1(n18637), .A2(n18383), .B1(n18635), .B2(n18373), .ZN(
        n18376) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18374), .B1(
        n18639), .B2(n18441), .ZN(n18375) );
  OAI211_X1 U21526 ( .C1(n18644), .C2(n18377), .A(n18376), .B(n18375), .ZN(
        P3_U2923) );
  NOR2_X1 U21527 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18378), .ZN(
        n18424) );
  AND2_X1 U21528 ( .A1(n18716), .A2(n18424), .ZN(n18396) );
  AOI22_X1 U21529 ( .A1(n18588), .A2(n18420), .B1(n18587), .B2(n18396), .ZN(
        n18382) );
  NAND2_X1 U21530 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18424), .ZN(
        n18464) );
  INV_X1 U21531 ( .A(n18464), .ZN(n18466) );
  OAI211_X1 U21532 ( .C1(n18466), .C2(n18810), .A(n18380), .B(n18379), .ZN(
        n18397) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18397), .B1(
        n18466), .B2(n18592), .ZN(n18381) );
  OAI211_X1 U21534 ( .C1(n18595), .C2(n18400), .A(n18382), .B(n18381), .ZN(
        P3_U2924) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18397), .B1(
        n18597), .B2(n18396), .ZN(n18385) );
  AOI22_X1 U21536 ( .A1(n18466), .A2(n18598), .B1(n18596), .B2(n18383), .ZN(
        n18384) );
  OAI211_X1 U21537 ( .C1(n18601), .C2(n18414), .A(n18385), .B(n18384), .ZN(
        P3_U2925) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18397), .B1(
        n18603), .B2(n18396), .ZN(n18387) );
  AOI22_X1 U21539 ( .A1(n18466), .A2(n18604), .B1(n18560), .B2(n18420), .ZN(
        n18386) );
  OAI211_X1 U21540 ( .C1(n18563), .C2(n18400), .A(n18387), .B(n18386), .ZN(
        P3_U2926) );
  AOI22_X1 U21541 ( .A1(n18564), .A2(n18420), .B1(n18609), .B2(n18396), .ZN(
        n18389) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18397), .B1(
        n18466), .B2(n18610), .ZN(n18388) );
  OAI211_X1 U21543 ( .C1(n18567), .C2(n18400), .A(n18389), .B(n18388), .ZN(
        P3_U2927) );
  AOI22_X1 U21544 ( .A1(n18568), .A2(n18420), .B1(n18614), .B2(n18396), .ZN(
        n18391) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18397), .B1(
        n18466), .B2(n18616), .ZN(n18390) );
  OAI211_X1 U21546 ( .C1(n18571), .C2(n18400), .A(n18391), .B(n18390), .ZN(
        P3_U2928) );
  AOI22_X1 U21547 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18397), .B1(
        n18620), .B2(n18396), .ZN(n18393) );
  AOI22_X1 U21548 ( .A1(n18466), .A2(n18622), .B1(n18621), .B2(n18420), .ZN(
        n18392) );
  OAI211_X1 U21549 ( .C1(n18625), .C2(n18400), .A(n18393), .B(n18392), .ZN(
        P3_U2929) );
  AOI22_X1 U21550 ( .A1(n18577), .A2(n18420), .B1(n18626), .B2(n18396), .ZN(
        n18395) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18397), .B1(
        n18466), .B2(n18629), .ZN(n18394) );
  OAI211_X1 U21552 ( .C1(n18580), .C2(n18400), .A(n18395), .B(n18394), .ZN(
        P3_U2930) );
  AOI22_X1 U21553 ( .A1(n18637), .A2(n18420), .B1(n18635), .B2(n18396), .ZN(
        n18399) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18397), .B1(
        n18466), .B2(n18639), .ZN(n18398) );
  OAI211_X1 U21555 ( .C1(n18644), .C2(n18400), .A(n18399), .B(n18398), .ZN(
        P3_U2931) );
  NAND2_X1 U21556 ( .A1(n18678), .A2(n18495), .ZN(n18481) );
  NAND2_X1 U21557 ( .A1(n18464), .A2(n18481), .ZN(n18446) );
  AOI22_X1 U21558 ( .A1(n18554), .A2(n18446), .B1(n18496), .B2(n18401), .ZN(
        n18402) );
  AOI21_X1 U21559 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18481), .A(n18402), 
        .ZN(n18405) );
  AND2_X1 U21560 ( .A1(n18716), .A2(n18446), .ZN(n18419) );
  AOI22_X1 U21561 ( .A1(n18549), .A2(n18420), .B1(n18587), .B2(n18419), .ZN(
        n18404) );
  INV_X1 U21562 ( .A(n18481), .ZN(n18491) );
  AOI22_X1 U21563 ( .A1(n18491), .A2(n18592), .B1(n18588), .B2(n18441), .ZN(
        n18403) );
  OAI211_X1 U21564 ( .C1(n18405), .C2(n20856), .A(n18404), .B(n18403), .ZN(
        P3_U2932) );
  AOI22_X1 U21565 ( .A1(n18597), .A2(n18419), .B1(n18596), .B2(n18420), .ZN(
        n18407) );
  INV_X1 U21566 ( .A(n18405), .ZN(n18421) );
  AOI22_X1 U21567 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18421), .B1(
        n18491), .B2(n18598), .ZN(n18406) );
  OAI211_X1 U21568 ( .C1(n18601), .C2(n18438), .A(n18407), .B(n18406), .ZN(
        P3_U2933) );
  AOI22_X1 U21569 ( .A1(n18560), .A2(n18441), .B1(n18603), .B2(n18419), .ZN(
        n18409) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18421), .B1(
        n18491), .B2(n18604), .ZN(n18408) );
  OAI211_X1 U21571 ( .C1(n18563), .C2(n18414), .A(n18409), .B(n18408), .ZN(
        P3_U2934) );
  AOI22_X1 U21572 ( .A1(n18564), .A2(n18441), .B1(n18609), .B2(n18419), .ZN(
        n18411) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18421), .B1(
        n18491), .B2(n18610), .ZN(n18410) );
  OAI211_X1 U21574 ( .C1(n18567), .C2(n18414), .A(n18411), .B(n18410), .ZN(
        P3_U2935) );
  AOI22_X1 U21575 ( .A1(n18568), .A2(n18441), .B1(n18614), .B2(n18419), .ZN(
        n18413) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18421), .B1(
        n18491), .B2(n18616), .ZN(n18412) );
  OAI211_X1 U21577 ( .C1(n18571), .C2(n18414), .A(n18413), .B(n18412), .ZN(
        P3_U2936) );
  AOI22_X1 U21578 ( .A1(n18573), .A2(n18420), .B1(n18620), .B2(n18419), .ZN(
        n18416) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18421), .B1(
        n18491), .B2(n18622), .ZN(n18415) );
  OAI211_X1 U21580 ( .C1(n18576), .C2(n18438), .A(n18416), .B(n18415), .ZN(
        P3_U2937) );
  AOI22_X1 U21581 ( .A1(n18628), .A2(n18420), .B1(n18626), .B2(n18419), .ZN(
        n18418) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18421), .B1(
        n18491), .B2(n18629), .ZN(n18417) );
  OAI211_X1 U21583 ( .C1(n18633), .C2(n18438), .A(n18418), .B(n18417), .ZN(
        P3_U2938) );
  AOI22_X1 U21584 ( .A1(n18542), .A2(n18420), .B1(n18635), .B2(n18419), .ZN(
        n18423) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18421), .B1(
        n18491), .B2(n18639), .ZN(n18422) );
  OAI211_X1 U21586 ( .C1(n18547), .C2(n18438), .A(n18423), .B(n18422), .ZN(
        P3_U2939) );
  INV_X1 U21587 ( .A(n18495), .ZN(n18471) );
  NOR2_X1 U21588 ( .A1(n18471), .A2(n18520), .ZN(n18474) );
  AOI22_X1 U21589 ( .A1(n18466), .A2(n18588), .B1(n18587), .B2(n18474), .ZN(
        n18427) );
  AOI22_X1 U21590 ( .A1(n18241), .A2(n18424), .B1(n18495), .B2(n18522), .ZN(
        n18442) );
  NAND2_X1 U21591 ( .A1(n18495), .A2(n18425), .ZN(n18502) );
  INV_X1 U21592 ( .A(n18502), .ZN(n18516) );
  AOI22_X1 U21593 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18442), .B1(
        n18516), .B2(n18592), .ZN(n18426) );
  OAI211_X1 U21594 ( .C1(n18595), .C2(n18438), .A(n18427), .B(n18426), .ZN(
        P3_U2940) );
  AOI22_X1 U21595 ( .A1(n18597), .A2(n18474), .B1(n18596), .B2(n18441), .ZN(
        n18429) );
  AOI22_X1 U21596 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18442), .B1(
        n18516), .B2(n18598), .ZN(n18428) );
  OAI211_X1 U21597 ( .C1(n18464), .C2(n18601), .A(n18429), .B(n18428), .ZN(
        P3_U2941) );
  AOI22_X1 U21598 ( .A1(n18603), .A2(n18474), .B1(n18602), .B2(n18441), .ZN(
        n18431) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18442), .B1(
        n18516), .B2(n18604), .ZN(n18430) );
  OAI211_X1 U21600 ( .C1(n18464), .C2(n18607), .A(n18431), .B(n18430), .ZN(
        P3_U2942) );
  AOI22_X1 U21601 ( .A1(n18466), .A2(n18564), .B1(n18609), .B2(n18474), .ZN(
        n18433) );
  AOI22_X1 U21602 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18442), .B1(
        n18516), .B2(n18610), .ZN(n18432) );
  OAI211_X1 U21603 ( .C1(n18567), .C2(n18438), .A(n18433), .B(n18432), .ZN(
        P3_U2943) );
  AOI22_X1 U21604 ( .A1(n18466), .A2(n18568), .B1(n18614), .B2(n18474), .ZN(
        n18435) );
  AOI22_X1 U21605 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18442), .B1(
        n18516), .B2(n18616), .ZN(n18434) );
  OAI211_X1 U21606 ( .C1(n18571), .C2(n18438), .A(n18435), .B(n18434), .ZN(
        P3_U2944) );
  AOI22_X1 U21607 ( .A1(n18466), .A2(n18621), .B1(n18620), .B2(n18474), .ZN(
        n18437) );
  AOI22_X1 U21608 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18442), .B1(
        n18516), .B2(n18622), .ZN(n18436) );
  OAI211_X1 U21609 ( .C1(n18625), .C2(n18438), .A(n18437), .B(n18436), .ZN(
        P3_U2945) );
  AOI22_X1 U21610 ( .A1(n18628), .A2(n18441), .B1(n18626), .B2(n18474), .ZN(
        n18440) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18442), .B1(
        n18516), .B2(n18629), .ZN(n18439) );
  OAI211_X1 U21612 ( .C1(n18464), .C2(n18633), .A(n18440), .B(n18439), .ZN(
        P3_U2946) );
  AOI22_X1 U21613 ( .A1(n18542), .A2(n18441), .B1(n18635), .B2(n18474), .ZN(
        n18444) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18442), .B1(
        n18516), .B2(n18639), .ZN(n18443) );
  OAI211_X1 U21615 ( .C1(n18464), .C2(n18547), .A(n18444), .B(n18443), .ZN(
        P3_U2947) );
  NAND2_X1 U21616 ( .A1(n18495), .A2(n18445), .ZN(n18541) );
  OAI221_X1 U21617 ( .B1(n18516), .B2(n18496), .C1(n18516), .C2(n18446), .A(
        n18810), .ZN(n18447) );
  AOI21_X1 U21618 ( .B1(n18541), .B2(n18447), .A(n18472), .ZN(n18470) );
  AOI22_X1 U21619 ( .A1(n18491), .A2(n18588), .B1(n18587), .B2(n18465), .ZN(
        n18449) );
  INV_X1 U21620 ( .A(n18541), .ZN(n18543) );
  AOI22_X1 U21621 ( .A1(n18549), .A2(n18466), .B1(n18543), .B2(n18592), .ZN(
        n18448) );
  OAI211_X1 U21622 ( .C1(n18470), .C2(n18450), .A(n18449), .B(n18448), .ZN(
        P3_U2948) );
  AOI22_X1 U21623 ( .A1(n18466), .A2(n18596), .B1(n18465), .B2(n18597), .ZN(
        n18452) );
  AOI22_X1 U21624 ( .A1(n18543), .A2(n18598), .B1(n18491), .B2(n18527), .ZN(
        n18451) );
  OAI211_X1 U21625 ( .C1(n18470), .C2(n20876), .A(n18452), .B(n18451), .ZN(
        P3_U2949) );
  AOI22_X1 U21626 ( .A1(n18466), .A2(n18602), .B1(n18465), .B2(n18603), .ZN(
        n18454) );
  INV_X1 U21627 ( .A(n18470), .ZN(n18461) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18461), .B1(
        n18543), .B2(n18604), .ZN(n18453) );
  OAI211_X1 U21629 ( .C1(n18481), .C2(n18607), .A(n18454), .B(n18453), .ZN(
        P3_U2950) );
  AOI22_X1 U21630 ( .A1(n18466), .A2(n18608), .B1(n18465), .B2(n18609), .ZN(
        n18456) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18461), .B1(
        n18543), .B2(n18610), .ZN(n18455) );
  OAI211_X1 U21632 ( .C1(n18481), .C2(n18613), .A(n18456), .B(n18455), .ZN(
        P3_U2951) );
  AOI22_X1 U21633 ( .A1(n18466), .A2(n18615), .B1(n18465), .B2(n18614), .ZN(
        n18458) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18461), .B1(
        n18543), .B2(n18616), .ZN(n18457) );
  OAI211_X1 U21635 ( .C1(n18481), .C2(n18619), .A(n18458), .B(n18457), .ZN(
        P3_U2952) );
  AOI22_X1 U21636 ( .A1(n18491), .A2(n18621), .B1(n18465), .B2(n18620), .ZN(
        n18460) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18461), .B1(
        n18543), .B2(n18622), .ZN(n18459) );
  OAI211_X1 U21638 ( .C1(n18464), .C2(n18625), .A(n18460), .B(n18459), .ZN(
        P3_U2953) );
  AOI22_X1 U21639 ( .A1(n18491), .A2(n18577), .B1(n18465), .B2(n18626), .ZN(
        n18463) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18461), .B1(
        n18543), .B2(n18629), .ZN(n18462) );
  OAI211_X1 U21641 ( .C1(n18464), .C2(n18580), .A(n18463), .B(n18462), .ZN(
        P3_U2954) );
  AOI22_X1 U21642 ( .A1(n18491), .A2(n18637), .B1(n18465), .B2(n18635), .ZN(
        n18468) );
  AOI22_X1 U21643 ( .A1(n18466), .A2(n18542), .B1(n18543), .B2(n18639), .ZN(
        n18467) );
  OAI211_X1 U21644 ( .C1(n18470), .C2(n18469), .A(n18468), .B(n18467), .ZN(
        P3_U2955) );
  NOR2_X1 U21645 ( .A1(n18675), .A2(n18471), .ZN(n18524) );
  AND2_X1 U21646 ( .A1(n18716), .A2(n18524), .ZN(n18490) );
  AOI22_X1 U21647 ( .A1(n18549), .A2(n18491), .B1(n18587), .B2(n18490), .ZN(
        n18476) );
  NOR2_X1 U21648 ( .A1(n18473), .A2(n18472), .ZN(n18589) );
  AOI22_X1 U21649 ( .A1(n18241), .A2(n18474), .B1(n18589), .B2(n18524), .ZN(
        n18492) );
  NAND2_X1 U21650 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18524), .ZN(
        n18586) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18492), .B1(
        n18592), .B2(n18572), .ZN(n18475) );
  OAI211_X1 U21652 ( .C1(n18502), .C2(n18557), .A(n18476), .B(n18475), .ZN(
        P3_U2956) );
  AOI22_X1 U21653 ( .A1(n18516), .A2(n18527), .B1(n18597), .B2(n18490), .ZN(
        n18478) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18492), .B1(
        n18598), .B2(n18572), .ZN(n18477) );
  OAI211_X1 U21655 ( .C1(n18481), .C2(n18530), .A(n18478), .B(n18477), .ZN(
        P3_U2957) );
  AOI22_X1 U21656 ( .A1(n18516), .A2(n18560), .B1(n18603), .B2(n18490), .ZN(
        n18480) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18492), .B1(
        n18604), .B2(n18572), .ZN(n18479) );
  OAI211_X1 U21658 ( .C1(n18481), .C2(n18563), .A(n18480), .B(n18479), .ZN(
        P3_U2958) );
  AOI22_X1 U21659 ( .A1(n18491), .A2(n18608), .B1(n18609), .B2(n18490), .ZN(
        n18483) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18492), .B1(
        n18610), .B2(n18572), .ZN(n18482) );
  OAI211_X1 U21661 ( .C1(n18502), .C2(n18613), .A(n18483), .B(n18482), .ZN(
        P3_U2959) );
  AOI22_X1 U21662 ( .A1(n18491), .A2(n18615), .B1(n18614), .B2(n18490), .ZN(
        n18485) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18492), .B1(
        n18616), .B2(n18572), .ZN(n18484) );
  OAI211_X1 U21664 ( .C1(n18502), .C2(n18619), .A(n18485), .B(n18484), .ZN(
        P3_U2960) );
  AOI22_X1 U21665 ( .A1(n18491), .A2(n18573), .B1(n18620), .B2(n18490), .ZN(
        n18487) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18492), .B1(
        n18622), .B2(n18572), .ZN(n18486) );
  OAI211_X1 U21667 ( .C1(n18502), .C2(n18576), .A(n18487), .B(n18486), .ZN(
        P3_U2961) );
  AOI22_X1 U21668 ( .A1(n18491), .A2(n18628), .B1(n18626), .B2(n18490), .ZN(
        n18489) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18492), .B1(
        n18629), .B2(n18572), .ZN(n18488) );
  OAI211_X1 U21670 ( .C1(n18502), .C2(n18633), .A(n18489), .B(n18488), .ZN(
        P3_U2962) );
  AOI22_X1 U21671 ( .A1(n18491), .A2(n18542), .B1(n18635), .B2(n18490), .ZN(
        n18494) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18492), .B1(
        n18639), .B2(n18572), .ZN(n18493) );
  OAI211_X1 U21673 ( .C1(n18502), .C2(n18547), .A(n18494), .B(n18493), .ZN(
        P3_U2963) );
  NAND2_X1 U21674 ( .A1(n18678), .A2(n18523), .ZN(n18643) );
  AOI21_X1 U21675 ( .B1(n18586), .B2(n18643), .A(n18548), .ZN(n18515) );
  AOI22_X1 U21676 ( .A1(n18543), .A2(n18588), .B1(n18587), .B2(n18515), .ZN(
        n18501) );
  INV_X1 U21677 ( .A(n18643), .ZN(n18627) );
  NAND2_X1 U21678 ( .A1(n18496), .A2(n18495), .ZN(n18497) );
  AOI221_X1 U21679 ( .B1(n18498), .B2(n18586), .C1(n18497), .C2(n18586), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18499) );
  OAI21_X1 U21680 ( .B1(n18627), .B2(n18499), .A(n18554), .ZN(n18517) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18517), .B1(
        n18592), .B2(n18627), .ZN(n18500) );
  OAI211_X1 U21682 ( .C1(n18595), .C2(n18502), .A(n18501), .B(n18500), .ZN(
        P3_U2964) );
  AOI22_X1 U21683 ( .A1(n18516), .A2(n18596), .B1(n18597), .B2(n18515), .ZN(
        n18504) );
  AOI22_X1 U21684 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18517), .B1(
        n18598), .B2(n18627), .ZN(n18503) );
  OAI211_X1 U21685 ( .C1(n18541), .C2(n18601), .A(n18504), .B(n18503), .ZN(
        P3_U2965) );
  AOI22_X1 U21686 ( .A1(n18516), .A2(n18602), .B1(n18603), .B2(n18515), .ZN(
        n18506) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18517), .B1(
        n18604), .B2(n18627), .ZN(n18505) );
  OAI211_X1 U21688 ( .C1(n18541), .C2(n18607), .A(n18506), .B(n18505), .ZN(
        P3_U2966) );
  AOI22_X1 U21689 ( .A1(n18516), .A2(n18608), .B1(n18609), .B2(n18515), .ZN(
        n18508) );
  AOI22_X1 U21690 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18517), .B1(
        n18610), .B2(n18627), .ZN(n18507) );
  OAI211_X1 U21691 ( .C1(n18541), .C2(n18613), .A(n18508), .B(n18507), .ZN(
        P3_U2967) );
  AOI22_X1 U21692 ( .A1(n18516), .A2(n18615), .B1(n18614), .B2(n18515), .ZN(
        n18510) );
  AOI22_X1 U21693 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18517), .B1(
        n18616), .B2(n18627), .ZN(n18509) );
  OAI211_X1 U21694 ( .C1(n18541), .C2(n18619), .A(n18510), .B(n18509), .ZN(
        P3_U2968) );
  AOI22_X1 U21695 ( .A1(n18516), .A2(n18573), .B1(n18620), .B2(n18515), .ZN(
        n18512) );
  AOI22_X1 U21696 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18517), .B1(
        n18622), .B2(n18627), .ZN(n18511) );
  OAI211_X1 U21697 ( .C1(n18541), .C2(n18576), .A(n18512), .B(n18511), .ZN(
        P3_U2969) );
  AOI22_X1 U21698 ( .A1(n18516), .A2(n18628), .B1(n18626), .B2(n18515), .ZN(
        n18514) );
  AOI22_X1 U21699 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18517), .B1(
        n18629), .B2(n18627), .ZN(n18513) );
  OAI211_X1 U21700 ( .C1(n18541), .C2(n18633), .A(n18514), .B(n18513), .ZN(
        P3_U2970) );
  AOI22_X1 U21701 ( .A1(n18516), .A2(n18542), .B1(n18635), .B2(n18515), .ZN(
        n18519) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18517), .B1(
        n18639), .B2(n18627), .ZN(n18518) );
  OAI211_X1 U21703 ( .C1(n18541), .C2(n18547), .A(n18519), .B(n18518), .ZN(
        P3_U2971) );
  NOR2_X1 U21704 ( .A1(n18521), .A2(n18520), .ZN(n18591) );
  AOI22_X1 U21705 ( .A1(n18588), .A2(n18572), .B1(n18587), .B2(n18591), .ZN(
        n18526) );
  AOI22_X1 U21706 ( .A1(n18241), .A2(n18524), .B1(n18523), .B2(n18522), .ZN(
        n18544) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18544), .B1(
        n18592), .B2(n18636), .ZN(n18525) );
  OAI211_X1 U21708 ( .C1(n18595), .C2(n18541), .A(n18526), .B(n18525), .ZN(
        P3_U2972) );
  AOI22_X1 U21709 ( .A1(n18527), .A2(n18572), .B1(n18597), .B2(n18591), .ZN(
        n18529) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18544), .B1(
        n18598), .B2(n18636), .ZN(n18528) );
  OAI211_X1 U21711 ( .C1(n18541), .C2(n18530), .A(n18529), .B(n18528), .ZN(
        P3_U2973) );
  AOI22_X1 U21712 ( .A1(n18560), .A2(n18572), .B1(n18603), .B2(n18591), .ZN(
        n18532) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18544), .B1(
        n18604), .B2(n18636), .ZN(n18531) );
  OAI211_X1 U21714 ( .C1(n18541), .C2(n18563), .A(n18532), .B(n18531), .ZN(
        P3_U2974) );
  AOI22_X1 U21715 ( .A1(n18543), .A2(n18608), .B1(n18609), .B2(n18591), .ZN(
        n18534) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18544), .B1(
        n18610), .B2(n18636), .ZN(n18533) );
  OAI211_X1 U21717 ( .C1(n18613), .C2(n18586), .A(n18534), .B(n18533), .ZN(
        P3_U2975) );
  AOI22_X1 U21718 ( .A1(n18568), .A2(n18572), .B1(n18614), .B2(n18591), .ZN(
        n18536) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18544), .B1(
        n18616), .B2(n18636), .ZN(n18535) );
  OAI211_X1 U21720 ( .C1(n18541), .C2(n18571), .A(n18536), .B(n18535), .ZN(
        P3_U2976) );
  AOI22_X1 U21721 ( .A1(n18621), .A2(n18572), .B1(n18620), .B2(n18591), .ZN(
        n18538) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18544), .B1(
        n18622), .B2(n18636), .ZN(n18537) );
  OAI211_X1 U21723 ( .C1(n18541), .C2(n18625), .A(n18538), .B(n18537), .ZN(
        P3_U2977) );
  AOI22_X1 U21724 ( .A1(n18577), .A2(n18572), .B1(n18626), .B2(n18591), .ZN(
        n18540) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18544), .B1(
        n18629), .B2(n18636), .ZN(n18539) );
  OAI211_X1 U21726 ( .C1(n18541), .C2(n18580), .A(n18540), .B(n18539), .ZN(
        P3_U2978) );
  AOI22_X1 U21727 ( .A1(n18543), .A2(n18542), .B1(n18635), .B2(n18591), .ZN(
        n18546) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18544), .B1(
        n18639), .B2(n18636), .ZN(n18545) );
  OAI211_X1 U21729 ( .C1(n18547), .C2(n18586), .A(n18546), .B(n18545), .ZN(
        P3_U2979) );
  NOR2_X1 U21730 ( .A1(n18548), .A2(n18550), .ZN(n18581) );
  AOI22_X1 U21731 ( .A1(n18549), .A2(n18572), .B1(n18587), .B2(n18581), .ZN(
        n18556) );
  NOR2_X1 U21732 ( .A1(n18572), .A2(n18627), .ZN(n18552) );
  OAI21_X1 U21733 ( .B1(n18552), .B2(n18551), .A(n18550), .ZN(n18553) );
  OAI211_X1 U21734 ( .C1(n9716), .C2(n18810), .A(n18554), .B(n18553), .ZN(
        n18583) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18583), .B1(
        n18592), .B2(n9716), .ZN(n18555) );
  OAI211_X1 U21736 ( .C1(n18557), .C2(n18643), .A(n18556), .B(n18555), .ZN(
        P3_U2980) );
  AOI22_X1 U21737 ( .A1(n18597), .A2(n18581), .B1(n18596), .B2(n18572), .ZN(
        n18559) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18583), .B1(
        n18598), .B2(n9716), .ZN(n18558) );
  OAI211_X1 U21739 ( .C1(n18601), .C2(n18643), .A(n18559), .B(n18558), .ZN(
        P3_U2981) );
  AOI22_X1 U21740 ( .A1(n18560), .A2(n18627), .B1(n18603), .B2(n18581), .ZN(
        n18562) );
  AOI22_X1 U21741 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18583), .B1(
        n18604), .B2(n9716), .ZN(n18561) );
  OAI211_X1 U21742 ( .C1(n18563), .C2(n18586), .A(n18562), .B(n18561), .ZN(
        P3_U2982) );
  AOI22_X1 U21743 ( .A1(n18564), .A2(n18627), .B1(n18609), .B2(n18581), .ZN(
        n18566) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18583), .B1(
        n18610), .B2(n9716), .ZN(n18565) );
  OAI211_X1 U21745 ( .C1(n18567), .C2(n18586), .A(n18566), .B(n18565), .ZN(
        P3_U2983) );
  AOI22_X1 U21746 ( .A1(n18568), .A2(n18627), .B1(n18614), .B2(n18581), .ZN(
        n18570) );
  AOI22_X1 U21747 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18583), .B1(
        n18616), .B2(n9716), .ZN(n18569) );
  OAI211_X1 U21748 ( .C1(n18571), .C2(n18586), .A(n18570), .B(n18569), .ZN(
        P3_U2984) );
  AOI22_X1 U21749 ( .A1(n18573), .A2(n18572), .B1(n18620), .B2(n18581), .ZN(
        n18575) );
  AOI22_X1 U21750 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18583), .B1(
        n18622), .B2(n9716), .ZN(n18574) );
  OAI211_X1 U21751 ( .C1(n18576), .C2(n18643), .A(n18575), .B(n18574), .ZN(
        P3_U2985) );
  AOI22_X1 U21752 ( .A1(n18577), .A2(n18627), .B1(n18626), .B2(n18581), .ZN(
        n18579) );
  AOI22_X1 U21753 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18583), .B1(
        n18629), .B2(n9716), .ZN(n18578) );
  OAI211_X1 U21754 ( .C1(n18580), .C2(n18586), .A(n18579), .B(n18578), .ZN(
        P3_U2986) );
  AOI22_X1 U21755 ( .A1(n18637), .A2(n18627), .B1(n18635), .B2(n18581), .ZN(
        n18585) );
  AOI22_X1 U21756 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18583), .B1(
        n18639), .B2(n9716), .ZN(n18584) );
  OAI211_X1 U21757 ( .C1(n18644), .C2(n18586), .A(n18585), .B(n18584), .ZN(
        P3_U2987) );
  AND2_X1 U21758 ( .A1(n18716), .A2(n18590), .ZN(n18634) );
  AOI22_X1 U21759 ( .A1(n18588), .A2(n18636), .B1(n18587), .B2(n18634), .ZN(
        n18594) );
  AOI22_X1 U21760 ( .A1(n18241), .A2(n18591), .B1(n18590), .B2(n18589), .ZN(
        n18640) );
  AOI22_X1 U21761 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18640), .B1(
        n18592), .B2(n18638), .ZN(n18593) );
  OAI211_X1 U21762 ( .C1(n18595), .C2(n18643), .A(n18594), .B(n18593), .ZN(
        P3_U2988) );
  AOI22_X1 U21763 ( .A1(n18597), .A2(n18634), .B1(n18596), .B2(n18627), .ZN(
        n18600) );
  AOI22_X1 U21764 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18640), .B1(
        n18598), .B2(n18638), .ZN(n18599) );
  OAI211_X1 U21765 ( .C1(n18601), .C2(n18632), .A(n18600), .B(n18599), .ZN(
        P3_U2989) );
  AOI22_X1 U21766 ( .A1(n18603), .A2(n18634), .B1(n18602), .B2(n18627), .ZN(
        n18606) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18640), .B1(
        n18604), .B2(n18638), .ZN(n18605) );
  OAI211_X1 U21768 ( .C1(n18607), .C2(n18632), .A(n18606), .B(n18605), .ZN(
        P3_U2990) );
  AOI22_X1 U21769 ( .A1(n18609), .A2(n18634), .B1(n18608), .B2(n18627), .ZN(
        n18612) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18640), .B1(
        n18610), .B2(n18638), .ZN(n18611) );
  OAI211_X1 U21771 ( .C1(n18613), .C2(n18632), .A(n18612), .B(n18611), .ZN(
        P3_U2991) );
  AOI22_X1 U21772 ( .A1(n18615), .A2(n18627), .B1(n18614), .B2(n18634), .ZN(
        n18618) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18640), .B1(
        n18616), .B2(n18638), .ZN(n18617) );
  OAI211_X1 U21774 ( .C1(n18619), .C2(n18632), .A(n18618), .B(n18617), .ZN(
        P3_U2992) );
  AOI22_X1 U21775 ( .A1(n18621), .A2(n18636), .B1(n18620), .B2(n18634), .ZN(
        n18624) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18640), .B1(
        n18622), .B2(n18638), .ZN(n18623) );
  OAI211_X1 U21777 ( .C1(n18625), .C2(n18643), .A(n18624), .B(n18623), .ZN(
        P3_U2993) );
  AOI22_X1 U21778 ( .A1(n18628), .A2(n18627), .B1(n18626), .B2(n18634), .ZN(
        n18631) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18640), .B1(
        n18629), .B2(n18638), .ZN(n18630) );
  OAI211_X1 U21780 ( .C1(n18633), .C2(n18632), .A(n18631), .B(n18630), .ZN(
        P3_U2994) );
  AOI22_X1 U21781 ( .A1(n18637), .A2(n18636), .B1(n18635), .B2(n18634), .ZN(
        n18642) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18640), .B1(
        n18639), .B2(n18638), .ZN(n18641) );
  OAI211_X1 U21783 ( .C1(n18644), .C2(n18643), .A(n18642), .B(n18641), .ZN(
        P3_U2995) );
  NOR2_X1 U21784 ( .A1(n18658), .A2(n9766), .ZN(n18647) );
  OAI222_X1 U21785 ( .A1(n18651), .A2(n18650), .B1(n18649), .B2(n18648), .C1(
        n18647), .C2(n18646), .ZN(n18853) );
  OAI21_X1 U21786 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18652), .ZN(n18653) );
  OAI211_X1 U21787 ( .C1(n18655), .C2(n18689), .A(n18654), .B(n18653), .ZN(
        n18701) );
  OAI21_X1 U21788 ( .B1(n21016), .B2(n18670), .A(n18656), .ZN(n18681) );
  OR2_X1 U21789 ( .A1(n18681), .A2(n18657), .ZN(n18671) );
  NAND2_X1 U21790 ( .A1(n18826), .A2(n18685), .ZN(n18663) );
  AOI22_X1 U21791 ( .A1(n18659), .A2(n18671), .B1(n18658), .B2(n18663), .ZN(
        n18814) );
  NOR2_X1 U21792 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18814), .ZN(
        n18668) );
  AOI21_X1 U21793 ( .B1(n18662), .B2(n18661), .A(n18660), .ZN(n18683) );
  OAI21_X1 U21794 ( .B1(n18664), .B2(n18683), .A(n18663), .ZN(n18665) );
  AOI21_X1 U21795 ( .B1(n18666), .B2(n18673), .A(n18665), .ZN(n18811) );
  NAND2_X1 U21796 ( .A1(n18689), .A2(n18811), .ZN(n18667) );
  AOI22_X1 U21797 ( .A1(n18689), .A2(n18668), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18667), .ZN(n18699) );
  NAND2_X1 U21798 ( .A1(n18670), .A2(n18669), .ZN(n18672) );
  AOI22_X1 U21799 ( .A1(n18832), .A2(n18672), .B1(n18834), .B2(n18671), .ZN(
        n18830) );
  AOI22_X1 U21800 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18673), .B1(
        n18672), .B2(n21016), .ZN(n18676) );
  INV_X1 U21801 ( .A(n18676), .ZN(n18836) );
  NOR3_X1 U21802 ( .A1(n18675), .A2(n18674), .A3(n18836), .ZN(n18677) );
  OAI22_X1 U21803 ( .A1(n18830), .A2(n18677), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18676), .ZN(n18679) );
  AOI21_X1 U21804 ( .B1(n18689), .B2(n18679), .A(n18678), .ZN(n18691) );
  NAND2_X1 U21805 ( .A1(n18834), .A2(n18826), .ZN(n18680) );
  OAI221_X1 U21806 ( .B1(n18834), .B2(n18826), .C1(n18682), .C2(n18681), .A(
        n18680), .ZN(n18687) );
  INV_X1 U21807 ( .A(n18683), .ZN(n18684) );
  NAND3_X1 U21808 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18685), .A3(
        n18684), .ZN(n18686) );
  OAI211_X1 U21809 ( .C1(n18822), .C2(n18688), .A(n18687), .B(n18686), .ZN(
        n18824) );
  AOI22_X1 U21810 ( .A1(n18690), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18824), .B2(n18689), .ZN(n18694) );
  OAI21_X1 U21811 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18691), .A(
        n18694), .ZN(n18693) );
  AOI21_X1 U21812 ( .B1(n18691), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18692) );
  NAND2_X1 U21813 ( .A1(n18693), .A2(n18692), .ZN(n18698) );
  INV_X1 U21814 ( .A(n18694), .ZN(n18695) );
  AOI21_X1 U21815 ( .B1(n20840), .B2(n18696), .A(n18695), .ZN(n18697) );
  AOI222_X1 U21816 ( .A1(n18699), .A2(n18698), .B1(n18699), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18698), .C2(n18697), .ZN(
        n18700) );
  NOR4_X1 U21817 ( .A1(n18702), .A2(n18853), .A3(n18701), .A4(n18700), .ZN(
        n18714) );
  INV_X1 U21818 ( .A(n18858), .ZN(n18703) );
  AOI22_X1 U21819 ( .A1(n18835), .A2(n18703), .B1(n18864), .B2(n17450), .ZN(
        n18704) );
  INV_X1 U21820 ( .A(n18704), .ZN(n18710) );
  OAI211_X1 U21821 ( .C1(n18706), .C2(n18705), .A(n18862), .B(n18714), .ZN(
        n18809) );
  OAI21_X1 U21822 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18707), .A(n18809), 
        .ZN(n18715) );
  NOR2_X1 U21823 ( .A1(n18708), .A2(n18715), .ZN(n18709) );
  MUX2_X1 U21824 ( .A(n18710), .B(n18709), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18712) );
  OAI211_X1 U21825 ( .C1(n18714), .C2(n18713), .A(n18712), .B(n18711), .ZN(
        P3_U2996) );
  NAND2_X1 U21826 ( .A1(n18864), .A2(n17450), .ZN(n18720) );
  NAND4_X1 U21827 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18864), .A4(n18856), .ZN(n18722) );
  INV_X1 U21828 ( .A(n18715), .ZN(n18717) );
  NAND3_X1 U21829 ( .A1(n18718), .A2(n18717), .A3(n18716), .ZN(n18719) );
  NAND4_X1 U21830 ( .A1(n18721), .A2(n18720), .A3(n18722), .A4(n18719), .ZN(
        P3_U2997) );
  AND4_X1 U21831 ( .A1(n18858), .A2(n18723), .A3(n18722), .A4(n18808), .ZN(
        P3_U2998) );
  AND2_X1 U21832 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18804), .ZN(
        P3_U2999) );
  AND2_X1 U21833 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18724), .ZN(
        P3_U3000) );
  AND2_X1 U21834 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18724), .ZN(
        P3_U3001) );
  AND2_X1 U21835 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18724), .ZN(
        P3_U3002) );
  AND2_X1 U21836 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18724), .ZN(
        P3_U3003) );
  AND2_X1 U21837 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18724), .ZN(
        P3_U3004) );
  AND2_X1 U21838 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18724), .ZN(
        P3_U3005) );
  AND2_X1 U21839 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18724), .ZN(
        P3_U3006) );
  AND2_X1 U21840 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18724), .ZN(
        P3_U3007) );
  AND2_X1 U21841 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18724), .ZN(
        P3_U3008) );
  AND2_X1 U21842 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18724), .ZN(
        P3_U3009) );
  AND2_X1 U21843 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18724), .ZN(
        P3_U3010) );
  INV_X1 U21844 ( .A(P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20904) );
  NOR2_X1 U21845 ( .A1(n20904), .A2(n18807), .ZN(P3_U3011) );
  AND2_X1 U21846 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18724), .ZN(
        P3_U3012) );
  AND2_X1 U21847 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18724), .ZN(
        P3_U3013) );
  INV_X1 U21848 ( .A(P3_DATAWIDTH_REG_16__SCAN_IN), .ZN(n21038) );
  NOR2_X1 U21849 ( .A1(n21038), .A2(n18807), .ZN(P3_U3014) );
  AND2_X1 U21850 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18724), .ZN(
        P3_U3015) );
  AND2_X1 U21851 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18724), .ZN(
        P3_U3016) );
  AND2_X1 U21852 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18724), .ZN(
        P3_U3017) );
  AND2_X1 U21853 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18724), .ZN(
        P3_U3018) );
  AND2_X1 U21854 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18724), .ZN(
        P3_U3019) );
  AND2_X1 U21855 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18724), .ZN(
        P3_U3020) );
  AND2_X1 U21856 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18724), .ZN(P3_U3021) );
  AND2_X1 U21857 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18724), .ZN(P3_U3022) );
  AND2_X1 U21858 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18724), .ZN(P3_U3023) );
  AND2_X1 U21859 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18724), .ZN(P3_U3024) );
  AND2_X1 U21860 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18804), .ZN(P3_U3025) );
  AND2_X1 U21861 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18804), .ZN(P3_U3026) );
  AND2_X1 U21862 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18804), .ZN(P3_U3027) );
  AND2_X1 U21863 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18804), .ZN(P3_U3028) );
  NAND2_X1 U21864 ( .A1(n18864), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18738) );
  OAI21_X1 U21865 ( .B1(n18725), .B2(n20717), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18726) );
  AOI22_X1 U21866 ( .A1(n18734), .A2(n21050), .B1(n18868), .B2(n18726), .ZN(
        n18728) );
  NAND3_X1 U21867 ( .A1(NA), .A2(n18734), .A3(n18729), .ZN(n18727) );
  OAI211_X1 U21868 ( .C1(P3_STATE_REG_2__SCAN_IN), .C2(n18738), .A(n18728), 
        .B(n18727), .ZN(P3_U3029) );
  NOR3_X1 U21869 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n18729), .A3(n20717), 
        .ZN(n18730) );
  AOI221_X1 U21870 ( .B1(n18731), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20717), .C2(P3_REQUESTPENDING_REG_SCAN_IN), .A(n18730), .ZN(n18733)
         );
  OAI211_X1 U21871 ( .C1(n18733), .C2(n18734), .A(n18738), .B(n18732), .ZN(
        P3_U3030) );
  INV_X1 U21872 ( .A(NA), .ZN(n20722) );
  OAI21_X1 U21873 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n20722), .A(n18734), 
        .ZN(n18737) );
  OAI222_X1 U21874 ( .A1(n20717), .A2(n21050), .B1(P3_STATE_REG_1__SCAN_IN), 
        .B2(P3_REQUESTPENDING_REG_SCAN_IN), .C1(n18738), .C2(NA), .ZN(n18735)
         );
  OAI211_X1 U21875 ( .C1(P3_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .B(n18735), .ZN(n18736) );
  OAI221_X1 U21876 ( .B1(n21050), .B2(n18738), .C1(n21050), .C2(n18737), .A(
        n18736), .ZN(P3_U3031) );
  INV_X1 U21877 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18740) );
  OAI222_X1 U21878 ( .A1(n18842), .A2(n18794), .B1(n18739), .B2(n18869), .C1(
        n18740), .C2(n18791), .ZN(P3_U3032) );
  OAI222_X1 U21879 ( .A1(n18791), .A2(n18742), .B1(n18741), .B2(n18800), .C1(
        n18740), .C2(n18794), .ZN(P3_U3033) );
  OAI222_X1 U21880 ( .A1(n18791), .A2(n18744), .B1(n18743), .B2(n18800), .C1(
        n18742), .C2(n18794), .ZN(P3_U3034) );
  INV_X1 U21881 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18747) );
  OAI222_X1 U21882 ( .A1(n18791), .A2(n18747), .B1(n18745), .B2(n18800), .C1(
        n18744), .C2(n18794), .ZN(P3_U3035) );
  OAI222_X1 U21883 ( .A1(n18747), .A2(n18794), .B1(n18746), .B2(n18800), .C1(
        n18748), .C2(n18791), .ZN(P3_U3036) );
  OAI222_X1 U21884 ( .A1(n18791), .A2(n18750), .B1(n18749), .B2(n18800), .C1(
        n18748), .C2(n18794), .ZN(P3_U3037) );
  OAI222_X1 U21885 ( .A1(n18791), .A2(n20903), .B1(n20855), .B2(n18800), .C1(
        n18750), .C2(n18794), .ZN(P3_U3038) );
  OAI222_X1 U21886 ( .A1(n20903), .A2(n18794), .B1(n20954), .B2(n18800), .C1(
        n18751), .C2(n18791), .ZN(P3_U3039) );
  OAI222_X1 U21887 ( .A1(n18791), .A2(n18753), .B1(n18752), .B2(n18800), .C1(
        n18751), .C2(n18794), .ZN(P3_U3040) );
  OAI222_X1 U21888 ( .A1(n18791), .A2(n18754), .B1(n21019), .B2(n18800), .C1(
        n18753), .C2(n18794), .ZN(P3_U3041) );
  OAI222_X1 U21889 ( .A1(n18791), .A2(n18756), .B1(n18755), .B2(n18800), .C1(
        n18754), .C2(n18794), .ZN(P3_U3042) );
  OAI222_X1 U21890 ( .A1(n18791), .A2(n18758), .B1(n18757), .B2(n18800), .C1(
        n18756), .C2(n18794), .ZN(P3_U3043) );
  OAI222_X1 U21891 ( .A1(n18791), .A2(n18761), .B1(n18759), .B2(n18800), .C1(
        n18758), .C2(n18794), .ZN(P3_U3044) );
  OAI222_X1 U21892 ( .A1(n18761), .A2(n18794), .B1(n18760), .B2(n18869), .C1(
        n18762), .C2(n18791), .ZN(P3_U3045) );
  OAI222_X1 U21893 ( .A1(n18791), .A2(n18763), .B1(n20829), .B2(n18869), .C1(
        n18762), .C2(n18794), .ZN(P3_U3046) );
  INV_X1 U21894 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18765) );
  OAI222_X1 U21895 ( .A1(n18791), .A2(n18765), .B1(n18764), .B2(n18869), .C1(
        n18763), .C2(n18794), .ZN(P3_U3047) );
  OAI222_X1 U21896 ( .A1(n18791), .A2(n18767), .B1(n18766), .B2(n18869), .C1(
        n18765), .C2(n18794), .ZN(P3_U3048) );
  OAI222_X1 U21897 ( .A1(n18791), .A2(n18770), .B1(n18768), .B2(n18869), .C1(
        n18767), .C2(n18794), .ZN(P3_U3049) );
  OAI222_X1 U21898 ( .A1(n18770), .A2(n18794), .B1(n18769), .B2(n18869), .C1(
        n18771), .C2(n18791), .ZN(P3_U3050) );
  OAI222_X1 U21899 ( .A1(n18791), .A2(n18774), .B1(n18772), .B2(n18869), .C1(
        n18771), .C2(n18794), .ZN(P3_U3051) );
  OAI222_X1 U21900 ( .A1(n18774), .A2(n18794), .B1(n18773), .B2(n18869), .C1(
        n18775), .C2(n18791), .ZN(P3_U3052) );
  OAI222_X1 U21901 ( .A1(n18791), .A2(n18778), .B1(n18776), .B2(n18869), .C1(
        n18775), .C2(n18794), .ZN(P3_U3053) );
  OAI222_X1 U21902 ( .A1(n18778), .A2(n18794), .B1(n18777), .B2(n18869), .C1(
        n18779), .C2(n18791), .ZN(P3_U3054) );
  OAI222_X1 U21903 ( .A1(n18791), .A2(n18781), .B1(n18780), .B2(n18869), .C1(
        n18779), .C2(n18794), .ZN(P3_U3055) );
  OAI222_X1 U21904 ( .A1(n18791), .A2(n18783), .B1(n18782), .B2(n18800), .C1(
        n18781), .C2(n18794), .ZN(P3_U3056) );
  OAI222_X1 U21905 ( .A1(n18791), .A2(n18785), .B1(n18784), .B2(n18800), .C1(
        n18783), .C2(n18794), .ZN(P3_U3057) );
  OAI222_X1 U21906 ( .A1(n18791), .A2(n18788), .B1(n18786), .B2(n18800), .C1(
        n18785), .C2(n18794), .ZN(P3_U3058) );
  OAI222_X1 U21907 ( .A1(n18788), .A2(n18794), .B1(n18787), .B2(n18800), .C1(
        n18789), .C2(n18791), .ZN(P3_U3059) );
  OAI222_X1 U21908 ( .A1(n18791), .A2(n18793), .B1(n18790), .B2(n18800), .C1(
        n18789), .C2(n18794), .ZN(P3_U3060) );
  OAI222_X1 U21909 ( .A1(n18794), .A2(n18793), .B1(n18792), .B2(n18800), .C1(
        n21051), .C2(n18791), .ZN(P3_U3061) );
  INV_X1 U21910 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18795) );
  AOI22_X1 U21911 ( .A1(n18869), .A2(n18796), .B1(n18795), .B2(n18868), .ZN(
        P3_U3274) );
  INV_X1 U21912 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18844) );
  INV_X1 U21913 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18797) );
  AOI22_X1 U21914 ( .A1(n18869), .A2(n18844), .B1(n18797), .B2(n18868), .ZN(
        P3_U3275) );
  INV_X1 U21915 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18798) );
  AOI22_X1 U21916 ( .A1(n18800), .A2(n18799), .B1(n18798), .B2(n18868), .ZN(
        P3_U3276) );
  INV_X1 U21917 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18850) );
  INV_X1 U21918 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18801) );
  AOI22_X1 U21919 ( .A1(n18869), .A2(n18850), .B1(n18801), .B2(n18868), .ZN(
        P3_U3277) );
  INV_X1 U21920 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18803) );
  INV_X1 U21921 ( .A(n18805), .ZN(n18802) );
  AOI21_X1 U21922 ( .B1(n18804), .B2(n18803), .A(n18802), .ZN(P3_U3280) );
  OAI21_X1 U21923 ( .B1(n18807), .B2(n18806), .A(n18805), .ZN(P3_U3281) );
  OAI221_X1 U21924 ( .B1(n18810), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18810), 
        .C2(n18809), .A(n18808), .ZN(P3_U3282) );
  NOR2_X1 U21925 ( .A1(n18811), .A2(n18829), .ZN(n18812) );
  NOR2_X1 U21926 ( .A1(n18812), .A2(n18841), .ZN(n18818) );
  INV_X1 U21927 ( .A(n18813), .ZN(n18816) );
  NOR3_X1 U21928 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18814), .A3(
        n18829), .ZN(n18815) );
  AOI21_X1 U21929 ( .B1(n18816), .B2(n18835), .A(n18815), .ZN(n18817) );
  OAI22_X1 U21930 ( .A1(n18819), .A2(n18818), .B1(n18841), .B2(n18817), .ZN(
        P3_U3285) );
  NAND2_X1 U21931 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18827) );
  INV_X1 U21932 ( .A(n18827), .ZN(n18823) );
  AOI22_X1 U21933 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n18821), .B2(n18820), .ZN(
        n18828) );
  AOI222_X1 U21934 ( .A1(n18824), .A2(n18837), .B1(n18823), .B2(n18828), .C1(
        n18835), .C2(n18822), .ZN(n18825) );
  AOI22_X1 U21935 ( .A1(n18841), .A2(n18826), .B1(n18825), .B2(n18839), .ZN(
        P3_U3288) );
  OAI22_X1 U21936 ( .A1(n18830), .A2(n18829), .B1(n18828), .B2(n18827), .ZN(
        n18831) );
  AOI21_X1 U21937 ( .B1(n18835), .B2(n18832), .A(n18831), .ZN(n18833) );
  AOI22_X1 U21938 ( .A1(n18841), .A2(n18834), .B1(n18833), .B2(n18839), .ZN(
        P3_U3289) );
  AOI222_X1 U21939 ( .A1(n18838), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18837), 
        .B2(n18836), .C1(n21016), .C2(n18835), .ZN(n18840) );
  AOI22_X1 U21940 ( .A1(n18841), .A2(n21016), .B1(n18840), .B2(n18839), .ZN(
        P3_U3290) );
  AOI21_X1 U21941 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18843) );
  AOI22_X1 U21942 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18843), .B2(n18842), .ZN(n18845) );
  AOI22_X1 U21943 ( .A1(n18846), .A2(n18845), .B1(n18844), .B2(n18849), .ZN(
        P3_U3292) );
  NOR2_X1 U21944 ( .A1(n18849), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18847) );
  AOI22_X1 U21945 ( .A1(n18850), .A2(n18849), .B1(n18848), .B2(n18847), .ZN(
        P3_U3293) );
  INV_X1 U21946 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18851) );
  AOI22_X1 U21947 ( .A1(n18869), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18851), 
        .B2(n18868), .ZN(P3_U3294) );
  MUX2_X1 U21948 ( .A(P3_MORE_REG_SCAN_IN), .B(n18853), .S(n18852), .Z(
        P3_U3295) );
  OAI21_X1 U21949 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18855), .A(n18854), 
        .ZN(n18857) );
  AOI211_X1 U21950 ( .C1(n18871), .C2(n18857), .A(n18864), .B(n18856), .ZN(
        n18860) );
  OAI21_X1 U21951 ( .B1(n18860), .B2(n18859), .A(n18858), .ZN(n18867) );
  OAI22_X1 U21952 ( .A1(n18864), .A2(n18863), .B1(n18862), .B2(n18861), .ZN(
        n18865) );
  NOR2_X1 U21953 ( .A1(n18873), .A2(n18865), .ZN(n18866) );
  MUX2_X1 U21954 ( .A(n18867), .B(P3_REQUESTPENDING_REG_SCAN_IN), .S(n18866), 
        .Z(P3_U3296) );
  INV_X1 U21955 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n21006) );
  AOI22_X1 U21956 ( .A1(n18869), .A2(n21006), .B1(n20937), .B2(n18868), .ZN(
        P3_U3297) );
  OAI21_X1 U21957 ( .B1(n18874), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n18872), 
        .ZN(n18870) );
  OAI21_X1 U21958 ( .B1(n18872), .B2(n18871), .A(n18870), .ZN(P3_U3298) );
  NOR3_X1 U21959 ( .A1(P3_MEMORYFETCH_REG_SCAN_IN), .A2(n18874), .A3(n18873), 
        .ZN(n18876) );
  NOR2_X1 U21960 ( .A1(n18876), .A2(n18875), .ZN(P3_U3299) );
  INV_X1 U21961 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18877) );
  NAND2_X1 U21962 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n21048), .ZN(n19753) );
  NAND2_X1 U21963 ( .A1(n19746), .A2(n19745), .ZN(n19750) );
  OAI21_X1 U21964 ( .B1(n19746), .B2(n19753), .A(n19750), .ZN(n19824) );
  OAI21_X1 U21965 ( .B1(n19746), .B2(n18877), .A(n19744), .ZN(P2_U2815) );
  AOI22_X1 U21966 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18878), .B1(n19875), 
        .B2(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18879) );
  INV_X1 U21967 ( .A(n18879), .ZN(P2_U2816) );
  NAND2_X1 U21968 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19746), .ZN(n19891) );
  AOI21_X1 U21969 ( .B1(n19746), .B2(n21048), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18880) );
  AOI22_X1 U21970 ( .A1(n19805), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18880), 
        .B2(n19891), .ZN(P2_U2817) );
  OAI21_X1 U21971 ( .B1(n19757), .B2(BS16), .A(n19824), .ZN(n19822) );
  OAI21_X1 U21972 ( .B1(n19824), .B2(n19882), .A(n19822), .ZN(P2_U2818) );
  NOR2_X1 U21973 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n21091) );
  AOI211_X1 U21974 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18881) );
  INV_X1 U21975 ( .A(P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n20842) );
  INV_X1 U21976 ( .A(P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20864) );
  AND4_X1 U21977 ( .A1(n21091), .A2(n18881), .A3(n20842), .A4(n20864), .ZN(
        n18889) );
  NOR4_X1 U21978 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18888) );
  NOR4_X1 U21979 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_6__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n18887) );
  NOR4_X1 U21980 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18885) );
  NOR4_X1 U21981 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18884) );
  NOR4_X1 U21982 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18883) );
  NOR4_X1 U21983 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18882) );
  AND4_X1 U21984 ( .A1(n18885), .A2(n18884), .A3(n18883), .A4(n18882), .ZN(
        n18886) );
  NAND4_X1 U21985 ( .A1(n18889), .A2(n18888), .A3(n18887), .A4(n18886), .ZN(
        n18895) );
  NOR2_X1 U21986 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18895), .ZN(n18890) );
  INV_X1 U21987 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19820) );
  AOI22_X1 U21988 ( .A1(n18890), .A2(n19060), .B1(n18895), .B2(n19820), .ZN(
        P2_U2820) );
  OR3_X1 U21989 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18894) );
  INV_X1 U21990 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19818) );
  AOI22_X1 U21991 ( .A1(n18890), .A2(n18894), .B1(n18895), .B2(n19818), .ZN(
        P2_U2821) );
  INV_X1 U21992 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19823) );
  NAND2_X1 U21993 ( .A1(n18890), .A2(n19823), .ZN(n18893) );
  INV_X1 U21994 ( .A(n18895), .ZN(n18896) );
  OAI21_X1 U21995 ( .B1(n19060), .B2(n19763), .A(n18896), .ZN(n18891) );
  OAI21_X1 U21996 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18896), .A(n18891), 
        .ZN(n18892) );
  OAI221_X1 U21997 ( .B1(n18893), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18893), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18892), .ZN(P2_U2822) );
  INV_X1 U21998 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19817) );
  OAI221_X1 U21999 ( .B1(n18896), .B2(n19817), .C1(n18895), .C2(n18894), .A(
        n18893), .ZN(P2_U2823) );
  NAND2_X1 U22000 ( .A1(n19032), .A2(n18897), .ZN(n18898) );
  XOR2_X1 U22001 ( .A(n18899), .B(n18898), .Z(n18908) );
  AOI22_X1 U22002 ( .A1(n18900), .A2(n19041), .B1(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19043), .ZN(n18901) );
  OAI211_X1 U22003 ( .C1(n19790), .C2(n19061), .A(n18901), .B(n19045), .ZN(
        n18902) );
  AOI21_X1 U22004 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19065), .A(n18902), .ZN(
        n18907) );
  INV_X1 U22005 ( .A(n18903), .ZN(n18904) );
  AOI22_X1 U22006 ( .A1(n18905), .A2(n19042), .B1(n18904), .B2(n19070), .ZN(
        n18906) );
  OAI211_X1 U22007 ( .C1(n19741), .C2(n18908), .A(n18907), .B(n18906), .ZN(
        P2_U2836) );
  NOR2_X1 U22008 ( .A1(n19052), .A2(n18909), .ZN(n18911) );
  XOR2_X1 U22009 ( .A(n18911), .B(n18910), .Z(n18920) );
  AOI22_X1 U22010 ( .A1(n18912), .A2(n19041), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19043), .ZN(n18913) );
  OAI211_X1 U22011 ( .C1(n19789), .C2(n19061), .A(n18913), .B(n19045), .ZN(
        n18914) );
  AOI21_X1 U22012 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n19065), .A(n18914), .ZN(
        n18919) );
  OAI22_X1 U22013 ( .A1(n18916), .A2(n19063), .B1(n18915), .B2(n19047), .ZN(
        n18917) );
  INV_X1 U22014 ( .A(n18917), .ZN(n18918) );
  OAI211_X1 U22015 ( .C1(n19741), .C2(n18920), .A(n18919), .B(n18918), .ZN(
        P2_U2837) );
  NAND2_X1 U22016 ( .A1(n19032), .A2(n18921), .ZN(n18922) );
  XOR2_X1 U22017 ( .A(n18923), .B(n18922), .Z(n18933) );
  OAI21_X1 U22018 ( .B1(n19787), .B2(n19061), .A(n19045), .ZN(n18927) );
  OAI22_X1 U22019 ( .A1(n18925), .A2(n19067), .B1(n18924), .B2(n19072), .ZN(
        n18926) );
  AOI211_X1 U22020 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19065), .A(n18927), .B(
        n18926), .ZN(n18932) );
  NOR2_X1 U22021 ( .A1(n18928), .A2(n19047), .ZN(n18929) );
  AOI21_X1 U22022 ( .B1(n18930), .B2(n19042), .A(n18929), .ZN(n18931) );
  OAI211_X1 U22023 ( .C1(n19741), .C2(n18933), .A(n18932), .B(n18931), .ZN(
        P2_U2838) );
  NOR2_X1 U22024 ( .A1(n19052), .A2(n18934), .ZN(n18936) );
  XOR2_X1 U22025 ( .A(n18936), .B(n18935), .Z(n18946) );
  OAI21_X1 U22026 ( .B1(n19785), .B2(n19061), .A(n19045), .ZN(n18941) );
  INV_X1 U22027 ( .A(n18937), .ZN(n18939) );
  OAI22_X1 U22028 ( .A1(n18939), .A2(n19067), .B1(n18938), .B2(n19072), .ZN(
        n18940) );
  AOI211_X1 U22029 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19065), .A(n18941), .B(
        n18940), .ZN(n18945) );
  NOR2_X1 U22030 ( .A1(n18942), .A2(n19047), .ZN(n18943) );
  AOI21_X1 U22031 ( .B1(n19088), .B2(n19042), .A(n18943), .ZN(n18944) );
  OAI211_X1 U22032 ( .C1(n19741), .C2(n18946), .A(n18945), .B(n18944), .ZN(
        P2_U2839) );
  XOR2_X1 U22033 ( .A(n18948), .B(n18947), .Z(n18956) );
  OAI21_X1 U22034 ( .B1(n19781), .B2(n19061), .A(n19045), .ZN(n18952) );
  INV_X1 U22035 ( .A(n18949), .ZN(n18950) );
  OAI22_X1 U22036 ( .A1(n18950), .A2(n19067), .B1(n10056), .B2(n19072), .ZN(
        n18951) );
  AOI211_X1 U22037 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n19065), .A(n18952), .B(
        n18951), .ZN(n18955) );
  AOI22_X1 U22038 ( .A1(n19092), .A2(n19042), .B1(n18953), .B2(n19070), .ZN(
        n18954) );
  OAI211_X1 U22039 ( .C1(n19741), .C2(n18956), .A(n18955), .B(n18954), .ZN(
        P2_U2841) );
  INV_X1 U22040 ( .A(n18957), .ZN(n18958) );
  AOI22_X1 U22041 ( .A1(n18958), .A2(n19041), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19043), .ZN(n18959) );
  OAI211_X1 U22042 ( .C1(n11549), .C2(n19061), .A(n18959), .B(n19045), .ZN(
        n18960) );
  AOI21_X1 U22043 ( .B1(P2_EBX_REG_12__SCAN_IN), .B2(n19065), .A(n18960), .ZN(
        n18967) );
  NOR2_X1 U22044 ( .A1(n19052), .A2(n18961), .ZN(n18963) );
  XNOR2_X1 U22045 ( .A(n18963), .B(n18962), .ZN(n18965) );
  AOI22_X1 U22046 ( .A1(n18965), .A2(n19036), .B1(n18964), .B2(n19070), .ZN(
        n18966) );
  OAI211_X1 U22047 ( .C1(n18968), .C2(n19063), .A(n18967), .B(n18966), .ZN(
        P2_U2843) );
  AOI22_X1 U22048 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19043), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n19065), .ZN(n18969) );
  OAI21_X1 U22049 ( .B1(n18970), .B2(n19067), .A(n18969), .ZN(n18971) );
  AOI211_X1 U22050 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19030), .A(n19029), 
        .B(n18971), .ZN(n18979) );
  NAND2_X1 U22051 ( .A1(n19032), .A2(n18972), .ZN(n18973) );
  XNOR2_X1 U22052 ( .A(n18974), .B(n18973), .ZN(n18977) );
  INV_X1 U22053 ( .A(n18975), .ZN(n18976) );
  AOI22_X1 U22054 ( .A1(n18977), .A2(n19036), .B1(n18976), .B2(n19070), .ZN(
        n18978) );
  OAI211_X1 U22055 ( .C1(n18980), .C2(n19063), .A(n18979), .B(n18978), .ZN(
        P2_U2844) );
  INV_X1 U22056 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18981) );
  OAI22_X1 U22057 ( .A1(n18982), .A2(n19067), .B1(n18981), .B2(n19072), .ZN(
        n18983) );
  INV_X1 U22058 ( .A(n18983), .ZN(n18984) );
  OAI211_X1 U22059 ( .C1(n11508), .C2(n19061), .A(n18984), .B(n19045), .ZN(
        n18985) );
  AOI21_X1 U22060 ( .B1(P2_EBX_REG_10__SCAN_IN), .B2(n19065), .A(n18985), .ZN(
        n18992) );
  NOR2_X1 U22061 ( .A1(n19052), .A2(n18986), .ZN(n18988) );
  XNOR2_X1 U22062 ( .A(n18988), .B(n18987), .ZN(n18990) );
  AOI22_X1 U22063 ( .A1(n18990), .A2(n19036), .B1(n18989), .B2(n19070), .ZN(
        n18991) );
  OAI211_X1 U22064 ( .C1(n19098), .C2(n19063), .A(n18992), .B(n18991), .ZN(
        P2_U2845) );
  NAND2_X1 U22065 ( .A1(n19032), .A2(n18993), .ZN(n18995) );
  XOR2_X1 U22066 ( .A(n18995), .B(n18994), .Z(n19003) );
  AOI22_X1 U22067 ( .A1(n18996), .A2(n19041), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19065), .ZN(n18997) );
  OAI211_X1 U22068 ( .C1(n19773), .C2(n19061), .A(n18997), .B(n19045), .ZN(
        n19001) );
  OAI22_X1 U22069 ( .A1(n18999), .A2(n19063), .B1(n18998), .B2(n19047), .ZN(
        n19000) );
  AOI211_X1 U22070 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19043), .A(
        n19001), .B(n19000), .ZN(n19002) );
  OAI21_X1 U22071 ( .B1(n19003), .B2(n19741), .A(n19002), .ZN(P2_U2846) );
  NOR2_X1 U22072 ( .A1(n19052), .A2(n19004), .ZN(n19006) );
  XOR2_X1 U22073 ( .A(n19006), .B(n19005), .Z(n19013) );
  AOI22_X1 U22074 ( .A1(n19007), .A2(n19041), .B1(n19043), .B2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19008) );
  OAI211_X1 U22075 ( .C1(n11468), .C2(n19061), .A(n19008), .B(n19045), .ZN(
        n19009) );
  AOI21_X1 U22076 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(n19065), .A(n19009), .ZN(
        n19012) );
  AOI22_X1 U22077 ( .A1(n19010), .A2(n19070), .B1(n19042), .B2(n19100), .ZN(
        n19011) );
  OAI211_X1 U22078 ( .C1(n19741), .C2(n19013), .A(n19012), .B(n19011), .ZN(
        P2_U2847) );
  OAI21_X1 U22079 ( .B1(n19769), .B2(n19061), .A(n19045), .ZN(n19017) );
  OAI22_X1 U22080 ( .A1(n19015), .A2(n19067), .B1(n19014), .B2(n13461), .ZN(
        n19016) );
  AOI211_X1 U22081 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19043), .A(
        n19017), .B(n19016), .ZN(n19024) );
  NOR2_X1 U22082 ( .A1(n19052), .A2(n19018), .ZN(n19020) );
  XNOR2_X1 U22083 ( .A(n19020), .B(n19019), .ZN(n19022) );
  AOI22_X1 U22084 ( .A1(n19022), .A2(n19036), .B1(n19021), .B2(n19070), .ZN(
        n19023) );
  OAI211_X1 U22085 ( .C1(n19063), .C2(n19025), .A(n19024), .B(n19023), .ZN(
        P2_U2849) );
  AOI22_X1 U22086 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19043), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19065), .ZN(n19026) );
  OAI21_X1 U22087 ( .B1(n19027), .B2(n19067), .A(n19026), .ZN(n19028) );
  AOI211_X1 U22088 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19030), .A(n19029), .B(
        n19028), .ZN(n19039) );
  NAND2_X1 U22089 ( .A1(n19032), .A2(n19031), .ZN(n19033) );
  XNOR2_X1 U22090 ( .A(n19034), .B(n19033), .ZN(n19037) );
  AOI22_X1 U22091 ( .A1(n19037), .A2(n19036), .B1(n19035), .B2(n19070), .ZN(
        n19038) );
  OAI211_X1 U22092 ( .C1(n19063), .C2(n19112), .A(n19039), .B(n19038), .ZN(
        P2_U2850) );
  AOI22_X1 U22093 ( .A1(n19041), .A2(n19040), .B1(n19065), .B2(
        P2_EBX_REG_4__SCAN_IN), .ZN(n19059) );
  AOI22_X1 U22094 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19043), .B1(
        n19042), .B2(n19185), .ZN(n19044) );
  OAI211_X1 U22095 ( .C1(n11438), .C2(n19061), .A(n19045), .B(n19044), .ZN(
        n19046) );
  INV_X1 U22096 ( .A(n19046), .ZN(n19058) );
  OAI22_X1 U22097 ( .A1(n19108), .A2(n19049), .B1(n19048), .B2(n19047), .ZN(
        n19050) );
  INV_X1 U22098 ( .A(n19050), .ZN(n19057) );
  INV_X1 U22099 ( .A(n19166), .ZN(n19055) );
  NOR2_X1 U22100 ( .A1(n19052), .A2(n19051), .ZN(n19054) );
  AOI21_X1 U22101 ( .B1(n19055), .B2(n19054), .A(n19741), .ZN(n19053) );
  OAI21_X1 U22102 ( .B1(n19055), .B2(n19054), .A(n19053), .ZN(n19056) );
  NAND4_X1 U22103 ( .A1(n19059), .A2(n19058), .A3(n19057), .A4(n19056), .ZN(
        P2_U2851) );
  OAI22_X1 U22104 ( .A1(n19063), .A2(n19062), .B1(n19061), .B2(n19060), .ZN(
        n19064) );
  AOI21_X1 U22105 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n19065), .A(n19064), .ZN(
        n19066) );
  OAI21_X1 U22106 ( .B1(n19068), .B2(n19067), .A(n19066), .ZN(n19069) );
  AOI21_X1 U22107 ( .B1(n19170), .B2(n19070), .A(n19069), .ZN(n19076) );
  INV_X1 U22108 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19183) );
  AOI21_X1 U22109 ( .B1(n19072), .B2(n19071), .A(n19183), .ZN(n19073) );
  AOI21_X1 U22110 ( .B1(n19248), .B2(n19074), .A(n19073), .ZN(n19075) );
  OAI211_X1 U22111 ( .C1(n19078), .C2(n19077), .A(n19076), .B(n19075), .ZN(
        P2_U2855) );
  AOI22_X1 U22112 ( .A1(n19084), .A2(BUF2_REG_31__SCAN_IN), .B1(n15992), .B2(
        n19087), .ZN(n19080) );
  AOI22_X1 U22113 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19104), .B1(n19083), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19079) );
  NAND2_X1 U22114 ( .A1(n19080), .A2(n19079), .ZN(P2_U2888) );
  AOI22_X1 U22115 ( .A1(n19082), .A2(n19081), .B1(n19104), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19091) );
  AOI22_X1 U22116 ( .A1(n19084), .A2(BUF2_REG_16__SCAN_IN), .B1(n19083), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19090) );
  NOR2_X1 U22117 ( .A1(n19085), .A2(n19107), .ZN(n19086) );
  AOI21_X1 U22118 ( .B1(n19088), .B2(n19087), .A(n19086), .ZN(n19089) );
  NAND3_X1 U22119 ( .A1(n19091), .A2(n19090), .A3(n19089), .ZN(P2_U2903) );
  INV_X1 U22120 ( .A(n19092), .ZN(n19095) );
  AOI22_X1 U22121 ( .A1(n19106), .A2(n19093), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19104), .ZN(n19094) );
  OAI21_X1 U22122 ( .B1(n19113), .B2(n19095), .A(n19094), .ZN(P2_U2905) );
  AOI22_X1 U22123 ( .A1(n19106), .A2(n19096), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19104), .ZN(n19097) );
  OAI21_X1 U22124 ( .B1(n19113), .B2(n19098), .A(n19097), .ZN(P2_U2909) );
  INV_X1 U22125 ( .A(n19113), .ZN(n19101) );
  AOI22_X1 U22126 ( .A1(n19101), .A2(n19100), .B1(n19106), .B2(n19099), .ZN(
        n19102) );
  OAI21_X1 U22127 ( .B1(n19103), .B2(n20860), .A(n19102), .ZN(P2_U2911) );
  AOI22_X1 U22128 ( .A1(n19106), .A2(n19105), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19104), .ZN(n19111) );
  OR3_X1 U22129 ( .A1(n19109), .A2(n19108), .A3(n19107), .ZN(n19110) );
  OAI211_X1 U22130 ( .C1(n19113), .C2(n19112), .A(n19111), .B(n19110), .ZN(
        P2_U2914) );
  NOR2_X1 U22131 ( .A1(n19150), .A2(n19114), .ZN(P2_U2920) );
  INV_X1 U22132 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n21031) );
  INV_X1 U22133 ( .A(n19115), .ZN(n19117) );
  AOI22_X1 U22134 ( .A1(n19143), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(n19117), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n19116) );
  OAI21_X1 U22135 ( .B1(n21031), .B2(n19877), .A(n19116), .ZN(P2_U2929) );
  AOI22_X1 U22136 ( .A1(n19117), .A2(P2_EAX_REG_16__SCAN_IN), .B1(
        P2_UWORD_REG_0__SCAN_IN), .B2(n19144), .ZN(n19118) );
  OAI21_X1 U22137 ( .B1(n21032), .B2(n19150), .A(n19118), .ZN(P2_U2935) );
  OAI222_X1 U22138 ( .A1(n19150), .A2(n20941), .B1(n19146), .B2(n19120), .C1(
        n19877), .C2(n19119), .ZN(P2_U2936) );
  AOI22_X1 U22139 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19148), .B1(n19147), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19121) );
  OAI21_X1 U22140 ( .B1(n20811), .B2(n19150), .A(n19121), .ZN(P2_U2937) );
  INV_X1 U22141 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n19122) );
  OAI222_X1 U22142 ( .A1(n19150), .A2(n20919), .B1(n19146), .B2(n19123), .C1(
        n19877), .C2(n19122), .ZN(P2_U2938) );
  AOI22_X1 U22143 ( .A1(n19144), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19124) );
  OAI21_X1 U22144 ( .B1(n19125), .B2(n19146), .A(n19124), .ZN(P2_U2939) );
  AOI22_X1 U22145 ( .A1(n19144), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19126) );
  OAI21_X1 U22146 ( .B1(n19127), .B2(n19146), .A(n19126), .ZN(P2_U2940) );
  AOI22_X1 U22147 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19148), .B1(n19143), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19128) );
  OAI21_X1 U22148 ( .B1(n20820), .B2(n19877), .A(n19128), .ZN(P2_U2941) );
  AOI22_X1 U22149 ( .A1(n19144), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19129) );
  OAI21_X1 U22150 ( .B1(n19130), .B2(n19146), .A(n19129), .ZN(P2_U2942) );
  AOI22_X1 U22151 ( .A1(n19144), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19131) );
  OAI21_X1 U22152 ( .B1(n20860), .B2(n19146), .A(n19131), .ZN(P2_U2943) );
  AOI22_X1 U22153 ( .A1(n19144), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19132) );
  OAI21_X1 U22154 ( .B1(n19133), .B2(n19146), .A(n19132), .ZN(P2_U2944) );
  INV_X1 U22155 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n20959) );
  OAI222_X1 U22156 ( .A1(n19877), .A2(n20959), .B1(n19146), .B2(n19135), .C1(
        n19150), .C2(n19134), .ZN(P2_U2945) );
  INV_X1 U22157 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19137) );
  AOI22_X1 U22158 ( .A1(n19144), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19136) );
  OAI21_X1 U22159 ( .B1(n19137), .B2(n19146), .A(n19136), .ZN(P2_U2946) );
  INV_X1 U22160 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19139) );
  AOI22_X1 U22161 ( .A1(n19144), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19138) );
  OAI21_X1 U22162 ( .B1(n19139), .B2(n19146), .A(n19138), .ZN(P2_U2947) );
  INV_X1 U22163 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n21041) );
  AOI22_X1 U22164 ( .A1(n19144), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19140) );
  OAI21_X1 U22165 ( .B1(n21041), .B2(n19146), .A(n19140), .ZN(P2_U2948) );
  INV_X1 U22166 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19142) );
  AOI22_X1 U22167 ( .A1(n19144), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19141) );
  OAI21_X1 U22168 ( .B1(n19142), .B2(n19146), .A(n19141), .ZN(P2_U2949) );
  AOI22_X1 U22169 ( .A1(n19144), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19143), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19145) );
  OAI21_X1 U22170 ( .B1(n13233), .B2(n19146), .A(n19145), .ZN(P2_U2950) );
  AOI22_X1 U22171 ( .A1(P2_EAX_REG_0__SCAN_IN), .A2(n19148), .B1(n19147), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n19149) );
  OAI21_X1 U22172 ( .B1(n20958), .B2(n19150), .A(n19149), .ZN(P2_U2951) );
  AOI22_X1 U22173 ( .A1(n19152), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n19151), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19154) );
  NAND2_X1 U22174 ( .A1(n19154), .A2(n19153), .ZN(P2_U2981) );
  AOI22_X1 U22175 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19169), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19029), .ZN(n19165) );
  INV_X1 U22176 ( .A(n19155), .ZN(n19156) );
  XNOR2_X1 U22177 ( .A(n19157), .B(n19156), .ZN(n19188) );
  INV_X1 U22178 ( .A(n19188), .ZN(n19162) );
  XNOR2_X1 U22179 ( .A(n19158), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19160) );
  XNOR2_X1 U22180 ( .A(n19160), .B(n19159), .ZN(n19197) );
  OAI22_X1 U22181 ( .A1(n19162), .A2(n19161), .B1(n19177), .B2(n19197), .ZN(
        n19163) );
  AOI21_X1 U22182 ( .B1(n19171), .B2(n19193), .A(n19163), .ZN(n19164) );
  OAI211_X1 U22183 ( .C1(n19167), .C2(n19166), .A(n19165), .B(n19164), .ZN(
        P2_U3010) );
  NOR2_X1 U22184 ( .A1(n19169), .A2(n19168), .ZN(n19184) );
  NAND2_X1 U22185 ( .A1(n19171), .A2(n19170), .ZN(n19181) );
  INV_X1 U22186 ( .A(n19172), .ZN(n19180) );
  INV_X1 U22187 ( .A(n19173), .ZN(n19174) );
  NAND2_X1 U22188 ( .A1(n19175), .A2(n19174), .ZN(n19179) );
  OR2_X1 U22189 ( .A1(n19177), .A2(n19176), .ZN(n19178) );
  AND4_X1 U22190 ( .A1(n19181), .A2(n19180), .A3(n19179), .A4(n19178), .ZN(
        n19182) );
  OAI21_X1 U22191 ( .B1(n19184), .B2(n19183), .A(n19182), .ZN(P2_U3014) );
  AOI22_X1 U22192 ( .A1(n19186), .A2(n19185), .B1(n19029), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n19200) );
  NAND2_X1 U22193 ( .A1(n19188), .A2(n19187), .ZN(n19195) );
  NOR2_X1 U22194 ( .A1(n19190), .A2(n19189), .ZN(n19191) );
  AOI21_X1 U22195 ( .B1(n19193), .B2(n19192), .A(n19191), .ZN(n19194) );
  OAI211_X1 U22196 ( .C1(n19197), .C2(n19196), .A(n19195), .B(n19194), .ZN(
        n19198) );
  INV_X1 U22197 ( .A(n19198), .ZN(n19199) );
  OAI211_X1 U22198 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n19201), .A(
        n19200), .B(n19199), .ZN(P2_U3042) );
  NAND2_X1 U22199 ( .A1(n13299), .A2(n19845), .ZN(n19309) );
  NOR2_X1 U22200 ( .A1(n19464), .A2(n19309), .ZN(n19242) );
  AOI22_X1 U22201 ( .A1(n19721), .A2(n19598), .B1(n19645), .B2(n19242), .ZN(
        n19211) );
  AOI21_X1 U22202 ( .B1(n19735), .B2(n19256), .A(n19882), .ZN(n19202) );
  INV_X1 U22203 ( .A(n19825), .ZN(n19835) );
  NOR2_X1 U22204 ( .A1(n19202), .A2(n19835), .ZN(n19207) );
  AOI21_X1 U22205 ( .B1(n19203), .B2(n19871), .A(n19825), .ZN(n19204) );
  AOI21_X1 U22206 ( .B1(n19207), .B2(n19205), .A(n19204), .ZN(n19206) );
  OAI21_X1 U22207 ( .B1(n19727), .B2(n19242), .A(n19207), .ZN(n19209) );
  OAI21_X1 U22208 ( .B1(n19203), .B2(n19242), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19208) );
  NAND2_X1 U22209 ( .A1(n19209), .A2(n19208), .ZN(n19244) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19245), .B1(
        n19658), .B2(n19244), .ZN(n19210) );
  OAI211_X1 U22211 ( .C1(n19601), .C2(n19256), .A(n19211), .B(n19210), .ZN(
        P2_U3048) );
  AOI22_X1 U22212 ( .A1(n19602), .A2(n19721), .B1(n19662), .B2(n19242), .ZN(
        n19213) );
  AOI22_X1 U22213 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19245), .B1(
        n19664), .B2(n19244), .ZN(n19212) );
  OAI211_X1 U22214 ( .C1(n19605), .C2(n19256), .A(n19213), .B(n19212), .ZN(
        P2_U3049) );
  AOI22_X1 U22215 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19235), .ZN(n19671) );
  AOI22_X1 U22216 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19235), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19234), .ZN(n19699) );
  NOR2_X2 U22217 ( .A1(n10689), .A2(n19240), .ZN(n19693) );
  AOI22_X1 U22218 ( .A1(n19721), .A2(n19668), .B1(n19693), .B2(n19242), .ZN(
        n19217) );
  INV_X1 U22219 ( .A(n19214), .ZN(n19215) );
  NOR2_X2 U22220 ( .A1(n19215), .A2(n19498), .ZN(n19694) );
  AOI22_X1 U22221 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19245), .B1(
        n19694), .B2(n19244), .ZN(n19216) );
  OAI211_X1 U22222 ( .C1(n19671), .C2(n19256), .A(n19217), .B(n19216), .ZN(
        P2_U3050) );
  AOI22_X1 U22223 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19235), .ZN(n19705) );
  AOI22_X1 U22224 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19235), .ZN(n19675) );
  NOR2_X2 U22225 ( .A1(n19218), .A2(n19240), .ZN(n19700) );
  AOI22_X1 U22226 ( .A1(n19702), .A2(n19721), .B1(n19700), .B2(n19242), .ZN(
        n19221) );
  NOR2_X2 U22227 ( .A1(n19219), .A2(n19498), .ZN(n19701) );
  AOI22_X1 U22228 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19245), .B1(
        n19701), .B2(n19244), .ZN(n19220) );
  OAI211_X1 U22229 ( .C1(n19705), .C2(n19256), .A(n19221), .B(n19220), .ZN(
        P2_U3051) );
  AOI22_X1 U22230 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19235), .ZN(n19613) );
  NOR2_X2 U22231 ( .A1(n19224), .A2(n19240), .ZN(n19706) );
  AOI22_X1 U22232 ( .A1(n19610), .A2(n19721), .B1(n19706), .B2(n19242), .ZN(
        n19227) );
  NOR2_X2 U22233 ( .A1(n19225), .A2(n19498), .ZN(n19707) );
  AOI22_X1 U22234 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19245), .B1(
        n19707), .B2(n19244), .ZN(n19226) );
  OAI211_X1 U22235 ( .C1(n19613), .C2(n19256), .A(n19227), .B(n19226), .ZN(
        P2_U3052) );
  AOI22_X1 U22236 ( .A1(n19679), .A2(n19721), .B1(n19712), .B2(n19242), .ZN(
        n19229) );
  AOI22_X1 U22237 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19245), .B1(
        n19713), .B2(n19244), .ZN(n19228) );
  OAI211_X1 U22238 ( .C1(n19682), .C2(n19256), .A(n19229), .B(n19228), .ZN(
        P2_U3053) );
  AOI22_X1 U22239 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19234), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19235), .ZN(n19619) );
  AOI22_X1 U22240 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19235), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19234), .ZN(n19725) );
  INV_X1 U22241 ( .A(n19725), .ZN(n19616) );
  NOR2_X2 U22242 ( .A1(n19230), .A2(n19240), .ZN(n19718) );
  AOI22_X1 U22243 ( .A1(n19616), .A2(n19721), .B1(n19718), .B2(n19242), .ZN(
        n19233) );
  NOR2_X2 U22244 ( .A1(n19231), .A2(n19498), .ZN(n19719) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19245), .B1(
        n19719), .B2(n19244), .ZN(n19232) );
  OAI211_X1 U22246 ( .C1(n19619), .C2(n19256), .A(n19233), .B(n19232), .ZN(
        P2_U3054) );
  AOI22_X1 U22247 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19235), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19234), .ZN(n19736) );
  NOR2_X2 U22248 ( .A1(n19241), .A2(n19240), .ZN(n19726) );
  AOI22_X1 U22249 ( .A1(n19730), .A2(n19721), .B1(n19726), .B2(n19242), .ZN(
        n19247) );
  NOR2_X2 U22250 ( .A1(n19243), .A2(n19498), .ZN(n19728) );
  AOI22_X1 U22251 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19245), .B1(
        n19728), .B2(n19244), .ZN(n19246) );
  OAI211_X1 U22252 ( .C1(n19736), .C2(n19256), .A(n19247), .B(n19246), .ZN(
        P2_U3055) );
  INV_X1 U22253 ( .A(n19309), .ZN(n19277) );
  NAND2_X1 U22254 ( .A1(n19277), .A2(n10893), .ZN(n19253) );
  NOR2_X1 U22255 ( .A1(n19861), .A2(n19253), .ZN(n19271) );
  OR3_X1 U22256 ( .A1(n19249), .A2(n19271), .A3(n19872), .ZN(n19254) );
  OAI21_X1 U22257 ( .B1(n19253), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19872), 
        .ZN(n19250) );
  AND2_X1 U22258 ( .A1(n19254), .A2(n19250), .ZN(n19272) );
  AOI22_X1 U22259 ( .A1(n19272), .A2(n19658), .B1(n19645), .B2(n19271), .ZN(
        n19258) );
  INV_X1 U22260 ( .A(n19463), .ZN(n19496) );
  NAND2_X1 U22261 ( .A1(n19251), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19439) );
  OR3_X1 U22262 ( .A1(n19496), .A2(n19439), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n19252) );
  OAI21_X1 U22263 ( .B1(n19858), .B2(n19253), .A(n19252), .ZN(n19255) );
  NAND3_X1 U22264 ( .A1(n19255), .A2(n19651), .A3(n19254), .ZN(n19274) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19598), .ZN(n19257) );
  OAI211_X1 U22266 ( .C1(n19601), .C2(n19308), .A(n19258), .B(n19257), .ZN(
        P2_U3056) );
  AOI22_X1 U22267 ( .A1(n19272), .A2(n19664), .B1(n19662), .B2(n19271), .ZN(
        n19260) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19602), .ZN(n19259) );
  OAI211_X1 U22269 ( .C1(n19605), .C2(n19308), .A(n19260), .B(n19259), .ZN(
        P2_U3057) );
  AOI22_X1 U22270 ( .A1(n19272), .A2(n19694), .B1(n19693), .B2(n19271), .ZN(
        n19262) );
  AOI22_X1 U22271 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19668), .ZN(n19261) );
  OAI211_X1 U22272 ( .C1(n19671), .C2(n19308), .A(n19262), .B(n19261), .ZN(
        P2_U3058) );
  AOI22_X1 U22273 ( .A1(n19272), .A2(n19701), .B1(n19700), .B2(n19271), .ZN(
        n19264) );
  AOI22_X1 U22274 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19702), .ZN(n19263) );
  OAI211_X1 U22275 ( .C1(n19705), .C2(n19308), .A(n19264), .B(n19263), .ZN(
        P2_U3059) );
  AOI22_X1 U22276 ( .A1(n19272), .A2(n19707), .B1(n19706), .B2(n19271), .ZN(
        n19266) );
  AOI22_X1 U22277 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19610), .ZN(n19265) );
  OAI211_X1 U22278 ( .C1(n19613), .C2(n19308), .A(n19266), .B(n19265), .ZN(
        P2_U3060) );
  AOI22_X1 U22279 ( .A1(n19272), .A2(n19713), .B1(n19712), .B2(n19271), .ZN(
        n19268) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19679), .ZN(n19267) );
  OAI211_X1 U22281 ( .C1(n19682), .C2(n19308), .A(n19268), .B(n19267), .ZN(
        P2_U3061) );
  AOI22_X1 U22282 ( .A1(n19272), .A2(n19719), .B1(n19718), .B2(n19271), .ZN(
        n19270) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19616), .ZN(n19269) );
  OAI211_X1 U22284 ( .C1(n19619), .C2(n19308), .A(n19270), .B(n19269), .ZN(
        P2_U3062) );
  AOI22_X1 U22285 ( .A1(n19272), .A2(n19728), .B1(n19726), .B2(n19271), .ZN(
        n19276) );
  AOI22_X1 U22286 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19274), .B1(
        n19273), .B2(n19730), .ZN(n19275) );
  OAI211_X1 U22287 ( .C1(n19736), .C2(n19308), .A(n19276), .B(n19275), .ZN(
        P2_U3063) );
  INV_X1 U22288 ( .A(n10941), .ZN(n19278) );
  NAND2_X1 U22289 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19277), .ZN(
        n19315) );
  NOR2_X1 U22290 ( .A1(n19315), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19303) );
  OAI21_X1 U22291 ( .B1(n19278), .B2(n19303), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19279) );
  OR2_X1 U22292 ( .A1(n19530), .A2(n19309), .ZN(n19284) );
  NAND2_X1 U22293 ( .A1(n19279), .A2(n19284), .ZN(n19304) );
  AOI22_X1 U22294 ( .A1(n19304), .A2(n19658), .B1(n19645), .B2(n19303), .ZN(
        n19290) );
  INV_X1 U22295 ( .A(n19303), .ZN(n19280) );
  OAI21_X1 U22296 ( .B1(n10941), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19280), 
        .ZN(n19287) );
  NAND2_X1 U22297 ( .A1(n19399), .A2(n19826), .ZN(n19337) );
  INV_X1 U22298 ( .A(n19308), .ZN(n19283) );
  OAI21_X1 U22299 ( .B1(n19329), .B2(n19283), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19285) );
  NAND2_X1 U22300 ( .A1(n19285), .A2(n19284), .ZN(n19286) );
  MUX2_X1 U22301 ( .A(n19287), .B(n19286), .S(n19825), .Z(n19288) );
  NAND2_X1 U22302 ( .A1(n19288), .A2(n19651), .ZN(n19305) );
  AOI22_X1 U22303 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19305), .B1(
        n19329), .B2(n19646), .ZN(n19289) );
  OAI211_X1 U22304 ( .C1(n19661), .C2(n19308), .A(n19290), .B(n19289), .ZN(
        P2_U3064) );
  AOI22_X1 U22305 ( .A1(n19304), .A2(n19664), .B1(n19662), .B2(n19303), .ZN(
        n19292) );
  AOI22_X1 U22306 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19305), .B1(
        n19329), .B2(n19663), .ZN(n19291) );
  OAI211_X1 U22307 ( .C1(n19667), .C2(n19308), .A(n19292), .B(n19291), .ZN(
        P2_U3065) );
  AOI22_X1 U22308 ( .A1(n19304), .A2(n19694), .B1(n19693), .B2(n19303), .ZN(
        n19294) );
  INV_X1 U22309 ( .A(n19671), .ZN(n19696) );
  AOI22_X1 U22310 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19305), .B1(
        n19329), .B2(n19696), .ZN(n19293) );
  OAI211_X1 U22311 ( .C1(n19699), .C2(n19308), .A(n19294), .B(n19293), .ZN(
        P2_U3066) );
  AOI22_X1 U22312 ( .A1(n19304), .A2(n19701), .B1(n19700), .B2(n19303), .ZN(
        n19296) );
  INV_X1 U22313 ( .A(n19705), .ZN(n19672) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19305), .B1(
        n19329), .B2(n19672), .ZN(n19295) );
  OAI211_X1 U22315 ( .C1(n19675), .C2(n19308), .A(n19296), .B(n19295), .ZN(
        P2_U3067) );
  AOI22_X1 U22316 ( .A1(n19304), .A2(n19707), .B1(n19706), .B2(n19303), .ZN(
        n19298) );
  INV_X1 U22317 ( .A(n19613), .ZN(n19708) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19305), .B1(
        n19329), .B2(n19708), .ZN(n19297) );
  OAI211_X1 U22319 ( .C1(n19711), .C2(n19308), .A(n19298), .B(n19297), .ZN(
        P2_U3068) );
  INV_X1 U22320 ( .A(n19679), .ZN(n19717) );
  AOI22_X1 U22321 ( .A1(n19304), .A2(n19713), .B1(n19712), .B2(n19303), .ZN(
        n19300) );
  AOI22_X1 U22322 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19305), .B1(
        n19329), .B2(n19714), .ZN(n19299) );
  OAI211_X1 U22323 ( .C1(n19717), .C2(n19308), .A(n19300), .B(n19299), .ZN(
        P2_U3069) );
  AOI22_X1 U22324 ( .A1(n19304), .A2(n19719), .B1(n19718), .B2(n19303), .ZN(
        n19302) );
  INV_X1 U22325 ( .A(n19619), .ZN(n19720) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19305), .B1(
        n19329), .B2(n19720), .ZN(n19301) );
  OAI211_X1 U22327 ( .C1(n19725), .C2(n19308), .A(n19302), .B(n19301), .ZN(
        P2_U3070) );
  AOI22_X1 U22328 ( .A1(n19304), .A2(n19728), .B1(n19726), .B2(n19303), .ZN(
        n19307) );
  INV_X1 U22329 ( .A(n19736), .ZN(n19686) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19305), .B1(
        n19329), .B2(n19686), .ZN(n19306) );
  OAI211_X1 U22331 ( .C1(n19692), .C2(n19308), .A(n19307), .B(n19306), .ZN(
        P2_U3071) );
  NOR2_X1 U22332 ( .A1(n19558), .A2(n19309), .ZN(n19332) );
  AOI22_X1 U22333 ( .A1(n19598), .A2(n19329), .B1(n19645), .B2(n19332), .ZN(
        n19318) );
  OAI21_X1 U22334 ( .B1(n19566), .B2(n19439), .A(n19825), .ZN(n19316) );
  INV_X1 U22335 ( .A(n19315), .ZN(n19310) );
  NOR2_X1 U22336 ( .A1(n19316), .A2(n19310), .ZN(n19311) );
  AOI211_X1 U22337 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n10950), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19311), .ZN(n19312) );
  OAI21_X1 U22338 ( .B1(n19332), .B2(n19312), .A(n19651), .ZN(n19334) );
  OAI21_X1 U22339 ( .B1(n19313), .B2(n19332), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19314) );
  OAI21_X1 U22340 ( .B1(n19316), .B2(n19315), .A(n19314), .ZN(n19333) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19334), .B1(
        n19658), .B2(n19333), .ZN(n19317) );
  OAI211_X1 U22342 ( .C1(n19601), .C2(n19342), .A(n19318), .B(n19317), .ZN(
        P2_U3072) );
  AOI22_X1 U22343 ( .A1(n19602), .A2(n19329), .B1(n19662), .B2(n19332), .ZN(
        n19320) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19334), .B1(
        n19664), .B2(n19333), .ZN(n19319) );
  OAI211_X1 U22345 ( .C1(n19605), .C2(n19342), .A(n19320), .B(n19319), .ZN(
        P2_U3073) );
  AOI22_X1 U22346 ( .A1(n19668), .A2(n19329), .B1(n19332), .B2(n19693), .ZN(
        n19322) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19334), .B1(
        n19694), .B2(n19333), .ZN(n19321) );
  OAI211_X1 U22348 ( .C1(n19671), .C2(n19342), .A(n19322), .B(n19321), .ZN(
        P2_U3074) );
  AOI22_X1 U22349 ( .A1(n19672), .A2(n19364), .B1(n19332), .B2(n19700), .ZN(
        n19324) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19334), .B1(
        n19701), .B2(n19333), .ZN(n19323) );
  OAI211_X1 U22351 ( .C1(n19675), .C2(n19337), .A(n19324), .B(n19323), .ZN(
        P2_U3075) );
  AOI22_X1 U22352 ( .A1(n19610), .A2(n19329), .B1(n19332), .B2(n19706), .ZN(
        n19326) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19334), .B1(
        n19707), .B2(n19333), .ZN(n19325) );
  OAI211_X1 U22354 ( .C1(n19613), .C2(n19342), .A(n19326), .B(n19325), .ZN(
        P2_U3076) );
  AOI22_X1 U22355 ( .A1(n19679), .A2(n19329), .B1(n19712), .B2(n19332), .ZN(
        n19328) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19334), .B1(
        n19713), .B2(n19333), .ZN(n19327) );
  OAI211_X1 U22357 ( .C1(n19682), .C2(n19342), .A(n19328), .B(n19327), .ZN(
        P2_U3077) );
  AOI22_X1 U22358 ( .A1(n19616), .A2(n19329), .B1(n19332), .B2(n19718), .ZN(
        n19331) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19334), .B1(
        n19719), .B2(n19333), .ZN(n19330) );
  OAI211_X1 U22360 ( .C1(n19619), .C2(n19342), .A(n19331), .B(n19330), .ZN(
        P2_U3078) );
  AOI22_X1 U22361 ( .A1(n19686), .A2(n19364), .B1(n19332), .B2(n19726), .ZN(
        n19336) );
  AOI22_X1 U22362 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19334), .B1(
        n19728), .B2(n19333), .ZN(n19335) );
  OAI211_X1 U22363 ( .C1(n19692), .C2(n19337), .A(n19336), .B(n19335), .ZN(
        P2_U3079) );
  NAND2_X1 U22364 ( .A1(n13299), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19435) );
  NOR2_X1 U22365 ( .A1(n19464), .A2(n19435), .ZN(n19362) );
  NOR3_X1 U22366 ( .A1(n19338), .A2(n19362), .A3(n19872), .ZN(n19343) );
  INV_X1 U22367 ( .A(n19402), .ZN(n19340) );
  NAND2_X1 U22368 ( .A1(n19340), .A2(n19339), .ZN(n19595) );
  NOR2_X1 U22369 ( .A1(n19595), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19347) );
  AOI21_X1 U22370 ( .B1(n19871), .B2(n19347), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19341) );
  NOR2_X1 U22371 ( .A1(n19343), .A2(n19341), .ZN(n19363) );
  AOI22_X1 U22372 ( .A1(n19363), .A2(n19658), .B1(n19645), .B2(n19362), .ZN(
        n19349) );
  AOI21_X1 U22373 ( .B1(n19342), .B2(n19398), .A(n19882), .ZN(n19346) );
  INV_X1 U22374 ( .A(n19362), .ZN(n19344) );
  AOI211_X1 U22375 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19344), .A(n19498), 
        .B(n19343), .ZN(n19345) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19365), .B1(
        n19364), .B2(n19598), .ZN(n19348) );
  OAI211_X1 U22377 ( .C1(n19601), .C2(n19398), .A(n19349), .B(n19348), .ZN(
        P2_U3080) );
  AOI22_X1 U22378 ( .A1(n19363), .A2(n19664), .B1(n19662), .B2(n19362), .ZN(
        n19351) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19365), .B1(
        n19364), .B2(n19602), .ZN(n19350) );
  OAI211_X1 U22380 ( .C1(n19605), .C2(n19398), .A(n19351), .B(n19350), .ZN(
        P2_U3081) );
  AOI22_X1 U22381 ( .A1(n19363), .A2(n19694), .B1(n19693), .B2(n19362), .ZN(
        n19353) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19365), .B1(
        n19364), .B2(n19668), .ZN(n19352) );
  OAI211_X1 U22383 ( .C1(n19671), .C2(n19398), .A(n19353), .B(n19352), .ZN(
        P2_U3082) );
  AOI22_X1 U22384 ( .A1(n19363), .A2(n19701), .B1(n19700), .B2(n19362), .ZN(
        n19355) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19365), .B1(
        n19364), .B2(n19702), .ZN(n19354) );
  OAI211_X1 U22386 ( .C1(n19705), .C2(n19398), .A(n19355), .B(n19354), .ZN(
        P2_U3083) );
  AOI22_X1 U22387 ( .A1(n19363), .A2(n19707), .B1(n19706), .B2(n19362), .ZN(
        n19357) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19365), .B1(
        n19364), .B2(n19610), .ZN(n19356) );
  OAI211_X1 U22389 ( .C1(n19613), .C2(n19398), .A(n19357), .B(n19356), .ZN(
        P2_U3084) );
  AOI22_X1 U22390 ( .A1(n19363), .A2(n19713), .B1(n19712), .B2(n19362), .ZN(
        n19359) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19365), .B1(
        n19364), .B2(n19679), .ZN(n19358) );
  OAI211_X1 U22392 ( .C1(n19682), .C2(n19398), .A(n19359), .B(n19358), .ZN(
        P2_U3085) );
  AOI22_X1 U22393 ( .A1(n19363), .A2(n19719), .B1(n19718), .B2(n19362), .ZN(
        n19361) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19365), .B1(
        n19364), .B2(n19616), .ZN(n19360) );
  OAI211_X1 U22395 ( .C1(n19619), .C2(n19398), .A(n19361), .B(n19360), .ZN(
        P2_U3086) );
  AOI22_X1 U22396 ( .A1(n19363), .A2(n19728), .B1(n19726), .B2(n19362), .ZN(
        n19367) );
  AOI22_X1 U22397 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19365), .B1(
        n19364), .B2(n19730), .ZN(n19366) );
  OAI211_X1 U22398 ( .C1(n19736), .C2(n19398), .A(n19367), .B(n19366), .ZN(
        P2_U3087) );
  INV_X1 U22399 ( .A(n19369), .ZN(n19370) );
  NOR2_X1 U22400 ( .A1(n19435), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19373) );
  INV_X1 U22401 ( .A(n19373), .ZN(n19376) );
  NOR2_X1 U22402 ( .A1(n19861), .A2(n19376), .ZN(n19393) );
  AOI22_X1 U22403 ( .A1(n19412), .A2(n19646), .B1(n19645), .B2(n19393), .ZN(
        n19379) );
  OAI21_X1 U22404 ( .B1(n19439), .B2(n19370), .A(n19825), .ZN(n19377) );
  INV_X1 U22405 ( .A(n19393), .ZN(n19371) );
  OAI211_X1 U22406 ( .C1(n10946), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19835), 
        .B(n19371), .ZN(n19372) );
  OAI211_X1 U22407 ( .C1(n19377), .C2(n19373), .A(n19651), .B(n19372), .ZN(
        n19395) );
  OAI21_X1 U22408 ( .B1(n19374), .B2(n19393), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19375) );
  OAI21_X1 U22409 ( .B1(n19377), .B2(n19376), .A(n19375), .ZN(n19394) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19395), .B1(
        n19658), .B2(n19394), .ZN(n19378) );
  OAI211_X1 U22411 ( .C1(n19661), .C2(n19398), .A(n19379), .B(n19378), .ZN(
        P2_U3088) );
  AOI22_X1 U22412 ( .A1(n19412), .A2(n19663), .B1(n19662), .B2(n19393), .ZN(
        n19381) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19395), .B1(
        n19664), .B2(n19394), .ZN(n19380) );
  OAI211_X1 U22414 ( .C1(n19667), .C2(n19398), .A(n19381), .B(n19380), .ZN(
        P2_U3089) );
  INV_X1 U22415 ( .A(n19398), .ZN(n19386) );
  AOI22_X1 U22416 ( .A1(n19668), .A2(n19386), .B1(n19693), .B2(n19393), .ZN(
        n19383) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19395), .B1(
        n19694), .B2(n19394), .ZN(n19382) );
  OAI211_X1 U22418 ( .C1(n19671), .C2(n19433), .A(n19383), .B(n19382), .ZN(
        P2_U3090) );
  AOI22_X1 U22419 ( .A1(n19412), .A2(n19672), .B1(n19393), .B2(n19700), .ZN(
        n19385) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19395), .B1(
        n19701), .B2(n19394), .ZN(n19384) );
  OAI211_X1 U22421 ( .C1(n19675), .C2(n19398), .A(n19385), .B(n19384), .ZN(
        P2_U3091) );
  AOI22_X1 U22422 ( .A1(n19610), .A2(n19386), .B1(n19393), .B2(n19706), .ZN(
        n19388) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19395), .B1(
        n19707), .B2(n19394), .ZN(n19387) );
  OAI211_X1 U22424 ( .C1(n19613), .C2(n19433), .A(n19388), .B(n19387), .ZN(
        P2_U3092) );
  AOI22_X1 U22425 ( .A1(n19412), .A2(n19714), .B1(n19712), .B2(n19393), .ZN(
        n19390) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19395), .B1(
        n19713), .B2(n19394), .ZN(n19389) );
  OAI211_X1 U22427 ( .C1(n19717), .C2(n19398), .A(n19390), .B(n19389), .ZN(
        P2_U3093) );
  AOI22_X1 U22428 ( .A1(n19412), .A2(n19720), .B1(n19393), .B2(n19718), .ZN(
        n19392) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19395), .B1(
        n19719), .B2(n19394), .ZN(n19391) );
  OAI211_X1 U22430 ( .C1(n19725), .C2(n19398), .A(n19392), .B(n19391), .ZN(
        P2_U3094) );
  AOI22_X1 U22431 ( .A1(n19412), .A2(n19686), .B1(n19393), .B2(n19726), .ZN(
        n19397) );
  AOI22_X1 U22432 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19395), .B1(
        n19728), .B2(n19394), .ZN(n19396) );
  OAI211_X1 U22433 ( .C1(n19692), .C2(n19398), .A(n19397), .B(n19396), .ZN(
        P2_U3095) );
  INV_X1 U22434 ( .A(n19399), .ZN(n19400) );
  OAI21_X1 U22435 ( .B1(n19412), .B2(n19459), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19404) );
  INV_X1 U22436 ( .A(n19435), .ZN(n19401) );
  NAND2_X1 U22437 ( .A1(n19402), .A2(n19401), .ZN(n19403) );
  NAND2_X1 U22438 ( .A1(n19404), .A2(n19403), .ZN(n19408) );
  NOR3_X2 U22439 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19644), .ZN(n19428) );
  NOR2_X1 U22440 ( .A1(n19825), .A2(n19428), .ZN(n19405) );
  OAI21_X1 U22441 ( .B1(n19409), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19405), 
        .ZN(n19406) );
  AND2_X1 U22442 ( .A1(n19406), .A2(n19651), .ZN(n19407) );
  INV_X1 U22443 ( .A(n19409), .ZN(n19410) );
  OAI21_X1 U22444 ( .B1(n19410), .B2(n19428), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19411) );
  OAI21_X1 U22445 ( .B1(n19435), .B2(n19530), .A(n19411), .ZN(n19429) );
  AOI22_X1 U22446 ( .A1(n19429), .A2(n19658), .B1(n19645), .B2(n19428), .ZN(
        n19414) );
  AOI22_X1 U22447 ( .A1(n19412), .A2(n19598), .B1(n19459), .B2(n19646), .ZN(
        n19413) );
  OAI211_X1 U22448 ( .C1(n19415), .C2(n11450), .A(n19414), .B(n19413), .ZN(
        P2_U3096) );
  AOI22_X1 U22449 ( .A1(n19429), .A2(n19664), .B1(n19662), .B2(n19428), .ZN(
        n19417) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19430), .B1(
        n19459), .B2(n19663), .ZN(n19416) );
  OAI211_X1 U22451 ( .C1(n19667), .C2(n19433), .A(n19417), .B(n19416), .ZN(
        P2_U3097) );
  AOI22_X1 U22452 ( .A1(n19429), .A2(n19694), .B1(n19693), .B2(n19428), .ZN(
        n19419) );
  AOI22_X1 U22453 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19430), .B1(
        n19459), .B2(n19696), .ZN(n19418) );
  OAI211_X1 U22454 ( .C1(n19699), .C2(n19433), .A(n19419), .B(n19418), .ZN(
        P2_U3098) );
  AOI22_X1 U22455 ( .A1(n19429), .A2(n19701), .B1(n19700), .B2(n19428), .ZN(
        n19421) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19430), .B1(
        n19459), .B2(n19672), .ZN(n19420) );
  OAI211_X1 U22457 ( .C1(n19675), .C2(n19433), .A(n19421), .B(n19420), .ZN(
        P2_U3099) );
  AOI22_X1 U22458 ( .A1(n19429), .A2(n19707), .B1(n19706), .B2(n19428), .ZN(
        n19423) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19430), .B1(
        n19459), .B2(n19708), .ZN(n19422) );
  OAI211_X1 U22460 ( .C1(n19711), .C2(n19433), .A(n19423), .B(n19422), .ZN(
        P2_U3100) );
  AOI22_X1 U22461 ( .A1(n19429), .A2(n19713), .B1(n19712), .B2(n19428), .ZN(
        n19425) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19430), .B1(
        n19459), .B2(n19714), .ZN(n19424) );
  OAI211_X1 U22463 ( .C1(n19717), .C2(n19433), .A(n19425), .B(n19424), .ZN(
        P2_U3101) );
  AOI22_X1 U22464 ( .A1(n19429), .A2(n19719), .B1(n19718), .B2(n19428), .ZN(
        n19427) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19430), .B1(
        n19459), .B2(n19720), .ZN(n19426) );
  OAI211_X1 U22466 ( .C1(n19725), .C2(n19433), .A(n19427), .B(n19426), .ZN(
        P2_U3102) );
  AOI22_X1 U22467 ( .A1(n19429), .A2(n19728), .B1(n19726), .B2(n19428), .ZN(
        n19432) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19430), .B1(
        n19459), .B2(n19686), .ZN(n19431) );
  OAI211_X1 U22469 ( .C1(n19692), .C2(n19433), .A(n19432), .B(n19431), .ZN(
        P2_U3103) );
  NOR2_X1 U22470 ( .A1(n19558), .A2(n19435), .ZN(n19467) );
  NOR2_X1 U22471 ( .A1(n19467), .A2(n19872), .ZN(n19436) );
  NAND2_X1 U22472 ( .A1(n10951), .A2(n19436), .ZN(n19440) );
  OR2_X1 U22473 ( .A1(n19644), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19442) );
  OAI21_X1 U22474 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19442), .A(n19872), 
        .ZN(n19437) );
  AND2_X1 U22475 ( .A1(n19440), .A2(n19437), .ZN(n19458) );
  AOI22_X1 U22476 ( .A1(n19458), .A2(n19658), .B1(n19645), .B2(n19467), .ZN(
        n19445) );
  OR2_X1 U22477 ( .A1(n19439), .A2(n19438), .ZN(n19836) );
  OAI211_X1 U22478 ( .C1(n19871), .C2(n19467), .A(n19440), .B(n19651), .ZN(
        n19441) );
  AOI21_X1 U22479 ( .B1(n19836), .B2(n19442), .A(n19441), .ZN(n19443) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19598), .ZN(n19444) );
  OAI211_X1 U22481 ( .C1(n19601), .C2(n19495), .A(n19445), .B(n19444), .ZN(
        P2_U3104) );
  AOI22_X1 U22482 ( .A1(n19458), .A2(n19664), .B1(n19662), .B2(n19467), .ZN(
        n19447) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19602), .ZN(n19446) );
  OAI211_X1 U22484 ( .C1(n19605), .C2(n19495), .A(n19447), .B(n19446), .ZN(
        P2_U3105) );
  AOI22_X1 U22485 ( .A1(n19458), .A2(n19694), .B1(n19467), .B2(n19693), .ZN(
        n19449) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19668), .ZN(n19448) );
  OAI211_X1 U22487 ( .C1(n19671), .C2(n19495), .A(n19449), .B(n19448), .ZN(
        P2_U3106) );
  AOI22_X1 U22488 ( .A1(n19458), .A2(n19701), .B1(n19467), .B2(n19700), .ZN(
        n19451) );
  AOI22_X1 U22489 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19702), .ZN(n19450) );
  OAI211_X1 U22490 ( .C1(n19705), .C2(n19495), .A(n19451), .B(n19450), .ZN(
        P2_U3107) );
  AOI22_X1 U22491 ( .A1(n19458), .A2(n19707), .B1(n19467), .B2(n19706), .ZN(
        n19453) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19610), .ZN(n19452) );
  OAI211_X1 U22493 ( .C1(n19613), .C2(n19495), .A(n19453), .B(n19452), .ZN(
        P2_U3108) );
  AOI22_X1 U22494 ( .A1(n19458), .A2(n19713), .B1(n19712), .B2(n19467), .ZN(
        n19455) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19679), .ZN(n19454) );
  OAI211_X1 U22496 ( .C1(n19682), .C2(n19495), .A(n19455), .B(n19454), .ZN(
        P2_U3109) );
  AOI22_X1 U22497 ( .A1(n19458), .A2(n19719), .B1(n19467), .B2(n19718), .ZN(
        n19457) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19616), .ZN(n19456) );
  OAI211_X1 U22499 ( .C1(n19619), .C2(n19495), .A(n19457), .B(n19456), .ZN(
        P2_U3110) );
  AOI22_X1 U22500 ( .A1(n19458), .A2(n19728), .B1(n19467), .B2(n19726), .ZN(
        n19462) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19460), .B1(
        n19459), .B2(n19730), .ZN(n19461) );
  OAI211_X1 U22502 ( .C1(n19736), .C2(n19495), .A(n19462), .B(n19461), .ZN(
        P2_U3111) );
  NAND2_X1 U22503 ( .A1(n19527), .A2(n19463), .ZN(n19516) );
  NAND2_X1 U22504 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19845), .ZN(
        n19557) );
  NOR2_X1 U22505 ( .A1(n19464), .A2(n19557), .ZN(n19490) );
  AOI22_X1 U22506 ( .A1(n19646), .A2(n19522), .B1(n19645), .B2(n19490), .ZN(
        n19477) );
  INV_X1 U22507 ( .A(n19495), .ZN(n19465) );
  OAI21_X1 U22508 ( .B1(n19522), .B2(n19465), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19466) );
  NAND2_X1 U22509 ( .A1(n19466), .A2(n19825), .ZN(n19475) );
  NOR2_X1 U22510 ( .A1(n19490), .A2(n19467), .ZN(n19473) );
  INV_X1 U22511 ( .A(n19473), .ZN(n19471) );
  INV_X1 U22512 ( .A(n19490), .ZN(n19468) );
  OAI211_X1 U22513 ( .C1(n19469), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19835), 
        .B(n19468), .ZN(n19470) );
  OAI211_X1 U22514 ( .C1(n19475), .C2(n19471), .A(n19651), .B(n19470), .ZN(
        n19492) );
  OAI21_X1 U22515 ( .B1(n19472), .B2(n19490), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19474) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19492), .B1(
        n19658), .B2(n19491), .ZN(n19476) );
  OAI211_X1 U22517 ( .C1(n19661), .C2(n19495), .A(n19477), .B(n19476), .ZN(
        P2_U3112) );
  AOI22_X1 U22518 ( .A1(n19663), .A2(n19522), .B1(n19662), .B2(n19490), .ZN(
        n19479) );
  AOI22_X1 U22519 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19492), .B1(
        n19664), .B2(n19491), .ZN(n19478) );
  OAI211_X1 U22520 ( .C1(n19667), .C2(n19495), .A(n19479), .B(n19478), .ZN(
        P2_U3113) );
  AOI22_X1 U22521 ( .A1(n19696), .A2(n19522), .B1(n19693), .B2(n19490), .ZN(
        n19481) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19492), .B1(
        n19694), .B2(n19491), .ZN(n19480) );
  OAI211_X1 U22523 ( .C1(n19699), .C2(n19495), .A(n19481), .B(n19480), .ZN(
        P2_U3114) );
  AOI22_X1 U22524 ( .A1(n19672), .A2(n19522), .B1(n19700), .B2(n19490), .ZN(
        n19483) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19492), .B1(
        n19701), .B2(n19491), .ZN(n19482) );
  OAI211_X1 U22526 ( .C1(n19675), .C2(n19495), .A(n19483), .B(n19482), .ZN(
        P2_U3115) );
  AOI22_X1 U22527 ( .A1(n19708), .A2(n19522), .B1(n19706), .B2(n19490), .ZN(
        n19485) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19492), .B1(
        n19707), .B2(n19491), .ZN(n19484) );
  OAI211_X1 U22529 ( .C1(n19711), .C2(n19495), .A(n19485), .B(n19484), .ZN(
        P2_U3116) );
  AOI22_X1 U22530 ( .A1(n19714), .A2(n19522), .B1(n19712), .B2(n19490), .ZN(
        n19487) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19492), .B1(
        n19713), .B2(n19491), .ZN(n19486) );
  OAI211_X1 U22532 ( .C1(n19717), .C2(n19495), .A(n19487), .B(n19486), .ZN(
        P2_U3117) );
  AOI22_X1 U22533 ( .A1(n19720), .A2(n19522), .B1(n19718), .B2(n19490), .ZN(
        n19489) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19492), .B1(
        n19719), .B2(n19491), .ZN(n19488) );
  OAI211_X1 U22535 ( .C1(n19725), .C2(n19495), .A(n19489), .B(n19488), .ZN(
        P2_U3118) );
  AOI22_X1 U22536 ( .A1(n19686), .A2(n19522), .B1(n19726), .B2(n19490), .ZN(
        n19494) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19492), .B1(
        n19728), .B2(n19491), .ZN(n19493) );
  OAI211_X1 U22538 ( .C1(n19692), .C2(n19495), .A(n19494), .B(n19493), .ZN(
        P2_U3119) );
  NOR3_X2 U22539 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19861), .A3(
        n19557), .ZN(n19521) );
  AOI22_X1 U22540 ( .A1(n19522), .A2(n19598), .B1(n19645), .B2(n19521), .ZN(
        n19507) );
  INV_X1 U22541 ( .A(n19561), .ZN(n19497) );
  OAI21_X1 U22542 ( .B1(n19497), .B2(n19496), .A(n19825), .ZN(n19505) );
  NOR2_X1 U22543 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19557), .ZN(
        n19501) );
  OAI21_X1 U22544 ( .B1(n19502), .B2(n19872), .A(n19871), .ZN(n19499) );
  INV_X1 U22545 ( .A(n19521), .ZN(n19531) );
  AOI21_X1 U22546 ( .B1(n19499), .B2(n19531), .A(n19498), .ZN(n19500) );
  OAI21_X1 U22547 ( .B1(n19505), .B2(n19501), .A(n19500), .ZN(n19524) );
  INV_X1 U22548 ( .A(n19501), .ZN(n19504) );
  OAI21_X1 U22549 ( .B1(n19502), .B2(n19521), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19503) );
  OAI21_X1 U22550 ( .B1(n19505), .B2(n19504), .A(n19503), .ZN(n19523) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19524), .B1(
        n19658), .B2(n19523), .ZN(n19506) );
  OAI211_X1 U22552 ( .C1(n19601), .C2(n19532), .A(n19507), .B(n19506), .ZN(
        P2_U3120) );
  AOI22_X1 U22553 ( .A1(n19602), .A2(n19522), .B1(n19662), .B2(n19521), .ZN(
        n19509) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19524), .B1(
        n19664), .B2(n19523), .ZN(n19508) );
  OAI211_X1 U22555 ( .C1(n19605), .C2(n19532), .A(n19509), .B(n19508), .ZN(
        P2_U3121) );
  AOI22_X1 U22556 ( .A1(n19696), .A2(n19552), .B1(n19693), .B2(n19521), .ZN(
        n19511) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19524), .B1(
        n19694), .B2(n19523), .ZN(n19510) );
  OAI211_X1 U22558 ( .C1(n19699), .C2(n19516), .A(n19511), .B(n19510), .ZN(
        P2_U3122) );
  AOI22_X1 U22559 ( .A1(n19702), .A2(n19522), .B1(n19700), .B2(n19521), .ZN(
        n19513) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19524), .B1(
        n19701), .B2(n19523), .ZN(n19512) );
  OAI211_X1 U22561 ( .C1(n19705), .C2(n19532), .A(n19513), .B(n19512), .ZN(
        P2_U3123) );
  AOI22_X1 U22562 ( .A1(n19708), .A2(n19552), .B1(n19706), .B2(n19521), .ZN(
        n19515) );
  AOI22_X1 U22563 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19524), .B1(
        n19707), .B2(n19523), .ZN(n19514) );
  OAI211_X1 U22564 ( .C1(n19711), .C2(n19516), .A(n19515), .B(n19514), .ZN(
        P2_U3124) );
  AOI22_X1 U22565 ( .A1(n19679), .A2(n19522), .B1(n19712), .B2(n19521), .ZN(
        n19518) );
  AOI22_X1 U22566 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19524), .B1(
        n19713), .B2(n19523), .ZN(n19517) );
  OAI211_X1 U22567 ( .C1(n19682), .C2(n19532), .A(n19518), .B(n19517), .ZN(
        P2_U3125) );
  AOI22_X1 U22568 ( .A1(n19616), .A2(n19522), .B1(n19718), .B2(n19521), .ZN(
        n19520) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19524), .B1(
        n19719), .B2(n19523), .ZN(n19519) );
  OAI211_X1 U22570 ( .C1(n19619), .C2(n19532), .A(n19520), .B(n19519), .ZN(
        P2_U3126) );
  AOI22_X1 U22571 ( .A1(n19730), .A2(n19522), .B1(n19726), .B2(n19521), .ZN(
        n19526) );
  AOI22_X1 U22572 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19524), .B1(
        n19728), .B2(n19523), .ZN(n19525) );
  OAI211_X1 U22573 ( .C1(n19736), .C2(n19532), .A(n19526), .B(n19525), .ZN(
        P2_U3127) );
  NOR3_X2 U22574 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10893), .A3(
        n19557), .ZN(n19550) );
  OAI21_X1 U22575 ( .B1(n19528), .B2(n19550), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19529) );
  OAI21_X1 U22576 ( .B1(n19557), .B2(n19530), .A(n19529), .ZN(n19551) );
  AOI22_X1 U22577 ( .A1(n19551), .A2(n19658), .B1(n19645), .B2(n19550), .ZN(
        n19537) );
  OAI221_X1 U22578 ( .B1(n19587), .B2(n19882), .C1(n19532), .C2(n19882), .A(
        n19531), .ZN(n19533) );
  OAI211_X1 U22579 ( .C1(n19528), .C2(n19872), .A(n19533), .B(n19871), .ZN(
        n19534) );
  INV_X1 U22580 ( .A(n19534), .ZN(n19535) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19598), .ZN(n19536) );
  OAI211_X1 U22582 ( .C1(n19601), .C2(n19587), .A(n19537), .B(n19536), .ZN(
        P2_U3128) );
  AOI22_X1 U22583 ( .A1(n19551), .A2(n19664), .B1(n19662), .B2(n19550), .ZN(
        n19539) );
  AOI22_X1 U22584 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19602), .ZN(n19538) );
  OAI211_X1 U22585 ( .C1(n19605), .C2(n19587), .A(n19539), .B(n19538), .ZN(
        P2_U3129) );
  AOI22_X1 U22586 ( .A1(n19551), .A2(n19694), .B1(n19693), .B2(n19550), .ZN(
        n19541) );
  AOI22_X1 U22587 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19668), .ZN(n19540) );
  OAI211_X1 U22588 ( .C1(n19671), .C2(n19587), .A(n19541), .B(n19540), .ZN(
        P2_U3130) );
  AOI22_X1 U22589 ( .A1(n19551), .A2(n19701), .B1(n19700), .B2(n19550), .ZN(
        n19543) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19702), .ZN(n19542) );
  OAI211_X1 U22591 ( .C1(n19705), .C2(n19587), .A(n19543), .B(n19542), .ZN(
        P2_U3131) );
  AOI22_X1 U22592 ( .A1(n19551), .A2(n19707), .B1(n19706), .B2(n19550), .ZN(
        n19545) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19610), .ZN(n19544) );
  OAI211_X1 U22594 ( .C1(n19613), .C2(n19587), .A(n19545), .B(n19544), .ZN(
        P2_U3132) );
  AOI22_X1 U22595 ( .A1(n19551), .A2(n19713), .B1(n19712), .B2(n19550), .ZN(
        n19547) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19679), .ZN(n19546) );
  OAI211_X1 U22597 ( .C1(n19682), .C2(n19587), .A(n19547), .B(n19546), .ZN(
        P2_U3133) );
  AOI22_X1 U22598 ( .A1(n19551), .A2(n19719), .B1(n19718), .B2(n19550), .ZN(
        n19549) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19616), .ZN(n19548) );
  OAI211_X1 U22600 ( .C1(n19619), .C2(n19587), .A(n19549), .B(n19548), .ZN(
        P2_U3134) );
  AOI22_X1 U22601 ( .A1(n19551), .A2(n19728), .B1(n19726), .B2(n19550), .ZN(
        n19555) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19553), .B1(
        n19552), .B2(n19730), .ZN(n19554) );
  OAI211_X1 U22603 ( .C1(n19736), .C2(n19587), .A(n19555), .B(n19554), .ZN(
        P2_U3135) );
  INV_X1 U22604 ( .A(n19557), .ZN(n19556) );
  NAND2_X1 U22605 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19556), .ZN(
        n19563) );
  OR2_X1 U22606 ( .A1(n19563), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19560) );
  NOR2_X1 U22607 ( .A1(n19558), .A2(n19557), .ZN(n19582) );
  NOR3_X1 U22608 ( .A1(n19559), .A2(n19582), .A3(n19872), .ZN(n19562) );
  AOI21_X1 U22609 ( .B1(n19872), .B2(n19560), .A(n19562), .ZN(n19583) );
  AOI22_X1 U22610 ( .A1(n19583), .A2(n19658), .B1(n19645), .B2(n19582), .ZN(
        n19569) );
  NAND2_X1 U22611 ( .A1(n19561), .A2(n19826), .ZN(n19564) );
  AOI21_X1 U22612 ( .B1(n19564), .B2(n19563), .A(n19562), .ZN(n19565) );
  OAI211_X1 U22613 ( .C1(n19582), .C2(n19871), .A(n19565), .B(n19651), .ZN(
        n19584) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19584), .B1(
        n19622), .B2(n19646), .ZN(n19568) );
  OAI211_X1 U22615 ( .C1(n19661), .C2(n19587), .A(n19569), .B(n19568), .ZN(
        P2_U3136) );
  AOI22_X1 U22616 ( .A1(n19583), .A2(n19664), .B1(n19662), .B2(n19582), .ZN(
        n19571) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19584), .B1(
        n19622), .B2(n19663), .ZN(n19570) );
  OAI211_X1 U22618 ( .C1(n19667), .C2(n19587), .A(n19571), .B(n19570), .ZN(
        P2_U3137) );
  AOI22_X1 U22619 ( .A1(n19583), .A2(n19694), .B1(n19693), .B2(n19582), .ZN(
        n19573) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19584), .B1(
        n19622), .B2(n19696), .ZN(n19572) );
  OAI211_X1 U22621 ( .C1(n19699), .C2(n19587), .A(n19573), .B(n19572), .ZN(
        P2_U3138) );
  AOI22_X1 U22622 ( .A1(n19583), .A2(n19701), .B1(n19700), .B2(n19582), .ZN(
        n19575) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19584), .B1(
        n19622), .B2(n19672), .ZN(n19574) );
  OAI211_X1 U22624 ( .C1(n19675), .C2(n19587), .A(n19575), .B(n19574), .ZN(
        P2_U3139) );
  AOI22_X1 U22625 ( .A1(n19583), .A2(n19707), .B1(n19706), .B2(n19582), .ZN(
        n19577) );
  AOI22_X1 U22626 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19584), .B1(
        n19622), .B2(n19708), .ZN(n19576) );
  OAI211_X1 U22627 ( .C1(n19711), .C2(n19587), .A(n19577), .B(n19576), .ZN(
        P2_U3140) );
  AOI22_X1 U22628 ( .A1(n19583), .A2(n19713), .B1(n19712), .B2(n19582), .ZN(
        n19579) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19584), .B1(
        n19622), .B2(n19714), .ZN(n19578) );
  OAI211_X1 U22630 ( .C1(n19717), .C2(n19587), .A(n19579), .B(n19578), .ZN(
        P2_U3141) );
  AOI22_X1 U22631 ( .A1(n19583), .A2(n19719), .B1(n19718), .B2(n19582), .ZN(
        n19581) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19584), .B1(
        n19622), .B2(n19720), .ZN(n19580) );
  OAI211_X1 U22633 ( .C1(n19725), .C2(n19587), .A(n19581), .B(n19580), .ZN(
        P2_U3142) );
  AOI22_X1 U22634 ( .A1(n19583), .A2(n19728), .B1(n19726), .B2(n19582), .ZN(
        n19586) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19584), .B1(
        n19622), .B2(n19686), .ZN(n19585) );
  OAI211_X1 U22636 ( .C1(n19692), .C2(n19587), .A(n19586), .B(n19585), .ZN(
        P2_U3143) );
  INV_X1 U22637 ( .A(n19588), .ZN(n19592) );
  NOR2_X1 U22638 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19589), .ZN(
        n19620) );
  OAI21_X1 U22639 ( .B1(n19590), .B2(n19620), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19591) );
  OAI21_X1 U22640 ( .B1(n19592), .B2(n19595), .A(n19591), .ZN(n19621) );
  AOI22_X1 U22641 ( .A1(n19621), .A2(n19658), .B1(n19645), .B2(n19620), .ZN(
        n19600) );
  AOI21_X1 U22642 ( .B1(n19593), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19597) );
  OAI21_X1 U22643 ( .B1(n19630), .B2(n19622), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19594) );
  OAI21_X1 U22644 ( .B1(n19595), .B2(n13299), .A(n19594), .ZN(n19596) );
  OAI211_X1 U22645 ( .C1(n19620), .C2(n19597), .A(n19596), .B(n19651), .ZN(
        n19623) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19598), .ZN(n19599) );
  OAI211_X1 U22647 ( .C1(n19601), .C2(n19643), .A(n19600), .B(n19599), .ZN(
        P2_U3144) );
  AOI22_X1 U22648 ( .A1(n19621), .A2(n19664), .B1(n19662), .B2(n19620), .ZN(
        n19604) );
  AOI22_X1 U22649 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19602), .ZN(n19603) );
  OAI211_X1 U22650 ( .C1(n19605), .C2(n19643), .A(n19604), .B(n19603), .ZN(
        P2_U3145) );
  AOI22_X1 U22651 ( .A1(n19621), .A2(n19694), .B1(n19693), .B2(n19620), .ZN(
        n19607) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19668), .ZN(n19606) );
  OAI211_X1 U22653 ( .C1(n19671), .C2(n19643), .A(n19607), .B(n19606), .ZN(
        P2_U3146) );
  AOI22_X1 U22654 ( .A1(n19621), .A2(n19701), .B1(n19700), .B2(n19620), .ZN(
        n19609) );
  AOI22_X1 U22655 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19702), .ZN(n19608) );
  OAI211_X1 U22656 ( .C1(n19705), .C2(n19643), .A(n19609), .B(n19608), .ZN(
        P2_U3147) );
  AOI22_X1 U22657 ( .A1(n19621), .A2(n19707), .B1(n19706), .B2(n19620), .ZN(
        n19612) );
  AOI22_X1 U22658 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19610), .ZN(n19611) );
  OAI211_X1 U22659 ( .C1(n19613), .C2(n19643), .A(n19612), .B(n19611), .ZN(
        P2_U3148) );
  AOI22_X1 U22660 ( .A1(n19621), .A2(n19713), .B1(n19712), .B2(n19620), .ZN(
        n19615) );
  AOI22_X1 U22661 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19679), .ZN(n19614) );
  OAI211_X1 U22662 ( .C1(n19682), .C2(n19643), .A(n19615), .B(n19614), .ZN(
        P2_U3149) );
  AOI22_X1 U22663 ( .A1(n19621), .A2(n19719), .B1(n19718), .B2(n19620), .ZN(
        n19618) );
  AOI22_X1 U22664 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19616), .ZN(n19617) );
  OAI211_X1 U22665 ( .C1(n19619), .C2(n19643), .A(n19618), .B(n19617), .ZN(
        P2_U3150) );
  AOI22_X1 U22666 ( .A1(n19621), .A2(n19728), .B1(n19726), .B2(n19620), .ZN(
        n19625) );
  AOI22_X1 U22667 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19623), .B1(
        n19622), .B2(n19730), .ZN(n19624) );
  OAI211_X1 U22668 ( .C1(n19736), .C2(n19643), .A(n19625), .B(n19624), .ZN(
        P2_U3151) );
  AOI22_X1 U22669 ( .A1(n19639), .A2(n19664), .B1(n19648), .B2(n19662), .ZN(
        n19627) );
  INV_X1 U22670 ( .A(n19634), .ZN(n19640) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19640), .B1(
        n19678), .B2(n19663), .ZN(n19626) );
  OAI211_X1 U22672 ( .C1(n19667), .C2(n19643), .A(n19627), .B(n19626), .ZN(
        P2_U3153) );
  INV_X1 U22673 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20970) );
  AOI22_X1 U22674 ( .A1(n19639), .A2(n19694), .B1(n19648), .B2(n19693), .ZN(
        n19629) );
  AOI22_X1 U22675 ( .A1(n19630), .A2(n19668), .B1(n19678), .B2(n19696), .ZN(
        n19628) );
  OAI211_X1 U22676 ( .C1(n19634), .C2(n20970), .A(n19629), .B(n19628), .ZN(
        P2_U3154) );
  AOI22_X1 U22677 ( .A1(n19639), .A2(n19701), .B1(n19648), .B2(n19700), .ZN(
        n19632) );
  AOI22_X1 U22678 ( .A1(n19630), .A2(n19702), .B1(n19678), .B2(n19672), .ZN(
        n19631) );
  OAI211_X1 U22679 ( .C1(n19634), .C2(n19633), .A(n19632), .B(n19631), .ZN(
        P2_U3155) );
  AOI22_X1 U22680 ( .A1(n19639), .A2(n19707), .B1(n19648), .B2(n19706), .ZN(
        n19636) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19640), .B1(
        n19678), .B2(n19708), .ZN(n19635) );
  OAI211_X1 U22682 ( .C1(n19711), .C2(n19643), .A(n19636), .B(n19635), .ZN(
        P2_U3156) );
  AOI22_X1 U22683 ( .A1(n19639), .A2(n19719), .B1(n19648), .B2(n19718), .ZN(
        n19638) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19640), .B1(
        n19678), .B2(n19720), .ZN(n19637) );
  OAI211_X1 U22685 ( .C1(n19725), .C2(n19643), .A(n19638), .B(n19637), .ZN(
        P2_U3158) );
  AOI22_X1 U22686 ( .A1(n19639), .A2(n19728), .B1(n19648), .B2(n19726), .ZN(
        n19642) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19640), .B1(
        n19678), .B2(n19686), .ZN(n19641) );
  OAI211_X1 U22688 ( .C1(n19692), .C2(n19643), .A(n19642), .B(n19641), .ZN(
        P2_U3159) );
  NOR3_X2 U22689 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13299), .A3(
        n19644), .ZN(n19685) );
  AOI22_X1 U22690 ( .A1(n19646), .A2(n19731), .B1(n19645), .B2(n19685), .ZN(
        n19660) );
  OAI21_X1 U22691 ( .B1(n19731), .B2(n19678), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19647) );
  NAND2_X1 U22692 ( .A1(n19647), .A2(n19825), .ZN(n19657) );
  NOR2_X1 U22693 ( .A1(n19685), .A2(n19648), .ZN(n19656) );
  INV_X1 U22694 ( .A(n19656), .ZN(n19652) );
  INV_X1 U22695 ( .A(n19685), .ZN(n19649) );
  OAI211_X1 U22696 ( .C1(n19653), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19835), 
        .B(n19649), .ZN(n19650) );
  OAI211_X1 U22697 ( .C1(n19657), .C2(n19652), .A(n19651), .B(n19650), .ZN(
        n19688) );
  INV_X1 U22698 ( .A(n19653), .ZN(n19654) );
  OAI21_X1 U22699 ( .B1(n19654), .B2(n19685), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19655) );
  AOI22_X1 U22700 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19688), .B1(
        n19658), .B2(n19687), .ZN(n19659) );
  OAI211_X1 U22701 ( .C1(n19661), .C2(n19691), .A(n19660), .B(n19659), .ZN(
        P2_U3160) );
  AOI22_X1 U22702 ( .A1(n19663), .A2(n19731), .B1(n19662), .B2(n19685), .ZN(
        n19666) );
  AOI22_X1 U22703 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19688), .B1(
        n19664), .B2(n19687), .ZN(n19665) );
  OAI211_X1 U22704 ( .C1(n19667), .C2(n19691), .A(n19666), .B(n19665), .ZN(
        P2_U3161) );
  AOI22_X1 U22705 ( .A1(n19678), .A2(n19668), .B1(n19693), .B2(n19685), .ZN(
        n19670) );
  AOI22_X1 U22706 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19688), .B1(
        n19694), .B2(n19687), .ZN(n19669) );
  OAI211_X1 U22707 ( .C1(n19671), .C2(n19724), .A(n19670), .B(n19669), .ZN(
        P2_U3162) );
  AOI22_X1 U22708 ( .A1(n19672), .A2(n19731), .B1(n19700), .B2(n19685), .ZN(
        n19674) );
  AOI22_X1 U22709 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19688), .B1(
        n19701), .B2(n19687), .ZN(n19673) );
  OAI211_X1 U22710 ( .C1(n19675), .C2(n19691), .A(n19674), .B(n19673), .ZN(
        P2_U3163) );
  AOI22_X1 U22711 ( .A1(n19708), .A2(n19731), .B1(n19706), .B2(n19685), .ZN(
        n19677) );
  AOI22_X1 U22712 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19688), .B1(
        n19707), .B2(n19687), .ZN(n19676) );
  OAI211_X1 U22713 ( .C1(n19711), .C2(n19691), .A(n19677), .B(n19676), .ZN(
        P2_U3164) );
  AOI22_X1 U22714 ( .A1(n19679), .A2(n19678), .B1(n19712), .B2(n19685), .ZN(
        n19681) );
  AOI22_X1 U22715 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19688), .B1(
        n19713), .B2(n19687), .ZN(n19680) );
  OAI211_X1 U22716 ( .C1(n19682), .C2(n19724), .A(n19681), .B(n19680), .ZN(
        P2_U3165) );
  AOI22_X1 U22717 ( .A1(n19720), .A2(n19731), .B1(n19718), .B2(n19685), .ZN(
        n19684) );
  AOI22_X1 U22718 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19688), .B1(
        n19719), .B2(n19687), .ZN(n19683) );
  OAI211_X1 U22719 ( .C1(n19725), .C2(n19691), .A(n19684), .B(n19683), .ZN(
        P2_U3166) );
  AOI22_X1 U22720 ( .A1(n19686), .A2(n19731), .B1(n19726), .B2(n19685), .ZN(
        n19690) );
  AOI22_X1 U22721 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19688), .B1(
        n19728), .B2(n19687), .ZN(n19689) );
  OAI211_X1 U22722 ( .C1(n19692), .C2(n19691), .A(n19690), .B(n19689), .ZN(
        P2_U3167) );
  AOI22_X1 U22723 ( .A1(n19729), .A2(n19694), .B1(n19727), .B2(n19693), .ZN(
        n19698) );
  INV_X1 U22724 ( .A(n19695), .ZN(n19732) );
  AOI22_X1 U22725 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19732), .B1(
        n19721), .B2(n19696), .ZN(n19697) );
  OAI211_X1 U22726 ( .C1(n19699), .C2(n19724), .A(n19698), .B(n19697), .ZN(
        P2_U3170) );
  AOI22_X1 U22727 ( .A1(n19729), .A2(n19701), .B1(n19727), .B2(n19700), .ZN(
        n19704) );
  AOI22_X1 U22728 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19732), .B1(
        n19731), .B2(n19702), .ZN(n19703) );
  OAI211_X1 U22729 ( .C1(n19705), .C2(n19735), .A(n19704), .B(n19703), .ZN(
        P2_U3171) );
  AOI22_X1 U22730 ( .A1(n19729), .A2(n19707), .B1(n19727), .B2(n19706), .ZN(
        n19710) );
  AOI22_X1 U22731 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19732), .B1(
        n19721), .B2(n19708), .ZN(n19709) );
  OAI211_X1 U22732 ( .C1(n19711), .C2(n19724), .A(n19710), .B(n19709), .ZN(
        P2_U3172) );
  AOI22_X1 U22733 ( .A1(n19729), .A2(n19713), .B1(n19727), .B2(n19712), .ZN(
        n19716) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19732), .B1(
        n19721), .B2(n19714), .ZN(n19715) );
  OAI211_X1 U22735 ( .C1(n19717), .C2(n19724), .A(n19716), .B(n19715), .ZN(
        P2_U3173) );
  AOI22_X1 U22736 ( .A1(n19729), .A2(n19719), .B1(n19727), .B2(n19718), .ZN(
        n19723) );
  AOI22_X1 U22737 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19732), .B1(
        n19721), .B2(n19720), .ZN(n19722) );
  OAI211_X1 U22738 ( .C1(n19725), .C2(n19724), .A(n19723), .B(n19722), .ZN(
        P2_U3174) );
  AOI22_X1 U22739 ( .A1(n19729), .A2(n19728), .B1(n19727), .B2(n19726), .ZN(
        n19734) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19732), .B1(
        n19731), .B2(n19730), .ZN(n19733) );
  OAI211_X1 U22741 ( .C1(n19736), .C2(n19735), .A(n19734), .B(n19733), .ZN(
        P2_U3175) );
  NOR2_X1 U22742 ( .A1(n19876), .A2(n19884), .ZN(n19738) );
  AOI21_X1 U22743 ( .B1(n19827), .B2(n19738), .A(n19737), .ZN(n19742) );
  NOR2_X1 U22744 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19884), .ZN(n19739) );
  OAI211_X1 U22745 ( .C1(n19743), .C2(n19739), .A(n19876), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19740) );
  OAI211_X1 U22746 ( .C1(n19743), .C2(n19742), .A(n19741), .B(n19740), .ZN(
        P2_U3177) );
  AND2_X1 U22747 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19744), .ZN(
        P2_U3179) );
  AND2_X1 U22748 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19744), .ZN(
        P2_U3180) );
  AND2_X1 U22749 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19744), .ZN(
        P2_U3181) );
  AND2_X1 U22750 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19744), .ZN(
        P2_U3182) );
  AND2_X1 U22751 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19744), .ZN(
        P2_U3183) );
  AND2_X1 U22752 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19744), .ZN(
        P2_U3184) );
  AND2_X1 U22753 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19744), .ZN(
        P2_U3185) );
  AND2_X1 U22754 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19744), .ZN(
        P2_U3186) );
  INV_X1 U22755 ( .A(P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20983) );
  NOR2_X1 U22756 ( .A1(n20983), .A2(n19824), .ZN(P2_U3187) );
  AND2_X1 U22757 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19744), .ZN(
        P2_U3188) );
  AND2_X1 U22758 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19744), .ZN(
        P2_U3189) );
  AND2_X1 U22759 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19744), .ZN(
        P2_U3190) );
  AND2_X1 U22760 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19744), .ZN(
        P2_U3191) );
  AND2_X1 U22761 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19744), .ZN(
        P2_U3192) );
  AND2_X1 U22762 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19744), .ZN(
        P2_U3193) );
  AND2_X1 U22763 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19744), .ZN(
        P2_U3194) );
  AND2_X1 U22764 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19744), .ZN(
        P2_U3195) );
  AND2_X1 U22765 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19744), .ZN(
        P2_U3196) );
  AND2_X1 U22766 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19744), .ZN(
        P2_U3197) );
  NOR2_X1 U22767 ( .A1(n20842), .A2(n19824), .ZN(P2_U3198) );
  AND2_X1 U22768 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19744), .ZN(
        P2_U3199) );
  NOR2_X1 U22769 ( .A1(n20864), .A2(n19824), .ZN(P2_U3200) );
  AND2_X1 U22770 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19744), .ZN(P2_U3201) );
  AND2_X1 U22771 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19744), .ZN(P2_U3202) );
  AND2_X1 U22772 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19744), .ZN(P2_U3203) );
  AND2_X1 U22773 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19744), .ZN(P2_U3204) );
  INV_X1 U22774 ( .A(P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n21053) );
  NOR2_X1 U22775 ( .A1(n21053), .A2(n19824), .ZN(P2_U3205) );
  AND2_X1 U22776 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19744), .ZN(P2_U3206) );
  AND2_X1 U22777 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19744), .ZN(P2_U3207) );
  AND2_X1 U22778 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19744), .ZN(P2_U3208) );
  NOR2_X1 U22779 ( .A1(n19880), .A2(n19745), .ZN(n19756) );
  INV_X1 U22780 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19889) );
  OR3_X1 U22781 ( .A1(n19756), .A2(n19889), .A3(n19746), .ZN(n19748) );
  AOI211_X1 U22782 ( .C1(n20717), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19757), .B(n19805), .ZN(n19747) );
  NOR2_X1 U22783 ( .A1(n20722), .A2(n19750), .ZN(n19762) );
  AOI211_X1 U22784 ( .C1(n21048), .C2(n19748), .A(n19747), .B(n19762), .ZN(
        n19749) );
  INV_X1 U22785 ( .A(n19749), .ZN(P2_U3209) );
  AOI21_X1 U22786 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20717), .A(n21048), 
        .ZN(n19754) );
  NOR2_X1 U22787 ( .A1(n19889), .A2(n19754), .ZN(n19751) );
  AOI21_X1 U22788 ( .B1(n19751), .B2(n19750), .A(n19756), .ZN(n19752) );
  OAI211_X1 U22789 ( .C1(n20717), .C2(n19753), .A(n19752), .B(n19881), .ZN(
        P2_U3210) );
  AOI21_X1 U22790 ( .B1(n19755), .B2(n19876), .A(n19754), .ZN(n19761) );
  AOI22_X1 U22791 ( .A1(n19889), .A2(n19757), .B1(n20722), .B2(n19756), .ZN(
        n19758) );
  INV_X1 U22792 ( .A(n19758), .ZN(n19759) );
  OAI211_X1 U22793 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19759), .ZN(n19760) );
  OAI21_X1 U22794 ( .B1(n19762), .B2(n19761), .A(n19760), .ZN(P2_U3211) );
  NAND2_X1 U22795 ( .A1(n19805), .A2(n21048), .ZN(n19815) );
  OAI222_X1 U22796 ( .A1(n19813), .A2(n19763), .B1(n20972), .B2(n19805), .C1(
        n20918), .C2(n19812), .ZN(P2_U3212) );
  OAI222_X1 U22797 ( .A1(n19813), .A2(n20918), .B1(n19764), .B2(n19805), .C1(
        n19766), .C2(n19812), .ZN(P2_U3213) );
  OAI222_X1 U22798 ( .A1(n19813), .A2(n19766), .B1(n19765), .B2(n19805), .C1(
        n11438), .C2(n19812), .ZN(P2_U3214) );
  OAI222_X1 U22799 ( .A1(n19812), .A2(n13782), .B1(n19767), .B2(n19805), .C1(
        n11438), .C2(n19813), .ZN(P2_U3215) );
  OAI222_X1 U22800 ( .A1(n19815), .A2(n19769), .B1(n19768), .B2(n19805), .C1(
        n13782), .C2(n19813), .ZN(P2_U3216) );
  OAI222_X1 U22801 ( .A1(n19815), .A2(n19771), .B1(n19770), .B2(n19805), .C1(
        n19769), .C2(n19813), .ZN(P2_U3217) );
  OAI222_X1 U22802 ( .A1(n19815), .A2(n11468), .B1(n19772), .B2(n19805), .C1(
        n19771), .C2(n19813), .ZN(P2_U3218) );
  OAI222_X1 U22803 ( .A1(n19815), .A2(n19773), .B1(n20982), .B2(n19805), .C1(
        n11468), .C2(n19813), .ZN(P2_U3219) );
  OAI222_X1 U22804 ( .A1(n19815), .A2(n11508), .B1(n19774), .B2(n19805), .C1(
        n19773), .C2(n19813), .ZN(P2_U3220) );
  INV_X1 U22805 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19776) );
  OAI222_X1 U22806 ( .A1(n19812), .A2(n19776), .B1(n19775), .B2(n19805), .C1(
        n11508), .C2(n19813), .ZN(P2_U3221) );
  OAI222_X1 U22807 ( .A1(n19812), .A2(n11549), .B1(n19777), .B2(n19805), .C1(
        n19776), .C2(n19813), .ZN(P2_U3222) );
  OAI222_X1 U22808 ( .A1(n19812), .A2(n19779), .B1(n19778), .B2(n19805), .C1(
        n11549), .C2(n19813), .ZN(P2_U3223) );
  OAI222_X1 U22809 ( .A1(n19812), .A2(n19781), .B1(n19780), .B2(n19805), .C1(
        n19779), .C2(n19813), .ZN(P2_U3224) );
  OAI222_X1 U22810 ( .A1(n19812), .A2(n19783), .B1(n19782), .B2(n19805), .C1(
        n19781), .C2(n19813), .ZN(P2_U3225) );
  OAI222_X1 U22811 ( .A1(n19812), .A2(n19785), .B1(n19784), .B2(n19805), .C1(
        n19783), .C2(n19813), .ZN(P2_U3226) );
  OAI222_X1 U22812 ( .A1(n19815), .A2(n19787), .B1(n19786), .B2(n19805), .C1(
        n19785), .C2(n19813), .ZN(P2_U3227) );
  OAI222_X1 U22813 ( .A1(n19815), .A2(n19789), .B1(n19788), .B2(n19805), .C1(
        n19787), .C2(n19813), .ZN(P2_U3228) );
  OAI222_X1 U22814 ( .A1(n19815), .A2(n19790), .B1(n20832), .B2(n19805), .C1(
        n19789), .C2(n19813), .ZN(P2_U3229) );
  OAI222_X1 U22815 ( .A1(n19815), .A2(n19792), .B1(n19791), .B2(n19805), .C1(
        n19790), .C2(n19813), .ZN(P2_U3230) );
  OAI222_X1 U22816 ( .A1(n19815), .A2(n19794), .B1(n19793), .B2(n19805), .C1(
        n19792), .C2(n19813), .ZN(P2_U3231) );
  OAI222_X1 U22817 ( .A1(n19815), .A2(n19796), .B1(n19795), .B2(n19805), .C1(
        n19794), .C2(n19813), .ZN(P2_U3232) );
  OAI222_X1 U22818 ( .A1(n19812), .A2(n19798), .B1(n19797), .B2(n19805), .C1(
        n19796), .C2(n19813), .ZN(P2_U3233) );
  OAI222_X1 U22819 ( .A1(n19812), .A2(n19800), .B1(n19799), .B2(n19805), .C1(
        n19798), .C2(n19813), .ZN(P2_U3234) );
  OAI222_X1 U22820 ( .A1(n19812), .A2(n19802), .B1(n19801), .B2(n19805), .C1(
        n19800), .C2(n19813), .ZN(P2_U3235) );
  INV_X1 U22821 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19804) );
  OAI222_X1 U22822 ( .A1(n19812), .A2(n19804), .B1(n19803), .B2(n19805), .C1(
        n19802), .C2(n19813), .ZN(P2_U3236) );
  OAI222_X1 U22823 ( .A1(n19812), .A2(n19807), .B1(n21007), .B2(n19805), .C1(
        n19804), .C2(n19813), .ZN(P2_U3237) );
  INV_X1 U22824 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19808) );
  OAI222_X1 U22825 ( .A1(n19813), .A2(n19807), .B1(n19806), .B2(n19805), .C1(
        n19808), .C2(n19812), .ZN(P2_U3238) );
  INV_X1 U22826 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19810) );
  OAI222_X1 U22827 ( .A1(n19812), .A2(n19810), .B1(n19809), .B2(n19805), .C1(
        n19808), .C2(n19813), .ZN(P2_U3239) );
  OAI222_X1 U22828 ( .A1(n19812), .A2(n20975), .B1(n19811), .B2(n19805), .C1(
        n19810), .C2(n19813), .ZN(P2_U3240) );
  OAI222_X1 U22829 ( .A1(n19815), .A2(n19814), .B1(n20956), .B2(n19805), .C1(
        n20975), .C2(n19813), .ZN(P2_U3241) );
  INV_X1 U22830 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19816) );
  AOI22_X1 U22831 ( .A1(n19805), .A2(n19817), .B1(n19816), .B2(n19891), .ZN(
        P2_U3585) );
  MUX2_X1 U22832 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19805), .Z(P2_U3586) );
  AOI22_X1 U22833 ( .A1(n19805), .A2(n19818), .B1(n20987), .B2(n19891), .ZN(
        P2_U3587) );
  INV_X1 U22834 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19819) );
  AOI22_X1 U22835 ( .A1(n19805), .A2(n19820), .B1(n19819), .B2(n19891), .ZN(
        P2_U3588) );
  OAI21_X1 U22836 ( .B1(n19824), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19822), 
        .ZN(n19821) );
  INV_X1 U22837 ( .A(n19821), .ZN(P2_U3591) );
  OAI21_X1 U22838 ( .B1(n19824), .B2(n19823), .A(n19822), .ZN(P2_U3592) );
  AND2_X1 U22839 ( .A1(n19825), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19850) );
  NAND2_X1 U22840 ( .A1(n19826), .A2(n19850), .ZN(n19839) );
  INV_X1 U22841 ( .A(n19827), .ZN(n19828) );
  NAND3_X1 U22842 ( .A1(n19848), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19828), 
        .ZN(n19829) );
  NAND2_X1 U22843 ( .A1(n19829), .A2(n19846), .ZN(n19840) );
  NAND2_X1 U22844 ( .A1(n19839), .A2(n19840), .ZN(n19831) );
  NAND2_X1 U22845 ( .A1(n19831), .A2(n19830), .ZN(n19834) );
  NAND2_X1 U22846 ( .A1(n19832), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19833) );
  OAI211_X1 U22847 ( .C1(n19836), .C2(n19835), .A(n19834), .B(n19833), .ZN(
        n19837) );
  INV_X1 U22848 ( .A(n19837), .ZN(n19838) );
  AOI22_X1 U22849 ( .A1(n19854), .A2(n13299), .B1(n19838), .B2(n19862), .ZN(
        P2_U3602) );
  OAI21_X1 U22850 ( .B1(n19841), .B2(n19840), .A(n19839), .ZN(n19842) );
  AOI21_X1 U22851 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19843), .A(n19842), 
        .ZN(n19844) );
  AOI22_X1 U22852 ( .A1(n19854), .A2(n19845), .B1(n19844), .B2(n19862), .ZN(
        P2_U3603) );
  INV_X1 U22853 ( .A(n19846), .ZN(n19856) );
  NOR2_X1 U22854 ( .A1(n19856), .A2(n19847), .ZN(n19849) );
  MUX2_X1 U22855 ( .A(n19850), .B(n19849), .S(n19848), .Z(n19851) );
  AOI21_X1 U22856 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19852), .A(n19851), 
        .ZN(n19853) );
  AOI22_X1 U22857 ( .A1(n19854), .A2(n10893), .B1(n19853), .B2(n19862), .ZN(
        P2_U3604) );
  OAI22_X1 U22858 ( .A1(n19857), .A2(n19856), .B1(n19872), .B2(n19855), .ZN(
        n19859) );
  OAI21_X1 U22859 ( .B1(n19859), .B2(n19858), .A(n19862), .ZN(n19860) );
  OAI21_X1 U22860 ( .B1(n19862), .B2(n19861), .A(n19860), .ZN(P2_U3605) );
  AOI22_X1 U22861 ( .A1(n19805), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19863), 
        .B2(n19891), .ZN(P2_U3608) );
  AOI22_X1 U22862 ( .A1(n19866), .A2(n19865), .B1(n10702), .B2(n19864), .ZN(
        n19868) );
  OAI21_X1 U22863 ( .B1(n19868), .B2(n11195), .A(n19867), .ZN(n19870) );
  MUX2_X1 U22864 ( .A(P2_MORE_REG_SCAN_IN), .B(n19870), .S(n19869), .Z(
        P2_U3609) );
  OAI21_X1 U22865 ( .B1(n19873), .B2(n19872), .A(n19871), .ZN(n19874) );
  OAI211_X1 U22866 ( .C1(n19877), .C2(n19876), .A(n19875), .B(n19874), .ZN(
        n19890) );
  NOR2_X1 U22867 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19878), .ZN(n19879) );
  AOI21_X1 U22868 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19880), .A(n19879), 
        .ZN(n19887) );
  AOI21_X1 U22869 ( .B1(n19883), .B2(n19882), .A(n19881), .ZN(n19885) );
  NOR3_X1 U22870 ( .A1(n11376), .A2(n19885), .A3(n19884), .ZN(n19886) );
  OAI21_X1 U22871 ( .B1(n19887), .B2(n19886), .A(n19890), .ZN(n19888) );
  OAI21_X1 U22872 ( .B1(n19890), .B2(n19889), .A(n19888), .ZN(P2_U3610) );
  OAI22_X1 U22873 ( .A1(n19891), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19805), .ZN(n19892) );
  INV_X1 U22874 ( .A(n19892), .ZN(P2_U3611) );
  AOI21_X1 U22875 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20877), .A(n12961), 
        .ZN(n20718) );
  INV_X1 U22876 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n19893) );
  INV_X2 U22877 ( .A(n20794), .ZN(n20809) );
  NOR2_X1 U22878 ( .A1(n20718), .A2(n20809), .ZN(n20786) );
  OAI21_X1 U22879 ( .B1(n20913), .B2(n12961), .A(n20783), .ZN(P1_U2802) );
  OAI21_X1 U22880 ( .B1(n19895), .B2(n19894), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19896) );
  OAI21_X1 U22881 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19897), .A(n19896), 
        .ZN(P1_U2803) );
  NOR2_X1 U22882 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19899) );
  OAI21_X1 U22883 ( .B1(n19899), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20794), .ZN(
        n19898) );
  OAI21_X1 U22884 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20794), .A(n19898), 
        .ZN(P1_U2804) );
  OAI21_X1 U22885 ( .B1(BS16), .B2(n19899), .A(n20786), .ZN(n20784) );
  OAI21_X1 U22886 ( .B1(n20786), .B2(n21079), .A(n20784), .ZN(P1_U2805) );
  OAI21_X1 U22887 ( .B1(n19902), .B2(n19901), .A(n19900), .ZN(P1_U2806) );
  NOR4_X1 U22888 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19906) );
  NOR4_X1 U22889 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19905) );
  NOR4_X1 U22890 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_27__SCAN_IN), .A3(P1_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_29__SCAN_IN), .ZN(n19904) );
  NOR4_X1 U22891 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19903) );
  NAND4_X1 U22892 ( .A1(n19906), .A2(n19905), .A3(n19904), .A4(n19903), .ZN(
        n19912) );
  NOR4_X1 U22893 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19910) );
  AOI211_X1 U22894 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_6__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19909) );
  NOR4_X1 U22895 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19908) );
  NOR4_X1 U22896 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19907) );
  NAND4_X1 U22897 ( .A1(n19910), .A2(n19909), .A3(n19908), .A4(n19907), .ZN(
        n19911) );
  NOR2_X1 U22898 ( .A1(n19912), .A2(n19911), .ZN(n20793) );
  INV_X1 U22899 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20781) );
  NOR3_X1 U22900 ( .A1(P1_DATAWIDTH_REG_0__SCAN_IN), .A2(
        P1_REIP_REG_0__SCAN_IN), .A3(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19914)
         );
  OAI21_X1 U22901 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19914), .A(n20793), .ZN(
        n19913) );
  OAI21_X1 U22902 ( .B1(n20793), .B2(n20781), .A(n19913), .ZN(P1_U2807) );
  INV_X1 U22903 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20788) );
  INV_X1 U22904 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20785) );
  AOI21_X1 U22905 ( .B1(n20788), .B2(n20785), .A(n19914), .ZN(n19915) );
  INV_X1 U22906 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20778) );
  INV_X1 U22907 ( .A(n20793), .ZN(n20790) );
  AOI22_X1 U22908 ( .A1(n20793), .A2(n19915), .B1(n20778), .B2(n20790), .ZN(
        P1_U2808) );
  AOI22_X1 U22909 ( .A1(n20003), .A2(n19949), .B1(n19982), .B2(n19916), .ZN(
        n19924) );
  INV_X1 U22910 ( .A(n20000), .ZN(n19917) );
  AOI22_X1 U22911 ( .A1(n19994), .A2(P1_EBX_REG_9__SCAN_IN), .B1(n19991), .B2(
        n19917), .ZN(n19918) );
  OAI211_X1 U22912 ( .C1(n19993), .C2(n19919), .A(n19918), .B(n19954), .ZN(
        n19920) );
  AOI221_X1 U22913 ( .B1(n19922), .B2(P1_REIP_REG_9__SCAN_IN), .C1(n19921), 
        .C2(n20946), .A(n19920), .ZN(n19923) );
  NAND2_X1 U22914 ( .A1(n19924), .A2(n19923), .ZN(P1_U2831) );
  NAND2_X1 U22915 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19925) );
  AND2_X1 U22916 ( .A1(n19989), .A2(n19925), .ZN(n19926) );
  OR2_X1 U22917 ( .A1(n19970), .A2(n19926), .ZN(n19940) );
  NAND2_X1 U22918 ( .A1(n19940), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n19935) );
  INV_X1 U22919 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20735) );
  NAND3_X1 U22920 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n20735), .ZN(n19932) );
  NAND2_X1 U22921 ( .A1(n19975), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n19927) );
  NAND2_X1 U22922 ( .A1(n19927), .A2(n19954), .ZN(n19928) );
  AOI21_X1 U22923 ( .B1(n19994), .B2(P1_EBX_REG_7__SCAN_IN), .A(n19928), .ZN(
        n19931) );
  NAND2_X1 U22924 ( .A1(n19991), .A2(n19929), .ZN(n19930) );
  OAI211_X1 U22925 ( .C1(n19932), .C2(n19959), .A(n19931), .B(n19930), .ZN(
        n19933) );
  INV_X1 U22926 ( .A(n19933), .ZN(n19934) );
  NAND2_X1 U22927 ( .A1(n19935), .A2(n19934), .ZN(n19936) );
  AOI21_X1 U22928 ( .B1(n19937), .B2(n19949), .A(n19936), .ZN(n19938) );
  OAI21_X1 U22929 ( .B1(n19939), .B2(n19992), .A(n19938), .ZN(P1_U2833) );
  INV_X1 U22930 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20731) );
  NOR3_X1 U22931 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20731), .A3(n19959), .ZN(
        n19948) );
  INV_X1 U22932 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19945) );
  AOI22_X1 U22933 ( .A1(n19991), .A2(n19941), .B1(P1_REIP_REG_6__SCAN_IN), 
        .B2(n19940), .ZN(n19942) );
  NAND2_X1 U22934 ( .A1(n19954), .A2(n19942), .ZN(n19943) );
  AOI21_X1 U22935 ( .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n19975), .A(
        n19943), .ZN(n19944) );
  OAI21_X1 U22936 ( .B1(n19946), .B2(n19945), .A(n19944), .ZN(n19947) );
  NOR2_X1 U22937 ( .A1(n19948), .A2(n19947), .ZN(n19952) );
  NAND2_X1 U22938 ( .A1(n19950), .A2(n19949), .ZN(n19951) );
  OAI211_X1 U22939 ( .C1(n19992), .C2(n19953), .A(n19952), .B(n19951), .ZN(
        P1_U2834) );
  INV_X1 U22940 ( .A(n19999), .ZN(n19971) );
  INV_X1 U22941 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19956) );
  AOI22_X1 U22942 ( .A1(n19991), .A2(n20006), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n19970), .ZN(n19955) );
  OAI211_X1 U22943 ( .C1(n19993), .C2(n19956), .A(n19955), .B(n19954), .ZN(
        n19957) );
  AOI21_X1 U22944 ( .B1(n19994), .B2(P1_EBX_REG_5__SCAN_IN), .A(n19957), .ZN(
        n19958) );
  OAI21_X1 U22945 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n19959), .A(n19958), .ZN(
        n19960) );
  AOI21_X1 U22946 ( .B1(n20009), .B2(n19971), .A(n19960), .ZN(n19961) );
  OAI21_X1 U22947 ( .B1(n19962), .B2(n19992), .A(n19961), .ZN(P1_U2835) );
  AOI22_X1 U22948 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19975), .B1(
        n19963), .B2(n19995), .ZN(n19969) );
  AOI21_X1 U22949 ( .B1(n19994), .B2(P1_EBX_REG_4__SCAN_IN), .A(n19964), .ZN(
        n19968) );
  NAND2_X1 U22950 ( .A1(n19991), .A2(n20088), .ZN(n19967) );
  INV_X1 U22951 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20729) );
  NAND3_X1 U22952 ( .A1(n19985), .A2(n20729), .A3(n19965), .ZN(n19966) );
  AND4_X1 U22953 ( .A1(n19969), .A2(n19968), .A3(n19967), .A4(n19966), .ZN(
        n19973) );
  AOI22_X1 U22954 ( .A1(n20080), .A2(n19971), .B1(n19970), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n19972) );
  OAI211_X1 U22955 ( .C1(n20084), .C2(n19992), .A(n19973), .B(n19972), .ZN(
        P1_U2836) );
  INV_X1 U22956 ( .A(n19995), .ZN(n19977) );
  AOI22_X1 U22957 ( .A1(n19975), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n19974), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n19976) );
  OAI21_X1 U22958 ( .B1(n19977), .B2(n20520), .A(n19976), .ZN(n19978) );
  AOI21_X1 U22959 ( .B1(n19994), .B2(P1_EBX_REG_2__SCAN_IN), .A(n19978), .ZN(
        n19979) );
  OAI21_X1 U22960 ( .B1(n19980), .B2(n19999), .A(n19979), .ZN(n19981) );
  AOI21_X1 U22961 ( .B1(n19983), .B2(n19982), .A(n19981), .ZN(n19987) );
  OAI211_X1 U22962 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), 
        .A(n19985), .B(n19984), .ZN(n19986) );
  OAI211_X1 U22963 ( .C1(n20108), .C2(n19988), .A(n19987), .B(n19986), .ZN(
        P1_U2838) );
  AOI22_X1 U22964 ( .A1(n19991), .A2(n19990), .B1(P1_REIP_REG_0__SCAN_IN), 
        .B2(n19989), .ZN(n19998) );
  NAND2_X1 U22965 ( .A1(n19993), .A2(n19992), .ZN(n19996) );
  AOI222_X1 U22966 ( .A1(n19996), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19995), .B2(n20256), .C1(P1_EBX_REG_0__SCAN_IN), .C2(n19994), .ZN(
        n19997) );
  OAI211_X1 U22967 ( .C1(n19999), .C2(n20017), .A(n19998), .B(n19997), .ZN(
        P1_U2840) );
  NOR2_X1 U22968 ( .A1(n20001), .A2(n20000), .ZN(n20002) );
  AOI21_X1 U22969 ( .B1(n20003), .B2(n20008), .A(n20002), .ZN(n20004) );
  OAI21_X1 U22970 ( .B1(n20012), .B2(n20005), .A(n20004), .ZN(P1_U2863) );
  AOI22_X1 U22971 ( .A1(n20009), .A2(n20008), .B1(n20007), .B2(n20006), .ZN(
        n20010) );
  OAI21_X1 U22972 ( .B1(n20012), .B2(n20011), .A(n20010), .ZN(P1_U2867) );
  INV_X1 U22973 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20052) );
  INV_X1 U22974 ( .A(n20141), .ZN(n20013) );
  OAI222_X1 U22975 ( .A1(n20017), .A2(n20016), .B1(n20052), .B2(n20015), .C1(
        n20014), .C2(n20013), .ZN(P1_U2904) );
  INV_X1 U22976 ( .A(n20018), .ZN(n20020) );
  AOI22_X1 U22977 ( .A1(n20020), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n20049), .ZN(n20019) );
  OAI21_X1 U22978 ( .B1(n20976), .B2(n20800), .A(n20019), .ZN(P1_U2910) );
  AOI22_X1 U22979 ( .A1(n20020), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n20049), .ZN(n20021) );
  OAI21_X1 U22980 ( .B1(n21024), .B2(n20800), .A(n20021), .ZN(P1_U2912) );
  OAI222_X1 U22981 ( .A1(n20800), .A2(n20023), .B1(n20051), .B2(n20022), .C1(
        n20953), .C2(n20044), .ZN(P1_U2921) );
  INV_X1 U22982 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20025) );
  AOI22_X1 U22983 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20024) );
  OAI21_X1 U22984 ( .B1(n20025), .B2(n20051), .A(n20024), .ZN(P1_U2922) );
  INV_X1 U22985 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20027) );
  AOI22_X1 U22986 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20026) );
  OAI21_X1 U22987 ( .B1(n20027), .B2(n20051), .A(n20026), .ZN(P1_U2923) );
  INV_X1 U22988 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20029) );
  AOI22_X1 U22989 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20028) );
  OAI21_X1 U22990 ( .B1(n20029), .B2(n20051), .A(n20028), .ZN(P1_U2924) );
  AOI22_X1 U22991 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20030) );
  OAI21_X1 U22992 ( .B1(n20896), .B2(n20051), .A(n20030), .ZN(P1_U2925) );
  INV_X1 U22993 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20032) );
  AOI22_X1 U22994 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20031) );
  OAI21_X1 U22995 ( .B1(n20032), .B2(n20051), .A(n20031), .ZN(P1_U2926) );
  INV_X1 U22996 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20034) );
  AOI22_X1 U22997 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20033) );
  OAI21_X1 U22998 ( .B1(n20034), .B2(n20051), .A(n20033), .ZN(P1_U2927) );
  AOI22_X1 U22999 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20035) );
  OAI21_X1 U23000 ( .B1(n20036), .B2(n20051), .A(n20035), .ZN(P1_U2928) );
  AOI22_X1 U23001 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20037) );
  OAI21_X1 U23002 ( .B1(n12112), .B2(n20051), .A(n20037), .ZN(P1_U2929) );
  AOI22_X1 U23003 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20038) );
  OAI21_X1 U23004 ( .B1(n20039), .B2(n20051), .A(n20038), .ZN(P1_U2930) );
  AOI22_X1 U23005 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20040) );
  OAI21_X1 U23006 ( .B1(n12080), .B2(n20051), .A(n20040), .ZN(P1_U2931) );
  AOI22_X1 U23007 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20041) );
  OAI21_X1 U23008 ( .B1(n20042), .B2(n20051), .A(n20041), .ZN(P1_U2932) );
  INV_X1 U23009 ( .A(P1_LWORD_REG_3__SCAN_IN), .ZN(n20817) );
  OAI222_X1 U23010 ( .A1(n20800), .A2(n20817), .B1(n20051), .B2(n20888), .C1(
        n20044), .C2(n20043), .ZN(P1_U2933) );
  AOI22_X1 U23011 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20045) );
  OAI21_X1 U23012 ( .B1(n20046), .B2(n20051), .A(n20045), .ZN(P1_U2934) );
  AOI22_X1 U23013 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20047) );
  OAI21_X1 U23014 ( .B1(n20048), .B2(n20051), .A(n20047), .ZN(P1_U2935) );
  AOI22_X1 U23015 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n9734), .B1(n20049), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20050) );
  OAI21_X1 U23016 ( .B1(n20052), .B2(n20051), .A(n20050), .ZN(P1_U2936) );
  AOI22_X1 U23017 ( .A1(n20073), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20072), .ZN(n20054) );
  NAND2_X1 U23018 ( .A1(n20060), .A2(n20053), .ZN(n20062) );
  NAND2_X1 U23019 ( .A1(n20054), .A2(n20062), .ZN(P1_U2946) );
  AOI22_X1 U23020 ( .A1(n20073), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20072), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20056) );
  NAND2_X1 U23021 ( .A1(n20060), .A2(n20055), .ZN(n20066) );
  NAND2_X1 U23022 ( .A1(n20056), .A2(n20066), .ZN(P1_U2948) );
  AOI22_X1 U23023 ( .A1(n20073), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20072), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20058) );
  NAND2_X1 U23024 ( .A1(n20060), .A2(n20057), .ZN(n20068) );
  NAND2_X1 U23025 ( .A1(n20058), .A2(n20068), .ZN(P1_U2949) );
  AOI22_X1 U23026 ( .A1(n20073), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20072), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20061) );
  NAND2_X1 U23027 ( .A1(n20060), .A2(n20059), .ZN(n20074) );
  NAND2_X1 U23028 ( .A1(n20061), .A2(n20074), .ZN(P1_U2951) );
  AOI22_X1 U23029 ( .A1(n20073), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20072), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20063) );
  NAND2_X1 U23030 ( .A1(n20063), .A2(n20062), .ZN(P1_U2961) );
  AOI22_X1 U23031 ( .A1(n20073), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20072), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20065) );
  NAND2_X1 U23032 ( .A1(n20065), .A2(n20064), .ZN(P1_U2962) );
  AOI22_X1 U23033 ( .A1(n20073), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20072), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20067) );
  NAND2_X1 U23034 ( .A1(n20067), .A2(n20066), .ZN(P1_U2963) );
  AOI22_X1 U23035 ( .A1(n20073), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20072), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20069) );
  NAND2_X1 U23036 ( .A1(n20069), .A2(n20068), .ZN(P1_U2964) );
  AOI22_X1 U23037 ( .A1(n20073), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20072), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20071) );
  NAND2_X1 U23038 ( .A1(n20071), .A2(n20070), .ZN(P1_U2965) );
  AOI22_X1 U23039 ( .A1(n20073), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20072), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20075) );
  NAND2_X1 U23040 ( .A1(n20075), .A2(n20074), .ZN(P1_U2966) );
  AOI22_X1 U23041 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n13397), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20083) );
  XOR2_X1 U23042 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n20077), .Z(
        n20078) );
  XNOR2_X1 U23043 ( .A(n20079), .B(n20078), .ZN(n20087) );
  AOI22_X1 U23044 ( .A1(n20087), .A2(n20081), .B1(n14666), .B2(n20080), .ZN(
        n20082) );
  OAI211_X1 U23045 ( .C1(n20085), .C2(n20084), .A(n20083), .B(n20082), .ZN(
        P1_U2995) );
  AOI211_X1 U23046 ( .C1(n20086), .C2(n20111), .A(n20105), .B(n20104), .ZN(
        n20102) );
  AOI222_X1 U23047 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n13397), .B1(n20126), 
        .B2(n20088), .C1(n20128), .C2(n20087), .ZN(n20091) );
  OAI211_X1 U23048 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20098), .B(n20089), .ZN(n20090) );
  OAI211_X1 U23049 ( .C1(n20102), .C2(n20092), .A(n20091), .B(n20090), .ZN(
        P1_U3027) );
  INV_X1 U23050 ( .A(n20093), .ZN(n20094) );
  AOI21_X1 U23051 ( .B1(n20126), .B2(n20095), .A(n20094), .ZN(n20100) );
  INV_X1 U23052 ( .A(n20096), .ZN(n20097) );
  AOI22_X1 U23053 ( .A1(n20098), .A2(n20101), .B1(n20097), .B2(n20128), .ZN(
        n20099) );
  OAI211_X1 U23054 ( .C1(n20102), .C2(n20101), .A(n20100), .B(n20099), .ZN(
        P1_U3028) );
  OR2_X1 U23055 ( .A1(n20135), .A2(n20103), .ZN(n20121) );
  NOR2_X1 U23056 ( .A1(n20105), .A2(n20104), .ZN(n20119) );
  INV_X1 U23057 ( .A(n20106), .ZN(n20117) );
  INV_X1 U23058 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20923) );
  OAI22_X1 U23059 ( .A1(n20109), .A2(n20108), .B1(n20923), .B2(n20107), .ZN(
        n20116) );
  NOR2_X1 U23060 ( .A1(n20110), .A2(n20135), .ZN(n20112) );
  AOI21_X1 U23061 ( .B1(n20112), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n20111), .ZN(n20113) );
  NOR2_X1 U23062 ( .A1(n20114), .A2(n20113), .ZN(n20115) );
  AOI211_X1 U23063 ( .C1(n20117), .C2(n20128), .A(n20116), .B(n20115), .ZN(
        n20118) );
  OAI221_X1 U23064 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20121), .C1(
        n20120), .C2(n20119), .A(n20118), .ZN(P1_U3029) );
  NAND3_X1 U23065 ( .A1(n20135), .A2(n20123), .A3(n20122), .ZN(n20131) );
  AOI21_X1 U23066 ( .B1(n20126), .B2(n20125), .A(n20124), .ZN(n20130) );
  NAND3_X1 U23067 ( .A1(n20128), .A2(n13314), .A3(n20127), .ZN(n20129) );
  AND3_X1 U23068 ( .A1(n20131), .A2(n20130), .A3(n20129), .ZN(n20132) );
  OAI221_X1 U23069 ( .B1(n20135), .B2(n20134), .C1(n20135), .C2(n20133), .A(
        n20132), .ZN(P1_U3030) );
  AND2_X1 U23070 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20136), .ZN(
        P1_U3032) );
  INV_X1 U23071 ( .A(n20222), .ZN(n20138) );
  NAND2_X1 U23072 ( .A1(n20223), .A2(n20138), .ZN(n20369) );
  NAND2_X1 U23073 ( .A1(n20656), .A2(n20649), .ZN(n20139) );
  NAND2_X1 U23074 ( .A1(n20649), .A2(n21079), .ZN(n20517) );
  OAI21_X1 U23075 ( .B1(n20218), .B2(n20139), .A(n20517), .ZN(n20149) );
  OR2_X1 U23076 ( .A1(n20140), .A2(n20399), .ZN(n20225) );
  NOR2_X1 U23077 ( .A1(n20225), .A2(n20598), .ZN(n20147) );
  AND2_X1 U23078 ( .A1(n20146), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20459) );
  INV_X1 U23079 ( .A(n20457), .ZN(n20401) );
  OR2_X1 U23080 ( .A1(n20400), .A2(n20401), .ZN(n20290) );
  INV_X1 U23081 ( .A(n20290), .ZN(n20151) );
  AOI22_X1 U23082 ( .A1(n20149), .A2(n20147), .B1(n20459), .B2(n20151), .ZN(
        n20196) );
  NAND2_X1 U23083 ( .A1(n20141), .A2(n20185), .ZN(n20536) );
  NOR2_X2 U23084 ( .A1(n20142), .A2(n12861), .ZN(n20192) );
  NOR2_X2 U23085 ( .A1(n20143), .A2(n20142), .ZN(n20191) );
  AOI22_X1 U23086 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20192), .B1(DATAI_24_), 
        .B2(n20191), .ZN(n20660) );
  NAND2_X1 U23087 ( .A1(n20185), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20170) );
  OR2_X1 U23088 ( .A1(n20144), .A2(n20170), .ZN(n20525) );
  NAND3_X1 U23089 ( .A1(n20488), .A2(n12539), .A3(n20524), .ZN(n20198) );
  INV_X1 U23090 ( .A(n20198), .ZN(n20201) );
  NAND2_X1 U23091 ( .A1(n20568), .A2(n20201), .ZN(n20189) );
  OAI22_X1 U23092 ( .A1(n20656), .A2(n20660), .B1(n20525), .B2(n20189), .ZN(
        n20145) );
  INV_X1 U23093 ( .A(n20145), .ZN(n20153) );
  NOR2_X1 U23094 ( .A1(n20146), .A2(n11980), .ZN(n20523) );
  NOR2_X1 U23095 ( .A1(n20294), .A2(n20523), .ZN(n20465) );
  INV_X1 U23096 ( .A(n20147), .ZN(n20148) );
  AOI22_X1 U23097 ( .A1(n20149), .A2(n20148), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20189), .ZN(n20150) );
  OAI211_X1 U23098 ( .C1(n20151), .C2(n11980), .A(n20465), .B(n20150), .ZN(
        n20193) );
  AOI22_X1 U23099 ( .A1(DATAI_16_), .A2(n20191), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20192), .ZN(n20610) );
  INV_X1 U23100 ( .A(n20610), .ZN(n20657) );
  AOI22_X1 U23101 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20193), .B1(
        n20218), .B2(n20657), .ZN(n20152) );
  OAI211_X1 U23102 ( .C1(n20196), .C2(n20536), .A(n20153), .B(n20152), .ZN(
        P1_U3033) );
  NAND2_X1 U23103 ( .A1(n20154), .A2(n20185), .ZN(n20541) );
  AOI22_X1 U23104 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20192), .B1(DATAI_25_), 
        .B2(n20191), .ZN(n20666) );
  AND2_X1 U23105 ( .A1(n20155), .A2(n20187), .ZN(n20661) );
  INV_X1 U23106 ( .A(n20661), .ZN(n20537) );
  OAI22_X1 U23107 ( .A1(n20656), .A2(n20666), .B1(n20537), .B2(n20189), .ZN(
        n20156) );
  INV_X1 U23108 ( .A(n20156), .ZN(n20158) );
  AOI22_X1 U23109 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20192), .B1(DATAI_17_), 
        .B2(n20191), .ZN(n20614) );
  INV_X1 U23110 ( .A(n20614), .ZN(n20663) );
  AOI22_X1 U23111 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20193), .B1(
        n20218), .B2(n20663), .ZN(n20157) );
  OAI211_X1 U23112 ( .C1(n20196), .C2(n20541), .A(n20158), .B(n20157), .ZN(
        P1_U3034) );
  NAND2_X1 U23113 ( .A1(n20159), .A2(n20185), .ZN(n20546) );
  AOI22_X1 U23114 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20192), .B1(DATAI_26_), 
        .B2(n20191), .ZN(n20672) );
  INV_X1 U23115 ( .A(n20667), .ZN(n20542) );
  OAI22_X1 U23116 ( .A1(n20656), .A2(n20672), .B1(n20542), .B2(n20189), .ZN(
        n20161) );
  INV_X1 U23117 ( .A(n20161), .ZN(n20163) );
  AOI22_X1 U23118 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20192), .B1(DATAI_18_), 
        .B2(n20191), .ZN(n20618) );
  INV_X1 U23119 ( .A(n20618), .ZN(n20669) );
  AOI22_X1 U23120 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20193), .B1(
        n20218), .B2(n20669), .ZN(n20162) );
  OAI211_X1 U23121 ( .C1(n20196), .C2(n20546), .A(n20163), .B(n20162), .ZN(
        P1_U3035) );
  NAND2_X1 U23122 ( .A1(n20164), .A2(n20185), .ZN(n20551) );
  AOI22_X1 U23123 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20192), .B1(DATAI_27_), 
        .B2(n20191), .ZN(n20678) );
  INV_X1 U23124 ( .A(n20673), .ZN(n20547) );
  OAI22_X1 U23125 ( .A1(n20656), .A2(n20678), .B1(n20547), .B2(n20189), .ZN(
        n20166) );
  INV_X1 U23126 ( .A(n20166), .ZN(n20168) );
  AOI22_X1 U23127 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20192), .B1(DATAI_19_), 
        .B2(n20191), .ZN(n20622) );
  INV_X1 U23128 ( .A(n20622), .ZN(n20675) );
  AOI22_X1 U23129 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20193), .B1(
        n20218), .B2(n20675), .ZN(n20167) );
  OAI211_X1 U23130 ( .C1(n20196), .C2(n20551), .A(n20168), .B(n20167), .ZN(
        P1_U3036) );
  NAND2_X1 U23131 ( .A1(n20169), .A2(n20185), .ZN(n20556) );
  AOI22_X1 U23132 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20192), .B1(DATAI_28_), 
        .B2(n20191), .ZN(n20684) );
  OR2_X1 U23133 ( .A1(n20171), .A2(n20170), .ZN(n20552) );
  OAI22_X1 U23134 ( .A1(n20656), .A2(n20684), .B1(n20552), .B2(n20189), .ZN(
        n20172) );
  INV_X1 U23135 ( .A(n20172), .ZN(n20174) );
  AOI22_X1 U23136 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20192), .B1(DATAI_20_), 
        .B2(n20191), .ZN(n20626) );
  INV_X1 U23137 ( .A(n20626), .ZN(n20681) );
  AOI22_X1 U23138 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20193), .B1(
        n20218), .B2(n20681), .ZN(n20173) );
  OAI211_X1 U23139 ( .C1(n20196), .C2(n20556), .A(n20174), .B(n20173), .ZN(
        P1_U3037) );
  NAND2_X1 U23140 ( .A1(n20175), .A2(n20185), .ZN(n20561) );
  AOI22_X1 U23141 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20192), .B1(DATAI_29_), 
        .B2(n20191), .ZN(n20690) );
  INV_X1 U23142 ( .A(n20685), .ZN(n20557) );
  OAI22_X1 U23143 ( .A1(n20656), .A2(n20690), .B1(n20557), .B2(n20189), .ZN(
        n20177) );
  INV_X1 U23144 ( .A(n20177), .ZN(n20179) );
  AOI22_X1 U23145 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20192), .B1(DATAI_21_), 
        .B2(n20191), .ZN(n20630) );
  INV_X1 U23146 ( .A(n20630), .ZN(n20687) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20193), .B1(
        n20218), .B2(n20687), .ZN(n20178) );
  OAI211_X1 U23148 ( .C1(n20196), .C2(n20561), .A(n20179), .B(n20178), .ZN(
        P1_U3038) );
  NAND2_X1 U23149 ( .A1(n20180), .A2(n20185), .ZN(n21074) );
  AOI22_X1 U23150 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20192), .B1(DATAI_30_), 
        .B2(n20191), .ZN(n21073) );
  INV_X1 U23151 ( .A(n20691), .ZN(n21069) );
  OAI22_X1 U23152 ( .A1(n20656), .A2(n21073), .B1(n21069), .B2(n20189), .ZN(
        n20182) );
  INV_X1 U23153 ( .A(n20182), .ZN(n20184) );
  AOI22_X1 U23154 ( .A1(DATAI_22_), .A2(n20191), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20192), .ZN(n21070) );
  INV_X1 U23155 ( .A(n21070), .ZN(n20693) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20193), .B1(
        n20218), .B2(n20693), .ZN(n20183) );
  OAI211_X1 U23157 ( .C1(n20196), .C2(n21074), .A(n20184), .B(n20183), .ZN(
        P1_U3039) );
  NAND2_X1 U23158 ( .A1(n20186), .A2(n20185), .ZN(n20567) );
  AOI22_X1 U23159 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20192), .B1(DATAI_31_), 
        .B2(n20191), .ZN(n20706) );
  INV_X1 U23160 ( .A(n20697), .ZN(n20562) );
  OAI22_X1 U23161 ( .A1(n20656), .A2(n20706), .B1(n20562), .B2(n20189), .ZN(
        n20190) );
  INV_X1 U23162 ( .A(n20190), .ZN(n20195) );
  AOI22_X1 U23163 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20192), .B1(DATAI_23_), 
        .B2(n20191), .ZN(n20641) );
  INV_X1 U23164 ( .A(n20641), .ZN(n20700) );
  AOI22_X1 U23165 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20193), .B1(
        n20218), .B2(n20700), .ZN(n20194) );
  OAI211_X1 U23166 ( .C1(n20196), .C2(n20567), .A(n20195), .B(n20194), .ZN(
        P1_U3040) );
  INV_X1 U23167 ( .A(n20225), .ZN(n20258) );
  INV_X1 U23168 ( .A(n20197), .ZN(n20569) );
  NOR2_X1 U23169 ( .A1(n20568), .A2(n20198), .ZN(n20216) );
  AOI21_X1 U23170 ( .B1(n20258), .B2(n20569), .A(n20216), .ZN(n20199) );
  OAI22_X1 U23171 ( .A1(n20199), .A2(n20644), .B1(n20198), .B2(n11980), .ZN(
        n20217) );
  AOI22_X1 U23172 ( .A1(n20217), .A2(n20646), .B1(n20645), .B2(n20216), .ZN(
        n20203) );
  AOI21_X1 U23173 ( .B1(n20568), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20294), 
        .ZN(n20653) );
  OAI211_X1 U23174 ( .C1(n20262), .C2(n20431), .A(n20654), .B(n20199), .ZN(
        n20200) );
  OAI211_X1 U23175 ( .C1(n20649), .C2(n20201), .A(n20653), .B(n20200), .ZN(
        n20219) );
  INV_X1 U23176 ( .A(n20660), .ZN(n20607) );
  AOI22_X1 U23177 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20607), .ZN(n20202) );
  OAI211_X1 U23178 ( .C1(n20610), .C2(n20250), .A(n20203), .B(n20202), .ZN(
        P1_U3041) );
  AOI22_X1 U23179 ( .A1(n20217), .A2(n20662), .B1(n20661), .B2(n20216), .ZN(
        n20205) );
  INV_X1 U23180 ( .A(n20666), .ZN(n20611) );
  AOI22_X1 U23181 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20611), .ZN(n20204) );
  OAI211_X1 U23182 ( .C1(n20614), .C2(n20250), .A(n20205), .B(n20204), .ZN(
        P1_U3042) );
  AOI22_X1 U23183 ( .A1(n20217), .A2(n20668), .B1(n20667), .B2(n20216), .ZN(
        n20207) );
  INV_X1 U23184 ( .A(n20672), .ZN(n20615) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20615), .ZN(n20206) );
  OAI211_X1 U23186 ( .C1(n20618), .C2(n20250), .A(n20207), .B(n20206), .ZN(
        P1_U3043) );
  AOI22_X1 U23187 ( .A1(n20217), .A2(n20674), .B1(n20673), .B2(n20216), .ZN(
        n20209) );
  INV_X1 U23188 ( .A(n20678), .ZN(n20619) );
  AOI22_X1 U23189 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20619), .ZN(n20208) );
  OAI211_X1 U23190 ( .C1(n20622), .C2(n20250), .A(n20209), .B(n20208), .ZN(
        P1_U3044) );
  AOI22_X1 U23191 ( .A1(n20217), .A2(n20680), .B1(n20679), .B2(n20216), .ZN(
        n20211) );
  INV_X1 U23192 ( .A(n20684), .ZN(n20623) );
  AOI22_X1 U23193 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20623), .ZN(n20210) );
  OAI211_X1 U23194 ( .C1(n20626), .C2(n20250), .A(n20211), .B(n20210), .ZN(
        P1_U3045) );
  AOI22_X1 U23195 ( .A1(n20217), .A2(n20686), .B1(n20685), .B2(n20216), .ZN(
        n20213) );
  INV_X1 U23196 ( .A(n20690), .ZN(n20627) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20627), .ZN(n20212) );
  OAI211_X1 U23198 ( .C1(n20630), .C2(n20250), .A(n20213), .B(n20212), .ZN(
        P1_U3046) );
  AOI22_X1 U23199 ( .A1(n20217), .A2(n20692), .B1(n20691), .B2(n20216), .ZN(
        n20215) );
  INV_X1 U23200 ( .A(n21073), .ZN(n20631) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20631), .ZN(n20214) );
  OAI211_X1 U23202 ( .C1(n21070), .C2(n20250), .A(n20215), .B(n20214), .ZN(
        P1_U3047) );
  AOI22_X1 U23203 ( .A1(n20217), .A2(n20698), .B1(n20697), .B2(n20216), .ZN(
        n20221) );
  INV_X1 U23204 ( .A(n20706), .ZN(n20636) );
  AOI22_X1 U23205 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20219), .B1(
        n20218), .B2(n20636), .ZN(n20220) );
  OAI211_X1 U23206 ( .C1(n20641), .C2(n20250), .A(n20221), .B(n20220), .ZN(
        P1_U3048) );
  NOR2_X2 U23207 ( .A1(n20262), .A2(n20455), .ZN(n20283) );
  NAND2_X1 U23208 ( .A1(n20250), .A2(n20649), .ZN(n20224) );
  OAI21_X1 U23209 ( .B1(n20283), .B2(n20224), .A(n20517), .ZN(n20227) );
  NOR2_X1 U23210 ( .A1(n20225), .A2(n20521), .ZN(n20229) );
  NOR3_X1 U23211 ( .A1(n20524), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20263) );
  NAND2_X1 U23212 ( .A1(n20568), .A2(n20263), .ZN(n20249) );
  OAI22_X1 U23213 ( .A1(n20250), .A2(n20660), .B1(n20525), .B2(n20249), .ZN(
        n20226) );
  INV_X1 U23214 ( .A(n20226), .ZN(n20232) );
  INV_X1 U23215 ( .A(n20227), .ZN(n20230) );
  NOR2_X1 U23216 ( .A1(n10220), .A2(n11980), .ZN(n20345) );
  AOI21_X1 U23217 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20249), .A(n20345), 
        .ZN(n20228) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20252), .B1(
        n20283), .B2(n20657), .ZN(n20231) );
  OAI211_X1 U23219 ( .C1(n20255), .C2(n20536), .A(n20232), .B(n20231), .ZN(
        P1_U3049) );
  INV_X1 U23220 ( .A(n20249), .ZN(n20242) );
  AOI22_X1 U23221 ( .A1(n20283), .A2(n20663), .B1(n20661), .B2(n20242), .ZN(
        n20234) );
  INV_X1 U23222 ( .A(n20250), .ZN(n20243) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20252), .B1(
        n20243), .B2(n20611), .ZN(n20233) );
  OAI211_X1 U23224 ( .C1(n20255), .C2(n20541), .A(n20234), .B(n20233), .ZN(
        P1_U3050) );
  AOI22_X1 U23225 ( .A1(n20283), .A2(n20669), .B1(n20242), .B2(n20667), .ZN(
        n20236) );
  AOI22_X1 U23226 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20252), .B1(
        n20243), .B2(n20615), .ZN(n20235) );
  OAI211_X1 U23227 ( .C1(n20255), .C2(n20546), .A(n20236), .B(n20235), .ZN(
        P1_U3051) );
  OAI22_X1 U23228 ( .A1(n20250), .A2(n20678), .B1(n20249), .B2(n20547), .ZN(
        n20237) );
  INV_X1 U23229 ( .A(n20237), .ZN(n20239) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20252), .B1(
        n20283), .B2(n20675), .ZN(n20238) );
  OAI211_X1 U23231 ( .C1(n20255), .C2(n20551), .A(n20239), .B(n20238), .ZN(
        P1_U3052) );
  AOI22_X1 U23232 ( .A1(n20283), .A2(n20681), .B1(n20242), .B2(n20679), .ZN(
        n20241) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20252), .B1(
        n20243), .B2(n20623), .ZN(n20240) );
  OAI211_X1 U23234 ( .C1(n20255), .C2(n20556), .A(n20241), .B(n20240), .ZN(
        P1_U3053) );
  AOI22_X1 U23235 ( .A1(n20283), .A2(n20687), .B1(n20242), .B2(n20685), .ZN(
        n20245) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20252), .B1(
        n20243), .B2(n20627), .ZN(n20244) );
  OAI211_X1 U23237 ( .C1(n20255), .C2(n20561), .A(n20245), .B(n20244), .ZN(
        P1_U3054) );
  OAI22_X1 U23238 ( .A1(n20250), .A2(n21073), .B1(n20249), .B2(n21069), .ZN(
        n20246) );
  INV_X1 U23239 ( .A(n20246), .ZN(n20248) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20252), .B1(
        n20283), .B2(n20693), .ZN(n20247) );
  OAI211_X1 U23241 ( .C1(n20255), .C2(n21074), .A(n20248), .B(n20247), .ZN(
        P1_U3055) );
  OAI22_X1 U23242 ( .A1(n20250), .A2(n20706), .B1(n20562), .B2(n20249), .ZN(
        n20251) );
  INV_X1 U23243 ( .A(n20251), .ZN(n20254) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20252), .B1(
        n20283), .B2(n20700), .ZN(n20253) );
  OAI211_X1 U23245 ( .C1(n20255), .C2(n20567), .A(n20254), .B(n20253), .ZN(
        P1_U3056) );
  AND2_X1 U23246 ( .A1(n20257), .A2(n20256), .ZN(n20642) );
  NOR2_X1 U23247 ( .A1(n20489), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20282) );
  AOI21_X1 U23248 ( .B1(n20258), .B2(n20642), .A(n20282), .ZN(n20265) );
  INV_X1 U23249 ( .A(n20265), .ZN(n20261) );
  INV_X1 U23250 ( .A(n20262), .ZN(n20260) );
  AOI21_X1 U23251 ( .B1(n20260), .B2(n20259), .A(n20644), .ZN(n20266) );
  AOI22_X1 U23252 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20263), .B1(n20261), 
        .B2(n20266), .ZN(n20287) );
  NOR2_X2 U23253 ( .A1(n20262), .A2(n20369), .ZN(n20312) );
  AOI22_X1 U23254 ( .A1(n20312), .A2(n20657), .B1(n20645), .B2(n20282), .ZN(
        n20269) );
  OAI21_X1 U23255 ( .B1(n20654), .B2(n20263), .A(n20653), .ZN(n20264) );
  AOI21_X1 U23256 ( .B1(n20266), .B2(n20265), .A(n20264), .ZN(n20267) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20284), .B1(
        n20283), .B2(n20607), .ZN(n20268) );
  OAI211_X1 U23258 ( .C1(n20287), .C2(n20536), .A(n20269), .B(n20268), .ZN(
        P1_U3057) );
  AOI22_X1 U23259 ( .A1(n20312), .A2(n20663), .B1(n20282), .B2(n20661), .ZN(
        n20271) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20284), .B1(
        n20283), .B2(n20611), .ZN(n20270) );
  OAI211_X1 U23261 ( .C1(n20287), .C2(n20541), .A(n20271), .B(n20270), .ZN(
        P1_U3058) );
  AOI22_X1 U23262 ( .A1(n20283), .A2(n20615), .B1(n20282), .B2(n20667), .ZN(
        n20273) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20284), .B1(
        n20312), .B2(n20669), .ZN(n20272) );
  OAI211_X1 U23264 ( .C1(n20287), .C2(n20546), .A(n20273), .B(n20272), .ZN(
        P1_U3059) );
  AOI22_X1 U23265 ( .A1(n20283), .A2(n20619), .B1(n20282), .B2(n20673), .ZN(
        n20275) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20284), .B1(
        n20312), .B2(n20675), .ZN(n20274) );
  OAI211_X1 U23267 ( .C1(n20287), .C2(n20551), .A(n20275), .B(n20274), .ZN(
        P1_U3060) );
  AOI22_X1 U23268 ( .A1(n20283), .A2(n20623), .B1(n20282), .B2(n20679), .ZN(
        n20277) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20284), .B1(
        n20312), .B2(n20681), .ZN(n20276) );
  OAI211_X1 U23270 ( .C1(n20287), .C2(n20556), .A(n20277), .B(n20276), .ZN(
        P1_U3061) );
  AOI22_X1 U23271 ( .A1(n20283), .A2(n20627), .B1(n20282), .B2(n20685), .ZN(
        n20279) );
  AOI22_X1 U23272 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20284), .B1(
        n20312), .B2(n20687), .ZN(n20278) );
  OAI211_X1 U23273 ( .C1(n20287), .C2(n20561), .A(n20279), .B(n20278), .ZN(
        P1_U3062) );
  AOI22_X1 U23274 ( .A1(n20283), .A2(n20631), .B1(n20282), .B2(n20691), .ZN(
        n20281) );
  AOI22_X1 U23275 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20284), .B1(
        n20312), .B2(n20693), .ZN(n20280) );
  OAI211_X1 U23276 ( .C1(n20287), .C2(n21074), .A(n20281), .B(n20280), .ZN(
        P1_U3063) );
  AOI22_X1 U23277 ( .A1(n20312), .A2(n20700), .B1(n20282), .B2(n20697), .ZN(
        n20286) );
  AOI22_X1 U23278 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20284), .B1(
        n20283), .B2(n20636), .ZN(n20285) );
  OAI211_X1 U23279 ( .C1(n20287), .C2(n20567), .A(n20286), .B(n20285), .ZN(
        P1_U3064) );
  INV_X1 U23280 ( .A(n20523), .ZN(n20599) );
  NOR2_X1 U23281 ( .A1(n20520), .A2(n20288), .ZN(n20372) );
  NAND3_X1 U23282 ( .A1(n20372), .A2(n20654), .A3(n20521), .ZN(n20289) );
  OAI21_X1 U23283 ( .B1(n20599), .B2(n20290), .A(n20289), .ZN(n20311) );
  NAND3_X1 U23284 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20488), .A3(
        n20524), .ZN(n20317) );
  NOR2_X1 U23285 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20317), .ZN(
        n20310) );
  AOI22_X1 U23286 ( .A1(n20311), .A2(n20646), .B1(n20645), .B2(n20310), .ZN(
        n20297) );
  INV_X1 U23287 ( .A(n20312), .ZN(n20291) );
  AOI21_X1 U23288 ( .B1(n20291), .B2(n20341), .A(n21079), .ZN(n20292) );
  AOI21_X1 U23289 ( .B1(n20372), .B2(n20521), .A(n20292), .ZN(n20293) );
  NOR2_X1 U23290 ( .A1(n20293), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20295) );
  NOR2_X1 U23291 ( .A1(n20294), .A2(n20459), .ZN(n20605) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20607), .ZN(n20296) );
  OAI211_X1 U23293 ( .C1(n20610), .C2(n20341), .A(n20297), .B(n20296), .ZN(
        P1_U3065) );
  AOI22_X1 U23294 ( .A1(n20311), .A2(n20662), .B1(n20661), .B2(n20310), .ZN(
        n20299) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20611), .ZN(n20298) );
  OAI211_X1 U23296 ( .C1(n20614), .C2(n20341), .A(n20299), .B(n20298), .ZN(
        P1_U3066) );
  AOI22_X1 U23297 ( .A1(n20311), .A2(n20668), .B1(n20667), .B2(n20310), .ZN(
        n20301) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20615), .ZN(n20300) );
  OAI211_X1 U23299 ( .C1(n20618), .C2(n20341), .A(n20301), .B(n20300), .ZN(
        P1_U3067) );
  AOI22_X1 U23300 ( .A1(n20311), .A2(n20674), .B1(n20673), .B2(n20310), .ZN(
        n20303) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20619), .ZN(n20302) );
  OAI211_X1 U23302 ( .C1(n20622), .C2(n20341), .A(n20303), .B(n20302), .ZN(
        P1_U3068) );
  AOI22_X1 U23303 ( .A1(n20311), .A2(n20680), .B1(n20679), .B2(n20310), .ZN(
        n20305) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20623), .ZN(n20304) );
  OAI211_X1 U23305 ( .C1(n20626), .C2(n20341), .A(n20305), .B(n20304), .ZN(
        P1_U3069) );
  AOI22_X1 U23306 ( .A1(n20311), .A2(n20686), .B1(n20685), .B2(n20310), .ZN(
        n20307) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20627), .ZN(n20306) );
  OAI211_X1 U23308 ( .C1(n20630), .C2(n20341), .A(n20307), .B(n20306), .ZN(
        P1_U3070) );
  AOI22_X1 U23309 ( .A1(n20311), .A2(n20692), .B1(n20691), .B2(n20310), .ZN(
        n20309) );
  AOI22_X1 U23310 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20631), .ZN(n20308) );
  OAI211_X1 U23311 ( .C1(n21070), .C2(n20341), .A(n20309), .B(n20308), .ZN(
        P1_U3071) );
  AOI22_X1 U23312 ( .A1(n20311), .A2(n20698), .B1(n20697), .B2(n20310), .ZN(
        n20315) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20636), .ZN(n20314) );
  OAI211_X1 U23314 ( .C1(n20641), .C2(n20341), .A(n20315), .B(n20314), .ZN(
        P1_U3072) );
  NOR2_X1 U23315 ( .A1(n20568), .A2(n20317), .ZN(n20336) );
  AOI21_X1 U23316 ( .B1(n20372), .B2(n20569), .A(n20336), .ZN(n20316) );
  OAI22_X1 U23317 ( .A1(n20316), .A2(n20644), .B1(n20317), .B2(n11980), .ZN(
        n20337) );
  AOI22_X1 U23318 ( .A1(n20337), .A2(n20646), .B1(n20645), .B2(n20336), .ZN(
        n20323) );
  INV_X1 U23319 ( .A(n20317), .ZN(n20320) );
  INV_X1 U23320 ( .A(n20370), .ZN(n20318) );
  NOR3_X1 U23321 ( .A1(n20318), .A2(n20644), .A3(n20431), .ZN(n20319) );
  OAI21_X1 U23322 ( .B1(n20320), .B2(n20319), .A(n20653), .ZN(n20338) );
  INV_X1 U23323 ( .A(n20576), .ZN(n20321) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20338), .B1(
        n20364), .B2(n20657), .ZN(n20322) );
  OAI211_X1 U23325 ( .C1(n20660), .C2(n20341), .A(n20323), .B(n20322), .ZN(
        P1_U3073) );
  AOI22_X1 U23326 ( .A1(n20337), .A2(n20662), .B1(n20661), .B2(n20336), .ZN(
        n20325) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20338), .B1(
        n20364), .B2(n20663), .ZN(n20324) );
  OAI211_X1 U23328 ( .C1(n20666), .C2(n20341), .A(n20325), .B(n20324), .ZN(
        P1_U3074) );
  AOI22_X1 U23329 ( .A1(n20337), .A2(n20668), .B1(n20667), .B2(n20336), .ZN(
        n20327) );
  AOI22_X1 U23330 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20338), .B1(
        n20364), .B2(n20669), .ZN(n20326) );
  OAI211_X1 U23331 ( .C1(n20672), .C2(n20341), .A(n20327), .B(n20326), .ZN(
        P1_U3075) );
  AOI22_X1 U23332 ( .A1(n20337), .A2(n20674), .B1(n20673), .B2(n20336), .ZN(
        n20329) );
  AOI22_X1 U23333 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20338), .B1(
        n20364), .B2(n20675), .ZN(n20328) );
  OAI211_X1 U23334 ( .C1(n20678), .C2(n20341), .A(n20329), .B(n20328), .ZN(
        P1_U3076) );
  AOI22_X1 U23335 ( .A1(n20337), .A2(n20680), .B1(n20679), .B2(n20336), .ZN(
        n20331) );
  AOI22_X1 U23336 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20338), .B1(
        n20364), .B2(n20681), .ZN(n20330) );
  OAI211_X1 U23337 ( .C1(n20684), .C2(n20341), .A(n20331), .B(n20330), .ZN(
        P1_U3077) );
  AOI22_X1 U23338 ( .A1(n20337), .A2(n20686), .B1(n20685), .B2(n20336), .ZN(
        n20333) );
  AOI22_X1 U23339 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20338), .B1(
        n20364), .B2(n20687), .ZN(n20332) );
  OAI211_X1 U23340 ( .C1(n20690), .C2(n20341), .A(n20333), .B(n20332), .ZN(
        P1_U3078) );
  AOI22_X1 U23341 ( .A1(n20337), .A2(n20692), .B1(n20691), .B2(n20336), .ZN(
        n20335) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20338), .B1(
        n20364), .B2(n20693), .ZN(n20334) );
  OAI211_X1 U23343 ( .C1(n21073), .C2(n20341), .A(n20335), .B(n20334), .ZN(
        P1_U3079) );
  AOI22_X1 U23344 ( .A1(n20337), .A2(n20698), .B1(n20697), .B2(n20336), .ZN(
        n20340) );
  AOI22_X1 U23345 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20338), .B1(
        n20364), .B2(n20700), .ZN(n20339) );
  OAI211_X1 U23346 ( .C1(n20706), .C2(n20341), .A(n20340), .B(n20339), .ZN(
        P1_U3080) );
  INV_X1 U23347 ( .A(n20364), .ZN(n20342) );
  NAND2_X1 U23348 ( .A1(n20342), .A2(n20654), .ZN(n20343) );
  INV_X1 U23349 ( .A(n20455), .ZN(n20596) );
  OAI21_X1 U23350 ( .B1(n20343), .B2(n20394), .A(n20517), .ZN(n20347) );
  AND2_X1 U23351 ( .A1(n20372), .A2(n20598), .ZN(n20344) );
  INV_X1 U23352 ( .A(n20377), .ZN(n20373) );
  NOR2_X1 U23353 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20373), .ZN(
        n20363) );
  AOI22_X1 U23354 ( .A1(n20394), .A2(n20657), .B1(n20645), .B2(n20363), .ZN(
        n20350) );
  INV_X1 U23355 ( .A(n20344), .ZN(n20346) );
  AOI21_X1 U23356 ( .B1(n20347), .B2(n20346), .A(n20345), .ZN(n20348) );
  OAI211_X1 U23357 ( .C1(n20363), .C2(n20532), .A(n20605), .B(n20348), .ZN(
        n20365) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20365), .B1(
        n20364), .B2(n20607), .ZN(n20349) );
  OAI211_X1 U23359 ( .C1(n20368), .C2(n20536), .A(n20350), .B(n20349), .ZN(
        P1_U3081) );
  AOI22_X1 U23360 ( .A1(n20394), .A2(n20663), .B1(n20661), .B2(n20363), .ZN(
        n20352) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20365), .B1(
        n20364), .B2(n20611), .ZN(n20351) );
  OAI211_X1 U23362 ( .C1(n20368), .C2(n20541), .A(n20352), .B(n20351), .ZN(
        P1_U3082) );
  AOI22_X1 U23363 ( .A1(n20364), .A2(n20615), .B1(n20667), .B2(n20363), .ZN(
        n20354) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20365), .B1(
        n20394), .B2(n20669), .ZN(n20353) );
  OAI211_X1 U23365 ( .C1(n20368), .C2(n20546), .A(n20354), .B(n20353), .ZN(
        P1_U3083) );
  AOI22_X1 U23366 ( .A1(n20394), .A2(n20675), .B1(n20673), .B2(n20363), .ZN(
        n20356) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20365), .B1(
        n20364), .B2(n20619), .ZN(n20355) );
  OAI211_X1 U23368 ( .C1(n20368), .C2(n20551), .A(n20356), .B(n20355), .ZN(
        P1_U3084) );
  AOI22_X1 U23369 ( .A1(n20364), .A2(n20623), .B1(n20679), .B2(n20363), .ZN(
        n20358) );
  AOI22_X1 U23370 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20365), .B1(
        n20394), .B2(n20681), .ZN(n20357) );
  OAI211_X1 U23371 ( .C1(n20368), .C2(n20556), .A(n20358), .B(n20357), .ZN(
        P1_U3085) );
  AOI22_X1 U23372 ( .A1(n20394), .A2(n20687), .B1(n20685), .B2(n20363), .ZN(
        n20360) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20365), .B1(
        n20364), .B2(n20627), .ZN(n20359) );
  OAI211_X1 U23374 ( .C1(n20368), .C2(n20561), .A(n20360), .B(n20359), .ZN(
        P1_U3086) );
  AOI22_X1 U23375 ( .A1(n20394), .A2(n20693), .B1(n20691), .B2(n20363), .ZN(
        n20362) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20365), .B1(
        n20364), .B2(n20631), .ZN(n20361) );
  OAI211_X1 U23377 ( .C1(n20368), .C2(n21074), .A(n20362), .B(n20361), .ZN(
        P1_U3087) );
  AOI22_X1 U23378 ( .A1(n20394), .A2(n20700), .B1(n20697), .B2(n20363), .ZN(
        n20367) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20365), .B1(
        n20364), .B2(n20636), .ZN(n20366) );
  OAI211_X1 U23380 ( .C1(n20368), .C2(n20567), .A(n20367), .B(n20366), .ZN(
        P1_U3088) );
  INV_X1 U23381 ( .A(n20371), .ZN(n20392) );
  AOI21_X1 U23382 ( .B1(n20372), .B2(n20642), .A(n20392), .ZN(n20374) );
  OAI22_X1 U23383 ( .A1(n20374), .A2(n20644), .B1(n20373), .B2(n11980), .ZN(
        n20393) );
  AOI22_X1 U23384 ( .A1(n20393), .A2(n20646), .B1(n20645), .B2(n20392), .ZN(
        n20379) );
  NAND2_X1 U23385 ( .A1(n20375), .A2(n20374), .ZN(n20376) );
  OAI221_X1 U23386 ( .B1(n20654), .B2(n20377), .C1(n20644), .C2(n20376), .A(
        n20653), .ZN(n20395) );
  AOI22_X1 U23387 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20607), .ZN(n20378) );
  OAI211_X1 U23388 ( .C1(n20610), .C2(n20404), .A(n20379), .B(n20378), .ZN(
        P1_U3089) );
  AOI22_X1 U23389 ( .A1(n20393), .A2(n20662), .B1(n20661), .B2(n20392), .ZN(
        n20381) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20611), .ZN(n20380) );
  OAI211_X1 U23391 ( .C1(n20614), .C2(n20404), .A(n20381), .B(n20380), .ZN(
        P1_U3090) );
  AOI22_X1 U23392 ( .A1(n20393), .A2(n20668), .B1(n20667), .B2(n20392), .ZN(
        n20383) );
  AOI22_X1 U23393 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20615), .ZN(n20382) );
  OAI211_X1 U23394 ( .C1(n20618), .C2(n20404), .A(n20383), .B(n20382), .ZN(
        P1_U3091) );
  AOI22_X1 U23395 ( .A1(n20393), .A2(n20674), .B1(n20673), .B2(n20392), .ZN(
        n20385) );
  AOI22_X1 U23396 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20619), .ZN(n20384) );
  OAI211_X1 U23397 ( .C1(n20622), .C2(n20404), .A(n20385), .B(n20384), .ZN(
        P1_U3092) );
  AOI22_X1 U23398 ( .A1(n20393), .A2(n20680), .B1(n20679), .B2(n20392), .ZN(
        n20387) );
  AOI22_X1 U23399 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20623), .ZN(n20386) );
  OAI211_X1 U23400 ( .C1(n20626), .C2(n20404), .A(n20387), .B(n20386), .ZN(
        P1_U3093) );
  AOI22_X1 U23401 ( .A1(n20393), .A2(n20686), .B1(n20685), .B2(n20392), .ZN(
        n20389) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20627), .ZN(n20388) );
  OAI211_X1 U23403 ( .C1(n20630), .C2(n20404), .A(n20389), .B(n20388), .ZN(
        P1_U3094) );
  AOI22_X1 U23404 ( .A1(n20393), .A2(n20692), .B1(n20691), .B2(n20392), .ZN(
        n20391) );
  AOI22_X1 U23405 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20631), .ZN(n20390) );
  OAI211_X1 U23406 ( .C1(n21070), .C2(n20404), .A(n20391), .B(n20390), .ZN(
        P1_U3095) );
  AOI22_X1 U23407 ( .A1(n20393), .A2(n20698), .B1(n20697), .B2(n20392), .ZN(
        n20397) );
  AOI22_X1 U23408 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20395), .B1(
        n20394), .B2(n20636), .ZN(n20396) );
  OAI211_X1 U23409 ( .C1(n20641), .C2(n20404), .A(n20397), .B(n20396), .ZN(
        P1_U3096) );
  AND2_X1 U23410 ( .A1(n20399), .A2(n20520), .ZN(n20490) );
  NAND3_X1 U23411 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12539), .A3(
        n20524), .ZN(n20429) );
  NOR2_X1 U23412 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20429), .ZN(
        n20423) );
  AOI21_X1 U23413 ( .B1(n20490), .B2(n20521), .A(n20423), .ZN(n20406) );
  INV_X1 U23414 ( .A(n20459), .ZN(n20403) );
  INV_X1 U23415 ( .A(n20400), .ZN(n20402) );
  NOR2_X1 U23416 ( .A1(n20402), .A2(n20401), .ZN(n20522) );
  INV_X1 U23417 ( .A(n20522), .ZN(n20528) );
  OAI22_X1 U23418 ( .A1(n20406), .A2(n20644), .B1(n20403), .B2(n20528), .ZN(
        n20424) );
  AOI22_X1 U23419 ( .A1(n20424), .A2(n20646), .B1(n20645), .B2(n20423), .ZN(
        n20410) );
  INV_X1 U23420 ( .A(n20453), .ZN(n20405) );
  OAI21_X1 U23421 ( .B1(n20405), .B2(n20425), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20407) );
  NAND2_X1 U23422 ( .A1(n20407), .A2(n20406), .ZN(n20408) );
  OAI211_X1 U23423 ( .C1(n20423), .C2(n20532), .A(n20465), .B(n20408), .ZN(
        n20426) );
  AOI22_X1 U23424 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20607), .ZN(n20409) );
  OAI211_X1 U23425 ( .C1(n20610), .C2(n20453), .A(n20410), .B(n20409), .ZN(
        P1_U3097) );
  AOI22_X1 U23426 ( .A1(n20424), .A2(n20662), .B1(n20661), .B2(n20423), .ZN(
        n20412) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20611), .ZN(n20411) );
  OAI211_X1 U23428 ( .C1(n20614), .C2(n20453), .A(n20412), .B(n20411), .ZN(
        P1_U3098) );
  AOI22_X1 U23429 ( .A1(n20424), .A2(n20668), .B1(n20667), .B2(n20423), .ZN(
        n20414) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20615), .ZN(n20413) );
  OAI211_X1 U23431 ( .C1(n20618), .C2(n20453), .A(n20414), .B(n20413), .ZN(
        P1_U3099) );
  AOI22_X1 U23432 ( .A1(n20424), .A2(n20674), .B1(n20673), .B2(n20423), .ZN(
        n20416) );
  AOI22_X1 U23433 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20619), .ZN(n20415) );
  OAI211_X1 U23434 ( .C1(n20622), .C2(n20453), .A(n20416), .B(n20415), .ZN(
        P1_U3100) );
  AOI22_X1 U23435 ( .A1(n20424), .A2(n20680), .B1(n20679), .B2(n20423), .ZN(
        n20418) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20623), .ZN(n20417) );
  OAI211_X1 U23437 ( .C1(n20626), .C2(n20453), .A(n20418), .B(n20417), .ZN(
        P1_U3101) );
  AOI22_X1 U23438 ( .A1(n20424), .A2(n20686), .B1(n20685), .B2(n20423), .ZN(
        n20420) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20627), .ZN(n20419) );
  OAI211_X1 U23440 ( .C1(n20630), .C2(n20453), .A(n20420), .B(n20419), .ZN(
        P1_U3102) );
  AOI22_X1 U23441 ( .A1(n20424), .A2(n20692), .B1(n20691), .B2(n20423), .ZN(
        n20422) );
  AOI22_X1 U23442 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20631), .ZN(n20421) );
  OAI211_X1 U23443 ( .C1(n21070), .C2(n20453), .A(n20422), .B(n20421), .ZN(
        P1_U3103) );
  AOI22_X1 U23444 ( .A1(n20424), .A2(n20698), .B1(n20697), .B2(n20423), .ZN(
        n20428) );
  AOI22_X1 U23445 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20636), .ZN(n20427) );
  OAI211_X1 U23446 ( .C1(n20641), .C2(n20453), .A(n20428), .B(n20427), .ZN(
        P1_U3104) );
  NOR2_X1 U23447 ( .A1(n20568), .A2(n20429), .ZN(n20448) );
  AOI21_X1 U23448 ( .B1(n20490), .B2(n20569), .A(n20448), .ZN(n20430) );
  OAI22_X1 U23449 ( .A1(n20430), .A2(n20644), .B1(n20429), .B2(n11980), .ZN(
        n20449) );
  AOI22_X1 U23450 ( .A1(n20449), .A2(n20646), .B1(n20645), .B2(n20448), .ZN(
        n20435) );
  INV_X1 U23451 ( .A(n20429), .ZN(n20433) );
  OAI211_X1 U23452 ( .C1(n20493), .C2(n20431), .A(n20649), .B(n20430), .ZN(
        n20432) );
  OAI211_X1 U23453 ( .C1(n20654), .C2(n20433), .A(n20653), .B(n20432), .ZN(
        n20450) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20450), .B1(
        n20481), .B2(n20657), .ZN(n20434) );
  OAI211_X1 U23455 ( .C1(n20660), .C2(n20453), .A(n20435), .B(n20434), .ZN(
        P1_U3105) );
  AOI22_X1 U23456 ( .A1(n20449), .A2(n20662), .B1(n20661), .B2(n20448), .ZN(
        n20437) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20450), .B1(
        n20481), .B2(n20663), .ZN(n20436) );
  OAI211_X1 U23458 ( .C1(n20666), .C2(n20453), .A(n20437), .B(n20436), .ZN(
        P1_U3106) );
  AOI22_X1 U23459 ( .A1(n20449), .A2(n20668), .B1(n20667), .B2(n20448), .ZN(
        n20439) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20450), .B1(
        n20481), .B2(n20669), .ZN(n20438) );
  OAI211_X1 U23461 ( .C1(n20672), .C2(n20453), .A(n20439), .B(n20438), .ZN(
        P1_U3107) );
  AOI22_X1 U23462 ( .A1(n20449), .A2(n20674), .B1(n20673), .B2(n20448), .ZN(
        n20441) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20450), .B1(
        n20481), .B2(n20675), .ZN(n20440) );
  OAI211_X1 U23464 ( .C1(n20678), .C2(n20453), .A(n20441), .B(n20440), .ZN(
        P1_U3108) );
  AOI22_X1 U23465 ( .A1(n20449), .A2(n20680), .B1(n20679), .B2(n20448), .ZN(
        n20443) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20450), .B1(
        n20481), .B2(n20681), .ZN(n20442) );
  OAI211_X1 U23467 ( .C1(n20684), .C2(n20453), .A(n20443), .B(n20442), .ZN(
        P1_U3109) );
  AOI22_X1 U23468 ( .A1(n20449), .A2(n20686), .B1(n20685), .B2(n20448), .ZN(
        n20445) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20450), .B1(
        n20481), .B2(n20687), .ZN(n20444) );
  OAI211_X1 U23470 ( .C1(n20690), .C2(n20453), .A(n20445), .B(n20444), .ZN(
        P1_U3110) );
  AOI22_X1 U23471 ( .A1(n20449), .A2(n20692), .B1(n20691), .B2(n20448), .ZN(
        n20447) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20450), .B1(
        n20481), .B2(n20693), .ZN(n20446) );
  OAI211_X1 U23473 ( .C1(n21073), .C2(n20453), .A(n20447), .B(n20446), .ZN(
        P1_U3111) );
  AOI22_X1 U23474 ( .A1(n20449), .A2(n20698), .B1(n20697), .B2(n20448), .ZN(
        n20452) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20450), .B1(
        n20481), .B2(n20700), .ZN(n20451) );
  OAI211_X1 U23476 ( .C1(n20706), .C2(n20453), .A(n20452), .B(n20451), .ZN(
        P1_U3112) );
  INV_X1 U23477 ( .A(n20481), .ZN(n20454) );
  NAND2_X1 U23478 ( .A1(n20454), .A2(n20654), .ZN(n20456) );
  OAI21_X1 U23479 ( .B1(n20456), .B2(n20512), .A(n20517), .ZN(n20463) );
  AND2_X1 U23480 ( .A1(n20490), .A2(n20598), .ZN(n20460) );
  OR2_X1 U23481 ( .A1(n20457), .A2(n20488), .ZN(n20600) );
  INV_X1 U23482 ( .A(n20600), .ZN(n20458) );
  NAND3_X1 U23483 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n12539), .ZN(n20491) );
  NOR2_X1 U23484 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20491), .ZN(
        n20480) );
  AOI22_X1 U23485 ( .A1(n20481), .A2(n20607), .B1(n20645), .B2(n20480), .ZN(
        n20467) );
  INV_X1 U23486 ( .A(n20460), .ZN(n20462) );
  INV_X1 U23487 ( .A(n20480), .ZN(n20461) );
  AOI22_X1 U23488 ( .A1(n20463), .A2(n20462), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20461), .ZN(n20464) );
  NAND2_X1 U23489 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20600), .ZN(n20604) );
  NAND3_X1 U23490 ( .A1(n20465), .A2(n20464), .A3(n20604), .ZN(n20482) );
  AOI22_X1 U23491 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20482), .B1(
        n20512), .B2(n20657), .ZN(n20466) );
  OAI211_X1 U23492 ( .C1(n20485), .C2(n20536), .A(n20467), .B(n20466), .ZN(
        P1_U3113) );
  AOI22_X1 U23493 ( .A1(n20481), .A2(n20611), .B1(n20661), .B2(n20480), .ZN(
        n20469) );
  AOI22_X1 U23494 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20482), .B1(
        n20512), .B2(n20663), .ZN(n20468) );
  OAI211_X1 U23495 ( .C1(n20485), .C2(n20541), .A(n20469), .B(n20468), .ZN(
        P1_U3114) );
  AOI22_X1 U23496 ( .A1(n20481), .A2(n20615), .B1(n20667), .B2(n20480), .ZN(
        n20471) );
  AOI22_X1 U23497 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20482), .B1(
        n20512), .B2(n20669), .ZN(n20470) );
  OAI211_X1 U23498 ( .C1(n20485), .C2(n20546), .A(n20471), .B(n20470), .ZN(
        P1_U3115) );
  AOI22_X1 U23499 ( .A1(n20481), .A2(n20619), .B1(n20673), .B2(n20480), .ZN(
        n20473) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20482), .B1(
        n20512), .B2(n20675), .ZN(n20472) );
  OAI211_X1 U23501 ( .C1(n20485), .C2(n20551), .A(n20473), .B(n20472), .ZN(
        P1_U3116) );
  AOI22_X1 U23502 ( .A1(n20512), .A2(n20681), .B1(n20679), .B2(n20480), .ZN(
        n20475) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20482), .B1(
        n20481), .B2(n20623), .ZN(n20474) );
  OAI211_X1 U23504 ( .C1(n20485), .C2(n20556), .A(n20475), .B(n20474), .ZN(
        P1_U3117) );
  AOI22_X1 U23505 ( .A1(n20481), .A2(n20627), .B1(n20685), .B2(n20480), .ZN(
        n20477) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20482), .B1(
        n20512), .B2(n20687), .ZN(n20476) );
  OAI211_X1 U23507 ( .C1(n20485), .C2(n20561), .A(n20477), .B(n20476), .ZN(
        P1_U3118) );
  AOI22_X1 U23508 ( .A1(n20512), .A2(n20693), .B1(n20691), .B2(n20480), .ZN(
        n20479) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20482), .B1(
        n20481), .B2(n20631), .ZN(n20478) );
  OAI211_X1 U23510 ( .C1(n20485), .C2(n21074), .A(n20479), .B(n20478), .ZN(
        P1_U3119) );
  AOI22_X1 U23511 ( .A1(n20481), .A2(n20636), .B1(n20697), .B2(n20480), .ZN(
        n20484) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20482), .B1(
        n20512), .B2(n20700), .ZN(n20483) );
  OAI211_X1 U23513 ( .C1(n20485), .C2(n20567), .A(n20484), .B(n20483), .ZN(
        P1_U3120) );
  NOR2_X1 U23514 ( .A1(n20489), .A2(n20488), .ZN(n20510) );
  AOI21_X1 U23515 ( .B1(n20490), .B2(n20642), .A(n20510), .ZN(n20492) );
  OAI22_X1 U23516 ( .A1(n20492), .A2(n20644), .B1(n20491), .B2(n11980), .ZN(
        n20511) );
  AOI22_X1 U23517 ( .A1(n20511), .A2(n20646), .B1(n20645), .B2(n20510), .ZN(
        n20497) );
  INV_X1 U23518 ( .A(n20491), .ZN(n20495) );
  OAI211_X1 U23519 ( .C1(n20493), .C2(n20650), .A(n20649), .B(n20492), .ZN(
        n20494) );
  OAI211_X1 U23520 ( .C1(n20649), .C2(n20495), .A(n20653), .B(n20494), .ZN(
        n20513) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20607), .ZN(n20496) );
  OAI211_X1 U23522 ( .C1(n20610), .C2(n21072), .A(n20497), .B(n20496), .ZN(
        P1_U3121) );
  AOI22_X1 U23523 ( .A1(n20511), .A2(n20662), .B1(n20661), .B2(n20510), .ZN(
        n20499) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20611), .ZN(n20498) );
  OAI211_X1 U23525 ( .C1(n20614), .C2(n21072), .A(n20499), .B(n20498), .ZN(
        P1_U3122) );
  AOI22_X1 U23526 ( .A1(n20511), .A2(n20668), .B1(n20667), .B2(n20510), .ZN(
        n20501) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20615), .ZN(n20500) );
  OAI211_X1 U23528 ( .C1(n20618), .C2(n21072), .A(n20501), .B(n20500), .ZN(
        P1_U3123) );
  AOI22_X1 U23529 ( .A1(n20511), .A2(n20674), .B1(n20673), .B2(n20510), .ZN(
        n20503) );
  AOI22_X1 U23530 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20619), .ZN(n20502) );
  OAI211_X1 U23531 ( .C1(n20622), .C2(n21072), .A(n20503), .B(n20502), .ZN(
        P1_U3124) );
  AOI22_X1 U23532 ( .A1(n20511), .A2(n20680), .B1(n20679), .B2(n20510), .ZN(
        n20505) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20623), .ZN(n20504) );
  OAI211_X1 U23534 ( .C1(n20626), .C2(n21072), .A(n20505), .B(n20504), .ZN(
        P1_U3125) );
  AOI22_X1 U23535 ( .A1(n20511), .A2(n20686), .B1(n20685), .B2(n20510), .ZN(
        n20507) );
  AOI22_X1 U23536 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20627), .ZN(n20506) );
  OAI211_X1 U23537 ( .C1(n20630), .C2(n21072), .A(n20507), .B(n20506), .ZN(
        P1_U3126) );
  AOI22_X1 U23538 ( .A1(n20511), .A2(n20692), .B1(n20691), .B2(n20510), .ZN(
        n20509) );
  AOI22_X1 U23539 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20631), .ZN(n20508) );
  OAI211_X1 U23540 ( .C1(n21070), .C2(n21072), .A(n20509), .B(n20508), .ZN(
        P1_U3127) );
  AOI22_X1 U23541 ( .A1(n20511), .A2(n20698), .B1(n20697), .B2(n20510), .ZN(
        n20515) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20513), .B1(
        n20512), .B2(n20636), .ZN(n20514) );
  OAI211_X1 U23543 ( .C1(n20641), .C2(n21072), .A(n20515), .B(n20514), .ZN(
        P1_U3128) );
  NAND3_X1 U23544 ( .A1(n21072), .A2(n20649), .A3(n21071), .ZN(n20518) );
  NAND2_X1 U23545 ( .A1(n20518), .A2(n20517), .ZN(n20530) );
  NOR2_X1 U23546 ( .A1(n20520), .A2(n20519), .ZN(n20643) );
  AND2_X1 U23547 ( .A1(n20643), .A2(n20521), .ZN(n20527) );
  NAND3_X1 U23548 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20524), .ZN(n20570) );
  NOR2_X1 U23549 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20570), .ZN(
        n20533) );
  INV_X1 U23550 ( .A(n20533), .ZN(n21068) );
  OAI22_X1 U23551 ( .A1(n21071), .A2(n20610), .B1(n20525), .B2(n21068), .ZN(
        n20526) );
  INV_X1 U23552 ( .A(n20526), .ZN(n20535) );
  INV_X1 U23553 ( .A(n20527), .ZN(n20529) );
  AOI22_X1 U23554 ( .A1(n20530), .A2(n20529), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20528), .ZN(n20531) );
  OAI211_X1 U23555 ( .C1(n20533), .C2(n20532), .A(n20605), .B(n20531), .ZN(
        n21078) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21078), .B1(
        n20564), .B2(n20607), .ZN(n20534) );
  OAI211_X1 U23557 ( .C1(n21075), .C2(n20536), .A(n20535), .B(n20534), .ZN(
        P1_U3129) );
  OAI22_X1 U23558 ( .A1(n21071), .A2(n20614), .B1(n20537), .B2(n21068), .ZN(
        n20538) );
  INV_X1 U23559 ( .A(n20538), .ZN(n20540) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21078), .B1(
        n20564), .B2(n20611), .ZN(n20539) );
  OAI211_X1 U23561 ( .C1(n21075), .C2(n20541), .A(n20540), .B(n20539), .ZN(
        P1_U3130) );
  OAI22_X1 U23562 ( .A1(n21071), .A2(n20618), .B1(n20542), .B2(n21068), .ZN(
        n20543) );
  INV_X1 U23563 ( .A(n20543), .ZN(n20545) );
  AOI22_X1 U23564 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21078), .B1(
        n20564), .B2(n20615), .ZN(n20544) );
  OAI211_X1 U23565 ( .C1(n21075), .C2(n20546), .A(n20545), .B(n20544), .ZN(
        P1_U3131) );
  OAI22_X1 U23566 ( .A1(n21071), .A2(n20622), .B1(n20547), .B2(n21068), .ZN(
        n20548) );
  INV_X1 U23567 ( .A(n20548), .ZN(n20550) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21078), .B1(
        n20564), .B2(n20619), .ZN(n20549) );
  OAI211_X1 U23569 ( .C1(n21075), .C2(n20551), .A(n20550), .B(n20549), .ZN(
        P1_U3132) );
  OAI22_X1 U23570 ( .A1(n21071), .A2(n20626), .B1(n20552), .B2(n21068), .ZN(
        n20553) );
  INV_X1 U23571 ( .A(n20553), .ZN(n20555) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21078), .B1(
        n20564), .B2(n20623), .ZN(n20554) );
  OAI211_X1 U23573 ( .C1(n21075), .C2(n20556), .A(n20555), .B(n20554), .ZN(
        P1_U3133) );
  OAI22_X1 U23574 ( .A1(n21071), .A2(n20630), .B1(n20557), .B2(n21068), .ZN(
        n20558) );
  INV_X1 U23575 ( .A(n20558), .ZN(n20560) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21078), .B1(
        n20564), .B2(n20627), .ZN(n20559) );
  OAI211_X1 U23577 ( .C1(n21075), .C2(n20561), .A(n20560), .B(n20559), .ZN(
        P1_U3134) );
  OAI22_X1 U23578 ( .A1(n21071), .A2(n20641), .B1(n20562), .B2(n21068), .ZN(
        n20563) );
  INV_X1 U23579 ( .A(n20563), .ZN(n20566) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21078), .B1(
        n20564), .B2(n20636), .ZN(n20565) );
  OAI211_X1 U23581 ( .C1(n21075), .C2(n20567), .A(n20566), .B(n20565), .ZN(
        P1_U3136) );
  NOR2_X1 U23582 ( .A1(n20568), .A2(n20570), .ZN(n20591) );
  AOI21_X1 U23583 ( .B1(n20643), .B2(n20569), .A(n20591), .ZN(n20572) );
  OAI22_X1 U23584 ( .A1(n20572), .A2(n20644), .B1(n20570), .B2(n11980), .ZN(
        n20592) );
  AOI22_X1 U23585 ( .A1(n20592), .A2(n20646), .B1(n20645), .B2(n20591), .ZN(
        n20578) );
  INV_X1 U23586 ( .A(n20570), .ZN(n20575) );
  INV_X1 U23587 ( .A(n20571), .ZN(n20573) );
  NAND2_X1 U23588 ( .A1(n20573), .A2(n20572), .ZN(n20574) );
  OAI221_X1 U23589 ( .B1(n20654), .B2(n20575), .C1(n20644), .C2(n20574), .A(
        n20653), .ZN(n20593) );
  NOR2_X2 U23590 ( .A1(n20651), .A2(n20576), .ZN(n20637) );
  AOI22_X1 U23591 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20593), .B1(
        n20637), .B2(n20657), .ZN(n20577) );
  OAI211_X1 U23592 ( .C1(n20660), .C2(n21071), .A(n20578), .B(n20577), .ZN(
        P1_U3137) );
  AOI22_X1 U23593 ( .A1(n20592), .A2(n20662), .B1(n20661), .B2(n20591), .ZN(
        n20580) );
  AOI22_X1 U23594 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20593), .B1(
        n20637), .B2(n20663), .ZN(n20579) );
  OAI211_X1 U23595 ( .C1(n20666), .C2(n21071), .A(n20580), .B(n20579), .ZN(
        P1_U3138) );
  AOI22_X1 U23596 ( .A1(n20592), .A2(n20668), .B1(n20667), .B2(n20591), .ZN(
        n20582) );
  AOI22_X1 U23597 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20593), .B1(
        n20637), .B2(n20669), .ZN(n20581) );
  OAI211_X1 U23598 ( .C1(n20672), .C2(n21071), .A(n20582), .B(n20581), .ZN(
        P1_U3139) );
  AOI22_X1 U23599 ( .A1(n20592), .A2(n20674), .B1(n20673), .B2(n20591), .ZN(
        n20584) );
  AOI22_X1 U23600 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20593), .B1(
        n20637), .B2(n20675), .ZN(n20583) );
  OAI211_X1 U23601 ( .C1(n20678), .C2(n21071), .A(n20584), .B(n20583), .ZN(
        P1_U3140) );
  AOI22_X1 U23602 ( .A1(n20592), .A2(n20680), .B1(n20679), .B2(n20591), .ZN(
        n20586) );
  AOI22_X1 U23603 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20593), .B1(
        n20637), .B2(n20681), .ZN(n20585) );
  OAI211_X1 U23604 ( .C1(n20684), .C2(n21071), .A(n20586), .B(n20585), .ZN(
        P1_U3141) );
  AOI22_X1 U23605 ( .A1(n20592), .A2(n20686), .B1(n20685), .B2(n20591), .ZN(
        n20588) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20593), .B1(
        n20637), .B2(n20687), .ZN(n20587) );
  OAI211_X1 U23607 ( .C1(n20690), .C2(n21071), .A(n20588), .B(n20587), .ZN(
        P1_U3142) );
  AOI22_X1 U23608 ( .A1(n20592), .A2(n20692), .B1(n20691), .B2(n20591), .ZN(
        n20590) );
  AOI22_X1 U23609 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20593), .B1(
        n20637), .B2(n20693), .ZN(n20589) );
  OAI211_X1 U23610 ( .C1(n21073), .C2(n21071), .A(n20590), .B(n20589), .ZN(
        P1_U3143) );
  AOI22_X1 U23611 ( .A1(n20592), .A2(n20698), .B1(n20697), .B2(n20591), .ZN(
        n20595) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20593), .B1(
        n20637), .B2(n20700), .ZN(n20594) );
  OAI211_X1 U23613 ( .C1(n20706), .C2(n21071), .A(n20595), .B(n20594), .ZN(
        P1_U3144) );
  INV_X1 U23614 ( .A(n20651), .ZN(n20597) );
  NAND2_X1 U23615 ( .A1(n20643), .A2(n20598), .ZN(n20602) );
  OAI22_X1 U23616 ( .A1(n20602), .A2(n20644), .B1(n20600), .B2(n20599), .ZN(
        n20635) );
  NOR2_X1 U23617 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20647), .ZN(
        n20634) );
  AOI22_X1 U23618 ( .A1(n20635), .A2(n20646), .B1(n20645), .B2(n20634), .ZN(
        n20609) );
  INV_X1 U23619 ( .A(n20705), .ZN(n20601) );
  OAI21_X1 U23620 ( .B1(n20601), .B2(n20637), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20603) );
  AOI21_X1 U23621 ( .B1(n20603), .B2(n20602), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20606) );
  AOI22_X1 U23622 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20607), .ZN(n20608) );
  OAI211_X1 U23623 ( .C1(n20610), .C2(n20705), .A(n20609), .B(n20608), .ZN(
        P1_U3145) );
  AOI22_X1 U23624 ( .A1(n20635), .A2(n20662), .B1(n20661), .B2(n20634), .ZN(
        n20613) );
  AOI22_X1 U23625 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20611), .ZN(n20612) );
  OAI211_X1 U23626 ( .C1(n20614), .C2(n20705), .A(n20613), .B(n20612), .ZN(
        P1_U3146) );
  AOI22_X1 U23627 ( .A1(n20635), .A2(n20668), .B1(n20667), .B2(n20634), .ZN(
        n20617) );
  AOI22_X1 U23628 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20615), .ZN(n20616) );
  OAI211_X1 U23629 ( .C1(n20618), .C2(n20705), .A(n20617), .B(n20616), .ZN(
        P1_U3147) );
  AOI22_X1 U23630 ( .A1(n20635), .A2(n20674), .B1(n20673), .B2(n20634), .ZN(
        n20621) );
  AOI22_X1 U23631 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20619), .ZN(n20620) );
  OAI211_X1 U23632 ( .C1(n20622), .C2(n20705), .A(n20621), .B(n20620), .ZN(
        P1_U3148) );
  AOI22_X1 U23633 ( .A1(n20635), .A2(n20680), .B1(n20679), .B2(n20634), .ZN(
        n20625) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20623), .ZN(n20624) );
  OAI211_X1 U23635 ( .C1(n20626), .C2(n20705), .A(n20625), .B(n20624), .ZN(
        P1_U3149) );
  AOI22_X1 U23636 ( .A1(n20635), .A2(n20686), .B1(n20685), .B2(n20634), .ZN(
        n20629) );
  AOI22_X1 U23637 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20627), .ZN(n20628) );
  OAI211_X1 U23638 ( .C1(n20630), .C2(n20705), .A(n20629), .B(n20628), .ZN(
        P1_U3150) );
  AOI22_X1 U23639 ( .A1(n20635), .A2(n20692), .B1(n20691), .B2(n20634), .ZN(
        n20633) );
  AOI22_X1 U23640 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20631), .ZN(n20632) );
  OAI211_X1 U23641 ( .C1(n21070), .C2(n20705), .A(n20633), .B(n20632), .ZN(
        P1_U3151) );
  AOI22_X1 U23642 ( .A1(n20635), .A2(n20698), .B1(n20697), .B2(n20634), .ZN(
        n20640) );
  AOI22_X1 U23643 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20638), .B1(
        n20637), .B2(n20636), .ZN(n20639) );
  OAI211_X1 U23644 ( .C1(n20641), .C2(n20705), .A(n20640), .B(n20639), .ZN(
        P1_U3152) );
  AOI21_X1 U23645 ( .B1(n20643), .B2(n20642), .A(n20696), .ZN(n20648) );
  OAI22_X1 U23646 ( .A1(n20648), .A2(n20644), .B1(n20647), .B2(n11980), .ZN(
        n20699) );
  AOI22_X1 U23647 ( .A1(n20699), .A2(n20646), .B1(n20645), .B2(n20696), .ZN(
        n20659) );
  INV_X1 U23648 ( .A(n20647), .ZN(n20655) );
  OAI211_X1 U23649 ( .C1(n20651), .C2(n20650), .A(n20649), .B(n20648), .ZN(
        n20652) );
  OAI211_X1 U23650 ( .C1(n20655), .C2(n20654), .A(n20653), .B(n20652), .ZN(
        n20702) );
  AOI22_X1 U23651 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20702), .B1(
        n20701), .B2(n20657), .ZN(n20658) );
  OAI211_X1 U23652 ( .C1(n20660), .C2(n20705), .A(n20659), .B(n20658), .ZN(
        P1_U3153) );
  AOI22_X1 U23653 ( .A1(n20699), .A2(n20662), .B1(n20661), .B2(n20696), .ZN(
        n20665) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20702), .B1(
        n20701), .B2(n20663), .ZN(n20664) );
  OAI211_X1 U23655 ( .C1(n20666), .C2(n20705), .A(n20665), .B(n20664), .ZN(
        P1_U3154) );
  AOI22_X1 U23656 ( .A1(n20699), .A2(n20668), .B1(n20667), .B2(n20696), .ZN(
        n20671) );
  AOI22_X1 U23657 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20702), .B1(
        n20701), .B2(n20669), .ZN(n20670) );
  OAI211_X1 U23658 ( .C1(n20672), .C2(n20705), .A(n20671), .B(n20670), .ZN(
        P1_U3155) );
  AOI22_X1 U23659 ( .A1(n20699), .A2(n20674), .B1(n20673), .B2(n20696), .ZN(
        n20677) );
  AOI22_X1 U23660 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20702), .B1(
        n20701), .B2(n20675), .ZN(n20676) );
  OAI211_X1 U23661 ( .C1(n20678), .C2(n20705), .A(n20677), .B(n20676), .ZN(
        P1_U3156) );
  AOI22_X1 U23662 ( .A1(n20699), .A2(n20680), .B1(n20679), .B2(n20696), .ZN(
        n20683) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20702), .B1(
        n20701), .B2(n20681), .ZN(n20682) );
  OAI211_X1 U23664 ( .C1(n20684), .C2(n20705), .A(n20683), .B(n20682), .ZN(
        P1_U3157) );
  AOI22_X1 U23665 ( .A1(n20699), .A2(n20686), .B1(n20685), .B2(n20696), .ZN(
        n20689) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20702), .B1(
        n20701), .B2(n20687), .ZN(n20688) );
  OAI211_X1 U23667 ( .C1(n20690), .C2(n20705), .A(n20689), .B(n20688), .ZN(
        P1_U3158) );
  AOI22_X1 U23668 ( .A1(n20699), .A2(n20692), .B1(n20691), .B2(n20696), .ZN(
        n20695) );
  AOI22_X1 U23669 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20702), .B1(
        n20701), .B2(n20693), .ZN(n20694) );
  OAI211_X1 U23670 ( .C1(n21073), .C2(n20705), .A(n20695), .B(n20694), .ZN(
        P1_U3159) );
  AOI22_X1 U23671 ( .A1(n20699), .A2(n20698), .B1(n20697), .B2(n20696), .ZN(
        n20704) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20702), .B1(
        n20701), .B2(n20700), .ZN(n20703) );
  OAI211_X1 U23673 ( .C1(n20706), .C2(n20705), .A(n20704), .B(n20703), .ZN(
        P1_U3160) );
  NOR2_X1 U23674 ( .A1(n20708), .A2(n20707), .ZN(n20711) );
  OAI21_X1 U23675 ( .B1(n20711), .B2(n11980), .A(n20709), .ZN(P1_U3163) );
  AND2_X1 U23676 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20783), .ZN(
        P1_U3164) );
  INV_X1 U23677 ( .A(P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n21021) );
  NOR2_X1 U23678 ( .A1(n20786), .A2(n21021), .ZN(P1_U3165) );
  AND2_X1 U23679 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20783), .ZN(
        P1_U3166) );
  AND2_X1 U23680 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20783), .ZN(
        P1_U3167) );
  AND2_X1 U23681 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20783), .ZN(
        P1_U3168) );
  AND2_X1 U23682 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20783), .ZN(
        P1_U3169) );
  AND2_X1 U23683 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20783), .ZN(
        P1_U3170) );
  AND2_X1 U23684 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20783), .ZN(
        P1_U3171) );
  AND2_X1 U23685 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20783), .ZN(
        P1_U3172) );
  AND2_X1 U23686 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20783), .ZN(
        P1_U3173) );
  AND2_X1 U23687 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20783), .ZN(
        P1_U3174) );
  AND2_X1 U23688 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20783), .ZN(
        P1_U3175) );
  AND2_X1 U23689 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20783), .ZN(
        P1_U3176) );
  AND2_X1 U23690 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20783), .ZN(
        P1_U3177) );
  AND2_X1 U23691 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20783), .ZN(
        P1_U3178) );
  AND2_X1 U23692 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20783), .ZN(
        P1_U3179) );
  AND2_X1 U23693 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20783), .ZN(
        P1_U3180) );
  AND2_X1 U23694 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20783), .ZN(
        P1_U3181) );
  AND2_X1 U23695 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20783), .ZN(
        P1_U3182) );
  AND2_X1 U23696 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20783), .ZN(
        P1_U3183) );
  AND2_X1 U23697 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20783), .ZN(
        P1_U3184) );
  AND2_X1 U23698 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20783), .ZN(
        P1_U3185) );
  AND2_X1 U23699 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20783), .ZN(P1_U3186) );
  AND2_X1 U23700 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20783), .ZN(P1_U3187) );
  AND2_X1 U23701 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20783), .ZN(P1_U3188) );
  INV_X1 U23702 ( .A(P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20910) );
  NOR2_X1 U23703 ( .A1(n20786), .A2(n20910), .ZN(P1_U3189) );
  AND2_X1 U23704 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20783), .ZN(P1_U3190) );
  AND2_X1 U23705 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20783), .ZN(P1_U3191) );
  AND2_X1 U23706 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20783), .ZN(P1_U3192) );
  AND2_X1 U23707 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20783), .ZN(P1_U3193) );
  NAND2_X1 U23708 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20716), .ZN(n20721) );
  INV_X1 U23709 ( .A(n20721), .ZN(n20715) );
  OAI21_X1 U23710 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20722), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20712) );
  AOI211_X1 U23711 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20713), .B(
        n20712), .ZN(n20714) );
  OAI22_X1 U23712 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20715), .B1(n20809), 
        .B2(n20714), .ZN(P1_U3194) );
  NOR3_X1 U23713 ( .A1(NA), .A2(n12961), .A3(n20716), .ZN(n20720) );
  AOI21_X1 U23714 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20877), .A(n20717), .ZN(n20719) );
  AOI222_X1 U23715 ( .A1(n20720), .A2(n20719), .B1(n20720), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .C1(n20719), .C2(n20718), .ZN(n20724)
         );
  OAI211_X1 U23716 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20722), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20721), .ZN(n20723) );
  NAND2_X1 U23717 ( .A1(n20724), .A2(n20723), .ZN(P1_U3196) );
  NAND2_X1 U23718 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20809), .ZN(n20771) );
  NAND2_X1 U23719 ( .A1(n20809), .A2(n20877), .ZN(n20775) );
  OAI222_X1 U23720 ( .A1(n20771), .A2(n20788), .B1(n20725), .B2(n20809), .C1(
        n20923), .C2(n20775), .ZN(P1_U3197) );
  INV_X1 U23721 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20726) );
  OAI222_X1 U23722 ( .A1(n20771), .A2(n20923), .B1(n20726), .B2(n20809), .C1(
        n20728), .C2(n20775), .ZN(P1_U3198) );
  INV_X1 U23723 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20727) );
  OAI222_X1 U23724 ( .A1(n20771), .A2(n20728), .B1(n20727), .B2(n20809), .C1(
        n20729), .C2(n20775), .ZN(P1_U3199) );
  INV_X1 U23725 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20730) );
  OAI222_X1 U23726 ( .A1(n20775), .A2(n20731), .B1(n20730), .B2(n20809), .C1(
        n20729), .C2(n20771), .ZN(P1_U3200) );
  INV_X1 U23727 ( .A(n20771), .ZN(n20773) );
  INV_X1 U23728 ( .A(n20775), .ZN(n20769) );
  AOI222_X1 U23729 ( .A1(n20773), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20794), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20769), .ZN(n20732) );
  INV_X1 U23730 ( .A(n20732), .ZN(P1_U3201) );
  AOI222_X1 U23731 ( .A1(n20773), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20794), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20769), .ZN(n20733) );
  INV_X1 U23732 ( .A(n20733), .ZN(P1_U3202) );
  INV_X1 U23733 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n20734) );
  OAI222_X1 U23734 ( .A1(n20771), .A2(n20735), .B1(n20734), .B2(n20809), .C1(
        n20737), .C2(n20775), .ZN(P1_U3203) );
  INV_X1 U23735 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n20736) );
  OAI222_X1 U23736 ( .A1(n20771), .A2(n20737), .B1(n20736), .B2(n20809), .C1(
        n20946), .C2(n20775), .ZN(P1_U3204) );
  INV_X1 U23737 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20738) );
  OAI222_X1 U23738 ( .A1(n20775), .A2(n21000), .B1(n20738), .B2(n20809), .C1(
        n20946), .C2(n20771), .ZN(P1_U3205) );
  INV_X1 U23739 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20739) );
  OAI222_X1 U23740 ( .A1(n20775), .A2(n15754), .B1(n20739), .B2(n20809), .C1(
        n21000), .C2(n20771), .ZN(P1_U3206) );
  INV_X1 U23741 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20740) );
  OAI222_X1 U23742 ( .A1(n20775), .A2(n20741), .B1(n20740), .B2(n20809), .C1(
        n15754), .C2(n20771), .ZN(P1_U3207) );
  INV_X1 U23743 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20742) );
  OAI222_X1 U23744 ( .A1(n20775), .A2(n20744), .B1(n20742), .B2(n20809), .C1(
        n20741), .C2(n20771), .ZN(P1_U3208) );
  AOI22_X1 U23745 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20794), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20769), .ZN(n20743) );
  OAI21_X1 U23746 ( .B1(n20744), .B2(n20771), .A(n20743), .ZN(P1_U3209) );
  INV_X1 U23747 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20746) );
  AOI22_X1 U23748 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20794), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20773), .ZN(n20745) );
  OAI21_X1 U23749 ( .B1(n20746), .B2(n20775), .A(n20745), .ZN(P1_U3210) );
  INV_X1 U23750 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20985) );
  OAI222_X1 U23751 ( .A1(n20771), .A2(n20746), .B1(n20985), .B2(n20809), .C1(
        n20748), .C2(n20775), .ZN(P1_U3211) );
  INV_X1 U23752 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20747) );
  OAI222_X1 U23753 ( .A1(n20771), .A2(n20748), .B1(n20747), .B2(n20809), .C1(
        n20749), .C2(n20775), .ZN(P1_U3212) );
  INV_X1 U23754 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20750) );
  OAI222_X1 U23755 ( .A1(n20775), .A2(n20752), .B1(n20750), .B2(n20809), .C1(
        n20749), .C2(n20771), .ZN(P1_U3213) );
  AOI22_X1 U23756 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20794), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20769), .ZN(n20751) );
  OAI21_X1 U23757 ( .B1(n20752), .B2(n20771), .A(n20751), .ZN(P1_U3214) );
  AOI22_X1 U23758 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20794), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20773), .ZN(n20753) );
  OAI21_X1 U23759 ( .B1(n20754), .B2(n20775), .A(n20753), .ZN(P1_U3215) );
  INV_X1 U23760 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n20755) );
  OAI222_X1 U23761 ( .A1(n20775), .A2(n20757), .B1(n20755), .B2(n20809), .C1(
        n20754), .C2(n20771), .ZN(P1_U3216) );
  INV_X1 U23762 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n20756) );
  OAI222_X1 U23763 ( .A1(n20771), .A2(n20757), .B1(n20756), .B2(n20809), .C1(
        n20759), .C2(n20775), .ZN(P1_U3217) );
  AOI22_X1 U23764 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20794), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20769), .ZN(n20758) );
  OAI21_X1 U23765 ( .B1(n20759), .B2(n20771), .A(n20758), .ZN(P1_U3218) );
  AOI22_X1 U23766 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20794), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20773), .ZN(n20760) );
  OAI21_X1 U23767 ( .B1(n20762), .B2(n20775), .A(n20760), .ZN(P1_U3219) );
  INV_X1 U23768 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20761) );
  OAI222_X1 U23769 ( .A1(n20771), .A2(n20762), .B1(n20761), .B2(n20809), .C1(
        n20764), .C2(n20775), .ZN(P1_U3220) );
  AOI22_X1 U23770 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n20769), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20794), .ZN(n20763) );
  OAI21_X1 U23771 ( .B1(n20764), .B2(n20771), .A(n20763), .ZN(P1_U3221) );
  AOI22_X1 U23772 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n20773), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20794), .ZN(n20765) );
  OAI21_X1 U23773 ( .B1(n20766), .B2(n20775), .A(n20765), .ZN(P1_U3222) );
  AOI222_X1 U23774 ( .A1(n20773), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20794), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20769), .ZN(n20767) );
  INV_X1 U23775 ( .A(n20767), .ZN(P1_U3223) );
  AOI222_X1 U23776 ( .A1(n20773), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20794), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20769), .ZN(n20768) );
  INV_X1 U23777 ( .A(n20768), .ZN(P1_U3224) );
  AOI22_X1 U23778 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20769), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20794), .ZN(n20770) );
  OAI21_X1 U23779 ( .B1(n20772), .B2(n20771), .A(n20770), .ZN(P1_U3225) );
  AOI22_X1 U23780 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20773), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20794), .ZN(n20774) );
  OAI21_X1 U23781 ( .B1(n20776), .B2(n20775), .A(n20774), .ZN(P1_U3226) );
  INV_X1 U23782 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20777) );
  AOI22_X1 U23783 ( .A1(n20809), .A2(n20778), .B1(n20777), .B2(n20794), .ZN(
        P1_U3458) );
  INV_X1 U23784 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20816) );
  INV_X1 U23785 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20779) );
  AOI22_X1 U23786 ( .A1(n20809), .A2(n20816), .B1(n20779), .B2(n20794), .ZN(
        P1_U3459) );
  INV_X1 U23787 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20780) );
  AOI22_X1 U23788 ( .A1(n20809), .A2(n20781), .B1(n20780), .B2(n20794), .ZN(
        P1_U3460) );
  INV_X1 U23789 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20791) );
  AOI22_X1 U23790 ( .A1(n20809), .A2(n20791), .B1(n20962), .B2(n20794), .ZN(
        P1_U3461) );
  INV_X1 U23791 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21022) );
  INV_X1 U23792 ( .A(n20784), .ZN(n20782) );
  AOI21_X1 U23793 ( .B1(n21022), .B2(n20783), .A(n20782), .ZN(P1_U3464) );
  OAI21_X1 U23794 ( .B1(n20786), .B2(n20785), .A(n20784), .ZN(P1_U3465) );
  AOI21_X1 U23795 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20787) );
  OAI22_X1 U23796 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(n20788), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(n20787), .ZN(n20789) );
  AOI22_X1 U23797 ( .A1(n20793), .A2(n20789), .B1(n20816), .B2(n20790), .ZN(
        P1_U3481) );
  NOR2_X1 U23798 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20792) );
  AOI22_X1 U23799 ( .A1(n20793), .A2(n20792), .B1(n20791), .B2(n20790), .ZN(
        P1_U3482) );
  INV_X1 U23800 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20795) );
  AOI22_X1 U23801 ( .A1(n20809), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20795), 
        .B2(n20794), .ZN(P1_U3483) );
  INV_X1 U23802 ( .A(n20796), .ZN(n20797) );
  OAI211_X1 U23803 ( .C1(n20800), .C2(n20799), .A(n20798), .B(n20797), .ZN(
        n20808) );
  INV_X1 U23804 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20807) );
  NOR2_X1 U23805 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20801), .ZN(n20806) );
  OAI211_X1 U23806 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20803), .A(n20802), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20804) );
  NAND2_X1 U23807 ( .A1(n20808), .A2(n20804), .ZN(n20805) );
  OAI22_X1 U23808 ( .A1(n20808), .A2(n20807), .B1(n20806), .B2(n20805), .ZN(
        P1_U3485) );
  MUX2_X1 U23809 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n20809), .Z(P1_U3486) );
  AOI22_X1 U23810 ( .A1(n14312), .A2(keyinput81), .B1(keyinput77), .B2(n20811), 
        .ZN(n20810) );
  OAI221_X1 U23811 ( .B1(n14312), .B2(keyinput81), .C1(n20811), .C2(keyinput77), .A(n20810), .ZN(n20824) );
  AOI22_X1 U23812 ( .A1(n20814), .A2(keyinput91), .B1(n20813), .B2(keyinput65), 
        .ZN(n20812) );
  OAI221_X1 U23813 ( .B1(n20814), .B2(keyinput91), .C1(n20813), .C2(keyinput65), .A(n20812), .ZN(n20823) );
  AOI22_X1 U23814 ( .A1(n20817), .A2(keyinput56), .B1(n20816), .B2(keyinput101), .ZN(n20815) );
  OAI221_X1 U23815 ( .B1(n20817), .B2(keyinput56), .C1(n20816), .C2(
        keyinput101), .A(n20815), .ZN(n20822) );
  AOI22_X1 U23816 ( .A1(n20820), .A2(keyinput39), .B1(n20819), .B2(keyinput124), .ZN(n20818) );
  OAI221_X1 U23817 ( .B1(n20820), .B2(keyinput39), .C1(n20819), .C2(
        keyinput124), .A(n20818), .ZN(n20821) );
  NOR4_X1 U23818 ( .A1(n20824), .A2(n20823), .A3(n20822), .A4(n20821), .ZN(
        n20872) );
  AOI22_X1 U23819 ( .A1(n20827), .A2(keyinput100), .B1(keyinput63), .B2(n20826), .ZN(n20825) );
  OAI221_X1 U23820 ( .B1(n20827), .B2(keyinput100), .C1(n20826), .C2(
        keyinput63), .A(n20825), .ZN(n20838) );
  AOI22_X1 U23821 ( .A1(n20829), .A2(keyinput117), .B1(n21105), .B2(keyinput6), 
        .ZN(n20828) );
  OAI221_X1 U23822 ( .B1(n20829), .B2(keyinput117), .C1(n21105), .C2(keyinput6), .A(n20828), .ZN(n20837) );
  AOI22_X1 U23823 ( .A1(n20832), .A2(keyinput60), .B1(keyinput10), .B2(n20831), 
        .ZN(n20830) );
  OAI221_X1 U23824 ( .B1(n20832), .B2(keyinput60), .C1(n20831), .C2(keyinput10), .A(n20830), .ZN(n20836) );
  AOI22_X1 U23825 ( .A1(n11294), .A2(keyinput76), .B1(n20834), .B2(keyinput52), 
        .ZN(n20833) );
  OAI221_X1 U23826 ( .B1(n11294), .B2(keyinput76), .C1(n20834), .C2(keyinput52), .A(n20833), .ZN(n20835) );
  NOR4_X1 U23827 ( .A1(n20838), .A2(n20837), .A3(n20836), .A4(n20835), .ZN(
        n20871) );
  AOI22_X1 U23828 ( .A1(n20841), .A2(keyinput47), .B1(n20840), .B2(keyinput127), .ZN(n20839) );
  OAI221_X1 U23829 ( .B1(n20841), .B2(keyinput47), .C1(n20840), .C2(
        keyinput127), .A(n20839), .ZN(n20845) );
  XOR2_X1 U23830 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B(keyinput27), .Z(
        n20844) );
  XNOR2_X1 U23831 ( .A(n20842), .B(keyinput66), .ZN(n20843) );
  OR3_X1 U23832 ( .A1(n20845), .A2(n20844), .A3(n20843), .ZN(n20853) );
  AOI22_X1 U23833 ( .A1(n20848), .A2(keyinput83), .B1(keyinput49), .B2(n20847), 
        .ZN(n20846) );
  OAI221_X1 U23834 ( .B1(n20848), .B2(keyinput83), .C1(n20847), .C2(keyinput49), .A(n20846), .ZN(n20852) );
  AOI22_X1 U23835 ( .A1(n21079), .A2(keyinput105), .B1(keyinput119), .B2(
        n20850), .ZN(n20849) );
  OAI221_X1 U23836 ( .B1(n21079), .B2(keyinput105), .C1(n20850), .C2(
        keyinput119), .A(n20849), .ZN(n20851) );
  NOR3_X1 U23837 ( .A1(n20853), .A2(n20852), .A3(n20851), .ZN(n20870) );
  AOI22_X1 U23838 ( .A1(n20856), .A2(keyinput4), .B1(keyinput78), .B2(n20855), 
        .ZN(n20854) );
  OAI221_X1 U23839 ( .B1(n20856), .B2(keyinput4), .C1(n20855), .C2(keyinput78), 
        .A(n20854), .ZN(n20868) );
  AOI22_X1 U23840 ( .A1(n15754), .A2(keyinput1), .B1(keyinput42), .B2(n20858), 
        .ZN(n20857) );
  OAI221_X1 U23841 ( .B1(n15754), .B2(keyinput1), .C1(n20858), .C2(keyinput42), 
        .A(n20857), .ZN(n20867) );
  INV_X1 U23842 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n20861) );
  AOI22_X1 U23843 ( .A1(n20861), .A2(keyinput46), .B1(n20860), .B2(keyinput51), 
        .ZN(n20859) );
  OAI221_X1 U23844 ( .B1(n20861), .B2(keyinput46), .C1(n20860), .C2(keyinput51), .A(n20859), .ZN(n20866) );
  INV_X1 U23845 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n20863) );
  AOI22_X1 U23846 ( .A1(n20864), .A2(keyinput98), .B1(n20863), .B2(keyinput26), 
        .ZN(n20862) );
  OAI221_X1 U23847 ( .B1(n20864), .B2(keyinput98), .C1(n20863), .C2(keyinput26), .A(n20862), .ZN(n20865) );
  NOR4_X1 U23848 ( .A1(n20868), .A2(n20867), .A3(n20866), .A4(n20865), .ZN(
        n20869) );
  NAND4_X1 U23849 ( .A1(n20872), .A2(n20871), .A3(n20870), .A4(n20869), .ZN(
        n21067) );
  AOI22_X1 U23850 ( .A1(n9963), .A2(keyinput48), .B1(keyinput115), .B2(n20874), 
        .ZN(n20873) );
  OAI221_X1 U23851 ( .B1(n9963), .B2(keyinput48), .C1(n20874), .C2(keyinput115), .A(n20873), .ZN(n20886) );
  AOI22_X1 U23852 ( .A1(n20877), .A2(keyinput29), .B1(keyinput94), .B2(n20876), 
        .ZN(n20875) );
  OAI221_X1 U23853 ( .B1(n20877), .B2(keyinput29), .C1(n20876), .C2(keyinput94), .A(n20875), .ZN(n20885) );
  AOI22_X1 U23854 ( .A1(n20879), .A2(keyinput41), .B1(keyinput113), .B2(n14610), .ZN(n20878) );
  OAI221_X1 U23855 ( .B1(n20879), .B2(keyinput41), .C1(n14610), .C2(
        keyinput113), .A(n20878), .ZN(n20884) );
  AOI22_X1 U23856 ( .A1(n20882), .A2(keyinput30), .B1(n20881), .B2(keyinput71), 
        .ZN(n20880) );
  OAI221_X1 U23857 ( .B1(n20882), .B2(keyinput30), .C1(n20881), .C2(keyinput71), .A(n20880), .ZN(n20883) );
  NOR4_X1 U23858 ( .A1(n20886), .A2(n20885), .A3(n20884), .A4(n20883), .ZN(
        n20935) );
  AOI22_X1 U23859 ( .A1(n20888), .A2(keyinput104), .B1(n21088), .B2(keyinput12), .ZN(n20887) );
  OAI221_X1 U23860 ( .B1(n20888), .B2(keyinput104), .C1(n21088), .C2(
        keyinput12), .A(n20887), .ZN(n20900) );
  INV_X1 U23861 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U23862 ( .A1(n20890), .A2(keyinput13), .B1(n21107), .B2(keyinput54), 
        .ZN(n20889) );
  OAI221_X1 U23863 ( .B1(n20890), .B2(keyinput13), .C1(n21107), .C2(keyinput54), .A(n20889), .ZN(n20899) );
  INV_X1 U23864 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U23865 ( .A1(n20893), .A2(keyinput79), .B1(keyinput57), .B2(n20892), 
        .ZN(n20891) );
  OAI221_X1 U23866 ( .B1(n20893), .B2(keyinput79), .C1(n20892), .C2(keyinput57), .A(n20891), .ZN(n20898) );
  AOI22_X1 U23867 ( .A1(n20896), .A2(keyinput7), .B1(keyinput67), .B2(n20895), 
        .ZN(n20894) );
  OAI221_X1 U23868 ( .B1(n20896), .B2(keyinput7), .C1(n20895), .C2(keyinput67), 
        .A(n20894), .ZN(n20897) );
  NOR4_X1 U23869 ( .A1(n20900), .A2(n20899), .A3(n20898), .A4(n20897), .ZN(
        n20934) );
  AOI22_X1 U23870 ( .A1(n20903), .A2(keyinput31), .B1(n20902), .B2(keyinput8), 
        .ZN(n20901) );
  OAI221_X1 U23871 ( .B1(n20903), .B2(keyinput31), .C1(n20902), .C2(keyinput8), 
        .A(n20901), .ZN(n20907) );
  XOR2_X1 U23872 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B(keyinput85), .Z(
        n20906) );
  XNOR2_X1 U23873 ( .A(n20904), .B(keyinput24), .ZN(n20905) );
  OR3_X1 U23874 ( .A1(n20907), .A2(n20906), .A3(n20905), .ZN(n20916) );
  AOI22_X1 U23875 ( .A1(n20910), .A2(keyinput86), .B1(n20909), .B2(keyinput43), 
        .ZN(n20908) );
  OAI221_X1 U23876 ( .B1(n20910), .B2(keyinput86), .C1(n20909), .C2(keyinput43), .A(n20908), .ZN(n20915) );
  AOI22_X1 U23877 ( .A1(n20913), .A2(keyinput40), .B1(n20912), .B2(keyinput72), 
        .ZN(n20911) );
  OAI221_X1 U23878 ( .B1(n20913), .B2(keyinput40), .C1(n20912), .C2(keyinput72), .A(n20911), .ZN(n20914) );
  NOR3_X1 U23879 ( .A1(n20916), .A2(n20915), .A3(n20914), .ZN(n20933) );
  AOI22_X1 U23880 ( .A1(n20919), .A2(keyinput92), .B1(n20918), .B2(keyinput62), 
        .ZN(n20917) );
  OAI221_X1 U23881 ( .B1(n20919), .B2(keyinput92), .C1(n20918), .C2(keyinput62), .A(n20917), .ZN(n20931) );
  AOI22_X1 U23882 ( .A1(n21080), .A2(keyinput21), .B1(keyinput116), .B2(n20921), .ZN(n20920) );
  OAI221_X1 U23883 ( .B1(n21080), .B2(keyinput21), .C1(n20921), .C2(
        keyinput116), .A(n20920), .ZN(n20930) );
  AOI22_X1 U23884 ( .A1(n20924), .A2(keyinput75), .B1(keyinput18), .B2(n20923), 
        .ZN(n20922) );
  OAI221_X1 U23885 ( .B1(n20924), .B2(keyinput75), .C1(n20923), .C2(keyinput18), .A(n20922), .ZN(n20929) );
  INV_X1 U23886 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20926) );
  AOI22_X1 U23887 ( .A1(n20927), .A2(keyinput3), .B1(n20926), .B2(keyinput17), 
        .ZN(n20925) );
  OAI221_X1 U23888 ( .B1(n20927), .B2(keyinput3), .C1(n20926), .C2(keyinput17), 
        .A(n20925), .ZN(n20928) );
  NOR4_X1 U23889 ( .A1(n20931), .A2(n20930), .A3(n20929), .A4(n20928), .ZN(
        n20932) );
  NAND4_X1 U23890 ( .A1(n20935), .A2(n20934), .A3(n20933), .A4(n20932), .ZN(
        n21066) );
  AOI22_X1 U23891 ( .A1(n20938), .A2(keyinput22), .B1(n20937), .B2(keyinput89), 
        .ZN(n20936) );
  OAI221_X1 U23892 ( .B1(n20938), .B2(keyinput22), .C1(n20937), .C2(keyinput89), .A(n20936), .ZN(n20951) );
  INV_X1 U23893 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n20940) );
  AOI22_X1 U23894 ( .A1(n20941), .A2(keyinput93), .B1(n20940), .B2(keyinput69), 
        .ZN(n20939) );
  OAI221_X1 U23895 ( .B1(n20941), .B2(keyinput93), .C1(n20940), .C2(keyinput69), .A(n20939), .ZN(n20950) );
  AOI22_X1 U23896 ( .A1(n20944), .A2(keyinput11), .B1(keyinput44), .B2(n20943), 
        .ZN(n20942) );
  OAI221_X1 U23897 ( .B1(n20944), .B2(keyinput11), .C1(n20943), .C2(keyinput44), .A(n20942), .ZN(n20949) );
  AOI22_X1 U23898 ( .A1(n20947), .A2(keyinput108), .B1(n20946), .B2(keyinput37), .ZN(n20945) );
  OAI221_X1 U23899 ( .B1(n20947), .B2(keyinput108), .C1(n20946), .C2(
        keyinput37), .A(n20945), .ZN(n20948) );
  NOR4_X1 U23900 ( .A1(n20951), .A2(n20950), .A3(n20949), .A4(n20948), .ZN(
        n20998) );
  AOI22_X1 U23901 ( .A1(n20954), .A2(keyinput110), .B1(keyinput111), .B2(
        n20953), .ZN(n20952) );
  OAI221_X1 U23902 ( .B1(n20954), .B2(keyinput110), .C1(n20953), .C2(
        keyinput111), .A(n20952), .ZN(n20966) );
  AOI22_X1 U23903 ( .A1(n20956), .A2(keyinput38), .B1(n10056), .B2(keyinput68), 
        .ZN(n20955) );
  OAI221_X1 U23904 ( .B1(n20956), .B2(keyinput38), .C1(n10056), .C2(keyinput68), .A(n20955), .ZN(n20965) );
  AOI22_X1 U23905 ( .A1(n20959), .A2(keyinput19), .B1(n20958), .B2(keyinput96), 
        .ZN(n20957) );
  OAI221_X1 U23906 ( .B1(n20959), .B2(keyinput19), .C1(n20958), .C2(keyinput96), .A(n20957), .ZN(n20964) );
  AOI22_X1 U23907 ( .A1(n20962), .A2(keyinput45), .B1(n20961), .B2(keyinput23), 
        .ZN(n20960) );
  OAI221_X1 U23908 ( .B1(n20962), .B2(keyinput45), .C1(n20961), .C2(keyinput23), .A(n20960), .ZN(n20963) );
  NOR4_X1 U23909 ( .A1(n20966), .A2(n20965), .A3(n20964), .A4(n20963), .ZN(
        n20997) );
  AOI22_X1 U23910 ( .A1(n20968), .A2(keyinput97), .B1(n14587), .B2(keyinput34), 
        .ZN(n20967) );
  OAI221_X1 U23911 ( .B1(n20968), .B2(keyinput97), .C1(n14587), .C2(keyinput34), .A(n20967), .ZN(n20980) );
  AOI22_X1 U23912 ( .A1(n11004), .A2(keyinput120), .B1(keyinput123), .B2(
        n20970), .ZN(n20969) );
  OAI221_X1 U23913 ( .B1(n11004), .B2(keyinput120), .C1(n20970), .C2(
        keyinput123), .A(n20969), .ZN(n20979) );
  AOI22_X1 U23914 ( .A1(n20973), .A2(keyinput2), .B1(n20972), .B2(keyinput32), 
        .ZN(n20971) );
  OAI221_X1 U23915 ( .B1(n20973), .B2(keyinput2), .C1(n20972), .C2(keyinput32), 
        .A(n20971), .ZN(n20978) );
  AOI22_X1 U23916 ( .A1(n20976), .A2(keyinput118), .B1(n20975), .B2(keyinput82), .ZN(n20974) );
  OAI221_X1 U23917 ( .B1(n20976), .B2(keyinput118), .C1(n20975), .C2(
        keyinput82), .A(n20974), .ZN(n20977) );
  NOR4_X1 U23918 ( .A1(n20980), .A2(n20979), .A3(n20978), .A4(n20977), .ZN(
        n20996) );
  AOI22_X1 U23919 ( .A1(n20983), .A2(keyinput90), .B1(n20982), .B2(keyinput9), 
        .ZN(n20981) );
  OAI221_X1 U23920 ( .B1(n20983), .B2(keyinput90), .C1(n20982), .C2(keyinput9), 
        .A(n20981), .ZN(n20994) );
  AOI22_X1 U23921 ( .A1(n20985), .A2(keyinput70), .B1(n14168), .B2(keyinput87), 
        .ZN(n20984) );
  OAI221_X1 U23922 ( .B1(n20985), .B2(keyinput70), .C1(n14168), .C2(keyinput87), .A(n20984), .ZN(n20993) );
  AOI22_X1 U23923 ( .A1(n20988), .A2(keyinput125), .B1(n20987), .B2(keyinput95), .ZN(n20986) );
  OAI221_X1 U23924 ( .B1(n20988), .B2(keyinput125), .C1(n20987), .C2(
        keyinput95), .A(n20986), .ZN(n20992) );
  AOI22_X1 U23925 ( .A1(n20990), .A2(keyinput122), .B1(n13461), .B2(
        keyinput103), .ZN(n20989) );
  NOR4_X1 U23926 ( .A1(n20994), .A2(n20993), .A3(n20992), .A4(n20991), .ZN(
        n20995) );
  NAND4_X1 U23927 ( .A1(n20998), .A2(n20997), .A3(n20996), .A4(n20995), .ZN(
        n21065) );
  AOI22_X1 U23928 ( .A1(n21001), .A2(keyinput80), .B1(n21000), .B2(keyinput35), 
        .ZN(n20999) );
  OAI221_X1 U23929 ( .B1(n21001), .B2(keyinput80), .C1(n21000), .C2(keyinput35), .A(n20999), .ZN(n21013) );
  AOI22_X1 U23930 ( .A1(n21004), .A2(keyinput0), .B1(n21003), .B2(keyinput114), 
        .ZN(n21002) );
  OAI221_X1 U23931 ( .B1(n21004), .B2(keyinput0), .C1(n21003), .C2(keyinput114), .A(n21002), .ZN(n21012) );
  AOI22_X1 U23932 ( .A1(n21007), .A2(keyinput25), .B1(keyinput102), .B2(n21006), .ZN(n21005) );
  OAI221_X1 U23933 ( .B1(n21007), .B2(keyinput25), .C1(n21006), .C2(
        keyinput102), .A(n21005), .ZN(n21011) );
  XNOR2_X1 U23934 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B(keyinput64), .ZN(
        n21009) );
  XNOR2_X1 U23935 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B(keyinput88), .ZN(
        n21008) );
  NAND2_X1 U23936 ( .A1(n21009), .A2(n21008), .ZN(n21010) );
  NOR4_X1 U23937 ( .A1(n21013), .A2(n21012), .A3(n21011), .A4(n21010), .ZN(
        n21063) );
  INV_X1 U23938 ( .A(P3_UWORD_REG_12__SCAN_IN), .ZN(n21015) );
  AOI22_X1 U23939 ( .A1(n21016), .A2(keyinput73), .B1(keyinput112), .B2(n21015), .ZN(n21014) );
  OAI221_X1 U23940 ( .B1(n21016), .B2(keyinput73), .C1(n21015), .C2(
        keyinput112), .A(n21014), .ZN(n21029) );
  AOI22_X1 U23941 ( .A1(n21019), .A2(keyinput16), .B1(n21018), .B2(keyinput121), .ZN(n21017) );
  OAI221_X1 U23942 ( .B1(n21019), .B2(keyinput16), .C1(n21018), .C2(
        keyinput121), .A(n21017), .ZN(n21028) );
  AOI22_X1 U23943 ( .A1(n21022), .A2(keyinput109), .B1(n21021), .B2(keyinput28), .ZN(n21020) );
  OAI221_X1 U23944 ( .B1(n21022), .B2(keyinput109), .C1(n21021), .C2(
        keyinput28), .A(n21020), .ZN(n21027) );
  AOI22_X1 U23945 ( .A1(n21025), .A2(keyinput59), .B1(keyinput36), .B2(n21024), 
        .ZN(n21023) );
  OAI221_X1 U23946 ( .B1(n21025), .B2(keyinput59), .C1(n21024), .C2(keyinput36), .A(n21023), .ZN(n21026) );
  NOR4_X1 U23947 ( .A1(n21029), .A2(n21028), .A3(n21027), .A4(n21026), .ZN(
        n21062) );
  AOI22_X1 U23948 ( .A1(n21032), .A2(keyinput50), .B1(keyinput58), .B2(n21031), 
        .ZN(n21030) );
  OAI221_X1 U23949 ( .B1(n21032), .B2(keyinput50), .C1(n21031), .C2(keyinput58), .A(n21030), .ZN(n21045) );
  AOI22_X1 U23950 ( .A1(n21035), .A2(keyinput55), .B1(n21034), .B2(keyinput5), 
        .ZN(n21033) );
  OAI221_X1 U23951 ( .B1(n21035), .B2(keyinput55), .C1(n21034), .C2(keyinput5), 
        .A(n21033), .ZN(n21044) );
  INV_X1 U23952 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n21037) );
  AOI22_X1 U23953 ( .A1(n21038), .A2(keyinput20), .B1(n21037), .B2(keyinput99), 
        .ZN(n21036) );
  OAI221_X1 U23954 ( .B1(n21038), .B2(keyinput20), .C1(n21037), .C2(keyinput99), .A(n21036), .ZN(n21043) );
  AOI22_X1 U23955 ( .A1(n21041), .A2(keyinput107), .B1(keyinput106), .B2(
        n21040), .ZN(n21039) );
  OAI221_X1 U23956 ( .B1(n21041), .B2(keyinput107), .C1(n21040), .C2(
        keyinput106), .A(n21039), .ZN(n21042) );
  NOR4_X1 U23957 ( .A1(n21045), .A2(n21044), .A3(n21043), .A4(n21042), .ZN(
        n21061) );
  AOI22_X1 U23958 ( .A1(n21048), .A2(keyinput14), .B1(keyinput126), .B2(n21047), .ZN(n21046) );
  OAI221_X1 U23959 ( .B1(n21048), .B2(keyinput14), .C1(n21047), .C2(
        keyinput126), .A(n21046), .ZN(n21059) );
  AOI22_X1 U23960 ( .A1(n21051), .A2(keyinput61), .B1(keyinput74), .B2(n21050), 
        .ZN(n21049) );
  OAI221_X1 U23961 ( .B1(n21051), .B2(keyinput61), .C1(n21050), .C2(keyinput74), .A(n21049), .ZN(n21058) );
  AOI22_X1 U23962 ( .A1(n21053), .A2(keyinput84), .B1(n18981), .B2(keyinput33), 
        .ZN(n21052) );
  OAI221_X1 U23963 ( .B1(n21053), .B2(keyinput84), .C1(n18981), .C2(keyinput33), .A(n21052), .ZN(n21057) );
  INV_X1 U23964 ( .A(DATAI_31_), .ZN(n21106) );
  AOI22_X1 U23965 ( .A1(n21055), .A2(keyinput53), .B1(keyinput15), .B2(n21106), 
        .ZN(n21054) );
  OAI221_X1 U23966 ( .B1(n21055), .B2(keyinput53), .C1(n21106), .C2(keyinput15), .A(n21054), .ZN(n21056) );
  NOR4_X1 U23967 ( .A1(n21059), .A2(n21058), .A3(n21057), .A4(n21056), .ZN(
        n21060) );
  NAND4_X1 U23968 ( .A1(n21063), .A2(n21062), .A3(n21061), .A4(n21060), .ZN(
        n21064) );
  NOR4_X1 U23969 ( .A1(n21067), .A2(n21066), .A3(n21065), .A4(n21064), .ZN(
        n21131) );
  OAI22_X1 U23970 ( .A1(n21071), .A2(n21070), .B1(n21069), .B2(n21068), .ZN(
        n21077) );
  OAI22_X1 U23971 ( .A1(n21075), .A2(n21074), .B1(n21073), .B2(n21072), .ZN(
        n21076) );
  AOI211_X1 U23972 ( .C1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .C2(n21078), .A(
        n21077), .B(n21076), .ZN(n21129) );
  NOR4_X1 U23973 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        n21079), .ZN(n21090) );
  NOR4_X1 U23974 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_11__2__SCAN_IN), .A3(P1_INSTQUEUE_REG_7__3__SCAN_IN), 
        .A4(n21080), .ZN(n21081) );
  NAND3_X1 U23975 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_14__4__SCAN_IN), .A3(n21081), .ZN(n21087) );
  NOR4_X1 U23976 ( .A1(P3_DATAO_REG_12__SCAN_IN), .A2(P3_DATAO_REG_20__SCAN_IN), .A3(P3_MEMORYFETCH_REG_SCAN_IN), .A4(P3_M_IO_N_REG_SCAN_IN), .ZN(n21085) );
  NOR4_X1 U23977 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(
        P1_BYTEENABLE_REG_2__SCAN_IN), .A3(P3_ADDRESS_REG_9__SCAN_IN), .A4(
        P3_DATAO_REG_11__SCAN_IN), .ZN(n21084) );
  NOR4_X1 U23978 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), .A3(P1_ADS_N_REG_SCAN_IN), .A4(P1_UWORD_REG_8__SCAN_IN), .ZN(n21083) );
  NOR4_X1 U23979 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_DATAO_REG_15__SCAN_IN), 
        .A3(P2_DATAO_REG_16__SCAN_IN), .A4(P2_DATAO_REG_25__SCAN_IN), .ZN(
        n21082) );
  NAND4_X1 U23980 ( .A1(n21085), .A2(n21084), .A3(n21083), .A4(n21082), .ZN(
        n21086) );
  NOR4_X1 U23981 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21088), .A3(
        n21087), .A4(n21086), .ZN(n21089) );
  NAND4_X1 U23982 ( .A1(n21092), .A2(n21091), .A3(n21090), .A4(n21089), .ZN(
        n21127) );
  NOR4_X1 U23983 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_12__1__SCAN_IN), .A3(P2_INSTQUEUE_REG_7__1__SCAN_IN), 
        .A4(BUF1_REG_29__SCAN_IN), .ZN(n21096) );
  NOR4_X1 U23984 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(P3_EBX_REG_8__SCAN_IN), .ZN(
        n21095) );
  NOR4_X1 U23985 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_EAX_REG_29__SCAN_IN), .A3(P1_REIP_REG_10__SCAN_IN), .A4(
        P1_REIP_REG_11__SCAN_IN), .ZN(n21094) );
  NOR4_X1 U23986 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A3(P1_EAX_REG_11__SCAN_IN), .A4(
        P1_REIP_REG_9__SCAN_IN), .ZN(n21093) );
  NAND4_X1 U23987 ( .A1(n21096), .A2(n21095), .A3(n21094), .A4(n21093), .ZN(
        n21126) );
  NOR4_X1 U23988 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .A3(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_16__SCAN_IN), .ZN(n21100) );
  NOR4_X1 U23989 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(
        P2_STATE_REG_2__SCAN_IN), .A3(P2_EAX_REG_3__SCAN_IN), .A4(
        BUF1_REG_3__SCAN_IN), .ZN(n21099) );
  NOR4_X1 U23990 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_8__5__SCAN_IN), .A3(P3_INSTQUEUE_REG_5__4__SCAN_IN), 
        .A4(P3_REIP_REG_8__SCAN_IN), .ZN(n21098) );
  NOR4_X1 U23991 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A4(BUF2_REG_5__SCAN_IN), .ZN(
        n21097) );
  NAND4_X1 U23992 ( .A1(n21100), .A2(n21099), .A3(n21098), .A4(n21097), .ZN(
        n21125) );
  NAND4_X1 U23993 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P1_EAX_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .A4(
        P2_LWORD_REG_10__SCAN_IN), .ZN(n21104) );
  NAND4_X1 U23994 ( .A1(P3_DATAO_REG_27__SCAN_IN), .A2(
        P1_UWORD_REG_10__SCAN_IN), .A3(P1_LWORD_REG_3__SCAN_IN), .A4(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n21103) );
  NAND4_X1 U23995 ( .A1(P2_EBX_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), 
        .A4(P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21102) );
  NAND4_X1 U23996 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(P2_UWORD_REG_6__SCAN_IN), 
        .A3(P2_LWORD_REG_6__SCAN_IN), .A4(P2_UWORD_REG_14__SCAN_IN), .ZN(
        n21101) );
  NOR4_X1 U23997 ( .A1(n21104), .A2(n21103), .A3(n21102), .A4(n21101), .ZN(
        n21123) );
  NAND4_X1 U23998 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), .A3(P2_DATAO_REG_13__SCAN_IN), .A4(P3_LWORD_REG_1__SCAN_IN), .ZN(n21111) );
  NAND4_X1 U23999 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n21107), .A3(n21106), 
        .A4(n21105), .ZN(n21110) );
  NAND4_X1 U24000 ( .A1(P3_ADDRESS_REG_6__SCAN_IN), .A2(
        P3_UWORD_REG_1__SCAN_IN), .A3(P2_DATAO_REG_0__SCAN_IN), .A4(
        P3_DATAO_REG_25__SCAN_IN), .ZN(n21109) );
  NAND4_X1 U24001 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(
        P3_ADDRESS_REG_14__SCAN_IN), .A3(P3_DATAO_REG_17__SCAN_IN), .A4(
        P3_ADDRESS_REG_7__SCAN_IN), .ZN(n21108) );
  NOR4_X1 U24002 ( .A1(n21111), .A2(n21110), .A3(n21109), .A4(n21108), .ZN(
        n21122) );
  NAND4_X1 U24003 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_13__2__SCAN_IN), .A3(P2_EAX_REG_20__SCAN_IN), .A4(
        BUF1_REG_19__SCAN_IN), .ZN(n21115) );
  NAND4_X1 U24004 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(P3_REIP_REG_31__SCAN_IN), 
        .A3(P3_EBX_REG_15__SCAN_IN), .A4(P3_EBX_REG_4__SCAN_IN), .ZN(n21114)
         );
  NAND4_X1 U24005 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(P1_EAX_REG_17__SCAN_IN), .A4(
        BUF1_REG_24__SCAN_IN), .ZN(n21113) );
  NAND4_X1 U24006 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .A3(P2_INSTQUEUE_REG_10__2__SCAN_IN), 
        .A4(BUF1_REG_25__SCAN_IN), .ZN(n21112) );
  NOR4_X1 U24007 ( .A1(n21115), .A2(n21114), .A3(n21113), .A4(n21112), .ZN(
        n21121) );
  NAND4_X1 U24008 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A4(P3_UWORD_REG_12__SCAN_IN), 
        .ZN(n21119) );
  NAND4_X1 U24009 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_0__4__SCAN_IN), .A3(P3_STATE_REG_2__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n21118) );
  NAND4_X1 U24010 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .A3(P3_INSTQUEUE_REG_14__5__SCAN_IN), 
        .A4(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n21117) );
  NAND4_X1 U24011 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .A3(P3_INSTQUEUE_REG_8__0__SCAN_IN), 
        .A4(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n21116) );
  NOR4_X1 U24012 ( .A1(n21119), .A2(n21118), .A3(n21117), .A4(n21116), .ZN(
        n21120) );
  NAND4_X1 U24013 ( .A1(n21123), .A2(n21122), .A3(n21121), .A4(n21120), .ZN(
        n21124) );
  NOR4_X1 U24014 ( .A1(n21127), .A2(n21126), .A3(n21125), .A4(n21124), .ZN(
        n21128) );
  XOR2_X1 U24015 ( .A(n21129), .B(n21128), .Z(n21130) );
  XNOR2_X1 U24016 ( .A(n21131), .B(n21130), .ZN(P1_U3135) );
  AND2_X2 U11188 ( .A1(n14669), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9900) );
  AOI21_X2 U11442 ( .B1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n12243), .A(
        n10017), .ZN(n10016) );
  NOR2_X4 U11847 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11723) );
  OAI21_X1 U11378 ( .B1(n12729), .B2(n12740), .A(n12728), .ZN(n13104) );
  NAND2_X1 U11238 ( .A1(n10108), .A2(n15794), .ZN(n14685) );
  NAND2_X2 U11242 ( .A1(n10120), .A2(n10119), .ZN(n14744) );
  AND2_X2 U11422 ( .A1(n11845), .A2(n20176), .ZN(n12733) );
  AND2_X2 U12786 ( .A1(n11728), .A2(n11732), .ZN(n11916) );
  AND4_X1 U11189 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11760) );
  AND4_X1 U11460 ( .A1(n11755), .A2(n11754), .A3(n11753), .A4(n11752), .ZN(
        n11761) );
  AND4_X2 U14925 ( .A1(n11763), .A2(n11762), .A3(n11761), .A4(n11760), .ZN(
        n20171) );
  INV_X2 U11284 ( .A(n10309), .ZN(n10267) );
  INV_X2 U11166 ( .A(n10267), .ZN(n17177) );
  INV_X1 U11665 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12543) );
  NAND2_X1 U11515 ( .A1(n12240), .A2(n12239), .ZN(n14451) );
  CLKBUF_X1 U11174 ( .A(n11965), .Z(n11902) );
  OR2_X1 U11214 ( .A1(n11909), .A2(n11908), .ZN(n12780) );
  AND2_X1 U11220 ( .A1(n13137), .A2(n12591), .ZN(n9886) );
  AND2_X2 U11232 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13346) );
  NOR2_X1 U11233 ( .A1(n12009), .A2(n12790), .ZN(n12787) );
  AND2_X1 U11234 ( .A1(n13346), .A2(n11728), .ZN(n11917) );
  AND4_X1 U11281 ( .A1(n11727), .A2(n11726), .A3(n11725), .A4(n11724), .ZN(
        n9803) );
  CLKBUF_X1 U11302 ( .A(n10728), .Z(n10740) );
  NAND2_X1 U11439 ( .A1(n14652), .A2(n14662), .ZN(n12809) );
  AND4_X1 U11498 ( .A1(n9822), .A2(n11775), .A3(n9774), .A4(n11774), .ZN(
        n12813) );
  BUF_X1 U11500 ( .A(n17031), .Z(n17038) );
  AND4_X2 U11505 ( .A1(n11813), .A2(n11812), .A3(n11811), .A4(n11810), .ZN(
        n20144) );
  INV_X1 U11506 ( .A(n13882), .ZN(n12240) );
  NAND2_X1 U11516 ( .A1(n12811), .A2(n12810), .ZN(n9885) );
  NAND2_X1 U11543 ( .A1(n12807), .A2(n15794), .ZN(n14662) );
  NAND2_X1 U11589 ( .A1(n14705), .A2(n10112), .ZN(n9892) );
  NAND2_X1 U11606 ( .A1(n13409), .A2(n12748), .ZN(n20079) );
  NAND2_X2 U11736 ( .A1(n9988), .A2(n9986), .ZN(n13814) );
  CLKBUF_X2 U12424 ( .A(n10371), .Z(n9719) );
  NAND2_X1 U12493 ( .A1(n9893), .A2(n9892), .ZN(n14692) );
  CLKBUF_X1 U12645 ( .A(n16473), .Z(n16481) );
endmodule

