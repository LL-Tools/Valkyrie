

module b22_C_SARLock_k_128_8 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6580, n6581, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620;

  INV_X4 U7329 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U7330 ( .A1(n13769), .A2(n7640), .ZN(n13849) );
  NAND2_X1 U7331 ( .A1(n9238), .A2(n9237), .ZN(n14266) );
  NAND2_X1 U7332 ( .A1(n8882), .A2(n8881), .ZN(n14270) );
  INV_X1 U7333 ( .A(n13151), .ZN(n13186) );
  NAND2_X1 U7334 ( .A1(n12018), .A2(n7404), .ZN(n10386) );
  BUF_X1 U7335 ( .A(n10158), .Z(n12592) );
  NAND2_X2 U7336 ( .A1(n9425), .A2(n7274), .ZN(n8478) );
  AND2_X1 U7337 ( .A1(n10014), .A2(n10013), .ZN(n12325) );
  INV_X1 U7338 ( .A(n9751), .ZN(n11844) );
  INV_X2 U7339 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7976) );
  CLKBUF_X1 U7340 ( .A(n15114), .Z(n6580) );
  OAI21_X1 U7341 ( .B1(n9019), .B2(n11795), .A(n9272), .ZN(n15114) );
  CLKBUF_X1 U7342 ( .A(n15327), .Z(n6581) );
  NOR2_X1 U7343 ( .A1(n15331), .A2(n9297), .ZN(n15327) );
  NOR4_X1 U7344 ( .A1(n12222), .A2(n7637), .A3(n12221), .A4(n12220), .ZN(
        n12225) );
  INV_X1 U7345 ( .A(n12417), .ZN(n12467) );
  NAND2_X1 U7346 ( .A1(n9020), .A2(n9019), .ZN(n9265) );
  NOR4_X1 U7347 ( .A1(n12520), .A2(n12519), .A3(n14600), .A4(n12518), .ZN(
        n12521) );
  AND2_X1 U7348 ( .A1(n13695), .A2(n12887), .ZN(n7637) );
  INV_X1 U7349 ( .A(n12183), .ZN(n12165) );
  CLKBUF_X2 U7350 ( .A(n12734), .Z(n6801) );
  OAI21_X1 U7351 ( .B1(n15448), .B2(n8267), .A(n8266), .ZN(n11401) );
  INV_X1 U7352 ( .A(n12592), .ZN(n13792) );
  INV_X1 U7353 ( .A(n12666), .ZN(n12708) );
  NAND2_X1 U7354 ( .A1(n14632), .A2(n14631), .ZN(n14630) );
  INV_X1 U7355 ( .A(n11695), .ZN(n14768) );
  NOR2_X1 U7356 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n7267) );
  INV_X1 U7357 ( .A(n12833), .ZN(n13601) );
  AND2_X1 U7358 ( .A1(n13621), .A2(n15569), .ZN(n6766) );
  INV_X1 U7359 ( .A(n8520), .ZN(n8983) );
  XNOR2_X1 U7360 ( .A(n14087), .B(n13896), .ZN(n14082) );
  INV_X2 U7361 ( .A(n11728), .ZN(n12710) );
  INV_X1 U7362 ( .A(n12289), .ZN(n11985) );
  NAND3_X1 U7363 ( .A1(n9330), .A2(n7268), .A3(n7267), .ZN(n9520) );
  INV_X1 U7364 ( .A(n7798), .ZN(n10629) );
  INV_X1 U7365 ( .A(n7819), .ZN(n12039) );
  INV_X1 U7366 ( .A(n10221), .ZN(n13038) );
  NOR2_X1 U7367 ( .A1(n13962), .A2(n13997), .ZN(n14174) );
  XNOR2_X1 U7368 ( .A(n8466), .B(n8465), .ZN(n9439) );
  AND2_X1 U7369 ( .A1(n9404), .A2(n9400), .ZN(n9323) );
  OR2_X1 U7370 ( .A1(n14338), .A2(n14337), .ZN(n14339) );
  NAND2_X1 U7371 ( .A1(n14339), .A2(n6808), .ZN(n14397) );
  AND2_X1 U7372 ( .A1(n6590), .A2(n12298), .ZN(n15233) );
  NAND2_X1 U7373 ( .A1(n15054), .A2(n6832), .ZN(n15175) );
  INV_X1 U7374 ( .A(n8938), .ZN(n9019) );
  OR2_X1 U7375 ( .A1(n6594), .A2(n14177), .ZN(P2_U3529) );
  BUF_X1 U7376 ( .A(n8937), .Z(n6585) );
  INV_X2 U7377 ( .A(n9914), .ZN(n10037) );
  INV_X2 U7378 ( .A(n9265), .ZN(n7523) );
  NAND2_X2 U7379 ( .A1(n8937), .A2(n11104), .ZN(n9898) );
  NOR2_X2 U7380 ( .A1(n11157), .A2(n15249), .ZN(n11158) );
  NAND2_X2 U7381 ( .A1(n12618), .A2(n12617), .ZN(n12622) );
  OR2_X2 U7382 ( .A1(n11739), .A2(n11740), .ZN(n12618) );
  NAND2_X1 U7383 ( .A1(n6602), .A2(n9750), .ZN(n7819) );
  NAND2_X2 U7384 ( .A1(n12763), .A2(n12762), .ZN(n12761) );
  AND2_X2 U7385 ( .A1(n6597), .A2(n6598), .ZN(n12763) );
  NAND2_X4 U7386 ( .A1(n7638), .A2(n7142), .ZN(n14166) );
  OAI21_X2 U7387 ( .B1(n13803), .B2(n13872), .A(n13791), .ZN(n13795) );
  NOR2_X2 U7388 ( .A1(n10435), .A2(n10434), .ZN(n11085) );
  NAND2_X2 U7389 ( .A1(n8980), .A2(n9439), .ZN(n9425) );
  INV_X4 U7390 ( .A(n8162), .ZN(n8134) );
  INV_X2 U7391 ( .A(n7834), .ZN(n8162) );
  OAI21_X1 U7392 ( .B1(n9527), .B2(n9526), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9530) );
  INV_X1 U7393 ( .A(n7868), .ZN(n6583) );
  CLKBUF_X1 U7394 ( .A(n15027), .Z(n6584) );
  XNOR2_X1 U7395 ( .A(n9530), .B(n9529), .ZN(n15027) );
  NOR2_X2 U7396 ( .A1(n10338), .A2(n12312), .ZN(n10849) );
  INV_X1 U7397 ( .A(n12312), .ZN(n12314) );
  NAND2_X2 U7398 ( .A1(n9795), .A2(n9794), .ZN(n12312) );
  AND2_X2 U7399 ( .A1(n8207), .A2(n8206), .ZN(n13703) );
  AND2_X2 U7400 ( .A1(n10256), .A2(n9310), .ZN(n9315) );
  BUF_X4 U7401 ( .A(n8484), .Z(n8738) );
  AOI21_X2 U7402 ( .B1(n6973), .B2(n6972), .A(n6687), .ZN(n6971) );
  NAND4_X2 U7403 ( .A1(n7789), .A2(n7788), .A3(n7787), .A4(n7786), .ZN(n7798)
         );
  OR2_X2 U7404 ( .A1(n11986), .A2(n9843), .ZN(n7410) );
  NAND2_X2 U7405 ( .A1(n11595), .A2(n6701), .ZN(n12240) );
  NAND2_X2 U7406 ( .A1(n6757), .A2(n6756), .ZN(n11595) );
  INV_X2 U7407 ( .A(n15023), .ZN(n9747) );
  NAND2_X2 U7408 ( .A1(n8472), .A2(n7634), .ZN(n9901) );
  NOR2_X2 U7409 ( .A1(n7513), .A2(n6638), .ZN(n12011) );
  NAND2_X2 U7410 ( .A1(n11817), .A2(n11816), .ZN(n14830) );
  OAI22_X1 U7411 ( .A1(n9800), .A2(n12315), .B1(n12314), .B2(n12665), .ZN(
        n10000) );
  XNOR2_X2 U7412 ( .A(n8880), .B(n8879), .ZN(n14307) );
  NOR2_X2 U7413 ( .A1(n14329), .A2(n7346), .ZN(n7345) );
  OAI22_X2 U7414 ( .A1(n10569), .A2(n7289), .B1(n12345), .B2(n10513), .ZN(
        n10723) );
  OAI21_X2 U7415 ( .B1(n7737), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n15180), .ZN(
        n15185) );
  XNOR2_X2 U7416 ( .A(n11192), .B(n11049), .ZN(n11052) );
  XNOR2_X2 U7417 ( .A(n7773), .B(n7772), .ZN(n10196) );
  NAND2_X2 U7418 ( .A1(n11048), .A2(n11047), .ZN(n11192) );
  INV_X1 U7419 ( .A(n15034), .ZN(n6590) );
  NOR2_X2 U7420 ( .A1(n9746), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n7323) );
  AND2_X2 U7421 ( .A1(n8174), .A2(n8173), .ZN(n13711) );
  AND2_X2 U7422 ( .A1(n14082), .A2(n7485), .ZN(n7484) );
  NAND2_X2 U7423 ( .A1(n8844), .A2(n8843), .ZN(n14031) );
  INV_X1 U7424 ( .A(n9748), .ZN(n15020) );
  AND4_X2 U7425 ( .A1(n7749), .A2(n7748), .A3(n7839), .A4(n7747), .ZN(n7750)
         );
  NOR2_X2 U7426 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n7748) );
  XNOR2_X2 U7427 ( .A(n9317), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9404) );
  XOR2_X2 U7428 ( .A(n14600), .B(n14597), .Z(n14876) );
  XNOR2_X1 U7429 ( .A(n12243), .B(n12241), .ZN(n12845) );
  NAND2_X1 U7430 ( .A1(n12240), .A2(n12239), .ZN(n12243) );
  OAI21_X2 U7431 ( .B1(n8244), .B2(P3_IR_REG_19__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8245) );
  OAI21_X2 U7432 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n7714), .A(n15040), .ZN(
        n15615) );
  OAI21_X2 U7433 ( .B1(n13204), .B2(n6999), .A(n7462), .ZN(n13181) );
  NAND2_X2 U7434 ( .A1(n8767), .A2(n8766), .ZN(n14233) );
  OAI22_X2 U7435 ( .A1(n13876), .A2(n13874), .B1(n12551), .B2(n12550), .ZN(
        n13830) );
  XNOR2_X2 U7436 ( .A(n12550), .B(n12551), .ZN(n13876) );
  NAND4_X4 U7437 ( .A1(n7803), .A2(n7802), .A3(n7801), .A4(n7800), .ZN(n12896)
         );
  NAND2_X2 U7438 ( .A1(n13224), .A2(n12147), .ZN(n13204) );
  OAI22_X2 U7439 ( .A1(n12770), .A2(n12769), .B1(n12768), .B2(n12888), .ZN(
        n12773) );
  NAND2_X2 U7440 ( .A1(n13747), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7761) );
  CLKBUF_X1 U7441 ( .A(n13038), .Z(n6586) );
  BUF_X8 U7442 ( .A(n13038), .Z(n6587) );
  NOR2_X2 U7443 ( .A1(n15415), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n7709) );
  AOI21_X1 U7444 ( .B1(n11994), .B2(n14939), .A(n11993), .ZN(n14624) );
  AND2_X1 U7445 ( .A1(n13849), .A2(n13850), .ZN(n13815) );
  NAND2_X1 U7446 ( .A1(n14368), .A2(n14369), .ZN(n14367) );
  CLKBUF_X1 U7447 ( .A(n11969), .Z(n6799) );
  NAND2_X2 U7448 ( .A1(n11811), .A2(n11810), .ZN(n14980) );
  AND2_X1 U7449 ( .A1(n7046), .A2(n6736), .ZN(n13032) );
  NAND2_X1 U7450 ( .A1(n7263), .A2(n6643), .ZN(n7048) );
  NAND2_X1 U7451 ( .A1(n14816), .A2(n11818), .ZN(n14800) );
  NAND2_X1 U7452 ( .A1(n7968), .A2(n6619), .ZN(n13685) );
  NAND2_X1 U7453 ( .A1(n11447), .A2(n7095), .ZN(n11640) );
  NAND2_X1 U7454 ( .A1(n7733), .A2(n15051), .ZN(n15056) );
  NAND2_X1 U7455 ( .A1(n15053), .A2(n15052), .ZN(n15051) );
  XNOR2_X1 U7456 ( .A(n7732), .B(n7118), .ZN(n15053) );
  INV_X1 U7457 ( .A(n14429), .ZN(n12341) );
  INV_X1 U7458 ( .A(n12895), .ZN(n11173) );
  INV_X1 U7459 ( .A(n15459), .ZN(n11035) );
  NAND2_X2 U7460 ( .A1(n10629), .A2(n10533), .ZN(n12055) );
  AND2_X1 U7461 ( .A1(n10849), .A2(n15236), .ZN(n10850) );
  AND2_X1 U7462 ( .A1(n12489), .A2(n15232), .ZN(n12487) );
  INV_X4 U7463 ( .A(n7523), .ZN(n9173) );
  CLKBUF_X3 U7464 ( .A(n9799), .Z(n12666) );
  INV_X4 U7465 ( .A(n10037), .ZN(n13997) );
  AND4_X1 U7466 ( .A1(n10018), .A2(n10017), .A3(n10016), .A4(n10015), .ZN(
        n12326) );
  CLKBUF_X2 U7467 ( .A(P2_U3947), .Z(n6589) );
  INV_X1 U7468 ( .A(n12450), .ZN(n11944) );
  INV_X1 U7469 ( .A(n13915), .ZN(n10135) );
  AND3_X1 U7470 ( .A1(n7785), .A2(n7784), .A3(n7783), .ZN(n10524) );
  INV_X2 U7471 ( .A(n12339), .ZN(n6588) );
  NAND2_X1 U7472 ( .A1(n15020), .A2(n9747), .ZN(n11649) );
  AND2_X2 U7474 ( .A1(n7764), .A2(n7765), .ZN(n7831) );
  NAND2_X1 U7475 ( .A1(n8473), .A2(n8477), .ZN(n9752) );
  CLKBUF_X1 U7476 ( .A(n9559), .Z(n14490) );
  XNOR2_X1 U7477 ( .A(n9716), .B(n9715), .ZN(n11165) );
  CLKBUF_X1 U7478 ( .A(n10298), .Z(n6753) );
  NAND2_X1 U7480 ( .A1(n7274), .A2(P3_U3151), .ZN(n12609) );
  INV_X1 U7481 ( .A(n6966), .ZN(n8710) );
  AND2_X1 U7482 ( .A1(n8545), .A2(n8362), .ZN(n8365) );
  NOR2_X1 U7483 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n8364) );
  NOR2_X1 U7484 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n8363) );
  NOR2_X4 U7485 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7160) );
  NAND2_X1 U7486 ( .A1(n6825), .A2(n6824), .ZN(n13620) );
  OAI211_X1 U7487 ( .C1(n14615), .C2(n15229), .A(n14624), .B(n14620), .ZN(
        n14979) );
  OR2_X1 U7488 ( .A1(n9275), .A2(n9270), .ZN(n6900) );
  NAND2_X1 U7489 ( .A1(n12686), .A2(n12685), .ZN(n14358) );
  NAND2_X1 U7490 ( .A1(n13764), .A2(n13763), .ZN(n13803) );
  NAND2_X1 U7491 ( .A1(n14347), .A2(n12663), .ZN(n14406) );
  NAND2_X1 U7492 ( .A1(n6930), .A2(n7373), .ZN(n13764) );
  INV_X1 U7493 ( .A(n13108), .ZN(n13102) );
  NAND2_X1 U7494 ( .A1(n6744), .A2(n6855), .ZN(n14188) );
  AND2_X1 U7495 ( .A1(n13096), .A2(n10799), .ZN(n7083) );
  NAND2_X1 U7496 ( .A1(n8222), .A2(n8221), .ZN(n13096) );
  NOR2_X1 U7497 ( .A1(n14591), .A2(n14602), .ZN(n14584) );
  OR2_X1 U7498 ( .A1(n14042), .A2(n9291), .ZN(n14043) );
  OR2_X1 U7499 ( .A1(n14266), .A2(n14173), .ZN(n6596) );
  NAND2_X1 U7500 ( .A1(n14367), .A2(n12632), .ZN(n14377) );
  NOR2_X1 U7501 ( .A1(n13021), .A2(n13022), .ZN(n13033) );
  AND2_X1 U7502 ( .A1(n14980), .A2(n14634), .ZN(n7312) );
  NAND2_X2 U7503 ( .A1(n12804), .A2(n13122), .ZN(n12169) );
  NAND2_X1 U7504 ( .A1(n6933), .A2(n6765), .ZN(n13807) );
  OR2_X1 U7505 ( .A1(n8203), .A2(n8202), .ZN(n8204) );
  NAND2_X1 U7506 ( .A1(n7048), .A2(n7047), .ZN(n7046) );
  NAND2_X1 U7507 ( .A1(n8870), .A2(n8869), .ZN(n14189) );
  NAND2_X1 U7508 ( .A1(n11943), .A2(n11942), .ZN(n14878) );
  AND2_X1 U7509 ( .A1(n6932), .A2(n13808), .ZN(n6765) );
  NAND2_X1 U7510 ( .A1(n7158), .A2(n7157), .ZN(n14689) );
  NAND2_X1 U7511 ( .A1(n14800), .A2(n11827), .ZN(n11829) );
  OR2_X1 U7512 ( .A1(n12949), .A2(n7196), .ZN(n7195) );
  NAND2_X1 U7513 ( .A1(n14052), .A2(n8993), .ZN(n14053) );
  NAND2_X1 U7514 ( .A1(n8856), .A2(n8855), .ZN(n14196) );
  NAND2_X1 U7515 ( .A1(n11931), .A2(n11930), .ZN(n14887) );
  NAND2_X1 U7516 ( .A1(n11965), .A2(n12388), .ZN(n14820) );
  AND2_X1 U7517 ( .A1(n12960), .A2(n12959), .ZN(n12984) );
  NAND2_X1 U7518 ( .A1(n14817), .A2(n14821), .ZN(n14816) );
  NAND2_X1 U7519 ( .A1(n11917), .A2(n11916), .ZN(n14987) );
  NAND2_X1 U7520 ( .A1(n7099), .A2(n11813), .ZN(n14817) );
  OAI21_X1 U7521 ( .B1(n8854), .B2(n13511), .A(n8852), .ZN(n8457) );
  NAND2_X1 U7522 ( .A1(n6877), .A2(n7633), .ZN(n6878) );
  NOR2_X2 U7523 ( .A1(n14085), .A2(n14210), .ZN(n14052) );
  NAND2_X1 U7524 ( .A1(n8167), .A2(n8153), .ZN(n8168) );
  AND2_X1 U7525 ( .A1(n12922), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6877) );
  OR2_X1 U7526 ( .A1(n8152), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8167) );
  NAND2_X1 U7527 ( .A1(n6843), .A2(n6842), .ZN(n12958) );
  NAND2_X1 U7528 ( .A1(n11892), .A2(n11891), .ZN(n14909) );
  NAND2_X1 U7529 ( .A1(n8819), .A2(n8818), .ZN(n14210) );
  AND2_X1 U7530 ( .A1(n7045), .A2(n12940), .ZN(n12943) );
  OR2_X1 U7531 ( .A1(n12911), .A2(n12932), .ZN(n7633) );
  NAND2_X1 U7532 ( .A1(n11427), .A2(n12505), .ZN(n11447) );
  NAND2_X1 U7533 ( .A1(n7260), .A2(n7259), .ZN(n7044) );
  NAND2_X1 U7534 ( .A1(n7149), .A2(n7152), .ZN(n14829) );
  NAND2_X1 U7535 ( .A1(n8110), .A2(n8109), .ZN(n8124) );
  OR2_X1 U7536 ( .A1(n8098), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8110) );
  AND2_X1 U7537 ( .A1(n11313), .A2(n11312), .ZN(n11319) );
  INV_X1 U7538 ( .A(n11657), .ZN(n7149) );
  NAND2_X1 U7539 ( .A1(n10516), .A2(n10515), .ZN(n10760) );
  XNOR2_X1 U7540 ( .A(n8444), .B(SI_22_), .ZN(n8804) );
  OR2_X1 U7541 ( .A1(n8096), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8097) );
  OAI211_X1 U7542 ( .C1(n8791), .C2(n8440), .A(n7578), .B(n8442), .ZN(n8444)
         );
  NAND2_X1 U7543 ( .A1(n8734), .A2(n8733), .ZN(n14293) );
  XNOR2_X1 U7544 ( .A(n8759), .B(n8758), .ZN(n11843) );
  NAND2_X1 U7545 ( .A1(n11452), .A2(n11451), .ZN(n11746) );
  NAND2_X1 U7546 ( .A1(n8681), .A2(n8680), .ZN(n15119) );
  XNOR2_X1 U7547 ( .A(n8729), .B(n8728), .ZN(n11819) );
  NAND2_X1 U7548 ( .A1(n8697), .A2(n8696), .ZN(n14257) );
  XNOR2_X1 U7549 ( .A(n8439), .B(SI_20_), .ZN(n8779) );
  OR2_X1 U7550 ( .A1(n8752), .A2(n8431), .ZN(n8755) );
  AND2_X1 U7551 ( .A1(n7184), .A2(n6888), .ZN(n11664) );
  CLKBUF_X1 U7552 ( .A(n12752), .Z(n6828) );
  OAI21_X1 U7553 ( .B1(n8708), .B2(n7574), .A(n7572), .ZN(n8753) );
  XNOR2_X1 U7554 ( .A(n8708), .B(n8707), .ZN(n11814) );
  NAND2_X1 U7555 ( .A1(n7119), .A2(n15047), .ZN(n7732) );
  NAND2_X1 U7556 ( .A1(n6982), .A2(n8427), .ZN(n8708) );
  NAND2_X1 U7557 ( .A1(n7982), .A2(n7981), .ZN(n13740) );
  OR2_X1 U7558 ( .A1(n10920), .A2(n12202), .ZN(n15462) );
  OAI21_X1 U7559 ( .B1(n8009), .B2(n7243), .A(n7240), .ZN(n8042) );
  XNOR2_X1 U7560 ( .A(n11373), .B(n11374), .ZN(n11255) );
  OAI21_X1 U7561 ( .B1(n11080), .B2(n7190), .A(n7189), .ZN(n11338) );
  NAND2_X1 U7562 ( .A1(n8624), .A2(n8623), .ZN(n10906) );
  OR2_X1 U7563 ( .A1(n8422), .A2(n9707), .ZN(n8424) );
  NAND2_X1 U7564 ( .A1(n7114), .A2(n11299), .ZN(n12375) );
  NAND2_X1 U7565 ( .A1(n10839), .A2(n12491), .ZN(n10841) );
  OR2_X1 U7566 ( .A1(n8102), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8116) );
  XNOR2_X1 U7567 ( .A(n11232), .B(n11251), .ZN(n11080) );
  OAI21_X2 U7568 ( .B1(n9831), .B2(n10822), .A(n14852), .ZN(n9832) );
  NOR2_X1 U7569 ( .A1(n11078), .A2(n11077), .ZN(n11232) );
  NAND2_X1 U7570 ( .A1(n6752), .A2(n6641), .ZN(n7043) );
  AND2_X2 U7571 ( .A1(n14607), .A2(n14852), .ZN(n14855) );
  NAND2_X1 U7572 ( .A1(n10573), .A2(n10572), .ZN(n12351) );
  INV_X1 U7573 ( .A(n8259), .ZN(n12204) );
  NAND2_X1 U7574 ( .A1(n8590), .A2(n8589), .ZN(n10704) );
  NAND2_X1 U7575 ( .A1(n10329), .A2(n10312), .ZN(n10839) );
  NAND2_X1 U7576 ( .A1(n8576), .A2(n8575), .ZN(n15326) );
  NOR2_X1 U7577 ( .A1(n10447), .A2(n10446), .ZN(n11078) );
  INV_X2 U7578 ( .A(n12734), .ZN(n12771) );
  NAND2_X1 U7579 ( .A1(n8586), .A2(n8408), .ZN(n8601) );
  CLKBUF_X1 U7580 ( .A(n12664), .Z(n6812) );
  AND2_X1 U7581 ( .A1(n7053), .A2(n7052), .ZN(n11250) );
  INV_X1 U7582 ( .A(n15493), .ZN(n9975) );
  AND2_X1 U7583 ( .A1(n8315), .A2(n8314), .ZN(n13743) );
  INV_X1 U7584 ( .A(n6973), .ZN(n6969) );
  INV_X1 U7585 ( .A(n9799), .ZN(n9802) );
  OR2_X1 U7586 ( .A1(n8032), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8050) );
  CLKBUF_X1 U7587 ( .A(n12665), .Z(n6749) );
  NAND2_X1 U7588 ( .A1(n8519), .A2(n8518), .ZN(n9941) );
  XNOR2_X1 U7589 ( .A(n10158), .B(n9900), .ZN(n9906) );
  AND2_X1 U7590 ( .A1(n7090), .A2(n6974), .ZN(n6973) );
  NAND2_X2 U7591 ( .A1(n9797), .A2(n9796), .ZN(n12665) );
  CLKBUF_X3 U7592 ( .A(n11649), .Z(n12454) );
  NAND2_X1 U7593 ( .A1(n9797), .A2(n12300), .ZN(n9799) );
  NAND2_X1 U7594 ( .A1(n7834), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7767) );
  AOI22_X1 U7595 ( .A1(n10229), .A2(n15411), .B1(n10228), .B2(n10227), .ZN(
        n10238) );
  NAND4_X1 U7596 ( .A1(n8497), .A2(n8496), .A3(n8495), .A4(n8494), .ZN(n13915)
         );
  XOR2_X1 U7597 ( .A(n7653), .B(P3_ADDR_REG_5__SCAN_IN), .Z(n7718) );
  CLKBUF_X3 U7598 ( .A(n7831), .Z(n6606) );
  OR2_X1 U7599 ( .A1(n7999), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8016) );
  INV_X2 U7600 ( .A(n8478), .ZN(n9235) );
  NAND2_X1 U7601 ( .A1(n8309), .A2(n8310), .ZN(n11591) );
  CLKBUF_X3 U7602 ( .A(n8485), .Z(n8871) );
  NAND2_X1 U7603 ( .A1(n6602), .A2(n7274), .ZN(n8205) );
  NAND2_X1 U7604 ( .A1(n8313), .A2(n8312), .ZN(n11638) );
  AND2_X1 U7605 ( .A1(n12230), .A2(n10353), .ZN(n10354) );
  AND2_X2 U7606 ( .A1(n7321), .A2(n7317), .ZN(n9748) );
  AND2_X1 U7607 ( .A1(n8925), .A2(n6929), .ZN(n8937) );
  XNOR2_X1 U7608 ( .A(n7763), .B(P3_IR_REG_29__SCAN_IN), .ZN(n7765) );
  OR2_X1 U7609 ( .A1(n7323), .A2(n7322), .ZN(n7321) );
  AND2_X1 U7610 ( .A1(n8331), .A2(n12060), .ZN(n12228) );
  MUX2_X1 U7611 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8307), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8309) );
  AND2_X2 U7612 ( .A1(n12236), .A2(n10352), .ZN(n12183) );
  NAND2_X1 U7613 ( .A1(n10784), .A2(n13060), .ZN(n12230) );
  INV_X1 U7614 ( .A(n9775), .ZN(n12298) );
  NAND2_X1 U7615 ( .A1(n8373), .A2(n11773), .ZN(n8520) );
  XNOR2_X1 U7616 ( .A(n9519), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U7617 ( .A1(n9721), .A2(n9720), .ZN(n11695) );
  XNOR2_X1 U7618 ( .A(n7515), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8373) );
  NAND2_X1 U7619 ( .A1(n7630), .A2(n8926), .ZN(n11104) );
  OR2_X1 U7620 ( .A1(n14299), .A2(n14300), .ZN(n7515) );
  NAND2_X1 U7621 ( .A1(n8925), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8923) );
  XNOR2_X1 U7622 ( .A(n8763), .B(n8762), .ZN(n11795) );
  XNOR2_X1 U7623 ( .A(n7647), .B(n7126), .ZN(n7705) );
  INV_X2 U7624 ( .A(n14304), .ZN(n14312) );
  AND2_X1 U7625 ( .A1(n9714), .A2(n7359), .ZN(n9324) );
  XNOR2_X1 U7626 ( .A(n8248), .B(n7755), .ZN(n12060) );
  NAND2_X1 U7627 ( .A1(n7613), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U7628 ( .A1(n8908), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8464) );
  AND2_X2 U7629 ( .A1(n7165), .A2(n7477), .ZN(n8338) );
  NAND2_X1 U7630 ( .A1(n7646), .A2(n6775), .ZN(n7647) );
  NOR2_X1 U7631 ( .A1(n8760), .A2(n7394), .ZN(n6807) );
  AND3_X1 U7632 ( .A1(n7750), .A2(n7751), .A3(n6803), .ZN(n7165) );
  NOR2_X1 U7633 ( .A1(n8369), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n7550) );
  AND2_X2 U7634 ( .A1(n7160), .A2(n7058), .ZN(n7751) );
  AND2_X1 U7635 ( .A1(n7757), .A2(n7758), .ZN(n7481) );
  AND3_X1 U7636 ( .A1(n7075), .A2(n7074), .A3(n7076), .ZN(n7752) );
  AND2_X1 U7637 ( .A1(n10255), .A2(n9311), .ZN(n9314) );
  INV_X1 U7638 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8045) );
  NOR2_X1 U7639 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_12__SCAN_IN), .ZN(
        n7074) );
  NOR2_X1 U7640 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7076) );
  NOR2_X1 U7641 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n10257) );
  INV_X1 U7642 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9407) );
  INV_X4 U7643 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  XNOR2_X1 U7644 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n7708) );
  NOR2_X1 U7645 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n7075) );
  INV_X1 U7646 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7839) );
  NOR2_X1 U7647 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n7167) );
  INV_X1 U7648 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8065) );
  INV_X1 U7649 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8079) );
  INV_X1 U7650 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7753) );
  NOR2_X1 U7651 ( .A1(P3_IR_REG_5__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7749) );
  OAI21_X1 U7652 ( .B1(n13132), .B2(n13135), .A(n12169), .ZN(n6591) );
  INV_X1 U7653 ( .A(n10629), .ZN(n6592) );
  NAND2_X2 U7654 ( .A1(n12171), .A2(n12169), .ZN(n13135) );
  NAND2_X1 U7655 ( .A1(n14426), .A2(n10509), .ZN(n10516) );
  NAND2_X1 U7656 ( .A1(n6593), .A2(n14115), .ZN(n14085) );
  NOR2_X1 U7657 ( .A1(n14087), .A2(n14222), .ZN(n6593) );
  AND2_X1 U7658 ( .A1(n14248), .A2(n14266), .ZN(n6594) );
  AND2_X1 U7659 ( .A1(n6595), .A2(n7139), .ZN(n11622) );
  NOR2_X1 U7660 ( .A1(n14257), .A2(n15119), .ZN(n6595) );
  NOR2_X1 U7661 ( .A1(n13967), .A2(n6596), .ZN(n7136) );
  NOR2_X1 U7662 ( .A1(n14126), .A2(n14116), .ZN(n14115) );
  MUX2_X1 U7663 ( .A(n7135), .B(P2_REG1_REG_30__SCAN_IN), .S(n6794), .Z(n14177) );
  NAND2_X1 U7664 ( .A1(n12262), .A2(n6600), .ZN(n6597) );
  OR2_X1 U7665 ( .A1(n6599), .A2(n7169), .ZN(n6598) );
  INV_X1 U7666 ( .A(n7168), .ZN(n6599) );
  AND2_X1 U7667 ( .A1(n12261), .A2(n7168), .ZN(n6600) );
  NAND2_X1 U7668 ( .A1(n12877), .A2(n12876), .ZN(n6601) );
  NAND2_X1 U7669 ( .A1(n12877), .A2(n12876), .ZN(n12875) );
  NAND2_X2 U7670 ( .A1(n7812), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7766) );
  OAI222_X1 U7671 ( .A1(P3_U3151), .A2(n12610), .B1(n12609), .B2(n12608), .C1(
        n13756), .C2(n12607), .ZN(P3_U3265) );
  NAND2_X1 U7672 ( .A1(n15607), .A2(n7721), .ZN(n7725) );
  NAND2_X2 U7673 ( .A1(n7180), .A2(n12247), .ZN(n12829) );
  NAND2_X1 U7674 ( .A1(n7305), .A2(n7307), .ZN(n11427) );
  AOI21_X2 U7675 ( .B1(n14650), .B2(n14649), .A(n11940), .ZN(n14626) );
  OAI21_X2 U7676 ( .B1(n10841), .B2(n12493), .A(n7302), .ZN(n11060) );
  NOR2_X4 U7677 ( .A1(n6630), .A2(n7271), .ZN(n12308) );
  OR2_X1 U7679 ( .A1(n7762), .A2(n7976), .ZN(n7763) );
  AND2_X4 U7680 ( .A1(n8338), .A2(n7088), .ZN(n8308) );
  NOR2_X2 U7681 ( .A1(n10684), .A2(n10372), .ZN(n10543) );
  AND4_X4 U7682 ( .A1(n7769), .A2(n7768), .A3(n7767), .A4(n7766), .ZN(n15493)
         );
  NAND2_X1 U7683 ( .A1(n9425), .A2(n7620), .ZN(n9236) );
  MUX2_X2 U7684 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14315), .S(n9425), .Z(n10143)
         );
  NAND2_X1 U7685 ( .A1(n11034), .A2(n11033), .ZN(n11170) );
  NAND2_X1 U7686 ( .A1(n8297), .A2(n8298), .ZN(n6602) );
  NAND2_X1 U7687 ( .A1(n10179), .A2(n9750), .ZN(n6603) );
  NAND2_X2 U7688 ( .A1(n10142), .A2(n11104), .ZN(n9914) );
  INV_X1 U7689 ( .A(n12734), .ZN(n6604) );
  INV_X1 U7690 ( .A(n12734), .ZN(n6605) );
  NAND2_X4 U7691 ( .A1(n10355), .A2(n10354), .ZN(n12734) );
  OAI222_X1 U7692 ( .A1(P3_U3151), .A2(n10784), .B1(n12609), .B2(n10783), .C1(
        n13756), .C2(n10782), .ZN(P3_U3275) );
  NAND2_X2 U7693 ( .A1(n7449), .A2(n12068), .ZN(n10359) );
  NAND2_X2 U7694 ( .A1(n9975), .A2(n8254), .ZN(n7449) );
  AND2_X1 U7695 ( .A1(n13754), .A2(n7764), .ZN(n6608) );
  INV_X1 U7696 ( .A(n6608), .ZN(n6609) );
  AND2_X1 U7697 ( .A1(n9022), .A2(n9021), .ZN(n9032) );
  OR2_X1 U7698 ( .A1(n13674), .A2(n12890), .ZN(n12135) );
  INV_X1 U7699 ( .A(n12060), .ZN(n10352) );
  NAND2_X1 U7700 ( .A1(n7390), .A2(n7392), .ZN(n7389) );
  OR2_X1 U7701 ( .A1(n13175), .A2(n13186), .ZN(n13148) );
  NOR2_X1 U7702 ( .A1(n6679), .A2(n7070), .ZN(n7069) );
  INV_X1 U7703 ( .A(n8291), .ZN(n7070) );
  OR2_X1 U7704 ( .A1(n13242), .A2(n13222), .ZN(n12139) );
  AND2_X1 U7705 ( .A1(n13865), .A2(n12558), .ZN(n7392) );
  NAND2_X1 U7706 ( .A1(n14049), .A2(n6649), .ZN(n6855) );
  NAND2_X1 U7707 ( .A1(n14048), .A2(n8840), .ZN(n7609) );
  NAND2_X1 U7708 ( .A1(n8790), .A2(n8789), .ZN(n14093) );
  NOR2_X1 U7709 ( .A1(n6678), .A2(n7615), .ZN(n7614) );
  OAI21_X1 U7710 ( .B1(n9032), .B2(n9033), .A(n9031), .ZN(n9035) );
  INV_X1 U7711 ( .A(n12334), .ZN(n12335) );
  NAND2_X1 U7712 ( .A1(n7419), .A2(n7418), .ZN(n7416) );
  NOR2_X1 U7713 ( .A1(n7419), .A2(n7418), .ZN(n7417) );
  INV_X1 U7714 ( .A(n9080), .ZN(n6915) );
  NAND2_X1 U7715 ( .A1(n12398), .A2(n7430), .ZN(n7429) );
  INV_X1 U7716 ( .A(n12388), .ZN(n7430) );
  OAI22_X1 U7717 ( .A1(n12377), .A2(n7448), .B1(n7447), .B2(n12378), .ZN(
        n12384) );
  INV_X1 U7718 ( .A(n12376), .ZN(n7447) );
  NOR2_X1 U7719 ( .A1(n12379), .A2(n12376), .ZN(n7448) );
  INV_X1 U7720 ( .A(n12418), .ZN(n7412) );
  INV_X1 U7721 ( .A(n6920), .ZN(n6918) );
  AOI21_X1 U7722 ( .B1(n7572), .B2(n7569), .A(n7568), .ZN(n7567) );
  NOR2_X1 U7723 ( .A1(n7575), .A2(n8437), .ZN(n7569) );
  INV_X1 U7724 ( .A(n8411), .ZN(n7094) );
  XNOR2_X1 U7725 ( .A(n10444), .B(n10307), .ZN(n10301) );
  INV_X1 U7726 ( .A(n11359), .ZN(n7186) );
  NOR2_X1 U7727 ( .A1(n13033), .A2(n13034), .ZN(n13036) );
  OR2_X1 U7728 ( .A1(n8343), .A2(n13094), .ZN(n12186) );
  OR2_X1 U7729 ( .A1(n13096), .A2(n13111), .ZN(n8295) );
  OR2_X1 U7730 ( .A1(n13108), .A2(n8217), .ZN(n7476) );
  OR2_X1 U7731 ( .A1(n12870), .A2(n13110), .ZN(n13103) );
  OR2_X1 U7732 ( .A1(n13187), .A2(n13197), .ZN(n12160) );
  NAND2_X1 U7733 ( .A1(n8056), .A2(n12135), .ZN(n13239) );
  OAI21_X1 U7734 ( .B1(n7946), .B2(n7233), .A(n7231), .ZN(n7972) );
  INV_X1 U7735 ( .A(n7232), .ZN(n7231) );
  OAI21_X1 U7736 ( .B1(n7238), .B2(n7233), .A(n7969), .ZN(n7232) );
  INV_X1 U7737 ( .A(n7235), .ZN(n7233) );
  INV_X1 U7738 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7747) );
  NAND2_X1 U7739 ( .A1(n9351), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7843) );
  NAND2_X1 U7740 ( .A1(n13807), .A2(n6763), .ZN(n12579) );
  NAND2_X1 U7741 ( .A1(n12568), .A2(n6764), .ZN(n6763) );
  INV_X1 U7742 ( .A(n12569), .ZN(n6764) );
  AND2_X1 U7743 ( .A1(n8372), .A2(n8373), .ZN(n8485) );
  NAND2_X1 U7744 ( .A1(n7494), .A2(n7496), .ZN(n6821) );
  XNOR2_X1 U7745 ( .A(n10890), .B(n13908), .ZN(n9283) );
  NOR2_X1 U7746 ( .A1(n6957), .A2(n6956), .ZN(n13979) );
  INV_X1 U7747 ( .A(n12701), .ZN(n7357) );
  INV_X1 U7748 ( .A(n11841), .ZN(n7106) );
  AOI21_X1 U7749 ( .B1(n7092), .B2(n7094), .A(n7091), .ZN(n7090) );
  INV_X1 U7750 ( .A(n8414), .ZN(n7091) );
  OAI21_X1 U7751 ( .B1(n7274), .B2(n9409), .A(n6778), .ZN(n8409) );
  NAND2_X1 U7752 ( .A1(n7274), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U7753 ( .A1(n8409), .A2(SI_9_), .ZN(n8411) );
  NAND2_X1 U7754 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6776), .ZN(n6775) );
  NAND2_X1 U7755 ( .A1(n7707), .A2(n7706), .ZN(n7646) );
  INV_X1 U7756 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6776) );
  OAI21_X1 U7757 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n7663), .A(n7662), .ZN(
        n7701) );
  INV_X1 U7758 ( .A(n8157), .ZN(n8156) );
  NAND2_X1 U7759 ( .A1(n13743), .A2(n12228), .ZN(n10355) );
  INV_X2 U7760 ( .A(n7868), .ZN(n12030) );
  INV_X1 U7761 ( .A(n7812), .ZN(n7868) );
  NAND2_X1 U7762 ( .A1(n6885), .A2(n6628), .ZN(n6884) );
  INV_X1 U7763 ( .A(n11338), .ZN(n6885) );
  NAND2_X1 U7764 ( .A1(n11338), .A2(n11259), .ZN(n6881) );
  OR2_X1 U7765 ( .A1(n12900), .A2(n12899), .ZN(n12901) );
  NAND2_X1 U7766 ( .A1(n12907), .A2(n12908), .ZN(n12931) );
  AND2_X1 U7767 ( .A1(n6880), .A2(n6879), .ZN(n12949) );
  INV_X1 U7768 ( .A(n12927), .ZN(n6879) );
  OR2_X1 U7769 ( .A1(n12952), .A2(n12953), .ZN(n7263) );
  AND2_X1 U7770 ( .A1(n13168), .A2(n6650), .ZN(n7067) );
  NAND2_X1 U7771 ( .A1(n13667), .A2(n6666), .ZN(n13224) );
  OAI21_X1 U7772 ( .B1(n13260), .B2(n8280), .A(n8279), .ZN(n13245) );
  AOI21_X1 U7773 ( .B1(n7010), .B2(n7013), .A(n7008), .ZN(n7007) );
  INV_X1 U7774 ( .A(n12107), .ZN(n7008) );
  INV_X1 U7775 ( .A(n12040), .ZN(n8082) );
  NAND2_X1 U7776 ( .A1(n12058), .A2(n12060), .ZN(n15559) );
  INV_X1 U7777 ( .A(n15517), .ZN(n15494) );
  NAND2_X1 U7778 ( .A1(n8126), .A2(n8125), .ZN(n8140) );
  NAND2_X1 U7779 ( .A1(n8124), .A2(n8123), .ZN(n8126) );
  AND2_X1 U7780 ( .A1(n8095), .A2(n8078), .ZN(n8093) );
  NAND2_X1 U7781 ( .A1(n8009), .A2(n7249), .ZN(n7246) );
  OAI21_X1 U7782 ( .B1(n7389), .B2(n7383), .A(n7388), .ZN(n6938) );
  INV_X1 U7783 ( .A(n13840), .ZN(n7383) );
  NAND2_X1 U7784 ( .A1(n7390), .A2(n7391), .ZN(n7388) );
  INV_X1 U7785 ( .A(n6730), .ZN(n6936) );
  AND2_X1 U7786 ( .A1(n8938), .A2(n6585), .ZN(n9921) );
  OR2_X1 U7787 ( .A1(n13850), .A2(n12591), .ZN(n7377) );
  NAND2_X1 U7788 ( .A1(n6807), .A2(n6806), .ZN(n8925) );
  INV_X1 U7789 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6806) );
  AOI21_X1 U7790 ( .B1(n7607), .B2(n7606), .A(n6647), .ZN(n7605) );
  INV_X1 U7791 ( .A(n8840), .ZN(n7606) );
  NAND2_X1 U7792 ( .A1(n14079), .A2(n7611), .ZN(n14061) );
  AND2_X1 U7793 ( .A1(n14068), .A2(n8814), .ZN(n7611) );
  NAND2_X1 U7794 ( .A1(n14093), .A2(n14095), .ZN(n6857) );
  NAND2_X1 U7795 ( .A1(n7491), .A2(n6654), .ZN(n7488) );
  NOR2_X1 U7796 ( .A1(n7618), .A2(n8776), .ZN(n7617) );
  INV_X1 U7797 ( .A(n8750), .ZN(n7618) );
  AND2_X1 U7798 ( .A1(n7595), .A2(n6863), .ZN(n6862) );
  OR2_X1 U7799 ( .A1(n7597), .A2(n8705), .ZN(n6863) );
  NAND2_X1 U7800 ( .A1(n7596), .A2(n8741), .ZN(n7595) );
  INV_X1 U7801 ( .A(n7598), .ZN(n7596) );
  NAND2_X1 U7802 ( .A1(n8726), .A2(n8741), .ZN(n7597) );
  OAI21_X1 U7803 ( .B1(n11184), .B2(n8673), .A(n8674), .ZN(n15118) );
  NOR2_X1 U7804 ( .A1(n15134), .A2(n6959), .ZN(n6958) );
  INV_X1 U7805 ( .A(n8954), .ZN(n6959) );
  NAND2_X1 U7806 ( .A1(n15352), .A2(n8935), .ZN(n14147) );
  NAND2_X1 U7807 ( .A1(n7512), .A2(n7612), .ZN(n7613) );
  NAND2_X1 U7808 ( .A1(n7334), .A2(n7337), .ZN(n14338) );
  AND2_X1 U7809 ( .A1(n7338), .A2(n12648), .ZN(n7337) );
  AND2_X1 U7810 ( .A1(n14316), .A2(n7356), .ZN(n7355) );
  OR2_X1 U7811 ( .A1(n14437), .A2(n7357), .ZN(n7356) );
  NAND2_X1 U7812 ( .A1(n14395), .A2(n6719), .ZN(n14347) );
  AND2_X1 U7813 ( .A1(n15034), .A2(n9775), .ZN(n12293) );
  OR2_X1 U7814 ( .A1(n12523), .A2(n12522), .ZN(n6788) );
  AND2_X1 U7815 ( .A1(n12514), .A2(n11901), .ZN(n7324) );
  NAND2_X1 U7816 ( .A1(n7151), .A2(n7150), .ZN(n11657) );
  INV_X1 U7817 ( .A(n11746), .ZN(n7150) );
  INV_X1 U7818 ( .A(n7281), .ZN(n7280) );
  NAND2_X1 U7819 ( .A1(n9751), .A2(n9750), .ZN(n11448) );
  NAND2_X1 U7820 ( .A1(n9766), .A2(n12455), .ZN(n14939) );
  INV_X2 U7821 ( .A(n11448), .ZN(n12456) );
  AND2_X1 U7822 ( .A1(n14789), .A2(n14946), .ZN(n15229) );
  AND2_X2 U7823 ( .A1(n9717), .A2(n9316), .ZN(n9714) );
  INV_X1 U7824 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9316) );
  OAI21_X1 U7825 ( .B1(n15049), .B2(n15048), .A(n7120), .ZN(n7119) );
  INV_X1 U7826 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7120) );
  INV_X1 U7827 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n13070) );
  NAND2_X1 U7828 ( .A1(n8143), .A2(n8142), .ZN(n13175) );
  NAND2_X1 U7829 ( .A1(n15049), .A2(n15048), .ZN(n15047) );
  NAND2_X1 U7830 ( .A1(n15185), .A2(n15186), .ZN(n15184) );
  NAND2_X1 U7831 ( .A1(n7408), .A2(n7407), .ZN(n12310) );
  AOI21_X1 U7832 ( .B1(n7417), .B2(n7416), .A(n7414), .ZN(n7413) );
  NAND2_X1 U7833 ( .A1(n6902), .A2(n9051), .ZN(n6901) );
  INV_X1 U7834 ( .A(n7449), .ZN(n12064) );
  NAND2_X1 U7835 ( .A1(n12368), .A2(n12365), .ZN(n7435) );
  NOR2_X1 U7836 ( .A1(n12368), .A2(n12365), .ZN(n7436) );
  INV_X1 U7837 ( .A(n9085), .ZN(n6909) );
  NAND2_X1 U7838 ( .A1(n6907), .A2(n6615), .ZN(n6906) );
  INV_X1 U7839 ( .A(n6911), .ZN(n6907) );
  NAND2_X1 U7840 ( .A1(n6635), .A2(n6915), .ZN(n6913) );
  NOR2_X1 U7841 ( .A1(n6914), .A2(n6912), .ZN(n6911) );
  NOR2_X1 U7842 ( .A1(n9076), .A2(n7532), .ZN(n6912) );
  NOR2_X1 U7843 ( .A1(n6635), .A2(n6915), .ZN(n6914) );
  OR2_X1 U7844 ( .A1(n9071), .A2(n9070), .ZN(n9077) );
  AOI21_X1 U7845 ( .B1(n9069), .B2(n9068), .A(n9067), .ZN(n9071) );
  INV_X1 U7846 ( .A(n12404), .ZN(n7428) );
  NAND2_X1 U7847 ( .A1(n6692), .A2(n7429), .ZN(n7425) );
  INV_X1 U7848 ( .A(n12386), .ZN(n7431) );
  AND3_X1 U7849 ( .A1(n14788), .A2(n6620), .A3(n11652), .ZN(n6813) );
  OAI21_X1 U7850 ( .B1(n12384), .B2(n12383), .A(n12382), .ZN(n6994) );
  INV_X1 U7851 ( .A(n12407), .ZN(n6990) );
  NAND2_X1 U7852 ( .A1(n6926), .A2(n6715), .ZN(n6924) );
  NOR2_X1 U7853 ( .A1(n6926), .A2(n6715), .ZN(n6925) );
  OAI22_X1 U7854 ( .A1(n7552), .A2(n9084), .B1(n9093), .B2(n9092), .ZN(n9097)
         );
  NAND2_X1 U7855 ( .A1(n6691), .A2(n7549), .ZN(n7548) );
  INV_X1 U7856 ( .A(n12414), .ZN(n6782) );
  NAND2_X1 U7857 ( .A1(n7537), .A2(n7536), .ZN(n7535) );
  NAND2_X1 U7858 ( .A1(n7519), .A2(n7516), .ZN(n9129) );
  NAND2_X1 U7859 ( .A1(n7521), .A2(n7520), .ZN(n7519) );
  AND2_X1 U7860 ( .A1(n9128), .A2(n9127), .ZN(n6923) );
  NOR2_X1 U7861 ( .A1(n9133), .A2(n6716), .ZN(n7537) );
  NAND2_X1 U7862 ( .A1(n9133), .A2(n6716), .ZN(n7536) );
  OR2_X1 U7863 ( .A1(n12431), .A2(n7442), .ZN(n6780) );
  NAND2_X1 U7864 ( .A1(n7441), .A2(n12430), .ZN(n7440) );
  NOR2_X1 U7865 ( .A1(n7441), .A2(n12430), .ZN(n7442) );
  NAND2_X1 U7866 ( .A1(n6748), .A2(n8275), .ZN(n8273) );
  NAND2_X1 U7867 ( .A1(n9148), .A2(n9147), .ZN(n6917) );
  NOR2_X1 U7868 ( .A1(n6636), .A2(n7529), .ZN(n7528) );
  NOR2_X1 U7869 ( .A1(n9225), .A2(n9215), .ZN(n9255) );
  NAND2_X1 U7870 ( .A1(n6636), .A2(n7529), .ZN(n7527) );
  NAND2_X1 U7871 ( .A1(n12299), .A2(n12298), .ZN(n12462) );
  INV_X1 U7872 ( .A(n8630), .ZN(n6974) );
  INV_X1 U7873 ( .A(n8270), .ZN(n7085) );
  AOI21_X1 U7874 ( .B1(n8139), .B2(n8141), .A(n7255), .ZN(n7254) );
  INV_X1 U7875 ( .A(n8150), .ZN(n7255) );
  INV_X1 U7876 ( .A(n8141), .ZN(n7252) );
  NOR2_X1 U7877 ( .A1(n8949), .A2(n7498), .ZN(n7497) );
  INV_X1 U7878 ( .A(n8948), .ZN(n7498) );
  NOR2_X1 U7879 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n8362) );
  NOR2_X1 U7880 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8361) );
  NOR2_X1 U7881 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8359) );
  NOR2_X1 U7882 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8360) );
  INV_X1 U7883 ( .A(n12469), .ZN(n7423) );
  AOI21_X1 U7884 ( .B1(n7575), .B2(n7573), .A(n6680), .ZN(n7572) );
  INV_X1 U7885 ( .A(n8707), .ZN(n7573) );
  NAND2_X1 U7886 ( .A1(n8423), .A2(n7593), .ZN(n7592) );
  NOR2_X1 U7887 ( .A1(n7474), .A2(n7473), .ZN(n7472) );
  AND2_X1 U7888 ( .A1(n7262), .A2(n7261), .ZN(n11373) );
  NAND2_X1 U7889 ( .A1(n11254), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7261) );
  AND2_X1 U7890 ( .A1(n12955), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7264) );
  NAND2_X1 U7891 ( .A1(n8176), .A2(n8175), .ZN(n8192) );
  INV_X1 U7892 ( .A(n12130), .ZN(n7005) );
  OAI21_X1 U7893 ( .B1(n13558), .B2(n7005), .A(n13259), .ZN(n7004) );
  INV_X1 U7894 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7775) );
  INV_X1 U7895 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7774) );
  AND2_X1 U7896 ( .A1(n12116), .A2(n13574), .ZN(n8271) );
  INV_X1 U7897 ( .A(n7018), .ZN(n7017) );
  OAI21_X1 U7898 ( .B1(n12207), .B2(n7019), .A(n12096), .ZN(n7018) );
  INV_X1 U7899 ( .A(n12090), .ZN(n7019) );
  NAND2_X1 U7900 ( .A1(n10631), .A2(n15495), .ZN(n12070) );
  INV_X1 U7901 ( .A(n7249), .ZN(n7242) );
  NOR2_X1 U7902 ( .A1(n8022), .A2(n7250), .ZN(n7249) );
  AND2_X1 U7903 ( .A1(n10265), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8022) );
  INV_X1 U7904 ( .A(n8008), .ZN(n7250) );
  NOR2_X1 U7905 ( .A1(n7957), .A2(n7239), .ZN(n7238) );
  INV_X1 U7906 ( .A(n7945), .ZN(n7239) );
  NOR2_X1 U7907 ( .A1(n9451), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7236) );
  AOI21_X1 U7908 ( .B1(n7224), .B2(n7222), .A(n6689), .ZN(n7221) );
  INV_X1 U7909 ( .A(n7226), .ZN(n7222) );
  NOR2_X1 U7910 ( .A1(n7804), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n7861) );
  XNOR2_X1 U7911 ( .A(n15326), .B(n12592), .ZN(n6940) );
  AND2_X1 U7912 ( .A1(n7505), .A2(n9278), .ZN(n7504) );
  OR2_X1 U7913 ( .A1(n14023), .A2(n7506), .ZN(n7505) );
  INV_X1 U7914 ( .A(n8974), .ZN(n7506) );
  NOR2_X1 U7915 ( .A1(n8967), .A2(n7490), .ZN(n7489) );
  INV_X1 U7916 ( .A(n8966), .ZN(n7490) );
  INV_X1 U7917 ( .A(n6946), .ZN(n6945) );
  OAI21_X1 U7918 ( .B1(n6949), .B2(n6947), .A(n8961), .ZN(n6946) );
  INV_X1 U7919 ( .A(n6948), .ZN(n6947) );
  NAND2_X1 U7920 ( .A1(n10606), .A2(n6662), .ZN(n10694) );
  INV_X1 U7921 ( .A(n8540), .ZN(n7604) );
  INV_X1 U7922 ( .A(n8525), .ZN(n7603) );
  OR2_X1 U7923 ( .A1(n9949), .A2(n10138), .ZN(n9946) );
  NAND2_X1 U7924 ( .A1(n7508), .A2(n7507), .ZN(n11630) );
  AOI21_X1 U7925 ( .B1(n7509), .B2(n8958), .A(n6673), .ZN(n7507) );
  OAI21_X1 U7926 ( .B1(n8925), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U7927 ( .A1(n8761), .A2(n8762), .ZN(n7396) );
  INV_X1 U7928 ( .A(n12709), .ZN(n12664) );
  NAND2_X1 U7929 ( .A1(n14734), .A2(n7286), .ZN(n7285) );
  INV_X1 U7930 ( .A(n11970), .ZN(n7286) );
  NOR2_X1 U7931 ( .A1(n12511), .A2(n7288), .ZN(n7287) );
  INV_X1 U7932 ( .A(n11968), .ZN(n7288) );
  INV_X1 U7933 ( .A(n11828), .ZN(n7112) );
  INV_X1 U7934 ( .A(n11639), .ZN(n7097) );
  OR2_X1 U7935 ( .A1(n14967), .A2(n14823), .ZN(n12388) );
  NOR2_X1 U7936 ( .A1(n7309), .A2(n12501), .ZN(n7306) );
  INV_X1 U7937 ( .A(n10313), .ZN(n7303) );
  NAND2_X1 U7938 ( .A1(n10311), .A2(n10310), .ZN(n10330) );
  NOR2_X1 U7939 ( .A1(n12394), .A2(n7294), .ZN(n7293) );
  INV_X1 U7940 ( .A(n11966), .ZN(n7294) );
  NAND2_X1 U7941 ( .A1(n7320), .A2(n9744), .ZN(n7318) );
  INV_X1 U7942 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7320) );
  NOR2_X1 U7943 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), .ZN(
        n7319) );
  INV_X1 U7944 ( .A(n7583), .ZN(n7582) );
  OAI21_X1 U7945 ( .B1(n8879), .B2(n7584), .A(n8460), .ZN(n7583) );
  INV_X1 U7946 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9742) );
  AOI21_X1 U7947 ( .B1(n7564), .B2(n7566), .A(n6733), .ZN(n7562) );
  NOR2_X1 U7948 ( .A1(n8791), .A2(n8778), .ZN(n7579) );
  AOI21_X1 U7949 ( .B1(n7556), .B2(n7558), .A(n6688), .ZN(n7554) );
  INV_X1 U7950 ( .A(n7093), .ZN(n7092) );
  OAI21_X1 U7951 ( .B1(n8600), .B2(n7094), .A(n8413), .ZN(n7093) );
  NAND2_X1 U7952 ( .A1(n8385), .A2(SI_2_), .ZN(n8510) );
  OAI21_X1 U7953 ( .B1(n8387), .B2(n9753), .A(n7594), .ZN(n8380) );
  NAND2_X1 U7954 ( .A1(n8387), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7594) );
  OAI21_X1 U7955 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n7670), .A(n7669), .ZN(
        n7696) );
  INV_X1 U7956 ( .A(n11543), .ZN(n6756) );
  OR2_X1 U7957 ( .A1(n12814), .A2(n12265), .ZN(n7170) );
  NOR3_X1 U7958 ( .A1(n12189), .A2(n12188), .A3(n12187), .ZN(n12194) );
  MUX2_X1 U7959 ( .A(n12185), .B(n12184), .S(n12183), .Z(n12189) );
  OAI21_X1 U7960 ( .B1(n7461), .B2(n12235), .A(n12237), .ZN(n7457) );
  INV_X1 U7961 ( .A(n8162), .ZN(n12029) );
  OR2_X1 U7962 ( .A1(n10196), .A2(n10195), .ZN(n7181) );
  NAND2_X1 U7963 ( .A1(n7192), .A2(n10224), .ZN(n7194) );
  INV_X1 U7964 ( .A(n10207), .ZN(n7055) );
  AOI21_X1 U7965 ( .B1(n10240), .B2(n10206), .A(n7258), .ZN(n10207) );
  AOI21_X1 U7966 ( .B1(n10437), .B2(n7050), .A(n10439), .ZN(n7049) );
  NAND2_X1 U7967 ( .A1(n10295), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10438) );
  NOR2_X1 U7968 ( .A1(n10445), .A2(n7642), .ZN(n10447) );
  NAND2_X1 U7969 ( .A1(n7043), .A2(n7042), .ZN(n7262) );
  INV_X1 U7970 ( .A(n11347), .ZN(n7042) );
  NOR2_X1 U7971 ( .A1(n11338), .A2(n6887), .ZN(n11355) );
  NOR2_X1 U7972 ( .A1(n7185), .A2(n6883), .ZN(n6882) );
  NAND2_X1 U7973 ( .A1(n7186), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7185) );
  INV_X1 U7974 ( .A(n6886), .ZN(n6883) );
  NAND2_X1 U7975 ( .A1(n11671), .A2(n11672), .ZN(n11673) );
  NAND2_X1 U7976 ( .A1(n11673), .A2(n11674), .ZN(n11763) );
  NAND2_X1 U7977 ( .A1(n6878), .A2(n12922), .ZN(n6880) );
  INV_X1 U7978 ( .A(n12934), .ZN(n6842) );
  XNOR2_X1 U7979 ( .A(n12991), .B(n12992), .ZN(n12952) );
  OR2_X1 U7980 ( .A1(n13004), .A2(n6893), .ZN(n6890) );
  OR2_X1 U7981 ( .A1(n13031), .A2(n13003), .ZN(n6893) );
  NAND2_X1 U7982 ( .A1(n13030), .A2(n6892), .ZN(n6891) );
  INV_X1 U7983 ( .A(n13031), .ZN(n6892) );
  INV_X1 U7984 ( .A(n7030), .ZN(n13106) );
  INV_X1 U7985 ( .A(n13152), .ZN(n13122) );
  OAI21_X1 U7986 ( .B1(n13122), .B2(n13711), .A(n13134), .ZN(n13121) );
  INV_X1 U7987 ( .A(n12196), .ZN(n13182) );
  AND2_X1 U7988 ( .A1(n8282), .A2(n8281), .ZN(n7065) );
  AND2_X1 U7989 ( .A1(n12125), .A2(n12130), .ZN(n13558) );
  INV_X1 U7990 ( .A(n13571), .ZN(n15068) );
  INV_X1 U7991 ( .A(n12893), .ZN(n15452) );
  NAND2_X1 U7992 ( .A1(n11015), .A2(n12207), .ZN(n11017) );
  INV_X1 U7993 ( .A(n11171), .ZN(n12207) );
  OR2_X1 U7994 ( .A1(n6603), .A2(n9375), .ZN(n7828) );
  NAND2_X1 U7995 ( .A1(n12070), .A2(n12071), .ZN(n15477) );
  NOR2_X1 U7996 ( .A1(n10182), .A2(n15559), .ZN(n10488) );
  AND2_X1 U7997 ( .A1(n8304), .A2(n12183), .ZN(n15517) );
  NAND2_X1 U7998 ( .A1(n8101), .A2(n8100), .ZN(n12271) );
  OR2_X1 U7999 ( .A1(n10782), .A2(n7819), .ZN(n8101) );
  INV_X1 U8000 ( .A(n13239), .ZN(n7027) );
  NAND2_X1 U8001 ( .A1(n8013), .A2(n8012), .ZN(n13680) );
  AND2_X1 U8002 ( .A1(n7178), .A2(n8337), .ZN(n9532) );
  NAND2_X1 U8003 ( .A1(n8234), .A2(n8233), .ZN(n12022) );
  XNOR2_X1 U8004 ( .A(n8247), .B(n8246), .ZN(n12058) );
  INV_X1 U8005 ( .A(n7754), .ZN(n7480) );
  AND2_X1 U8006 ( .A1(n8076), .A2(n8059), .ZN(n8060) );
  NAND2_X1 U8007 ( .A1(n8058), .A2(n8057), .ZN(n8061) );
  NAND2_X1 U8008 ( .A1(n8061), .A2(n8060), .ZN(n8077) );
  NAND2_X1 U8009 ( .A1(n8042), .A2(n8041), .ZN(n8058) );
  AND2_X1 U8010 ( .A1(n7245), .A2(n7247), .ZN(n7244) );
  INV_X1 U8011 ( .A(n8025), .ZN(n7245) );
  NAND2_X1 U8012 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n7248), .ZN(n7247) );
  NAND2_X1 U8013 ( .A1(n8007), .A2(n8006), .ZN(n8009) );
  NAND2_X1 U8014 ( .A1(n7992), .A2(n7991), .ZN(n8007) );
  NOR2_X1 U8015 ( .A1(n7960), .A2(n7236), .ZN(n7235) );
  NAND2_X1 U8016 ( .A1(n7946), .A2(n7238), .ZN(n7237) );
  INV_X1 U8017 ( .A(n7236), .ZN(n7234) );
  INV_X1 U8018 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7963) );
  AOI21_X1 U8019 ( .B1(n7226), .B2(n7878), .A(n7225), .ZN(n7224) );
  INV_X1 U8020 ( .A(n7897), .ZN(n7225) );
  OR2_X1 U8021 ( .A1(n7879), .A2(n7878), .ZN(n7230) );
  NAND2_X1 U8022 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n7229), .ZN(n7228) );
  INV_X1 U8023 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7229) );
  AND2_X1 U8024 ( .A1(n7227), .A2(n7228), .ZN(n7226) );
  INV_X1 U8025 ( .A(n7881), .ZN(n7227) );
  NAND2_X1 U8026 ( .A1(n7214), .A2(n7843), .ZN(n7213) );
  OR2_X1 U8027 ( .A1(n7820), .A2(n7216), .ZN(n7215) );
  OR2_X1 U8028 ( .A1(n7861), .A2(n7976), .ZN(n7840) );
  AND2_X1 U8029 ( .A1(n7218), .A2(n7822), .ZN(n7217) );
  INV_X1 U8030 ( .A(n7824), .ZN(n7218) );
  NAND2_X1 U8031 ( .A1(n7821), .A2(n7636), .ZN(n7219) );
  NAND2_X1 U8032 ( .A1(n9342), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7793) );
  XNOR2_X1 U8033 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7792) );
  OR2_X1 U8034 ( .A1(n13759), .A2(n13758), .ZN(n13760) );
  INV_X1 U8035 ( .A(n6935), .ZN(n6934) );
  OAI21_X1 U8036 ( .B1(n10388), .B2(n7380), .A(n7378), .ZN(n7381) );
  AND2_X1 U8037 ( .A1(n7379), .A2(n10872), .ZN(n7378) );
  OR2_X1 U8038 ( .A1(n10387), .A2(n7380), .ZN(n7379) );
  INV_X1 U8039 ( .A(n10640), .ZN(n7380) );
  INV_X1 U8040 ( .A(n7389), .ZN(n7385) );
  NAND2_X1 U8041 ( .A1(n15103), .A2(n12549), .ZN(n12550) );
  NAND2_X1 U8042 ( .A1(n9267), .A2(n9266), .ZN(n9275) );
  AOI21_X1 U8043 ( .B1(n6610), .B2(n7605), .A(n6674), .ZN(n6856) );
  NAND2_X1 U8044 ( .A1(n14024), .A2(n14023), .ZN(n14022) );
  NAND2_X1 U8045 ( .A1(n14061), .A2(n8827), .ZN(n14049) );
  NAND2_X1 U8046 ( .A1(n7610), .A2(n9291), .ZN(n14051) );
  INV_X1 U8047 ( .A(n14049), .ZN(n7610) );
  NAND2_X1 U8048 ( .A1(n6857), .A2(n6663), .ZN(n14079) );
  NAND2_X1 U8049 ( .A1(n14109), .A2(n7489), .ZN(n7483) );
  NAND2_X1 U8050 ( .A1(n7486), .A2(n7488), .ZN(n7485) );
  INV_X1 U8051 ( .A(n7489), .ZN(n7486) );
  INV_X1 U8052 ( .A(n7488), .ZN(n7487) );
  OAI21_X1 U8053 ( .B1(n14132), .B2(n8962), .A(n8963), .ZN(n14110) );
  AOI21_X1 U8054 ( .B1(n6862), .B2(n7597), .A(n6860), .ZN(n6859) );
  INV_X1 U8055 ( .A(n14142), .ZN(n6860) );
  NAND2_X1 U8056 ( .A1(n11620), .A2(n8726), .ZN(n11700) );
  AND2_X1 U8057 ( .A1(n7599), .A2(n11703), .ZN(n7598) );
  NAND2_X1 U8058 ( .A1(n11629), .A2(n8726), .ZN(n7599) );
  NAND2_X1 U8059 ( .A1(n11621), .A2(n8725), .ZN(n11620) );
  AND2_X1 U8060 ( .A1(n8706), .A2(n8705), .ZN(n11621) );
  AND2_X1 U8061 ( .A1(n11513), .A2(n8959), .ZN(n7509) );
  OR2_X1 U8062 ( .A1(n15112), .A2(n8958), .ZN(n7510) );
  AND2_X1 U8063 ( .A1(n7510), .A2(n8959), .ZN(n11514) );
  OAI22_X1 U8064 ( .A1(n15118), .A2(n8691), .B1(n15119), .B2(n13904), .ZN(
        n11511) );
  NAND2_X1 U8065 ( .A1(n7139), .A2(n7138), .ZN(n15121) );
  NAND2_X1 U8066 ( .A1(n6868), .A2(n8661), .ZN(n11184) );
  NOR2_X1 U8067 ( .A1(n6962), .A2(n10981), .ZN(n6961) );
  INV_X1 U8068 ( .A(n8952), .ZN(n6962) );
  AND2_X1 U8069 ( .A1(n6821), .A2(n9283), .ZN(n7493) );
  NAND2_X1 U8070 ( .A1(n10543), .A2(n10562), .ZN(n10609) );
  NAND2_X1 U8071 ( .A1(n8942), .A2(n8508), .ZN(n10040) );
  AND2_X1 U8072 ( .A1(n9921), .A2(n9439), .ZN(n14027) );
  AND2_X1 U8073 ( .A1(n11264), .A2(n9019), .ZN(n10142) );
  NAND2_X1 U8074 ( .A1(n13969), .A2(n14176), .ZN(n7134) );
  AND2_X1 U8075 ( .A1(n13982), .A2(n13981), .ZN(n14184) );
  OR3_X1 U8076 ( .A1(n13980), .A2(n13979), .A3(n15125), .ZN(n13982) );
  NAND2_X1 U8077 ( .A1(n8794), .A2(n8793), .ZN(n14222) );
  AND2_X1 U8078 ( .A1(n9918), .A2(n8929), .ZN(n9964) );
  NOR2_X1 U8079 ( .A1(n14314), .A2(n8916), .ZN(n15340) );
  AND2_X1 U8080 ( .A1(n11722), .A2(n8915), .ZN(n8916) );
  MUX2_X1 U8081 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8924), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6929) );
  AND2_X1 U8082 ( .A1(n8651), .A2(n8665), .ZN(n10064) );
  AND2_X1 U8083 ( .A1(n8547), .A2(n8711), .ZN(n9490) );
  BUF_X1 U8084 ( .A(n8480), .Z(n8481) );
  AOI21_X1 U8085 ( .B1(n7355), .B2(n7357), .A(n6670), .ZN(n7353) );
  AND2_X1 U8086 ( .A1(n14323), .A2(n7331), .ZN(n7330) );
  NAND2_X1 U8087 ( .A1(n7332), .A2(n12672), .ZN(n7331) );
  INV_X1 U8088 ( .A(n14407), .ZN(n7332) );
  NAND2_X1 U8089 ( .A1(n12450), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7409) );
  NAND2_X1 U8090 ( .A1(n14377), .A2(n14379), .ZN(n14376) );
  OR2_X1 U8091 ( .A1(n11432), .A2(n11431), .ZN(n11647) );
  NOR2_X1 U8092 ( .A1(n12517), .A2(n7311), .ZN(n7310) );
  INV_X1 U8093 ( .A(n11951), .ZN(n7311) );
  CLKBUF_X1 U8094 ( .A(n14686), .Z(n6802) );
  INV_X1 U8095 ( .A(n7158), .ZN(n14703) );
  NAND2_X1 U8096 ( .A1(n14721), .A2(n11888), .ZN(n14698) );
  NAND2_X1 U8097 ( .A1(n6799), .A2(n7287), .ZN(n14746) );
  OAI21_X2 U8098 ( .B1(n11829), .B2(n7108), .A(n6639), .ZN(n14749) );
  INV_X1 U8099 ( .A(n7109), .ZN(n7108) );
  AND2_X1 U8100 ( .A1(n12511), .A2(n11856), .ZN(n7327) );
  NOR2_X1 U8101 ( .A1(n14763), .A2(n7106), .ZN(n7109) );
  NAND2_X1 U8102 ( .A1(n11829), .A2(n7111), .ZN(n7110) );
  OR2_X1 U8103 ( .A1(n14820), .A2(n14821), .ZN(n14818) );
  NOR2_X2 U8104 ( .A1(n14829), .A2(n14830), .ZN(n14827) );
  NOR2_X1 U8105 ( .A1(n11652), .A2(n7098), .ZN(n7095) );
  INV_X1 U8106 ( .A(n11446), .ZN(n7098) );
  AOI21_X1 U8107 ( .B1(n6616), .B2(n7279), .A(n6672), .ZN(n7275) );
  NAND2_X1 U8108 ( .A1(n11429), .A2(n7309), .ZN(n7277) );
  INV_X1 U8109 ( .A(n14464), .ZN(n11611) );
  NAND2_X1 U8110 ( .A1(n11156), .A2(n11155), .ZN(n11302) );
  NAND2_X1 U8111 ( .A1(n7314), .A2(n7313), .ZN(n11117) );
  NAND2_X1 U8112 ( .A1(n10743), .A2(n11058), .ZN(n11157) );
  NAND2_X1 U8113 ( .A1(n10576), .A2(n12498), .ZN(n10733) );
  INV_X1 U8114 ( .A(n14826), .ZN(n14850) );
  NAND2_X1 U8115 ( .A1(n9740), .A2(n9739), .ZN(n9788) );
  NAND2_X1 U8116 ( .A1(n12460), .A2(n12459), .ZN(n14591) );
  AND2_X1 U8117 ( .A1(n11871), .A2(n11870), .ZN(n14925) );
  AND2_X2 U8118 ( .A1(n10007), .A2(n10006), .ZN(n15236) );
  NAND2_X1 U8119 ( .A1(n9782), .A2(n10822), .ZN(n14966) );
  NOR2_X1 U8120 ( .A1(n8865), .A2(SI_27_), .ZN(n7589) );
  NAND2_X1 U8121 ( .A1(n8865), .A2(SI_27_), .ZN(n7588) );
  INV_X1 U8122 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9529) );
  NAND2_X1 U8123 ( .A1(n8817), .A2(n8815), .ZN(n7563) );
  XNOR2_X1 U8124 ( .A(n9327), .B(n9326), .ZN(n9820) );
  NAND2_X1 U8125 ( .A1(n7555), .A2(n8419), .ZN(n8663) );
  NAND2_X1 U8126 ( .A1(n8647), .A2(n8646), .ZN(n7555) );
  NAND2_X1 U8127 ( .A1(n8603), .A2(n8411), .ZN(n8618) );
  NAND2_X1 U8128 ( .A1(n8600), .A2(n8601), .ZN(n8603) );
  INV_X1 U8129 ( .A(n8401), .ZN(n8556) );
  NAND2_X1 U8130 ( .A1(n7100), .A2(n7101), .ZN(n8557) );
  AOI21_X1 U8131 ( .B1(n8541), .B2(n7103), .A(n7102), .ZN(n7101) );
  INV_X1 U8132 ( .A(n8396), .ZN(n7103) );
  NAND2_X1 U8133 ( .A1(n8557), .A2(n8556), .ZN(n8559) );
  XNOR2_X1 U8134 ( .A(n6838), .B(n7709), .ZN(n7711) );
  INV_X1 U8135 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7126) );
  NOR2_X1 U8136 ( .A1(n15044), .A2(n7726), .ZN(n7727) );
  OAI21_X1 U8137 ( .B1(n15175), .B2(n15174), .A(n7123), .ZN(n7122) );
  OR2_X1 U8138 ( .A1(n7692), .A2(n7691), .ZN(n7676) );
  INV_X1 U8139 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6835) );
  INV_X1 U8140 ( .A(n13703), .ZN(n12741) );
  INV_X1 U8141 ( .A(n10625), .ZN(n6742) );
  AOI21_X1 U8142 ( .B1(n7169), .B2(n12265), .A(n6720), .ZN(n7168) );
  OR2_X1 U8143 ( .A1(n6603), .A2(n9344), .ZN(n7900) );
  AND3_X1 U8144 ( .A1(n8137), .A2(n8136), .A3(n8135), .ZN(n13197) );
  NAND2_X1 U8145 ( .A1(n8113), .A2(n8112), .ZN(n13198) );
  NOR2_X1 U8146 ( .A1(n6626), .A2(n12872), .ZN(n7172) );
  NOR2_X1 U8147 ( .A1(n12279), .A2(n13151), .ZN(n7174) );
  AOI21_X1 U8148 ( .B1(n12279), .B2(n13186), .A(n12726), .ZN(n7175) );
  NAND2_X1 U8149 ( .A1(n8129), .A2(n8128), .ZN(n13187) );
  AND4_X1 U8150 ( .A1(n7943), .A2(n7942), .A3(n7941), .A4(n7940), .ZN(n15435)
         );
  INV_X1 U8151 ( .A(n12890), .ZN(n13263) );
  OR2_X1 U8152 ( .A1(n12735), .A2(n13152), .ZN(n6760) );
  NAND2_X1 U8153 ( .A1(n10620), .A2(n12235), .ZN(n12882) );
  OAI211_X1 U8154 ( .C1(n8162), .C2(n8161), .A(n8160), .B(n8159), .ZN(n13171)
         );
  INV_X1 U8155 ( .A(n13197), .ZN(n13170) );
  INV_X1 U8156 ( .A(n12901), .ZN(n7260) );
  NAND2_X1 U8157 ( .A1(n12901), .A2(n12932), .ZN(n12940) );
  XNOR2_X1 U8158 ( .A(n7195), .B(n12959), .ZN(n12950) );
  INV_X1 U8159 ( .A(n7195), .ZN(n12976) );
  NOR2_X1 U8160 ( .A1(n12950), .A2(n12962), .ZN(n12977) );
  INV_X1 U8161 ( .A(n7048), .ZN(n12996) );
  INV_X1 U8162 ( .A(n7046), .ZN(n13018) );
  OAI21_X1 U8163 ( .B1(n12950), .B2(n6898), .A(n6896), .ZN(n13002) );
  OR2_X1 U8164 ( .A1(n12979), .A2(n12962), .ZN(n6898) );
  NAND2_X1 U8165 ( .A1(n12978), .A2(n6897), .ZN(n6896) );
  INV_X1 U8166 ( .A(n12979), .ZN(n6897) );
  OR2_X1 U8167 ( .A1(n13004), .A2(n13003), .ZN(n6895) );
  NOR2_X1 U8168 ( .A1(n13050), .A2(n6841), .ZN(n6840) );
  NAND2_X1 U8169 ( .A1(n13048), .A2(n6737), .ZN(n6841) );
  NAND2_X1 U8170 ( .A1(n6891), .A2(n6890), .ZN(n13066) );
  NAND2_X1 U8171 ( .A1(n7203), .A2(n15425), .ZN(n6846) );
  XNOR2_X1 U8172 ( .A(n13068), .B(n13067), .ZN(n7203) );
  AND3_X1 U8173 ( .A1(n6890), .A2(n6891), .A3(n13065), .ZN(n13068) );
  NAND2_X1 U8174 ( .A1(n15421), .A2(n13073), .ZN(n7202) );
  INV_X1 U8175 ( .A(n13071), .ZN(n7201) );
  AOI21_X1 U8176 ( .B1(n7475), .B2(n7474), .A(n7473), .ZN(n7467) );
  NAND2_X1 U8177 ( .A1(n7080), .A2(n7077), .ZN(n13082) );
  NOR2_X1 U8178 ( .A1(n7079), .A2(n7078), .ZN(n7077) );
  NOR2_X1 U8179 ( .A1(n13111), .A2(n15492), .ZN(n7079) );
  INV_X1 U8180 ( .A(n13095), .ZN(n6824) );
  NAND2_X1 U8181 ( .A1(n6827), .A2(n6826), .ZN(n6825) );
  AOI21_X1 U8182 ( .B1(n11588), .B2(n12039), .A(n8154), .ZN(n13640) );
  OR2_X1 U8183 ( .A1(n13150), .A2(n13149), .ZN(n13638) );
  NAND2_X1 U8184 ( .A1(n8031), .A2(n8030), .ZN(n13676) );
  NAND2_X1 U8185 ( .A1(n7072), .A2(n12039), .ZN(n8031) );
  INV_X1 U8186 ( .A(n9887), .ZN(n7072) );
  NAND2_X1 U8187 ( .A1(n8084), .A2(n8083), .ZN(n13729) );
  INV_X1 U8188 ( .A(n7024), .ZN(n7023) );
  INV_X1 U8189 ( .A(n6800), .ZN(n8064) );
  OR3_X1 U8190 ( .A1(n11719), .A2(n11722), .A3(n14314), .ZN(n9934) );
  NAND2_X1 U8191 ( .A1(n7375), .A2(n6612), .ZN(n13814) );
  OR2_X1 U8192 ( .A1(n13849), .A2(n12591), .ZN(n7375) );
  NAND2_X1 U8193 ( .A1(n8719), .A2(n8718), .ZN(n14251) );
  NAND2_X1 U8194 ( .A1(n8781), .A2(n8780), .ZN(n14116) );
  NAND2_X1 U8195 ( .A1(n8635), .A2(n8634), .ZN(n11229) );
  NAND2_X1 U8196 ( .A1(n13849), .A2(n6612), .ZN(n7372) );
  AOI21_X1 U8197 ( .B1(n6612), .B2(n12591), .A(n6690), .ZN(n7376) );
  NAND2_X1 U8198 ( .A1(n9940), .A2(n14147), .ZN(n15107) );
  INV_X1 U8199 ( .A(n15104), .ZN(n13872) );
  NAND2_X1 U8200 ( .A1(n8877), .A2(n8876), .ZN(n13893) );
  OAI21_X1 U8201 ( .B1(n14035), .B2(n8887), .A(n8850), .ZN(n13894) );
  NAND2_X1 U8202 ( .A1(n6773), .A2(n6772), .ZN(n9430) );
  NAND2_X1 U8203 ( .A1(n9463), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6772) );
  OR2_X1 U8204 ( .A1(n9463), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6773) );
  INV_X1 U8205 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U8206 ( .A1(n11792), .A2(n15319), .ZN(n6770) );
  NOR2_X1 U8207 ( .A1(n11791), .A2(n6769), .ZN(n6768) );
  OR2_X1 U8208 ( .A1(n15300), .A2(n11795), .ZN(n6769) );
  INV_X1 U8209 ( .A(n9230), .ZN(n14264) );
  NAND2_X1 U8210 ( .A1(n8988), .A2(n8987), .ZN(n8989) );
  OR2_X1 U8211 ( .A1(n13974), .A2(n6956), .ZN(n13975) );
  INV_X1 U8212 ( .A(n8990), .ZN(n14163) );
  INV_X1 U8213 ( .A(n14264), .ZN(n6792) );
  OAI21_X1 U8214 ( .B1(n7619), .B2(n6621), .A(n9425), .ZN(n7142) );
  NOR2_X1 U8215 ( .A1(n9752), .A2(n7620), .ZN(n7619) );
  NAND2_X1 U8216 ( .A1(n9200), .A2(n9199), .ZN(n9230) );
  NAND2_X1 U8217 ( .A1(n7134), .A2(n15393), .ZN(n7133) );
  NAND2_X1 U8218 ( .A1(n7366), .A2(n7362), .ZN(n11739) );
  AOI21_X1 U8219 ( .B1(n7364), .B2(n7369), .A(n7363), .ZN(n7362) );
  NOR2_X1 U8220 ( .A1(n11734), .A2(n11735), .ZN(n7363) );
  NAND2_X1 U8221 ( .A1(n14397), .A2(n14396), .ZN(n14395) );
  NAND2_X1 U8222 ( .A1(n11141), .A2(n11140), .ZN(n12369) );
  OAI211_X1 U8223 ( .C1(n12526), .C2(n12524), .A(n6786), .B(n6785), .ZN(n6784)
         );
  AND2_X1 U8224 ( .A1(n6788), .A2(n6787), .ZN(n6786) );
  NAND2_X1 U8225 ( .A1(n12526), .A2(n12527), .ZN(n6785) );
  OR2_X1 U8226 ( .A1(n9830), .A2(n9819), .ZN(n12528) );
  OR2_X1 U8227 ( .A1(n9774), .A2(n14490), .ZN(n14824) );
  OR2_X1 U8228 ( .A1(n11449), .A2(n11448), .ZN(n11452) );
  NAND2_X1 U8229 ( .A1(n14979), .A2(n15264), .ZN(n6823) );
  CLKBUF_X1 U8230 ( .A(n15267), .Z(n15264) );
  OAI22_X1 U8231 ( .A1(n12458), .A2(n9362), .B1(n9751), .B2(n14504), .ZN(n9793) );
  INV_X1 U8232 ( .A(n14963), .ZN(n14900) );
  NAND2_X1 U8233 ( .A1(n14873), .A2(n7147), .ZN(n7146) );
  AND2_X1 U8234 ( .A1(n14872), .A2(n14871), .ZN(n7147) );
  NAND2_X1 U8235 ( .A1(n9714), .A2(n7361), .ZN(n9516) );
  XNOR2_X1 U8236 ( .A(n7711), .B(n7712), .ZN(n15619) );
  NOR2_X1 U8237 ( .A1(n15045), .A2(n15046), .ZN(n15044) );
  INV_X1 U8238 ( .A(n7731), .ZN(n7118) );
  OAI21_X1 U8239 ( .B1(n15185), .B2(n15186), .A(n7116), .ZN(n7115) );
  INV_X1 U8240 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7116) );
  NAND2_X1 U8241 ( .A1(n6759), .A2(n6758), .ZN(n7129) );
  INV_X1 U8242 ( .A(n15037), .ZN(n6758) );
  NAND2_X1 U8243 ( .A1(n7131), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7130) );
  NAND2_X1 U8244 ( .A1(n6815), .A2(n6814), .ZN(n12313) );
  NAND2_X1 U8245 ( .A1(n12339), .A2(n12312), .ZN(n6814) );
  NAND2_X1 U8246 ( .A1(n14475), .A2(n6588), .ZN(n6815) );
  NAND2_X1 U8247 ( .A1(n7523), .A2(n10143), .ZN(n9024) );
  INV_X1 U8248 ( .A(n12327), .ZN(n6817) );
  INV_X1 U8249 ( .A(n12342), .ZN(n7419) );
  INV_X1 U8250 ( .A(n12343), .ZN(n7418) );
  INV_X1 U8251 ( .A(n12350), .ZN(n7414) );
  NAND2_X1 U8252 ( .A1(n7540), .A2(n7539), .ZN(n7538) );
  INV_X1 U8253 ( .A(n9042), .ZN(n9043) );
  NAND2_X1 U8254 ( .A1(n9048), .A2(n9049), .ZN(n6905) );
  INV_X1 U8255 ( .A(n12352), .ZN(n7445) );
  NOR2_X1 U8256 ( .A1(n12355), .A2(n12352), .ZN(n7446) );
  NAND2_X1 U8257 ( .A1(n12068), .A2(n12183), .ZN(n7450) );
  OR2_X1 U8258 ( .A1(n9058), .A2(n9057), .ZN(n9064) );
  OAI21_X1 U8259 ( .B1(n12366), .B2(n7436), .A(n6683), .ZN(n12373) );
  NAND2_X1 U8260 ( .A1(n6615), .A2(n7531), .ZN(n6908) );
  NAND2_X1 U8261 ( .A1(n6910), .A2(n6913), .ZN(n9086) );
  OAI21_X1 U8262 ( .B1(n9077), .B2(n7530), .A(n6911), .ZN(n6910) );
  OAI21_X1 U8263 ( .B1(n12397), .B2(n7425), .A(n7428), .ZN(n7427) );
  INV_X1 U8264 ( .A(n9103), .ZN(n9106) );
  NAND2_X1 U8265 ( .A1(n7547), .A2(n9111), .ZN(n7546) );
  INV_X1 U8266 ( .A(n6691), .ZN(n7547) );
  AND2_X1 U8267 ( .A1(n9117), .A2(n9116), .ZN(n9119) );
  NAND2_X1 U8268 ( .A1(n6998), .A2(n7412), .ZN(n6997) );
  OR2_X1 U8269 ( .A1(n6998), .A2(n7412), .ZN(n6996) );
  INV_X1 U8270 ( .A(n9122), .ZN(n7517) );
  NOR2_X1 U8271 ( .A1(n9128), .A2(n9127), .ZN(n6920) );
  AND2_X1 U8272 ( .A1(n7535), .A2(n9136), .ZN(n7534) );
  OAI21_X1 U8273 ( .B1(n9129), .B2(n6921), .A(n6919), .ZN(n9141) );
  NAND2_X1 U8274 ( .A1(n7536), .A2(n6922), .ZN(n6921) );
  OAI21_X1 U8275 ( .B1(n7537), .B2(n6920), .A(n7536), .ZN(n6919) );
  INV_X1 U8276 ( .A(n6923), .ZN(n6922) );
  NAND2_X1 U8277 ( .A1(n6780), .A2(n6779), .ZN(n12436) );
  AND2_X1 U8278 ( .A1(n7440), .A2(n7439), .ZN(n6779) );
  AOI21_X1 U8279 ( .B1(n7442), .B2(n7440), .A(n7439), .ZN(n7438) );
  NAND2_X1 U8280 ( .A1(n6988), .A2(n12437), .ZN(n6987) );
  INV_X1 U8281 ( .A(n8437), .ZN(n7571) );
  INV_X1 U8282 ( .A(n8436), .ZN(n7568) );
  INV_X1 U8283 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7758) );
  INV_X1 U8284 ( .A(n7211), .ZN(n7210) );
  OAI21_X1 U8285 ( .B1(n8060), .B2(n7212), .A(n8093), .ZN(n7211) );
  INV_X1 U8286 ( .A(n8076), .ZN(n7212) );
  INV_X1 U8287 ( .A(n9152), .ZN(n7544) );
  NAND2_X1 U8288 ( .A1(n9224), .A2(n6669), .ZN(n7525) );
  NAND2_X1 U8289 ( .A1(n6640), .A2(n7528), .ZN(n7526) );
  AND2_X1 U8290 ( .A1(n9224), .A2(n6640), .ZN(n7524) );
  OAI22_X1 U8291 ( .A1(n12441), .A2(n7444), .B1(n12442), .B2(n7443), .ZN(
        n12445) );
  INV_X1 U8292 ( .A(n12440), .ZN(n7443) );
  NOR2_X1 U8293 ( .A1(n12440), .A2(n12443), .ZN(n7444) );
  OAI21_X1 U8294 ( .B1(n6986), .B2(n6681), .A(n6987), .ZN(n12441) );
  NOR2_X1 U8295 ( .A1(n14677), .A2(n7296), .ZN(n7295) );
  INV_X1 U8296 ( .A(n11975), .ZN(n7296) );
  NOR2_X1 U8297 ( .A1(n14807), .A2(n14786), .ZN(n7154) );
  NAND2_X1 U8298 ( .A1(n7589), .A2(n7588), .ZN(n7584) );
  NOR2_X1 U8299 ( .A1(n8879), .A2(n7587), .ZN(n7586) );
  INV_X1 U8300 ( .A(n7588), .ZN(n7587) );
  INV_X1 U8301 ( .A(n7565), .ZN(n7564) );
  OAI21_X1 U8302 ( .B1(n8815), .B2(n7566), .A(n8828), .ZN(n7565) );
  INV_X1 U8303 ( .A(n8449), .ZN(n7566) );
  INV_X1 U8304 ( .A(n8429), .ZN(n7576) );
  INV_X1 U8305 ( .A(n8692), .ZN(n7590) );
  INV_X1 U8306 ( .A(n7557), .ZN(n7556) );
  OAI21_X1 U8307 ( .B1(n8646), .B2(n7558), .A(n8662), .ZN(n7557) );
  INV_X1 U8308 ( .A(n8419), .ZN(n7558) );
  INV_X1 U8309 ( .A(n7092), .ZN(n6972) );
  NAND2_X1 U8310 ( .A1(n7125), .A2(n7648), .ZN(n7649) );
  NAND2_X1 U8311 ( .A1(n7705), .A2(n14509), .ZN(n7125) );
  MUX2_X1 U8312 ( .A(n12177), .B(n12176), .S(n12183), .Z(n12178) );
  NAND2_X1 U8313 ( .A1(n10300), .A2(n10299), .ZN(n10444) );
  NAND2_X1 U8314 ( .A1(n11093), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7052) );
  INV_X1 U8315 ( .A(n6712), .ZN(n7038) );
  AND2_X1 U8316 ( .A1(n7183), .A2(n6728), .ZN(n6888) );
  INV_X1 U8317 ( .A(n11756), .ZN(n7198) );
  NAND2_X1 U8318 ( .A1(n7197), .A2(n12910), .ZN(n12911) );
  AOI21_X1 U8319 ( .B1(n8287), .B2(n12151), .A(n7465), .ZN(n7464) );
  INV_X1 U8320 ( .A(n12156), .ZN(n7465) );
  INV_X1 U8321 ( .A(n12155), .ZN(n7463) );
  NAND2_X1 U8322 ( .A1(n8115), .A2(n8114), .ZN(n8132) );
  NOR2_X1 U8323 ( .A1(n7938), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7949) );
  AOI21_X1 U8324 ( .B1(n7012), .B2(n12103), .A(n7011), .ZN(n7010) );
  INV_X1 U8325 ( .A(n15439), .ZN(n7012) );
  INV_X1 U8326 ( .A(n12103), .ZN(n7013) );
  INV_X1 U8327 ( .A(n7063), .ZN(n7062) );
  INV_X1 U8328 ( .A(n8264), .ZN(n7064) );
  AOI21_X1 U8329 ( .B1(n7087), .B2(n7085), .A(n6684), .ZN(n7084) );
  NOR2_X1 U8330 ( .A1(n6637), .A2(n6614), .ZN(n7087) );
  INV_X1 U8331 ( .A(n10784), .ZN(n8331) );
  NAND2_X1 U8332 ( .A1(n9984), .A2(n9990), .ZN(n10182) );
  AND2_X1 U8333 ( .A1(n7756), .A2(n7089), .ZN(n7088) );
  INV_X1 U8334 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7089) );
  AND2_X1 U8335 ( .A1(n7167), .A2(n8246), .ZN(n6803) );
  INV_X1 U8336 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7757) );
  INV_X1 U8337 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7756) );
  AOI21_X1 U8338 ( .B1(n7254), .B2(n7252), .A(n6731), .ZN(n7251) );
  INV_X1 U8339 ( .A(n7254), .ZN(n7253) );
  INV_X1 U8340 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8246) );
  NAND2_X1 U8341 ( .A1(n7209), .A2(n7207), .ZN(n8096) );
  AOI21_X1 U8342 ( .B1(n7210), .B2(n7212), .A(n7208), .ZN(n7207) );
  NAND2_X1 U8343 ( .A1(n8061), .A2(n7210), .ZN(n7209) );
  INV_X1 U8344 ( .A(n8095), .ZN(n7208) );
  NAND2_X1 U8345 ( .A1(n8096), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8109) );
  NAND2_X1 U8346 ( .A1(n7843), .A2(n7636), .ZN(n7216) );
  INV_X1 U8347 ( .A(n7751), .ZN(n7804) );
  NAND2_X1 U8348 ( .A1(n9200), .A2(n7559), .ZN(n9263) );
  NOR2_X1 U8349 ( .A1(n13963), .A2(n7560), .ZN(n7559) );
  INV_X1 U8350 ( .A(n9199), .ZN(n7560) );
  OR2_X1 U8351 ( .A1(n8833), .A2(n13852), .ZN(n8845) );
  OR2_X1 U8352 ( .A1(n8845), .A2(n13821), .ZN(n8858) );
  INV_X1 U8353 ( .A(n8777), .ZN(n7615) );
  AND2_X1 U8354 ( .A1(n6613), .A2(n8960), .ZN(n6949) );
  AOI21_X1 U8355 ( .B1(n7497), .B2(n7495), .A(n6623), .ZN(n7494) );
  INV_X1 U8356 ( .A(n8947), .ZN(n7495) );
  INV_X1 U8357 ( .A(n7497), .ZN(n7496) );
  NOR2_X1 U8358 ( .A1(n8592), .A2(n8591), .ZN(n8610) );
  NAND2_X1 U8359 ( .A1(n7141), .A2(n7140), .ZN(n10608) );
  INV_X1 U8360 ( .A(n10609), .ZN(n7141) );
  AND2_X1 U8361 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8549) );
  OAI21_X1 U8362 ( .B1(n6964), .B2(n6963), .A(n7482), .ZN(n14069) );
  AOI21_X1 U8363 ( .B1(n7484), .B2(n7487), .A(n6675), .ZN(n7482) );
  INV_X1 U8364 ( .A(n7484), .ZN(n6963) );
  NAND2_X1 U8365 ( .A1(n10142), .A2(n10146), .ZN(n9931) );
  AND2_X1 U8366 ( .A1(n7612), .A2(n8465), .ZN(n7511) );
  INV_X1 U8367 ( .A(n8369), .ZN(n7612) );
  INV_X1 U8368 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8465) );
  INV_X1 U8369 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8462) );
  INV_X1 U8370 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8919) );
  NAND2_X1 U8371 ( .A1(n7395), .A2(n8912), .ZN(n7394) );
  INV_X1 U8372 ( .A(n7396), .ZN(n7395) );
  NOR2_X2 U8373 ( .A1(n6967), .A2(n6966), .ZN(n7551) );
  OR2_X1 U8374 ( .A1(n8587), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8604) );
  NOR2_X1 U8375 ( .A1(n7340), .A2(n7336), .ZN(n7335) );
  INV_X1 U8376 ( .A(n14379), .ZN(n7336) );
  INV_X1 U8377 ( .A(n14417), .ZN(n7340) );
  NAND2_X1 U8378 ( .A1(n14417), .A2(n7339), .ZN(n7338) );
  INV_X1 U8379 ( .A(n12665), .ZN(n10503) );
  NOR2_X1 U8380 ( .A1(n6659), .A2(n7421), .ZN(n7420) );
  AND2_X1 U8381 ( .A1(n7423), .A2(n7422), .ZN(n7421) );
  NOR2_X2 U8382 ( .A1(n14724), .A2(n14909), .ZN(n7158) );
  AND2_X1 U8383 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n11895), .ZN(n11906) );
  INV_X1 U8384 ( .A(n11867), .ZN(n7326) );
  NAND2_X1 U8385 ( .A1(n12510), .A2(n7105), .ZN(n7107) );
  NOR2_X1 U8386 ( .A1(n7106), .A2(n7111), .ZN(n7105) );
  OR2_X1 U8387 ( .A1(n11746), .A2(n11730), .ZN(n12387) );
  OR2_X1 U8388 ( .A1(n7309), .A2(n7279), .ZN(n7278) );
  INV_X1 U8389 ( .A(n11430), .ZN(n7279) );
  INV_X1 U8390 ( .A(n11136), .ZN(n7282) );
  OAI21_X1 U8391 ( .B1(n7283), .B2(n7282), .A(n12501), .ZN(n7281) );
  AND2_X1 U8392 ( .A1(n12500), .A2(n11105), .ZN(n7283) );
  INV_X1 U8393 ( .A(n10732), .ZN(n7315) );
  XNOR2_X1 U8394 ( .A(n12314), .B(n12315), .ZN(n12309) );
  INV_X1 U8395 ( .A(n7156), .ZN(n14668) );
  NAND2_X1 U8396 ( .A1(n7154), .A2(n7153), .ZN(n14767) );
  INV_X1 U8397 ( .A(n7154), .ZN(n14781) );
  NOR2_X2 U8398 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n10256) );
  AND2_X1 U8399 ( .A1(n7361), .A2(n7360), .ZN(n7359) );
  INV_X1 U8400 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7360) );
  INV_X1 U8401 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9326) );
  INV_X1 U8402 ( .A(n8399), .ZN(n7102) );
  NAND2_X1 U8403 ( .A1(n8393), .A2(SI_4_), .ZN(n8396) );
  AND2_X2 U8404 ( .A1(n6873), .A2(n6872), .ZN(n8387) );
  XNOR2_X1 U8405 ( .A(n7649), .B(n7124), .ZN(n7704) );
  OAI21_X1 U8406 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n7657), .A(n7656), .ZN(
        n7658) );
  OAI21_X1 U8407 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n7665), .A(n7664), .ZN(
        n7666) );
  NAND2_X1 U8408 ( .A1(n6805), .A2(n6804), .ZN(n10361) );
  NAND2_X1 U8409 ( .A1(n12068), .A2(n12734), .ZN(n6804) );
  INV_X1 U8410 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n13440) );
  NAND2_X1 U8411 ( .A1(n10790), .A2(n10791), .ZN(n10911) );
  NAND2_X1 U8412 ( .A1(n8086), .A2(n8085), .ZN(n8102) );
  AND2_X1 U8413 ( .A1(n12856), .A2(n12264), .ZN(n7169) );
  OR2_X1 U8414 ( .A1(n8069), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U8415 ( .A1(n8049), .A2(n13351), .ZN(n8069) );
  INV_X1 U8416 ( .A(n8050), .ZN(n8049) );
  NAND2_X1 U8417 ( .A1(n8015), .A2(n8014), .ZN(n8032) );
  INV_X1 U8418 ( .A(n12230), .ZN(n7459) );
  INV_X1 U8419 ( .A(n7470), .ZN(n7469) );
  OAI21_X1 U8420 ( .B1(n7475), .B2(n7473), .A(n12186), .ZN(n7470) );
  AND2_X1 U8421 ( .A1(n12190), .A2(n7625), .ZN(n12045) );
  OAI22_X1 U8422 ( .A1(n10238), .A2(n10239), .B1(n10231), .B2(n10230), .ZN(
        n15420) );
  INV_X1 U8423 ( .A(n7194), .ZN(n10214) );
  NAND2_X1 U8424 ( .A1(n6876), .A2(n6875), .ZN(n10300) );
  INV_X1 U8425 ( .A(n10215), .ZN(n6875) );
  INV_X1 U8426 ( .A(n10216), .ZN(n6876) );
  NOR2_X1 U8427 ( .A1(n11341), .A2(n11342), .ZN(n11340) );
  NOR2_X1 U8428 ( .A1(n11340), .A2(n11244), .ZN(n11362) );
  NAND2_X1 U8429 ( .A1(n6887), .A2(n11259), .ZN(n6886) );
  OR2_X1 U8430 ( .A1(n11237), .A2(n11236), .ZN(n7188) );
  NAND2_X1 U8431 ( .A1(n11356), .A2(n7186), .ZN(n7184) );
  AOI22_X1 U8432 ( .A1(n7036), .A2(n7038), .B1(n6625), .B2(n11378), .ZN(n7035)
         );
  NOR2_X1 U8433 ( .A1(n11375), .A2(n11376), .ZN(n11379) );
  INV_X1 U8434 ( .A(n6878), .ZN(n12923) );
  NAND2_X1 U8435 ( .A1(n12931), .A2(n6844), .ZN(n12935) );
  NAND2_X1 U8436 ( .A1(n6845), .A2(n7259), .ZN(n6844) );
  INV_X1 U8437 ( .A(n12933), .ZN(n6845) );
  NOR2_X1 U8438 ( .A1(n12984), .A2(n12961), .ZN(n12966) );
  AND2_X1 U8439 ( .A1(n12966), .A2(n12965), .ZN(n12983) );
  AND2_X1 U8440 ( .A1(n12955), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7196) );
  INV_X1 U8441 ( .A(n12995), .ZN(n7047) );
  NOR2_X1 U8442 ( .A1(n12983), .A2(n12984), .ZN(n12985) );
  NOR2_X1 U8443 ( .A1(n13042), .A2(n13041), .ZN(n13056) );
  AOI21_X1 U8444 ( .B1(n7476), .B2(n12180), .A(n12187), .ZN(n7475) );
  INV_X1 U8445 ( .A(n12180), .ZN(n7474) );
  INV_X1 U8446 ( .A(n12181), .ZN(n7473) );
  INV_X1 U8447 ( .A(n7475), .ZN(n7468) );
  NOR2_X1 U8448 ( .A1(n12047), .A2(n13074), .ZN(n7078) );
  AOI21_X1 U8449 ( .B1(n13092), .B2(n13093), .A(n15497), .ZN(n6826) );
  NAND2_X1 U8450 ( .A1(n13103), .A2(n12174), .ZN(n13127) );
  AND2_X1 U8451 ( .A1(n13147), .A2(n13148), .ZN(n13146) );
  NAND2_X1 U8452 ( .A1(n13181), .A2(n12159), .ZN(n8138) );
  AOI21_X1 U8453 ( .B1(n7464), .B2(n7466), .A(n7463), .ZN(n7462) );
  INV_X1 U8454 ( .A(n7464), .ZN(n6999) );
  INV_X1 U8455 ( .A(n12151), .ZN(n7466) );
  NAND2_X1 U8456 ( .A1(n8108), .A2(n13207), .ZN(n13206) );
  INV_X1 U8457 ( .A(n13204), .ZN(n8108) );
  AOI21_X1 U8458 ( .B1(n7003), .B2(n7005), .A(n12127), .ZN(n7001) );
  INV_X1 U8459 ( .A(n7004), .ZN(n7003) );
  INV_X1 U8460 ( .A(n12214), .ZN(n13254) );
  INV_X1 U8461 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n13347) );
  NAND2_X1 U8462 ( .A1(n7627), .A2(n8274), .ZN(n13578) );
  NAND2_X1 U8463 ( .A1(n15436), .A2(n8270), .ZN(n13569) );
  OR2_X1 U8464 ( .A1(n15438), .A2(n15439), .ZN(n15436) );
  OR2_X1 U8465 ( .A1(n7917), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U8466 ( .A1(n7028), .A2(n12039), .ZN(n7936) );
  INV_X1 U8467 ( .A(n9394), .ZN(n7028) );
  OR2_X1 U8468 ( .A1(n7819), .A2(n9377), .ZN(n7914) );
  AOI21_X1 U8469 ( .B1(n7017), .B2(n7019), .A(n7016), .ZN(n7015) );
  INV_X1 U8470 ( .A(n12095), .ZN(n7016) );
  NAND2_X1 U8471 ( .A1(n7903), .A2(n7902), .ZN(n7917) );
  INV_X1 U8472 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n7886) );
  AND2_X1 U8473 ( .A1(n7887), .A2(n7886), .ZN(n7903) );
  NOR2_X1 U8474 ( .A1(n7869), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7887) );
  NAND2_X1 U8475 ( .A1(n15463), .A2(n8264), .ZN(n11010) );
  OR2_X1 U8476 ( .A1(n7854), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7869) );
  NAND2_X1 U8477 ( .A1(n15462), .A2(n8263), .ZN(n15463) );
  AND2_X1 U8478 ( .A1(n15477), .A2(n15475), .ZN(n7059) );
  OR2_X1 U8479 ( .A1(n6603), .A2(n9381), .ZN(n7809) );
  INV_X1 U8480 ( .A(n12896), .ZN(n15495) );
  NAND2_X1 U8481 ( .A1(n8253), .A2(n9006), .ZN(n15502) );
  NAND2_X1 U8482 ( .A1(n10487), .A2(n10486), .ZN(n10489) );
  INV_X1 U8483 ( .A(n10357), .ZN(n15512) );
  NAND2_X1 U8484 ( .A1(n7968), .A2(n12112), .ZN(n13605) );
  NAND2_X1 U8485 ( .A1(n7071), .A2(n12039), .ZN(n7948) );
  INV_X1 U8486 ( .A(n9393), .ZN(n7071) );
  INV_X1 U8487 ( .A(n15569), .ZN(n15532) );
  OR2_X1 U8488 ( .A1(n9013), .A2(n8330), .ZN(n9987) );
  NAND2_X1 U8489 ( .A1(n7177), .A2(n11638), .ZN(n7178) );
  NAND2_X1 U8490 ( .A1(n12024), .A2(n12023), .ZN(n12038) );
  NAND2_X1 U8491 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), 
        .ZN(n7026) );
  OAI21_X1 U8492 ( .B1(n6632), .B2(n7026), .A(n7025), .ZN(n7024) );
  NAND2_X1 U8493 ( .A1(n7770), .A2(n7976), .ZN(n7025) );
  NAND2_X1 U8494 ( .A1(n8219), .A2(n8218), .ZN(n8232) );
  XNOR2_X1 U8495 ( .A(n7179), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U8496 ( .A1(n8312), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U8497 ( .A1(n8186), .A2(n8185), .ZN(n8189) );
  NAND2_X1 U8498 ( .A1(n8308), .A2(n7757), .ZN(n8312) );
  NOR2_X1 U8499 ( .A1(n8044), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U8500 ( .A1(n6800), .A2(n8065), .ZN(n8244) );
  INV_X1 U8501 ( .A(n7244), .ZN(n7243) );
  AOI21_X1 U8502 ( .B1(n7242), .B2(n7244), .A(n7241), .ZN(n7240) );
  INV_X1 U8503 ( .A(n8038), .ZN(n7241) );
  OR2_X1 U8504 ( .A1(n7995), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8028) );
  NAND2_X1 U8505 ( .A1(n6747), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6746) );
  INV_X1 U8506 ( .A(n7224), .ZN(n7223) );
  OR2_X1 U8507 ( .A1(n7875), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7893) );
  XNOR2_X1 U8508 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n7877) );
  XNOR2_X1 U8509 ( .A(n7840), .B(P3_IR_REG_4__SCAN_IN), .ZN(n10298) );
  NOR2_X1 U8510 ( .A1(n7623), .A2(n7205), .ZN(n7204) );
  XNOR2_X1 U8511 ( .A(n6940), .B(n10638), .ZN(n10387) );
  NAND2_X1 U8512 ( .A1(n9201), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7514) );
  NAND2_X1 U8513 ( .A1(n10639), .A2(n6940), .ZN(n10640) );
  NAND2_X1 U8514 ( .A1(n7381), .A2(n6939), .ZN(n10898) );
  AND2_X1 U8515 ( .A1(n10875), .A2(n10874), .ZN(n6939) );
  INV_X1 U8516 ( .A(n10878), .ZN(n10875) );
  NAND2_X1 U8517 ( .A1(n11319), .A2(n11320), .ZN(n11413) );
  NAND2_X1 U8518 ( .A1(n7399), .A2(n7397), .ZN(n11313) );
  NOR2_X1 U8519 ( .A1(n11222), .A2(n7398), .ZN(n7397) );
  INV_X1 U8520 ( .A(n11213), .ZN(n7398) );
  NAND2_X1 U8521 ( .A1(n10898), .A2(n7400), .ZN(n7399) );
  NOR2_X1 U8522 ( .A1(n11214), .A2(n7401), .ZN(n7400) );
  INV_X1 U8523 ( .A(n10897), .ZN(n7401) );
  INV_X1 U8524 ( .A(n10565), .ZN(n10382) );
  AND2_X1 U8525 ( .A1(n8549), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8563) );
  AND2_X1 U8526 ( .A1(n8563), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8577) );
  NOR2_X1 U8527 ( .A1(n8373), .A2(n11773), .ZN(n8484) );
  AOI21_X1 U8528 ( .B1(n9470), .B2(P2_REG2_REG_2__SCAN_IN), .A(n9469), .ZN(
        n15284) );
  AOI21_X1 U8529 ( .B1(n9484), .B2(P2_REG2_REG_3__SCAN_IN), .A(n15282), .ZN(
        n9598) );
  OAI21_X1 U8530 ( .B1(n9612), .B2(n9475), .A(n9474), .ZN(n9502) );
  AOI21_X1 U8531 ( .B1(n9586), .B2(P2_REG2_REG_7__SCAN_IN), .A(n9580), .ZN(
        n9583) );
  AOI21_X1 U8532 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n9861), .A(n9854), .ZN(
        n13922) );
  AOI21_X1 U8533 ( .B1(n10060), .B2(P2_REG2_REG_10__SCAN_IN), .A(n10059), .ZN(
        n13936) );
  NAND2_X1 U8534 ( .A1(n11781), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6848) );
  NAND2_X1 U8535 ( .A1(n6850), .A2(n6849), .ZN(n13956) );
  NAND2_X1 U8536 ( .A1(n11779), .A2(n13952), .ZN(n6849) );
  NOR2_X1 U8537 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13956), .ZN(n13955) );
  INV_X1 U8538 ( .A(n8995), .ZN(n13985) );
  NOR2_X1 U8539 ( .A1(n13979), .A2(n6656), .ZN(n6955) );
  INV_X1 U8540 ( .A(n9294), .ZN(n8977) );
  AOI21_X1 U8541 ( .B1(n7504), .B2(n7506), .A(n7503), .ZN(n7502) );
  INV_X1 U8542 ( .A(n9277), .ZN(n7503) );
  INV_X1 U8543 ( .A(n8782), .ZN(n8354) );
  AOI21_X1 U8544 ( .B1(n6945), .B2(n6947), .A(n6652), .ZN(n6942) );
  NAND2_X1 U8545 ( .A1(n6613), .A2(n6644), .ZN(n6948) );
  NAND2_X1 U8546 ( .A1(n11628), .A2(n6949), .ZN(n6944) );
  NAND2_X1 U8547 ( .A1(n11628), .A2(n8960), .ZN(n11704) );
  NAND2_X1 U8548 ( .A1(n8953), .A2(n8952), .ZN(n10982) );
  INV_X1 U8549 ( .A(n9285), .ZN(n10803) );
  INV_X1 U8550 ( .A(n9283), .ZN(n10770) );
  OAI21_X1 U8551 ( .B1(n10611), .B2(n7496), .A(n7494), .ZN(n10771) );
  NAND2_X1 U8552 ( .A1(n7499), .A2(n8948), .ZN(n10696) );
  NAND2_X1 U8553 ( .A1(n10611), .A2(n8947), .ZN(n7499) );
  NAND2_X1 U8554 ( .A1(n10606), .A2(n8582), .ZN(n10692) );
  NAND2_X1 U8555 ( .A1(n10541), .A2(n8569), .ZN(n10607) );
  NAND2_X1 U8556 ( .A1(n10607), .A2(n10610), .ZN(n10606) );
  NAND2_X1 U8557 ( .A1(n6951), .A2(n6950), .ZN(n10547) );
  AND2_X1 U8558 ( .A1(n6952), .A2(n9280), .ZN(n6950) );
  NAND2_X1 U8559 ( .A1(n10665), .A2(n6655), .ZN(n6951) );
  NAND2_X1 U8560 ( .A1(n10681), .A2(n10272), .ZN(n6952) );
  NOR2_X1 U8561 ( .A1(n6858), .A2(n9280), .ZN(n6774) );
  NOR2_X1 U8562 ( .A1(n7604), .A2(n7603), .ZN(n7602) );
  NAND2_X1 U8563 ( .A1(n10665), .A2(n8943), .ZN(n10678) );
  NAND2_X1 U8564 ( .A1(n10678), .A2(n10677), .ZN(n10676) );
  NAND2_X1 U8565 ( .A1(n10662), .A2(n8525), .ZN(n10682) );
  NAND2_X1 U8566 ( .A1(n9946), .A2(n8493), .ZN(n10036) );
  NAND2_X1 U8567 ( .A1(n8941), .A2(n6941), .ZN(n10043) );
  NAND2_X1 U8568 ( .A1(n10041), .A2(n10039), .ZN(n6941) );
  XNOR2_X1 U8569 ( .A(n9901), .B(n14166), .ZN(n9949) );
  NAND2_X1 U8570 ( .A1(n9950), .A2(n9949), .ZN(n10041) );
  XNOR2_X1 U8571 ( .A(n8938), .B(n9898), .ZN(n7403) );
  NAND2_X1 U8572 ( .A1(n8468), .A2(n8467), .ZN(n14179) );
  INV_X1 U8574 ( .A(n15386), .ZN(n14258) );
  INV_X1 U8575 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U8576 ( .A1(n7551), .A2(n7550), .ZN(n8910) );
  INV_X1 U8577 ( .A(n6807), .ZN(n8926) );
  OR2_X1 U8578 ( .A1(n8712), .A2(n8711), .ZN(n8714) );
  AND2_X1 U8579 ( .A1(n7368), .A2(n7369), .ZN(n7367) );
  INV_X1 U8580 ( .A(n11736), .ZN(n7368) );
  NOR2_X1 U8581 ( .A1(n11736), .A2(n7365), .ZN(n7364) );
  INV_X1 U8582 ( .A(n7370), .ZN(n7365) );
  INV_X1 U8583 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n13417) );
  NAND2_X1 U8584 ( .A1(n10760), .A2(n6660), .ZN(n11048) );
  OR2_X1 U8585 ( .A1(n11562), .A2(n11563), .ZN(n11561) );
  NOR2_X1 U8586 ( .A1(n11144), .A2(n11143), .ZN(n11287) );
  AND3_X1 U8587 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n10114) );
  INV_X1 U8588 ( .A(n9818), .ZN(n7344) );
  NOR2_X1 U8589 ( .A1(n11861), .A2(n14401), .ZN(n11872) );
  NAND2_X1 U8590 ( .A1(n6634), .A2(n7371), .ZN(n7370) );
  INV_X1 U8591 ( .A(n11479), .ZN(n7371) );
  NAND2_X1 U8592 ( .A1(n11561), .A2(n6634), .ZN(n7369) );
  INV_X1 U8593 ( .A(n11882), .ZN(n11883) );
  NAND2_X1 U8594 ( .A1(n14406), .A2(n14407), .ZN(n14405) );
  OR2_X1 U8595 ( .A1(n10736), .A2(n13417), .ZN(n11121) );
  OR2_X1 U8596 ( .A1(n11121), .A2(n11120), .ZN(n11144) );
  AND2_X1 U8597 ( .A1(n10114), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10412) );
  INV_X1 U8598 ( .A(n12525), .ZN(n6787) );
  INV_X1 U8599 ( .A(n11986), .ZN(n11878) );
  NAND2_X1 U8600 ( .A1(n12449), .A2(n12448), .ZN(n14870) );
  INV_X1 U8601 ( .A(n14887), .ZN(n7155) );
  AND2_X1 U8602 ( .A1(n14681), .A2(n11914), .ZN(n14667) );
  NAND2_X1 U8603 ( .A1(n14667), .A2(n14677), .ZN(n14666) );
  NAND2_X1 U8604 ( .A1(n7285), .A2(n6658), .ZN(n7284) );
  NOR2_X2 U8605 ( .A1(n14767), .A2(n14754), .ZN(n14753) );
  AOI21_X1 U8606 ( .B1(n7293), .B2(n14821), .A(n7291), .ZN(n7290) );
  INV_X1 U8607 ( .A(n12393), .ZN(n7291) );
  NOR2_X1 U8608 ( .A1(n11647), .A2(n11646), .ZN(n11823) );
  NAND2_X1 U8609 ( .A1(n11640), .A2(n7096), .ZN(n7099) );
  NOR2_X1 U8610 ( .A1(n11963), .A2(n7097), .ZN(n7096) );
  AOI21_X1 U8611 ( .B1(n11303), .B2(n7308), .A(n6671), .ZN(n7307) );
  INV_X1 U8612 ( .A(n11301), .ZN(n7308) );
  NAND2_X1 U8613 ( .A1(n11137), .A2(n11136), .ZN(n11294) );
  NAND2_X1 U8614 ( .A1(n11106), .A2(n11105), .ZN(n11111) );
  INV_X1 U8615 ( .A(n14824), .ZN(n14791) );
  NAND2_X1 U8616 ( .A1(n11106), .A2(n7283), .ZN(n11137) );
  INV_X1 U8617 ( .A(n10743), .ZN(n10744) );
  NOR2_X1 U8618 ( .A1(n10522), .A2(n14470), .ZN(n7289) );
  NAND2_X1 U8619 ( .A1(n10461), .A2(n10460), .ZN(n10462) );
  INV_X1 U8620 ( .A(n10474), .ZN(n10475) );
  NAND2_X1 U8621 ( .A1(n11059), .A2(n10401), .ZN(n10406) );
  NAND2_X1 U8622 ( .A1(n6789), .A2(n12341), .ZN(n10474) );
  INV_X1 U8623 ( .A(n11069), .ZN(n6789) );
  OAI21_X1 U8624 ( .B1(n10100), .B2(n11448), .A(n10102), .ZN(n12330) );
  AOI21_X1 U8626 ( .B1(n10322), .B2(n7303), .A(n6667), .ZN(n7302) );
  OR2_X1 U8627 ( .A1(n9774), .A2(n14494), .ZN(n14826) );
  OAI21_X1 U8628 ( .B1(n7273), .B2(n6622), .A(n9751), .ZN(n7272) );
  NAND2_X1 U8629 ( .A1(n12287), .A2(n12286), .ZN(n14583) );
  NAND2_X1 U8630 ( .A1(n14818), .A2(n7293), .ZN(n14803) );
  NAND2_X1 U8631 ( .A1(n14818), .A2(n11966), .ZN(n14801) );
  NAND2_X1 U8632 ( .A1(n11814), .A2(n12456), .ZN(n11817) );
  NAND2_X1 U8633 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), 
        .ZN(n7322) );
  XNOR2_X1 U8634 ( .A(n9234), .B(n9233), .ZN(n12457) );
  XNOR2_X1 U8635 ( .A(n9189), .B(n9188), .ZN(n12447) );
  NAND2_X1 U8636 ( .A1(n8446), .A2(n8445), .ZN(n8817) );
  NOR2_X1 U8637 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7361) );
  NAND2_X1 U8638 ( .A1(n9714), .A2(n9715), .ZN(n9518) );
  INV_X1 U8639 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U8640 ( .A1(n7577), .A2(n8429), .ZN(n8729) );
  OR2_X1 U8641 ( .A1(n10263), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n10494) );
  NAND2_X1 U8642 ( .A1(n7592), .A2(n8424), .ZN(n8693) );
  NAND2_X1 U8643 ( .A1(n7090), .A2(n6975), .ZN(n8631) );
  NAND2_X1 U8644 ( .A1(n7092), .A2(n8601), .ZN(n6975) );
  INV_X1 U8645 ( .A(n8410), .ZN(n8600) );
  NAND2_X1 U8646 ( .A1(n7104), .A2(n8396), .ZN(n8542) );
  NAND2_X1 U8647 ( .A1(n8395), .A2(n8527), .ZN(n7104) );
  CLKBUF_X1 U8648 ( .A(n9330), .Z(n9358) );
  NAND2_X1 U8649 ( .A1(n7645), .A2(n6754), .ZN(n7707) );
  NAND2_X1 U8650 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6755), .ZN(n6754) );
  INV_X1 U8651 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6755) );
  XNOR2_X1 U8652 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n7706) );
  XOR2_X1 U8653 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n7704), .Z(n7716) );
  OAI22_X1 U8654 ( .A1(n7675), .A2(P1_ADDR_REG_13__SCAN_IN), .B1(n7693), .B2(
        n7674), .ZN(n7691) );
  AOI21_X1 U8655 ( .B1(n13097), .B2(n6606), .A(n8229), .ZN(n13111) );
  AND4_X1 U8656 ( .A1(n7990), .A2(n7989), .A3(n7988), .A4(n7987), .ZN(n12830)
         );
  NAND2_X1 U8657 ( .A1(n11595), .A2(n11594), .ZN(n11597) );
  INV_X1 U8658 ( .A(n15483), .ZN(n10631) );
  AND2_X1 U8659 ( .A1(n8198), .A2(n8197), .ZN(n13110) );
  NAND2_X1 U8660 ( .A1(n10911), .A2(n10910), .ZN(n11032) );
  NAND2_X1 U8661 ( .A1(n12262), .A2(n12261), .ZN(n12814) );
  NAND2_X1 U8662 ( .A1(n11540), .A2(n11539), .ZN(n11542) );
  AND2_X1 U8663 ( .A1(n7170), .A2(n12264), .ZN(n12857) );
  NAND2_X1 U8664 ( .A1(n7170), .A2(n7169), .ZN(n12855) );
  NAND2_X1 U8665 ( .A1(n10910), .A2(n6611), .ZN(n7162) );
  NAND2_X1 U8666 ( .A1(n7163), .A2(n6611), .ZN(n7161) );
  INV_X1 U8667 ( .A(n12888), .ZN(n13123) );
  NAND2_X1 U8668 ( .A1(n7256), .A2(n8191), .ZN(n12870) );
  NAND2_X1 U8669 ( .A1(n11716), .A2(n12039), .ZN(n7256) );
  NAND2_X1 U8670 ( .A1(n9977), .A2(n10488), .ZN(n12885) );
  NAND2_X1 U8671 ( .A1(n10363), .A2(n15515), .ZN(n12880) );
  INV_X1 U8672 ( .A(n12052), .ZN(n7460) );
  NAND2_X1 U8673 ( .A1(n12231), .A2(n7459), .ZN(n7458) );
  NAND2_X1 U8674 ( .A1(n8184), .A2(n8183), .ZN(n13152) );
  INV_X1 U8675 ( .A(n12830), .ZN(n15065) );
  OR2_X1 U8676 ( .A1(n7868), .A2(n7813), .ZN(n7818) );
  OR2_X2 U8677 ( .A1(n9984), .A2(n13742), .ZN(n12897) );
  INV_X1 U8678 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n15415) );
  NAND2_X1 U8679 ( .A1(n7181), .A2(n10211), .ZN(n7182) );
  NAND2_X1 U8680 ( .A1(n7055), .A2(n7056), .ZN(n15427) );
  NOR2_X1 U8681 ( .A1(n10198), .A2(n10197), .ZN(n15425) );
  NAND2_X1 U8682 ( .A1(n7054), .A2(n7055), .ZN(n10208) );
  NAND2_X1 U8683 ( .A1(n7056), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7054) );
  AND2_X1 U8684 ( .A1(n10438), .A2(n10437), .ZN(n10440) );
  NOR2_X1 U8685 ( .A1(n11080), .A2(n11079), .ZN(n11233) );
  INV_X1 U8686 ( .A(n7043), .ZN(n11348) );
  INV_X1 U8687 ( .A(n7262), .ZN(n11346) );
  NAND2_X1 U8688 ( .A1(n7191), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7190) );
  NAND2_X1 U8689 ( .A1(n11234), .A2(n7191), .ZN(n7189) );
  INV_X1 U8690 ( .A(n11339), .ZN(n7191) );
  NAND2_X1 U8691 ( .A1(n7184), .A2(n7183), .ZN(n11663) );
  NOR2_X1 U8692 ( .A1(n11752), .A2(n11751), .ZN(n12900) );
  NAND2_X1 U8693 ( .A1(n11763), .A2(n6729), .ZN(n11766) );
  INV_X1 U8694 ( .A(n7263), .ZN(n12993) );
  AOI21_X1 U8695 ( .B1(n13750), .B2(n12039), .A(n12028), .ZN(n13079) );
  AND2_X1 U8696 ( .A1(n7068), .A2(n6650), .ZN(n13169) );
  NAND2_X1 U8697 ( .A1(n8292), .A2(n8291), .ZN(n13183) );
  AND2_X1 U8698 ( .A1(n13214), .A2(n13213), .ZN(n13657) );
  NAND2_X1 U8699 ( .A1(n7066), .A2(n8281), .ZN(n13232) );
  NAND2_X1 U8700 ( .A1(n8068), .A2(n8067), .ZN(n13242) );
  INV_X1 U8701 ( .A(n13667), .ZN(n8075) );
  NAND2_X1 U8702 ( .A1(n8048), .A2(n8047), .ZN(n13674) );
  NAND2_X1 U8703 ( .A1(n13556), .A2(n13558), .ZN(n7002) );
  NAND2_X1 U8704 ( .A1(n15434), .A2(n15439), .ZN(n7009) );
  NAND2_X1 U8705 ( .A1(n11017), .A2(n12090), .ZN(n15447) );
  NOR2_X1 U8706 ( .A1(n10489), .A2(n15527), .ZN(n15485) );
  AND2_X2 U8707 ( .A1(n10488), .A2(n15527), .ZN(n15508) );
  INV_X1 U8708 ( .A(n15504), .ZN(n15527) );
  NAND2_X1 U8709 ( .A1(n10489), .A2(n15525), .ZN(n15530) );
  NAND2_X1 U8710 ( .A1(n15485), .A2(n15523), .ZN(n13587) );
  NAND2_X1 U8711 ( .A1(n8237), .A2(n8236), .ZN(n8343) );
  NOR2_X1 U8712 ( .A1(n13082), .A2(n6648), .ZN(n9018) );
  INV_X1 U8713 ( .A(n13096), .ZN(n13699) );
  NOR2_X1 U8714 ( .A1(n13620), .A2(n6766), .ZN(n13696) );
  OR2_X1 U8715 ( .A1(n8205), .A2(n12612), .ZN(n8206) );
  NAND2_X1 U8716 ( .A1(n7073), .A2(n12039), .ZN(n8207) );
  INV_X1 U8717 ( .A(n12611), .ZN(n7073) );
  INV_X1 U8718 ( .A(n12870), .ZN(n13707) );
  OR2_X1 U8719 ( .A1(n13642), .A2(n13641), .ZN(n13712) );
  NAND2_X1 U8720 ( .A1(n10180), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13742) );
  AND2_X1 U8721 ( .A1(n8190), .A2(n8200), .ZN(n11716) );
  OR2_X1 U8722 ( .A1(n8189), .A2(n8188), .ZN(n8190) );
  INV_X1 U8723 ( .A(SI_26_), .ZN(n13511) );
  AND2_X1 U8724 ( .A1(n8186), .A2(n8172), .ZN(n11636) );
  OR2_X1 U8725 ( .A1(n8171), .A2(n8170), .ZN(n8172) );
  OAI21_X1 U8726 ( .B1(n8140), .B2(n8139), .A(n8141), .ZN(n8151) );
  AND2_X1 U8727 ( .A1(n7752), .A2(n7480), .ZN(n7479) );
  INV_X1 U8728 ( .A(SI_19_), .ZN(n10425) );
  NAND2_X1 U8729 ( .A1(n8077), .A2(n8076), .ZN(n8094) );
  INV_X1 U8730 ( .A(SI_16_), .ZN(n9886) );
  NAND2_X1 U8731 ( .A1(n7246), .A2(n7244), .ZN(n8039) );
  NAND2_X1 U8732 ( .A1(n7246), .A2(n7247), .ZN(n8026) );
  NAND2_X1 U8733 ( .A1(n8009), .A2(n8008), .ZN(n8023) );
  XNOR2_X1 U8734 ( .A(n8007), .B(n7993), .ZN(n9706) );
  INV_X1 U8735 ( .A(SI_13_), .ZN(n9578) );
  NAND2_X1 U8736 ( .A1(n7237), .A2(n7235), .ZN(n7970) );
  NAND2_X1 U8737 ( .A1(n7237), .A2(n7234), .ZN(n7961) );
  INV_X1 U8738 ( .A(SI_11_), .ZN(n13401) );
  NAND2_X1 U8739 ( .A1(n7220), .A2(n7224), .ZN(n7910) );
  NAND2_X1 U8740 ( .A1(n7879), .A2(n7226), .ZN(n7220) );
  NAND2_X1 U8741 ( .A1(n7230), .A2(n7226), .ZN(n7898) );
  NAND2_X1 U8742 ( .A1(n7230), .A2(n7228), .ZN(n7882) );
  INV_X1 U8743 ( .A(n10451), .ZN(n11093) );
  XNOR2_X1 U8744 ( .A(n7842), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10307) );
  NAND2_X1 U8745 ( .A1(n7219), .A2(n7217), .ZN(n7844) );
  NAND2_X1 U8746 ( .A1(n7219), .A2(n7822), .ZN(n7825) );
  NAND2_X1 U8747 ( .A1(n7794), .A2(n7793), .ZN(n7206) );
  NAND2_X1 U8748 ( .A1(n7058), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7057) );
  NAND2_X1 U8749 ( .A1(n7976), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7266) );
  NAND2_X1 U8750 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7772) );
  NAND2_X1 U8751 ( .A1(n10388), .A2(n10387), .ZN(n10641) );
  NAND2_X1 U8752 ( .A1(n7374), .A2(n13760), .ZN(n7373) );
  NAND2_X1 U8753 ( .A1(n13849), .A2(n6657), .ZN(n6930) );
  INV_X1 U8754 ( .A(n7376), .ZN(n7374) );
  NAND2_X1 U8755 ( .A1(n12542), .A2(n12541), .ZN(n15101) );
  AND2_X1 U8756 ( .A1(n12548), .A2(n12541), .ZN(n7405) );
  INV_X1 U8757 ( .A(n15100), .ZN(n12548) );
  NAND2_X1 U8758 ( .A1(n10898), .A2(n10897), .ZN(n11215) );
  INV_X1 U8759 ( .A(n7386), .ZN(n13780) );
  OAI21_X1 U8760 ( .B1(n13839), .B2(n7387), .A(n7393), .ZN(n7386) );
  INV_X1 U8761 ( .A(n7392), .ZN(n7387) );
  INV_X1 U8762 ( .A(n6938), .ZN(n7382) );
  NAND2_X1 U8763 ( .A1(n10641), .A2(n10640), .ZN(n10873) );
  NAND2_X1 U8764 ( .A1(n6934), .A2(n6936), .ZN(n6932) );
  OAI21_X1 U8765 ( .B1(n7384), .B2(n6936), .A(n6934), .ZN(n13809) );
  NAND2_X1 U8766 ( .A1(n7381), .A2(n10874), .ZN(n10877) );
  NAND2_X1 U8767 ( .A1(n8668), .A2(n8667), .ZN(n15148) );
  AND2_X1 U8768 ( .A1(n9939), .A2(n9923), .ZN(n15104) );
  AND2_X1 U8769 ( .A1(n15104), .A2(n13997), .ZN(n13875) );
  NAND2_X1 U8770 ( .A1(n7399), .A2(n11213), .ZN(n11223) );
  NAND2_X1 U8771 ( .A1(n9939), .A2(n9929), .ZN(n13853) );
  INV_X1 U8772 ( .A(n9903), .ZN(n9904) );
  NOR2_X1 U8773 ( .A1(n13839), .A2(n12559), .ZN(n13866) );
  OR2_X1 U8774 ( .A1(n9299), .A2(n8937), .ZN(n9300) );
  NAND2_X1 U8775 ( .A1(n8864), .A2(n8863), .ZN(n14028) );
  AND2_X1 U8776 ( .A1(n6856), .A2(n6854), .ZN(n6744) );
  INV_X1 U8777 ( .A(n14003), .ZN(n6854) );
  NAND2_X1 U8778 ( .A1(n6855), .A2(n6856), .ZN(n14004) );
  NAND2_X1 U8779 ( .A1(n14022), .A2(n8974), .ZN(n14016) );
  OAI21_X1 U8780 ( .B1(n14049), .B2(n7608), .A(n7605), .ZN(n14007) );
  NAND2_X1 U8781 ( .A1(n14051), .A2(n8840), .ZN(n14021) );
  AND2_X1 U8782 ( .A1(n14079), .A2(n8814), .ZN(n14062) );
  NAND2_X1 U8783 ( .A1(n6857), .A2(n8803), .ZN(n14077) );
  NAND2_X1 U8784 ( .A1(n7483), .A2(n7488), .ZN(n14081) );
  NAND2_X1 U8785 ( .A1(n14109), .A2(n8966), .ZN(n14096) );
  NAND2_X1 U8786 ( .A1(n7616), .A2(n8777), .ZN(n14108) );
  INV_X1 U8787 ( .A(n14233), .ZN(n8992) );
  NAND2_X1 U8788 ( .A1(n14144), .A2(n8750), .ZN(n14124) );
  OAI21_X1 U8789 ( .B1(n8706), .B2(n7597), .A(n6862), .ZN(n14141) );
  OAI21_X1 U8790 ( .B1(n11621), .B2(n7600), .A(n7598), .ZN(n11702) );
  NAND2_X1 U8791 ( .A1(n7510), .A2(n7509), .ZN(n11512) );
  NAND2_X1 U8792 ( .A1(n6960), .A2(n8954), .ZN(n15126) );
  NAND2_X1 U8793 ( .A1(n8653), .A2(n8652), .ZN(n15135) );
  OR2_X1 U8794 ( .A1(n8990), .A2(n8998), .ZN(n15334) );
  INV_X1 U8795 ( .A(n15334), .ZN(n15132) );
  NOR2_X1 U8796 ( .A1(n15331), .A2(n10148), .ZN(n14168) );
  INV_X1 U8797 ( .A(n7134), .ZN(n7132) );
  NAND2_X1 U8798 ( .A1(n8609), .A2(n8608), .ZN(n10890) );
  OR2_X1 U8799 ( .A1(n10726), .A2(n8478), .ZN(n8609) );
  NAND2_X1 U8800 ( .A1(n8548), .A2(n6869), .ZN(n10372) );
  OR2_X1 U8801 ( .A1(n10100), .A2(n8478), .ZN(n6869) );
  INV_X1 U8802 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6866) );
  AND2_X1 U8803 ( .A1(n9934), .A2(n9308), .ZN(n15352) );
  INV_X1 U8804 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n14300) );
  INV_X1 U8805 ( .A(n8373), .ZN(n12001) );
  INV_X1 U8806 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11721) );
  XNOR2_X1 U8807 ( .A(n8914), .B(n8913), .ZN(n11719) );
  INV_X1 U8808 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10529) );
  INV_X1 U8809 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9673) );
  INV_X1 U8810 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9418) );
  INV_X1 U8811 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9412) );
  INV_X1 U8812 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9392) );
  INV_X1 U8813 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9387) );
  INV_X1 U8814 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9365) );
  INV_X1 U8815 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9364) );
  INV_X1 U8816 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9367) );
  INV_X1 U8817 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9368) );
  NAND2_X1 U8818 ( .A1(n8483), .A2(n8482), .ZN(n9463) );
  MUX2_X1 U8819 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8479), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8483) );
  INV_X1 U8820 ( .A(n14316), .ZN(n6810) );
  NAND2_X1 U8821 ( .A1(n14405), .A2(n12672), .ZN(n14322) );
  NAND2_X1 U8822 ( .A1(n11110), .A2(n11109), .ZN(n15249) );
  NAND2_X1 U8823 ( .A1(n10003), .A2(n10004), .ZN(n14330) );
  NAND2_X1 U8824 ( .A1(n12714), .A2(n7351), .ZN(n7350) );
  INV_X1 U8825 ( .A(n7355), .ZN(n7351) );
  NAND2_X1 U8826 ( .A1(n7353), .A2(n12714), .ZN(n7352) );
  NAND2_X1 U8827 ( .A1(n10760), .A2(n10759), .ZN(n10763) );
  NAND2_X1 U8828 ( .A1(n14395), .A2(n12656), .ZN(n14349) );
  AOI21_X1 U8829 ( .B1(n7330), .B2(n7333), .A(n6668), .ZN(n7328) );
  INV_X1 U8830 ( .A(n12672), .ZN(n7333) );
  NAND2_X1 U8831 ( .A1(n12649), .A2(n6809), .ZN(n6808) );
  INV_X1 U8832 ( .A(n12650), .ZN(n6809) );
  OAI21_X1 U8833 ( .B1(n6839), .B2(n7370), .A(n7369), .ZN(n11737) );
  NAND2_X1 U8834 ( .A1(n15033), .A2(n9751), .ZN(n14917) );
  NOR2_X1 U8835 ( .A1(n6839), .A2(n11479), .ZN(n11564) );
  CLKBUF_X1 U8836 ( .A(n11478), .Z(n6839) );
  NAND2_X1 U8837 ( .A1(n14416), .A2(n14417), .ZN(n14415) );
  NAND2_X1 U8838 ( .A1(n14376), .A2(n14378), .ZN(n14416) );
  INV_X1 U8839 ( .A(n14456), .ZN(n14425) );
  INV_X1 U8840 ( .A(n10331), .ZN(n14474) );
  INV_X1 U8841 ( .A(n14870), .ZN(n14611) );
  NAND2_X1 U8842 ( .A1(n6802), .A2(n11975), .ZN(n14678) );
  NAND2_X1 U8843 ( .A1(n14700), .A2(n11901), .ZN(n14683) );
  NAND2_X1 U8844 ( .A1(n14749), .A2(n11867), .ZN(n14735) );
  NAND2_X1 U8845 ( .A1(n14746), .A2(n11970), .ZN(n14733) );
  NAND2_X1 U8846 ( .A1(n11857), .A2(n11856), .ZN(n14751) );
  NAND2_X1 U8847 ( .A1(n7110), .A2(n7109), .ZN(n11857) );
  NAND2_X1 U8848 ( .A1(n7110), .A2(n11841), .ZN(n14764) );
  NAND2_X1 U8849 ( .A1(n11829), .A2(n11828), .ZN(n14777) );
  NAND2_X1 U8850 ( .A1(n11640), .A2(n11639), .ZN(n11812) );
  NAND2_X1 U8851 ( .A1(n7277), .A2(n11430), .ZN(n11467) );
  NAND2_X1 U8852 ( .A1(n11426), .A2(n11425), .ZN(n12380) );
  NAND2_X1 U8853 ( .A1(n14840), .A2(n10823), .ZN(n14831) );
  NAND2_X1 U8854 ( .A1(n11304), .A2(n11303), .ZN(n11422) );
  NAND2_X1 U8855 ( .A1(n11302), .A2(n11301), .ZN(n11304) );
  NAND2_X1 U8856 ( .A1(n10734), .A2(n12499), .ZN(n11115) );
  NAND2_X1 U8857 ( .A1(n10733), .A2(n10732), .ZN(n10734) );
  NAND2_X1 U8858 ( .A1(n10314), .A2(n10322), .ZN(n10400) );
  NAND2_X1 U8859 ( .A1(n10841), .A2(n10313), .ZN(n10314) );
  OR2_X1 U8860 ( .A1(n9830), .A2(n9829), .ZN(n14852) );
  INV_X1 U8861 ( .A(n14838), .ZN(n14857) );
  AND2_X1 U8862 ( .A1(n14840), .A2(n14939), .ZN(n14856) );
  NAND2_X1 U8863 ( .A1(n11297), .A2(n12456), .ZN(n7114) );
  NAND2_X1 U8864 ( .A1(n10728), .A2(n10727), .ZN(n12356) );
  INV_X1 U8865 ( .A(n14583), .ZN(n14973) );
  INV_X1 U8866 ( .A(n14591), .ZN(n14977) );
  INV_X1 U8867 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7300) );
  OR3_X1 U8868 ( .A1(n14914), .A2(n14913), .A3(n14912), .ZN(n14993) );
  INV_X1 U8869 ( .A(n14830), .ZN(n15012) );
  INV_X2 U8870 ( .A(n15257), .ZN(n15259) );
  AND2_X1 U8871 ( .A1(n9320), .A2(n9321), .ZN(n9400) );
  NAND2_X1 U8872 ( .A1(n6831), .A2(n6829), .ZN(n9320) );
  NAND2_X1 U8873 ( .A1(n6830), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6829) );
  OAI21_X1 U8874 ( .B1(n9319), .B2(n9318), .A(P1_IR_REG_24__SCAN_IN), .ZN(
        n6831) );
  INV_X1 U8875 ( .A(n9396), .ZN(n9403) );
  INV_X1 U8876 ( .A(n7323), .ZN(n7629) );
  NAND2_X1 U8877 ( .A1(n9746), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U8878 ( .A1(n7581), .A2(n7588), .ZN(n8880) );
  INV_X1 U8879 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n13373) );
  INV_X1 U8880 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10496) );
  NAND2_X1 U8881 ( .A1(n8424), .A2(n7591), .ZN(n8678) );
  INV_X1 U8882 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n13505) );
  INV_X1 U8883 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9451) );
  INV_X1 U8884 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9424) );
  NAND2_X1 U8885 ( .A1(n8603), .A2(n8602), .ZN(n10726) );
  OR2_X1 U8886 ( .A1(n8601), .A2(n8600), .ZN(n8602) );
  INV_X1 U8887 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9391) );
  INV_X1 U8888 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U8889 ( .A1(n8559), .A2(n6931), .ZN(n8571) );
  NOR2_X1 U8890 ( .A1(n8570), .A2(n6981), .ZN(n6931) );
  NAND2_X1 U8891 ( .A1(n6871), .A2(n6870), .ZN(n10100) );
  NAND2_X1 U8892 ( .A1(n8542), .A2(n8541), .ZN(n6870) );
  NAND2_X1 U8893 ( .A1(n7148), .A2(n8398), .ZN(n6871) );
  INV_X1 U8894 ( .A(n8542), .ZN(n7148) );
  INV_X1 U8895 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9340) );
  INV_X1 U8896 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9351) );
  INV_X1 U8897 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9355) );
  INV_X1 U8898 ( .A(n8498), .ZN(n8500) );
  NOR2_X1 U8899 ( .A1(n7713), .A2(n15618), .ZN(n15041) );
  AOI21_X1 U8900 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n7715), .A(n15614), .ZN(
        n15606) );
  XNOR2_X1 U8901 ( .A(n7117), .B(n7720), .ZN(n15609) );
  NAND2_X1 U8902 ( .A1(n15609), .A2(n15608), .ZN(n15607) );
  XNOR2_X1 U8903 ( .A(n7725), .B(n7724), .ZN(n15045) );
  NAND2_X1 U8904 ( .A1(n15611), .A2(n7730), .ZN(n15049) );
  OAI21_X1 U8905 ( .B1(n15056), .B2(n15055), .A(n6833), .ZN(n6832) );
  INV_X1 U8906 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n6833) );
  INV_X1 U8907 ( .A(n7734), .ZN(n7121) );
  AOI21_X1 U8908 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n7738), .A(n15188), .ZN(
        n15193) );
  NOR2_X1 U8909 ( .A1(n7741), .A2(n7740), .ZN(n15059) );
  NAND2_X1 U8910 ( .A1(n6627), .A2(n12874), .ZN(n7173) );
  NAND2_X1 U8911 ( .A1(n7044), .A2(n12940), .ZN(n12902) );
  NOR2_X1 U8912 ( .A1(n12977), .A2(n12978), .ZN(n12980) );
  AND2_X1 U8913 ( .A1(n13047), .A2(n6840), .ZN(n13051) );
  AND2_X1 U8914 ( .A1(n7202), .A2(n7201), .ZN(n7200) );
  NAND2_X1 U8915 ( .A1(n11800), .A2(n9913), .ZN(n9927) );
  NAND2_X1 U8916 ( .A1(n7372), .A2(n7376), .ZN(n13761) );
  NAND2_X1 U8917 ( .A1(n6771), .A2(n6767), .ZN(n11797) );
  NAND2_X1 U8918 ( .A1(n6770), .A2(n6768), .ZN(n6767) );
  NAND2_X1 U8919 ( .A1(n11796), .A2(n11795), .ZN(n6771) );
  AOI21_X1 U8920 ( .B1(n14178), .B2(n6581), .A(n9002), .ZN(n9003) );
  AOI21_X1 U8921 ( .B1(n6792), .B2(n14248), .A(n6791), .ZN(n6790) );
  NOR2_X1 U8922 ( .A1(n15404), .A2(n14175), .ZN(n6791) );
  AND2_X1 U8923 ( .A1(n14270), .A2(n14248), .ZN(n6743) );
  AOI21_X1 U8924 ( .B1(n9230), .B2(n14294), .A(n6796), .ZN(n6795) );
  NOR2_X1 U8925 ( .A1(n15393), .A2(n14263), .ZN(n6796) );
  OAI21_X1 U8926 ( .B1(n7136), .B2(n7133), .A(n7137), .ZN(n14265) );
  NAND2_X1 U8927 ( .A1(n15391), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U8928 ( .A1(n6867), .A2(n6864), .ZN(P2_U3495) );
  AOI21_X1 U8929 ( .B1(n14270), .B2(n14294), .A(n6865), .ZN(n6864) );
  NAND2_X1 U8930 ( .A1(n14269), .A2(n15393), .ZN(n6867) );
  NOR2_X1 U8931 ( .A1(n15393), .A2(n6866), .ZN(n6865) );
  INV_X1 U8932 ( .A(n6784), .ZN(n12532) );
  NAND2_X1 U8933 ( .A1(n15265), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7143) );
  OR2_X1 U8934 ( .A1(n15264), .A2(n11952), .ZN(n6822) );
  NAND2_X1 U8935 ( .A1(n7301), .A2(n7298), .ZN(P1_U3524) );
  AOI21_X1 U8936 ( .B1(n14980), .B2(n14988), .A(n7299), .ZN(n7298) );
  NAND2_X1 U8937 ( .A1(n14979), .A2(n15259), .ZN(n7301) );
  NOR2_X1 U8938 ( .A1(n15259), .A2(n7300), .ZN(n7299) );
  INV_X1 U8939 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n6836) );
  AND2_X1 U8940 ( .A1(n6777), .A2(n7129), .ZN(n6837) );
  NAND2_X1 U8941 ( .A1(n15036), .A2(n15037), .ZN(n6777) );
  XNOR2_X1 U8942 ( .A(n7128), .B(n7127), .ZN(SUB_1596_U4) );
  XNOR2_X1 U8943 ( .A(n7746), .B(n6741), .ZN(n7127) );
  NAND2_X1 U8944 ( .A1(n7129), .A2(n7130), .ZN(n7128) );
  AND2_X1 U8945 ( .A1(n7608), .A2(n6617), .ZN(n6610) );
  OR2_X1 U8946 ( .A1(n11030), .A2(n15459), .ZN(n6611) );
  AND2_X1 U8947 ( .A1(n7377), .A2(n13816), .ZN(n6612) );
  OR2_X1 U8948 ( .A1(n14293), .A2(n13834), .ZN(n6613) );
  INV_X1 U8949 ( .A(n8298), .ZN(n10221) );
  XNOR2_X1 U8950 ( .A(n12375), .B(n7113), .ZN(n11303) );
  INV_X1 U8951 ( .A(n11303), .ZN(n7309) );
  INV_X1 U8952 ( .A(n12514), .ZN(n7297) );
  NAND2_X1 U8953 ( .A1(n13568), .A2(n8273), .ZN(n6614) );
  AND2_X1 U8954 ( .A1(n6913), .A2(n6909), .ZN(n6615) );
  CLKBUF_X3 U8955 ( .A(n7523), .Z(n9208) );
  AND2_X1 U8956 ( .A1(n11466), .A2(n7278), .ZN(n6616) );
  NAND2_X1 U8957 ( .A1(n14196), .A2(n14028), .ZN(n6617) );
  XOR2_X1 U8958 ( .A(n13729), .B(n13212), .Z(n6618) );
  INV_X1 U8959 ( .A(n9111), .ZN(n7549) );
  AND2_X1 U8960 ( .A1(n13598), .A2(n12112), .ZN(n6619) );
  AND2_X1 U8961 ( .A1(n7424), .A2(n7429), .ZN(n6620) );
  AND2_X1 U8962 ( .A1(n7620), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6621) );
  AND2_X1 U8963 ( .A1(n7274), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6622) );
  AND2_X1 U8964 ( .A1(n7500), .A2(n13909), .ZN(n6623) );
  AND2_X1 U8965 ( .A1(n12499), .A2(n7315), .ZN(n6624) );
  INV_X1 U8966 ( .A(n11764), .ZN(n7041) );
  AND2_X1 U8967 ( .A1(n6712), .A2(n7041), .ZN(n6625) );
  OAI211_X1 U8968 ( .C1(n7868), .C2(n8148), .A(n8147), .B(n8146), .ZN(n13151)
         );
  XOR2_X1 U8969 ( .A(n6711), .B(n7174), .Z(n6626) );
  XOR2_X1 U8970 ( .A(n6711), .B(n7175), .Z(n6627) );
  AND2_X1 U8971 ( .A1(n6889), .A2(n11374), .ZN(n6628) );
  INV_X1 U8972 ( .A(n15119), .ZN(n7138) );
  CLKBUF_X3 U8973 ( .A(n10503), .Z(n10103) );
  OR2_X1 U8974 ( .A1(n14008), .A2(n14189), .ZN(n6629) );
  NOR2_X1 U8975 ( .A1(n9751), .A2(n14484), .ZN(n6630) );
  OR2_X2 U8976 ( .A1(n11708), .A2(n14293), .ZN(n6631) );
  INV_X1 U8977 ( .A(n14465), .ZN(n7113) );
  INV_X1 U8978 ( .A(n6606), .ZN(n8238) );
  INV_X1 U8979 ( .A(n12208), .ZN(n7011) );
  NAND2_X1 U8980 ( .A1(n8491), .A2(n8490), .ZN(n9026) );
  AND2_X1 U8981 ( .A1(n7481), .A2(n7759), .ZN(n6632) );
  NAND2_X1 U8982 ( .A1(n12117), .A2(n12118), .ZN(n8272) );
  XNOR2_X1 U8983 ( .A(n14765), .B(n14792), .ZN(n14763) );
  OR2_X1 U8984 ( .A1(n14651), .A2(n14878), .ZN(n6633) );
  XNOR2_X1 U8985 ( .A(n8370), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8372) );
  INV_X1 U8986 ( .A(n8372), .ZN(n11773) );
  INV_X1 U8987 ( .A(n12714), .ZN(n7358) );
  NAND2_X1 U8988 ( .A1(n11609), .A2(n11608), .ZN(n6634) );
  AND2_X1 U8989 ( .A1(n9079), .A2(n9078), .ZN(n6635) );
  AND2_X1 U8990 ( .A1(n9163), .A2(n9162), .ZN(n6636) );
  AND2_X1 U8991 ( .A1(n15439), .A2(n8270), .ZN(n6637) );
  NAND2_X1 U8992 ( .A1(n7931), .A2(n7932), .ZN(n7946) );
  AND2_X1 U8993 ( .A1(n8871), .A2(n10686), .ZN(n6638) );
  AND2_X1 U8994 ( .A1(n11860), .A2(n11859), .ZN(n14999) );
  INV_X1 U8995 ( .A(n7608), .ZN(n7607) );
  AND2_X1 U8996 ( .A1(n7107), .A2(n7327), .ZN(n6639) );
  AND3_X1 U8997 ( .A1(n7751), .A2(n7750), .A3(n7167), .ZN(n7925) );
  NAND2_X1 U8998 ( .A1(n13206), .A2(n12151), .ZN(n13193) );
  XNOR2_X1 U8999 ( .A(n7876), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11251) );
  AND2_X1 U9000 ( .A1(n7641), .A2(n7527), .ZN(n6640) );
  OR2_X1 U9001 ( .A1(n11251), .A2(n11250), .ZN(n6641) );
  AND2_X1 U9002 ( .A1(n8295), .A2(n12181), .ZN(n13093) );
  AND2_X1 U9003 ( .A1(n12499), .A2(n12498), .ZN(n6642) );
  OR2_X1 U9004 ( .A1(n12992), .A2(n12991), .ZN(n6643) );
  AND2_X1 U9005 ( .A1(n14293), .A2(n13834), .ZN(n6644) );
  INV_X1 U9006 ( .A(n13977), .ZN(n6956) );
  AND3_X1 U9007 ( .A1(n7751), .A2(n7750), .A3(n7166), .ZN(n6645) );
  AND2_X1 U9008 ( .A1(n15460), .A2(n11176), .ZN(n6646) );
  INV_X1 U9009 ( .A(n7258), .ZN(n10224) );
  XNOR2_X1 U9010 ( .A(n7805), .B(P3_IR_REG_3__SCAN_IN), .ZN(n7258) );
  INV_X1 U9011 ( .A(n6964), .ZN(n14109) );
  AND2_X1 U9012 ( .A1(n14031), .A2(n13894), .ZN(n6647) );
  AND2_X1 U9013 ( .A1(n13087), .A2(n15569), .ZN(n6648) );
  AND2_X1 U9014 ( .A1(n7605), .A2(n6617), .ZN(n6649) );
  OR2_X1 U9015 ( .A1(n13187), .A2(n13170), .ZN(n6650) );
  INV_X1 U9016 ( .A(n12372), .ZN(n7433) );
  AND2_X1 U9017 ( .A1(n7287), .A2(n14734), .ZN(n6651) );
  AND2_X1 U9018 ( .A1(n14237), .A2(n13842), .ZN(n6652) );
  AND2_X1 U9019 ( .A1(n7034), .A2(n7036), .ZN(n6653) );
  INV_X1 U9020 ( .A(n9291), .ZN(n14048) );
  XNOR2_X1 U9021 ( .A(n14205), .B(n13822), .ZN(n9291) );
  NOR2_X1 U9022 ( .A1(n14222), .A2(n14114), .ZN(n6654) );
  XNOR2_X1 U9023 ( .A(n10687), .B(n12011), .ZN(n10681) );
  AND2_X1 U9024 ( .A1(n8943), .A2(n10272), .ZN(n6655) );
  AND2_X1 U9025 ( .A1(n13988), .A2(n13892), .ZN(n6656) );
  INV_X1 U9026 ( .A(n7575), .ZN(n7574) );
  NOR2_X1 U9027 ( .A1(n8430), .A2(n7576), .ZN(n7575) );
  AND2_X1 U9028 ( .A1(n6612), .A2(n13760), .ZN(n6657) );
  INV_X1 U9029 ( .A(n12432), .ZN(n7441) );
  INV_X1 U9030 ( .A(n12438), .ZN(n6988) );
  NAND2_X1 U9031 ( .A1(n14925), .A2(n14459), .ZN(n6658) );
  NOR2_X1 U9032 ( .A1(n12471), .A2(n12472), .ZN(n6659) );
  AND2_X1 U9033 ( .A1(n10761), .A2(n10759), .ZN(n6660) );
  AND2_X1 U9034 ( .A1(n9258), .A2(n7525), .ZN(n6661) );
  AND2_X1 U9035 ( .A1(n8598), .A2(n8582), .ZN(n6662) );
  AND2_X1 U9036 ( .A1(n8813), .A2(n8803), .ZN(n6663) );
  AND2_X1 U9037 ( .A1(n6928), .A2(n9063), .ZN(n6664) );
  OR2_X1 U9038 ( .A1(n8760), .A2(n7396), .ZN(n6665) );
  AND2_X1 U9039 ( .A1(n6618), .A2(n12139), .ZN(n6666) );
  AND2_X1 U9040 ( .A1(n12139), .A2(n12142), .ZN(n13233) );
  AND2_X1 U9041 ( .A1(n12325), .A2(n12326), .ZN(n6667) );
  AND2_X1 U9042 ( .A1(n12678), .A2(n12677), .ZN(n6668) );
  INV_X1 U9043 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9744) );
  INV_X1 U9044 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U9045 ( .A1(n7628), .A2(n7526), .ZN(n6669) );
  AND2_X1 U9046 ( .A1(n12707), .A2(n12706), .ZN(n6670) );
  NAND2_X1 U9047 ( .A1(n12911), .A2(n12932), .ZN(n12922) );
  NOR2_X1 U9048 ( .A1(n11842), .A2(n7112), .ZN(n7111) );
  NOR2_X1 U9049 ( .A1(n12375), .A2(n14465), .ZN(n6671) );
  NOR2_X1 U9050 ( .A1(n12380), .A2(n11611), .ZN(n6672) );
  NOR2_X1 U9051 ( .A1(n14257), .A2(n15099), .ZN(n6673) );
  NOR2_X1 U9052 ( .A1(n14196), .A2(n14028), .ZN(n6674) );
  NOR2_X1 U9053 ( .A1(n14087), .A2(n12570), .ZN(n6675) );
  INV_X1 U9054 ( .A(n7531), .ZN(n7530) );
  NAND2_X1 U9055 ( .A1(n7532), .A2(n9076), .ZN(n7531) );
  AND2_X1 U9056 ( .A1(n14707), .A2(n11973), .ZN(n6676) );
  AND2_X1 U9057 ( .A1(n6799), .A2(n11968), .ZN(n6677) );
  INV_X1 U9058 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9342) );
  AND2_X1 U9059 ( .A1(n14116), .A2(n13898), .ZN(n6678) );
  AND2_X1 U9060 ( .A1(n13187), .A2(n13170), .ZN(n6679) );
  AND2_X1 U9061 ( .A1(n8727), .A2(SI_17_), .ZN(n6680) );
  AND2_X1 U9062 ( .A1(n12434), .A2(n12433), .ZN(n6681) );
  AND2_X1 U9063 ( .A1(n9047), .A2(n7644), .ZN(n6682) );
  AND2_X1 U9064 ( .A1(n7435), .A2(n7433), .ZN(n6683) );
  NOR2_X1 U9065 ( .A1(n8277), .A2(n8276), .ZN(n6684) );
  INV_X1 U9066 ( .A(n8726), .ZN(n7600) );
  NAND2_X1 U9067 ( .A1(n7925), .A2(n7477), .ZN(n6685) );
  INV_X1 U9068 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8461) );
  OR2_X1 U9069 ( .A1(n12416), .A2(n12415), .ZN(n6686) );
  AND2_X1 U9070 ( .A1(n8416), .A2(n13401), .ZN(n6687) );
  AND2_X1 U9071 ( .A1(n8421), .A2(n9578), .ZN(n6688) );
  AND2_X1 U9072 ( .A1(n9392), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n6689) );
  INV_X1 U9073 ( .A(n10910), .ZN(n7164) );
  NAND2_X1 U9074 ( .A1(n12596), .A2(n12593), .ZN(n6690) );
  AND2_X1 U9075 ( .A1(n9110), .A2(n9109), .ZN(n6691) );
  OAI21_X1 U9076 ( .B1(n10791), .B2(n7164), .A(n11031), .ZN(n7163) );
  NAND2_X1 U9077 ( .A1(n7431), .A2(n12398), .ZN(n6692) );
  INV_X1 U9078 ( .A(n8272), .ZN(n13598) );
  INV_X1 U9079 ( .A(n12435), .ZN(n7439) );
  INV_X1 U9080 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9357) );
  INV_X1 U9081 ( .A(n12470), .ZN(n7422) );
  AND2_X1 U9082 ( .A1(n7572), .A2(n7571), .ZN(n6693) );
  XNOR2_X1 U9083 ( .A(n14786), .B(n14802), .ZN(n14788) );
  OAI21_X1 U9084 ( .B1(n9208), .B2(n12011), .A(n9050), .ZN(n9051) );
  INV_X1 U9085 ( .A(n9051), .ZN(n7522) );
  OR2_X1 U9086 ( .A1(n15193), .A2(n15194), .ZN(n6694) );
  NOR2_X1 U9087 ( .A1(n12356), .A2(n14468), .ZN(n6695) );
  OR2_X1 U9088 ( .A1(n8760), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n6696) );
  AND2_X1 U9089 ( .A1(n10206), .A2(n7258), .ZN(n6697) );
  NAND2_X1 U9090 ( .A1(n7925), .A2(n7479), .ZN(n6698) );
  AND2_X1 U9091 ( .A1(n6632), .A2(n7770), .ZN(n7022) );
  OR2_X1 U9092 ( .A1(n13969), .A2(n13970), .ZN(n6699) );
  AND2_X1 U9093 ( .A1(n7297), .A2(n11973), .ZN(n6700) );
  AND2_X1 U9094 ( .A1(n7176), .A2(n11594), .ZN(n6701) );
  OR2_X1 U9095 ( .A1(n12437), .A2(n6988), .ZN(n6702) );
  NAND2_X1 U9096 ( .A1(n10093), .A2(n10092), .ZN(n6703) );
  AND2_X1 U9097 ( .A1(n6895), .A2(n6894), .ZN(n6704) );
  AND2_X1 U9098 ( .A1(n7358), .A2(n7355), .ZN(n6705) );
  AND2_X1 U9099 ( .A1(n7088), .A2(n7481), .ZN(n6706) );
  AND2_X1 U9100 ( .A1(n14598), .A2(n11961), .ZN(n12517) );
  AND2_X1 U9101 ( .A1(n6846), .A2(n6750), .ZN(n6707) );
  INV_X1 U9102 ( .A(n12419), .ZN(n6998) );
  INV_X1 U9103 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7058) );
  OR2_X1 U9104 ( .A1(n7423), .A2(n7422), .ZN(n6708) );
  INV_X1 U9105 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6830) );
  AND3_X1 U9106 ( .A1(n8461), .A2(n8462), .A3(n8463), .ZN(n6709) );
  AND2_X1 U9107 ( .A1(n9093), .A2(n9092), .ZN(n6710) );
  XOR2_X1 U9108 ( .A(n12730), .B(n13171), .Z(n6711) );
  NAND2_X1 U9109 ( .A1(n11644), .A2(n11643), .ZN(n14967) );
  INV_X1 U9110 ( .A(n14967), .ZN(n7152) );
  NAND2_X1 U9111 ( .A1(n11905), .A2(n11904), .ZN(n14691) );
  INV_X1 U9112 ( .A(n14691), .ZN(n7157) );
  NAND2_X1 U9113 ( .A1(n11670), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U9114 ( .A1(n7750), .A2(n7751), .ZN(n7895) );
  INV_X1 U9115 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U9116 ( .A1(n7002), .A2(n12130), .ZN(n13257) );
  INV_X1 U9117 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7166) );
  AND2_X1 U9118 ( .A1(n6944), .A2(n6948), .ZN(n6713) );
  AND2_X1 U9119 ( .A1(n7384), .A2(n6937), .ZN(n6714) );
  INV_X1 U9120 ( .A(n11378), .ZN(n7039) );
  AND2_X1 U9121 ( .A1(n9095), .A2(n9094), .ZN(n6715) );
  AND2_X1 U9122 ( .A1(n9131), .A2(n9130), .ZN(n6716) );
  AND2_X1 U9123 ( .A1(n13667), .A2(n12139), .ZN(n6717) );
  AND2_X1 U9124 ( .A1(n11447), .A2(n11446), .ZN(n6718) );
  AND2_X1 U9125 ( .A1(n12658), .A2(n12656), .ZN(n6719) );
  AND2_X1 U9126 ( .A1(n12267), .A2(n13247), .ZN(n6720) );
  OR2_X1 U9127 ( .A1(n9152), .A2(n9154), .ZN(n6721) );
  AND2_X1 U9128 ( .A1(n9115), .A2(n9114), .ZN(n6722) );
  INV_X1 U9129 ( .A(n7393), .ZN(n7391) );
  OR2_X1 U9130 ( .A1(n11564), .A2(n11561), .ZN(n6723) );
  INV_X1 U9131 ( .A(n6889), .ZN(n6887) );
  NAND2_X1 U9132 ( .A1(n11254), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6889) );
  INV_X1 U9133 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10265) );
  OR2_X1 U9134 ( .A1(n12570), .A2(n10037), .ZN(n6724) );
  INV_X1 U9135 ( .A(n7037), .ZN(n7036) );
  OAI21_X1 U9136 ( .B1(n7039), .B2(n7038), .A(n11764), .ZN(n7037) );
  OR2_X1 U9137 ( .A1(n9148), .A2(n9147), .ZN(n6725) );
  OR2_X1 U9138 ( .A1(n7544), .A2(n9153), .ZN(n6726) );
  AND2_X1 U9139 ( .A1(n6721), .A2(n6917), .ZN(n6727) );
  NAND2_X1 U9140 ( .A1(n11670), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6728) );
  INV_X1 U9141 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9713) );
  AND2_X2 U9142 ( .A1(n9964), .A2(n9963), .ZN(n15404) );
  INV_X1 U9143 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7248) );
  AND2_X1 U9144 ( .A1(n8936), .A2(n14147), .ZN(n8990) );
  INV_X1 U9145 ( .A(n12932), .ZN(n7259) );
  NAND2_X1 U9146 ( .A1(n11847), .A2(n11846), .ZN(n14765) );
  INV_X1 U9147 ( .A(n14765), .ZN(n7153) );
  INV_X1 U9148 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n7050) );
  OR2_X1 U9149 ( .A1(n11765), .A2(n11764), .ZN(n6729) );
  OAI21_X1 U9150 ( .B1(n10980), .B2(n8644), .A(n8645), .ZN(n15133) );
  NAND2_X1 U9151 ( .A1(n7009), .A2(n12103), .ZN(n11582) );
  OR2_X1 U9152 ( .A1(n12567), .A2(n12566), .ZN(n6730) );
  INV_X1 U9153 ( .A(n14378), .ZN(n7339) );
  NAND2_X1 U9154 ( .A1(n12018), .A2(n10377), .ZN(n10563) );
  NAND2_X1 U9155 ( .A1(n7925), .A2(n7752), .ZN(n8044) );
  INV_X1 U9156 ( .A(n7151), .ZN(n11462) );
  NOR2_X2 U9157 ( .A1(n11440), .A2(n12380), .ZN(n7151) );
  AND2_X1 U9158 ( .A1(n11578), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6731) );
  OR2_X1 U9159 ( .A1(n8760), .A2(n8369), .ZN(n6732) );
  AND2_X1 U9160 ( .A1(n8451), .A2(SI_24_), .ZN(n6733) );
  INV_X1 U9161 ( .A(n7139), .ZN(n15120) );
  NOR2_X2 U9162 ( .A1(n15137), .A2(n15148), .ZN(n7139) );
  AND2_X1 U9163 ( .A1(n7188), .A2(n7187), .ZN(n6734) );
  AND2_X1 U9164 ( .A1(n7040), .A2(n7039), .ZN(n6735) );
  OR2_X1 U9165 ( .A1(n13011), .A2(n12994), .ZN(n6736) );
  INV_X1 U9166 ( .A(n15267), .ZN(n15265) );
  INV_X1 U9167 ( .A(n12872), .ZN(n12874) );
  INV_X1 U9168 ( .A(n13020), .ZN(n7265) );
  NAND2_X1 U9169 ( .A1(n7403), .A2(n11795), .ZN(n9899) );
  INV_X1 U9170 ( .A(n10704), .ZN(n7500) );
  NAND2_X1 U9171 ( .A1(n9905), .A2(n9904), .ZN(n10131) );
  INV_X1 U9172 ( .A(SI_27_), .ZN(n12612) );
  AND2_X2 U9173 ( .A1(n9964), .A2(n9958), .ZN(n15393) );
  INV_X1 U9174 ( .A(n14230), .ZN(n14248) );
  INV_X1 U9175 ( .A(n15326), .ZN(n7140) );
  AND2_X1 U9176 ( .A1(n8296), .A2(n12052), .ZN(n15497) );
  INV_X1 U9177 ( .A(n15497), .ZN(n15513) );
  NAND2_X1 U9178 ( .A1(n9909), .A2(n11802), .ZN(n11800) );
  OR2_X1 U9179 ( .A1(n15414), .A2(n13049), .ZN(n6737) );
  NOR2_X1 U9180 ( .A1(n11233), .A2(n11234), .ZN(n6738) );
  INV_X1 U9181 ( .A(n6874), .ZN(n10445) );
  NAND2_X1 U9182 ( .A1(n10301), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n6874) );
  AND2_X1 U9183 ( .A1(n9899), .A2(n10605), .ZN(n14261) );
  AND2_X1 U9184 ( .A1(n11274), .A2(n6848), .ZN(n6739) );
  XNOR2_X1 U9185 ( .A(n8080), .B(n8079), .ZN(n13060) );
  INV_X1 U9186 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7123) );
  AND2_X1 U9187 ( .A1(n12231), .A2(n7460), .ZN(n6740) );
  INV_X1 U9188 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7971) );
  XOR2_X1 U9189 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n6741) );
  INV_X1 U9190 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7124) );
  AOI21_X1 U9191 ( .B1(n6954), .B2(n6580), .A(n8989), .ZN(n14181) );
  INV_X1 U9192 ( .A(n6580), .ZN(n15125) );
  NAND2_X1 U9193 ( .A1(n9838), .A2(n9816), .ZN(n9817) );
  NAND2_X1 U9194 ( .A1(n9839), .A2(n9840), .ZN(n9838) );
  XNOR2_X1 U9195 ( .A(n9197), .B(n9196), .ZN(n14298) );
  NAND2_X1 U9196 ( .A1(n7585), .A2(n7582), .ZN(n9189) );
  NAND2_X1 U9197 ( .A1(n9192), .A2(n9191), .ZN(n9234) );
  OAI21_X2 U9198 ( .B1(n12829), .B2(n12248), .A(n12250), .ZN(n12746) );
  NAND2_X1 U9199 ( .A1(n10361), .A2(n10358), .ZN(n10531) );
  NAND3_X1 U9200 ( .A1(n10627), .A2(n6742), .A3(n10626), .ZN(n10789) );
  OAI21_X2 U9201 ( .B1(n10790), .B2(n7162), .A(n7161), .ZN(n11034) );
  INV_X1 U9202 ( .A(n11542), .ZN(n6757) );
  NAND2_X1 U9203 ( .A1(n8338), .A2(n7756), .ZN(n8306) );
  AOI21_X2 U9204 ( .B1(n12733), .B2(n12732), .A(n12731), .ZN(n12799) );
  INV_X1 U9205 ( .A(n6820), .ZN(n6819) );
  OR2_X1 U9206 ( .A1(n14186), .A2(n6743), .ZN(P2_U3527) );
  NAND2_X1 U9207 ( .A1(n7609), .A2(n8851), .ZN(n7608) );
  NAND2_X1 U9208 ( .A1(n7563), .A2(n8449), .ZN(n8830) );
  NAND2_X1 U9209 ( .A1(n10320), .A2(n12493), .ZN(n11063) );
  NAND2_X1 U9210 ( .A1(n11065), .A2(n10409), .ZN(n10457) );
  NAND2_X1 U9211 ( .A1(n10334), .A2(n10318), .ZN(n10843) );
  NAND2_X1 U9212 ( .A1(n14707), .A2(n6700), .ZN(n14686) );
  NAND2_X1 U9213 ( .A1(n11978), .A2(n11977), .ZN(n14654) );
  NOR2_X2 U9214 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9330) );
  OAI21_X1 U9215 ( .B1(n11106), .B2(n7282), .A(n7280), .ZN(n11296) );
  AOI21_X1 U9216 ( .B1(n11969), .B2(n6651), .A(n7284), .ZN(n14719) );
  AOI21_X1 U9217 ( .B1(n14787), .B2(n14788), .A(n11967), .ZN(n14761) );
  NAND3_X1 U9218 ( .A1(n7270), .A2(n7269), .A3(n9529), .ZN(n9741) );
  AOI21_X1 U9219 ( .B1(n14875), .B2(n14939), .A(n7146), .ZN(n7145) );
  NAND2_X1 U9220 ( .A1(n14709), .A2(n14708), .ZN(n14707) );
  NAND2_X1 U9221 ( .A1(n14761), .A2(n14763), .ZN(n11969) );
  NAND2_X1 U9222 ( .A1(n7292), .A2(n7290), .ZN(n14787) );
  NAND2_X1 U9223 ( .A1(n14978), .A2(n15267), .ZN(n7144) );
  NAND2_X1 U9224 ( .A1(n11193), .A2(n7643), .ZN(n11473) );
  NAND2_X1 U9225 ( .A1(n10099), .A2(n10098), .ZN(n10499) );
  NAND2_X1 U9226 ( .A1(n13195), .A2(n8290), .ZN(n8292) );
  NAND2_X1 U9227 ( .A1(n6745), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7992) );
  INV_X1 U9228 ( .A(n13578), .ZN(n6748) );
  NAND2_X1 U9229 ( .A1(n13155), .A2(n13154), .ZN(n13153) );
  NAND2_X1 U9230 ( .A1(n13230), .A2(n8283), .ZN(n13220) );
  AOI21_X1 U9231 ( .B1(n7929), .B2(n7639), .A(n7632), .ZN(n7931) );
  NAND2_X1 U9232 ( .A1(n7864), .A2(n7863), .ZN(n7879) );
  NAND2_X1 U9233 ( .A1(n6746), .A2(n7991), .ZN(n7973) );
  NAND2_X1 U9234 ( .A1(n7912), .A2(n7911), .ZN(n7928) );
  NOR2_X1 U9235 ( .A1(n13091), .A2(n7083), .ZN(n7082) );
  INV_X1 U9236 ( .A(n7973), .ZN(n6745) );
  INV_X1 U9237 ( .A(n7972), .ZN(n6747) );
  OR2_X1 U9238 ( .A1(n9848), .A2(n9847), .ZN(n9850) );
  NAND2_X1 U9239 ( .A1(n7998), .A2(n7997), .ZN(n12752) );
  NOR2_X1 U9240 ( .A1(n13092), .A2(n13093), .ZN(n13091) );
  XNOR2_X1 U9241 ( .A(n7082), .B(n12221), .ZN(n7081) );
  NAND2_X1 U9242 ( .A1(n7081), .A2(n15513), .ZN(n7080) );
  NAND2_X1 U9243 ( .A1(n6751), .A2(n15429), .ZN(n6750) );
  XNOR2_X1 U9244 ( .A(n13055), .B(n13062), .ZN(n6751) );
  INV_X1 U9245 ( .A(n11252), .ZN(n6752) );
  NAND2_X1 U9246 ( .A1(n14115), .A2(n14105), .ZN(n14099) );
  INV_X1 U9247 ( .A(n10437), .ZN(n7051) );
  NAND2_X1 U9248 ( .A1(n7032), .A2(n7031), .ZN(n11662) );
  OAI21_X1 U9249 ( .B1(n11379), .B2(n7037), .A(n7035), .ZN(n7033) );
  OAI211_X1 U9250 ( .C1(n13072), .C2(n15406), .A(n7200), .B(n6707), .ZN(
        P3_U3201) );
  NOR2_X1 U9251 ( .A1(n12951), .A2(n7264), .ZN(n12991) );
  NAND3_X1 U9252 ( .A1(n7551), .A2(n8462), .A3(n7550), .ZN(n8908) );
  NAND2_X1 U9253 ( .A1(n11060), .A2(n11062), .ZN(n11059) );
  NOR2_X2 U9254 ( .A1(n14596), .A2(n7312), .ZN(n14597) );
  NAND2_X1 U9255 ( .A1(n8473), .A2(n8384), .ZN(n8498) );
  XNOR2_X1 U9256 ( .A(n8529), .B(n8528), .ZN(n10011) );
  NAND2_X1 U9257 ( .A1(n7144), .A2(n7143), .ZN(P1_U3557) );
  NAND2_X1 U9258 ( .A1(n7329), .A2(n7328), .ZN(n14388) );
  NAND2_X1 U9259 ( .A1(n7354), .A2(n12701), .ZN(n6811) );
  NAND2_X1 U9260 ( .A1(n15179), .A2(n15178), .ZN(n15177) );
  INV_X1 U9261 ( .A(n15036), .ZN(n6759) );
  AOI21_X1 U9262 ( .B1(n6694), .B2(n6835), .A(n6834), .ZN(n7741) );
  XNOR2_X1 U9263 ( .A(n6837), .B(n6836), .ZN(SUB_1596_U62) );
  XNOR2_X1 U9264 ( .A(n10787), .B(n12896), .ZN(n10625) );
  NAND2_X1 U9265 ( .A1(n10359), .A2(n6605), .ZN(n6805) );
  NAND2_X1 U9266 ( .A1(n9319), .A2(n6830), .ZN(n9321) );
  NAND2_X1 U9267 ( .A1(n10531), .A2(n10530), .ZN(n10622) );
  OAI21_X2 U9268 ( .B1(n12799), .B2(n12800), .A(n6760), .ZN(n12862) );
  AOI21_X2 U9269 ( .B1(n14446), .B2(n14445), .A(n6761), .ZN(n14368) );
  NOR2_X1 U9270 ( .A1(n12622), .A2(n6762), .ZN(n6761) );
  INV_X1 U9271 ( .A(n12623), .ZN(n6762) );
  XNOR2_X1 U9272 ( .A(n6811), .B(n6810), .ZN(n14321) );
  XNOR2_X2 U9273 ( .A(n12307), .B(n14844), .ZN(n12490) );
  AND4_X4 U9274 ( .A1(n7410), .A2(n9749), .A3(n7411), .A4(n7409), .ZN(n12307)
         );
  NAND2_X1 U9275 ( .A1(n10406), .A2(n10410), .ZN(n10461) );
  NAND2_X1 U9276 ( .A1(n10575), .A2(n10574), .ZN(n10576) );
  OAI211_X1 U9277 ( .C1(n14876), .C2(n15229), .A(n14874), .B(n7145), .ZN(
        n14978) );
  NAND2_X1 U9278 ( .A1(n10371), .A2(n10370), .ZN(n10373) );
  NAND2_X1 U9279 ( .A1(n10160), .A2(n10161), .ZN(n10371) );
  NOR2_X2 U9280 ( .A1(n13829), .A2(n12555), .ZN(n13841) );
  NOR2_X2 U9281 ( .A1(n13830), .A2(n13831), .ZN(n13829) );
  NOR2_X1 U9282 ( .A1(n12571), .A2(n6724), .ZN(n12581) );
  NAND2_X1 U9283 ( .A1(n7570), .A2(n7567), .ZN(n8439) );
  NAND2_X1 U9284 ( .A1(n9276), .A2(n9211), .ZN(n9225) );
  NAND2_X1 U9285 ( .A1(n9274), .A2(n6900), .ZN(n6899) );
  OAI21_X1 U9286 ( .B1(n9158), .B2(n9161), .A(n7524), .ZN(n6927) );
  NAND2_X1 U9287 ( .A1(n6927), .A2(n6661), .ZN(n9262) );
  AOI21_X1 U9288 ( .B1(n8338), .B2(n6706), .A(n7976), .ZN(n7771) );
  NOR2_X1 U9289 ( .A1(n12905), .A2(n12906), .ZN(n12907) );
  AOI21_X1 U9290 ( .B1(n13012), .B2(n13011), .A(n13010), .ZN(n13013) );
  NAND2_X2 U9291 ( .A1(n15493), .A2(n15524), .ZN(n12068) );
  NAND2_X1 U9292 ( .A1(n7972), .A2(n7971), .ZN(n7991) );
  INV_X1 U9293 ( .A(n7217), .ZN(n7214) );
  NAND2_X1 U9294 ( .A1(n7215), .A2(n7213), .ZN(n7846) );
  OAI21_X1 U9295 ( .B1(n7879), .B2(n7223), .A(n7221), .ZN(n7912) );
  INV_X1 U9296 ( .A(n13091), .ZN(n6827) );
  NAND2_X1 U9297 ( .A1(n11269), .A2(n11270), .ZN(n11271) );
  NAND2_X1 U9298 ( .A1(n11775), .A2(n6848), .ZN(n15322) );
  INV_X1 U9299 ( .A(n11780), .ZN(n6850) );
  AOI21_X1 U9300 ( .B1(n10063), .B2(n11000), .A(n10993), .ZN(n15291) );
  NOR2_X2 U9301 ( .A1(n8371), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n14299) );
  NAND2_X1 U9302 ( .A1(n7512), .A2(n7511), .ZN(n8371) );
  NAND2_X1 U9303 ( .A1(n6861), .A2(n6859), .ZN(n14144) );
  NAND2_X1 U9304 ( .A1(n14184), .A2(n6819), .ZN(n14269) );
  NAND2_X1 U9305 ( .A1(n10542), .A2(n10546), .ZN(n10541) );
  NAND2_X1 U9306 ( .A1(n7601), .A2(n6774), .ZN(n10269) );
  NAND2_X1 U9307 ( .A1(n11276), .A2(n6739), .ZN(n11775) );
  NAND2_X1 U9308 ( .A1(n6852), .A2(n8629), .ZN(n10980) );
  NAND2_X1 U9309 ( .A1(n6853), .A2(n8616), .ZN(n10802) );
  NAND2_X1 U9310 ( .A1(n15133), .A2(n15134), .ZN(n6868) );
  OAI21_X1 U9311 ( .B1(n14185), .B2(n14261), .A(n14183), .ZN(n6820) );
  NAND2_X1 U9312 ( .A1(n15175), .A2(n15174), .ZN(n15173) );
  NAND2_X1 U9313 ( .A1(n7709), .A2(n7708), .ZN(n7645) );
  XNOR2_X1 U9314 ( .A(n7727), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15613) );
  INV_X1 U9315 ( .A(n15192), .ZN(n6834) );
  INV_X1 U9316 ( .A(n7719), .ZN(n7117) );
  NAND2_X1 U9317 ( .A1(n7115), .A2(n15184), .ZN(n15189) );
  NAND2_X1 U9318 ( .A1(n7122), .A2(n15173), .ZN(n7735) );
  XNOR2_X1 U9319 ( .A(n7735), .B(n7121), .ZN(n15179) );
  NAND2_X1 U9320 ( .A1(n6783), .A2(n6782), .ZN(n6781) );
  OR2_X1 U9321 ( .A1(n12426), .A2(n12425), .ZN(n12429) );
  INV_X1 U9322 ( .A(n9741), .ZN(n9743) );
  NAND3_X1 U9323 ( .A1(n6686), .A2(n6996), .A3(n6781), .ZN(n6995) );
  NAND2_X1 U9324 ( .A1(n12416), .A2(n12415), .ZN(n6783) );
  OR2_X1 U9325 ( .A1(n12445), .A2(n12446), .ZN(n6983) );
  NOR2_X2 U9326 ( .A1(n6633), .A2(n14980), .ZN(n14603) );
  NOR2_X1 U9327 ( .A1(n6624), .A2(n6695), .ZN(n7313) );
  INV_X2 U9328 ( .A(n8387), .ZN(n9750) );
  INV_X8 U9329 ( .A(n9750), .ZN(n7274) );
  AOI21_X1 U9330 ( .B1(n14628), .B2(n11951), .A(n11983), .ZN(n11962) );
  INV_X1 U9331 ( .A(n6980), .ZN(n6979) );
  XNOR2_X1 U9332 ( .A(n12356), .B(n11201), .ZN(n12499) );
  NOR2_X2 U9333 ( .A1(n10775), .A2(n10906), .ZN(n10809) );
  NAND2_X1 U9334 ( .A1(n10701), .A2(n10893), .ZN(n10775) );
  NAND2_X1 U9335 ( .A1(n6793), .A2(n6790), .ZN(P2_U3530) );
  OR2_X1 U9336 ( .A1(n14262), .A2(n6794), .ZN(n6793) );
  INV_X2 U9337 ( .A(n15404), .ZN(n6794) );
  NAND2_X1 U9338 ( .A1(n6797), .A2(n6795), .ZN(P2_U3498) );
  OR2_X1 U9339 ( .A1(n14262), .A2(n15391), .ZN(n6797) );
  INV_X1 U9340 ( .A(n7551), .ZN(n8760) );
  OR2_X1 U9341 ( .A1(n14166), .A2(n10143), .ZN(n10038) );
  NAND2_X1 U9342 ( .A1(n14034), .A2(n14013), .ZN(n14008) );
  OR2_X1 U9343 ( .A1(n10683), .A2(n10687), .ZN(n10684) );
  NAND2_X1 U9344 ( .A1(n6798), .A2(n7420), .ZN(n12476) );
  NAND3_X1 U9345 ( .A1(n6984), .A2(n6983), .A3(n6708), .ZN(n6798) );
  OR2_X1 U9346 ( .A1(n12421), .A2(n12424), .ZN(n12426) );
  INV_X1 U9347 ( .A(n12397), .ZN(n7424) );
  NAND2_X1 U9348 ( .A1(n12329), .A2(n12328), .ZN(n6818) );
  NAND2_X1 U9349 ( .A1(n12322), .A2(n12323), .ZN(n12329) );
  AOI21_X1 U9350 ( .B1(n12423), .B2(n12422), .A(n12420), .ZN(n12421) );
  NAND2_X1 U9351 ( .A1(n6992), .A2(n6813), .ZN(n6991) );
  NAND2_X2 U9352 ( .A1(n9748), .A2(n15023), .ZN(n12289) );
  NAND2_X1 U9353 ( .A1(n10459), .A2(n10458), .ZN(n10569) );
  NAND2_X1 U9354 ( .A1(n11296), .A2(n11295), .ZN(n11429) );
  INV_X1 U9355 ( .A(n9526), .ZN(n7270) );
  NAND2_X1 U9356 ( .A1(n6823), .A2(n6822), .ZN(n11997) );
  NAND2_X1 U9357 ( .A1(n7276), .A2(n7275), .ZN(n11653) );
  OAI21_X1 U9358 ( .B1(n10457), .B2(n14429), .A(n12340), .ZN(n10459) );
  OAI22_X1 U9359 ( .A1(n12487), .A2(n10316), .B1(n12307), .B2(n14844), .ZN(
        n10332) );
  NAND2_X1 U9360 ( .A1(n12788), .A2(n12789), .ZN(n7180) );
  OR2_X1 U9361 ( .A1(n6603), .A2(n9333), .ZN(n7776) );
  NAND2_X1 U9362 ( .A1(n10373), .A2(n12012), .ZN(n12018) );
  NAND2_X1 U9363 ( .A1(n12542), .A2(n7405), .ZN(n15103) );
  NAND2_X1 U9364 ( .A1(n11478), .A2(n7367), .ZN(n7366) );
  XNOR2_X1 U9365 ( .A(n10009), .B(n10010), .ZN(n14329) );
  OAI21_X1 U9366 ( .B1(n10295), .B2(n7051), .A(n7049), .ZN(n7053) );
  NAND2_X1 U9367 ( .A1(n7257), .A2(n10294), .ZN(n10436) );
  NAND3_X1 U9368 ( .A1(n7044), .A2(P3_REG1_REG_13__SCAN_IN), .A3(n12940), .ZN(
        n7045) );
  NOR2_X1 U9369 ( .A1(n11094), .A2(n15594), .ZN(n11252) );
  NAND2_X1 U9370 ( .A1(n11379), .A2(n6712), .ZN(n7034) );
  NAND2_X1 U9371 ( .A1(n12359), .A2(n12360), .ZN(n12358) );
  OAI21_X1 U9372 ( .B1(n12329), .B2(n12328), .A(n6816), .ZN(n12333) );
  NAND2_X1 U9373 ( .A1(n6818), .A2(n6817), .ZN(n6816) );
  NAND2_X4 U9374 ( .A1(n9748), .A2(n9747), .ZN(n11986) );
  NAND2_X1 U9375 ( .A1(n12426), .A2(n12425), .ZN(n7406) );
  NAND2_X1 U9376 ( .A1(n7406), .A2(n12427), .ZN(n12428) );
  NAND2_X1 U9377 ( .A1(n6943), .A2(n6942), .ZN(n14132) );
  NAND2_X1 U9378 ( .A1(n6960), .A2(n6958), .ZN(n15129) );
  NAND2_X1 U9379 ( .A1(n6979), .A2(n6981), .ZN(n6977) );
  OAI21_X1 U9380 ( .B1(n8556), .B2(n6981), .A(n8570), .ZN(n6980) );
  NOR2_X1 U9381 ( .A1(n14110), .A2(n14111), .ZN(n6964) );
  NAND2_X1 U9382 ( .A1(n14069), .A2(n8968), .ZN(n8971) );
  NAND2_X1 U9383 ( .A1(n7384), .A2(n6934), .ZN(n6933) );
  OAI21_X1 U9384 ( .B1(n6937), .B2(n6936), .A(n13858), .ZN(n6935) );
  NOR2_X2 U9385 ( .A1(n12581), .A2(n12580), .ZN(n12585) );
  NAND2_X1 U9386 ( .A1(n6971), .A2(n6969), .ZN(n6968) );
  INV_X1 U9387 ( .A(n13781), .ZN(n7390) );
  INV_X1 U9388 ( .A(n7478), .ZN(n7477) );
  AOI22_X2 U9389 ( .A1(n12862), .A2(n12863), .B1(n13110), .B2(n12737), .ZN(
        n12770) );
  NAND2_X1 U9390 ( .A1(n13210), .A2(n8289), .ZN(n13195) );
  NAND2_X1 U9391 ( .A1(n8381), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U9392 ( .A1(n13245), .A2(n12214), .ZN(n7066) );
  NAND2_X1 U9393 ( .A1(n8271), .A2(n7622), .ZN(n8274) );
  NAND2_X1 U9394 ( .A1(n7807), .A2(n7806), .ZN(n7820) );
  NAND2_X1 U9395 ( .A1(n7068), .A2(n7067), .ZN(n13167) );
  INV_X1 U9396 ( .A(n7087), .ZN(n7086) );
  OAI22_X1 U9397 ( .A1(n13557), .A2(n8278), .B1(n13582), .B2(n13680), .ZN(
        n13260) );
  OAI21_X2 U9398 ( .B1(n10499), .B2(n10498), .A(n10497), .ZN(n14428) );
  NAND2_X1 U9399 ( .A1(n11477), .A2(n11476), .ZN(n11478) );
  AOI21_X1 U9400 ( .B1(n7345), .B2(n7344), .A(n6703), .ZN(n7341) );
  NOR2_X1 U9401 ( .A1(n15189), .A2(n15190), .ZN(n15188) );
  NAND2_X1 U9402 ( .A1(n11154), .A2(n11153), .ZN(n11156) );
  NOR2_X2 U9403 ( .A1(n15604), .A2(n7717), .ZN(n7720) );
  INV_X1 U9404 ( .A(n7708), .ZN(n6838) );
  NAND2_X1 U9405 ( .A1(n11368), .A2(n11367), .ZN(n11671) );
  AND3_X1 U9406 ( .A1(n9806), .A2(n9805), .A3(n9804), .ZN(n9847) );
  NAND2_X2 U9407 ( .A1(n12694), .A2(n12693), .ZN(n14436) );
  INV_X1 U9408 ( .A(n12935), .ZN(n6843) );
  AOI21_X1 U9409 ( .B1(n10429), .B2(n10428), .A(n10427), .ZN(n10435) );
  NAND2_X2 U9410 ( .A1(n9323), .A2(n9733), .ZN(n9797) );
  XNOR2_X2 U9411 ( .A(n9322), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9733) );
  NOR2_X1 U9412 ( .A1(n11767), .A2(n11766), .ZN(n12905) );
  NOR2_X1 U9413 ( .A1(n11086), .A2(n11085), .ZN(n11087) );
  INV_X1 U9414 ( .A(n13009), .ZN(n13010) );
  NAND2_X1 U9415 ( .A1(n12985), .A2(n12986), .ZN(n13009) );
  NAND2_X1 U9416 ( .A1(n7156), .A2(n7155), .ZN(n14651) );
  OR2_X2 U9417 ( .A1(n11306), .A2(n12375), .ZN(n11440) );
  INV_X1 U9418 ( .A(n15232), .ZN(n12303) );
  NOR2_X1 U9419 ( .A1(n10587), .A2(n12351), .ZN(n10743) );
  NAND2_X1 U9420 ( .A1(n14125), .A2(n8992), .ZN(n14126) );
  NAND2_X1 U9421 ( .A1(n10809), .A2(n8991), .ZN(n15136) );
  NAND2_X1 U9422 ( .A1(n11622), .A2(n11626), .ZN(n11708) );
  INV_X1 U9423 ( .A(n9941), .ZN(n15360) );
  NOR2_X1 U9424 ( .A1(n7136), .A2(n7132), .ZN(n7135) );
  XNOR2_X2 U9425 ( .A(n8245), .B(n7753), .ZN(n10784) );
  NAND2_X1 U9426 ( .A1(n10996), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11269) );
  XNOR2_X1 U9427 ( .A(n6851), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n11794) );
  OR2_X1 U9428 ( .A1(n13955), .A2(n11780), .ZN(n6851) );
  NAND2_X1 U9429 ( .A1(n10802), .A2(n10803), .ZN(n6852) );
  NAND2_X1 U9430 ( .A1(n10769), .A2(n10770), .ZN(n6853) );
  NAND2_X1 U9431 ( .A1(n14188), .A2(n8878), .ZN(n13974) );
  NOR2_X1 U9432 ( .A1(n7604), .A2(n10681), .ZN(n6858) );
  NAND2_X1 U9433 ( .A1(n8706), .A2(n6862), .ZN(n6861) );
  MUX2_X1 U9434 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8387), .Z(n8385) );
  NAND4_X1 U9435 ( .A1(n13070), .A2(n7775), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n6872) );
  NAND4_X1 U9436 ( .A1(n11799), .A2(n7774), .A3(n11699), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U9437 ( .A1(n7633), .A2(n12922), .ZN(n12912) );
  INV_X1 U9438 ( .A(n6880), .ZN(n12924) );
  NAND3_X1 U9439 ( .A1(n6884), .A2(n6886), .A3(n6881), .ZN(n11237) );
  NAND3_X1 U9440 ( .A1(n6884), .A2(n6882), .A3(n6881), .ZN(n7183) );
  INV_X1 U9441 ( .A(n6895), .ZN(n13029) );
  INV_X1 U9442 ( .A(n13030), .ZN(n6894) );
  OAI21_X1 U9443 ( .B1(n9302), .B2(n6899), .A(n9303), .ZN(n9307) );
  NAND3_X1 U9444 ( .A1(n8361), .A2(n8360), .A3(n8359), .ZN(n6966) );
  NAND2_X1 U9445 ( .A1(n6709), .A2(n8710), .ZN(n6965) );
  NAND2_X1 U9446 ( .A1(n6903), .A2(n6901), .ZN(n9056) );
  INV_X1 U9447 ( .A(n6905), .ZN(n6902) );
  NAND2_X1 U9448 ( .A1(n6682), .A2(n6904), .ZN(n6903) );
  NAND2_X1 U9449 ( .A1(n6905), .A2(n7522), .ZN(n6904) );
  OAI21_X1 U9450 ( .B1(n9077), .B2(n6908), .A(n6906), .ZN(n9087) );
  NAND2_X1 U9451 ( .A1(n6916), .A2(n6727), .ZN(n7543) );
  NAND3_X1 U9452 ( .A1(n9142), .A2(n9143), .A3(n6725), .ZN(n6916) );
  OAI21_X1 U9453 ( .B1(n9129), .B2(n6923), .A(n6918), .ZN(n9134) );
  OAI21_X1 U9454 ( .B1(n9097), .B2(n6925), .A(n6924), .ZN(n9103) );
  INV_X1 U9455 ( .A(n9096), .ZN(n6926) );
  OAI22_X1 U9456 ( .A1(n9064), .A2(n6664), .B1(n9063), .B2(n6928), .ZN(n9069)
         );
  INV_X1 U9457 ( .A(n9062), .ZN(n6928) );
  NOR2_X1 U9458 ( .A1(n9898), .A2(n11795), .ZN(n9020) );
  NAND2_X1 U9459 ( .A1(n7384), .A2(n7382), .ZN(n13779) );
  NOR2_X1 U9460 ( .A1(n6938), .A2(n13782), .ZN(n6937) );
  MUX2_X1 U9461 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8387), .Z(n8397) );
  NAND2_X1 U9462 ( .A1(n11628), .A2(n6945), .ZN(n6943) );
  INV_X1 U9463 ( .A(n9280), .ZN(n6953) );
  XNOR2_X1 U9464 ( .A(n6955), .B(n8977), .ZN(n6954) );
  INV_X1 U9465 ( .A(n13978), .ZN(n6957) );
  NAND2_X1 U9466 ( .A1(n8953), .A2(n6961), .ZN(n6960) );
  NAND3_X2 U9467 ( .A1(n8516), .A2(n8709), .A3(n8365), .ZN(n6967) );
  NOR2_X2 U9468 ( .A1(n6965), .A2(n6967), .ZN(n7512) );
  OAI21_X1 U9469 ( .B1(n8601), .B2(n6969), .A(n6971), .ZN(n8647) );
  NAND3_X1 U9470 ( .A1(n6970), .A2(n6968), .A3(n7556), .ZN(n7553) );
  NAND2_X1 U9471 ( .A1(n8601), .A2(n6971), .ZN(n6970) );
  INV_X1 U9472 ( .A(n8402), .ZN(n6981) );
  NAND2_X1 U9473 ( .A1(n6976), .A2(n6979), .ZN(n8572) );
  OR2_X1 U9474 ( .A1(n8557), .A2(n6981), .ZN(n6976) );
  NAND3_X1 U9475 ( .A1(n6978), .A2(n6977), .A3(n8405), .ZN(n8584) );
  NAND2_X1 U9476 ( .A1(n8557), .A2(n6979), .ZN(n6978) );
  NAND3_X1 U9477 ( .A1(n8424), .A2(n7592), .A3(n7590), .ZN(n6982) );
  NAND2_X1 U9478 ( .A1(n6985), .A2(n12444), .ZN(n6984) );
  NAND2_X1 U9479 ( .A1(n12445), .A2(n12446), .ZN(n6985) );
  NAND2_X1 U9480 ( .A1(n12436), .A2(n6702), .ZN(n6986) );
  INV_X1 U9481 ( .A(n14788), .ZN(n7426) );
  NAND2_X1 U9482 ( .A1(n6991), .A2(n6989), .ZN(n12408) );
  AOI21_X1 U9483 ( .B1(n7427), .B2(n14788), .A(n6990), .ZN(n6989) );
  NAND2_X1 U9484 ( .A1(n6994), .A2(n6993), .ZN(n6992) );
  NAND2_X1 U9485 ( .A1(n12384), .A2(n12383), .ZN(n6993) );
  NAND2_X1 U9486 ( .A1(n6995), .A2(n6997), .ZN(n12423) );
  MUX2_X1 U9487 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8387), .Z(n8393) );
  NAND2_X1 U9488 ( .A1(n13556), .A2(n7003), .ZN(n7000) );
  NAND2_X1 U9489 ( .A1(n7000), .A2(n7001), .ZN(n13253) );
  NAND2_X1 U9490 ( .A1(n15434), .A2(n7010), .ZN(n7006) );
  NAND2_X1 U9491 ( .A1(n7006), .A2(n7007), .ZN(n15069) );
  NAND2_X1 U9492 ( .A1(n11015), .A2(n7017), .ZN(n7014) );
  NAND2_X1 U9493 ( .A1(n7014), .A2(n7015), .ZN(n11400) );
  NAND2_X4 U9494 ( .A1(n8297), .A2(n8298), .ZN(n10179) );
  NAND3_X2 U9495 ( .A1(n7021), .A2(n7020), .A3(n7023), .ZN(n8297) );
  NAND2_X1 U9496 ( .A1(n8308), .A2(n7022), .ZN(n7020) );
  OR2_X1 U9497 ( .A1(n8308), .A2(n7026), .ZN(n7021) );
  NAND2_X2 U9498 ( .A1(n7027), .A2(n13233), .ZN(n13667) );
  XNOR2_X2 U9499 ( .A(n7029), .B(n13093), .ZN(n13621) );
  NAND2_X2 U9500 ( .A1(n7030), .A2(n12180), .ZN(n7029) );
  OR2_X2 U9501 ( .A1(n13629), .A2(n7476), .ZN(n7030) );
  INV_X1 U9502 ( .A(n11379), .ZN(n7040) );
  NAND2_X1 U9503 ( .A1(n11379), .A2(n6625), .ZN(n7031) );
  INV_X1 U9504 ( .A(n7033), .ZN(n7032) );
  INV_X1 U9505 ( .A(n7045), .ZN(n12941) );
  XNOR2_X2 U9506 ( .A(n13032), .B(n7265), .ZN(n13021) );
  INV_X1 U9507 ( .A(n7053), .ZN(n11092) );
  NAND2_X1 U9508 ( .A1(n6697), .A2(n10240), .ZN(n7056) );
  OAI211_X2 U9509 ( .C1(n7160), .C2(n7057), .A(n7159), .B(n7266), .ZN(n10252)
         );
  NAND2_X1 U9510 ( .A1(n15499), .A2(n7059), .ZN(n15476) );
  NAND2_X1 U9511 ( .A1(n15462), .A2(n7062), .ZN(n7060) );
  NAND2_X1 U9512 ( .A1(n7061), .A2(n7060), .ZN(n15448) );
  AOI21_X1 U9513 ( .B1(n7062), .B2(n7064), .A(n6646), .ZN(n7061) );
  OAI21_X1 U9514 ( .B1(n8263), .B2(n7064), .A(n11171), .ZN(n7063) );
  NAND2_X1 U9515 ( .A1(n7066), .A2(n7065), .ZN(n13230) );
  NAND2_X1 U9516 ( .A1(n8292), .A2(n7069), .ZN(n7068) );
  OR2_X1 U9517 ( .A1(n7819), .A2(n9369), .ZN(n7852) );
  OR2_X1 U9518 ( .A1(n7819), .A2(n9379), .ZN(n7865) );
  OR2_X1 U9519 ( .A1(n6603), .A2(n9371), .ZN(n7885) );
  NAND3_X1 U9520 ( .A1(n7752), .A2(n7480), .A3(n7755), .ZN(n7478) );
  OAI21_X1 U9521 ( .B1(n15438), .B2(n7086), .A(n7084), .ZN(n13557) );
  NAND3_X1 U9522 ( .A1(n8395), .A2(n8541), .A3(n8527), .ZN(n7100) );
  NAND2_X1 U9523 ( .A1(n15036), .A2(n15037), .ZN(n7131) );
  NOR2_X2 U9524 ( .A1(n14053), .A2(n14031), .ZN(n14034) );
  NOR2_X2 U9525 ( .A1(n13967), .A2(n14266), .ZN(n13970) );
  NOR2_X2 U9526 ( .A1(n6631), .A2(n14237), .ZN(n14125) );
  NOR2_X2 U9527 ( .A1(n10608), .A2(n10704), .ZN(n10701) );
  INV_X1 U9528 ( .A(n14166), .ZN(n9900) );
  NOR2_X2 U9529 ( .A1(n14689), .A2(n14987), .ZN(n7156) );
  NAND2_X2 U9530 ( .A1(n7274), .A2(P1_U3086), .ZN(n15024) );
  MUX2_X1 U9531 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7620), .Z(n8415) );
  MUX2_X1 U9532 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n7620), .Z(n8432) );
  MUX2_X1 U9533 ( .A(n11578), .B(n11890), .S(n7620), .Z(n8447) );
  MUX2_X1 U9534 ( .A(n11723), .B(n13373), .S(n7620), .Z(n8452) );
  MUX2_X1 U9535 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n7620), .Z(n8865) );
  NAND2_X1 U9536 ( .A1(n7160), .A2(P3_IR_REG_2__SCAN_IN), .ZN(n7159) );
  NAND2_X1 U9537 ( .A1(n12280), .A2(n7172), .ZN(n7171) );
  OAI211_X1 U9538 ( .C1(n12280), .C2(n7173), .A(n7171), .B(n12284), .ZN(
        P3_U3169) );
  XNOR2_X1 U9539 ( .A(n12280), .B(n12279), .ZN(n12755) );
  INV_X1 U9540 ( .A(n11596), .ZN(n7176) );
  XNOR2_X1 U9541 ( .A(n11591), .B(P3_B_REG_SCAN_IN), .ZN(n7177) );
  NAND3_X1 U9542 ( .A1(n7178), .A2(n13503), .A3(n8337), .ZN(n8315) );
  NAND3_X1 U9543 ( .A1(n10211), .A2(P3_REG2_REG_1__SCAN_IN), .A3(n7181), .ZN(
        n10212) );
  NAND2_X1 U9544 ( .A1(n7182), .A2(n10175), .ZN(n10199) );
  INV_X1 U9545 ( .A(n7188), .ZN(n11357) );
  INV_X1 U9546 ( .A(n11356), .ZN(n7187) );
  NAND2_X1 U9547 ( .A1(n10244), .A2(n10213), .ZN(n7192) );
  NAND2_X1 U9548 ( .A1(n7193), .A2(n7194), .ZN(n15426) );
  NAND3_X1 U9549 ( .A1(n10244), .A2(n10213), .A3(n7258), .ZN(n7193) );
  INV_X1 U9550 ( .A(n7199), .ZN(n11755) );
  INV_X1 U9551 ( .A(n7197), .ZN(n12909) );
  NAND2_X1 U9552 ( .A1(n7199), .A2(n7198), .ZN(n7197) );
  OR2_X1 U9553 ( .A1(n11753), .A2(n11754), .ZN(n7199) );
  INV_X1 U9554 ( .A(n7793), .ZN(n7205) );
  NAND2_X1 U9555 ( .A1(n7204), .A2(n7794), .ZN(n7807) );
  XNOR2_X1 U9556 ( .A(n7206), .B(n7795), .ZN(n9373) );
  NAND2_X1 U9557 ( .A1(n7946), .A2(n7945), .ZN(n7958) );
  OAI21_X1 U9558 ( .B1(n8140), .B2(n7253), .A(n7251), .ZN(n8152) );
  NOR2_X1 U9559 ( .A1(n11667), .A2(n11668), .ZN(n11753) );
  AOI21_X1 U9560 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n13019), .A(n13002), .ZN(
        n13028) );
  NAND2_X1 U9561 ( .A1(n10212), .A2(n10211), .ZN(n10245) );
  NAND2_X1 U9562 ( .A1(n8109), .A2(n8097), .ZN(n8098) );
  NOR2_X1 U9563 ( .A1(n11664), .A2(n7041), .ZN(n11754) );
  NAND2_X1 U9564 ( .A1(n11666), .A2(n11665), .ZN(n11668) );
  NOR2_X1 U9565 ( .A1(n15426), .A2(n15487), .ZN(n15424) );
  INV_X1 U9566 ( .A(n11754), .ZN(n11666) );
  AND2_X2 U9567 ( .A1(n12325), .A2(n10850), .ZN(n11070) );
  OAI21_X1 U9568 ( .B1(SI_1_), .B2(n8380), .A(n8384), .ZN(n8476) );
  INV_X1 U9569 ( .A(n12044), .ZN(n13695) );
  OAI21_X1 U9570 ( .B1(n10208), .B2(n10209), .A(n7257), .ZN(n10220) );
  NAND2_X1 U9571 ( .A1(n10208), .A2(n10209), .ZN(n7257) );
  NOR2_X2 U9572 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n7268) );
  INV_X1 U9573 ( .A(n9527), .ZN(n7269) );
  NOR2_X1 U9574 ( .A1(n9752), .A2(n7274), .ZN(n7273) );
  NAND2_X2 U9575 ( .A1(n9559), .A2(n15027), .ZN(n9751) );
  INV_X1 U9576 ( .A(n7272), .ZN(n7271) );
  NAND2_X2 U9577 ( .A1(n9751), .A2(n7274), .ZN(n12458) );
  NAND2_X1 U9578 ( .A1(n11429), .A2(n6616), .ZN(n7276) );
  NAND2_X1 U9579 ( .A1(n10723), .A2(n10722), .ZN(n10725) );
  NAND2_X1 U9580 ( .A1(n14820), .A2(n7293), .ZN(n7292) );
  NAND2_X1 U9581 ( .A1(n14686), .A2(n7295), .ZN(n11978) );
  NAND2_X1 U9582 ( .A1(n11156), .A2(n7306), .ZN(n7305) );
  AND2_X2 U9583 ( .A1(n14628), .A2(n7310), .ZN(n14596) );
  NAND2_X1 U9584 ( .A1(n14626), .A2(n14625), .ZN(n14628) );
  NAND2_X1 U9585 ( .A1(n10576), .A2(n6642), .ZN(n7314) );
  NOR2_X1 U9586 ( .A1(n7316), .A2(n7319), .ZN(n7317) );
  NOR2_X1 U9587 ( .A1(n9746), .A2(n7318), .ZN(n7316) );
  NAND2_X1 U9588 ( .A1(n14700), .A2(n7324), .ZN(n14681) );
  NAND2_X1 U9589 ( .A1(n14749), .A2(n7325), .ZN(n11880) );
  NOR2_X1 U9590 ( .A1(n14734), .A2(n7326), .ZN(n7325) );
  NAND2_X1 U9591 ( .A1(n14406), .A2(n7330), .ZN(n7329) );
  NAND2_X1 U9592 ( .A1(n14377), .A2(n7335), .ZN(n7334) );
  NAND2_X1 U9593 ( .A1(n7342), .A2(n7341), .ZN(n10099) );
  NAND2_X1 U9594 ( .A1(n7343), .A2(n7345), .ZN(n7342) );
  INV_X1 U9595 ( .A(n9817), .ZN(n7343) );
  INV_X1 U9596 ( .A(n10003), .ZN(n7346) );
  NAND2_X1 U9597 ( .A1(n10004), .A2(n7345), .ZN(n10094) );
  NAND2_X1 U9598 ( .A1(n9817), .A2(n9818), .ZN(n10004) );
  NAND2_X1 U9599 ( .A1(n14436), .A2(n14437), .ZN(n7354) );
  OAI211_X1 U9600 ( .C1(n14436), .C2(n7352), .A(n7348), .B(n7347), .ZN(n12719)
         );
  NAND2_X1 U9601 ( .A1(n14436), .A2(n6705), .ZN(n7347) );
  OAI21_X1 U9602 ( .B1(n7353), .B2(n7358), .A(n7349), .ZN(n7348) );
  NAND2_X1 U9603 ( .A1(n7353), .A2(n7350), .ZN(n7349) );
  NAND3_X1 U9604 ( .A1(n11800), .A2(n9913), .A3(n9924), .ZN(n10161) );
  NOR2_X1 U9605 ( .A1(n13841), .A2(n13840), .ZN(n13839) );
  NAND2_X1 U9606 ( .A1(n13841), .A2(n7385), .ZN(n7384) );
  NAND2_X1 U9607 ( .A1(n12561), .A2(n12562), .ZN(n7393) );
  NAND2_X2 U9608 ( .A1(n7402), .A2(n9898), .ZN(n10158) );
  NAND3_X1 U9609 ( .A1(n8938), .A2(n11795), .A3(n9898), .ZN(n7402) );
  XNOR2_X2 U9610 ( .A(n8923), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8938) );
  AND2_X1 U9611 ( .A1(n10382), .A2(n10377), .ZN(n7404) );
  NAND3_X1 U9612 ( .A1(n12307), .A2(n14844), .A3(n12339), .ZN(n7407) );
  NAND3_X1 U9613 ( .A1(n14851), .A2(n6588), .A3(n12308), .ZN(n7408) );
  OAI21_X2 U9614 ( .B1(n12299), .B2(n11165), .A(n12462), .ZN(n12339) );
  XNOR2_X1 U9615 ( .A(n6590), .B(n14768), .ZN(n12299) );
  OR2_X1 U9616 ( .A1(n11649), .A2(n14479), .ZN(n7411) );
  OAI21_X1 U9617 ( .B1(n12344), .B2(n7417), .A(n7416), .ZN(n12349) );
  NAND2_X1 U9618 ( .A1(n7415), .A2(n7413), .ZN(n12347) );
  NAND2_X1 U9619 ( .A1(n12344), .A2(n7416), .ZN(n7415) );
  NAND2_X1 U9620 ( .A1(n7434), .A2(n7432), .ZN(n12371) );
  AOI21_X1 U9621 ( .B1(n7436), .B2(n7435), .A(n7433), .ZN(n7432) );
  NAND2_X1 U9622 ( .A1(n12366), .A2(n7435), .ZN(n7434) );
  NAND2_X1 U9623 ( .A1(n12431), .A2(n7440), .ZN(n7437) );
  NAND2_X1 U9624 ( .A1(n7437), .A2(n7438), .ZN(n12434) );
  OAI22_X1 U9625 ( .A1(n12353), .A2(n7446), .B1(n7445), .B2(n12354), .ZN(
        n12359) );
  NAND2_X1 U9626 ( .A1(n7449), .A2(n15520), .ZN(n10356) );
  OAI21_X1 U9627 ( .B1(n12064), .B2(n12183), .A(n7450), .ZN(n12069) );
  NAND2_X1 U9628 ( .A1(n7453), .A2(n7451), .ZN(P3_U3296) );
  NAND2_X1 U9629 ( .A1(n7452), .A2(n6740), .ZN(n7451) );
  XNOR2_X1 U9630 ( .A(n12051), .B(n13073), .ZN(n7452) );
  INV_X1 U9631 ( .A(n7454), .ZN(n7453) );
  OAI211_X1 U9632 ( .C1(n12229), .C2(n7458), .A(n7456), .B(n7455), .ZN(n7454)
         );
  NAND3_X1 U9633 ( .A1(n12229), .A2(n12231), .A3(n15527), .ZN(n7455) );
  INV_X1 U9634 ( .A(n7457), .ZN(n7456) );
  NAND2_X1 U9635 ( .A1(n12227), .A2(n12228), .ZN(n7461) );
  OAI21_X1 U9636 ( .B1(n13629), .B2(n7468), .A(n7467), .ZN(n12019) );
  NAND2_X1 U9637 ( .A1(n7471), .A2(n7469), .ZN(n12046) );
  NAND2_X1 U9638 ( .A1(n13629), .A2(n7472), .ZN(n7471) );
  AND2_X2 U9639 ( .A1(n13685), .A2(n12118), .ZN(n13586) );
  AND2_X2 U9640 ( .A1(n8308), .A2(n7022), .ZN(n7762) );
  NOR2_X2 U9641 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n8546) );
  AND2_X2 U9642 ( .A1(n8480), .A2(n8546), .ZN(n8516) );
  NOR2_X2 U9643 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8480) );
  OAI21_X1 U9644 ( .B1(n14109), .B2(n7487), .A(n7484), .ZN(n14080) );
  INV_X1 U9645 ( .A(n8967), .ZN(n7491) );
  NAND2_X1 U9646 ( .A1(n7493), .A2(n7492), .ZN(n8951) );
  NAND2_X1 U9647 ( .A1(n10611), .A2(n7494), .ZN(n7492) );
  NAND2_X1 U9648 ( .A1(n14024), .A2(n7504), .ZN(n7501) );
  NAND2_X1 U9649 ( .A1(n7501), .A2(n7502), .ZN(n13993) );
  NAND2_X1 U9650 ( .A1(n15112), .A2(n7509), .ZN(n7508) );
  INV_X1 U9651 ( .A(n12011), .ZN(n13913) );
  NAND3_X1 U9652 ( .A1(n8539), .A2(n8538), .A3(n7514), .ZN(n7513) );
  INV_X1 U9653 ( .A(n8520), .ZN(n8486) );
  NAND2_X1 U9654 ( .A1(n7518), .A2(n7517), .ZN(n7516) );
  NAND2_X1 U9655 ( .A1(n9124), .A2(n9123), .ZN(n7518) );
  INV_X1 U9656 ( .A(n9123), .ZN(n7520) );
  INV_X1 U9657 ( .A(n9124), .ZN(n7521) );
  AOI21_X1 U9658 ( .B1(n9056), .B2(n9055), .A(n9054), .ZN(n9058) );
  INV_X1 U9659 ( .A(n9164), .ZN(n7529) );
  INV_X1 U9660 ( .A(n9075), .ZN(n7532) );
  NAND2_X1 U9661 ( .A1(n9134), .A2(n7536), .ZN(n7533) );
  NAND2_X1 U9662 ( .A1(n7533), .A2(n7534), .ZN(n9139) );
  NAND2_X1 U9663 ( .A1(n9039), .A2(n9038), .ZN(n7542) );
  NAND2_X1 U9664 ( .A1(n7541), .A2(n7538), .ZN(n9046) );
  INV_X1 U9665 ( .A(n9039), .ZN(n7539) );
  INV_X1 U9666 ( .A(n9038), .ZN(n7540) );
  NAND3_X1 U9667 ( .A1(n7542), .A2(n9034), .A3(n9035), .ZN(n7541) );
  NAND2_X1 U9668 ( .A1(n7543), .A2(n6726), .ZN(n9160) );
  NAND2_X1 U9669 ( .A1(n7545), .A2(n7548), .ZN(n9117) );
  NAND3_X1 U9670 ( .A1(n9108), .A2(n7546), .A3(n9107), .ZN(n7545) );
  OR2_X1 U9671 ( .A1(n9087), .A2(n6710), .ZN(n7552) );
  NAND2_X1 U9672 ( .A1(n7553), .A2(n7554), .ZN(n8422) );
  NAND2_X1 U9673 ( .A1(n9206), .A2(n9263), .ZN(n9276) );
  NAND2_X1 U9674 ( .A1(n8817), .A2(n7564), .ZN(n7561) );
  NAND2_X1 U9675 ( .A1(n7561), .A2(n7562), .ZN(n8842) );
  NAND2_X1 U9676 ( .A1(n8708), .A2(n6693), .ZN(n7570) );
  NAND2_X1 U9677 ( .A1(n8708), .A2(n8707), .ZN(n7577) );
  NAND2_X1 U9678 ( .A1(n8779), .A2(n7579), .ZN(n7578) );
  NAND2_X1 U9679 ( .A1(n7580), .A2(n8440), .ZN(n8792) );
  NAND2_X1 U9680 ( .A1(n8779), .A2(n8438), .ZN(n7580) );
  OR2_X1 U9681 ( .A1(n8868), .A2(n7589), .ZN(n7581) );
  NAND2_X1 U9682 ( .A1(n8868), .A2(n7586), .ZN(n7585) );
  NAND2_X1 U9683 ( .A1(n8424), .A2(n8423), .ZN(n8676) );
  INV_X1 U9684 ( .A(n7592), .ZN(n7591) );
  INV_X1 U9685 ( .A(n8675), .ZN(n7593) );
  NAND2_X1 U9686 ( .A1(n10662), .A2(n7602), .ZN(n7601) );
  NAND2_X1 U9687 ( .A1(n10680), .A2(n8540), .ZN(n10267) );
  NAND2_X1 U9688 ( .A1(n10682), .A2(n10681), .ZN(n10680) );
  NAND2_X1 U9689 ( .A1(n14144), .A2(n7617), .ZN(n7616) );
  NAND2_X1 U9690 ( .A1(n7616), .A2(n7614), .ZN(n8790) );
  INV_X1 U9691 ( .A(n12746), .ZN(n12252) );
  OAI21_X1 U9692 ( .B1(n14181), .B2(n15331), .A(n9003), .ZN(n9004) );
  INV_X1 U9693 ( .A(n12618), .ZN(n11738) );
  CLKBUF_X1 U9694 ( .A(n9447), .Z(n10258) );
  AND2_X1 U9695 ( .A1(n9816), .A2(n9815), .ZN(n9840) );
  CLKBUF_X1 U9696 ( .A(n14761), .Z(n14762) );
  NAND2_X1 U9697 ( .A1(n11473), .A2(n11472), .ZN(n11477) );
  NAND2_X1 U9698 ( .A1(n10317), .A2(n12309), .ZN(n10334) );
  AOI21_X2 U9699 ( .B1(n12839), .B2(n13197), .A(n12278), .ZN(n12280) );
  INV_X1 U9700 ( .A(n12359), .ZN(n12362) );
  NAND2_X1 U9701 ( .A1(n9516), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9517) );
  AOI21_X1 U9702 ( .B1(n12709), .B2(n14851), .A(n9810), .ZN(n9812) );
  AND4_X2 U9703 ( .A1(n9773), .A2(n9772), .A3(n9771), .A4(n9770), .ZN(n12315)
         );
  CLKBUF_X1 U9704 ( .A(n10371), .Z(n12013) );
  OAI211_X1 U9705 ( .C1(P1_B_REG_SCAN_IN), .C2(n9397), .A(n9733), .B(n9398), 
        .ZN(n9738) );
  XNOR2_X1 U9706 ( .A(n9294), .B(n8897), .ZN(n14182) );
  INV_X1 U9707 ( .A(n10130), .ZN(n9905) );
  NAND2_X1 U9708 ( .A1(n9102), .A2(n9101), .ZN(n9108) );
  AND2_X1 U9709 ( .A1(n11104), .A2(n9297), .ZN(n10146) );
  NAND2_X1 U9710 ( .A1(n8908), .A2(n8907), .ZN(n14314) );
  XNOR2_X1 U9711 ( .A(n12579), .B(n12578), .ZN(n12571) );
  NAND2_X1 U9712 ( .A1(n9026), .A2(n9265), .ZN(n9025) );
  AOI21_X1 U9713 ( .B1(n9301), .B2(n10146), .A(n9300), .ZN(n9302) );
  NAND2_X1 U9714 ( .A1(n9275), .A2(n9273), .ZN(n9274) );
  INV_X1 U9715 ( .A(n8536), .ZN(n9204) );
  INV_X2 U9716 ( .A(n15530), .ZN(n15489) );
  AND2_X2 U9717 ( .A1(n9014), .A2(n10487), .ZN(n15603) );
  AND2_X1 U9718 ( .A1(n8347), .A2(n8346), .ZN(n7621) );
  NAND2_X1 U9719 ( .A1(n15582), .A2(n15523), .ZN(n13741) );
  NAND2_X1 U9720 ( .A1(n13572), .A2(n8272), .ZN(n7622) );
  AND2_X1 U9721 ( .A1(n9368), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7623) );
  AND2_X1 U9722 ( .A1(n12223), .A2(n12049), .ZN(n7624) );
  OR2_X1 U9723 ( .A1(n13695), .A2(n12886), .ZN(n7625) );
  OR2_X1 U9724 ( .A1(n13640), .A2(n12725), .ZN(n7626) );
  NAND2_X1 U9725 ( .A1(n13571), .A2(n8271), .ZN(n7627) );
  XNOR2_X1 U9726 ( .A(n12752), .B(n13601), .ZN(n12116) );
  AND2_X1 U9727 ( .A1(n9187), .A2(n9186), .ZN(n7628) );
  AND2_X1 U9728 ( .A1(n8928), .A2(n8927), .ZN(n7630) );
  OR2_X1 U9729 ( .A1(n9005), .A2(n9004), .ZN(P2_U3236) );
  AND2_X1 U9730 ( .A1(n9412), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7632) );
  INV_X1 U9731 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8761) );
  AND3_X1 U9732 ( .A1(n8471), .A2(n8470), .A3(n8469), .ZN(n7634) );
  AND4_X1 U9733 ( .A1(n9524), .A2(n9523), .A3(n9522), .A4(n9521), .ZN(n7635)
         );
  INV_X1 U9734 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U9735 ( .A1(n9355), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7636) );
  OR2_X1 U9736 ( .A1(n9425), .A2(n9463), .ZN(n7638) );
  NAND2_X1 U9737 ( .A1(n9409), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7639) );
  OR2_X1 U9738 ( .A1(n12585), .A2(n12584), .ZN(n7640) );
  AND2_X1 U9739 ( .A1(n9185), .A2(n9171), .ZN(n7641) );
  AND2_X1 U9740 ( .A1(n10444), .A2(n10443), .ZN(n7642) );
  INV_X1 U9741 ( .A(n9400), .ZN(n9397) );
  OR2_X1 U9742 ( .A1(n11192), .A2(n11191), .ZN(n7643) );
  INV_X1 U9743 ( .A(n11229), .ZN(n8991) );
  OR2_X1 U9744 ( .A1(n9046), .A2(n9045), .ZN(n7644) );
  OAI21_X1 U9745 ( .B1(n9025), .B2(n10143), .A(n9023), .ZN(n9028) );
  INV_X1 U9746 ( .A(n9104), .ZN(n9105) );
  NAND2_X1 U9747 ( .A1(n9106), .A2(n9105), .ZN(n9107) );
  OR2_X1 U9748 ( .A1(n9117), .A2(n9116), .ZN(n9118) );
  OAI21_X1 U9749 ( .B1(n14113), .B2(n9265), .A(n9137), .ZN(n9138) );
  INV_X1 U9750 ( .A(n13963), .ZN(n9205) );
  INV_X1 U9751 ( .A(n13079), .ZN(n12048) );
  AND2_X1 U9752 ( .A1(n9255), .A2(n9223), .ZN(n9224) );
  NAND2_X1 U9753 ( .A1(n7637), .A2(n12048), .ZN(n12049) );
  INV_X1 U9754 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7755) );
  INV_X1 U9755 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9312) );
  INV_X1 U9756 ( .A(n13207), .ZN(n8287) );
  NAND3_X1 U9757 ( .A1(n9419), .A2(n9407), .A3(n9312), .ZN(n9447) );
  INV_X1 U9758 ( .A(n8116), .ZN(n8115) );
  INV_X1 U9759 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U9760 ( .A1(n11664), .A2(n7041), .ZN(n11665) );
  OR2_X1 U9761 ( .A1(n8192), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8210) );
  OR2_X1 U9762 ( .A1(n8132), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8144) );
  OR2_X1 U9763 ( .A1(n13597), .A2(n13598), .ZN(n13595) );
  INV_X1 U9764 ( .A(n13168), .ZN(n13164) );
  INV_X1 U9765 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7759) );
  INV_X1 U9766 ( .A(n7928), .ZN(n7929) );
  INV_X1 U9767 ( .A(n8736), .ZN(n8352) );
  NAND2_X1 U9768 ( .A1(n14043), .A2(n8972), .ZN(n14024) );
  INV_X1 U9769 ( .A(n14205), .ZN(n8993) );
  XNOR2_X1 U9770 ( .A(n14591), .B(n12486), .ZN(n12519) );
  INV_X1 U9771 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11120) );
  AND2_X1 U9772 ( .A1(n11906), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11919) );
  INV_X1 U9773 ( .A(SI_12_), .ZN(n8417) );
  INV_X1 U9774 ( .A(n8087), .ZN(n8086) );
  INV_X1 U9775 ( .A(n15524), .ZN(n8254) );
  INV_X1 U9776 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n13351) );
  INV_X1 U9777 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7902) );
  AND3_X1 U9778 ( .A1(n8196), .A2(n8195), .A3(n8194), .ZN(n8197) );
  OR2_X1 U9779 ( .A1(n8144), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8157) );
  INV_X1 U9780 ( .A(n13741), .ZN(n8344) );
  INV_X1 U9781 ( .A(n12116), .ZN(n8005) );
  INV_X1 U9782 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7760) );
  OAI21_X1 U9783 ( .B1(n8168), .B2(n11721), .A(n8167), .ZN(n8171) );
  AND2_X1 U9784 ( .A1(n7945), .A2(n7930), .ZN(n7932) );
  OR2_X1 U9785 ( .A1(n8858), .A2(n8857), .ZN(n8885) );
  NAND2_X1 U9786 ( .A1(n8354), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U9787 ( .A1(n8352), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8746) );
  INV_X1 U9788 ( .A(n14179), .ZN(n8994) );
  INV_X1 U9789 ( .A(n14052), .ZN(n14064) );
  INV_X1 U9790 ( .A(n10809), .ZN(n10987) );
  OR2_X1 U9791 ( .A1(n12647), .A2(n12646), .ZN(n12648) );
  INV_X1 U9792 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11431) );
  AND2_X1 U9793 ( .A1(n11919), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11932) );
  INV_X1 U9794 ( .A(n11894), .ZN(n11895) );
  INV_X1 U9795 ( .A(n12309), .ZN(n10328) );
  OR2_X1 U9796 ( .A1(n8439), .A2(n10783), .ZN(n8440) );
  OR2_X1 U9797 ( .A1(n9670), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9671) );
  INV_X1 U9798 ( .A(n9520), .ZN(n10260) );
  INV_X1 U9799 ( .A(n12726), .ZN(n12279) );
  INV_X1 U9800 ( .A(n15474), .ZN(n10912) );
  NAND2_X1 U9801 ( .A1(n8156), .A2(n8155), .ZN(n8177) );
  NAND2_X1 U9802 ( .A1(n7984), .A2(n7983), .ZN(n7999) );
  INV_X1 U9803 ( .A(n12878), .ZN(n12867) );
  NAND2_X1 U9804 ( .A1(n12252), .A2(n12251), .ZN(n12744) );
  AND2_X1 U9805 ( .A1(n12035), .A2(n8242), .ZN(n13094) );
  INV_X1 U9806 ( .A(n13093), .ZN(n13090) );
  INV_X1 U9807 ( .A(n13211), .ZN(n13185) );
  INV_X1 U9808 ( .A(n12197), .ZN(n13194) );
  INV_X1 U9809 ( .A(n13582), .ZN(n13262) );
  INV_X1 U9810 ( .A(n12891), .ZN(n13600) );
  INV_X1 U9811 ( .A(n11402), .ZN(n12203) );
  OR2_X1 U9812 ( .A1(n13075), .A2(n13074), .ZN(n13615) );
  OR2_X1 U9813 ( .A1(n8205), .A2(n8127), .ZN(n8128) );
  INV_X1 U9814 ( .A(n10179), .ZN(n8081) );
  INV_X1 U9815 ( .A(n15515), .ZN(n15492) );
  AND2_X1 U9816 ( .A1(n12082), .A2(n12081), .ZN(n12202) );
  OR2_X1 U9817 ( .A1(n15504), .A2(n12236), .ZN(n13644) );
  INV_X1 U9818 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7770) );
  AND2_X1 U9819 ( .A1(n8057), .A2(n8040), .ZN(n8041) );
  AND2_X1 U9820 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n8350) );
  OR2_X1 U9821 ( .A1(n8769), .A2(n8768), .ZN(n8782) );
  OR2_X1 U9822 ( .A1(n8795), .A2(n13810), .ZN(n8820) );
  OR2_X1 U9823 ( .A1(n11212), .A2(n11211), .ZN(n11213) );
  NOR2_X1 U9824 ( .A1(n9930), .A2(n9920), .ZN(n9939) );
  AND2_X1 U9825 ( .A1(n8885), .A2(n8859), .ZN(n14011) );
  OR2_X1 U9826 ( .A1(n8721), .A2(n8720), .ZN(n8736) );
  INV_X1 U9827 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n13485) );
  INV_X1 U9828 ( .A(n15319), .ZN(n15281) );
  NAND2_X1 U9829 ( .A1(n8995), .A2(n8994), .ZN(n13967) );
  INV_X1 U9830 ( .A(n14082), .ZN(n8813) );
  INV_X1 U9831 ( .A(n14125), .ZN(n14145) );
  INV_X1 U9832 ( .A(n11629), .ZN(n8725) );
  NOR2_X1 U9833 ( .A1(n8654), .A2(n13485), .ZN(n8682) );
  INV_X1 U9834 ( .A(n15096), .ZN(n14025) );
  INV_X1 U9835 ( .A(n11795), .ZN(n9297) );
  OR3_X1 U9836 ( .A1(n14246), .A2(n14245), .A3(n14244), .ZN(n14291) );
  INV_X1 U9837 ( .A(n13905), .ZN(n11417) );
  NAND2_X1 U9838 ( .A1(n10142), .A2(n9928), .ZN(n15386) );
  AND2_X1 U9839 ( .A1(n15352), .A2(n9932), .ZN(n8929) );
  OR2_X1 U9840 ( .A1(n8650), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8665) );
  OR2_X1 U9841 ( .A1(n11849), .A2(n11848), .ZN(n11861) );
  OR2_X1 U9842 ( .A1(n9823), .A2(n12528), .ZN(n14410) );
  INV_X1 U9843 ( .A(n14438), .ZN(n14449) );
  OR2_X1 U9844 ( .A1(n12474), .A2(n12473), .ZN(n12475) );
  AND2_X1 U9845 ( .A1(n11823), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11834) );
  INV_X1 U9846 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14509) );
  INV_X1 U9847 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9638) );
  INV_X1 U9848 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n11143) );
  INV_X1 U9849 ( .A(n12507), .ZN(n14821) );
  OR2_X1 U9850 ( .A1(n14607), .A2(n14768), .ZN(n14783) );
  OR2_X1 U9851 ( .A1(n15034), .A2(n12522), .ZN(n10822) );
  INV_X1 U9852 ( .A(n12501), .ZN(n11155) );
  INV_X1 U9853 ( .A(n12500), .ZN(n11116) );
  INV_X1 U9854 ( .A(n14888), .ZN(n14828) );
  NAND2_X1 U9855 ( .A1(n14888), .A2(n14768), .ZN(n9829) );
  OAI21_X1 U9856 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n7677), .A(n7676), .ZN(
        n7690) );
  INV_X1 U9857 ( .A(n10786), .ZN(n10795) );
  AND2_X1 U9858 ( .A1(n10363), .A2(n15517), .ZN(n12878) );
  INV_X1 U9859 ( .A(n12885), .ZN(n12869) );
  INV_X1 U9860 ( .A(n13110), .ZN(n13133) );
  INV_X1 U9861 ( .A(n15406), .ZN(n15422) );
  INV_X1 U9862 ( .A(n13060), .ZN(n13073) );
  AND2_X1 U9863 ( .A1(n8305), .A2(n12183), .ZN(n15515) );
  AND2_X1 U9864 ( .A1(n15530), .A2(n15521), .ZN(n15071) );
  AND2_X1 U9865 ( .A1(n15530), .A2(n15505), .ZN(n15444) );
  INV_X1 U9866 ( .A(n15508), .ZN(n15525) );
  AND2_X1 U9867 ( .A1(n9013), .A2(n9012), .ZN(n10487) );
  INV_X1 U9868 ( .A(n15559), .ZN(n15523) );
  OR2_X1 U9869 ( .A1(n15502), .A2(n15579), .ZN(n15569) );
  INV_X1 U9870 ( .A(n13644), .ZN(n15579) );
  AND2_X1 U9871 ( .A1(n8317), .A2(n8316), .ZN(n10482) );
  INV_X1 U9872 ( .A(n12058), .ZN(n12236) );
  INV_X1 U9873 ( .A(n15111), .ZN(n13855) );
  OR2_X1 U9874 ( .A1(n13983), .A2(n8887), .ZN(n8894) );
  INV_X1 U9875 ( .A(n8738), .ZN(n8891) );
  INV_X1 U9876 ( .A(n8871), .ZN(n8887) );
  AND2_X1 U9877 ( .A1(n9441), .A2(n9440), .ZN(n15300) );
  OAI21_X1 U9878 ( .B1(n9934), .B2(n9428), .A(n9427), .ZN(n9441) );
  INV_X1 U9879 ( .A(n14137), .ZN(n15337) );
  INV_X1 U9880 ( .A(n14261), .ZN(n15372) );
  INV_X1 U9881 ( .A(n10605), .ZN(n15390) );
  AND2_X1 U9882 ( .A1(n9933), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9308) );
  INV_X1 U9883 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8913) );
  OR2_X1 U9884 ( .A1(n8665), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n8694) );
  AND2_X1 U9885 ( .A1(n9820), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9396) );
  NAND2_X1 U9886 ( .A1(n10028), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14441) );
  INV_X1 U9887 ( .A(n14441), .ZN(n14454) );
  AND4_X1 U9888 ( .A1(n11887), .A2(n11886), .A3(n11885), .A4(n11884), .ZN(
        n14351) );
  INV_X1 U9889 ( .A(n15208), .ZN(n14565) );
  INV_X1 U9890 ( .A(n15210), .ZN(n14576) );
  INV_X1 U9891 ( .A(n12515), .ZN(n14677) );
  INV_X1 U9892 ( .A(n14783), .ZN(n14835) );
  INV_X2 U9893 ( .A(n14855), .ZN(n14840) );
  INV_X1 U9894 ( .A(n14831), .ZN(n14858) );
  INV_X1 U9895 ( .A(n14939), .ZN(n15228) );
  INV_X1 U9896 ( .A(n15229), .ZN(n15256) );
  NAND2_X1 U9897 ( .A1(n9797), .A2(n9396), .ZN(n9830) );
  OR2_X1 U9898 ( .A1(n10494), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n11021) );
  AND2_X1 U9899 ( .A1(n10191), .A2(n10190), .ZN(n15417) );
  INV_X1 U9900 ( .A(n12882), .ZN(n11604) );
  NAND2_X1 U9901 ( .A1(n9974), .A2(n9973), .ZN(n12872) );
  NAND2_X1 U9902 ( .A1(n8216), .A2(n8215), .ZN(n12888) );
  INV_X1 U9903 ( .A(n15417), .ZN(n15414) );
  INV_X1 U9904 ( .A(n15425), .ZN(n15408) );
  NAND2_X1 U9905 ( .A1(n10183), .A2(n6587), .ZN(n15407) );
  INV_X1 U9906 ( .A(n15071), .ZN(n13606) );
  AND2_X1 U9907 ( .A1(n11408), .A2(n11407), .ZN(n15574) );
  AND2_X1 U9908 ( .A1(n10718), .A2(n10717), .ZN(n15550) );
  AOI21_X1 U9909 ( .B1(n8343), .B2(n13614), .A(n9016), .ZN(n9017) );
  NAND2_X1 U9910 ( .A1(n15603), .A2(n15523), .ZN(n13689) );
  INV_X1 U9911 ( .A(n15603), .ZN(n15600) );
  INV_X1 U9912 ( .A(n15582), .ZN(n8348) );
  INV_X1 U9913 ( .A(n12271), .ZN(n13725) );
  AND2_X1 U9914 ( .A1(n15550), .A2(n15549), .ZN(n15590) );
  AND2_X2 U9915 ( .A1(n8342), .A2(n9973), .ZN(n15582) );
  INV_X1 U9916 ( .A(n7765), .ZN(n13754) );
  INV_X1 U9917 ( .A(SI_14_), .ZN(n9707) );
  INV_X1 U9918 ( .A(n13749), .ZN(n13756) );
  NAND2_X1 U9919 ( .A1(n9993), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15111) );
  NAND2_X1 U9920 ( .A1(n8894), .A2(n8893), .ZN(n13892) );
  OR2_X1 U9921 ( .A1(n8703), .A2(n8702), .ZN(n13903) );
  INV_X1 U9922 ( .A(n15300), .ZN(n15311) );
  INV_X1 U9923 ( .A(n6581), .ZN(n14152) );
  OR2_X1 U9924 ( .A1(n8990), .A2(n8939), .ZN(n14137) );
  INV_X1 U9925 ( .A(n14163), .ZN(n15331) );
  OR3_X1 U9926 ( .A1(n14242), .A2(n14241), .A3(n14240), .ZN(n14290) );
  INV_X1 U9927 ( .A(n15393), .ZN(n15391) );
  NOR2_X1 U9928 ( .A1(n15349), .A2(n15340), .ZN(n15345) );
  INV_X1 U9929 ( .A(n15345), .ZN(n15346) );
  INV_X1 U9930 ( .A(n6585), .ZN(n11264) );
  INV_X1 U9931 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9897) );
  NAND2_X1 U9932 ( .A1(n9790), .A2(n9789), .ZN(n14456) );
  OR2_X1 U9933 ( .A1(n11437), .A2(n11436), .ZN(n14463) );
  CLKBUF_X2 U9934 ( .A(P1_U4016), .Z(n14496) );
  OR2_X1 U9935 ( .A1(n15201), .A2(n9566), .ZN(n15210) );
  OR2_X1 U9936 ( .A1(n15201), .A2(n14494), .ZN(n15212) );
  NAND2_X1 U9937 ( .A1(n14840), .A2(n10830), .ZN(n14838) );
  NAND2_X1 U9938 ( .A1(n15264), .A2(n14966), .ZN(n14963) );
  NAND2_X1 U9939 ( .A1(n15259), .A2(n14966), .ZN(n15011) );
  OR2_X1 U9940 ( .A1(n9967), .A2(n10817), .ZN(n15257) );
  OR2_X1 U9941 ( .A1(n9830), .A2(n9399), .ZN(n15224) );
  INV_X1 U9942 ( .A(n9404), .ZN(n11725) );
  INV_X1 U9943 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11100) );
  INV_X1 U9944 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9894) );
  INV_X1 U9945 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9409) );
  INV_X1 U9946 ( .A(n12897), .ZN(P3_U3897) );
  OAI21_X1 U9947 ( .B1(n9018), .B2(n8348), .A(n7621), .ZN(P3_U3456) );
  NOR2_X1 U9948 ( .A1(n9797), .A2(n9403), .ZN(P1_U4016) );
  INV_X1 U9949 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7679) );
  INV_X1 U9950 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n12970) );
  INV_X1 U9951 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15217) );
  NOR2_X1 U9952 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15217), .ZN(n7678) );
  INV_X1 U9953 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7677) );
  XNOR2_X1 U9954 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n7677), .ZN(n7692) );
  INV_X1 U9955 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n7675) );
  INV_X1 U9956 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n7672) );
  XNOR2_X1 U9957 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(P3_ADDR_REG_12__SCAN_IN), 
        .ZN(n7695) );
  INV_X1 U9958 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n7670) );
  XNOR2_X1 U9959 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7697) );
  INV_X1 U9960 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n7665) );
  XNOR2_X1 U9961 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7700) );
  INV_X1 U9962 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n7663) );
  XNOR2_X1 U9963 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7702) );
  INV_X1 U9964 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n7657) );
  XNOR2_X1 U9965 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n7722) );
  NAND2_X1 U9966 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n7647), .ZN(n7648) );
  NAND2_X1 U9967 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n7649), .ZN(n7652) );
  INV_X1 U9968 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7650) );
  NAND2_X1 U9969 ( .A1(n7704), .A2(n7650), .ZN(n7651) );
  NAND2_X1 U9970 ( .A1(n7652), .A2(n7651), .ZN(n7653) );
  NAND2_X1 U9971 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n7653), .ZN(n7655) );
  INV_X1 U9972 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U9973 ( .A1(n7718), .A2(n9683), .ZN(n7654) );
  NAND2_X1 U9974 ( .A1(n7655), .A2(n7654), .ZN(n7723) );
  NAND2_X1 U9975 ( .A1(n7722), .A2(n7723), .ZN(n7656) );
  NAND2_X1 U9976 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n7658), .ZN(n7661) );
  XOR2_X1 U9977 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n7658), .Z(n7729) );
  INV_X1 U9978 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7659) );
  NAND2_X1 U9979 ( .A1(n7729), .A2(n7659), .ZN(n7660) );
  NAND2_X1 U9980 ( .A1(n7661), .A2(n7660), .ZN(n7703) );
  NAND2_X1 U9981 ( .A1(n7702), .A2(n7703), .ZN(n7662) );
  NAND2_X1 U9982 ( .A1(n7700), .A2(n7701), .ZN(n7664) );
  NAND2_X1 U9983 ( .A1(n9638), .A2(n7666), .ZN(n7668) );
  XOR2_X1 U9984 ( .A(n9638), .B(n7666), .Z(n7699) );
  NAND2_X1 U9985 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n7699), .ZN(n7667) );
  NAND2_X1 U9986 ( .A1(n7668), .A2(n7667), .ZN(n7698) );
  NAND2_X1 U9987 ( .A1(n7697), .A2(n7698), .ZN(n7669) );
  NAND2_X1 U9988 ( .A1(n7695), .A2(n7696), .ZN(n7671) );
  OAI21_X1 U9989 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n7672), .A(n7671), .ZN(
        n7673) );
  INV_X1 U9990 ( .A(n7673), .ZN(n7693) );
  AND2_X1 U9991 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n7675), .ZN(n7674) );
  OAI22_X1 U9992 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n12970), .B1(n7678), .B2(
        n7690), .ZN(n7680) );
  NOR2_X1 U9993 ( .A1(n7679), .A2(n7680), .ZN(n7682) );
  XOR2_X1 U9994 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n7680), .Z(n7739) );
  NOR2_X1 U9995 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n7739), .ZN(n7681) );
  NOR2_X1 U9996 ( .A1(n7682), .A2(n7681), .ZN(n7684) );
  INV_X1 U9997 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7683) );
  NAND2_X1 U9998 ( .A1(n7684), .A2(n7683), .ZN(n7686) );
  XNOR2_X1 U9999 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n7684), .ZN(n7688) );
  NAND2_X1 U10000 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n7688), .ZN(n7685) );
  NAND2_X1 U10001 ( .A1(n7686), .A2(n7685), .ZN(n7742) );
  INV_X1 U10002 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n13049) );
  NOR2_X1 U10003 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n13049), .ZN(n7687) );
  AOI21_X1 U10004 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n13049), .A(n7687), .ZN(
        n7743) );
  XOR2_X1 U10005 ( .A(n7742), .B(n7743), .Z(n15037) );
  XNOR2_X1 U10006 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n7688), .ZN(n7740) );
  XOR2_X1 U10007 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .Z(n7689) );
  XOR2_X1 U10008 ( .A(n7690), .B(n7689), .Z(n15190) );
  XNOR2_X1 U10009 ( .A(n7692), .B(n7691), .ZN(n15186) );
  XNOR2_X1 U10010 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7694) );
  XNOR2_X1 U10011 ( .A(n7694), .B(n7693), .ZN(n15181) );
  XOR2_X1 U10012 ( .A(n7696), .B(n7695), .Z(n7734) );
  XOR2_X1 U10013 ( .A(n7698), .B(n7697), .Z(n15174) );
  XOR2_X1 U10014 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n7699), .Z(n15055) );
  XOR2_X1 U10015 ( .A(n7701), .B(n7700), .Z(n7731) );
  XOR2_X1 U10016 ( .A(n7703), .B(n7702), .Z(n15048) );
  AND2_X1 U10017 ( .A1(n7716), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n7717) );
  XNOR2_X1 U10018 ( .A(n7705), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15616) );
  XOR2_X1 U10019 ( .A(n7707), .B(n7706), .Z(n15042) );
  INV_X1 U10020 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7712) );
  NOR2_X1 U10021 ( .A1(n7711), .A2(n7712), .ZN(n7713) );
  AOI21_X1 U10022 ( .B1(n15415), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n7709), .ZN(
        n15610) );
  INV_X1 U10023 ( .A(n15610), .ZN(n7710) );
  NAND2_X1 U10024 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n7710), .ZN(n15620) );
  NOR2_X1 U10025 ( .A1(n15620), .A2(n15619), .ZN(n15618) );
  NOR2_X1 U10026 ( .A1(n15042), .A2(n15041), .ZN(n7714) );
  NAND2_X1 U10027 ( .A1(n15042), .A2(n15041), .ZN(n15040) );
  NAND2_X1 U10028 ( .A1(n15616), .A2(n15615), .ZN(n7715) );
  NOR2_X1 U10029 ( .A1(n15616), .A2(n15615), .ZN(n15614) );
  XNOR2_X1 U10030 ( .A(P2_ADDR_REG_4__SCAN_IN), .B(n7716), .ZN(n15605) );
  NOR2_X1 U10031 ( .A1(n15606), .A2(n15605), .ZN(n15604) );
  XNOR2_X1 U10032 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n7718), .ZN(n7719) );
  NAND2_X1 U10033 ( .A1(n7720), .A2(n7719), .ZN(n7721) );
  INV_X1 U10034 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15608) );
  INV_X1 U10035 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7724) );
  NOR2_X1 U10036 ( .A1(n7725), .A2(n7724), .ZN(n7726) );
  XOR2_X1 U10037 ( .A(n7723), .B(n7722), .Z(n15046) );
  INV_X1 U10038 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7728) );
  NAND2_X1 U10039 ( .A1(n7727), .A2(n7728), .ZN(n7730) );
  XNOR2_X1 U10040 ( .A(n7729), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15612) );
  NAND2_X1 U10041 ( .A1(n15613), .A2(n15612), .ZN(n15611) );
  NAND2_X1 U10042 ( .A1(n7731), .A2(n7732), .ZN(n7733) );
  INV_X1 U10043 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n15052) );
  NAND2_X1 U10044 ( .A1(n15055), .A2(n15056), .ZN(n15054) );
  NAND2_X1 U10045 ( .A1(n7734), .A2(n7735), .ZN(n7736) );
  INV_X1 U10046 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15178) );
  NAND2_X1 U10047 ( .A1(n7736), .A2(n15177), .ZN(n15182) );
  NOR2_X1 U10048 ( .A1(n15181), .A2(n15182), .ZN(n7737) );
  NAND2_X1 U10049 ( .A1(n15181), .A2(n15182), .ZN(n15180) );
  NAND2_X1 U10050 ( .A1(n15190), .A2(n15189), .ZN(n7738) );
  XNOR2_X1 U10051 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n7739), .ZN(n15194) );
  NAND2_X1 U10052 ( .A1(n15193), .A2(n15194), .ZN(n15192) );
  INV_X1 U10053 ( .A(n15059), .ZN(n15060) );
  INV_X1 U10054 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15062) );
  NAND2_X1 U10055 ( .A1(n7741), .A2(n7740), .ZN(n15061) );
  NAND2_X1 U10056 ( .A1(n15062), .A2(n15061), .ZN(n15058) );
  NAND2_X1 U10057 ( .A1(n15060), .A2(n15058), .ZN(n15036) );
  NAND2_X1 U10058 ( .A1(n7743), .A2(n7742), .ZN(n7744) );
  OAI21_X1 U10059 ( .B1(n13049), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n7744), .ZN(
        n7745) );
  XNOR2_X1 U10060 ( .A(n7745), .B(n13070), .ZN(n7746) );
  NAND4_X1 U10061 ( .A1(n8065), .A2(n8045), .A3(n8079), .A4(n7753), .ZN(n7754)
         );
  NAND2_X1 U10062 ( .A1(n7762), .A2(n7760), .ZN(n13747) );
  XNOR2_X2 U10063 ( .A(n7761), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7764) );
  NAND2_X1 U10064 ( .A1(n7831), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7769) );
  AND2_X4 U10065 ( .A1(n13754), .A2(n7764), .ZN(n7830) );
  NAND2_X1 U10066 ( .A1(n6608), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7768) );
  INV_X1 U10067 ( .A(n7764), .ZN(n12610) );
  AND2_X2 U10068 ( .A1(n12610), .A2(n7765), .ZN(n7834) );
  AND2_X2 U10069 ( .A1(n12610), .A2(n13754), .ZN(n7812) );
  XNOR2_X2 U10070 ( .A(n7771), .B(P3_IR_REG_27__SCAN_IN), .ZN(n8298) );
  INV_X1 U10071 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7773) );
  INV_X1 U10072 ( .A(SI_1_), .ZN(n9334) );
  OR2_X1 U10073 ( .A1(n8205), .A2(n9334), .ZN(n7777) );
  INV_X1 U10074 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8381) );
  XNOR2_X1 U10075 ( .A(n7790), .B(n7792), .ZN(n9333) );
  OAI211_X1 U10076 ( .C1(n10179), .C2(n10196), .A(n7777), .B(n7776), .ZN(
        n15524) );
  NAND2_X1 U10077 ( .A1(n7834), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7781) );
  NAND2_X1 U10078 ( .A1(n7812), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7780) );
  NAND2_X1 U10079 ( .A1(n7830), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7779) );
  NAND2_X1 U10080 ( .A1(n6606), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7778) );
  NAND4_X2 U10081 ( .A1(n7781), .A2(n7780), .A3(n7779), .A4(n7778), .ZN(n15516) );
  INV_X1 U10082 ( .A(SI_0_), .ZN(n9760) );
  OR2_X1 U10083 ( .A1(n8205), .A2(n9760), .ZN(n7785) );
  INV_X1 U10084 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U10085 ( .A1(n9761), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7782) );
  AND2_X1 U10086 ( .A1(n7790), .A2(n7782), .ZN(n9343) );
  OR2_X1 U10087 ( .A1(n7819), .A2(n9343), .ZN(n7784) );
  INV_X1 U10088 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10184) );
  OR2_X1 U10089 ( .A1(n10179), .A2(n10184), .ZN(n7783) );
  NOR2_X2 U10090 ( .A1(n15516), .A2(n10524), .ZN(n15520) );
  NAND2_X1 U10091 ( .A1(n10356), .A2(n12068), .ZN(n15491) );
  NAND2_X1 U10092 ( .A1(n6606), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U10093 ( .A1(n7830), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7788) );
  NAND2_X1 U10094 ( .A1(n7834), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U10095 ( .A1(n7812), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7786) );
  INV_X1 U10096 ( .A(n7790), .ZN(n7791) );
  NAND2_X1 U10097 ( .A1(n7792), .A2(n7791), .ZN(n7794) );
  XNOR2_X1 U10098 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7795) );
  OR2_X1 U10099 ( .A1(n7819), .A2(n9373), .ZN(n7797) );
  OR2_X1 U10100 ( .A1(n8205), .A2(SI_2_), .ZN(n7796) );
  OAI211_X1 U10101 ( .C1(n10252), .C2(n10179), .A(n7797), .B(n7796), .ZN(n7799) );
  INV_X1 U10102 ( .A(n7799), .ZN(n10533) );
  NAND2_X1 U10103 ( .A1(n7798), .A2(n7799), .ZN(n12054) );
  NAND2_X1 U10104 ( .A1(n12055), .A2(n12054), .ZN(n8255) );
  INV_X2 U10105 ( .A(n8255), .ZN(n12067) );
  NAND2_X1 U10106 ( .A1(n15491), .A2(n12067), .ZN(n15490) );
  NAND2_X1 U10107 ( .A1(n15490), .A2(n12055), .ZN(n15473) );
  NAND2_X1 U10108 ( .A1(n6607), .A2(n15484), .ZN(n7803) );
  NAND2_X1 U10109 ( .A1(n7830), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U10110 ( .A1(n8134), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7801) );
  NAND2_X1 U10111 ( .A1(n7812), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U10112 ( .A1(n7804), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7805) );
  OR2_X1 U10113 ( .A1(n8205), .A2(SI_3_), .ZN(n7810) );
  NAND2_X1 U10114 ( .A1(n9362), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7806) );
  XNOR2_X1 U10115 ( .A(n9367), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n7808) );
  XNOR2_X1 U10116 ( .A(n7820), .B(n7808), .ZN(n9381) );
  OAI211_X1 U10117 ( .C1(n7258), .C2(n10179), .A(n7810), .B(n7809), .ZN(n15483) );
  NAND2_X1 U10118 ( .A1(n12896), .A2(n15483), .ZN(n12071) );
  INV_X1 U10119 ( .A(n15477), .ZN(n12201) );
  NAND2_X1 U10120 ( .A1(n15473), .A2(n12201), .ZN(n7811) );
  NAND2_X1 U10121 ( .A1(n7811), .A2(n12070), .ZN(n10710) );
  INV_X1 U10122 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U10123 ( .A1(n7830), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7817) );
  AND2_X1 U10124 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7814) );
  NOR2_X1 U10125 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7832) );
  OR2_X1 U10126 ( .A1(n7814), .A2(n7832), .ZN(n10785) );
  NAND2_X1 U10127 ( .A1(n6606), .A2(n10785), .ZN(n7816) );
  NAND2_X1 U10128 ( .A1(n8134), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7815) );
  NAND4_X1 U10129 ( .A1(n7818), .A2(n7817), .A3(n7816), .A4(n7815), .ZN(n15474) );
  INV_X1 U10130 ( .A(n7820), .ZN(n7821) );
  NAND2_X1 U10131 ( .A1(n9367), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7822) );
  NAND2_X1 U10132 ( .A1(n9364), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7823) );
  NAND2_X1 U10133 ( .A1(n7843), .A2(n7823), .ZN(n7824) );
  NAND2_X1 U10134 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  AND2_X1 U10135 ( .A1(n7844), .A2(n7826), .ZN(n9375) );
  OR2_X1 U10136 ( .A1(n12040), .A2(SI_4_), .ZN(n7827) );
  OAI211_X1 U10137 ( .C1(n6753), .C2(n10179), .A(n7828), .B(n7827), .ZN(n10786) );
  NAND2_X1 U10138 ( .A1(n10912), .A2(n10795), .ZN(n12073) );
  NAND2_X1 U10139 ( .A1(n15474), .A2(n10786), .ZN(n12074) );
  NAND2_X1 U10140 ( .A1(n12073), .A2(n12074), .ZN(n8259) );
  NAND2_X1 U10141 ( .A1(n10710), .A2(n12204), .ZN(n7829) );
  NAND2_X1 U10142 ( .A1(n7829), .A2(n12073), .ZN(n10921) );
  NAND2_X1 U10143 ( .A1(n12030), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7838) );
  NAND2_X1 U10144 ( .A1(n7830), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U10145 ( .A1(n7832), .A2(n13440), .ZN(n7854) );
  OR2_X1 U10146 ( .A1(n13440), .A2(n7832), .ZN(n7833) );
  NAND2_X1 U10147 ( .A1(n7854), .A2(n7833), .ZN(n10926) );
  NAND2_X1 U10148 ( .A1(n6607), .A2(n10926), .ZN(n7836) );
  NAND2_X1 U10149 ( .A1(n8134), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7835) );
  NAND4_X1 U10150 ( .A1(n7838), .A2(n7837), .A3(n7836), .A4(n7835), .ZN(n15459) );
  NAND2_X1 U10151 ( .A1(n7840), .A2(n7839), .ZN(n7841) );
  NAND2_X1 U10152 ( .A1(n7841), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7842) );
  NAND2_X1 U10153 ( .A1(n9340), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U10154 ( .A1(n9365), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U10155 ( .A1(n7863), .A2(n7845), .ZN(n7847) );
  NAND2_X1 U10156 ( .A1(n7846), .A2(n7847), .ZN(n7850) );
  INV_X1 U10157 ( .A(n7846), .ZN(n7849) );
  INV_X1 U10158 ( .A(n7847), .ZN(n7848) );
  NAND2_X1 U10159 ( .A1(n7849), .A2(n7848), .ZN(n7864) );
  AND2_X1 U10160 ( .A1(n7850), .A2(n7864), .ZN(n9369) );
  OR2_X1 U10161 ( .A1(n12040), .A2(SI_5_), .ZN(n7851) );
  OAI211_X1 U10162 ( .C1(n10307), .C2(n6602), .A(n7852), .B(n7851), .ZN(n10925) );
  INV_X1 U10163 ( .A(n10925), .ZN(n10915) );
  NAND2_X1 U10164 ( .A1(n11035), .A2(n10915), .ZN(n12082) );
  NAND2_X1 U10165 ( .A1(n15459), .A2(n10925), .ZN(n12081) );
  NAND2_X1 U10166 ( .A1(n10921), .A2(n12202), .ZN(n7853) );
  NAND2_X1 U10167 ( .A1(n7853), .A2(n12082), .ZN(n15458) );
  NAND2_X1 U10168 ( .A1(n6583), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7859) );
  NAND2_X1 U10169 ( .A1(n7830), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U10170 ( .A1(n7854), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7855) );
  NAND2_X1 U10171 ( .A1(n7869), .A2(n7855), .ZN(n15470) );
  NAND2_X1 U10172 ( .A1(n6607), .A2(n15470), .ZN(n7857) );
  NAND2_X1 U10173 ( .A1(n8134), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7856) );
  NAND4_X1 U10174 ( .A1(n7859), .A2(n7858), .A3(n7857), .A4(n7856), .ZN(n12895) );
  NOR2_X1 U10175 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n7860) );
  NAND2_X1 U10176 ( .A1(n7861), .A2(n7860), .ZN(n7875) );
  NAND2_X1 U10177 ( .A1(n7875), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7862) );
  XNOR2_X1 U10178 ( .A(n7862), .B(P3_IR_REG_6__SCAN_IN), .ZN(n10451) );
  INV_X1 U10179 ( .A(SI_6_), .ZN(n9380) );
  OR2_X1 U10180 ( .A1(n12040), .A2(n9380), .ZN(n7866) );
  XNOR2_X1 U10181 ( .A(n7879), .B(n7877), .ZN(n9379) );
  OAI211_X1 U10182 ( .C1(n10179), .C2(n11093), .A(n7866), .B(n7865), .ZN(
        n11038) );
  NAND2_X1 U10183 ( .A1(n11173), .A2(n11038), .ZN(n12087) );
  INV_X1 U10184 ( .A(n11038), .ZN(n15469) );
  NAND2_X1 U10185 ( .A1(n12895), .A2(n15469), .ZN(n12088) );
  NAND2_X1 U10186 ( .A1(n12087), .A2(n12088), .ZN(n15464) );
  INV_X1 U10187 ( .A(n15464), .ZN(n12199) );
  NAND2_X1 U10188 ( .A1(n15458), .A2(n12199), .ZN(n7867) );
  NAND2_X1 U10189 ( .A1(n7867), .A2(n12087), .ZN(n11015) );
  NAND2_X1 U10190 ( .A1(n12030), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U10191 ( .A1(n7830), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7873) );
  AND2_X1 U10192 ( .A1(n7869), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7870) );
  OR2_X1 U10193 ( .A1(n7870), .A2(n7887), .ZN(n11166) );
  NAND2_X1 U10194 ( .A1(n6607), .A2(n11166), .ZN(n7872) );
  NAND2_X1 U10195 ( .A1(n8134), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7871) );
  NAND4_X1 U10196 ( .A1(n7874), .A2(n7873), .A3(n7872), .A4(n7871), .ZN(n15460) );
  NAND2_X1 U10197 ( .A1(n7893), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7876) );
  INV_X1 U10198 ( .A(n7877), .ZN(n7878) );
  NAND2_X1 U10199 ( .A1(n9386), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U10200 ( .A1(n9387), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n7880) );
  NAND2_X1 U10201 ( .A1(n7897), .A2(n7880), .ZN(n7881) );
  NAND2_X1 U10202 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  AND2_X1 U10203 ( .A1(n7898), .A2(n7883), .ZN(n9371) );
  OR2_X1 U10204 ( .A1(n12040), .A2(SI_7_), .ZN(n7884) );
  OAI211_X1 U10205 ( .C1(n11251), .C2(n10179), .A(n7885), .B(n7884), .ZN(
        n15560) );
  XNOR2_X1 U10206 ( .A(n15460), .B(n15560), .ZN(n11171) );
  INV_X1 U10207 ( .A(n15460), .ZN(n15451) );
  INV_X1 U10208 ( .A(n15560), .ZN(n11176) );
  NAND2_X1 U10209 ( .A1(n15451), .A2(n11176), .ZN(n12090) );
  NAND2_X1 U10210 ( .A1(n7830), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7892) );
  NAND2_X1 U10211 ( .A1(n12030), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7891) );
  NOR2_X1 U10212 ( .A1(n7887), .A2(n7886), .ZN(n7888) );
  OR2_X1 U10213 ( .A1(n7903), .A2(n7888), .ZN(n15454) );
  NAND2_X1 U10214 ( .A1(n6606), .A2(n15454), .ZN(n7890) );
  NAND2_X1 U10215 ( .A1(n8134), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7889) );
  NAND4_X1 U10216 ( .A1(n7892), .A2(n7891), .A3(n7890), .A4(n7889), .ZN(n12894) );
  OAI21_X1 U10217 ( .B1(n7893), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7894) );
  MUX2_X1 U10218 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7894), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n7896) );
  NAND2_X1 U10219 ( .A1(n7896), .A2(n7895), .ZN(n11254) );
  INV_X1 U10220 ( .A(SI_8_), .ZN(n9345) );
  OR2_X1 U10221 ( .A1(n12040), .A2(n9345), .ZN(n7901) );
  XNOR2_X1 U10222 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7899) );
  XNOR2_X1 U10223 ( .A(n7910), .B(n7899), .ZN(n9344) );
  OAI211_X1 U10224 ( .C1(n10179), .C2(n11254), .A(n7901), .B(n7900), .ZN(
        n15453) );
  INV_X1 U10225 ( .A(n15453), .ZN(n8265) );
  NAND2_X1 U10226 ( .A1(n12894), .A2(n8265), .ZN(n12096) );
  INV_X1 U10227 ( .A(n12894), .ZN(n11544) );
  NAND2_X1 U10228 ( .A1(n11544), .A2(n15453), .ZN(n12095) );
  NAND2_X1 U10229 ( .A1(n12030), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7908) );
  NAND2_X1 U10230 ( .A1(n7830), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7907) );
  OR2_X1 U10231 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  NAND2_X1 U10232 ( .A1(n7917), .A2(n7904), .ZN(n11549) );
  NAND2_X1 U10233 ( .A1(n6606), .A2(n11549), .ZN(n7906) );
  NAND2_X1 U10234 ( .A1(n8134), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7905) );
  NAND4_X1 U10235 ( .A1(n7908), .A2(n7907), .A3(n7906), .A4(n7905), .ZN(n12893) );
  NAND2_X1 U10236 ( .A1(n7895), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7909) );
  XNOR2_X1 U10237 ( .A(n7909), .B(n7166), .ZN(n11259) );
  INV_X1 U10238 ( .A(n11259), .ZN(n11374) );
  OR2_X1 U10239 ( .A1(n8205), .A2(SI_9_), .ZN(n7915) );
  NAND2_X1 U10240 ( .A1(n9391), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7911) );
  XNOR2_X1 U10241 ( .A(n9412), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n7913) );
  XNOR2_X1 U10242 ( .A(n7928), .B(n7913), .ZN(n9377) );
  OAI211_X1 U10243 ( .C1(n11374), .C2(n6602), .A(n7915), .B(n7914), .ZN(n11536) );
  INV_X1 U10244 ( .A(n11536), .ZN(n11548) );
  NAND2_X1 U10245 ( .A1(n15452), .A2(n11548), .ZN(n12099) );
  NAND2_X1 U10246 ( .A1(n12893), .A2(n11536), .ZN(n12100) );
  NAND2_X1 U10247 ( .A1(n12099), .A2(n12100), .ZN(n11402) );
  NAND2_X1 U10248 ( .A1(n11400), .A2(n12203), .ZN(n7916) );
  NAND2_X1 U10249 ( .A1(n7916), .A2(n12099), .ZN(n15434) );
  NAND2_X1 U10250 ( .A1(n7830), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7922) );
  NAND2_X1 U10251 ( .A1(n8134), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U10252 ( .A1(n12030), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U10253 ( .A1(n7917), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7918) );
  NAND2_X1 U10254 ( .A1(n7938), .A2(n7918), .ZN(n15442) );
  NAND2_X1 U10255 ( .A1(n6607), .A2(n15442), .ZN(n7919) );
  NAND4_X1 U10256 ( .A1(n7922), .A2(n7921), .A3(n7920), .A4(n7919), .ZN(n12892) );
  NOR2_X1 U10257 ( .A1(n6645), .A2(n7976), .ZN(n7923) );
  MUX2_X1 U10258 ( .A(n7976), .B(n7923), .S(P3_IR_REG_10__SCAN_IN), .Z(n7924)
         );
  INV_X1 U10259 ( .A(n7924), .ZN(n7927) );
  INV_X1 U10260 ( .A(n7925), .ZN(n7926) );
  NAND2_X1 U10261 ( .A1(n7927), .A2(n7926), .ZN(n11670) );
  INV_X1 U10262 ( .A(n11670), .ZN(n11383) );
  OR2_X1 U10263 ( .A1(n12040), .A2(SI_10_), .ZN(n7937) );
  NAND2_X1 U10264 ( .A1(n9424), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U10265 ( .A1(n9418), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n7930) );
  INV_X1 U10266 ( .A(n7931), .ZN(n7934) );
  INV_X1 U10267 ( .A(n7932), .ZN(n7933) );
  NAND2_X1 U10268 ( .A1(n7934), .A2(n7933), .ZN(n7935) );
  AND2_X1 U10269 ( .A1(n7946), .A2(n7935), .ZN(n9394) );
  OAI211_X1 U10270 ( .C1(n11383), .C2(n10179), .A(n7937), .B(n7936), .ZN(
        n15443) );
  INV_X1 U10271 ( .A(n15443), .ZN(n11601) );
  XNOR2_X1 U10272 ( .A(n12892), .B(n11601), .ZN(n15439) );
  INV_X1 U10273 ( .A(n12892), .ZN(n11545) );
  NAND2_X1 U10274 ( .A1(n11545), .A2(n11601), .ZN(n12103) );
  NAND2_X1 U10275 ( .A1(n7830), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U10276 ( .A1(n12030), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7942) );
  INV_X1 U10277 ( .A(n7949), .ZN(n7950) );
  NAND2_X1 U10278 ( .A1(n7938), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7939) );
  NAND2_X1 U10279 ( .A1(n7950), .A2(n7939), .ZN(n12846) );
  NAND2_X1 U10280 ( .A1(n6607), .A2(n12846), .ZN(n7941) );
  NAND2_X1 U10281 ( .A1(n12029), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7940) );
  OR2_X1 U10282 ( .A1(n7925), .A2(n7976), .ZN(n7944) );
  XNOR2_X1 U10283 ( .A(n7944), .B(n7963), .ZN(n11764) );
  XNOR2_X1 U10284 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n7956) );
  XNOR2_X1 U10285 ( .A(n7958), .B(n7956), .ZN(n9393) );
  OR2_X1 U10286 ( .A1(n12040), .A2(n13401), .ZN(n7947) );
  OAI211_X1 U10287 ( .C1(n10179), .C2(n11764), .A(n7948), .B(n7947), .ZN(
        n15085) );
  INV_X1 U10288 ( .A(n15085), .ZN(n11584) );
  XNOR2_X1 U10289 ( .A(n15435), .B(n11584), .ZN(n12208) );
  NAND2_X1 U10290 ( .A1(n15435), .A2(n15085), .ZN(n12107) );
  NAND2_X1 U10291 ( .A1(n7949), .A2(n13347), .ZN(n7985) );
  NAND2_X1 U10292 ( .A1(n7950), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U10293 ( .A1(n7985), .A2(n7951), .ZN(n15067) );
  NAND2_X1 U10294 ( .A1(n6606), .A2(n15067), .ZN(n7955) );
  NAND2_X1 U10295 ( .A1(n7830), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7954) );
  NAND2_X1 U10296 ( .A1(n8134), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7953) );
  NAND2_X1 U10297 ( .A1(n12030), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7952) );
  NAND4_X1 U10298 ( .A1(n7955), .A2(n7954), .A3(n7953), .A4(n7952), .ZN(n12891) );
  INV_X1 U10299 ( .A(n7956), .ZN(n7957) );
  NAND2_X1 U10300 ( .A1(n13505), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U10301 ( .A1(n9673), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7959) );
  NAND2_X1 U10302 ( .A1(n7969), .A2(n7959), .ZN(n7960) );
  NAND2_X1 U10303 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  AND2_X1 U10304 ( .A1(n7970), .A2(n7962), .ZN(n9415) );
  NAND2_X1 U10305 ( .A1(n9415), .A2(n12039), .ZN(n7967) );
  NAND2_X1 U10306 ( .A1(n7925), .A2(n7963), .ZN(n7975) );
  NAND2_X1 U10307 ( .A1(n7975), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7965) );
  INV_X1 U10308 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7964) );
  XNOR2_X1 U10309 ( .A(n7965), .B(n7964), .ZN(n12898) );
  INV_X1 U10310 ( .A(n12898), .ZN(n11770) );
  AOI22_X1 U10311 ( .A1(n8082), .A2(SI_12_), .B1(n8081), .B2(n11770), .ZN(
        n7966) );
  NAND2_X1 U10312 ( .A1(n7967), .A2(n7966), .ZN(n12791) );
  NAND2_X1 U10313 ( .A1(n13600), .A2(n12791), .ZN(n12112) );
  INV_X1 U10314 ( .A(n12791), .ZN(n15070) );
  NAND2_X1 U10315 ( .A1(n15070), .A2(n12891), .ZN(n12110) );
  NAND2_X1 U10316 ( .A1(n12112), .A2(n12110), .ZN(n13571) );
  NAND2_X1 U10317 ( .A1(n15069), .A2(n15068), .ZN(n7968) );
  NAND2_X1 U10318 ( .A1(n7973), .A2(n9713), .ZN(n7974) );
  NAND2_X1 U10319 ( .A1(n7992), .A2(n7974), .ZN(n9579) );
  NAND2_X1 U10320 ( .A1(n9579), .A2(n12039), .ZN(n7982) );
  NOR2_X1 U10321 ( .A1(n7975), .A2(P3_IR_REG_12__SCAN_IN), .ZN(n7979) );
  OR2_X1 U10322 ( .A1(n7979), .A2(n7976), .ZN(n7977) );
  INV_X1 U10323 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7978) );
  MUX2_X1 U10324 ( .A(n7977), .B(P3_IR_REG_31__SCAN_IN), .S(n7978), .Z(n7980)
         );
  NAND2_X1 U10325 ( .A1(n7979), .A2(n7978), .ZN(n7995) );
  NAND2_X1 U10326 ( .A1(n7980), .A2(n7995), .ZN(n12932) );
  AOI22_X1 U10327 ( .A1(n8082), .A2(n9578), .B1(n8081), .B2(n12932), .ZN(n7981) );
  NAND2_X1 U10328 ( .A1(n12030), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7990) );
  NAND2_X1 U10329 ( .A1(n7830), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7989) );
  INV_X1 U10330 ( .A(n7985), .ZN(n7984) );
  INV_X1 U10331 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7983) );
  NAND2_X1 U10332 ( .A1(n7985), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U10333 ( .A1(n7999), .A2(n7986), .ZN(n13602) );
  NAND2_X1 U10334 ( .A1(n6607), .A2(n13602), .ZN(n7988) );
  NAND2_X1 U10335 ( .A1(n8134), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7987) );
  OR2_X1 U10336 ( .A1(n13740), .A2(n15065), .ZN(n12117) );
  NAND2_X1 U10337 ( .A1(n13740), .A2(n15065), .ZN(n12118) );
  XNOR2_X1 U10338 ( .A(n9897), .B(P2_DATAO_REG_14__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U10339 ( .A1(n9706), .A2(n12039), .ZN(n7998) );
  NAND2_X1 U10340 ( .A1(n7995), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7994) );
  MUX2_X1 U10341 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7994), .S(
        P3_IR_REG_14__SCAN_IN), .Z(n7996) );
  NAND2_X1 U10342 ( .A1(n7996), .A2(n8028), .ZN(n12955) );
  INV_X1 U10343 ( .A(n12955), .ZN(n12947) );
  AOI22_X1 U10344 ( .A1(n8082), .A2(SI_14_), .B1(n8081), .B2(n12947), .ZN(
        n7997) );
  NAND2_X1 U10345 ( .A1(n7830), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8004) );
  NAND2_X1 U10346 ( .A1(n6583), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U10347 ( .A1(n7999), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10348 ( .A1(n8016), .A2(n8000), .ZN(n13588) );
  NAND2_X1 U10349 ( .A1(n6606), .A2(n13588), .ZN(n8002) );
  NAND2_X1 U10350 ( .A1(n8134), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8001) );
  NAND4_X1 U10351 ( .A1(n8004), .A2(n8003), .A3(n8002), .A4(n8001), .ZN(n12833) );
  NAND2_X1 U10352 ( .A1(n13586), .A2(n8005), .ZN(n13585) );
  NAND2_X1 U10353 ( .A1(n6828), .A2(n13601), .ZN(n12122) );
  NAND2_X1 U10354 ( .A1(n13585), .A2(n12122), .ZN(n13556) );
  NAND2_X1 U10355 ( .A1(n9897), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8006) );
  NAND2_X1 U10356 ( .A1(n9894), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8008) );
  XNOR2_X1 U10357 ( .A(n7248), .B(P2_DATAO_REG_15__SCAN_IN), .ZN(n8010) );
  XNOR2_X1 U10358 ( .A(n8023), .B(n8010), .ZN(n9882) );
  NAND2_X1 U10359 ( .A1(n9882), .A2(n12039), .ZN(n8013) );
  NAND2_X1 U10360 ( .A1(n8028), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8011) );
  XNOR2_X1 U10361 ( .A(n8011), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U10362 ( .A1(n8082), .A2(SI_15_), .B1(n8081), .B2(n12992), .ZN(
        n8012) );
  NAND2_X1 U10363 ( .A1(n12030), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U10364 ( .A1(n7830), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8020) );
  INV_X1 U10365 ( .A(n8016), .ZN(n8015) );
  INV_X1 U10366 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10367 ( .A1(n8016), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8017) );
  NAND2_X1 U10368 ( .A1(n8032), .A2(n8017), .ZN(n13561) );
  NAND2_X1 U10369 ( .A1(n6606), .A2(n13561), .ZN(n8019) );
  NAND2_X1 U10370 ( .A1(n12029), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8018) );
  NAND4_X1 U10371 ( .A1(n8021), .A2(n8020), .A3(n8019), .A4(n8018), .ZN(n13582) );
  OR2_X1 U10372 ( .A1(n13680), .A2(n13262), .ZN(n12125) );
  NAND2_X1 U10373 ( .A1(n13680), .A2(n13262), .ZN(n12130) );
  NAND2_X1 U10374 ( .A1(n10496), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U10375 ( .A1(n10529), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8024) );
  NAND2_X1 U10376 ( .A1(n8038), .A2(n8024), .ZN(n8025) );
  NAND2_X1 U10377 ( .A1(n8026), .A2(n8025), .ZN(n8027) );
  NAND2_X1 U10378 ( .A1(n8039), .A2(n8027), .ZN(n9887) );
  OAI21_X1 U10379 ( .B1(n8028), .B2(P3_IR_REG_15__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8029) );
  XNOR2_X1 U10380 ( .A(n8029), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U10381 ( .A1(n8082), .A2(SI_16_), .B1(n8081), .B2(n13011), .ZN(
        n8030) );
  NAND2_X1 U10382 ( .A1(n7830), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U10383 ( .A1(n12029), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8036) );
  NAND2_X1 U10384 ( .A1(n8032), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U10385 ( .A1(n8050), .A2(n8033), .ZN(n13264) );
  NAND2_X1 U10386 ( .A1(n6606), .A2(n13264), .ZN(n8035) );
  NAND2_X1 U10387 ( .A1(n12030), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8034) );
  NAND4_X1 U10388 ( .A1(n8037), .A2(n8036), .A3(n8035), .A4(n8034), .ZN(n13246) );
  XNOR2_X1 U10389 ( .A(n13676), .B(n13246), .ZN(n13259) );
  INV_X1 U10390 ( .A(n13246), .ZN(n13560) );
  NAND2_X1 U10391 ( .A1(n13676), .A2(n13560), .ZN(n12131) );
  INV_X1 U10392 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10540) );
  NAND2_X1 U10393 ( .A1(n10540), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8057) );
  INV_X1 U10394 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n13533) );
  NAND2_X1 U10395 ( .A1(n13533), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8040) );
  OR2_X1 U10396 ( .A1(n8042), .A2(n8041), .ZN(n8043) );
  NAND2_X1 U10397 ( .A1(n8058), .A2(n8043), .ZN(n10075) );
  NAND2_X1 U10398 ( .A1(n10075), .A2(n12039), .ZN(n8048) );
  INV_X1 U10399 ( .A(SI_17_), .ZN(n13366) );
  NAND2_X1 U10400 ( .A1(n8044), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8046) );
  XNOR2_X1 U10401 ( .A(n8046), .B(n8045), .ZN(n13020) );
  AOI22_X1 U10402 ( .A1(n8082), .A2(n13366), .B1(n8081), .B2(n13020), .ZN(
        n8047) );
  NAND2_X1 U10403 ( .A1(n7830), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8055) );
  NAND2_X1 U10404 ( .A1(n12029), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8054) );
  NAND2_X1 U10405 ( .A1(n8050), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8051) );
  NAND2_X1 U10406 ( .A1(n8069), .A2(n8051), .ZN(n13249) );
  NAND2_X1 U10407 ( .A1(n6606), .A2(n13249), .ZN(n8053) );
  NAND2_X1 U10408 ( .A1(n12030), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8052) );
  NAND4_X1 U10409 ( .A1(n8055), .A2(n8054), .A3(n8053), .A4(n8052), .ZN(n12890) );
  NAND2_X1 U10410 ( .A1(n13674), .A2(n12890), .ZN(n12136) );
  NAND2_X1 U10411 ( .A1(n12135), .A2(n12136), .ZN(n12214) );
  NAND2_X1 U10412 ( .A1(n13253), .A2(n13254), .ZN(n8056) );
  INV_X1 U10413 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n13404) );
  NAND2_X1 U10414 ( .A1(n13404), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8076) );
  INV_X1 U10415 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11025) );
  NAND2_X1 U10416 ( .A1(n11025), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8059) );
  OR2_X1 U10417 ( .A1(n8061), .A2(n8060), .ZN(n8062) );
  AND2_X1 U10418 ( .A1(n8077), .A2(n8062), .ZN(n10349) );
  NAND2_X1 U10419 ( .A1(n10349), .A2(n12039), .ZN(n8068) );
  NAND2_X1 U10420 ( .A1(n8064), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8063) );
  MUX2_X1 U10421 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8063), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n8066) );
  NAND2_X1 U10422 ( .A1(n8066), .A2(n8244), .ZN(n13054) );
  INV_X1 U10423 ( .A(n13054), .ZN(n13057) );
  AOI22_X1 U10424 ( .A1(n8082), .A2(SI_18_), .B1(n8081), .B2(n13057), .ZN(
        n8067) );
  NAND2_X1 U10425 ( .A1(n12030), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10426 ( .A1(n7830), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10427 ( .A1(n8069), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8070) );
  NAND2_X1 U10428 ( .A1(n8087), .A2(n8070), .ZN(n13236) );
  NAND2_X1 U10429 ( .A1(n6607), .A2(n13236), .ZN(n8072) );
  NAND2_X1 U10430 ( .A1(n12029), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8071) );
  NAND4_X1 U10431 ( .A1(n8074), .A2(n8073), .A3(n8072), .A4(n8071), .ZN(n13247) );
  INV_X1 U10432 ( .A(n13247), .ZN(n13222) );
  NAND2_X1 U10433 ( .A1(n13242), .A2(n13222), .ZN(n12142) );
  NAND2_X1 U10434 ( .A1(n11100), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8095) );
  INV_X1 U10435 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11102) );
  NAND2_X1 U10436 ( .A1(n11102), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8078) );
  XNOR2_X1 U10437 ( .A(n8094), .B(n8093), .ZN(n10426) );
  NAND2_X1 U10438 ( .A1(n10426), .A2(n12039), .ZN(n8084) );
  NAND2_X1 U10439 ( .A1(n8244), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8080) );
  AOI22_X1 U10440 ( .A1(n8082), .A2(n10425), .B1(n8081), .B2(n13060), .ZN(
        n8083) );
  NAND2_X1 U10441 ( .A1(n12030), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10442 ( .A1(n7830), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8091) );
  INV_X1 U10443 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8085) );
  NAND2_X1 U10444 ( .A1(n8087), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U10445 ( .A1(n8102), .A2(n8088), .ZN(n13225) );
  NAND2_X1 U10446 ( .A1(n6607), .A2(n13225), .ZN(n8090) );
  NAND2_X1 U10447 ( .A1(n12029), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8089) );
  NAND4_X1 U10448 ( .A1(n8092), .A2(n8091), .A3(n8090), .A4(n8089), .ZN(n13212) );
  OR2_X1 U10449 ( .A1(n13729), .A2(n13212), .ZN(n12147) );
  NAND2_X1 U10450 ( .A1(n8098), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U10451 ( .A1(n8110), .A2(n8099), .ZN(n10782) );
  INV_X1 U10452 ( .A(SI_20_), .ZN(n10783) );
  OR2_X1 U10453 ( .A1(n12040), .A2(n10783), .ZN(n8100) );
  NAND2_X1 U10454 ( .A1(n7830), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8107) );
  NAND2_X1 U10455 ( .A1(n12029), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8106) );
  NAND2_X1 U10456 ( .A1(n8102), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U10457 ( .A1(n8116), .A2(n8103), .ZN(n13215) );
  NAND2_X1 U10458 ( .A1(n6607), .A2(n13215), .ZN(n8105) );
  NAND2_X1 U10459 ( .A1(n12030), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8104) );
  NAND4_X1 U10460 ( .A1(n8107), .A2(n8106), .A3(n8105), .A4(n8104), .ZN(n12889) );
  XNOR2_X1 U10461 ( .A(n12271), .B(n12889), .ZN(n13207) );
  NAND2_X1 U10462 ( .A1(n13725), .A2(n12889), .ZN(n12151) );
  INV_X1 U10463 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11869) );
  NAND2_X1 U10464 ( .A1(n11869), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8125) );
  INV_X1 U10465 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11266) );
  NAND2_X1 U10466 ( .A1(n11266), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8111) );
  NAND2_X1 U10467 ( .A1(n8125), .A2(n8111), .ZN(n8122) );
  XNOR2_X1 U10468 ( .A(n8124), .B(n8122), .ZN(n11026) );
  NAND2_X1 U10469 ( .A1(n11026), .A2(n12039), .ZN(n8113) );
  INV_X1 U10470 ( .A(SI_21_), .ZN(n11027) );
  OR2_X1 U10471 ( .A1(n12040), .A2(n11027), .ZN(n8112) );
  NAND2_X1 U10472 ( .A1(n12030), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n8121) );
  NAND2_X1 U10473 ( .A1(n7830), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8120) );
  INV_X1 U10474 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8114) );
  NAND2_X1 U10475 ( .A1(n8116), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U10476 ( .A1(n8132), .A2(n8117), .ZN(n13199) );
  NAND2_X1 U10477 ( .A1(n6606), .A2(n13199), .ZN(n8119) );
  NAND2_X1 U10478 ( .A1(n12029), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8118) );
  NAND4_X1 U10479 ( .A1(n8121), .A2(n8120), .A3(n8119), .A4(n8118), .ZN(n13211) );
  NAND2_X1 U10480 ( .A1(n13198), .A2(n13185), .ZN(n12156) );
  OR2_X1 U10481 ( .A1(n13185), .A2(n13198), .ZN(n12155) );
  INV_X1 U10482 ( .A(n8122), .ZN(n8123) );
  INV_X1 U10483 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n12605) );
  XNOR2_X1 U10484 ( .A(n12605), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8139) );
  XNOR2_X1 U10485 ( .A(n8140), .B(n8139), .ZN(n11042) );
  NAND2_X1 U10486 ( .A1(n11042), .A2(n12039), .ZN(n8129) );
  INV_X1 U10487 ( .A(SI_22_), .ZN(n8127) );
  NAND2_X1 U10488 ( .A1(n7830), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8131) );
  NAND2_X1 U10489 ( .A1(n12030), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8130) );
  AND2_X1 U10490 ( .A1(n8131), .A2(n8130), .ZN(n8137) );
  NAND2_X1 U10491 ( .A1(n8132), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8133) );
  NAND2_X1 U10492 ( .A1(n8144), .A2(n8133), .ZN(n13188) );
  NAND2_X1 U10493 ( .A1(n13188), .A2(n6607), .ZN(n8136) );
  NAND2_X1 U10494 ( .A1(n12029), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8135) );
  NAND2_X1 U10495 ( .A1(n13187), .A2(n13197), .ZN(n12159) );
  NAND2_X1 U10496 ( .A1(n8138), .A2(n12160), .ZN(n13145) );
  NAND2_X1 U10497 ( .A1(n12605), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8141) );
  XNOR2_X1 U10498 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8150) );
  XNOR2_X1 U10499 ( .A(n8151), .B(n8150), .ZN(n11208) );
  NAND2_X1 U10500 ( .A1(n11208), .A2(n12039), .ZN(n8143) );
  INV_X1 U10501 ( .A(SI_23_), .ZN(n11210) );
  OR2_X1 U10502 ( .A1(n12040), .A2(n11210), .ZN(n8142) );
  INV_X1 U10503 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n8148) );
  NAND2_X1 U10504 ( .A1(n8144), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8145) );
  NAND2_X1 U10505 ( .A1(n8157), .A2(n8145), .ZN(n13174) );
  NAND2_X1 U10506 ( .A1(n13174), .A2(n6606), .ZN(n8147) );
  AOI22_X1 U10507 ( .A1(n7830), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n12029), 
        .B2(P3_REG1_REG_23__SCAN_IN), .ZN(n8146) );
  NAND2_X1 U10508 ( .A1(n13175), .A2(n13186), .ZN(n8149) );
  NAND2_X1 U10509 ( .A1(n13148), .A2(n8149), .ZN(n13168) );
  INV_X1 U10510 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11578) );
  NAND2_X1 U10511 ( .A1(n8152), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8153) );
  XNOR2_X1 U10512 ( .A(n8168), .B(P1_DATAO_REG_24__SCAN_IN), .ZN(n11588) );
  INV_X1 U10513 ( .A(SI_24_), .ZN(n11590) );
  NOR2_X1 U10514 ( .A1(n12040), .A2(n11590), .ZN(n8154) );
  INV_X1 U10515 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n8161) );
  INV_X1 U10516 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U10517 ( .A1(n8157), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8158) );
  NAND2_X1 U10518 ( .A1(n8177), .A2(n8158), .ZN(n13159) );
  NAND2_X1 U10519 ( .A1(n13159), .A2(n6607), .ZN(n8160) );
  AOI22_X1 U10520 ( .A1(n7830), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n6583), .B2(
        P3_REG0_REG_24__SCAN_IN), .ZN(n8159) );
  NOR2_X1 U10521 ( .A1(n13640), .A2(n13171), .ZN(n12053) );
  INV_X1 U10522 ( .A(n12053), .ZN(n8163) );
  AND2_X1 U10523 ( .A1(n13164), .A2(n8163), .ZN(n8164) );
  NAND2_X1 U10524 ( .A1(n13145), .A2(n8164), .ZN(n8166) );
  XNOR2_X1 U10525 ( .A(n13640), .B(n13171), .ZN(n13154) );
  INV_X1 U10526 ( .A(n13154), .ZN(n13147) );
  OR2_X1 U10527 ( .A1(n12053), .A2(n13146), .ZN(n8165) );
  NAND2_X1 U10528 ( .A1(n8166), .A2(n8165), .ZN(n13132) );
  NAND2_X1 U10529 ( .A1(n13373), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8185) );
  INV_X1 U10530 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11723) );
  NAND2_X1 U10531 ( .A1(n11723), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8169) );
  AND2_X1 U10532 ( .A1(n8185), .A2(n8169), .ZN(n8170) );
  NAND2_X1 U10533 ( .A1(n8171), .A2(n8170), .ZN(n8186) );
  NAND2_X1 U10534 ( .A1(n11636), .A2(n12039), .ZN(n8174) );
  INV_X1 U10535 ( .A(SI_25_), .ZN(n13365) );
  OR2_X1 U10536 ( .A1(n12040), .A2(n13365), .ZN(n8173) );
  INV_X1 U10537 ( .A(n8177), .ZN(n8176) );
  INV_X1 U10538 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U10539 ( .A1(n8177), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8178) );
  NAND2_X1 U10540 ( .A1(n8192), .A2(n8178), .ZN(n13140) );
  NAND2_X1 U10541 ( .A1(n13140), .A2(n6606), .ZN(n8184) );
  INV_X1 U10542 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U10543 ( .A1(n12030), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8180) );
  NAND2_X1 U10544 ( .A1(n12029), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8179) );
  OAI211_X1 U10545 ( .C1(n6609), .C2(n8181), .A(n8180), .B(n8179), .ZN(n8182)
         );
  INV_X1 U10546 ( .A(n8182), .ZN(n8183) );
  NAND2_X1 U10547 ( .A1(n13711), .A2(n13152), .ZN(n12171) );
  INV_X1 U10548 ( .A(n13711), .ZN(n12804) );
  OAI21_X2 U10549 ( .B1(n13132), .B2(n13135), .A(n12169), .ZN(n13128) );
  INV_X1 U10550 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n15028) );
  NAND2_X1 U10551 ( .A1(n15028), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8199) );
  INV_X1 U10552 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n14313) );
  NAND2_X1 U10553 ( .A1(n14313), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8187) );
  AND2_X1 U10554 ( .A1(n8199), .A2(n8187), .ZN(n8188) );
  NAND2_X1 U10555 ( .A1(n8189), .A2(n8188), .ZN(n8200) );
  OR2_X1 U10556 ( .A1(n12040), .A2(n13511), .ZN(n8191) );
  NAND2_X1 U10557 ( .A1(n8192), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8193) );
  NAND2_X1 U10558 ( .A1(n8210), .A2(n8193), .ZN(n13125) );
  NAND2_X1 U10559 ( .A1(n13125), .A2(n6607), .ZN(n8198) );
  NAND2_X1 U10560 ( .A1(n12029), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8196) );
  NAND2_X1 U10561 ( .A1(n7830), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10562 ( .A1(n6583), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U10563 ( .A1(n12870), .A2(n13110), .ZN(n12174) );
  NOR2_X2 U10564 ( .A1(n13128), .A2(n13127), .ZN(n13629) );
  INV_X1 U10565 ( .A(n13103), .ZN(n8217) );
  NAND2_X1 U10566 ( .A1(n8200), .A2(n8199), .ZN(n8203) );
  INV_X1 U10567 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15025) );
  NAND2_X1 U10568 ( .A1(n15025), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8218) );
  INV_X1 U10569 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n11774) );
  NAND2_X1 U10570 ( .A1(n11774), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8201) );
  AND2_X1 U10571 ( .A1(n8218), .A2(n8201), .ZN(n8202) );
  NAND2_X1 U10572 ( .A1(n8203), .A2(n8202), .ZN(n8219) );
  NAND2_X1 U10573 ( .A1(n8219), .A2(n8204), .ZN(n12611) );
  INV_X1 U10574 ( .A(n8210), .ZN(n8209) );
  INV_X1 U10575 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8208) );
  NAND2_X1 U10576 ( .A1(n8209), .A2(n8208), .ZN(n8224) );
  NAND2_X1 U10577 ( .A1(n8210), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8211) );
  NAND2_X1 U10578 ( .A1(n8224), .A2(n8211), .ZN(n13116) );
  NAND2_X1 U10579 ( .A1(n13116), .A2(n6607), .ZN(n8216) );
  NAND2_X1 U10580 ( .A1(n12029), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U10581 ( .A1(n7830), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U10582 ( .A1(n6583), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8212) );
  AND3_X1 U10583 ( .A1(n8214), .A2(n8213), .A3(n8212), .ZN(n8215) );
  NAND2_X1 U10584 ( .A1(n13703), .A2(n12888), .ZN(n12179) );
  NAND2_X1 U10585 ( .A1(n12741), .A2(n13123), .ZN(n12180) );
  NAND2_X1 U10586 ( .A1(n12179), .A2(n12180), .ZN(n13108) );
  INV_X1 U10587 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11999) );
  NAND2_X1 U10588 ( .A1(n11999), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8233) );
  INV_X1 U10589 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14310) );
  NAND2_X1 U10590 ( .A1(n14310), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8220) );
  NAND2_X1 U10591 ( .A1(n8233), .A2(n8220), .ZN(n8230) );
  XNOR2_X1 U10592 ( .A(n8232), .B(n8230), .ZN(n12533) );
  NAND2_X1 U10593 ( .A1(n12533), .A2(n12039), .ZN(n8222) );
  INV_X1 U10594 ( .A(SI_28_), .ZN(n12535) );
  OR2_X1 U10595 ( .A1(n12040), .A2(n12535), .ZN(n8221) );
  INV_X1 U10596 ( .A(n8224), .ZN(n8223) );
  NAND2_X1 U10597 ( .A1(n8223), .A2(n13534), .ZN(n13076) );
  NAND2_X1 U10598 ( .A1(n8224), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8225) );
  NAND2_X1 U10599 ( .A1(n13076), .A2(n8225), .ZN(n13097) );
  NAND2_X1 U10600 ( .A1(n12029), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8228) );
  NAND2_X1 U10601 ( .A1(n12030), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8227) );
  NAND2_X1 U10602 ( .A1(n7830), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8226) );
  NAND3_X1 U10603 ( .A1(n8228), .A2(n8227), .A3(n8226), .ZN(n8229) );
  INV_X1 U10604 ( .A(n8295), .ZN(n12187) );
  NAND2_X1 U10605 ( .A1(n13096), .A2(n13111), .ZN(n12181) );
  INV_X1 U10606 ( .A(n8230), .ZN(n8231) );
  NAND2_X1 U10607 ( .A1(n8232), .A2(n8231), .ZN(n8234) );
  INV_X1 U10608 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n12020) );
  XNOR2_X1 U10609 ( .A(n12020), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n8235) );
  XNOR2_X1 U10610 ( .A(n12022), .B(n8235), .ZN(n13752) );
  NAND2_X1 U10611 ( .A1(n13752), .A2(n12039), .ZN(n8237) );
  INV_X1 U10612 ( .A(SI_29_), .ZN(n13753) );
  OR2_X1 U10613 ( .A1(n12040), .A2(n13753), .ZN(n8236) );
  OR2_X1 U10614 ( .A1(n13076), .A2(n8238), .ZN(n12035) );
  NAND2_X1 U10615 ( .A1(n12029), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U10616 ( .A1(n12030), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U10617 ( .A1(n7830), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8239) );
  AND3_X1 U10618 ( .A1(n8241), .A2(n8240), .A3(n8239), .ZN(n8242) );
  NAND2_X1 U10619 ( .A1(n8343), .A2(n13094), .ZN(n12043) );
  NAND2_X1 U10620 ( .A1(n12186), .A2(n12043), .ZN(n12221) );
  INV_X1 U10621 ( .A(n12221), .ZN(n8243) );
  XNOR2_X1 U10622 ( .A(n12019), .B(n8243), .ZN(n13087) );
  NAND2_X1 U10623 ( .A1(n6685), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8247) );
  OAI21_X1 U10624 ( .B1(n8331), .B2(n12058), .A(n13073), .ZN(n8249) );
  NAND2_X1 U10625 ( .A1(n6698), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8248) );
  NAND2_X1 U10626 ( .A1(n8249), .A2(n12060), .ZN(n8251) );
  NAND2_X1 U10627 ( .A1(n10784), .A2(n12060), .ZN(n9007) );
  NAND2_X1 U10628 ( .A1(n9007), .A2(n12058), .ZN(n8250) );
  NAND2_X1 U10629 ( .A1(n8251), .A2(n8250), .ZN(n9980) );
  NOR2_X1 U10630 ( .A1(n12230), .A2(n15523), .ZN(n8252) );
  NAND2_X1 U10631 ( .A1(n9980), .A2(n8252), .ZN(n8253) );
  AND2_X1 U10632 ( .A1(n13073), .A2(n12236), .ZN(n8332) );
  INV_X1 U10633 ( .A(n8332), .ZN(n8296) );
  NAND2_X1 U10634 ( .A1(n8296), .A2(n12230), .ZN(n9008) );
  OR2_X1 U10635 ( .A1(n9008), .A2(n12058), .ZN(n9006) );
  NAND2_X1 U10636 ( .A1(n10784), .A2(n13073), .ZN(n15504) );
  INV_X1 U10637 ( .A(n13111), .ZN(n10799) );
  INV_X1 U10638 ( .A(n10524), .ZN(n9978) );
  AND2_X1 U10639 ( .A1(n15516), .A2(n9978), .ZN(n10357) );
  NAND2_X1 U10640 ( .A1(n10359), .A2(n15512), .ZN(n15511) );
  NAND2_X1 U10641 ( .A1(n15493), .A2(n8254), .ZN(n15496) );
  NAND2_X1 U10642 ( .A1(n15511), .A2(n15496), .ZN(n8256) );
  NAND2_X1 U10643 ( .A1(n8256), .A2(n8255), .ZN(n15499) );
  NAND2_X1 U10644 ( .A1(n10629), .A2(n7799), .ZN(n15475) );
  NAND2_X1 U10645 ( .A1(n12896), .A2(n10631), .ZN(n10711) );
  NAND2_X1 U10646 ( .A1(n15474), .A2(n10795), .ZN(n8258) );
  AND2_X1 U10647 ( .A1(n10711), .A2(n8258), .ZN(n8257) );
  NAND2_X1 U10648 ( .A1(n15476), .A2(n8257), .ZN(n8262) );
  INV_X1 U10649 ( .A(n8258), .ZN(n8260) );
  OR2_X1 U10650 ( .A1(n8260), .A2(n8259), .ZN(n8261) );
  AND2_X1 U10651 ( .A1(n8262), .A2(n8261), .ZN(n10920) );
  NAND2_X1 U10652 ( .A1(n11035), .A2(n10925), .ZN(n15461) );
  AND2_X1 U10653 ( .A1(n15464), .A2(n15461), .ZN(n8263) );
  NAND2_X1 U10654 ( .A1(n12895), .A2(n11038), .ZN(n8264) );
  AND2_X1 U10655 ( .A1(n12894), .A2(n15453), .ZN(n8267) );
  NAND2_X1 U10656 ( .A1(n11544), .A2(n8265), .ZN(n8266) );
  NAND2_X1 U10657 ( .A1(n11401), .A2(n11402), .ZN(n8269) );
  NAND2_X1 U10658 ( .A1(n15452), .A2(n11536), .ZN(n8268) );
  NAND2_X1 U10659 ( .A1(n8269), .A2(n8268), .ZN(n15438) );
  NAND2_X1 U10660 ( .A1(n12892), .A2(n11601), .ZN(n8270) );
  NAND2_X1 U10661 ( .A1(n15435), .A2(n11584), .ZN(n13568) );
  NAND2_X1 U10662 ( .A1(n6828), .A2(n12833), .ZN(n8275) );
  NAND2_X1 U10663 ( .A1(n13740), .A2(n12830), .ZN(n13574) );
  NAND2_X1 U10664 ( .A1(n12891), .A2(n12791), .ZN(n13572) );
  INV_X1 U10665 ( .A(n8273), .ZN(n8277) );
  OR2_X1 U10666 ( .A1(n15435), .A2(n11584), .ZN(n13570) );
  AND2_X1 U10667 ( .A1(n13570), .A2(n8274), .ZN(n13576) );
  AND2_X1 U10668 ( .A1(n13576), .A2(n8275), .ZN(n8276) );
  AND2_X1 U10669 ( .A1(n13680), .A2(n13582), .ZN(n8278) );
  NOR2_X1 U10670 ( .A1(n13676), .A2(n13246), .ZN(n8280) );
  NAND2_X1 U10671 ( .A1(n13676), .A2(n13246), .ZN(n8279) );
  OR2_X1 U10672 ( .A1(n13674), .A2(n13263), .ZN(n8281) );
  INV_X1 U10673 ( .A(n13233), .ZN(n8282) );
  OR2_X1 U10674 ( .A1(n13242), .A2(n13247), .ZN(n8283) );
  INV_X1 U10675 ( .A(n13212), .ZN(n13235) );
  OR2_X1 U10676 ( .A1(n13729), .A2(n13235), .ZN(n8284) );
  NAND2_X1 U10677 ( .A1(n13220), .A2(n8284), .ZN(n8286) );
  NAND2_X1 U10678 ( .A1(n13729), .A2(n13235), .ZN(n8285) );
  NAND2_X1 U10679 ( .A1(n8286), .A2(n8285), .ZN(n13208) );
  INV_X1 U10680 ( .A(n13208), .ZN(n8288) );
  NAND2_X1 U10681 ( .A1(n8288), .A2(n8287), .ZN(n13210) );
  NAND2_X1 U10682 ( .A1(n12271), .A2(n12889), .ZN(n8289) );
  OR2_X1 U10683 ( .A1(n13198), .A2(n13211), .ZN(n8290) );
  NAND2_X1 U10684 ( .A1(n13198), .A2(n13211), .ZN(n8291) );
  NAND2_X1 U10685 ( .A1(n13175), .A2(n13151), .ZN(n8293) );
  NAND2_X1 U10686 ( .A1(n13167), .A2(n8293), .ZN(n13155) );
  INV_X1 U10687 ( .A(n13171), .ZN(n12725) );
  NAND2_X1 U10688 ( .A1(n13153), .A2(n7626), .ZN(n13136) );
  NAND2_X1 U10689 ( .A1(n13136), .A2(n13135), .ZN(n13134) );
  NAND2_X1 U10690 ( .A1(n13707), .A2(n13110), .ZN(n8294) );
  AOI22_X1 U10691 ( .A1(n13121), .A2(n8294), .B1(n13133), .B2(n12870), .ZN(
        n13109) );
  NAND2_X1 U10692 ( .A1(n13109), .A2(n13108), .ZN(n13107) );
  OAI21_X1 U10693 ( .B1(n12888), .B2(n12741), .A(n13107), .ZN(n13092) );
  NAND2_X1 U10694 ( .A1(n8331), .A2(n10352), .ZN(n12052) );
  INV_X1 U10695 ( .A(n8297), .ZN(n12232) );
  NAND2_X1 U10696 ( .A1(n12232), .A2(n10221), .ZN(n10197) );
  NAND2_X1 U10697 ( .A1(n10179), .A2(n10197), .ZN(n8304) );
  INV_X1 U10698 ( .A(P3_B_REG_SCAN_IN), .ZN(n8299) );
  OR2_X1 U10699 ( .A1(n8297), .A2(n8299), .ZN(n8300) );
  NAND2_X1 U10700 ( .A1(n15517), .A2(n8300), .ZN(n13074) );
  AOI22_X1 U10701 ( .A1(n7830), .A2(P3_REG2_REG_30__SCAN_IN), .B1(n12030), 
        .B2(P3_REG0_REG_30__SCAN_IN), .ZN(n8301) );
  INV_X1 U10702 ( .A(n8301), .ZN(n8303) );
  INV_X1 U10703 ( .A(n12035), .ZN(n8302) );
  AOI211_X1 U10704 ( .C1(n12029), .C2(P3_REG1_REG_30__SCAN_IN), .A(n8303), .B(
        n8302), .ZN(n12047) );
  INV_X1 U10705 ( .A(n8304), .ZN(n8305) );
  INV_X1 U10706 ( .A(n9980), .ZN(n8335) );
  NAND2_X1 U10707 ( .A1(n8306), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8307) );
  INV_X1 U10708 ( .A(n8308), .ZN(n8310) );
  NAND2_X1 U10709 ( .A1(n8310), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8311) );
  MUX2_X1 U10710 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8311), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8313) );
  INV_X1 U10711 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n13503) );
  INV_X1 U10712 ( .A(n8337), .ZN(n11718) );
  NAND2_X1 U10713 ( .A1(n11718), .A2(n11591), .ZN(n8314) );
  INV_X1 U10714 ( .A(n13743), .ZN(n8319) );
  INV_X1 U10715 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U10716 ( .A1(n9532), .A2(n9414), .ZN(n8317) );
  NAND2_X1 U10717 ( .A1(n11718), .A2(n11638), .ZN(n8316) );
  INV_X1 U10718 ( .A(n10482), .ZN(n8318) );
  NAND2_X1 U10719 ( .A1(n8319), .A2(n8318), .ZN(n9013) );
  NOR4_X1 U10720 ( .A1(P3_D_REG_23__SCAN_IN), .A2(P3_D_REG_15__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8328) );
  INV_X1 U10721 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n13391) );
  INV_X1 U10722 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n13474) );
  INV_X1 U10723 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n13473) );
  INV_X1 U10724 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n13512) );
  NAND4_X1 U10725 ( .A1(n13391), .A2(n13474), .A3(n13473), .A4(n13512), .ZN(
        n8325) );
  NOR4_X1 U10726 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n8323) );
  NOR4_X1 U10727 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n8322) );
  NOR4_X1 U10728 ( .A1(P3_D_REG_28__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8321) );
  NOR4_X1 U10729 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_30__SCAN_IN), .A4(P3_D_REG_13__SCAN_IN), .ZN(n8320) );
  NAND4_X1 U10730 ( .A1(n8323), .A2(n8322), .A3(n8321), .A4(n8320), .ZN(n8324)
         );
  NOR4_X1 U10731 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        n8325), .A4(n8324), .ZN(n8327) );
  NOR4_X1 U10732 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8326) );
  NAND3_X1 U10733 ( .A1(n8328), .A2(n8327), .A3(n8326), .ZN(n8329) );
  NAND2_X1 U10734 ( .A1(n9532), .A2(n8329), .ZN(n9011) );
  INV_X1 U10735 ( .A(n9011), .ZN(n8330) );
  NAND3_X1 U10736 ( .A1(n13743), .A2(n10482), .A3(n9011), .ZN(n9981) );
  OR2_X1 U10737 ( .A1(n12230), .A2(n12165), .ZN(n10152) );
  INV_X1 U10738 ( .A(n10152), .ZN(n8333) );
  AND2_X1 U10739 ( .A1(n12228), .A2(n8332), .ZN(n9979) );
  NOR2_X1 U10740 ( .A1(n8333), .A2(n9979), .ZN(n8334) );
  OAI22_X1 U10741 ( .A1(n8335), .A2(n9987), .B1(n9981), .B2(n8334), .ZN(n8342)
         );
  NOR2_X1 U10742 ( .A1(n11638), .A2(n11591), .ZN(n8336) );
  NAND2_X1 U10743 ( .A1(n8337), .A2(n8336), .ZN(n9984) );
  INV_X1 U10744 ( .A(n8338), .ZN(n8339) );
  NAND2_X1 U10745 ( .A1(n8339), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8340) );
  MUX2_X1 U10746 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8340), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n8341) );
  NAND2_X1 U10747 ( .A1(n8341), .A2(n8306), .ZN(n10180) );
  INV_X1 U10748 ( .A(n13742), .ZN(n9990) );
  INV_X1 U10749 ( .A(n10182), .ZN(n9973) );
  INV_X1 U10750 ( .A(n8343), .ZN(n13085) );
  NAND2_X1 U10751 ( .A1(n8343), .A2(n8344), .ZN(n8347) );
  INV_X1 U10752 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8345) );
  OR2_X1 U10753 ( .A1(n15582), .A2(n8345), .ZN(n8346) );
  NAND2_X1 U10754 ( .A1(n8577), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8592) );
  INV_X1 U10755 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U10756 ( .A1(n8610), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U10757 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n8349) );
  OR2_X1 U10758 ( .A1(n8638), .A2(n8349), .ZN(n8654) );
  NAND2_X1 U10759 ( .A1(n8682), .A2(n8350), .ZN(n8699) );
  INV_X1 U10760 ( .A(n8699), .ZN(n8351) );
  NAND2_X1 U10761 ( .A1(n8351), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8721) );
  INV_X1 U10762 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8720) );
  INV_X1 U10763 ( .A(n8746), .ZN(n8353) );
  NAND2_X1 U10764 ( .A1(n8353), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8769) );
  INV_X1 U10765 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8768) );
  INV_X1 U10766 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13810) );
  INV_X1 U10767 ( .A(n8820), .ZN(n8356) );
  AND2_X1 U10768 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n8355) );
  NAND2_X1 U10769 ( .A1(n8356), .A2(n8355), .ZN(n8833) );
  INV_X1 U10770 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13852) );
  INV_X1 U10771 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13821) );
  INV_X1 U10772 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8857) );
  INV_X1 U10773 ( .A(n8885), .ZN(n8358) );
  AND2_X1 U10774 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8357) );
  NAND2_X1 U10775 ( .A1(n8358), .A2(n8357), .ZN(n9001) );
  NOR2_X2 U10776 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n8545) );
  NOR2_X1 U10778 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n8368) );
  NOR2_X1 U10779 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8367) );
  NOR2_X1 U10780 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8366) );
  NAND4_X1 U10781 ( .A1(n8368), .A2(n8367), .A3(n8366), .A4(n8913), .ZN(n8369)
         );
  NAND2_X1 U10782 ( .A1(n8371), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8370) );
  OR2_X1 U10783 ( .A1(n9001), .A2(n8887), .ZN(n8379) );
  INV_X1 U10784 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8376) );
  AND2_X4 U10785 ( .A1(n12001), .A2(n11773), .ZN(n8536) );
  NAND2_X1 U10786 ( .A1(n8536), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8375) );
  INV_X2 U10787 ( .A(n8520), .ZN(n9201) );
  NAND2_X1 U10788 ( .A1(n9201), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8374) );
  OAI211_X1 U10789 ( .C1(n8376), .C2(n8891), .A(n8375), .B(n8374), .ZN(n8377)
         );
  INV_X1 U10790 ( .A(n8377), .ZN(n8378) );
  NAND2_X1 U10791 ( .A1(n8379), .A2(n8378), .ZN(n13891) );
  NAND2_X1 U10792 ( .A1(n8380), .A2(SI_1_), .ZN(n8384) );
  INV_X1 U10793 ( .A(n8476), .ZN(n8383) );
  MUX2_X1 U10794 ( .A(n9761), .B(n8381), .S(n8387), .Z(n8382) );
  NOR2_X1 U10795 ( .A1(n8382), .A2(n9760), .ZN(n8474) );
  NAND2_X1 U10796 ( .A1(n8383), .A2(n8474), .ZN(n8473) );
  OAI21_X1 U10797 ( .B1(n8385), .B2(SI_2_), .A(n8510), .ZN(n8499) );
  INV_X1 U10798 ( .A(n8499), .ZN(n8386) );
  NAND2_X1 U10799 ( .A1(n8498), .A2(n8386), .ZN(n8511) );
  MUX2_X1 U10800 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8387), .Z(n8390) );
  NAND2_X1 U10801 ( .A1(n8390), .A2(SI_3_), .ZN(n8389) );
  AND2_X1 U10802 ( .A1(n8510), .A2(n8389), .ZN(n8388) );
  NAND2_X1 U10803 ( .A1(n8511), .A2(n8388), .ZN(n8527) );
  INV_X1 U10804 ( .A(n8389), .ZN(n8392) );
  OAI21_X1 U10805 ( .B1(SI_3_), .B2(n8390), .A(n8389), .ZN(n8512) );
  INV_X1 U10806 ( .A(n8512), .ZN(n8391) );
  OR2_X1 U10807 ( .A1(n8392), .A2(n8391), .ZN(n8526) );
  OAI21_X1 U10808 ( .B1(n8393), .B2(SI_4_), .A(n8396), .ZN(n8528) );
  INV_X1 U10809 ( .A(n8528), .ZN(n8394) );
  AND2_X1 U10810 ( .A1(n8526), .A2(n8394), .ZN(n8395) );
  NAND2_X1 U10811 ( .A1(n8397), .A2(SI_5_), .ZN(n8399) );
  OAI21_X1 U10812 ( .B1(n8397), .B2(SI_5_), .A(n8399), .ZN(n8398) );
  INV_X1 U10813 ( .A(n8398), .ZN(n8541) );
  MUX2_X1 U10814 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n8387), .Z(n8400) );
  NAND2_X1 U10815 ( .A1(n8400), .A2(SI_6_), .ZN(n8402) );
  OAI21_X1 U10816 ( .B1(SI_6_), .B2(n8400), .A(n8402), .ZN(n8401) );
  MUX2_X1 U10817 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n7274), .Z(n8403) );
  NAND2_X1 U10818 ( .A1(n8403), .A2(SI_7_), .ZN(n8405) );
  OAI21_X1 U10819 ( .B1(n8403), .B2(SI_7_), .A(n8405), .ZN(n8404) );
  INV_X1 U10820 ( .A(n8404), .ZN(n8570) );
  MUX2_X1 U10821 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n7274), .Z(n8406) );
  NAND2_X1 U10822 ( .A1(n8406), .A2(SI_8_), .ZN(n8408) );
  OAI21_X1 U10823 ( .B1(SI_8_), .B2(n8406), .A(n8408), .ZN(n8407) );
  INV_X1 U10824 ( .A(n8407), .ZN(n8583) );
  NAND2_X1 U10825 ( .A1(n8584), .A2(n8583), .ZN(n8586) );
  OAI21_X1 U10826 ( .B1(n8409), .B2(SI_9_), .A(n8411), .ZN(n8410) );
  MUX2_X1 U10827 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n7274), .Z(n8412) );
  NAND2_X1 U10828 ( .A1(n8412), .A2(SI_10_), .ZN(n8414) );
  OAI21_X1 U10829 ( .B1(n8412), .B2(SI_10_), .A(n8414), .ZN(n8617) );
  INV_X1 U10830 ( .A(n8617), .ZN(n8413) );
  XNOR2_X1 U10831 ( .A(n8415), .B(SI_11_), .ZN(n8630) );
  INV_X1 U10832 ( .A(n8415), .ZN(n8416) );
  MUX2_X1 U10833 ( .A(n13505), .B(n9673), .S(n7274), .Z(n8418) );
  XNOR2_X1 U10834 ( .A(n8418), .B(SI_12_), .ZN(n8646) );
  NAND2_X1 U10835 ( .A1(n8418), .A2(n8417), .ZN(n8419) );
  MUX2_X1 U10836 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n7274), .Z(n8420) );
  XNOR2_X1 U10837 ( .A(n8420), .B(n9578), .ZN(n8662) );
  INV_X1 U10838 ( .A(n8420), .ZN(n8421) );
  NAND2_X1 U10839 ( .A1(n8422), .A2(n9707), .ZN(n8423) );
  MUX2_X1 U10840 ( .A(n9894), .B(n9897), .S(n7274), .Z(n8675) );
  MUX2_X1 U10841 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n7274), .Z(n8425) );
  XNOR2_X1 U10842 ( .A(n8425), .B(SI_15_), .ZN(n8692) );
  INV_X1 U10843 ( .A(n8425), .ZN(n8426) );
  INV_X1 U10844 ( .A(SI_15_), .ZN(n9884) );
  NAND2_X1 U10845 ( .A1(n8426), .A2(n9884), .ZN(n8427) );
  MUX2_X1 U10846 ( .A(n10496), .B(n10529), .S(n7274), .Z(n8428) );
  XNOR2_X1 U10847 ( .A(n8428), .B(SI_16_), .ZN(n8707) );
  NAND2_X1 U10848 ( .A1(n8428), .A2(n9886), .ZN(n8429) );
  MUX2_X1 U10849 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n7274), .Z(n8727) );
  NOR2_X1 U10850 ( .A1(n8727), .A2(SI_17_), .ZN(n8430) );
  INV_X1 U10851 ( .A(SI_18_), .ZN(n10350) );
  MUX2_X1 U10852 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n7274), .Z(n8751) );
  INV_X1 U10853 ( .A(n8751), .ZN(n8431) );
  NAND2_X1 U10854 ( .A1(n8432), .A2(SI_19_), .ZN(n8757) );
  OAI21_X1 U10855 ( .B1(n10350), .B2(n8431), .A(n8757), .ZN(n8437) );
  NOR2_X1 U10856 ( .A1(n8751), .A2(SI_18_), .ZN(n8435) );
  INV_X1 U10857 ( .A(n8432), .ZN(n8433) );
  NAND2_X1 U10858 ( .A1(n8433), .A2(n10425), .ZN(n8756) );
  INV_X1 U10859 ( .A(n8756), .ZN(n8434) );
  AOI21_X1 U10860 ( .B1(n8435), .B2(n8757), .A(n8434), .ZN(n8436) );
  INV_X1 U10861 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n13338) );
  INV_X1 U10862 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11103) );
  MUX2_X1 U10863 ( .A(n13338), .B(n11103), .S(n7274), .Z(n8778) );
  INV_X1 U10864 ( .A(n8778), .ZN(n8438) );
  MUX2_X1 U10865 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n7274), .Z(n8441) );
  XNOR2_X1 U10866 ( .A(n8441), .B(SI_21_), .ZN(n8791) );
  NAND2_X1 U10867 ( .A1(n8441), .A2(SI_21_), .ZN(n8442) );
  INV_X1 U10868 ( .A(n8804), .ZN(n8443) );
  MUX2_X1 U10869 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n7274), .Z(n8805) );
  NAND2_X1 U10870 ( .A1(n8443), .A2(n8805), .ZN(n8446) );
  NAND2_X1 U10871 ( .A1(n8444), .A2(SI_22_), .ZN(n8445) );
  INV_X1 U10872 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11890) );
  XNOR2_X1 U10873 ( .A(n8447), .B(SI_23_), .ZN(n8815) );
  INV_X1 U10874 ( .A(n8447), .ZN(n8448) );
  NAND2_X1 U10875 ( .A1(n8448), .A2(SI_23_), .ZN(n8449) );
  INV_X1 U10876 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11903) );
  MUX2_X1 U10877 ( .A(n11903), .B(n11721), .S(n7274), .Z(n8450) );
  XNOR2_X1 U10878 ( .A(n8450), .B(SI_24_), .ZN(n8828) );
  INV_X1 U10879 ( .A(n8450), .ZN(n8451) );
  NAND2_X1 U10880 ( .A1(n8452), .A2(n13365), .ZN(n8455) );
  INV_X1 U10881 ( .A(n8452), .ZN(n8453) );
  NAND2_X1 U10882 ( .A1(n8453), .A2(SI_25_), .ZN(n8454) );
  NAND2_X1 U10883 ( .A1(n8455), .A2(n8454), .ZN(n8841) );
  OAI21_X2 U10884 ( .B1(n8842), .B2(n8841), .A(n8455), .ZN(n8854) );
  MUX2_X1 U10885 ( .A(n15028), .B(n14313), .S(n7274), .Z(n8852) );
  NAND2_X1 U10886 ( .A1(n8854), .A2(n13511), .ZN(n8456) );
  NAND2_X1 U10887 ( .A1(n8457), .A2(n8456), .ZN(n8868) );
  MUX2_X1 U10888 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n7274), .Z(n8458) );
  XNOR2_X1 U10889 ( .A(n8458), .B(SI_28_), .ZN(n8879) );
  INV_X1 U10890 ( .A(n8458), .ZN(n8459) );
  NAND2_X1 U10891 ( .A1(n8459), .A2(n12535), .ZN(n8460) );
  INV_X1 U10892 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15021) );
  MUX2_X1 U10893 ( .A(n15021), .B(n12020), .S(n7274), .Z(n9190) );
  XNOR2_X1 U10894 ( .A(n9190), .B(SI_29_), .ZN(n9188) );
  XNOR2_X2 U10895 ( .A(n8464), .B(n8463), .ZN(n8980) );
  NAND2_X1 U10896 ( .A1(n12447), .A2(n9235), .ZN(n8468) );
  OR2_X1 U10897 ( .A1(n6847), .A2(n12020), .ZN(n8467) );
  XOR2_X1 U10898 ( .A(n13891), .B(n14179), .Z(n9294) );
  NAND2_X1 U10899 ( .A1(n8536), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U10900 ( .A1(n8484), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U10901 ( .A1(n8486), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8470) );
  NAND2_X1 U10902 ( .A1(n8485), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8469) );
  INV_X1 U10903 ( .A(n8474), .ZN(n8475) );
  NAND2_X1 U10904 ( .A1(n8476), .A2(n8475), .ZN(n8477) );
  NAND2_X1 U10905 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8479) );
  INV_X1 U10906 ( .A(n8481), .ZN(n8482) );
  NAND2_X1 U10907 ( .A1(n8484), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U10908 ( .A1(n8485), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U10909 ( .A1(n8486), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8487) );
  AND3_X1 U10910 ( .A1(n8489), .A2(n8488), .A3(n8487), .ZN(n8491) );
  NAND2_X1 U10911 ( .A1(n8536), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8490) );
  NAND2_X1 U10912 ( .A1(n7274), .A2(SI_0_), .ZN(n8492) );
  XNOR2_X1 U10913 ( .A(n8492), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n14315) );
  NAND2_X1 U10914 ( .A1(n9026), .A2(n10143), .ZN(n9902) );
  INV_X1 U10915 ( .A(n9902), .ZN(n10138) );
  INV_X1 U10916 ( .A(n9901), .ZN(n11801) );
  NAND2_X1 U10917 ( .A1(n11801), .A2(n9900), .ZN(n8493) );
  NAND2_X1 U10918 ( .A1(n8536), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8497) );
  NAND2_X1 U10919 ( .A1(n8871), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U10920 ( .A1(n9201), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U10921 ( .A1(n8738), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U10922 ( .A1(n8500), .A2(n8499), .ZN(n8501) );
  NAND2_X1 U10923 ( .A1(n8501), .A2(n8511), .ZN(n9791) );
  NOR2_X1 U10924 ( .A1(n9791), .A2(n8478), .ZN(n8507) );
  NOR2_X1 U10925 ( .A1(n8481), .A2(n14300), .ZN(n8502) );
  MUX2_X1 U10926 ( .A(n14300), .B(n8502), .S(P2_IR_REG_2__SCAN_IN), .Z(n8503)
         );
  INV_X1 U10927 ( .A(n8503), .ZN(n8505) );
  INV_X1 U10928 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8504) );
  NAND2_X1 U10929 ( .A1(n8481), .A2(n8504), .ZN(n8514) );
  NAND2_X1 U10930 ( .A1(n8505), .A2(n8514), .ZN(n9480) );
  OAI22_X1 U10931 ( .A1(n9236), .A2(n9368), .B1(n9425), .B2(n9480), .ZN(n8506)
         );
  OR2_X2 U10932 ( .A1(n8507), .A2(n8506), .ZN(n14158) );
  NAND2_X1 U10933 ( .A1(n10135), .A2(n14158), .ZN(n8942) );
  INV_X1 U10934 ( .A(n14158), .ZN(n10048) );
  NAND2_X1 U10935 ( .A1(n10048), .A2(n13915), .ZN(n8508) );
  NAND2_X1 U10936 ( .A1(n10036), .A2(n10040), .ZN(n10035) );
  NAND2_X1 U10937 ( .A1(n10135), .A2(n10048), .ZN(n8509) );
  NAND2_X1 U10938 ( .A1(n10035), .A2(n8509), .ZN(n10664) );
  NAND2_X1 U10939 ( .A1(n8511), .A2(n8510), .ZN(n8513) );
  XNOR2_X1 U10940 ( .A(n8513), .B(n8512), .ZN(n10005) );
  NAND2_X1 U10941 ( .A1(n10005), .A2(n9235), .ZN(n8519) );
  INV_X2 U10942 ( .A(n9236), .ZN(n8765) );
  INV_X2 U10943 ( .A(n9425), .ZN(n8764) );
  NAND2_X1 U10944 ( .A1(n8514), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8515) );
  MUX2_X1 U10945 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8515), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8517) );
  INV_X1 U10946 ( .A(n8516), .ZN(n8531) );
  AND2_X1 U10947 ( .A1(n8517), .A2(n8531), .ZN(n9484) );
  AOI22_X1 U10948 ( .A1(n8765), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8764), .B2(
        n9484), .ZN(n8518) );
  NAND2_X1 U10949 ( .A1(n8536), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n8524) );
  INV_X1 U10950 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U10951 ( .A1(n8871), .A2(n9937), .ZN(n8523) );
  NAND2_X1 U10952 ( .A1(n8983), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U10953 ( .A1(n8738), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8521) );
  NAND4_X1 U10954 ( .A1(n8524), .A2(n8523), .A3(n8522), .A4(n8521), .ZN(n13914) );
  XNOR2_X1 U10955 ( .A(n9941), .B(n13914), .ZN(n10666) );
  INV_X1 U10956 ( .A(n10666), .ZN(n10663) );
  NAND2_X1 U10957 ( .A1(n10664), .A2(n10663), .ZN(n10662) );
  OR2_X1 U10958 ( .A1(n9941), .A2(n13914), .ZN(n8525) );
  AND2_X1 U10959 ( .A1(n8527), .A2(n8526), .ZN(n8529) );
  NAND2_X1 U10960 ( .A1(n10011), .A2(n9235), .ZN(n8535) );
  NAND2_X1 U10961 ( .A1(n8531), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8530) );
  MUX2_X1 U10962 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8530), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8533) );
  INV_X1 U10963 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U10964 ( .A1(n8516), .A2(n8532), .ZN(n8543) );
  NAND2_X1 U10965 ( .A1(n8533), .A2(n8543), .ZN(n9608) );
  INV_X1 U10966 ( .A(n9608), .ZN(n9487) );
  AOI22_X1 U10967 ( .A1(n8765), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8764), .B2(
        n9487), .ZN(n8534) );
  NAND2_X1 U10968 ( .A1(n8535), .A2(n8534), .ZN(n10687) );
  NAND2_X1 U10969 ( .A1(n8738), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U10970 ( .A1(n8536), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n8538) );
  NOR2_X1 U10971 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8537) );
  NOR2_X1 U10972 ( .A1(n8549), .A2(n8537), .ZN(n10686) );
  OR2_X1 U10973 ( .A1(n10687), .A2(n13913), .ZN(n8540) );
  NAND2_X1 U10974 ( .A1(n8543), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8544) );
  MUX2_X1 U10975 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8544), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8547) );
  AND3_X1 U10976 ( .A1(n8481), .A2(n8546), .A3(n8545), .ZN(n8648) );
  INV_X1 U10977 ( .A(n8648), .ZN(n8711) );
  AOI22_X1 U10978 ( .A1(n8765), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8764), .B2(
        n9490), .ZN(n8548) );
  NAND2_X1 U10979 ( .A1(n8738), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U10980 ( .A1(n8536), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8553) );
  NOR2_X1 U10981 ( .A1(n8549), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8550) );
  NOR2_X1 U10982 ( .A1(n8563), .A2(n8550), .ZN(n12004) );
  NAND2_X1 U10983 ( .A1(n8871), .A2(n12004), .ZN(n8552) );
  NAND2_X1 U10984 ( .A1(n9201), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8551) );
  NAND4_X1 U10985 ( .A1(n8554), .A2(n8553), .A3(n8552), .A4(n8551), .ZN(n13912) );
  XNOR2_X1 U10986 ( .A(n10372), .B(n13912), .ZN(n9280) );
  INV_X1 U10987 ( .A(n10372), .ZN(n12003) );
  INV_X1 U10988 ( .A(n13912), .ZN(n10544) );
  NAND2_X1 U10989 ( .A1(n12003), .A2(n10544), .ZN(n8555) );
  NAND2_X1 U10990 ( .A1(n10269), .A2(n8555), .ZN(n10542) );
  OR2_X1 U10991 ( .A1(n8557), .A2(n8556), .ZN(n8558) );
  NAND2_X1 U10992 ( .A1(n8559), .A2(n8558), .ZN(n10402) );
  OR2_X1 U10993 ( .A1(n10402), .A2(n8478), .ZN(n8562) );
  OR2_X1 U10994 ( .A1(n8648), .A2(n14300), .ZN(n8560) );
  XNOR2_X1 U10995 ( .A(n8560), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9506) );
  AOI22_X1 U10996 ( .A1(n8765), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8764), .B2(
        n9506), .ZN(n8561) );
  NAND2_X1 U10997 ( .A1(n8562), .A2(n8561), .ZN(n10655) );
  NAND2_X1 U10998 ( .A1(n8738), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8568) );
  NAND2_X1 U10999 ( .A1(n8536), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n8567) );
  NOR2_X1 U11000 ( .A1(n8563), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8564) );
  NOR2_X1 U11001 ( .A1(n8577), .A2(n8564), .ZN(n10654) );
  NAND2_X1 U11002 ( .A1(n8871), .A2(n10654), .ZN(n8566) );
  NAND2_X1 U11003 ( .A1(n8983), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n8565) );
  NAND4_X1 U11004 ( .A1(n8568), .A2(n8567), .A3(n8566), .A4(n8565), .ZN(n13911) );
  INV_X1 U11005 ( .A(n13911), .ZN(n12006) );
  XNOR2_X1 U11006 ( .A(n10655), .B(n12006), .ZN(n10546) );
  OR2_X1 U11007 ( .A1(n10655), .A2(n13911), .ZN(n8569) );
  NAND2_X1 U11008 ( .A1(n8572), .A2(n8571), .ZN(n10454) );
  OR2_X1 U11009 ( .A1(n10454), .A2(n8478), .ZN(n8576) );
  INV_X1 U11010 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11011 ( .A1(n8648), .A2(n8573), .ZN(n8587) );
  NAND2_X1 U11012 ( .A1(n8587), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8574) );
  XNOR2_X1 U11013 ( .A(n8574), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9586) );
  AOI22_X1 U11014 ( .A1(n8765), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8764), .B2(
        n9586), .ZN(n8575) );
  NAND2_X1 U11015 ( .A1(n8738), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U11016 ( .A1(n8536), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8580) );
  OAI21_X1 U11017 ( .B1(n8577), .B2(P2_REG3_REG_7__SCAN_IN), .A(n8592), .ZN(
        n10391) );
  INV_X1 U11018 ( .A(n10391), .ZN(n15330) );
  NAND2_X1 U11019 ( .A1(n8871), .A2(n15330), .ZN(n8579) );
  NAND2_X1 U11020 ( .A1(n8983), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8578) );
  NAND4_X1 U11021 ( .A1(n8581), .A2(n8580), .A3(n8579), .A4(n8578), .ZN(n13910) );
  INV_X1 U11022 ( .A(n13910), .ZN(n10645) );
  XNOR2_X1 U11023 ( .A(n15326), .B(n10645), .ZN(n10610) );
  OR2_X1 U11024 ( .A1(n15326), .A2(n13910), .ZN(n8582) );
  OR2_X1 U11025 ( .A1(n8584), .A2(n8583), .ZN(n8585) );
  NAND2_X1 U11026 ( .A1(n8586), .A2(n8585), .ZN(n10570) );
  OR2_X1 U11027 ( .A1(n10570), .A2(n8478), .ZN(n8590) );
  NAND2_X1 U11028 ( .A1(n8604), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8588) );
  XNOR2_X1 U11029 ( .A(n8588), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9861) );
  AOI22_X1 U11030 ( .A1(n8765), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8764), .B2(
        n9861), .ZN(n8589) );
  NAND2_X1 U11031 ( .A1(n8536), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11032 ( .A1(n8983), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8596) );
  AND2_X1 U11033 ( .A1(n8592), .A2(n8591), .ZN(n8593) );
  NOR2_X1 U11034 ( .A1(n8610), .A2(n8593), .ZN(n10703) );
  NAND2_X1 U11035 ( .A1(n8871), .A2(n10703), .ZN(n8595) );
  NAND2_X1 U11036 ( .A1(n8738), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8594) );
  NAND4_X1 U11037 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), .ZN(n13909) );
  XNOR2_X1 U11038 ( .A(n10704), .B(n13909), .ZN(n10695) );
  INV_X1 U11039 ( .A(n10695), .ZN(n8598) );
  NAND2_X1 U11040 ( .A1(n10704), .A2(n13909), .ZN(n8599) );
  NAND2_X1 U11041 ( .A1(n10694), .A2(n8599), .ZN(n10769) );
  INV_X1 U11042 ( .A(n8604), .ZN(n8606) );
  INV_X1 U11043 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U11044 ( .A1(n8606), .A2(n8605), .ZN(n8619) );
  NAND2_X1 U11045 ( .A1(n8619), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8607) );
  XNOR2_X1 U11046 ( .A(n8607), .B(P2_IR_REG_9__SCAN_IN), .ZN(n13925) );
  AOI22_X1 U11047 ( .A1(n8765), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8764), .B2(
        n13925), .ZN(n8608) );
  NAND2_X1 U11048 ( .A1(n8536), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8615) );
  NAND2_X1 U11049 ( .A1(n8983), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n8614) );
  OR2_X1 U11050 ( .A1(n8610), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8611) );
  AND2_X1 U11051 ( .A1(n8638), .A2(n8611), .ZN(n10879) );
  NAND2_X1 U11052 ( .A1(n8871), .A2(n10879), .ZN(n8613) );
  NAND2_X1 U11053 ( .A1(n8738), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8612) );
  NAND4_X1 U11054 ( .A1(n8615), .A2(n8614), .A3(n8613), .A4(n8612), .ZN(n13908) );
  NAND2_X1 U11055 ( .A1(n10890), .A2(n13908), .ZN(n8616) );
  XNOR2_X1 U11056 ( .A(n8618), .B(n8617), .ZN(n11107) );
  NAND2_X1 U11057 ( .A1(n11107), .A2(n9235), .ZN(n8624) );
  INV_X1 U11058 ( .A(n8619), .ZN(n8621) );
  INV_X1 U11059 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U11060 ( .A1(n8621), .A2(n8620), .ZN(n8632) );
  NAND2_X1 U11061 ( .A1(n8632), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8622) );
  XNOR2_X1 U11062 ( .A(n8622), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10060) );
  AOI22_X1 U11063 ( .A1(n8765), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n8764), 
        .B2(n10060), .ZN(n8623) );
  NAND2_X1 U11064 ( .A1(n8738), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U11065 ( .A1(n8536), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8627) );
  XNOR2_X1 U11066 ( .A(n8638), .B(P2_REG3_REG_10__SCAN_IN), .ZN(n10899) );
  NAND2_X1 U11067 ( .A1(n8871), .A2(n10899), .ZN(n8626) );
  NAND2_X1 U11068 ( .A1(n8983), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8625) );
  NAND4_X1 U11069 ( .A1(n8628), .A2(n8627), .A3(n8626), .A4(n8625), .ZN(n13907) );
  XNOR2_X1 U11070 ( .A(n10906), .B(n13907), .ZN(n9285) );
  NAND2_X1 U11071 ( .A1(n10906), .A2(n13907), .ZN(n8629) );
  XNOR2_X1 U11072 ( .A(n8631), .B(n8630), .ZN(n11138) );
  NAND2_X1 U11073 ( .A1(n11138), .A2(n9235), .ZN(n8635) );
  OAI21_X1 U11074 ( .B1(n8632), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8633) );
  XNOR2_X1 U11075 ( .A(n8633), .B(P2_IR_REG_11__SCAN_IN), .ZN(n13942) );
  AOI22_X1 U11076 ( .A1(n8765), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8764), 
        .B2(n13942), .ZN(n8634) );
  NAND2_X1 U11077 ( .A1(n8738), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U11078 ( .A1(n8536), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8642) );
  INV_X1 U11079 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8637) );
  INV_X1 U11080 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8636) );
  OAI21_X1 U11081 ( .B1(n8638), .B2(n8637), .A(n8636), .ZN(n8639) );
  AND2_X1 U11082 ( .A1(n8639), .A2(n8654), .ZN(n11224) );
  NAND2_X1 U11083 ( .A1(n8871), .A2(n11224), .ZN(n8641) );
  NAND2_X1 U11084 ( .A1(n8983), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8640) );
  NAND4_X1 U11085 ( .A1(n8643), .A2(n8642), .A3(n8641), .A4(n8640), .ZN(n13906) );
  AND2_X1 U11086 ( .A1(n11229), .A2(n13906), .ZN(n8644) );
  OR2_X1 U11087 ( .A1(n11229), .A2(n13906), .ZN(n8645) );
  XNOR2_X1 U11088 ( .A(n8647), .B(n8646), .ZN(n11297) );
  NAND2_X1 U11089 ( .A1(n11297), .A2(n9235), .ZN(n8653) );
  NAND2_X1 U11090 ( .A1(n8648), .A2(n8710), .ZN(n8650) );
  NAND2_X1 U11091 ( .A1(n8650), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8649) );
  MUX2_X1 U11092 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8649), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8651) );
  AOI22_X1 U11093 ( .A1(n8765), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8764), 
        .B2(n10064), .ZN(n8652) );
  NAND2_X1 U11094 ( .A1(n8738), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U11095 ( .A1(n8536), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n8658) );
  AND2_X1 U11096 ( .A1(n8654), .A2(n13485), .ZN(n8655) );
  NOR2_X1 U11097 ( .A1(n8682), .A2(n8655), .ZN(n15131) );
  NAND2_X1 U11098 ( .A1(n8871), .A2(n15131), .ZN(n8657) );
  NAND2_X1 U11099 ( .A1(n8983), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8656) );
  NAND4_X1 U11100 ( .A1(n8659), .A2(n8658), .A3(n8657), .A4(n8656), .ZN(n13905) );
  OR2_X1 U11101 ( .A1(n15135), .A2(n11417), .ZN(n8955) );
  NAND2_X1 U11102 ( .A1(n15135), .A2(n11417), .ZN(n8660) );
  NAND2_X1 U11103 ( .A1(n8955), .A2(n8660), .ZN(n15134) );
  OR2_X1 U11104 ( .A1(n15135), .A2(n13905), .ZN(n8661) );
  XNOR2_X1 U11105 ( .A(n8663), .B(n8662), .ZN(n11423) );
  NAND2_X1 U11106 ( .A1(n11423), .A2(n9235), .ZN(n8668) );
  NAND2_X1 U11107 ( .A1(n8665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8664) );
  MUX2_X1 U11108 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8664), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n8666) );
  NAND2_X1 U11109 ( .A1(n8666), .A2(n8694), .ZN(n11002) );
  INV_X1 U11110 ( .A(n11002), .ZN(n15292) );
  AOI22_X1 U11111 ( .A1(n8765), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8764), 
        .B2(n15292), .ZN(n8667) );
  NAND2_X1 U11112 ( .A1(n8536), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n8672) );
  INV_X1 U11113 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8684) );
  XNOR2_X1 U11114 ( .A(n8682), .B(n8684), .ZN(n11415) );
  NAND2_X1 U11115 ( .A1(n8871), .A2(n11415), .ZN(n8671) );
  NAND2_X1 U11116 ( .A1(n9201), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11117 ( .A1(n8738), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8669) );
  NAND4_X1 U11118 ( .A1(n8672), .A2(n8671), .A3(n8670), .A4(n8669), .ZN(n11414) );
  NOR2_X1 U11119 ( .A1(n15148), .A2(n11414), .ZN(n8673) );
  NAND2_X1 U11120 ( .A1(n15148), .A2(n11414), .ZN(n8674) );
  NAND2_X1 U11121 ( .A1(n8676), .A2(n8675), .ZN(n8677) );
  NAND2_X1 U11122 ( .A1(n8678), .A2(n8677), .ZN(n11449) );
  OR2_X1 U11123 ( .A1(n11449), .A2(n8478), .ZN(n8681) );
  NAND2_X1 U11124 ( .A1(n8694), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8679) );
  XNOR2_X1 U11125 ( .A(n8679), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11268) );
  AOI22_X1 U11126 ( .A1(n8765), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8764), 
        .B2(n11268), .ZN(n8680) );
  INV_X1 U11127 ( .A(n8682), .ZN(n8685) );
  INV_X1 U11128 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8683) );
  OAI21_X1 U11129 ( .B1(n8685), .B2(n8684), .A(n8683), .ZN(n8686) );
  NAND2_X1 U11130 ( .A1(n8699), .A2(n8686), .ZN(n15110) );
  INV_X1 U11131 ( .A(n15110), .ZN(n15116) );
  NAND2_X1 U11132 ( .A1(n15116), .A2(n8871), .ZN(n8690) );
  NAND2_X1 U11133 ( .A1(n8536), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U11134 ( .A1(n8983), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8688) );
  NAND2_X1 U11135 ( .A1(n8738), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8687) );
  NAND4_X1 U11136 ( .A1(n8690), .A2(n8689), .A3(n8688), .A4(n8687), .ZN(n13904) );
  AND2_X1 U11137 ( .A1(n15119), .A2(n13904), .ZN(n8691) );
  XNOR2_X1 U11138 ( .A(n8693), .B(n8692), .ZN(n11641) );
  NAND2_X1 U11139 ( .A1(n11641), .A2(n9235), .ZN(n8697) );
  OAI21_X1 U11140 ( .B1(n8694), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8695) );
  XNOR2_X1 U11141 ( .A(n8695), .B(P2_IR_REG_15__SCAN_IN), .ZN(n15301) );
  AOI22_X1 U11142 ( .A1(n8765), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8764), 
        .B2(n15301), .ZN(n8696) );
  INV_X1 U11143 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11519) );
  INV_X1 U11144 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n13339) );
  OAI22_X1 U11145 ( .A1(n8520), .A2(n11519), .B1(n9204), .B2(n13339), .ZN(
        n8703) );
  INV_X1 U11146 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8698) );
  NAND2_X1 U11147 ( .A1(n8699), .A2(n8698), .ZN(n8700) );
  NAND2_X1 U11148 ( .A1(n8721), .A2(n8700), .ZN(n13879) );
  INV_X1 U11149 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8701) );
  OAI22_X1 U11150 ( .A1(n13879), .A2(n8887), .B1(n8891), .B2(n8701), .ZN(n8702) );
  XNOR2_X1 U11151 ( .A(n14257), .B(n13903), .ZN(n11513) );
  INV_X1 U11152 ( .A(n11513), .ZN(n8704) );
  NAND2_X1 U11153 ( .A1(n11511), .A2(n8704), .ZN(n8706) );
  OR2_X1 U11154 ( .A1(n14257), .A2(n13903), .ZN(n8705) );
  NAND2_X1 U11155 ( .A1(n11814), .A2(n9235), .ZN(n8719) );
  NAND2_X1 U11156 ( .A1(n8710), .A2(n8709), .ZN(n8712) );
  NAND2_X1 U11157 ( .A1(n8714), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8713) );
  MUX2_X1 U11158 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8713), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8717) );
  INV_X1 U11159 ( .A(n8714), .ZN(n8716) );
  INV_X1 U11160 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U11161 ( .A1(n8716), .A2(n8715), .ZN(n8730) );
  NAND2_X1 U11162 ( .A1(n8717), .A2(n8730), .ZN(n11776) );
  INV_X1 U11163 ( .A(n11776), .ZN(n11781) );
  AOI22_X1 U11164 ( .A1(n8765), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8764), 
        .B2(n11781), .ZN(n8718) );
  NAND2_X1 U11165 ( .A1(n8721), .A2(n8720), .ZN(n8722) );
  NAND2_X1 U11166 ( .A1(n8736), .A2(n8722), .ZN(n13833) );
  AOI22_X1 U11167 ( .A1(n8738), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n8536), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U11168 ( .A1(n8983), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8723) );
  OAI211_X1 U11169 ( .C1(n13833), .C2(n8887), .A(n8724), .B(n8723), .ZN(n13902) );
  XNOR2_X1 U11170 ( .A(n14251), .B(n13902), .ZN(n11629) );
  NAND2_X1 U11171 ( .A1(n14251), .A2(n13902), .ZN(n8726) );
  XNOR2_X1 U11172 ( .A(n8727), .B(n13366), .ZN(n8728) );
  NAND2_X1 U11173 ( .A1(n11819), .A2(n9235), .ZN(n8734) );
  NAND2_X1 U11174 ( .A1(n8730), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8731) );
  MUX2_X1 U11175 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8731), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8732) );
  AND2_X1 U11176 ( .A1(n8732), .A2(n8760), .ZN(n11784) );
  AOI22_X1 U11177 ( .A1(n8765), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8764), 
        .B2(n11784), .ZN(n8733) );
  INV_X1 U11178 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n11777) );
  INV_X1 U11179 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8735) );
  NAND2_X1 U11180 ( .A1(n8736), .A2(n8735), .ZN(n8737) );
  NAND2_X1 U11181 ( .A1(n8746), .A2(n8737), .ZN(n11710) );
  OR2_X1 U11182 ( .A1(n11710), .A2(n8887), .ZN(n8740) );
  AOI22_X1 U11183 ( .A1(n8738), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n8536), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n8739) );
  OAI211_X1 U11184 ( .C1(n8520), .C2(n11777), .A(n8740), .B(n8739), .ZN(n13901) );
  INV_X1 U11185 ( .A(n13901), .ZN(n13834) );
  XNOR2_X1 U11186 ( .A(n14293), .B(n13834), .ZN(n11703) );
  NAND2_X1 U11187 ( .A1(n14293), .A2(n13901), .ZN(n8741) );
  XNOR2_X1 U11188 ( .A(n8753), .B(SI_18_), .ZN(n8752) );
  XNOR2_X1 U11189 ( .A(n8752), .B(n8751), .ZN(n11830) );
  NAND2_X1 U11190 ( .A1(n11830), .A2(n9235), .ZN(n8744) );
  NAND2_X1 U11191 ( .A1(n8760), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8742) );
  XNOR2_X1 U11192 ( .A(n8742), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13952) );
  AOI22_X1 U11193 ( .A1(n8765), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8764), 
        .B2(n13952), .ZN(n8743) );
  NAND2_X2 U11194 ( .A1(n8744), .A2(n8743), .ZN(n14237) );
  INV_X1 U11195 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n11786) );
  INV_X1 U11196 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U11197 ( .A1(n8746), .A2(n8745), .ZN(n8747) );
  NAND2_X1 U11198 ( .A1(n8769), .A2(n8747), .ZN(n14148) );
  OR2_X1 U11199 ( .A1(n14148), .A2(n8887), .ZN(n8749) );
  AOI22_X1 U11200 ( .A1(n9201), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8536), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n8748) );
  OAI211_X1 U11201 ( .C1(n8891), .C2(n11786), .A(n8749), .B(n8748), .ZN(n13900) );
  INV_X1 U11202 ( .A(n13900), .ZN(n13842) );
  XNOR2_X1 U11203 ( .A(n14237), .B(n13842), .ZN(n14142) );
  OR2_X1 U11204 ( .A1(n14237), .A2(n13900), .ZN(n8750) );
  NAND2_X1 U11205 ( .A1(n8753), .A2(SI_18_), .ZN(n8754) );
  NAND2_X1 U11206 ( .A1(n8755), .A2(n8754), .ZN(n8759) );
  NAND2_X1 U11207 ( .A1(n8757), .A2(n8756), .ZN(n8758) );
  NAND2_X1 U11208 ( .A1(n11843), .A2(n9235), .ZN(n8767) );
  NAND2_X1 U11209 ( .A1(n6696), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8763) );
  AOI22_X1 U11210 ( .A1(n8765), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9297), 
        .B2(n8764), .ZN(n8766) );
  NAND2_X1 U11211 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  AND2_X1 U11212 ( .A1(n8782), .A2(n8770), .ZN(n14128) );
  NAND2_X1 U11213 ( .A1(n14128), .A2(n8871), .ZN(n8775) );
  INV_X1 U11214 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13336) );
  NAND2_X1 U11215 ( .A1(n9201), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U11216 ( .A1(n8536), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8771) );
  OAI211_X1 U11217 ( .C1(n8891), .C2(n13336), .A(n8772), .B(n8771), .ZN(n8773)
         );
  INV_X1 U11218 ( .A(n8773), .ZN(n8774) );
  NAND2_X1 U11219 ( .A1(n8775), .A2(n8774), .ZN(n13899) );
  NOR2_X1 U11220 ( .A1(n14233), .A2(n13899), .ZN(n8776) );
  NAND2_X1 U11221 ( .A1(n14233), .A2(n13899), .ZN(n8777) );
  XNOR2_X1 U11222 ( .A(n8779), .B(n8778), .ZN(n11858) );
  NAND2_X1 U11223 ( .A1(n11858), .A2(n9235), .ZN(n8781) );
  OR2_X1 U11224 ( .A1(n6847), .A2(n11103), .ZN(n8780) );
  INV_X1 U11225 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13860) );
  NAND2_X1 U11226 ( .A1(n8782), .A2(n13860), .ZN(n8783) );
  NAND2_X1 U11227 ( .A1(n8795), .A2(n8783), .ZN(n14117) );
  OR2_X1 U11228 ( .A1(n14117), .A2(n8887), .ZN(n8788) );
  INV_X1 U11229 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n14228) );
  NAND2_X1 U11230 ( .A1(n9201), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U11231 ( .A1(n8536), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8784) );
  OAI211_X1 U11232 ( .C1(n8891), .C2(n14228), .A(n8785), .B(n8784), .ZN(n8786)
         );
  INV_X1 U11233 ( .A(n8786), .ZN(n8787) );
  NAND2_X1 U11234 ( .A1(n8788), .A2(n8787), .ZN(n13898) );
  OR2_X1 U11235 ( .A1(n14116), .A2(n13898), .ZN(n8789) );
  XNOR2_X1 U11236 ( .A(n8792), .B(n8791), .ZN(n11868) );
  NAND2_X1 U11237 ( .A1(n11868), .A2(n9235), .ZN(n8794) );
  OR2_X1 U11238 ( .A1(n6847), .A2(n11266), .ZN(n8793) );
  NAND2_X1 U11239 ( .A1(n8795), .A2(n13810), .ZN(n8796) );
  AND2_X1 U11240 ( .A1(n8820), .A2(n8796), .ZN(n14102) );
  NAND2_X1 U11241 ( .A1(n14102), .A2(n8871), .ZN(n8802) );
  INV_X1 U11242 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8799) );
  NAND2_X1 U11243 ( .A1(n8983), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8798) );
  NAND2_X1 U11244 ( .A1(n8536), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8797) );
  OAI211_X1 U11245 ( .C1(n8891), .C2(n8799), .A(n8798), .B(n8797), .ZN(n8800)
         );
  INV_X1 U11246 ( .A(n8800), .ZN(n8801) );
  NAND2_X1 U11247 ( .A1(n8802), .A2(n8801), .ZN(n13897) );
  XNOR2_X1 U11248 ( .A(n14222), .B(n13897), .ZN(n14094) );
  INV_X1 U11249 ( .A(n14094), .ZN(n14095) );
  OR2_X1 U11250 ( .A1(n14222), .A2(n13897), .ZN(n8803) );
  XNOR2_X1 U11251 ( .A(n8804), .B(n8805), .ZN(n12603) );
  NAND2_X1 U11252 ( .A1(n12603), .A2(n9235), .ZN(n8807) );
  OR2_X1 U11253 ( .A1(n6847), .A2(n12605), .ZN(n8806) );
  NAND2_X2 U11254 ( .A1(n8807), .A2(n8806), .ZN(n14087) );
  XNOR2_X1 U11255 ( .A(n8820), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n14088) );
  NAND2_X1 U11256 ( .A1(n14088), .A2(n8871), .ZN(n8812) );
  INV_X1 U11257 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n14218) );
  NAND2_X1 U11258 ( .A1(n9201), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8809) );
  NAND2_X1 U11259 ( .A1(n8536), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8808) );
  OAI211_X1 U11260 ( .C1(n8891), .C2(n14218), .A(n8809), .B(n8808), .ZN(n8810)
         );
  INV_X1 U11261 ( .A(n8810), .ZN(n8811) );
  NAND2_X1 U11262 ( .A1(n8812), .A2(n8811), .ZN(n13896) );
  NAND2_X1 U11263 ( .A1(n14087), .A2(n13896), .ZN(n8814) );
  INV_X1 U11264 ( .A(n8815), .ZN(n8816) );
  XNOR2_X1 U11265 ( .A(n8817), .B(n8816), .ZN(n11889) );
  NAND2_X1 U11266 ( .A1(n11889), .A2(n9235), .ZN(n8819) );
  OR2_X1 U11267 ( .A1(n6847), .A2(n11578), .ZN(n8818) );
  INV_X1 U11268 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12573) );
  INV_X1 U11269 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13771) );
  OAI21_X1 U11270 ( .B1(n8820), .B2(n12573), .A(n13771), .ZN(n8821) );
  NAND2_X1 U11271 ( .A1(n8821), .A2(n8833), .ZN(n14073) );
  OR2_X1 U11272 ( .A1(n14073), .A2(n8887), .ZN(n8826) );
  INV_X1 U11273 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n13405) );
  NAND2_X1 U11274 ( .A1(n8738), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8823) );
  NAND2_X1 U11275 ( .A1(n9201), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8822) );
  OAI211_X1 U11276 ( .C1(n9204), .C2(n13405), .A(n8823), .B(n8822), .ZN(n8824)
         );
  INV_X1 U11277 ( .A(n8824), .ZN(n8825) );
  NAND2_X1 U11278 ( .A1(n8826), .A2(n8825), .ZN(n13895) );
  INV_X1 U11279 ( .A(n13895), .ZN(n8969) );
  XNOR2_X1 U11280 ( .A(n14210), .B(n8969), .ZN(n14068) );
  OR2_X1 U11281 ( .A1(n14210), .A2(n13895), .ZN(n8827) );
  INV_X1 U11282 ( .A(n8828), .ZN(n8829) );
  XNOR2_X1 U11283 ( .A(n8830), .B(n8829), .ZN(n11902) );
  NAND2_X1 U11284 ( .A1(n11902), .A2(n9235), .ZN(n8832) );
  OR2_X1 U11285 ( .A1(n6847), .A2(n11721), .ZN(n8831) );
  NAND2_X2 U11286 ( .A1(n8832), .A2(n8831), .ZN(n14205) );
  NAND2_X1 U11287 ( .A1(n8833), .A2(n13852), .ZN(n8834) );
  NAND2_X1 U11288 ( .A1(n8845), .A2(n8834), .ZN(n13851) );
  OR2_X1 U11289 ( .A1(n13851), .A2(n8887), .ZN(n8839) );
  INV_X1 U11290 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13430) );
  NAND2_X1 U11291 ( .A1(n8738), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U11292 ( .A1(n9201), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8835) );
  OAI211_X1 U11293 ( .C1(n9204), .C2(n13430), .A(n8836), .B(n8835), .ZN(n8837)
         );
  INV_X1 U11294 ( .A(n8837), .ZN(n8838) );
  NAND2_X1 U11295 ( .A1(n8839), .A2(n8838), .ZN(n14026) );
  INV_X1 U11296 ( .A(n14026), .ZN(n13822) );
  NAND2_X1 U11297 ( .A1(n14205), .A2(n14026), .ZN(n8840) );
  XNOR2_X1 U11298 ( .A(n8842), .B(n8841), .ZN(n11915) );
  NAND2_X1 U11299 ( .A1(n11915), .A2(n9235), .ZN(n8844) );
  OR2_X1 U11300 ( .A1(n6847), .A2(n11723), .ZN(n8843) );
  NAND2_X1 U11301 ( .A1(n8845), .A2(n13821), .ZN(n8846) );
  NAND2_X1 U11302 ( .A1(n8858), .A2(n8846), .ZN(n14035) );
  INV_X1 U11303 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n14202) );
  NAND2_X1 U11304 ( .A1(n9201), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U11305 ( .A1(n8536), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8847) );
  OAI211_X1 U11306 ( .C1(n8891), .C2(n14202), .A(n8848), .B(n8847), .ZN(n8849)
         );
  INV_X1 U11307 ( .A(n8849), .ZN(n8850) );
  OR2_X1 U11308 ( .A1(n14031), .A2(n13894), .ZN(n8851) );
  XNOR2_X1 U11309 ( .A(n8852), .B(SI_26_), .ZN(n8853) );
  XNOR2_X1 U11310 ( .A(n8854), .B(n8853), .ZN(n14311) );
  NAND2_X1 U11311 ( .A1(n14311), .A2(n9235), .ZN(n8856) );
  OR2_X1 U11312 ( .A1(n6847), .A2(n14313), .ZN(n8855) );
  NAND2_X1 U11313 ( .A1(n8858), .A2(n8857), .ZN(n8859) );
  NAND2_X1 U11314 ( .A1(n14011), .A2(n8871), .ZN(n8864) );
  INV_X1 U11315 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n13443) );
  NAND2_X1 U11316 ( .A1(n8738), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8861) );
  NAND2_X1 U11317 ( .A1(n8983), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8860) );
  OAI211_X1 U11318 ( .C1(n9204), .C2(n13443), .A(n8861), .B(n8860), .ZN(n8862)
         );
  INV_X1 U11319 ( .A(n8862), .ZN(n8863) );
  INV_X1 U11320 ( .A(n8865), .ZN(n8866) );
  XNOR2_X1 U11321 ( .A(n8866), .B(SI_27_), .ZN(n8867) );
  XNOR2_X1 U11322 ( .A(n8868), .B(n8867), .ZN(n11941) );
  NAND2_X1 U11323 ( .A1(n11941), .A2(n9235), .ZN(n8870) );
  OR2_X1 U11324 ( .A1(n6847), .A2(n11774), .ZN(n8869) );
  XNOR2_X1 U11325 ( .A(n8885), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13999) );
  NAND2_X1 U11326 ( .A1(n13999), .A2(n8871), .ZN(n8877) );
  INV_X1 U11327 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8874) );
  NAND2_X1 U11328 ( .A1(n9201), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8873) );
  NAND2_X1 U11329 ( .A1(n8536), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8872) );
  OAI211_X1 U11330 ( .C1(n8891), .C2(n8874), .A(n8873), .B(n8872), .ZN(n8875)
         );
  INV_X1 U11331 ( .A(n8875), .ZN(n8876) );
  XNOR2_X1 U11332 ( .A(n14189), .B(n13893), .ZN(n14003) );
  NAND2_X1 U11333 ( .A1(n14189), .A2(n13893), .ZN(n8878) );
  NAND2_X1 U11334 ( .A1(n14307), .A2(n9235), .ZN(n8882) );
  OR2_X1 U11335 ( .A1(n6847), .A2(n14310), .ZN(n8881) );
  INV_X1 U11336 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8884) );
  INV_X1 U11337 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8883) );
  OAI21_X1 U11338 ( .B1(n8885), .B2(n8884), .A(n8883), .ZN(n8886) );
  NAND2_X1 U11339 ( .A1(n8886), .A2(n9001), .ZN(n13983) );
  INV_X1 U11340 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8890) );
  NAND2_X1 U11341 ( .A1(n9201), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U11342 ( .A1(n8536), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8888) );
  OAI211_X1 U11343 ( .C1(n8891), .C2(n8890), .A(n8889), .B(n8888), .ZN(n8892)
         );
  INV_X1 U11344 ( .A(n8892), .ZN(n8893) );
  NAND2_X1 U11345 ( .A1(n14270), .A2(n13892), .ZN(n8896) );
  OR2_X1 U11346 ( .A1(n14270), .A2(n13892), .ZN(n8895) );
  NAND2_X1 U11347 ( .A1(n8896), .A2(n8895), .ZN(n13977) );
  NAND2_X1 U11348 ( .A1(n13974), .A2(n6956), .ZN(n13976) );
  NAND2_X1 U11349 ( .A1(n13976), .A2(n8896), .ZN(n8897) );
  NOR4_X1 U11350 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8901) );
  NOR4_X1 U11351 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n8900) );
  NOR4_X1 U11352 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8899) );
  NOR4_X1 U11353 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n8898) );
  NAND4_X1 U11354 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(n8918)
         );
  NOR2_X1 U11355 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .ZN(
        n8905) );
  NOR4_X1 U11356 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n8904) );
  NOR4_X1 U11357 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n8903) );
  NOR4_X1 U11358 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8902) );
  NAND4_X1 U11359 ( .A1(n8905), .A2(n8904), .A3(n8903), .A4(n8902), .ZN(n8917)
         );
  NAND2_X1 U11360 ( .A1(n8910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8906) );
  MUX2_X1 U11361 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8906), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8907) );
  NAND2_X1 U11362 ( .A1(n6732), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8909) );
  MUX2_X1 U11363 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8909), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8911) );
  NAND2_X1 U11364 ( .A1(n8911), .A2(n8910), .ZN(n11722) );
  NAND2_X1 U11365 ( .A1(n8920), .A2(n8919), .ZN(n8922) );
  NAND2_X1 U11366 ( .A1(n8922), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8914) );
  XNOR2_X1 U11367 ( .A(n11719), .B(P2_B_REG_SCAN_IN), .ZN(n8915) );
  OAI21_X1 U11368 ( .B1(n8918), .B2(n8917), .A(n15340), .ZN(n9918) );
  OR2_X1 U11369 ( .A1(n8920), .A2(n8919), .ZN(n8921) );
  NAND2_X1 U11370 ( .A1(n8922), .A2(n8921), .ZN(n9933) );
  NAND2_X1 U11371 ( .A1(n8926), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8924) );
  NAND3_X1 U11372 ( .A1(n6665), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_20__SCAN_IN), .ZN(n8928) );
  NAND2_X1 U11373 ( .A1(n14300), .A2(n8912), .ZN(n8927) );
  NAND2_X1 U11374 ( .A1(n11104), .A2(n11795), .ZN(n9928) );
  NAND2_X1 U11375 ( .A1(n9921), .A2(n9928), .ZN(n9932) );
  NAND2_X1 U11376 ( .A1(n11719), .A2(n14314), .ZN(n8931) );
  INV_X1 U11377 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15347) );
  NAND2_X1 U11378 ( .A1(n15340), .A2(n15347), .ZN(n8930) );
  NAND2_X1 U11379 ( .A1(n8931), .A2(n8930), .ZN(n15348) );
  INV_X1 U11380 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15350) );
  NAND2_X1 U11381 ( .A1(n15340), .A2(n15350), .ZN(n8933) );
  NAND2_X1 U11382 ( .A1(n14314), .A2(n11722), .ZN(n8932) );
  NAND2_X1 U11383 ( .A1(n8933), .A2(n8932), .ZN(n15351) );
  INV_X1 U11384 ( .A(n15351), .ZN(n9919) );
  AND2_X1 U11385 ( .A1(n15348), .A2(n9919), .ZN(n8934) );
  NAND2_X1 U11386 ( .A1(n9964), .A2(n8934), .ZN(n8936) );
  INV_X1 U11387 ( .A(n9931), .ZN(n8935) );
  INV_X1 U11388 ( .A(n9020), .ZN(n10148) );
  AND2_X1 U11389 ( .A1(n9899), .A2(n10148), .ZN(n8939) );
  NOR2_X1 U11390 ( .A1(n14182), .A2(n14137), .ZN(n9005) );
  INV_X1 U11391 ( .A(n14270), .ZN(n13988) );
  INV_X1 U11392 ( .A(n10143), .ZN(n8940) );
  NOR2_X1 U11393 ( .A1(n8940), .A2(n9026), .ZN(n9950) );
  OR2_X1 U11394 ( .A1(n9901), .A2(n9900), .ZN(n10039) );
  INV_X1 U11395 ( .A(n10040), .ZN(n8941) );
  NAND2_X1 U11396 ( .A1(n10043), .A2(n8942), .ZN(n10667) );
  NAND2_X1 U11397 ( .A1(n10667), .A2(n10666), .ZN(n10665) );
  INV_X1 U11398 ( .A(n13914), .ZN(n10165) );
  NAND2_X1 U11399 ( .A1(n9941), .A2(n10165), .ZN(n8943) );
  INV_X1 U11400 ( .A(n10681), .ZN(n10677) );
  NAND2_X1 U11401 ( .A1(n10687), .A2(n12011), .ZN(n10272) );
  NAND2_X1 U11402 ( .A1(n10372), .A2(n10544), .ZN(n10545) );
  NAND2_X1 U11403 ( .A1(n10547), .A2(n10545), .ZN(n8945) );
  INV_X1 U11404 ( .A(n10546), .ZN(n8944) );
  NAND2_X1 U11405 ( .A1(n8945), .A2(n8944), .ZN(n10549) );
  NAND2_X1 U11406 ( .A1(n10655), .A2(n12006), .ZN(n8946) );
  NAND2_X1 U11407 ( .A1(n10549), .A2(n8946), .ZN(n10611) );
  OR2_X1 U11408 ( .A1(n15326), .A2(n10645), .ZN(n8947) );
  NAND2_X1 U11409 ( .A1(n15326), .A2(n10645), .ZN(n8948) );
  INV_X1 U11410 ( .A(n13909), .ZN(n10881) );
  AND2_X1 U11411 ( .A1(n10704), .A2(n10881), .ZN(n8949) );
  INV_X1 U11412 ( .A(n13908), .ZN(n10902) );
  OR2_X1 U11413 ( .A1(n10890), .A2(n10902), .ZN(n8950) );
  NAND2_X1 U11414 ( .A1(n8951), .A2(n8950), .ZN(n10804) );
  NAND2_X1 U11415 ( .A1(n10804), .A2(n9285), .ZN(n8953) );
  INV_X1 U11416 ( .A(n13907), .ZN(n11226) );
  OR2_X1 U11417 ( .A1(n10906), .A2(n11226), .ZN(n8952) );
  INV_X1 U11418 ( .A(n13906), .ZN(n10903) );
  XNOR2_X1 U11419 ( .A(n11229), .B(n10903), .ZN(n10981) );
  NAND2_X1 U11420 ( .A1(n11229), .A2(n10903), .ZN(n8954) );
  NAND2_X1 U11421 ( .A1(n15129), .A2(n8955), .ZN(n11181) );
  INV_X1 U11422 ( .A(n11414), .ZN(n15097) );
  XNOR2_X1 U11423 ( .A(n15148), .B(n15097), .ZN(n11183) );
  INV_X1 U11424 ( .A(n11183), .ZN(n11180) );
  NAND2_X1 U11425 ( .A1(n11181), .A2(n11180), .ZN(n8957) );
  OR2_X1 U11426 ( .A1(n15148), .A2(n15097), .ZN(n8956) );
  NAND2_X1 U11427 ( .A1(n8957), .A2(n8956), .ZN(n15112) );
  INV_X1 U11428 ( .A(n13904), .ZN(n13880) );
  NOR2_X1 U11429 ( .A1(n15119), .A2(n13880), .ZN(n8958) );
  NAND2_X1 U11430 ( .A1(n15119), .A2(n13880), .ZN(n8959) );
  INV_X1 U11431 ( .A(n13903), .ZN(n15099) );
  NAND2_X1 U11432 ( .A1(n11630), .A2(n11629), .ZN(n11628) );
  INV_X1 U11433 ( .A(n13902), .ZN(n13882) );
  OR2_X1 U11434 ( .A1(n14251), .A2(n13882), .ZN(n8960) );
  OR2_X1 U11435 ( .A1(n14237), .A2(n13842), .ZN(n8961) );
  INV_X1 U11436 ( .A(n13899), .ZN(n14113) );
  AND2_X1 U11437 ( .A1(n14233), .A2(n14113), .ZN(n8962) );
  OR2_X1 U11438 ( .A1(n14233), .A2(n14113), .ZN(n8963) );
  INV_X1 U11439 ( .A(n13898), .ZN(n8964) );
  NAND2_X1 U11440 ( .A1(n14116), .A2(n8964), .ZN(n8966) );
  OR2_X1 U11441 ( .A1(n14116), .A2(n8964), .ZN(n8965) );
  NAND2_X1 U11442 ( .A1(n8966), .A2(n8965), .ZN(n14111) );
  INV_X1 U11443 ( .A(n13897), .ZN(n14114) );
  AND2_X1 U11444 ( .A1(n14222), .A2(n14114), .ZN(n8967) );
  INV_X1 U11445 ( .A(n13896), .ZN(n12570) );
  NAND2_X1 U11446 ( .A1(n14210), .A2(n8969), .ZN(n8968) );
  OR2_X1 U11447 ( .A1(n14210), .A2(n8969), .ZN(n8970) );
  NAND2_X1 U11448 ( .A1(n8971), .A2(n8970), .ZN(n14042) );
  NAND2_X1 U11449 ( .A1(n14205), .A2(n13822), .ZN(n8972) );
  XNOR2_X1 U11450 ( .A(n14031), .B(n13894), .ZN(n14023) );
  INV_X1 U11451 ( .A(n13894), .ZN(n8973) );
  NAND2_X1 U11452 ( .A1(n14031), .A2(n8973), .ZN(n8974) );
  INV_X1 U11453 ( .A(n14028), .ZN(n13823) );
  OR2_X1 U11454 ( .A1(n14196), .A2(n13823), .ZN(n9278) );
  NAND2_X1 U11455 ( .A1(n14196), .A2(n13823), .ZN(n9277) );
  INV_X1 U11456 ( .A(n13893), .ZN(n8975) );
  AND2_X1 U11457 ( .A1(n14189), .A2(n8975), .ZN(n8976) );
  AOI21_X1 U11458 ( .B1(n14003), .B2(n13993), .A(n8976), .ZN(n13978) );
  INV_X1 U11459 ( .A(n11104), .ZN(n8978) );
  NAND2_X1 U11460 ( .A1(n8978), .A2(n6585), .ZN(n9272) );
  INV_X1 U11461 ( .A(n9439), .ZN(n8979) );
  NAND2_X1 U11462 ( .A1(n9921), .A2(n8979), .ZN(n15096) );
  NAND2_X1 U11463 ( .A1(n13892), .A2(n14025), .ZN(n8988) );
  INV_X1 U11464 ( .A(P2_B_REG_SCAN_IN), .ZN(n8981) );
  OR2_X1 U11465 ( .A1(n8980), .A2(n8981), .ZN(n8982) );
  AND2_X1 U11466 ( .A1(n14027), .A2(n8982), .ZN(n13964) );
  NAND2_X1 U11467 ( .A1(n8738), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8986) );
  NAND2_X1 U11468 ( .A1(n8983), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8985) );
  NAND2_X1 U11469 ( .A1(n8536), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8984) );
  AND3_X1 U11470 ( .A1(n8986), .A2(n8985), .A3(n8984), .ZN(n9240) );
  INV_X1 U11471 ( .A(n9240), .ZN(n13890) );
  NAND2_X1 U11472 ( .A1(n13964), .A2(n13890), .ZN(n8987) );
  INV_X1 U11473 ( .A(n14196), .ZN(n14013) );
  INV_X1 U11474 ( .A(n14251), .ZN(n11626) );
  INV_X1 U11475 ( .A(n10890), .ZN(n10893) );
  INV_X1 U11476 ( .A(n10655), .ZN(n10562) );
  NOR2_X1 U11477 ( .A1(n10038), .A2(n14158), .ZN(n10672) );
  NAND2_X1 U11478 ( .A1(n10672), .A2(n15360), .ZN(n10683) );
  OR2_X2 U11479 ( .A1(n15136), .A2(n15135), .ZN(n15137) );
  INV_X1 U11480 ( .A(n14222), .ZN(n14105) );
  NOR2_X2 U11481 ( .A1(n6629), .A2(n14270), .ZN(n8995) );
  AOI21_X1 U11482 ( .B1(n14179), .B2(n13985), .A(n13997), .ZN(n8996) );
  AND2_X1 U11483 ( .A1(n8996), .A2(n13967), .ZN(n14178) );
  INV_X1 U11484 ( .A(n10142), .ZN(n8997) );
  NOR2_X1 U11485 ( .A1(n8997), .A2(n11104), .ZN(n9938) );
  INV_X1 U11486 ( .A(n9938), .ZN(n8998) );
  NAND2_X1 U11487 ( .A1(n14179), .A2(n15132), .ZN(n9000) );
  NAND2_X1 U11488 ( .A1(n8990), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8999) );
  OAI211_X1 U11489 ( .C1(n14147), .C2(n9001), .A(n9000), .B(n8999), .ZN(n9002)
         );
  NAND2_X1 U11490 ( .A1(n9006), .A2(n12165), .ZN(n10481) );
  NOR2_X1 U11491 ( .A1(n9008), .A2(n9007), .ZN(n9009) );
  OR2_X1 U11492 ( .A1(n10481), .A2(n9009), .ZN(n9010) );
  NAND2_X1 U11493 ( .A1(n12230), .A2(n12183), .ZN(n9982) );
  NAND2_X1 U11494 ( .A1(n10481), .A2(n9982), .ZN(n10483) );
  OAI22_X1 U11495 ( .A1(n10482), .A2(n9010), .B1(n13743), .B2(n10483), .ZN(
        n9014) );
  AND2_X1 U11496 ( .A1(n9973), .A2(n9011), .ZN(n9012) );
  INV_X1 U11497 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9015) );
  NOR2_X1 U11498 ( .A1(n15603), .A2(n9015), .ZN(n9016) );
  OAI21_X1 U11499 ( .B1(n9018), .B2(n15600), .A(n9017), .ZN(P3_U3488) );
  NAND2_X1 U11500 ( .A1(n9265), .A2(n9901), .ZN(n9022) );
  NAND2_X1 U11501 ( .A1(n7523), .A2(n14166), .ZN(n9021) );
  AOI21_X1 U11502 ( .B1(n9297), .B2(n9019), .A(n9898), .ZN(n9023) );
  OAI211_X1 U11503 ( .C1(n9026), .C2(n10143), .A(n9025), .B(n9024), .ZN(n9027)
         );
  NAND2_X1 U11504 ( .A1(n9028), .A2(n9027), .ZN(n9033) );
  NAND2_X1 U11505 ( .A1(n9265), .A2(n14166), .ZN(n9030) );
  NAND2_X1 U11506 ( .A1(n9901), .A2(n7523), .ZN(n9029) );
  NAND2_X1 U11507 ( .A1(n9030), .A2(n9029), .ZN(n9031) );
  NAND2_X1 U11508 ( .A1(n9033), .A2(n9032), .ZN(n9034) );
  NAND2_X1 U11509 ( .A1(n9265), .A2(n14158), .ZN(n9037) );
  NAND2_X1 U11510 ( .A1(n13915), .A2(n7523), .ZN(n9036) );
  NAND2_X1 U11511 ( .A1(n9037), .A2(n9036), .ZN(n9039) );
  AOI22_X1 U11512 ( .A1(n9265), .A2(n13915), .B1(n7523), .B2(n14158), .ZN(
        n9038) );
  NAND2_X1 U11513 ( .A1(n9941), .A2(n7523), .ZN(n9041) );
  NAND2_X1 U11514 ( .A1(n9173), .A2(n13914), .ZN(n9040) );
  NAND2_X1 U11515 ( .A1(n9041), .A2(n9040), .ZN(n9045) );
  NAND2_X1 U11516 ( .A1(n9046), .A2(n9045), .ZN(n9044) );
  AOI22_X1 U11517 ( .A1(n9941), .A2(n9173), .B1(n9208), .B2(n13914), .ZN(n9042) );
  NAND2_X1 U11518 ( .A1(n9044), .A2(n9043), .ZN(n9047) );
  NAND2_X1 U11519 ( .A1(n10687), .A2(n9173), .ZN(n9049) );
  NAND2_X1 U11520 ( .A1(n13913), .A2(n9208), .ZN(n9048) );
  NAND2_X1 U11521 ( .A1(n10687), .A2(n7523), .ZN(n9050) );
  NAND2_X1 U11522 ( .A1(n10372), .A2(n9208), .ZN(n9053) );
  NAND2_X1 U11523 ( .A1(n9173), .A2(n13912), .ZN(n9052) );
  NAND2_X1 U11524 ( .A1(n9053), .A2(n9052), .ZN(n9055) );
  AOI22_X1 U11525 ( .A1(n10372), .A2(n9173), .B1(n9208), .B2(n13912), .ZN(
        n9054) );
  NOR2_X1 U11526 ( .A1(n9056), .A2(n9055), .ZN(n9057) );
  NAND2_X1 U11527 ( .A1(n10655), .A2(n9173), .ZN(n9060) );
  NAND2_X1 U11528 ( .A1(n13911), .A2(n9208), .ZN(n9059) );
  NAND2_X1 U11529 ( .A1(n9060), .A2(n9059), .ZN(n9063) );
  NAND2_X1 U11530 ( .A1(n10655), .A2(n9208), .ZN(n9061) );
  OAI21_X1 U11531 ( .B1(n9208), .B2(n12006), .A(n9061), .ZN(n9062) );
  NAND2_X1 U11532 ( .A1(n15326), .A2(n9208), .ZN(n9066) );
  NAND2_X1 U11533 ( .A1(n9173), .A2(n13910), .ZN(n9065) );
  NAND2_X1 U11534 ( .A1(n9066), .A2(n9065), .ZN(n9068) );
  AOI22_X1 U11535 ( .A1(n15326), .A2(n9173), .B1(n9208), .B2(n13910), .ZN(
        n9067) );
  NOR2_X1 U11536 ( .A1(n9069), .A2(n9068), .ZN(n9070) );
  NAND2_X1 U11537 ( .A1(n10704), .A2(n9173), .ZN(n9073) );
  NAND2_X1 U11538 ( .A1(n13909), .A2(n9208), .ZN(n9072) );
  NAND2_X1 U11539 ( .A1(n9073), .A2(n9072), .ZN(n9076) );
  NAND2_X1 U11540 ( .A1(n10704), .A2(n9208), .ZN(n9074) );
  OAI21_X1 U11541 ( .B1(n9208), .B2(n10881), .A(n9074), .ZN(n9075) );
  NAND2_X1 U11542 ( .A1(n10890), .A2(n9208), .ZN(n9079) );
  NAND2_X1 U11543 ( .A1(n9173), .A2(n13908), .ZN(n9078) );
  AOI22_X1 U11544 ( .A1(n10890), .A2(n9173), .B1(n9208), .B2(n13908), .ZN(
        n9080) );
  NAND2_X1 U11545 ( .A1(n10906), .A2(n9173), .ZN(n9082) );
  NAND2_X1 U11546 ( .A1(n13907), .A2(n9208), .ZN(n9081) );
  NAND2_X1 U11547 ( .A1(n9082), .A2(n9081), .ZN(n9085) );
  AOI22_X1 U11548 ( .A1(n10906), .A2(n9208), .B1(n9173), .B2(n13907), .ZN(
        n9083) );
  AOI21_X1 U11549 ( .B1(n9086), .B2(n9085), .A(n9083), .ZN(n9084) );
  NAND2_X1 U11550 ( .A1(n11229), .A2(n9208), .ZN(n9089) );
  NAND2_X1 U11551 ( .A1(n9173), .A2(n13906), .ZN(n9088) );
  NAND2_X1 U11552 ( .A1(n9089), .A2(n9088), .ZN(n9092) );
  NAND2_X1 U11553 ( .A1(n11229), .A2(n9173), .ZN(n9090) );
  OAI21_X1 U11554 ( .B1(n10903), .B2(n9265), .A(n9090), .ZN(n9091) );
  INV_X1 U11555 ( .A(n9091), .ZN(n9093) );
  NAND2_X1 U11556 ( .A1(n15135), .A2(n9173), .ZN(n9095) );
  NAND2_X1 U11557 ( .A1(n13905), .A2(n9208), .ZN(n9094) );
  AOI22_X1 U11558 ( .A1(n15135), .A2(n9208), .B1(n9173), .B2(n13905), .ZN(
        n9096) );
  NAND2_X1 U11559 ( .A1(n15148), .A2(n9208), .ZN(n9099) );
  NAND2_X1 U11560 ( .A1(n9173), .A2(n11414), .ZN(n9098) );
  NAND2_X1 U11561 ( .A1(n9099), .A2(n9098), .ZN(n9104) );
  NAND2_X1 U11562 ( .A1(n9103), .A2(n9104), .ZN(n9102) );
  NAND2_X1 U11563 ( .A1(n15148), .A2(n9173), .ZN(n9100) );
  OAI21_X1 U11564 ( .B1(n15097), .B2(n9265), .A(n9100), .ZN(n9101) );
  NAND2_X1 U11565 ( .A1(n15119), .A2(n9173), .ZN(n9110) );
  NAND2_X1 U11566 ( .A1(n13904), .A2(n9208), .ZN(n9109) );
  AOI22_X1 U11567 ( .A1(n15119), .A2(n9208), .B1(n9173), .B2(n13904), .ZN(
        n9111) );
  NAND2_X1 U11568 ( .A1(n14257), .A2(n9208), .ZN(n9113) );
  NAND2_X1 U11569 ( .A1(n13903), .A2(n9173), .ZN(n9112) );
  NAND2_X1 U11570 ( .A1(n9113), .A2(n9112), .ZN(n9116) );
  NAND2_X1 U11571 ( .A1(n14257), .A2(n9173), .ZN(n9115) );
  NAND2_X1 U11572 ( .A1(n13903), .A2(n9208), .ZN(n9114) );
  OAI21_X1 U11573 ( .B1(n9119), .B2(n6722), .A(n9118), .ZN(n9124) );
  NAND2_X1 U11574 ( .A1(n14251), .A2(n9173), .ZN(n9121) );
  NAND2_X1 U11575 ( .A1(n13902), .A2(n9208), .ZN(n9120) );
  NAND2_X1 U11576 ( .A1(n9121), .A2(n9120), .ZN(n9123) );
  AOI22_X1 U11577 ( .A1(n14251), .A2(n9208), .B1(n9173), .B2(n13902), .ZN(
        n9122) );
  NAND2_X1 U11578 ( .A1(n14293), .A2(n9208), .ZN(n9126) );
  NAND2_X1 U11579 ( .A1(n13901), .A2(n9173), .ZN(n9125) );
  NAND2_X1 U11580 ( .A1(n9126), .A2(n9125), .ZN(n9128) );
  AOI22_X1 U11581 ( .A1(n14293), .A2(n9173), .B1(n9208), .B2(n13901), .ZN(
        n9127) );
  NAND2_X1 U11582 ( .A1(n14237), .A2(n9173), .ZN(n9131) );
  NAND2_X1 U11583 ( .A1(n13900), .A2(n9208), .ZN(n9130) );
  AOI22_X1 U11584 ( .A1(n14237), .A2(n9208), .B1(n9173), .B2(n13900), .ZN(
        n9132) );
  INV_X1 U11585 ( .A(n9132), .ZN(n9133) );
  AND2_X1 U11586 ( .A1(n13899), .A2(n9173), .ZN(n9135) );
  AOI21_X1 U11587 ( .B1(n14233), .B2(n9208), .A(n9135), .ZN(n9140) );
  INV_X1 U11588 ( .A(n9140), .ZN(n9136) );
  NAND2_X1 U11589 ( .A1(n14233), .A2(n9173), .ZN(n9137) );
  NAND2_X1 U11590 ( .A1(n9139), .A2(n9138), .ZN(n9143) );
  NAND2_X1 U11591 ( .A1(n9141), .A2(n9140), .ZN(n9142) );
  AND2_X1 U11592 ( .A1(n13898), .A2(n9208), .ZN(n9144) );
  AOI21_X1 U11593 ( .B1(n14116), .B2(n9173), .A(n9144), .ZN(n9148) );
  NAND2_X1 U11594 ( .A1(n14116), .A2(n9208), .ZN(n9146) );
  NAND2_X1 U11595 ( .A1(n13898), .A2(n9173), .ZN(n9145) );
  NAND2_X1 U11596 ( .A1(n9146), .A2(n9145), .ZN(n9147) );
  NAND2_X1 U11597 ( .A1(n14222), .A2(n9208), .ZN(n9150) );
  NAND2_X1 U11598 ( .A1(n13897), .A2(n9173), .ZN(n9149) );
  NAND2_X1 U11599 ( .A1(n9150), .A2(n9149), .ZN(n9153) );
  NAND2_X1 U11600 ( .A1(n14222), .A2(n9173), .ZN(n9151) );
  OAI21_X1 U11601 ( .B1(n14114), .B2(n9265), .A(n9151), .ZN(n9152) );
  INV_X1 U11602 ( .A(n9153), .ZN(n9154) );
  NAND2_X1 U11603 ( .A1(n14087), .A2(n9173), .ZN(n9156) );
  NAND2_X1 U11604 ( .A1(n13896), .A2(n9208), .ZN(n9155) );
  NAND2_X1 U11605 ( .A1(n9156), .A2(n9155), .ZN(n9159) );
  AOI22_X1 U11606 ( .A1(n14087), .A2(n9208), .B1(n9173), .B2(n13896), .ZN(
        n9157) );
  AOI21_X1 U11607 ( .B1(n9160), .B2(n9159), .A(n9157), .ZN(n9158) );
  NOR2_X1 U11608 ( .A1(n9160), .A2(n9159), .ZN(n9161) );
  NAND2_X1 U11609 ( .A1(n14210), .A2(n9208), .ZN(n9163) );
  NAND2_X1 U11610 ( .A1(n13895), .A2(n9173), .ZN(n9162) );
  AOI22_X1 U11611 ( .A1(n14210), .A2(n9173), .B1(n9208), .B2(n13895), .ZN(
        n9164) );
  AND2_X1 U11612 ( .A1(n13894), .A2(n9173), .ZN(n9165) );
  AOI21_X1 U11613 ( .B1(n14031), .B2(n9208), .A(n9165), .ZN(n9181) );
  NAND2_X1 U11614 ( .A1(n14031), .A2(n9173), .ZN(n9167) );
  NAND2_X1 U11615 ( .A1(n13894), .A2(n9208), .ZN(n9166) );
  NAND2_X1 U11616 ( .A1(n9167), .A2(n9166), .ZN(n9180) );
  NAND2_X1 U11617 ( .A1(n9181), .A2(n9180), .ZN(n9185) );
  AND2_X1 U11618 ( .A1(n14026), .A2(n9173), .ZN(n9168) );
  AOI21_X1 U11619 ( .B1(n14205), .B2(n9208), .A(n9168), .ZN(n9177) );
  NAND2_X1 U11620 ( .A1(n14205), .A2(n9173), .ZN(n9170) );
  NAND2_X1 U11621 ( .A1(n14026), .A2(n9208), .ZN(n9169) );
  NAND2_X1 U11622 ( .A1(n9170), .A2(n9169), .ZN(n9176) );
  NAND2_X1 U11623 ( .A1(n9177), .A2(n9176), .ZN(n9171) );
  AND2_X1 U11624 ( .A1(n14028), .A2(n9208), .ZN(n9172) );
  AOI21_X1 U11625 ( .B1(n14196), .B2(n9173), .A(n9172), .ZN(n9220) );
  NAND2_X1 U11626 ( .A1(n14196), .A2(n7523), .ZN(n9175) );
  NAND2_X1 U11627 ( .A1(n14028), .A2(n9173), .ZN(n9174) );
  NAND2_X1 U11628 ( .A1(n9175), .A2(n9174), .ZN(n9219) );
  NAND2_X1 U11629 ( .A1(n9220), .A2(n9219), .ZN(n9187) );
  INV_X1 U11630 ( .A(n9176), .ZN(n9179) );
  INV_X1 U11631 ( .A(n9177), .ZN(n9178) );
  AND2_X1 U11632 ( .A1(n9179), .A2(n9178), .ZN(n9184) );
  INV_X1 U11633 ( .A(n9180), .ZN(n9183) );
  INV_X1 U11634 ( .A(n9181), .ZN(n9182) );
  AOI22_X1 U11635 ( .A1(n9185), .A2(n9184), .B1(n9183), .B2(n9182), .ZN(n9186)
         );
  NAND2_X1 U11636 ( .A1(n9189), .A2(n9188), .ZN(n9192) );
  NAND2_X1 U11637 ( .A1(n9190), .A2(n13753), .ZN(n9191) );
  MUX2_X1 U11638 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7274), .Z(n9193) );
  XNOR2_X1 U11639 ( .A(n9193), .B(SI_30_), .ZN(n9232) );
  NAND2_X1 U11640 ( .A1(n9193), .A2(SI_30_), .ZN(n9194) );
  OAI21_X1 U11641 ( .B1(n9234), .B2(n9232), .A(n9194), .ZN(n9197) );
  MUX2_X1 U11642 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7274), .Z(n9195) );
  XNOR2_X1 U11643 ( .A(n9195), .B(SI_31_), .ZN(n9196) );
  NAND2_X1 U11644 ( .A1(n14298), .A2(n9235), .ZN(n9200) );
  INV_X1 U11645 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9198) );
  OR2_X1 U11646 ( .A1(n6847), .A2(n9198), .ZN(n9199) );
  INV_X1 U11647 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14263) );
  NAND2_X1 U11648 ( .A1(n8738), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U11649 ( .A1(n9201), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9202) );
  OAI211_X1 U11650 ( .C1(n9204), .C2(n14263), .A(n9203), .B(n9202), .ZN(n13963) );
  NAND2_X1 U11651 ( .A1(n9230), .A2(n13963), .ZN(n9206) );
  AND2_X1 U11652 ( .A1(n13891), .A2(n9173), .ZN(n9207) );
  AOI21_X1 U11653 ( .B1(n14179), .B2(n9208), .A(n9207), .ZN(n9246) );
  NAND2_X1 U11654 ( .A1(n14179), .A2(n9173), .ZN(n9210) );
  NAND2_X1 U11655 ( .A1(n13891), .A2(n9208), .ZN(n9209) );
  NAND2_X1 U11656 ( .A1(n9210), .A2(n9209), .ZN(n9245) );
  NAND2_X1 U11657 ( .A1(n9246), .A2(n9245), .ZN(n9211) );
  AND2_X1 U11658 ( .A1(n13892), .A2(n9173), .ZN(n9212) );
  AOI21_X1 U11659 ( .B1(n14270), .B2(n9208), .A(n9212), .ZN(n9227) );
  NAND2_X1 U11660 ( .A1(n14270), .A2(n9173), .ZN(n9214) );
  NAND2_X1 U11661 ( .A1(n13892), .A2(n9208), .ZN(n9213) );
  NAND2_X1 U11662 ( .A1(n9214), .A2(n9213), .ZN(n9226) );
  AND2_X1 U11663 ( .A1(n9227), .A2(n9226), .ZN(n9215) );
  AND2_X1 U11664 ( .A1(n13893), .A2(n9173), .ZN(n9216) );
  AOI21_X1 U11665 ( .B1(n14189), .B2(n7523), .A(n9216), .ZN(n9251) );
  NAND2_X1 U11666 ( .A1(n14189), .A2(n9173), .ZN(n9218) );
  NAND2_X1 U11667 ( .A1(n13893), .A2(n7523), .ZN(n9217) );
  NAND2_X1 U11668 ( .A1(n9218), .A2(n9217), .ZN(n9252) );
  INV_X1 U11669 ( .A(n9219), .ZN(n9222) );
  INV_X1 U11670 ( .A(n9220), .ZN(n9221) );
  AOI22_X1 U11671 ( .A1(n9251), .A2(n9252), .B1(n9222), .B2(n9221), .ZN(n9223)
         );
  INV_X1 U11672 ( .A(n9225), .ZN(n9250) );
  INV_X1 U11673 ( .A(n9226), .ZN(n9229) );
  INV_X1 U11674 ( .A(n9227), .ZN(n9228) );
  AND2_X1 U11675 ( .A1(n9229), .A2(n9228), .ZN(n9249) );
  NAND2_X1 U11676 ( .A1(n6792), .A2(n9173), .ZN(n9231) );
  OAI211_X1 U11677 ( .C1(n9205), .C2(n9265), .A(n9263), .B(n9231), .ZN(n9248)
         );
  INV_X1 U11678 ( .A(n9232), .ZN(n9233) );
  NAND2_X1 U11679 ( .A1(n12457), .A2(n9235), .ZN(n9238) );
  INV_X1 U11680 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12036) );
  OR2_X1 U11681 ( .A1(n6847), .A2(n12036), .ZN(n9237) );
  NAND2_X1 U11682 ( .A1(n9173), .A2(n13963), .ZN(n9264) );
  NAND2_X1 U11683 ( .A1(n10146), .A2(n8938), .ZN(n9271) );
  AND2_X1 U11684 ( .A1(n9928), .A2(n6585), .ZN(n9239) );
  AND2_X1 U11685 ( .A1(n9271), .A2(n9239), .ZN(n9241) );
  AOI21_X1 U11686 ( .B1(n9264), .B2(n9241), .A(n9240), .ZN(n9242) );
  AOI21_X1 U11687 ( .B1(n14266), .B2(n9208), .A(n9242), .ZN(n9260) );
  NAND2_X1 U11688 ( .A1(n14266), .A2(n9173), .ZN(n9244) );
  NAND2_X1 U11689 ( .A1(n9208), .A2(n13890), .ZN(n9243) );
  NAND2_X1 U11690 ( .A1(n9244), .A2(n9243), .ZN(n9259) );
  OAI22_X1 U11691 ( .A1(n9260), .A2(n9259), .B1(n9246), .B2(n9245), .ZN(n9247)
         );
  AOI22_X1 U11692 ( .A1(n9250), .A2(n9249), .B1(n9248), .B2(n9247), .ZN(n9257)
         );
  INV_X1 U11693 ( .A(n9251), .ZN(n9254) );
  INV_X1 U11694 ( .A(n9252), .ZN(n9253) );
  NAND3_X1 U11695 ( .A1(n9255), .A2(n9254), .A3(n9253), .ZN(n9256) );
  AND2_X1 U11696 ( .A1(n9257), .A2(n9256), .ZN(n9258) );
  NAND2_X1 U11697 ( .A1(n9260), .A2(n9259), .ZN(n9261) );
  NAND2_X1 U11698 ( .A1(n9262), .A2(n9261), .ZN(n9267) );
  OAI211_X1 U11699 ( .C1(n14264), .C2(n9265), .A(n9264), .B(n9263), .ZN(n9266)
         );
  NAND2_X1 U11700 ( .A1(n6585), .A2(n11795), .ZN(n9268) );
  OAI211_X1 U11701 ( .C1(n9898), .C2(n8938), .A(n9268), .B(n9928), .ZN(n9269)
         );
  INV_X1 U11702 ( .A(n9269), .ZN(n9270) );
  OAI21_X1 U11703 ( .B1(n9272), .B2(n11795), .A(n9271), .ZN(n9273) );
  INV_X1 U11704 ( .A(n9275), .ZN(n9301) );
  INV_X1 U11705 ( .A(n9276), .ZN(n9296) );
  XOR2_X1 U11706 ( .A(n13890), .B(n14266), .Z(n9295) );
  NAND2_X1 U11707 ( .A1(n9278), .A2(n9277), .ZN(n14015) );
  OR2_X1 U11708 ( .A1(n9026), .A2(n10143), .ZN(n9279) );
  AND2_X1 U11709 ( .A1(n9279), .A2(n9902), .ZN(n15357) );
  NOR3_X1 U11710 ( .A1(n15357), .A2(n11104), .A3(n10040), .ZN(n9281) );
  NAND4_X1 U11711 ( .A1(n10666), .A2(n9281), .A3(n9280), .A4(n9949), .ZN(n9282) );
  NOR4_X1 U11712 ( .A1(n10610), .A2(n10546), .A3(n10681), .A4(n9282), .ZN(
        n9284) );
  NAND4_X1 U11713 ( .A1(n9285), .A2(n9284), .A3(n9283), .A4(n10695), .ZN(n9286) );
  NOR4_X1 U11714 ( .A1(n11183), .A2(n10981), .A3(n15134), .A4(n9286), .ZN(
        n9287) );
  XNOR2_X1 U11715 ( .A(n15119), .B(n13904), .ZN(n15117) );
  NAND4_X1 U11716 ( .A1(n11629), .A2(n9287), .A3(n11513), .A4(n15117), .ZN(
        n9288) );
  NOR4_X1 U11717 ( .A1(n14111), .A2(n14142), .A3(n11703), .A4(n9288), .ZN(
        n9289) );
  XNOR2_X1 U11718 ( .A(n14233), .B(n13899), .ZN(n14131) );
  NAND4_X1 U11719 ( .A1(n14082), .A2(n9289), .A3(n14094), .A4(n14131), .ZN(
        n9290) );
  NOR4_X1 U11720 ( .A1(n14015), .A2(n14068), .A3(n9291), .A4(n9290), .ZN(n9292) );
  NAND4_X1 U11721 ( .A1(n13977), .A2(n9292), .A3(n14003), .A4(n14023), .ZN(
        n9293) );
  NOR4_X1 U11722 ( .A1(n9296), .A2(n9295), .A3(n9294), .A4(n9293), .ZN(n9298)
         );
  XNOR2_X1 U11723 ( .A(n9298), .B(n9297), .ZN(n9299) );
  NOR2_X1 U11724 ( .A1(n9933), .A2(P2_U3088), .ZN(n9303) );
  INV_X1 U11725 ( .A(n15352), .ZN(n15349) );
  NOR4_X1 U11726 ( .A1(n15349), .A2(n15096), .A3(n8980), .A4(n9928), .ZN(n9305) );
  INV_X1 U11727 ( .A(n9303), .ZN(n11576) );
  OAI21_X1 U11728 ( .B1(n11576), .B2(n8938), .A(P2_B_REG_SCAN_IN), .ZN(n9304)
         );
  OR2_X1 U11729 ( .A1(n9305), .A2(n9304), .ZN(n9306) );
  NAND2_X1 U11730 ( .A1(n9307), .A2(n9306), .ZN(P2_U3328) );
  INV_X1 U11731 ( .A(n9308), .ZN(n9309) );
  NOR2_X1 U11732 ( .A1(n9934), .A2(n9309), .ZN(P2_U3947) );
  NOR2_X1 U11733 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), 
        .ZN(n9310) );
  NOR2_X2 U11734 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n10255) );
  NOR2_X1 U11735 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .ZN(n9311) );
  INV_X2 U11736 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9419) );
  INV_X1 U11737 ( .A(n9447), .ZN(n9313) );
  NAND4_X2 U11738 ( .A1(n9314), .A2(n9315), .A3(n9313), .A4(n10257), .ZN(n9527) );
  NOR2_X2 U11739 ( .A1(n9527), .A2(n9520), .ZN(n9717) );
  AND2_X2 U11740 ( .A1(n9324), .A2(n9326), .ZN(n9319) );
  NAND2_X1 U11741 ( .A1(n9321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9317) );
  INV_X1 U11742 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9318) );
  OAI21_X2 U11743 ( .B1(n9321), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9322) );
  INV_X1 U11744 ( .A(n9324), .ZN(n9325) );
  NAND2_X1 U11745 ( .A1(n9325), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9327) );
  INV_X2 U11746 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U11747 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9329) );
  MUX2_X1 U11748 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9329), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9332) );
  INV_X1 U11749 ( .A(n9358), .ZN(n9331) );
  NAND2_X1 U11750 ( .A1(n9332), .A2(n9331), .ZN(n14484) );
  AND2_X1 U11751 ( .A1(n7620), .A2(P1_U3086), .ZN(n11574) );
  INV_X2 U11752 ( .A(n11574), .ZN(n15030) );
  INV_X1 U11753 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9753) );
  OAI222_X1 U11754 ( .A1(P1_U3086), .A2(n14484), .B1(n15030), .B2(n9752), .C1(
        n9753), .C2(n15024), .ZN(P1_U3354) );
  NOR2_X2 U11755 ( .A1(n7274), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13749) );
  OAI222_X1 U11756 ( .A1(P3_U3151), .A2(n10196), .B1(n12609), .B2(n9334), .C1(
        n13756), .C2(n9333), .ZN(P3_U3294) );
  INV_X1 U11757 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9335) );
  AND2_X1 U11758 ( .A1(n9358), .A2(n9335), .ZN(n9360) );
  INV_X1 U11759 ( .A(n9360), .ZN(n9352) );
  OR2_X1 U11760 ( .A1(n9352), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9347) );
  INV_X1 U11761 ( .A(n9347), .ZN(n9337) );
  INV_X1 U11762 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U11763 ( .A1(n9337), .A2(n9336), .ZN(n9349) );
  NAND2_X1 U11764 ( .A1(n9349), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9338) );
  MUX2_X1 U11765 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9338), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9339) );
  AND2_X1 U11766 ( .A1(n9520), .A2(n9339), .ZN(n10101) );
  INV_X1 U11767 ( .A(n10101), .ZN(n9341) );
  OAI222_X1 U11768 ( .A1(P1_U3086), .A2(n9341), .B1(n15030), .B2(n10100), .C1(
        n9340), .C2(n15024), .ZN(P1_U3350) );
  NOR2_X1 U11769 ( .A1(n7274), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14304) );
  AND2_X1 U11770 ( .A1(n7274), .A2(P2_U3088), .ZN(n14306) );
  INV_X2 U11771 ( .A(n14306), .ZN(n10596) );
  OAI222_X1 U11772 ( .A1(n14312), .A2(n9342), .B1(n9463), .B2(P2_U3088), .C1(
        n10596), .C2(n9752), .ZN(P2_U3326) );
  OAI222_X1 U11773 ( .A1(n10184), .A2(P3_U3151), .B1(n13756), .B2(n9343), .C1(
        n9760), .C2(n12609), .ZN(P3_U3295) );
  OAI222_X1 U11774 ( .A1(P3_U3151), .A2(n11254), .B1(n12609), .B2(n9345), .C1(
        n13756), .C2(n9344), .ZN(P3_U3287) );
  AOI22_X1 U11775 ( .A1(n9506), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n14304), .ZN(n9346) );
  OAI21_X1 U11776 ( .B1(n10402), .B2(n10596), .A(n9346), .ZN(P2_U3321) );
  INV_X1 U11777 ( .A(n15024), .ZN(n15015) );
  INV_X1 U11778 ( .A(n10011), .ZN(n9363) );
  NAND2_X1 U11779 ( .A1(n9347), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9348) );
  MUX2_X1 U11780 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9348), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9350) );
  NAND2_X1 U11781 ( .A1(n9350), .A2(n9349), .ZN(n14525) );
  OAI222_X1 U11782 ( .A1(n15024), .A2(n9351), .B1(n15030), .B2(n9363), .C1(
        n14525), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U11783 ( .A(n10005), .ZN(n9366) );
  NAND2_X1 U11784 ( .A1(n9352), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9353) );
  XNOR2_X1 U11785 ( .A(n9353), .B(P1_IR_REG_3__SCAN_IN), .ZN(n14515) );
  INV_X1 U11786 ( .A(n14515), .ZN(n9354) );
  OAI222_X1 U11787 ( .A1(n15024), .A2(n9355), .B1(n15030), .B2(n9366), .C1(
        n9354), .C2(P1_U3086), .ZN(P1_U3352) );
  OR2_X1 U11788 ( .A1(n10260), .A2(n9318), .ZN(n9356) );
  XNOR2_X1 U11789 ( .A(n9356), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10403) );
  INV_X1 U11790 ( .A(n10403), .ZN(n9630) );
  OAI222_X1 U11791 ( .A1(P1_U3086), .A2(n9630), .B1(n15030), .B2(n10402), .C1(
        n9357), .C2(n15024), .ZN(P1_U3349) );
  NOR2_X1 U11792 ( .A1(n9358), .A2(n9318), .ZN(n9359) );
  MUX2_X1 U11793 ( .A(n9318), .B(n9359), .S(P1_IR_REG_2__SCAN_IN), .Z(n9361)
         );
  NOR2_X1 U11794 ( .A1(n9361), .A2(n9360), .ZN(n9792) );
  INV_X1 U11795 ( .A(n9792), .ZN(n14504) );
  OAI222_X1 U11796 ( .A1(P1_U3086), .A2(n14504), .B1(n15030), .B2(n9791), .C1(
        n9362), .C2(n15024), .ZN(P1_U3353) );
  OAI222_X1 U11797 ( .A1(n14312), .A2(n9364), .B1(n10596), .B2(n9363), .C1(
        P2_U3088), .C2(n9608), .ZN(P2_U3323) );
  INV_X1 U11798 ( .A(n9490), .ZN(n9621) );
  OAI222_X1 U11799 ( .A1(n14312), .A2(n9365), .B1(n9621), .B2(P2_U3088), .C1(
        n10596), .C2(n10100), .ZN(P2_U3322) );
  INV_X1 U11800 ( .A(n9484), .ZN(n15276) );
  OAI222_X1 U11801 ( .A1(n14312), .A2(n9367), .B1(n10596), .B2(n9366), .C1(
        P2_U3088), .C2(n15276), .ZN(P2_U3324) );
  OAI222_X1 U11802 ( .A1(n14312), .A2(n9368), .B1(n9480), .B2(P2_U3088), .C1(
        n10596), .C2(n9791), .ZN(P2_U3325) );
  INV_X1 U11803 ( .A(n12609), .ZN(n9883) );
  AOI222_X1 U11804 ( .A1(n9369), .A2(n13749), .B1(SI_5_), .B2(n9883), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n10307), .ZN(n9370) );
  INV_X1 U11805 ( .A(n9370), .ZN(P3_U3290) );
  AOI222_X1 U11806 ( .A1(n9371), .A2(n13749), .B1(SI_7_), .B2(n9883), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n11251), .ZN(n9372) );
  INV_X1 U11807 ( .A(n9372), .ZN(P3_U3288) );
  AOI222_X1 U11808 ( .A1(n9373), .A2(n13749), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10252), .C1(SI_2_), .C2(n9883), .ZN(n9374) );
  INV_X1 U11809 ( .A(n9374), .ZN(P3_U3293) );
  AOI222_X1 U11810 ( .A1(n9375), .A2(n13749), .B1(n6753), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n9883), .ZN(n9376) );
  INV_X1 U11811 ( .A(n9376), .ZN(P3_U3291) );
  AOI222_X1 U11812 ( .A1(n9377), .A2(n13749), .B1(SI_9_), .B2(n9883), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n11374), .ZN(n9378) );
  INV_X1 U11813 ( .A(n9378), .ZN(P3_U3286) );
  OAI222_X1 U11814 ( .A1(P3_U3151), .A2(n11093), .B1(n12609), .B2(n9380), .C1(
        n13756), .C2(n9379), .ZN(P3_U3289) );
  INV_X1 U11815 ( .A(n9381), .ZN(n9383) );
  INV_X1 U11816 ( .A(SI_3_), .ZN(n9382) );
  OAI222_X1 U11817 ( .A1(n13756), .A2(n9383), .B1(n12609), .B2(n9382), .C1(
        P3_U3151), .C2(n10224), .ZN(P3_U3292) );
  INV_X1 U11818 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U11819 ( .A1(n10260), .A2(n9384), .ZN(n9385) );
  NAND2_X1 U11820 ( .A1(n9385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9389) );
  XNOR2_X1 U11821 ( .A(n9389), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14552) );
  INV_X1 U11822 ( .A(n14552), .ZN(n14543) );
  OAI222_X1 U11823 ( .A1(P1_U3086), .A2(n14543), .B1(n15030), .B2(n10454), 
        .C1(n9386), .C2(n15024), .ZN(P1_U3348) );
  INV_X1 U11824 ( .A(n9586), .ZN(n9515) );
  OAI222_X1 U11825 ( .A1(n14312), .A2(n9387), .B1(n9515), .B2(P2_U3088), .C1(
        n10596), .C2(n10454), .ZN(P2_U3320) );
  INV_X1 U11826 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9388) );
  NAND2_X1 U11827 ( .A1(n9389), .A2(n9388), .ZN(n9390) );
  NAND2_X1 U11828 ( .A1(n9390), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9449) );
  XNOR2_X1 U11829 ( .A(n9449), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10571) );
  INV_X1 U11830 ( .A(n10571), .ZN(n9645) );
  OAI222_X1 U11831 ( .A1(n15024), .A2(n9391), .B1(n15030), .B2(n10570), .C1(
        P1_U3086), .C2(n9645), .ZN(P1_U3347) );
  INV_X1 U11832 ( .A(n9861), .ZN(n9595) );
  OAI222_X1 U11833 ( .A1(n14312), .A2(n9392), .B1(n9595), .B2(P2_U3088), .C1(
        n10596), .C2(n10570), .ZN(P2_U3319) );
  OAI222_X1 U11834 ( .A1(n13756), .A2(n9393), .B1(n11764), .B2(P3_U3151), .C1(
        n13401), .C2(n12609), .ZN(P3_U3284) );
  AOI222_X1 U11835 ( .A1(n9394), .A2(n13749), .B1(SI_10_), .B2(n9883), .C1(
        P3_STATE_REG_SCAN_IN), .C2(n11383), .ZN(n9395) );
  INV_X1 U11836 ( .A(n9395), .ZN(P3_U3285) );
  NAND3_X1 U11837 ( .A1(n11725), .A2(P1_B_REG_SCAN_IN), .A3(n9397), .ZN(n9398)
         );
  INV_X1 U11838 ( .A(n9738), .ZN(n9399) );
  INV_X1 U11839 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9402) );
  NOR3_X1 U11840 ( .A1(n9733), .A2(n9400), .A3(n9403), .ZN(n9401) );
  AOI21_X1 U11841 ( .B1(n15224), .B2(n9402), .A(n9401), .ZN(P1_U3445) );
  INV_X1 U11842 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9406) );
  NOR3_X1 U11843 ( .A1(n9733), .A2(n9404), .A3(n9403), .ZN(n9405) );
  AOI21_X1 U11844 ( .B1(n15224), .B2(n9406), .A(n9405), .ZN(P1_U3446) );
  NAND2_X1 U11845 ( .A1(n9449), .A2(n9407), .ZN(n9408) );
  NAND2_X1 U11846 ( .A1(n9408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9420) );
  XNOR2_X1 U11847 ( .A(n9420), .B(P1_IR_REG_9__SCAN_IN), .ZN(n14572) );
  INV_X1 U11848 ( .A(n14572), .ZN(n9410) );
  OAI222_X1 U11849 ( .A1(P1_U3086), .A2(n9410), .B1(n15030), .B2(n10726), .C1(
        n9409), .C2(n15024), .ZN(P1_U3346) );
  INV_X1 U11850 ( .A(n13925), .ZN(n9411) );
  OAI222_X1 U11851 ( .A1(n14312), .A2(n9412), .B1(n9411), .B2(P2_U3088), .C1(
        n10596), .C2(n10726), .ZN(P2_U3318) );
  NAND2_X1 U11852 ( .A1(n10482), .A2(n9990), .ZN(n9413) );
  OAI21_X1 U11853 ( .B1(n9990), .B2(n9414), .A(n9413), .ZN(P3_U3377) );
  AOI222_X1 U11854 ( .A1(n9415), .A2(n13749), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11770), .C1(SI_12_), .C2(n9883), .ZN(n9416) );
  INV_X1 U11855 ( .A(n9416), .ZN(P3_U3283) );
  NAND2_X1 U11856 ( .A1(n6589), .A2(n11414), .ZN(n9417) );
  OAI21_X1 U11857 ( .B1(n6589), .B2(n7971), .A(n9417), .ZN(P2_U3544) );
  INV_X1 U11858 ( .A(n11107), .ZN(n9423) );
  INV_X1 U11859 ( .A(n10060), .ZN(n10054) );
  OAI222_X1 U11860 ( .A1(n14312), .A2(n9418), .B1(n10596), .B2(n9423), .C1(
        P2_U3088), .C2(n10054), .ZN(P2_U3317) );
  NAND2_X1 U11861 ( .A1(n9420), .A2(n9419), .ZN(n9421) );
  NAND2_X1 U11862 ( .A1(n9421), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9422) );
  XNOR2_X1 U11863 ( .A(n9422), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11108) );
  INV_X1 U11864 ( .A(n11108), .ZN(n9660) );
  OAI222_X1 U11865 ( .A1(n15024), .A2(n9424), .B1(n15030), .B2(n9423), .C1(
        n9660), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U11866 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n14165) );
  NAND3_X1 U11867 ( .A1(n9430), .A2(P2_REG2_REG_0__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n9457) );
  INV_X1 U11868 ( .A(n9457), .ZN(n9446) );
  INV_X1 U11869 ( .A(n9933), .ZN(n9428) );
  NAND2_X1 U11870 ( .A1(n9921), .A2(n9933), .ZN(n9426) );
  NAND2_X1 U11871 ( .A1(n9426), .A2(n9425), .ZN(n9427) );
  OR2_X1 U11872 ( .A1(n9439), .A2(P2_U3088), .ZN(n14308) );
  NOR2_X1 U11873 ( .A1(n8980), .A2(n14308), .ZN(n9429) );
  AND2_X1 U11874 ( .A1(n9441), .A2(n9429), .ZN(n15319) );
  INV_X1 U11875 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10151) );
  NOR2_X1 U11876 ( .A1(n15281), .A2(n10151), .ZN(n15268) );
  AOI22_X1 U11877 ( .A1(n15268), .A2(P2_IR_REG_0__SCAN_IN), .B1(n15319), .B2(
        n9430), .ZN(n9445) );
  INV_X1 U11878 ( .A(n14308), .ZN(n9431) );
  AND2_X1 U11879 ( .A1(n9431), .A2(n8980), .ZN(n9432) );
  NAND2_X1 U11880 ( .A1(n9441), .A2(n9432), .ZN(n15269) );
  INV_X1 U11881 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15394) );
  INV_X1 U11882 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9434) );
  INV_X1 U11883 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n13426) );
  MUX2_X1 U11884 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n13426), .S(n9463), .Z(n9433) );
  OAI21_X1 U11885 ( .B1(n15394), .B2(n9434), .A(n9433), .ZN(n9437) );
  MUX2_X1 U11886 ( .A(n13426), .B(P2_REG1_REG_1__SCAN_IN), .S(n9463), .Z(n9436) );
  AND2_X1 U11887 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9435) );
  NAND2_X1 U11888 ( .A1(n9436), .A2(n9435), .ZN(n9462) );
  NAND2_X1 U11889 ( .A1(n9437), .A2(n9462), .ZN(n9438) );
  NOR2_X1 U11890 ( .A1(n15269), .A2(n9438), .ZN(n9443) );
  AND2_X1 U11891 ( .A1(n9439), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9440) );
  OR2_X1 U11892 ( .A1(n9441), .A2(P2_U3088), .ZN(n11798) );
  OAI22_X1 U11893 ( .A1(n15311), .A2(n9463), .B1(n11798), .B2(n7712), .ZN(
        n9442) );
  AOI211_X1 U11894 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(P2_U3088), .A(n9443), 
        .B(n9442), .ZN(n9444) );
  OAI21_X1 U11895 ( .B1(n9446), .B2(n9445), .A(n9444), .ZN(P2_U3215) );
  INV_X1 U11896 ( .A(n11138), .ZN(n9452) );
  NAND2_X1 U11897 ( .A1(n10258), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9448) );
  NAND2_X1 U11898 ( .A1(n9449), .A2(n9448), .ZN(n9670) );
  INV_X1 U11899 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9450) );
  XNOR2_X1 U11900 ( .A(n9670), .B(n9450), .ZN(n11139) );
  INV_X1 U11901 ( .A(n11139), .ZN(n9692) );
  OAI222_X1 U11902 ( .A1(n15024), .A2(n9451), .B1(n15030), .B2(n9452), .C1(
        P1_U3086), .C2(n9692), .ZN(P1_U3344) );
  INV_X1 U11903 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9453) );
  INV_X1 U11904 ( .A(n13942), .ZN(n13939) );
  OAI222_X1 U11905 ( .A1(n14312), .A2(n9453), .B1(n10596), .B2(n9452), .C1(
        P2_U3088), .C2(n13939), .ZN(P2_U3316) );
  INV_X1 U11906 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n9468) );
  NOR2_X1 U11907 ( .A1(n15311), .A2(n9480), .ZN(n9460) );
  INV_X1 U11908 ( .A(n9463), .ZN(n9454) );
  NAND2_X1 U11909 ( .A1(n9454), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9456) );
  INV_X1 U11910 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n13398) );
  MUX2_X1 U11911 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n13398), .S(n9480), .Z(n9455) );
  AOI21_X1 U11912 ( .B1(n9457), .B2(n9456), .A(n9455), .ZN(n9469) );
  AND3_X1 U11913 ( .A1(n9457), .A2(n9456), .A3(n9455), .ZN(n9458) );
  NOR3_X1 U11914 ( .A1(n15281), .A2(n9469), .A3(n9458), .ZN(n9459) );
  AOI211_X1 U11915 ( .C1(P2_REG3_REG_2__SCAN_IN), .C2(P2_U3088), .A(n9460), 
        .B(n9459), .ZN(n9467) );
  INV_X1 U11916 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9461) );
  MUX2_X1 U11917 ( .A(n9461), .B(P2_REG1_REG_2__SCAN_IN), .S(n9480), .Z(n9465)
         );
  OAI21_X1 U11918 ( .B1(n13426), .B2(n9463), .A(n9462), .ZN(n9464) );
  INV_X1 U11919 ( .A(n15269), .ZN(n15317) );
  NAND2_X1 U11920 ( .A1(n9465), .A2(n9464), .ZN(n9482) );
  OAI211_X1 U11921 ( .C1(n9465), .C2(n9464), .A(n15317), .B(n9482), .ZN(n9466)
         );
  OAI211_X1 U11922 ( .C1(n9468), .C2(n11798), .A(n9467), .B(n9466), .ZN(
        P2_U3216) );
  NAND2_X1 U11923 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n10560) );
  INV_X1 U11924 ( .A(n10560), .ZN(n9479) );
  INV_X1 U11925 ( .A(n9480), .ZN(n9470) );
  INV_X1 U11926 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9471) );
  MUX2_X1 U11927 ( .A(n9471), .B(P2_REG2_REG_3__SCAN_IN), .S(n9484), .Z(n15283) );
  NOR2_X1 U11928 ( .A1(n15284), .A2(n15283), .ZN(n15282) );
  INV_X1 U11929 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9472) );
  MUX2_X1 U11930 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9472), .S(n9608), .Z(n9597)
         );
  NOR2_X1 U11931 ( .A1(n9598), .A2(n9597), .ZN(n9596) );
  AOI21_X1 U11932 ( .B1(n9487), .B2(P2_REG2_REG_4__SCAN_IN), .A(n9596), .ZN(
        n9614) );
  INV_X1 U11933 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9473) );
  MUX2_X1 U11934 ( .A(n9473), .B(P2_REG2_REG_5__SCAN_IN), .S(n9490), .Z(n9613)
         );
  NOR2_X1 U11935 ( .A1(n9614), .A2(n9613), .ZN(n9612) );
  NOR2_X1 U11936 ( .A1(n9621), .A2(n9473), .ZN(n9475) );
  INV_X1 U11937 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10653) );
  MUX2_X1 U11938 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10653), .S(n9506), .Z(n9474) );
  INV_X1 U11939 ( .A(n9502), .ZN(n9477) );
  NOR3_X1 U11940 ( .A1(n9612), .A2(n9475), .A3(n9474), .ZN(n9476) );
  NOR3_X1 U11941 ( .A1(n9477), .A2(n9476), .A3(n15281), .ZN(n9478) );
  AOI211_X1 U11942 ( .C1(n15300), .C2(n9506), .A(n9479), .B(n9478), .ZN(n9498)
         );
  OR2_X1 U11943 ( .A1(n9480), .A2(n9461), .ZN(n9481) );
  NAND2_X1 U11944 ( .A1(n9482), .A2(n9481), .ZN(n15280) );
  INV_X1 U11945 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9483) );
  MUX2_X1 U11946 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9483), .S(n9484), .Z(n15279) );
  NAND2_X1 U11947 ( .A1(n15280), .A2(n15279), .ZN(n15278) );
  NAND2_X1 U11948 ( .A1(n9484), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9485) );
  NAND2_X1 U11949 ( .A1(n15278), .A2(n9485), .ZN(n9602) );
  INV_X1 U11950 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9486) );
  MUX2_X1 U11951 ( .A(n9486), .B(P2_REG1_REG_4__SCAN_IN), .S(n9608), .Z(n9601)
         );
  NAND2_X1 U11952 ( .A1(n9602), .A2(n9601), .ZN(n9600) );
  NAND2_X1 U11953 ( .A1(n9487), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9488) );
  NAND2_X1 U11954 ( .A1(n9600), .A2(n9488), .ZN(n9611) );
  INV_X1 U11955 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9489) );
  MUX2_X1 U11956 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9489), .S(n9490), .Z(n9610)
         );
  NAND2_X1 U11957 ( .A1(n9611), .A2(n9610), .ZN(n9609) );
  NAND2_X1 U11958 ( .A1(n9490), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U11959 ( .A1(n9609), .A2(n9495), .ZN(n9493) );
  INV_X1 U11960 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9491) );
  MUX2_X1 U11961 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9491), .S(n9506), .Z(n9492)
         );
  NAND2_X1 U11962 ( .A1(n9493), .A2(n9492), .ZN(n9510) );
  MUX2_X1 U11963 ( .A(n9491), .B(P2_REG1_REG_6__SCAN_IN), .S(n9506), .Z(n9494)
         );
  NAND3_X1 U11964 ( .A1(n9609), .A2(n9495), .A3(n9494), .ZN(n9496) );
  NAND3_X1 U11965 ( .A1(n15317), .A2(n9510), .A3(n9496), .ZN(n9497) );
  OAI211_X1 U11966 ( .C1(n7724), .C2(n11798), .A(n9498), .B(n9497), .ZN(
        P2_U3220) );
  INV_X1 U11967 ( .A(n11798), .ZN(n15314) );
  NAND2_X1 U11968 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10394) );
  INV_X1 U11969 ( .A(n10394), .ZN(n9505) );
  NAND2_X1 U11970 ( .A1(n9506), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9501) );
  INV_X1 U11971 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9499) );
  MUX2_X1 U11972 ( .A(n9499), .B(P2_REG2_REG_7__SCAN_IN), .S(n9586), .Z(n9500)
         );
  AOI21_X1 U11973 ( .B1(n9502), .B2(n9501), .A(n9500), .ZN(n9580) );
  AND3_X1 U11974 ( .A1(n9502), .A2(n9501), .A3(n9500), .ZN(n9503) );
  NOR3_X1 U11975 ( .A1(n9580), .A2(n9503), .A3(n15281), .ZN(n9504) );
  AOI211_X1 U11976 ( .C1(n15314), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n9505), .B(
        n9504), .ZN(n9514) );
  NAND2_X1 U11977 ( .A1(n9506), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9509) );
  INV_X1 U11978 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9507) );
  MUX2_X1 U11979 ( .A(n9507), .B(P2_REG1_REG_7__SCAN_IN), .S(n9586), .Z(n9508)
         );
  AOI21_X1 U11980 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9585) );
  INV_X1 U11981 ( .A(n9585), .ZN(n9512) );
  NAND3_X1 U11982 ( .A1(n9510), .A2(n9509), .A3(n9508), .ZN(n9511) );
  NAND3_X1 U11983 ( .A1(n15317), .A2(n9512), .A3(n9511), .ZN(n9513) );
  OAI211_X1 U11984 ( .C1(n15311), .C2(n9515), .A(n9514), .B(n9513), .ZN(
        P2_U3221) );
  OR2_X1 U11985 ( .A1(n9820), .A2(P1_U3086), .ZN(n12531) );
  NAND2_X1 U11986 ( .A1(n9830), .A2(n12531), .ZN(n9558) );
  XNOR2_X2 U11987 ( .A(n9517), .B(P1_IR_REG_22__SCAN_IN), .ZN(n15034) );
  NAND2_X1 U11988 ( .A1(n9518), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9519) );
  INV_X1 U11989 ( .A(n9520), .ZN(n9525) );
  NOR2_X1 U11990 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n9524) );
  NOR2_X1 U11991 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n9523) );
  NOR2_X1 U11992 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9522) );
  NOR2_X1 U11993 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n9521) );
  NAND2_X1 U11994 ( .A1(n9525), .A2(n7635), .ZN(n9526) );
  NAND2_X1 U11995 ( .A1(n9741), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9528) );
  XNOR2_X1 U11996 ( .A(n9528), .B(n9742), .ZN(n9559) );
  AOI21_X1 U11997 ( .B1(n9820), .B2(n12293), .A(n11844), .ZN(n9557) );
  INV_X1 U11998 ( .A(n9557), .ZN(n9531) );
  AND2_X1 U11999 ( .A1(n9558), .A2(n9531), .ZN(n15199) );
  NOR2_X1 U12000 ( .A1(n15199), .A2(n14496), .ZN(P1_U3085) );
  NOR2_X1 U12001 ( .A1(n9532), .A2(n13742), .ZN(n9535) );
  CLKBUF_X1 U12002 ( .A(n9535), .Z(n9556) );
  INV_X1 U12003 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9533) );
  NOR2_X1 U12004 ( .A1(n9556), .A2(n9533), .ZN(P3_U3245) );
  INV_X1 U12005 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9534) );
  NOR2_X1 U12006 ( .A1(n9556), .A2(n9534), .ZN(P3_U3244) );
  INV_X1 U12007 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9536) );
  NOR2_X1 U12008 ( .A1(n9556), .A2(n9536), .ZN(P3_U3248) );
  INV_X1 U12009 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9537) );
  NOR2_X1 U12010 ( .A1(n9556), .A2(n9537), .ZN(P3_U3243) );
  INV_X1 U12011 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n13349) );
  NOR2_X1 U12012 ( .A1(n9535), .A2(n13349), .ZN(P3_U3250) );
  INV_X1 U12013 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9538) );
  NOR2_X1 U12014 ( .A1(n9535), .A2(n9538), .ZN(P3_U3251) );
  INV_X1 U12015 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9539) );
  NOR2_X1 U12016 ( .A1(n9535), .A2(n9539), .ZN(P3_U3252) );
  INV_X1 U12017 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n13402) );
  NOR2_X1 U12018 ( .A1(n9535), .A2(n13402), .ZN(P3_U3253) );
  NOR2_X1 U12019 ( .A1(n9535), .A2(n13473), .ZN(P3_U3246) );
  INV_X1 U12020 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9540) );
  NOR2_X1 U12021 ( .A1(n9535), .A2(n9540), .ZN(P3_U3247) );
  INV_X1 U12022 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9541) );
  NOR2_X1 U12023 ( .A1(n9535), .A2(n9541), .ZN(P3_U3256) );
  INV_X1 U12024 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9542) );
  NOR2_X1 U12025 ( .A1(n9535), .A2(n9542), .ZN(P3_U3257) );
  INV_X1 U12026 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9543) );
  NOR2_X1 U12027 ( .A1(n9556), .A2(n9543), .ZN(P3_U3258) );
  INV_X1 U12028 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n13478) );
  NOR2_X1 U12029 ( .A1(n9535), .A2(n13478), .ZN(P3_U3259) );
  INV_X1 U12030 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9544) );
  NOR2_X1 U12031 ( .A1(n9556), .A2(n9544), .ZN(P3_U3241) );
  INV_X1 U12032 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n13488) );
  NOR2_X1 U12033 ( .A1(n9556), .A2(n13488), .ZN(P3_U3242) );
  INV_X1 U12034 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9545) );
  NOR2_X1 U12035 ( .A1(n9535), .A2(n9545), .ZN(P3_U3262) );
  INV_X1 U12036 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9546) );
  NOR2_X1 U12037 ( .A1(n9556), .A2(n9546), .ZN(P3_U3263) );
  INV_X1 U12038 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9547) );
  NOR2_X1 U12039 ( .A1(n9556), .A2(n9547), .ZN(P3_U3240) );
  NOR2_X1 U12040 ( .A1(n9556), .A2(n13474), .ZN(P3_U3260) );
  INV_X1 U12041 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9548) );
  NOR2_X1 U12042 ( .A1(n9535), .A2(n9548), .ZN(P3_U3261) );
  INV_X1 U12043 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9549) );
  NOR2_X1 U12044 ( .A1(n9556), .A2(n9549), .ZN(P3_U3235) );
  NOR2_X1 U12045 ( .A1(n9556), .A2(n13512), .ZN(P3_U3249) );
  INV_X1 U12046 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9550) );
  NOR2_X1 U12047 ( .A1(n9556), .A2(n9550), .ZN(P3_U3234) );
  INV_X1 U12048 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9551) );
  NOR2_X1 U12049 ( .A1(n9556), .A2(n9551), .ZN(P3_U3254) );
  NOR2_X1 U12050 ( .A1(n9556), .A2(n13391), .ZN(P3_U3236) );
  INV_X1 U12051 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9552) );
  NOR2_X1 U12052 ( .A1(n9556), .A2(n9552), .ZN(P3_U3237) );
  INV_X1 U12053 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9553) );
  NOR2_X1 U12054 ( .A1(n9556), .A2(n9553), .ZN(P3_U3255) );
  INV_X1 U12055 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9554) );
  NOR2_X1 U12056 ( .A1(n9556), .A2(n9554), .ZN(P3_U3239) );
  INV_X1 U12057 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9555) );
  NOR2_X1 U12058 ( .A1(n9556), .A2(n9555), .ZN(P3_U3238) );
  NAND2_X1 U12059 ( .A1(n9558), .A2(n9557), .ZN(n15201) );
  INV_X1 U12060 ( .A(n14490), .ZN(n14494) );
  INV_X1 U12061 ( .A(n14525), .ZN(n10012) );
  INV_X1 U12062 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9769) );
  MUX2_X1 U12063 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9769), .S(n9792), .Z(n14499) );
  INV_X1 U12064 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14479) );
  MUX2_X1 U12065 ( .A(n14479), .B(P1_REG1_REG_1__SCAN_IN), .S(n14484), .Z(
        n9561) );
  AND2_X1 U12066 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9560) );
  NAND2_X1 U12067 ( .A1(n9561), .A2(n9560), .ZN(n14483) );
  OAI21_X1 U12068 ( .B1(n14479), .B2(n14484), .A(n14483), .ZN(n14498) );
  NAND2_X1 U12069 ( .A1(n14499), .A2(n14498), .ZN(n14513) );
  NAND2_X1 U12070 ( .A1(n9792), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n14512) );
  NAND2_X1 U12071 ( .A1(n14513), .A2(n14512), .ZN(n9563) );
  INV_X1 U12072 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9824) );
  MUX2_X1 U12073 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9824), .S(n14515), .Z(n9562) );
  NAND2_X1 U12074 ( .A1(n9563), .A2(n9562), .ZN(n14530) );
  NAND2_X1 U12075 ( .A1(n14515), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n14529) );
  INV_X1 U12076 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n13501) );
  MUX2_X1 U12077 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n13501), .S(n14525), .Z(
        n14528) );
  AOI21_X1 U12078 ( .B1(n14530), .B2(n14529), .A(n14528), .ZN(n14527) );
  AOI21_X1 U12079 ( .B1(n10012), .B2(P1_REG1_REG_4__SCAN_IN), .A(n14527), .ZN(
        n9675) );
  INV_X1 U12080 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15262) );
  MUX2_X1 U12081 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n15262), .S(n10101), .Z(
        n9676) );
  NAND2_X1 U12082 ( .A1(n9675), .A2(n9676), .ZN(n9674) );
  OAI21_X1 U12083 ( .B1(n10101), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9674), .ZN(
        n9565) );
  INV_X1 U12084 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9629) );
  MUX2_X1 U12085 ( .A(n9629), .B(P1_REG1_REG_6__SCAN_IN), .S(n10403), .Z(n9564) );
  NOR2_X1 U12086 ( .A1(n9565), .A2(n9564), .ZN(n14548) );
  INV_X1 U12087 ( .A(n6584), .ZN(n15197) );
  OR2_X1 U12088 ( .A1(n15201), .A2(n15197), .ZN(n15208) );
  AOI211_X1 U12089 ( .C1(n9565), .C2(n9564), .A(n14548), .B(n15208), .ZN(n9575) );
  OR2_X1 U12090 ( .A1(n14490), .A2(n6584), .ZN(n9566) );
  INV_X1 U12091 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10857) );
  MUX2_X1 U12092 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10857), .S(n9792), .Z(
        n14501) );
  INV_X1 U12093 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9567) );
  MUX2_X1 U12094 ( .A(n9567), .B(P1_REG2_REG_1__SCAN_IN), .S(n14484), .Z(
        n14478) );
  AND2_X1 U12095 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14492) );
  NAND2_X1 U12096 ( .A1(n14478), .A2(n14492), .ZN(n14477) );
  OAI21_X1 U12097 ( .B1(n9567), .B2(n14484), .A(n14477), .ZN(n14500) );
  NAND2_X1 U12098 ( .A1(n14501), .A2(n14500), .ZN(n14518) );
  NAND2_X1 U12099 ( .A1(n9792), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14517) );
  NAND2_X1 U12100 ( .A1(n14518), .A2(n14517), .ZN(n9569) );
  INV_X1 U12101 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10848) );
  MUX2_X1 U12102 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10848), .S(n14515), .Z(
        n9568) );
  NAND2_X1 U12103 ( .A1(n9569), .A2(n9568), .ZN(n14536) );
  NAND2_X1 U12104 ( .A1(n14515), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14535) );
  INV_X1 U12105 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9570) );
  MUX2_X1 U12106 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9570), .S(n14525), .Z(
        n14534) );
  AOI21_X1 U12107 ( .B1(n14536), .B2(n14535), .A(n14534), .ZN(n14533) );
  NOR2_X1 U12108 ( .A1(n14525), .A2(n9570), .ZN(n9679) );
  INV_X1 U12109 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11068) );
  MUX2_X1 U12110 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n11068), .S(n10101), .Z(
        n9678) );
  OAI21_X1 U12111 ( .B1(n14533), .B2(n9679), .A(n9678), .ZN(n9677) );
  NAND2_X1 U12112 ( .A1(n10101), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9572) );
  INV_X1 U12113 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9622) );
  MUX2_X1 U12114 ( .A(n9622), .B(P1_REG2_REG_6__SCAN_IN), .S(n10403), .Z(n9571) );
  AOI21_X1 U12115 ( .B1(n9677), .B2(n9572), .A(n9571), .ZN(n14557) );
  AND3_X1 U12116 ( .A1(n9677), .A2(n9572), .A3(n9571), .ZN(n9573) );
  NOR3_X1 U12117 ( .A1(n15210), .A2(n14557), .A3(n9573), .ZN(n9574) );
  NOR2_X1 U12118 ( .A1(n9575), .A2(n9574), .ZN(n9577) );
  AND2_X1 U12119 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14430) );
  AOI21_X1 U12120 ( .B1(n15199), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n14430), .ZN(
        n9576) );
  OAI211_X1 U12121 ( .C1(n9630), .C2(n15212), .A(n9577), .B(n9576), .ZN(
        P1_U3249) );
  OAI222_X1 U12122 ( .A1(n13756), .A2(n9579), .B1(n12609), .B2(n9578), .C1(
        n12932), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U12123 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9581) );
  MUX2_X1 U12124 ( .A(n9581), .B(P2_REG2_REG_8__SCAN_IN), .S(n9861), .Z(n9582)
         );
  NOR2_X1 U12125 ( .A1(n9583), .A2(n9582), .ZN(n9854) );
  AOI211_X1 U12126 ( .C1(n9583), .C2(n9582), .A(n9854), .B(n15281), .ZN(n9584)
         );
  INV_X1 U12127 ( .A(n9584), .ZN(n9591) );
  AOI21_X1 U12128 ( .B1(n9586), .B2(P2_REG1_REG_7__SCAN_IN), .A(n9585), .ZN(
        n9588) );
  INV_X1 U12129 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n15398) );
  MUX2_X1 U12130 ( .A(n15398), .B(P2_REG1_REG_8__SCAN_IN), .S(n9861), .Z(n9587) );
  NOR2_X1 U12131 ( .A1(n9588), .A2(n9587), .ZN(n9860) );
  AOI211_X1 U12132 ( .C1(n9588), .C2(n9587), .A(n9860), .B(n15269), .ZN(n9589)
         );
  INV_X1 U12133 ( .A(n9589), .ZN(n9590) );
  NAND2_X1 U12134 ( .A1(n9591), .A2(n9590), .ZN(n9593) );
  NAND2_X1 U12135 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n10643) );
  INV_X1 U12136 ( .A(n10643), .ZN(n9592) );
  AOI211_X1 U12137 ( .C1(n15314), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n9593), .B(
        n9592), .ZN(n9594) );
  OAI21_X1 U12138 ( .B1(n9595), .B2(n15311), .A(n9594), .ZN(P2_U3222) );
  AOI211_X1 U12139 ( .C1(n9598), .C2(n9597), .A(n9596), .B(n15281), .ZN(n9599)
         );
  INV_X1 U12140 ( .A(n9599), .ZN(n9604) );
  OAI211_X1 U12141 ( .C1(n9602), .C2(n9601), .A(n15317), .B(n9600), .ZN(n9603)
         );
  NAND2_X1 U12142 ( .A1(n9604), .A2(n9603), .ZN(n9606) );
  NAND2_X1 U12143 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n10168) );
  INV_X1 U12144 ( .A(n10168), .ZN(n9605) );
  AOI211_X1 U12145 ( .C1(n15314), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n9606), .B(
        n9605), .ZN(n9607) );
  OAI21_X1 U12146 ( .B1(n9608), .B2(n15311), .A(n9607), .ZN(P2_U3218) );
  OAI211_X1 U12147 ( .C1(n9611), .C2(n9610), .A(n15317), .B(n9609), .ZN(n9617)
         );
  AOI211_X1 U12148 ( .C1(n9614), .C2(n9613), .A(n9612), .B(n15281), .ZN(n9615)
         );
  INV_X1 U12149 ( .A(n9615), .ZN(n9616) );
  NAND2_X1 U12150 ( .A1(n9617), .A2(n9616), .ZN(n9619) );
  NAND2_X1 U12151 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n12002) );
  INV_X1 U12152 ( .A(n12002), .ZN(n9618) );
  AOI211_X1 U12153 ( .C1(n15314), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n9619), .B(
        n9618), .ZN(n9620) );
  OAI21_X1 U12154 ( .B1(n9621), .B2(n15311), .A(n9620), .ZN(P2_U3219) );
  NOR2_X1 U12155 ( .A1(n9630), .A2(n9622), .ZN(n14551) );
  INV_X1 U12156 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10950) );
  MUX2_X1 U12157 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10950), .S(n14552), .Z(
        n9623) );
  OAI21_X1 U12158 ( .B1(n14557), .B2(n14551), .A(n9623), .ZN(n14555) );
  NAND2_X1 U12159 ( .A1(n14552), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9649) );
  INV_X1 U12160 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n13476) );
  MUX2_X1 U12161 ( .A(n13476), .B(P1_REG2_REG_8__SCAN_IN), .S(n10571), .Z(
        n9648) );
  AOI21_X1 U12162 ( .B1(n14555), .B2(n9649), .A(n9648), .ZN(n14579) );
  NOR2_X1 U12163 ( .A1(n9645), .A2(n13476), .ZN(n14573) );
  INV_X1 U12164 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10960) );
  MUX2_X1 U12165 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10960), .S(n14572), .Z(
        n9624) );
  OAI21_X1 U12166 ( .B1(n14579), .B2(n14573), .A(n9624), .ZN(n14577) );
  NAND2_X1 U12167 ( .A1(n14572), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9627) );
  INV_X1 U12168 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9625) );
  MUX2_X1 U12169 ( .A(n9625), .B(P1_REG2_REG_10__SCAN_IN), .S(n11108), .Z(
        n9626) );
  AOI21_X1 U12170 ( .B1(n14577), .B2(n9627), .A(n9626), .ZN(n9666) );
  NAND3_X1 U12171 ( .A1(n14577), .A2(n9627), .A3(n9626), .ZN(n9628) );
  NAND2_X1 U12172 ( .A1(n9628), .A2(n14576), .ZN(n9642) );
  INV_X1 U12173 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9631) );
  NOR2_X1 U12174 ( .A1(n9630), .A2(n9629), .ZN(n14547) );
  MUX2_X1 U12175 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9631), .S(n14552), .Z(
        n14546) );
  OAI21_X1 U12176 ( .B1(n14548), .B2(n14547), .A(n14546), .ZN(n14550) );
  OAI21_X1 U12177 ( .B1(n9631), .B2(n14543), .A(n14550), .ZN(n9643) );
  INV_X1 U12178 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9632) );
  NAND2_X1 U12179 ( .A1(n9645), .A2(n9632), .ZN(n9633) );
  OAI21_X1 U12180 ( .B1(n9645), .B2(n9632), .A(n9633), .ZN(n9644) );
  NOR2_X1 U12181 ( .A1(n9643), .A2(n9644), .ZN(n14564) );
  INV_X1 U12182 ( .A(n9633), .ZN(n14562) );
  INV_X1 U12183 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n13354) );
  MUX2_X1 U12184 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n13354), .S(n14572), .Z(
        n14563) );
  OAI21_X1 U12185 ( .B1(n14564), .B2(n14562), .A(n14563), .ZN(n14561) );
  OAI21_X1 U12186 ( .B1(n14572), .B2(P1_REG1_REG_9__SCAN_IN), .A(n14561), .ZN(
        n9635) );
  INV_X1 U12187 ( .A(n9635), .ZN(n9637) );
  INV_X1 U12188 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10738) );
  MUX2_X1 U12189 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10738), .S(n11108), .Z(
        n9636) );
  MUX2_X1 U12190 ( .A(n10738), .B(P1_REG1_REG_10__SCAN_IN), .S(n11108), .Z(
        n9634) );
  OR2_X1 U12191 ( .A1(n9635), .A2(n9634), .ZN(n9655) );
  OAI211_X1 U12192 ( .C1(n9637), .C2(n9636), .A(n14565), .B(n9655), .ZN(n9641)
         );
  INV_X1 U12193 ( .A(n15212), .ZN(n14571) );
  INV_X1 U12194 ( .A(n15199), .ZN(n15216) );
  NAND2_X1 U12195 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11200)
         );
  OAI21_X1 U12196 ( .B1(n15216), .B2(n9638), .A(n11200), .ZN(n9639) );
  AOI21_X1 U12197 ( .B1(n11108), .B2(n14571), .A(n9639), .ZN(n9640) );
  OAI211_X1 U12198 ( .C1(n9666), .C2(n9642), .A(n9641), .B(n9640), .ZN(
        P1_U3253) );
  AOI21_X1 U12199 ( .B1(n9644), .B2(n9643), .A(n14564), .ZN(n9654) );
  AND2_X1 U12200 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9647) );
  NOR2_X1 U12201 ( .A1(n15212), .A2(n9645), .ZN(n9646) );
  AOI211_X1 U12202 ( .C1(n15199), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9647), .B(
        n9646), .ZN(n9653) );
  INV_X1 U12203 ( .A(n14579), .ZN(n9651) );
  NAND3_X1 U12204 ( .A1(n14555), .A2(n9649), .A3(n9648), .ZN(n9650) );
  NAND3_X1 U12205 ( .A1(n14576), .A2(n9651), .A3(n9650), .ZN(n9652) );
  OAI211_X1 U12206 ( .C1(n9654), .C2(n15208), .A(n9653), .B(n9652), .ZN(
        P1_U3251) );
  INV_X1 U12207 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11123) );
  MUX2_X1 U12208 ( .A(n11123), .B(P1_REG1_REG_11__SCAN_IN), .S(n11139), .Z(
        n9657) );
  OAI21_X1 U12209 ( .B1(n10738), .B2(n9660), .A(n9655), .ZN(n9656) );
  NOR2_X1 U12210 ( .A1(n9656), .A2(n9657), .ZN(n9698) );
  AOI21_X1 U12211 ( .B1(n9657), .B2(n9656), .A(n9698), .ZN(n9669) );
  INV_X1 U12212 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9658) );
  NAND2_X1 U12213 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11480)
         );
  OAI21_X1 U12214 ( .B1(n15216), .B2(n9658), .A(n11480), .ZN(n9659) );
  AOI21_X1 U12215 ( .B1(n14571), .B2(n11139), .A(n9659), .ZN(n9668) );
  NOR2_X1 U12216 ( .A1(n9660), .A2(n9625), .ZN(n9664) );
  INV_X1 U12217 ( .A(n9664), .ZN(n9662) );
  INV_X1 U12218 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9691) );
  MUX2_X1 U12219 ( .A(n9691), .B(P1_REG2_REG_11__SCAN_IN), .S(n11139), .Z(
        n9661) );
  NAND2_X1 U12220 ( .A1(n9662), .A2(n9661), .ZN(n9665) );
  MUX2_X1 U12221 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n9691), .S(n11139), .Z(
        n9663) );
  OAI21_X1 U12222 ( .B1(n9666), .B2(n9664), .A(n9663), .ZN(n9690) );
  OAI211_X1 U12223 ( .C1(n9666), .C2(n9665), .A(n9690), .B(n14576), .ZN(n9667)
         );
  OAI211_X1 U12224 ( .C1(n9669), .C2(n15208), .A(n9668), .B(n9667), .ZN(
        P1_U3254) );
  INV_X1 U12225 ( .A(n11297), .ZN(n9672) );
  NAND2_X1 U12226 ( .A1(n9671), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9710) );
  XNOR2_X1 U12227 ( .A(n9710), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11298) );
  INV_X1 U12228 ( .A(n11298), .ZN(n9872) );
  OAI222_X1 U12229 ( .A1(n15024), .A2(n13505), .B1(n15030), .B2(n9672), .C1(
        P1_U3086), .C2(n9872), .ZN(P1_U3343) );
  INV_X1 U12230 ( .A(n10064), .ZN(n11000) );
  OAI222_X1 U12231 ( .A1(n14312), .A2(n9673), .B1(n11000), .B2(P2_U3088), .C1(
        n10596), .C2(n9672), .ZN(P2_U3315) );
  OAI21_X1 U12232 ( .B1(n9676), .B2(n9675), .A(n9674), .ZN(n9686) );
  INV_X1 U12233 ( .A(n9677), .ZN(n9681) );
  NOR3_X1 U12234 ( .A1(n14533), .A2(n9679), .A3(n9678), .ZN(n9680) );
  NOR3_X1 U12235 ( .A1(n15210), .A2(n9681), .A3(n9680), .ZN(n9685) );
  NAND2_X1 U12236 ( .A1(n14571), .A2(n10101), .ZN(n9682) );
  NAND2_X1 U12237 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10123) );
  OAI211_X1 U12238 ( .C1(n9683), .C2(n15216), .A(n9682), .B(n10123), .ZN(n9684) );
  AOI211_X1 U12239 ( .C1(n14565), .C2(n9686), .A(n9685), .B(n9684), .ZN(n9687)
         );
  INV_X1 U12240 ( .A(n9687), .ZN(P1_U3248) );
  INV_X1 U12241 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9688) );
  MUX2_X1 U12242 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9688), .S(n11298), .Z(
        n9689) );
  INV_X1 U12243 ( .A(n9689), .ZN(n9694) );
  OAI21_X1 U12244 ( .B1(n9692), .B2(n9691), .A(n9690), .ZN(n9693) );
  NOR2_X1 U12245 ( .A1(n9693), .A2(n9694), .ZN(n9871) );
  AOI21_X1 U12246 ( .B1(n9694), .B2(n9693), .A(n9871), .ZN(n9705) );
  NOR2_X1 U12247 ( .A1(n11139), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9696) );
  INV_X1 U12248 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9695) );
  MUX2_X1 U12249 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9695), .S(n11298), .Z(
        n9697) );
  OAI21_X1 U12250 ( .B1(n9698), .B2(n9696), .A(n9697), .ZN(n9870) );
  INV_X1 U12251 ( .A(n9870), .ZN(n9700) );
  NOR3_X1 U12252 ( .A1(n9698), .A2(n9697), .A3(n9696), .ZN(n9699) );
  OAI21_X1 U12253 ( .B1(n9700), .B2(n9699), .A(n14565), .ZN(n9704) );
  NOR2_X1 U12254 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11143), .ZN(n9702) );
  NOR2_X1 U12255 ( .A1(n15212), .A2(n9872), .ZN(n9701) );
  AOI211_X1 U12256 ( .C1(n15199), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n9702), .B(
        n9701), .ZN(n9703) );
  OAI211_X1 U12257 ( .C1(n9705), .C2(n15210), .A(n9704), .B(n9703), .ZN(
        P1_U3255) );
  INV_X1 U12258 ( .A(n9706), .ZN(n9708) );
  OAI222_X1 U12259 ( .A1(n13756), .A2(n9708), .B1(n12609), .B2(n9707), .C1(
        n12955), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12260 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9709) );
  NAND2_X1 U12261 ( .A1(n9710), .A2(n9709), .ZN(n9711) );
  NAND2_X1 U12262 ( .A1(n9711), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9891) );
  XNOR2_X1 U12263 ( .A(n9891), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11424) );
  INV_X1 U12264 ( .A(n11424), .ZN(n10079) );
  INV_X1 U12265 ( .A(n11423), .ZN(n9712) );
  OAI222_X1 U12266 ( .A1(n10079), .A2(P1_U3086), .B1(n15024), .B2(n7971), .C1(
        n9712), .C2(n15030), .ZN(P1_U3342) );
  OAI222_X1 U12267 ( .A1(n14312), .A2(n9713), .B1(n11002), .B2(P2_U3088), .C1(
        n10596), .C2(n9712), .ZN(P2_U3314) );
  INV_X1 U12268 ( .A(n9714), .ZN(n9720) );
  NAND2_X1 U12269 ( .A1(n9720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9716) );
  INV_X1 U12270 ( .A(n9717), .ZN(n9718) );
  NAND2_X1 U12271 ( .A1(n9718), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9719) );
  MUX2_X1 U12272 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9719), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9721) );
  NAND2_X1 U12273 ( .A1(n11165), .A2(n11695), .ZN(n9722) );
  AND2_X1 U12274 ( .A1(n12293), .A2(n9722), .ZN(n9819) );
  INV_X1 U12275 ( .A(n12528), .ZN(n9737) );
  NOR4_X1 U12276 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9731) );
  NOR4_X1 U12277 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9730) );
  INV_X1 U12278 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15220) );
  INV_X1 U12279 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15221) );
  INV_X1 U12280 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n15218) );
  INV_X1 U12281 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n15222) );
  NAND4_X1 U12282 ( .A1(n15220), .A2(n15221), .A3(n15218), .A4(n15222), .ZN(
        n9728) );
  NOR4_X1 U12283 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n9726) );
  NOR4_X1 U12284 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n9725) );
  NOR4_X1 U12285 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9724) );
  NOR4_X1 U12286 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n9723) );
  NAND4_X1 U12287 ( .A1(n9726), .A2(n9725), .A3(n9724), .A4(n9723), .ZN(n9727)
         );
  NOR4_X1 U12288 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9728), .A4(n9727), .ZN(n9729) );
  AND3_X1 U12289 ( .A1(n9731), .A2(n9730), .A3(n9729), .ZN(n9732) );
  NOR2_X1 U12290 ( .A1(n9738), .A2(n9732), .ZN(n9787) );
  INV_X1 U12291 ( .A(n9787), .ZN(n9736) );
  AND2_X2 U12292 ( .A1(n15233), .A2(n11165), .ZN(n14888) );
  OR2_X1 U12293 ( .A1(n9738), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9735) );
  INV_X1 U12294 ( .A(n9733), .ZN(n15032) );
  NAND2_X1 U12295 ( .A1(n15032), .A2(n11725), .ZN(n9734) );
  NAND2_X1 U12296 ( .A1(n9735), .A2(n9734), .ZN(n9786) );
  NAND4_X1 U12297 ( .A1(n9737), .A2(n9736), .A3(n9829), .A4(n9786), .ZN(n9967)
         );
  OR2_X1 U12298 ( .A1(n9738), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9740) );
  NAND2_X1 U12299 ( .A1(n15032), .A2(n9397), .ZN(n9739) );
  NOR2_X2 U12300 ( .A1(n9967), .A2(n9788), .ZN(n15267) );
  NAND2_X1 U12301 ( .A1(n9743), .A2(n9742), .ZN(n9746) );
  XNOR2_X2 U12302 ( .A(n9745), .B(n9744), .ZN(n15023) );
  INV_X1 U12303 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9843) );
  AND2_X4 U12304 ( .A1(n15020), .A2(n15023), .ZN(n12450) );
  OR2_X1 U12305 ( .A1(n12289), .A2(n9567), .ZN(n9749) );
  INV_X1 U12306 ( .A(n12308), .ZN(n14844) );
  INV_X1 U12307 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n14853) );
  OR2_X1 U12308 ( .A1(n11986), .A2(n14853), .ZN(n9759) );
  NAND2_X1 U12309 ( .A1(n12450), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9758) );
  INV_X1 U12310 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9754) );
  OR2_X1 U12311 ( .A1(n11649), .A2(n9754), .ZN(n9757) );
  INV_X1 U12312 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9755) );
  OR2_X1 U12313 ( .A1(n12289), .A2(n9755), .ZN(n9756) );
  AND4_X2 U12314 ( .A1(n9759), .A2(n9758), .A3(n9757), .A4(n9756), .ZN(n12489)
         );
  NOR2_X1 U12315 ( .A1(n12490), .A2(n12489), .ZN(n9767) );
  INV_X1 U12316 ( .A(n9767), .ZN(n9764) );
  NOR2_X1 U12317 ( .A1(n7274), .A2(n9760), .ZN(n9762) );
  XNOR2_X1 U12318 ( .A(n9762), .B(n9761), .ZN(n15035) );
  MUX2_X1 U12319 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15035), .S(n9751), .Z(n15232)
         );
  OR2_X1 U12320 ( .A1(n12489), .A2(n12303), .ZN(n9763) );
  NAND2_X1 U12321 ( .A1(n12490), .A2(n9763), .ZN(n10311) );
  OAI21_X1 U12322 ( .B1(n9764), .B2(n12303), .A(n10311), .ZN(n14845) );
  INV_X1 U12323 ( .A(n14845), .ZN(n9784) );
  NAND2_X1 U12324 ( .A1(n11165), .A2(n14768), .ZN(n9765) );
  OR2_X1 U12325 ( .A1(n15034), .A2(n9765), .ZN(n14946) );
  NAND2_X1 U12326 ( .A1(n15034), .A2(n14768), .ZN(n9766) );
  INV_X1 U12327 ( .A(n11165), .ZN(n12296) );
  NAND2_X1 U12328 ( .A1(n9775), .A2(n12296), .ZN(n12455) );
  INV_X1 U12329 ( .A(n12293), .ZN(n9774) );
  OAI21_X1 U12330 ( .B1(n9767), .B2(n15228), .A(n14824), .ZN(n9779) );
  NAND2_X1 U12331 ( .A1(n12308), .A2(n12303), .ZN(n10338) );
  OAI21_X1 U12332 ( .B1(n12308), .B2(n12303), .A(n10338), .ZN(n9780) );
  XNOR2_X1 U12333 ( .A(n9780), .B(n12307), .ZN(n9768) );
  OAI21_X1 U12334 ( .B1(n9768), .B2(n15228), .A(n12489), .ZN(n9778) );
  NAND2_X1 U12335 ( .A1(n12450), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9773) );
  INV_X1 U12336 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10858) );
  OR2_X1 U12337 ( .A1(n11986), .A2(n10858), .ZN(n9772) );
  OR2_X1 U12338 ( .A1(n11649), .A2(n9769), .ZN(n9771) );
  OR2_X1 U12339 ( .A1(n12289), .A2(n10857), .ZN(n9770) );
  INV_X1 U12340 ( .A(n12315), .ZN(n14475) );
  NAND2_X1 U12341 ( .A1(n15034), .A2(n11695), .ZN(n9776) );
  NAND2_X1 U12342 ( .A1(n9775), .A2(n11165), .ZN(n12300) );
  AND2_X2 U12343 ( .A1(n9776), .A2(n12300), .ZN(n11728) );
  NOR2_X1 U12344 ( .A1(n9776), .A2(n12300), .ZN(n9777) );
  NOR2_X1 U12345 ( .A1(n11728), .A2(n9777), .ZN(n10830) );
  NAND2_X1 U12346 ( .A1(n10830), .A2(n11695), .ZN(n14789) );
  INV_X1 U12347 ( .A(n14789), .ZN(n14629) );
  AOI222_X1 U12348 ( .A1(n9779), .A2(n9778), .B1(n14475), .B2(n14850), .C1(
        n14845), .C2(n14629), .ZN(n14841) );
  INV_X1 U12349 ( .A(n9780), .ZN(n14843) );
  INV_X1 U12350 ( .A(n15233), .ZN(n9781) );
  OR2_X1 U12351 ( .A1(n9781), .A2(n11695), .ZN(n9782) );
  NAND2_X1 U12352 ( .A1(n12298), .A2(n12296), .ZN(n12522) );
  AOI22_X1 U12353 ( .A1(n14843), .A2(n14888), .B1(n14844), .B2(n14966), .ZN(
        n9783) );
  OAI211_X1 U12354 ( .C1(n9784), .C2(n14946), .A(n14841), .B(n9783), .ZN(n9968) );
  NAND2_X1 U12355 ( .A1(n9968), .A2(n15267), .ZN(n9785) );
  OAI21_X1 U12356 ( .B1(n15267), .B2(n14479), .A(n9785), .ZN(P1_U3529) );
  NOR2_X1 U12357 ( .A1(n9787), .A2(n9786), .ZN(n10818) );
  INV_X1 U12358 ( .A(n9788), .ZN(n10817) );
  NAND2_X1 U12359 ( .A1(n10818), .A2(n10817), .ZN(n9823) );
  OR2_X1 U12360 ( .A1(n9823), .A2(n9830), .ZN(n9831) );
  INV_X1 U12361 ( .A(n9831), .ZN(n9790) );
  NOR2_X1 U12362 ( .A1(n14966), .A2(n12293), .ZN(n9789) );
  OR2_X1 U12363 ( .A1(n9791), .A2(n11448), .ZN(n9795) );
  INV_X1 U12364 ( .A(n9793), .ZN(n9794) );
  INV_X1 U12365 ( .A(n12300), .ZN(n9796) );
  OAI22_X1 U12366 ( .A1(n12314), .A2(n12666), .B1(n12665), .B2(n12315), .ZN(
        n9798) );
  XNOR2_X1 U12367 ( .A(n9798), .B(n11728), .ZN(n10002) );
  NAND2_X1 U12368 ( .A1(n14888), .A2(n11695), .ZN(n14659) );
  AND2_X4 U12369 ( .A1(n9802), .A2(n14659), .ZN(n12709) );
  INV_X1 U12370 ( .A(n12709), .ZN(n9800) );
  XNOR2_X1 U12371 ( .A(n10002), .B(n10000), .ZN(n9818) );
  INV_X1 U12372 ( .A(n9797), .ZN(n9803) );
  AOI22_X1 U12373 ( .A1(n10503), .A2(n15232), .B1(n9803), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9801) );
  OAI21_X1 U12374 ( .B1(n9800), .B2(n12489), .A(n9801), .ZN(n9848) );
  INV_X1 U12375 ( .A(n12489), .ZN(n14476) );
  NAND2_X1 U12376 ( .A1(n10503), .A2(n14476), .ZN(n9806) );
  NAND2_X1 U12377 ( .A1(n9802), .A2(n15232), .ZN(n9805) );
  NAND2_X1 U12378 ( .A1(n9803), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9804) );
  INV_X1 U12379 ( .A(n9847), .ZN(n9807) );
  OR2_X1 U12380 ( .A1(n9807), .A2(n11728), .ZN(n9808) );
  NAND2_X1 U12381 ( .A1(n9850), .A2(n9808), .ZN(n9839) );
  OAI22_X1 U12382 ( .A1(n12308), .A2(n12666), .B1(n12665), .B2(n12307), .ZN(
        n9809) );
  XNOR2_X1 U12383 ( .A(n9809), .B(n11728), .ZN(n9811) );
  INV_X1 U12384 ( .A(n12307), .ZN(n14851) );
  NOR2_X1 U12385 ( .A1(n12665), .A2(n12308), .ZN(n9810) );
  NAND2_X1 U12386 ( .A1(n9811), .A2(n9812), .ZN(n9816) );
  INV_X1 U12387 ( .A(n9811), .ZN(n9814) );
  INV_X1 U12388 ( .A(n9812), .ZN(n9813) );
  NAND2_X1 U12389 ( .A1(n9814), .A2(n9813), .ZN(n9815) );
  OAI21_X1 U12390 ( .B1(n9818), .B2(n9817), .A(n10004), .ZN(n9836) );
  OAI21_X1 U12391 ( .B1(n9823), .B2(n9819), .A(n9829), .ZN(n9822) );
  AND2_X1 U12392 ( .A1(n9797), .A2(n9820), .ZN(n9821) );
  NAND2_X1 U12393 ( .A1(n9822), .A2(n9821), .ZN(n10028) );
  NOR2_X1 U12394 ( .A1(n10028), .A2(P1_U3086), .ZN(n9853) );
  NOR2_X2 U12395 ( .A1(n14410), .A2(n14824), .ZN(n14447) );
  NOR2_X2 U12396 ( .A1(n14410), .A2(n14826), .ZN(n14438) );
  NAND2_X1 U12397 ( .A1(n12450), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9828) );
  OR2_X1 U12398 ( .A1(n11649), .A2(n9824), .ZN(n9827) );
  OR2_X1 U12399 ( .A1(n12289), .A2(n10848), .ZN(n9826) );
  OR2_X1 U12400 ( .A1(n11986), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9825) );
  AND4_X2 U12401 ( .A1(n9828), .A2(n9827), .A3(n9826), .A4(n9825), .ZN(n10331)
         );
  AOI22_X1 U12402 ( .A1(n14447), .A2(n14851), .B1(n14438), .B2(n14474), .ZN(
        n9834) );
  NAND2_X1 U12403 ( .A1(n9832), .A2(n12312), .ZN(n9833) );
  OAI211_X1 U12404 ( .C1(n9853), .C2(n10858), .A(n9834), .B(n9833), .ZN(n9835)
         );
  AOI21_X1 U12405 ( .B1(n14425), .B2(n9836), .A(n9835), .ZN(n9837) );
  INV_X1 U12406 ( .A(n9837), .ZN(P1_U3237) );
  OAI21_X1 U12407 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(n9845) );
  AOI22_X1 U12408 ( .A1(n14447), .A2(n14476), .B1(n14438), .B2(n14475), .ZN(
        n9842) );
  NAND2_X1 U12409 ( .A1(n9832), .A2(n14844), .ZN(n9841) );
  OAI211_X1 U12410 ( .C1(n9853), .C2(n9843), .A(n9842), .B(n9841), .ZN(n9844)
         );
  AOI21_X1 U12411 ( .B1(n14425), .B2(n9845), .A(n9844), .ZN(n9846) );
  INV_X1 U12412 ( .A(n9846), .ZN(P1_U3222) );
  NAND2_X1 U12413 ( .A1(n9848), .A2(n9847), .ZN(n9849) );
  AND2_X1 U12414 ( .A1(n9850), .A2(n9849), .ZN(n14493) );
  OAI22_X1 U12415 ( .A1(n14449), .A2(n12307), .B1(n14493), .B2(n14456), .ZN(
        n9851) );
  AOI21_X1 U12416 ( .B1(n15232), .B2(n9832), .A(n9851), .ZN(n9852) );
  OAI21_X1 U12417 ( .B1(n9853), .B2(n14853), .A(n9852), .ZN(P1_U3232) );
  INV_X1 U12418 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n13916) );
  MUX2_X1 U12419 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n13916), .S(n13925), .Z(
        n9855) );
  NAND2_X1 U12420 ( .A1(n13922), .A2(n9855), .ZN(n13920) );
  OR2_X1 U12421 ( .A1(n13925), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n13921) );
  NAND2_X1 U12422 ( .A1(n13920), .A2(n13921), .ZN(n9858) );
  INV_X1 U12423 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9856) );
  MUX2_X1 U12424 ( .A(n9856), .B(P2_REG2_REG_10__SCAN_IN), .S(n10060), .Z(
        n9857) );
  NOR2_X1 U12425 ( .A1(n9858), .A2(n9857), .ZN(n10059) );
  AOI211_X1 U12426 ( .C1(n9858), .C2(n9857), .A(n15281), .B(n10059), .ZN(n9859) );
  INV_X1 U12427 ( .A(n9859), .ZN(n9869) );
  NAND2_X1 U12428 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10900)
         );
  INV_X1 U12429 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n15400) );
  MUX2_X1 U12430 ( .A(n15400), .B(P2_REG1_REG_10__SCAN_IN), .S(n10060), .Z(
        n9864) );
  AOI21_X1 U12431 ( .B1(n9861), .B2(P2_REG1_REG_8__SCAN_IN), .A(n9860), .ZN(
        n13926) );
  INV_X1 U12432 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n13917) );
  MUX2_X1 U12433 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n13917), .S(n13925), .Z(
        n9862) );
  NAND2_X1 U12434 ( .A1(n13926), .A2(n9862), .ZN(n13927) );
  OAI21_X1 U12435 ( .B1(n13925), .B2(P2_REG1_REG_9__SCAN_IN), .A(n13927), .ZN(
        n9863) );
  NOR2_X1 U12436 ( .A1(n9863), .A2(n9864), .ZN(n13947) );
  AOI211_X1 U12437 ( .C1(n9864), .C2(n9863), .A(n13947), .B(n15269), .ZN(n9865) );
  INV_X1 U12438 ( .A(n9865), .ZN(n9866) );
  NAND2_X1 U12439 ( .A1(n10900), .A2(n9866), .ZN(n9867) );
  AOI21_X1 U12440 ( .B1(n15314), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9867), .ZN(
        n9868) );
  OAI211_X1 U12441 ( .C1(n15311), .C2(n10054), .A(n9869), .B(n9868), .ZN(
        P2_U3224) );
  OAI21_X1 U12442 ( .B1(n11298), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9870), .ZN(
        n10077) );
  INV_X1 U12443 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11501) );
  MUX2_X1 U12444 ( .A(n11501), .B(P1_REG1_REG_13__SCAN_IN), .S(n11424), .Z(
        n10076) );
  XNOR2_X1 U12445 ( .A(n10077), .B(n10076), .ZN(n9881) );
  NAND2_X1 U12446 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11614)
         );
  AOI21_X1 U12447 ( .B1(n9872), .B2(n9688), .A(n9871), .ZN(n9876) );
  INV_X1 U12448 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9873) );
  MUX2_X1 U12449 ( .A(n9873), .B(P1_REG2_REG_13__SCAN_IN), .S(n11424), .Z(
        n9874) );
  INV_X1 U12450 ( .A(n9874), .ZN(n9875) );
  NAND2_X1 U12451 ( .A1(n9876), .A2(n9875), .ZN(n10084) );
  OAI211_X1 U12452 ( .C1(n9876), .C2(n9875), .A(n14576), .B(n10084), .ZN(n9877) );
  NAND2_X1 U12453 ( .A1(n11614), .A2(n9877), .ZN(n9879) );
  NOR2_X1 U12454 ( .A1(n15212), .A2(n10079), .ZN(n9878) );
  AOI211_X1 U12455 ( .C1(n15199), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n9879), .B(
        n9878), .ZN(n9880) );
  OAI21_X1 U12456 ( .B1(n9881), .B2(n15208), .A(n9880), .ZN(P1_U3256) );
  INV_X1 U12457 ( .A(n9882), .ZN(n9885) );
  INV_X1 U12458 ( .A(n12992), .ZN(n12959) );
  AOI222_X1 U12459 ( .A1(n9885), .A2(n13749), .B1(n12959), .B2(
        P3_STATE_REG_SCAN_IN), .C1(n9884), .C2(n9883), .ZN(P3_U3280) );
  INV_X1 U12460 ( .A(n13011), .ZN(n13019) );
  OAI222_X1 U12461 ( .A1(n13756), .A2(n9887), .B1(n13019), .B2(P3_U3151), .C1(
        n9886), .C2(n12609), .ZN(P3_U3279) );
  INV_X1 U12462 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n9889) );
  NAND2_X1 U12463 ( .A1(n12833), .A2(P3_U3897), .ZN(n9888) );
  OAI21_X1 U12464 ( .B1(P3_U3897), .B2(n9889), .A(n9888), .ZN(P3_U3505) );
  INV_X1 U12465 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9890) );
  NAND2_X1 U12466 ( .A1(n9891), .A2(n9890), .ZN(n9892) );
  NAND2_X1 U12467 ( .A1(n9892), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9893) );
  XNOR2_X1 U12468 ( .A(n9893), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11450) );
  INV_X1 U12469 ( .A(n11450), .ZN(n10939) );
  OAI222_X1 U12470 ( .A1(P1_U3086), .A2(n10939), .B1(n15030), .B2(n11449), 
        .C1(n9894), .C2(n15024), .ZN(P1_U3341) );
  INV_X1 U12471 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n9896) );
  NAND2_X1 U12472 ( .A1(n13582), .A2(P3_U3897), .ZN(n9895) );
  OAI21_X1 U12473 ( .B1(P3_U3897), .B2(n9896), .A(n9895), .ZN(P3_U3506) );
  INV_X1 U12474 ( .A(n11268), .ZN(n11278) );
  OAI222_X1 U12475 ( .A1(n14312), .A2(n9897), .B1(n11278), .B2(P2_U3088), .C1(
        n10596), .C2(n11449), .ZN(P2_U3313) );
  NAND2_X1 U12476 ( .A1(n9901), .A2(n9914), .ZN(n9907) );
  XNOR2_X1 U12477 ( .A(n9906), .B(n9907), .ZN(n10130) );
  OR2_X1 U12478 ( .A1(n10158), .A2(n10143), .ZN(n10129) );
  OAI21_X1 U12479 ( .B1(n9902), .B2(n10037), .A(n10129), .ZN(n9903) );
  NAND2_X1 U12480 ( .A1(n9906), .A2(n9907), .ZN(n9908) );
  NAND2_X1 U12481 ( .A1(n10131), .A2(n9908), .ZN(n9909) );
  XNOR2_X1 U12482 ( .A(n10158), .B(n14158), .ZN(n9910) );
  NAND2_X1 U12483 ( .A1(n13915), .A2(n9914), .ZN(n9911) );
  XNOR2_X1 U12484 ( .A(n9910), .B(n9911), .ZN(n11802) );
  INV_X1 U12485 ( .A(n9910), .ZN(n9912) );
  NAND2_X1 U12486 ( .A1(n9912), .A2(n9911), .ZN(n9913) );
  XNOR2_X1 U12487 ( .A(n9941), .B(n10158), .ZN(n10163) );
  AND2_X1 U12488 ( .A1(n13914), .A2(n9914), .ZN(n9915) );
  NAND2_X1 U12489 ( .A1(n10163), .A2(n9915), .ZN(n10159) );
  OR2_X1 U12490 ( .A1(n10163), .A2(n9915), .ZN(n9916) );
  NAND2_X1 U12491 ( .A1(n10159), .A2(n9916), .ZN(n9926) );
  INV_X1 U12492 ( .A(n15348), .ZN(n9917) );
  NAND2_X1 U12493 ( .A1(n9918), .A2(n9917), .ZN(n9930) );
  NAND2_X1 U12494 ( .A1(n15352), .A2(n9919), .ZN(n9920) );
  INV_X1 U12495 ( .A(n9921), .ZN(n9922) );
  AND2_X1 U12496 ( .A1(n15386), .A2(n9922), .ZN(n9923) );
  INV_X1 U12497 ( .A(n9926), .ZN(n9924) );
  INV_X1 U12498 ( .A(n10161), .ZN(n9925) );
  AOI211_X1 U12499 ( .C1(n9927), .C2(n9926), .A(n13872), .B(n9925), .ZN(n9945)
         );
  INV_X1 U12500 ( .A(n9928), .ZN(n9929) );
  INV_X1 U12501 ( .A(n13853), .ZN(n15106) );
  NAND2_X1 U12502 ( .A1(n15106), .A2(n14027), .ZN(n13883) );
  OR2_X1 U12503 ( .A1(n13853), .A2(n15096), .ZN(n13881) );
  INV_X1 U12504 ( .A(n13881), .ZN(n12009) );
  NAND2_X1 U12505 ( .A1(n9930), .A2(n9931), .ZN(n9936) );
  NAND2_X1 U12506 ( .A1(n9931), .A2(n15351), .ZN(n9962) );
  AND4_X1 U12507 ( .A1(n9934), .A2(n9933), .A3(n9932), .A4(n9962), .ZN(n9935)
         );
  NAND2_X1 U12508 ( .A1(n9936), .A2(n9935), .ZN(n9993) );
  AOI22_X1 U12509 ( .A1(n12009), .A2(n13915), .B1(n13855), .B2(n9937), .ZN(
        n9943) );
  NAND2_X1 U12510 ( .A1(n9939), .A2(n9938), .ZN(n9940) );
  NOR2_X1 U12511 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9937), .ZN(n15274) );
  AOI21_X1 U12512 ( .B1(n15107), .B2(n9941), .A(n15274), .ZN(n9942) );
  OAI211_X1 U12513 ( .C1(n12011), .C2(n13883), .A(n9943), .B(n9942), .ZN(n9944) );
  OR2_X1 U12514 ( .A1(n9945), .A2(n9944), .ZN(P2_U3190) );
  NAND2_X1 U12515 ( .A1(n10146), .A2(n9019), .ZN(n10605) );
  INV_X1 U12516 ( .A(n9946), .ZN(n9947) );
  AOI21_X1 U12517 ( .B1(n10138), .B2(n9949), .A(n9947), .ZN(n9952) );
  INV_X1 U12518 ( .A(n9952), .ZN(n14167) );
  INV_X1 U12519 ( .A(n10038), .ZN(n9948) );
  AOI211_X1 U12520 ( .C1(n10143), .C2(n14166), .A(n13997), .B(n9948), .ZN(
        n14169) );
  OAI21_X1 U12521 ( .B1(n9950), .B2(n9949), .A(n10041), .ZN(n9955) );
  INV_X1 U12522 ( .A(n14027), .ZN(n15098) );
  INV_X1 U12523 ( .A(n9026), .ZN(n9951) );
  OAI22_X1 U12524 ( .A1(n10135), .A2(n15098), .B1(n9951), .B2(n15096), .ZN(
        n9954) );
  NOR2_X1 U12525 ( .A1(n9952), .A2(n9899), .ZN(n9953) );
  AOI211_X1 U12526 ( .C1(n6580), .C2(n9955), .A(n9954), .B(n9953), .ZN(n14164)
         );
  INV_X1 U12527 ( .A(n14164), .ZN(n9956) );
  AOI211_X1 U12528 ( .C1(n15390), .C2(n14167), .A(n14169), .B(n9956), .ZN(
        n9966) );
  INV_X1 U12529 ( .A(n9962), .ZN(n9957) );
  AND2_X1 U12530 ( .A1(n15348), .A2(n9957), .ZN(n9958) );
  NAND2_X1 U12531 ( .A1(n15393), .A2(n14258), .ZN(n14287) );
  INV_X1 U12532 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9959) );
  OAI22_X1 U12533 ( .A1(n14287), .A2(n9900), .B1(n15393), .B2(n9959), .ZN(
        n9960) );
  INV_X1 U12534 ( .A(n9960), .ZN(n9961) );
  OAI21_X1 U12535 ( .B1(n9966), .B2(n15391), .A(n9961), .ZN(P2_U3433) );
  NOR2_X1 U12536 ( .A1(n15348), .A2(n9962), .ZN(n9963) );
  NAND2_X1 U12537 ( .A1(n15404), .A2(n14258), .ZN(n14230) );
  AOI22_X1 U12538 ( .A1(n14248), .A2(n14166), .B1(n6794), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n9965) );
  OAI21_X1 U12539 ( .B1(n9966), .B2(n6794), .A(n9965), .ZN(P2_U3500) );
  INV_X1 U12540 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9970) );
  NAND2_X1 U12541 ( .A1(n9968), .A2(n15259), .ZN(n9969) );
  OAI21_X1 U12542 ( .B1(n15259), .B2(n9970), .A(n9969), .ZN(P1_U3462) );
  NAND2_X1 U12543 ( .A1(n15516), .A2(n10524), .ZN(n12059) );
  INV_X1 U12544 ( .A(n12059), .ZN(n12063) );
  NOR2_X1 U12545 ( .A1(n15520), .A2(n12063), .ZN(n12200) );
  INV_X1 U12546 ( .A(n9979), .ZN(n9972) );
  NAND2_X1 U12547 ( .A1(n9980), .A2(n15559), .ZN(n9971) );
  OAI22_X1 U12548 ( .A1(n9972), .A2(n9987), .B1(n9981), .B2(n9971), .ZN(n9974)
         );
  OR2_X1 U12549 ( .A1(n10182), .A2(n12230), .ZN(n9976) );
  NOR2_X1 U12550 ( .A1(n9987), .A2(n9976), .ZN(n10363) );
  NAND2_X1 U12551 ( .A1(n9981), .A2(n15504), .ZN(n9977) );
  AOI22_X1 U12552 ( .A1(n9975), .A2(n12878), .B1(n12869), .B2(n9978), .ZN(
        n9992) );
  NAND2_X1 U12553 ( .A1(n9987), .A2(n9979), .ZN(n9985) );
  NAND2_X1 U12554 ( .A1(n9981), .A2(n9980), .ZN(n9983) );
  NAND4_X1 U12555 ( .A1(n9985), .A2(n9984), .A3(n9983), .A4(n9982), .ZN(n9986)
         );
  NAND2_X1 U12556 ( .A1(n9986), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9989) );
  NOR2_X1 U12557 ( .A1(n10182), .A2(n10152), .ZN(n12233) );
  NAND2_X1 U12558 ( .A1(n9987), .A2(n12233), .ZN(n9988) );
  AND2_X1 U12559 ( .A1(n9989), .A2(n9988), .ZN(n10620) );
  NAND2_X1 U12560 ( .A1(n10620), .A2(n9990), .ZN(n10532) );
  NAND2_X1 U12561 ( .A1(n10532), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9991) );
  OAI211_X1 U12562 ( .C1(n12200), .C2(n12872), .A(n9992), .B(n9991), .ZN(
        P3_U3172) );
  NOR2_X1 U12563 ( .A1(n9993), .A2(P2_U3088), .ZN(n11806) );
  INV_X1 U12564 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9999) );
  NAND2_X1 U12565 ( .A1(n13875), .A2(n9026), .ZN(n9996) );
  AOI21_X1 U12566 ( .B1(n9026), .B2(n13997), .A(n13872), .ZN(n9994) );
  NOR2_X1 U12567 ( .A1(n9994), .A2(n15107), .ZN(n9995) );
  MUX2_X1 U12568 ( .A(n9996), .B(n9995), .S(n10143), .Z(n9998) );
  INV_X1 U12569 ( .A(n13883), .ZN(n10167) );
  NAND2_X1 U12570 ( .A1(n10167), .A2(n9901), .ZN(n9997) );
  OAI211_X1 U12571 ( .C1(n11806), .C2(n9999), .A(n9998), .B(n9997), .ZN(
        P2_U3204) );
  INV_X1 U12572 ( .A(n10000), .ZN(n10001) );
  NAND2_X1 U12573 ( .A1(n10002), .A2(n10001), .ZN(n10003) );
  NAND2_X1 U12574 ( .A1(n10005), .A2(n12456), .ZN(n10007) );
  INV_X2 U12575 ( .A(n12458), .ZN(n11845) );
  AOI22_X1 U12576 ( .A1(n11845), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n11844), 
        .B2(n14515), .ZN(n10006) );
  OAI22_X1 U12577 ( .A1(n15236), .A2(n12666), .B1(n12665), .B2(n10331), .ZN(
        n10008) );
  XNOR2_X1 U12578 ( .A(n10008), .B(n12710), .ZN(n10010) );
  OAI22_X1 U12579 ( .A1(n12664), .A2(n10331), .B1(n15236), .B2(n12665), .ZN(
        n10009) );
  NAND2_X1 U12580 ( .A1(n10010), .A2(n10009), .ZN(n10093) );
  NAND2_X1 U12581 ( .A1(n10094), .A2(n10093), .ZN(n10021) );
  NAND2_X1 U12582 ( .A1(n10011), .A2(n12456), .ZN(n10014) );
  AOI22_X1 U12583 ( .A1(n11845), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11844), 
        .B2(n10012), .ZN(n10013) );
  NAND2_X1 U12584 ( .A1(n12450), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10018) );
  OR2_X1 U12585 ( .A1(n11649), .A2(n13501), .ZN(n10017) );
  XNOR2_X1 U12586 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10833) );
  OR2_X1 U12587 ( .A1(n11986), .A2(n10833), .ZN(n10016) );
  OR2_X1 U12588 ( .A1(n12289), .A2(n9570), .ZN(n10015) );
  OAI22_X1 U12589 ( .A1(n12325), .A2(n12666), .B1(n12665), .B2(n12326), .ZN(
        n10019) );
  XNOR2_X1 U12590 ( .A(n10019), .B(n12710), .ZN(n10095) );
  OAI22_X1 U12591 ( .A1(n12664), .A2(n12326), .B1(n12325), .B2(n12665), .ZN(
        n10091) );
  INV_X1 U12592 ( .A(n10091), .ZN(n10096) );
  XNOR2_X1 U12593 ( .A(n10095), .B(n10096), .ZN(n10020) );
  XNOR2_X1 U12594 ( .A(n10021), .B(n10020), .ZN(n10032) );
  INV_X1 U12595 ( .A(n12325), .ZN(n12324) );
  AOI22_X1 U12596 ( .A1(n12324), .A2(n9832), .B1(n14447), .B2(n14474), .ZN(
        n10031) );
  AOI21_X1 U12597 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10022) );
  NOR2_X1 U12598 ( .A1(n10022), .A2(n10114), .ZN(n11071) );
  NAND2_X1 U12599 ( .A1(n11878), .A2(n11071), .ZN(n10027) );
  OR2_X1 U12600 ( .A1(n12289), .A2(n11068), .ZN(n10026) );
  INV_X1 U12601 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10023) );
  OR2_X1 U12602 ( .A1(n11944), .A2(n10023), .ZN(n10025) );
  OR2_X1 U12603 ( .A1(n12454), .A2(n15262), .ZN(n10024) );
  NAND4_X1 U12604 ( .A1(n10027), .A2(n10026), .A3(n10025), .A4(n10024), .ZN(
        n14472) );
  INV_X1 U12605 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n13455) );
  NOR2_X1 U12606 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13455), .ZN(n14523) );
  NOR2_X1 U12607 ( .A1(n14441), .A2(n10833), .ZN(n10029) );
  AOI211_X1 U12608 ( .C1(n14438), .C2(n14472), .A(n14523), .B(n10029), .ZN(
        n10030) );
  OAI211_X1 U12609 ( .C1(n10032), .C2(n14456), .A(n10031), .B(n10030), .ZN(
        P1_U3230) );
  INV_X1 U12610 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n10034) );
  INV_X1 U12611 ( .A(n15435), .ZN(n15064) );
  NAND2_X1 U12612 ( .A1(n15064), .A2(P3_U3897), .ZN(n10033) );
  OAI21_X1 U12613 ( .B1(P3_U3897), .B2(n10034), .A(n10033), .ZN(P3_U3502) );
  OAI21_X1 U12614 ( .B1(n10036), .B2(n10040), .A(n10035), .ZN(n14156) );
  AOI211_X1 U12615 ( .C1(n14158), .C2(n10038), .A(n13997), .B(n10672), .ZN(
        n14157) );
  INV_X1 U12616 ( .A(n9899), .ZN(n10551) );
  AOI22_X1 U12617 ( .A1(n14025), .A2(n9901), .B1(n13914), .B2(n14027), .ZN(
        n11805) );
  INV_X1 U12618 ( .A(n11805), .ZN(n10045) );
  NAND3_X1 U12619 ( .A1(n10041), .A2(n10040), .A3(n10039), .ZN(n10042) );
  AOI21_X1 U12620 ( .B1(n10043), .B2(n10042), .A(n15125), .ZN(n10044) );
  AOI211_X1 U12621 ( .C1(n10551), .C2(n14156), .A(n10045), .B(n10044), .ZN(
        n14159) );
  INV_X1 U12622 ( .A(n14159), .ZN(n10046) );
  AOI211_X1 U12623 ( .C1(n15390), .C2(n14156), .A(n14157), .B(n10046), .ZN(
        n10052) );
  INV_X1 U12624 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10047) );
  OAI22_X1 U12625 ( .A1(n14287), .A2(n10048), .B1(n15393), .B2(n10047), .ZN(
        n10049) );
  INV_X1 U12626 ( .A(n10049), .ZN(n10050) );
  OAI21_X1 U12627 ( .B1(n10052), .B2(n15391), .A(n10050), .ZN(P2_U3436) );
  AOI22_X1 U12628 ( .A1(n14248), .A2(n14158), .B1(n6794), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10051) );
  OAI21_X1 U12629 ( .B1(n10052), .B2(n6794), .A(n10051), .ZN(P2_U3501) );
  INV_X1 U12630 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n15160) );
  NOR2_X1 U12631 ( .A1(n10064), .A2(n15160), .ZN(n10053) );
  AOI21_X1 U12632 ( .B1(n15160), .B2(n10064), .A(n10053), .ZN(n10058) );
  INV_X1 U12633 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n15402) );
  NOR2_X1 U12634 ( .A1(n10054), .A2(n15400), .ZN(n13941) );
  MUX2_X1 U12635 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n15402), .S(n13942), .Z(
        n10055) );
  OAI21_X1 U12636 ( .B1(n13947), .B2(n13941), .A(n10055), .ZN(n13945) );
  OAI21_X1 U12637 ( .B1(n15402), .B2(n13939), .A(n13945), .ZN(n10057) );
  NOR2_X1 U12638 ( .A1(n10064), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10056) );
  AOI211_X1 U12639 ( .C1(n10064), .C2(P2_REG1_REG_12__SCAN_IN), .A(n10056), 
        .B(n10057), .ZN(n10999) );
  AOI21_X1 U12640 ( .B1(n10058), .B2(n10057), .A(n10999), .ZN(n10073) );
  INV_X1 U12641 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10061) );
  MUX2_X1 U12642 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10061), .S(n13942), .Z(
        n13935) );
  NAND2_X1 U12643 ( .A1(n13936), .A2(n13935), .ZN(n13934) );
  NAND2_X1 U12644 ( .A1(n13939), .A2(n10061), .ZN(n10066) );
  INV_X1 U12645 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U12646 ( .A1(n10064), .A2(n10063), .ZN(n10062) );
  OAI21_X1 U12647 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(n10065) );
  INV_X1 U12648 ( .A(n10065), .ZN(n10067) );
  AOI21_X1 U12649 ( .B1(n13934), .B2(n10066), .A(n10067), .ZN(n10993) );
  AND3_X1 U12650 ( .A1(n13934), .A2(n10067), .A3(n10066), .ZN(n10068) );
  OAI21_X1 U12651 ( .B1(n10993), .B2(n10068), .A(n15319), .ZN(n10072) );
  NOR2_X1 U12652 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13485), .ZN(n10070) );
  NOR2_X1 U12653 ( .A1(n15311), .A2(n11000), .ZN(n10069) );
  AOI211_X1 U12654 ( .C1(n15314), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n10070), 
        .B(n10069), .ZN(n10071) );
  OAI211_X1 U12655 ( .C1(n10073), .C2(n15269), .A(n10072), .B(n10071), .ZN(
        P2_U3226) );
  OAI22_X1 U12656 ( .A1(n7265), .A2(P3_U3151), .B1(SI_17_), .B2(n12609), .ZN(
        n10074) );
  AOI21_X1 U12657 ( .B1(n10075), .B2(n13749), .A(n10074), .ZN(P3_U3278) );
  INV_X1 U12658 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U12659 ( .A1(n11450), .A2(n11434), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n10939), .ZN(n10081) );
  OR2_X1 U12660 ( .A1(n10077), .A2(n10076), .ZN(n10078) );
  OAI21_X1 U12661 ( .B1(n10079), .B2(n11501), .A(n10078), .ZN(n10080) );
  NOR2_X1 U12662 ( .A1(n10081), .A2(n10080), .ZN(n10938) );
  AOI21_X1 U12663 ( .B1(n10081), .B2(n10080), .A(n10938), .ZN(n10090) );
  NAND2_X1 U12664 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n11741)
         );
  NAND2_X1 U12665 ( .A1(n15199), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n10082) );
  OAI211_X1 U12666 ( .C1(n15212), .C2(n10939), .A(n11741), .B(n10082), .ZN(
        n10083) );
  INV_X1 U12667 ( .A(n10083), .ZN(n10089) );
  NAND2_X1 U12668 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n11424), .ZN(n10085) );
  NAND2_X1 U12669 ( .A1(n10085), .A2(n10084), .ZN(n10087) );
  INV_X1 U12670 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11461) );
  XNOR2_X1 U12671 ( .A(n11450), .B(n11461), .ZN(n10086) );
  NAND2_X1 U12672 ( .A1(n10086), .A2(n10087), .ZN(n10932) );
  OAI211_X1 U12673 ( .C1(n10087), .C2(n10086), .A(n10932), .B(n14576), .ZN(
        n10088) );
  OAI211_X1 U12674 ( .C1(n10090), .C2(n15208), .A(n10089), .B(n10088), .ZN(
        P1_U3257) );
  NAND2_X1 U12675 ( .A1(n10095), .A2(n10091), .ZN(n10092) );
  INV_X1 U12676 ( .A(n10095), .ZN(n10097) );
  NAND2_X1 U12677 ( .A1(n10097), .A2(n10096), .ZN(n10098) );
  AOI22_X1 U12678 ( .A1(n11845), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11844), 
        .B2(n10101), .ZN(n10102) );
  AOI22_X1 U12679 ( .A1(n12709), .A2(n14472), .B1(n10103), .B2(n12330), .ZN(
        n10108) );
  NAND2_X1 U12680 ( .A1(n12708), .A2(n12330), .ZN(n10105) );
  NAND2_X1 U12681 ( .A1(n10103), .A2(n14472), .ZN(n10104) );
  NAND2_X1 U12682 ( .A1(n10105), .A2(n10104), .ZN(n10106) );
  XNOR2_X1 U12683 ( .A(n10106), .B(n11728), .ZN(n10107) );
  AND2_X1 U12684 ( .A1(n10108), .A2(n10107), .ZN(n10498) );
  INV_X1 U12685 ( .A(n10498), .ZN(n10111) );
  INV_X1 U12686 ( .A(n10107), .ZN(n10110) );
  INV_X1 U12687 ( .A(n10108), .ZN(n10109) );
  NAND2_X1 U12688 ( .A1(n10110), .A2(n10109), .ZN(n10497) );
  NAND2_X1 U12689 ( .A1(n10111), .A2(n10497), .ZN(n10112) );
  XNOR2_X1 U12690 ( .A(n10499), .B(n10112), .ZN(n10128) );
  NAND2_X1 U12691 ( .A1(n11985), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10122) );
  INV_X1 U12692 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10113) );
  OR2_X1 U12693 ( .A1(n11944), .A2(n10113), .ZN(n10121) );
  INV_X1 U12694 ( .A(n10412), .ZN(n10118) );
  INV_X1 U12695 ( .A(n10114), .ZN(n10116) );
  INV_X1 U12696 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10115) );
  NAND2_X1 U12697 ( .A1(n10116), .A2(n10115), .ZN(n10117) );
  NAND2_X1 U12698 ( .A1(n10118), .A2(n10117), .ZN(n14431) );
  OR2_X1 U12699 ( .A1(n11986), .A2(n14431), .ZN(n10120) );
  OR2_X1 U12700 ( .A1(n12454), .A2(n9629), .ZN(n10119) );
  NAND4_X1 U12701 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n14471) );
  NAND2_X1 U12702 ( .A1(n14438), .A2(n14471), .ZN(n10124) );
  NAND2_X1 U12703 ( .A1(n10124), .A2(n10123), .ZN(n10126) );
  INV_X1 U12704 ( .A(n12330), .ZN(n15243) );
  INV_X1 U12705 ( .A(n9832), .ZN(n14450) );
  INV_X1 U12706 ( .A(n14447), .ZN(n11567) );
  OAI22_X1 U12707 ( .A1(n15243), .A2(n14450), .B1(n11567), .B2(n12326), .ZN(
        n10125) );
  AOI211_X1 U12708 ( .C1(n11071), .C2(n14454), .A(n10126), .B(n10125), .ZN(
        n10127) );
  OAI21_X1 U12709 ( .B1(n10128), .B2(n14456), .A(n10127), .ZN(P1_U3227) );
  INV_X1 U12710 ( .A(n10129), .ZN(n10133) );
  INV_X1 U12711 ( .A(n10131), .ZN(n10132) );
  AOI21_X1 U12712 ( .B1(n10133), .B2(n10130), .A(n10132), .ZN(n10141) );
  INV_X1 U12713 ( .A(n15107), .ZN(n13888) );
  INV_X1 U12714 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10134) );
  OAI22_X1 U12715 ( .A1(n13888), .A2(n9900), .B1(n11806), .B2(n10134), .ZN(
        n10137) );
  NOR2_X1 U12716 ( .A1(n13883), .A2(n10135), .ZN(n10136) );
  AOI211_X1 U12717 ( .C1(n12009), .C2(n9026), .A(n10137), .B(n10136), .ZN(
        n10140) );
  NAND3_X1 U12718 ( .A1(n13875), .A2(n10138), .A3(n10130), .ZN(n10139) );
  OAI211_X1 U12719 ( .C1(n10141), .C2(n13872), .A(n10140), .B(n10139), .ZN(
        P2_U3194) );
  NAND2_X1 U12720 ( .A1(n10143), .A2(n10142), .ZN(n15353) );
  NAND2_X1 U12721 ( .A1(n9899), .A2(n15125), .ZN(n10145) );
  AND2_X1 U12722 ( .A1(n9901), .A2(n14027), .ZN(n10144) );
  AOI21_X1 U12723 ( .B1(n15357), .B2(n10145), .A(n10144), .ZN(n15354) );
  OAI21_X1 U12724 ( .B1(n10146), .B2(n15353), .A(n15354), .ZN(n10147) );
  INV_X1 U12725 ( .A(n14147), .ZN(n15329) );
  AOI22_X1 U12726 ( .A1(n14163), .A2(n10147), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n15329), .ZN(n10150) );
  NAND2_X1 U12727 ( .A1(n14168), .A2(n15357), .ZN(n10149) );
  OAI211_X1 U12728 ( .C1(n14163), .C2(n10151), .A(n10150), .B(n10149), .ZN(
        P2_U3265) );
  NAND2_X1 U12729 ( .A1(n10152), .A2(n15559), .ZN(n10153) );
  OR2_X1 U12730 ( .A1(n12200), .A2(n10153), .ZN(n10155) );
  OR2_X1 U12731 ( .A1(n15493), .A2(n15494), .ZN(n10154) );
  NAND2_X1 U12732 ( .A1(n10155), .A2(n10154), .ZN(n10526) );
  INV_X1 U12733 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10174) );
  OAI22_X1 U12734 ( .A1(n13689), .A2(n10524), .B1(n15603), .B2(n10174), .ZN(
        n10156) );
  AOI21_X1 U12735 ( .B1(n10526), .B2(n15603), .A(n10156), .ZN(n10157) );
  INV_X1 U12736 ( .A(n10157), .ZN(P3_U3459) );
  XNOR2_X1 U12737 ( .A(n10687), .B(n10158), .ZN(n10368) );
  NAND2_X1 U12738 ( .A1(n13913), .A2(n9914), .ZN(n10369) );
  XNOR2_X1 U12739 ( .A(n10368), .B(n10369), .ZN(n10162) );
  AND2_X1 U12740 ( .A1(n10162), .A2(n10159), .ZN(n10160) );
  OAI21_X1 U12741 ( .B1(n10162), .B2(n10161), .A(n12013), .ZN(n10172) );
  INV_X1 U12742 ( .A(n10162), .ZN(n10164) );
  NAND3_X1 U12743 ( .A1(n13875), .A2(n10164), .A3(n10163), .ZN(n10166) );
  AOI21_X1 U12744 ( .B1(n10166), .B2(n13881), .A(n10165), .ZN(n10171) );
  INV_X1 U12745 ( .A(n10687), .ZN(n15367) );
  AOI22_X1 U12746 ( .A1(n10167), .A2(n13912), .B1(n13855), .B2(n10686), .ZN(
        n10169) );
  OAI211_X1 U12747 ( .C1(n15367), .C2(n13888), .A(n10169), .B(n10168), .ZN(
        n10170) );
  AOI211_X1 U12748 ( .C1(n15104), .C2(n10172), .A(n10171), .B(n10170), .ZN(
        n10173) );
  INV_X1 U12749 ( .A(n10173), .ZN(P2_U3202) );
  INV_X1 U12750 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10194) );
  MUX2_X1 U12751 ( .A(n10194), .B(n10174), .S(n6586), .Z(n15405) );
  AND2_X1 U12752 ( .A1(n15405), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15411) );
  INV_X1 U12753 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10175) );
  OR2_X1 U12754 ( .A1(n6586), .A2(n10175), .ZN(n10177) );
  NAND2_X1 U12755 ( .A1(n6586), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10176) );
  NAND2_X1 U12756 ( .A1(n10177), .A2(n10176), .ZN(n10226) );
  XOR2_X1 U12757 ( .A(n10196), .B(n10226), .Z(n10229) );
  XOR2_X1 U12758 ( .A(n15411), .B(n10229), .Z(n10203) );
  NAND2_X1 U12759 ( .A1(P3_U3897), .A2(n8297), .ZN(n15406) );
  NAND2_X1 U12760 ( .A1(n10180), .A2(n12183), .ZN(n10178) );
  NAND2_X1 U12761 ( .A1(n6602), .A2(n10178), .ZN(n10191) );
  INV_X1 U12762 ( .A(n10180), .ZN(n10181) );
  NAND2_X1 U12763 ( .A1(n10181), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12235) );
  AND2_X1 U12764 ( .A1(n10182), .A2(n12235), .ZN(n10189) );
  OR2_X1 U12765 ( .A1(n10191), .A2(n10189), .ZN(n10198) );
  INV_X1 U12766 ( .A(n10198), .ZN(n10183) );
  MUX2_X1 U12767 ( .A(P3_U3897), .B(n10183), .S(n8297), .Z(n15421) );
  INV_X1 U12768 ( .A(n10196), .ZN(n10228) );
  INV_X1 U12769 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15583) );
  NAND2_X1 U12770 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10184), .ZN(n10185) );
  INV_X1 U12771 ( .A(n10185), .ZN(n10186) );
  OR2_X1 U12772 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10185), .ZN(n10204) );
  OAI21_X1 U12773 ( .B1(n10196), .B2(n10186), .A(n10204), .ZN(n10188) );
  OR2_X1 U12774 ( .A1(n10188), .A2(n15583), .ZN(n10205) );
  INV_X1 U12775 ( .A(n10205), .ZN(n10187) );
  AOI21_X1 U12776 ( .B1(n15583), .B2(n10188), .A(n10187), .ZN(n10193) );
  INV_X1 U12777 ( .A(n10189), .ZN(n10190) );
  AOI22_X1 U12778 ( .A1(n15417), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10192) );
  OAI21_X1 U12779 ( .B1(n15407), .B2(n10193), .A(n10192), .ZN(n10201) );
  NOR2_X1 U12780 ( .A1(n10194), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10195) );
  OR3_X1 U12781 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n10194), .ZN(n10211) );
  AOI21_X1 U12782 ( .B1(n10212), .B2(n10199), .A(n15408), .ZN(n10200) );
  AOI211_X1 U12783 ( .C1(n15421), .C2(n10228), .A(n10201), .B(n10200), .ZN(
        n10202) );
  OAI21_X1 U12784 ( .B1(n10203), .B2(n15406), .A(n10202), .ZN(P3_U3183) );
  INV_X1 U12785 ( .A(n15421), .ZN(n12916) );
  INV_X1 U12786 ( .A(n6753), .ZN(n10286) );
  INV_X1 U12787 ( .A(n15407), .ZN(n15429) );
  INV_X1 U12788 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15589) );
  MUX2_X1 U12789 ( .A(n15589), .B(P3_REG1_REG_4__SCAN_IN), .S(n10298), .Z(
        n10209) );
  INV_X1 U12790 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15585) );
  MUX2_X1 U12791 ( .A(n15585), .B(P3_REG1_REG_2__SCAN_IN), .S(n10252), .Z(
        n10242) );
  NAND2_X1 U12792 ( .A1(n10205), .A2(n10204), .ZN(n10241) );
  NAND2_X1 U12793 ( .A1(n10242), .A2(n10241), .ZN(n10240) );
  INV_X1 U12794 ( .A(n10252), .ZN(n10230) );
  NAND2_X1 U12795 ( .A1(n10230), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10206) );
  INV_X1 U12796 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15587) );
  AND2_X1 U12797 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10794) );
  INV_X1 U12798 ( .A(n10794), .ZN(n10210) );
  OAI21_X1 U12799 ( .B1(n15414), .B2(n7124), .A(n10210), .ZN(n10219) );
  INV_X1 U12800 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15510) );
  MUX2_X1 U12801 ( .A(n15510), .B(P3_REG2_REG_2__SCAN_IN), .S(n10252), .Z(
        n10246) );
  NAND2_X1 U12802 ( .A1(n10246), .A2(n10245), .ZN(n10244) );
  NAND2_X1 U12803 ( .A1(n10230), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10213) );
  INV_X1 U12804 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n15487) );
  NOR2_X1 U12805 ( .A1(n15424), .A2(n10214), .ZN(n10216) );
  INV_X1 U12806 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10297) );
  MUX2_X1 U12807 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n10297), .S(n10298), .Z(
        n10215) );
  NAND2_X1 U12808 ( .A1(n10216), .A2(n10215), .ZN(n10217) );
  AOI21_X1 U12809 ( .B1(n10300), .B2(n10217), .A(n15408), .ZN(n10218) );
  AOI211_X1 U12810 ( .C1(n15429), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        n10237) );
  MUX2_X1 U12811 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n6587), .Z(n10287) );
  XNOR2_X1 U12812 ( .A(n10287), .B(n6753), .ZN(n10234) );
  OR2_X1 U12813 ( .A1(n6587), .A2(n15487), .ZN(n10223) );
  NAND2_X1 U12814 ( .A1(n6587), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10222) );
  NAND2_X1 U12815 ( .A1(n10223), .A2(n10222), .ZN(n10225) );
  OR2_X1 U12816 ( .A1(n10224), .A2(n10225), .ZN(n10232) );
  XNOR2_X1 U12817 ( .A(n10225), .B(n7258), .ZN(n15419) );
  INV_X1 U12818 ( .A(n10226), .ZN(n10227) );
  MUX2_X1 U12819 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n6587), .Z(n10231) );
  XOR2_X1 U12820 ( .A(n10252), .B(n10231), .Z(n10239) );
  NAND2_X1 U12821 ( .A1(n15419), .A2(n15420), .ZN(n15418) );
  NAND2_X1 U12822 ( .A1(n10232), .A2(n15418), .ZN(n10233) );
  NAND2_X1 U12823 ( .A1(n10234), .A2(n10233), .ZN(n10285) );
  OAI21_X1 U12824 ( .B1(n10234), .B2(n10233), .A(n10285), .ZN(n10235) );
  NAND2_X1 U12825 ( .A1(n10235), .A2(n15422), .ZN(n10236) );
  OAI211_X1 U12826 ( .C1(n12916), .C2(n10286), .A(n10237), .B(n10236), .ZN(
        P3_U3186) );
  XOR2_X1 U12827 ( .A(n10239), .B(n10238), .Z(n10254) );
  OAI21_X1 U12828 ( .B1(n10242), .B2(n10241), .A(n10240), .ZN(n10243) );
  NAND2_X1 U12829 ( .A1(n15429), .A2(n10243), .ZN(n10250) );
  AOI22_X1 U12830 ( .A1(n15417), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10249) );
  OAI21_X1 U12831 ( .B1(n10246), .B2(n10245), .A(n10244), .ZN(n10247) );
  NAND2_X1 U12832 ( .A1(n15425), .A2(n10247), .ZN(n10248) );
  NAND3_X1 U12833 ( .A1(n10250), .A2(n10249), .A3(n10248), .ZN(n10251) );
  AOI21_X1 U12834 ( .B1(n10252), .B2(n15421), .A(n10251), .ZN(n10253) );
  OAI21_X1 U12835 ( .B1(n10254), .B2(n15406), .A(n10253), .ZN(P3_U3184) );
  NAND3_X1 U12836 ( .A1(n10257), .A2(n10256), .A3(n10255), .ZN(n10259) );
  NOR2_X1 U12837 ( .A1(n10259), .A2(n10258), .ZN(n10261) );
  NAND2_X1 U12838 ( .A1(n10261), .A2(n10260), .ZN(n10263) );
  NAND2_X1 U12839 ( .A1(n10263), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10262) );
  MUX2_X1 U12840 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10262), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n10264) );
  AND2_X1 U12841 ( .A1(n10264), .A2(n10494), .ZN(n11642) );
  INV_X1 U12842 ( .A(n11642), .ZN(n15211) );
  INV_X1 U12843 ( .A(n11641), .ZN(n10266) );
  OAI222_X1 U12844 ( .A1(n15211), .A2(P1_U3086), .B1(n15030), .B2(n10266), 
        .C1(n10265), .C2(n15024), .ZN(P1_U3340) );
  INV_X1 U12845 ( .A(n15301), .ZN(n11279) );
  OAI222_X1 U12846 ( .A1(n14312), .A2(n7248), .B1(n10596), .B2(n10266), .C1(
        P2_U3088), .C2(n11279), .ZN(P2_U3312) );
  OR2_X1 U12847 ( .A1(n10267), .A2(n6953), .ZN(n10268) );
  NAND2_X1 U12848 ( .A1(n10269), .A2(n10268), .ZN(n10603) );
  NAND2_X1 U12849 ( .A1(n10684), .A2(n10372), .ZN(n10270) );
  NAND2_X1 U12850 ( .A1(n10270), .A2(n10037), .ZN(n10271) );
  NOR2_X1 U12851 ( .A1(n10543), .A2(n10271), .ZN(n10597) );
  NAND3_X1 U12852 ( .A1(n10676), .A2(n6953), .A3(n10272), .ZN(n10273) );
  NAND2_X1 U12853 ( .A1(n10547), .A2(n10273), .ZN(n10277) );
  NAND2_X1 U12854 ( .A1(n13913), .A2(n14025), .ZN(n10275) );
  NAND2_X1 U12855 ( .A1(n13911), .A2(n14027), .ZN(n10274) );
  NAND2_X1 U12856 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  AOI21_X1 U12857 ( .B1(n10277), .B2(n6580), .A(n10276), .ZN(n10279) );
  NAND2_X1 U12858 ( .A1(n10603), .A2(n10551), .ZN(n10278) );
  NAND2_X1 U12859 ( .A1(n10279), .A2(n10278), .ZN(n10600) );
  AOI211_X1 U12860 ( .C1(n15390), .C2(n10603), .A(n10597), .B(n10600), .ZN(
        n10284) );
  INV_X1 U12861 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10280) );
  OAI22_X1 U12862 ( .A1(n14287), .A2(n12003), .B1(n15393), .B2(n10280), .ZN(
        n10281) );
  INV_X1 U12863 ( .A(n10281), .ZN(n10282) );
  OAI21_X1 U12864 ( .B1(n10284), .B2(n15391), .A(n10282), .ZN(P2_U3445) );
  AOI22_X1 U12865 ( .A1(n14248), .A2(n10372), .B1(n6794), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n10283) );
  OAI21_X1 U12866 ( .B1(n10284), .B2(n6794), .A(n10283), .ZN(P2_U3504) );
  OAI21_X1 U12867 ( .B1(n10287), .B2(n10286), .A(n10285), .ZN(n10429) );
  OR2_X1 U12868 ( .A1(n6587), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n10289) );
  NAND2_X1 U12869 ( .A1(n6587), .A2(n7050), .ZN(n10288) );
  NAND2_X1 U12870 ( .A1(n10289), .A2(n10288), .ZN(n10290) );
  AND2_X1 U12871 ( .A1(n10290), .A2(n10307), .ZN(n10427) );
  INV_X1 U12872 ( .A(n10427), .ZN(n10292) );
  INV_X1 U12873 ( .A(n10290), .ZN(n10291) );
  INV_X1 U12874 ( .A(n10307), .ZN(n10443) );
  NAND2_X1 U12875 ( .A1(n10291), .A2(n10443), .ZN(n10428) );
  NAND2_X1 U12876 ( .A1(n10292), .A2(n10428), .ZN(n10293) );
  XNOR2_X1 U12877 ( .A(n10429), .B(n10293), .ZN(n10309) );
  OR2_X1 U12878 ( .A1(n6753), .A2(n15589), .ZN(n10294) );
  XNOR2_X1 U12879 ( .A(n10436), .B(n10307), .ZN(n10295) );
  OAI21_X1 U12880 ( .B1(n10295), .B2(P3_REG1_REG_5__SCAN_IN), .A(n10438), .ZN(
        n10296) );
  NAND2_X1 U12881 ( .A1(n15429), .A2(n10296), .ZN(n10305) );
  NOR2_X1 U12882 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13440), .ZN(n10914) );
  AOI21_X1 U12883 ( .B1(n15417), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n10914), .ZN(
        n10304) );
  OR2_X1 U12884 ( .A1(n6753), .A2(n10297), .ZN(n10299) );
  OAI21_X1 U12885 ( .B1(n10301), .B2(P3_REG2_REG_5__SCAN_IN), .A(n6874), .ZN(
        n10302) );
  NAND2_X1 U12886 ( .A1(n15425), .A2(n10302), .ZN(n10303) );
  NAND3_X1 U12887 ( .A1(n10305), .A2(n10304), .A3(n10303), .ZN(n10306) );
  AOI21_X1 U12888 ( .B1(n10307), .B2(n15421), .A(n10306), .ZN(n10308) );
  OAI21_X1 U12889 ( .B1(n15406), .B2(n10309), .A(n10308), .ZN(P3_U3187) );
  NAND2_X1 U12890 ( .A1(n12307), .A2(n12308), .ZN(n10310) );
  NAND2_X1 U12891 ( .A1(n10330), .A2(n10328), .ZN(n10329) );
  NAND2_X1 U12892 ( .A1(n12315), .A2(n12314), .ZN(n10312) );
  XNOR2_X1 U12893 ( .A(n15236), .B(n10331), .ZN(n12317) );
  INV_X1 U12894 ( .A(n12317), .ZN(n12491) );
  NAND2_X1 U12895 ( .A1(n15236), .A2(n10331), .ZN(n10313) );
  XNOR2_X1 U12896 ( .A(n12325), .B(n12326), .ZN(n12493) );
  INV_X1 U12897 ( .A(n12493), .ZN(n10322) );
  OAI21_X1 U12898 ( .B1(n10314), .B2(n10322), .A(n10400), .ZN(n10829) );
  INV_X1 U12899 ( .A(n10850), .ZN(n10315) );
  AOI211_X1 U12900 ( .C1(n12324), .C2(n10315), .A(n14828), .B(n11070), .ZN(
        n10835) );
  INV_X1 U12901 ( .A(n14472), .ZN(n10417) );
  AND2_X1 U12902 ( .A1(n12307), .A2(n14844), .ZN(n10316) );
  INV_X1 U12903 ( .A(n10332), .ZN(n10317) );
  NAND2_X1 U12904 ( .A1(n12315), .A2(n12312), .ZN(n10318) );
  NAND2_X1 U12905 ( .A1(n10843), .A2(n12317), .ZN(n10842) );
  NOR2_X1 U12906 ( .A1(n15236), .A2(n14474), .ZN(n12319) );
  INV_X1 U12907 ( .A(n12319), .ZN(n10319) );
  NAND2_X1 U12908 ( .A1(n10842), .A2(n10319), .ZN(n10320) );
  INV_X1 U12909 ( .A(n10320), .ZN(n10323) );
  INV_X1 U12910 ( .A(n11063), .ZN(n10321) );
  AOI21_X1 U12911 ( .B1(n10323), .B2(n10322), .A(n10321), .ZN(n10324) );
  OAI222_X1 U12912 ( .A1(n14826), .A2(n10417), .B1(n14824), .B2(n10331), .C1(
        n15228), .C2(n10324), .ZN(n10831) );
  AOI211_X1 U12913 ( .C1(n15256), .C2(n10829), .A(n10835), .B(n10831), .ZN(
        n10344) );
  INV_X1 U12914 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10325) );
  OAI22_X1 U12915 ( .A1(n15011), .A2(n12325), .B1(n15259), .B2(n10325), .ZN(
        n10326) );
  INV_X1 U12916 ( .A(n10326), .ZN(n10327) );
  OAI21_X1 U12917 ( .B1(n10344), .B2(n15257), .A(n10327), .ZN(P1_U3471) );
  OAI21_X1 U12918 ( .B1(n10330), .B2(n10328), .A(n10329), .ZN(n10337) );
  INV_X1 U12919 ( .A(n10337), .ZN(n10863) );
  OAI22_X1 U12920 ( .A1(n10331), .A2(n14826), .B1(n12307), .B2(n14824), .ZN(
        n10336) );
  NAND2_X1 U12921 ( .A1(n10332), .A2(n10328), .ZN(n10333) );
  AOI21_X1 U12922 ( .B1(n10334), .B2(n10333), .A(n15228), .ZN(n10335) );
  AOI211_X1 U12923 ( .C1(n14629), .C2(n10337), .A(n10336), .B(n10335), .ZN(
        n10856) );
  NAND2_X1 U12924 ( .A1(n10338), .A2(n12312), .ZN(n10339) );
  NAND2_X1 U12925 ( .A1(n10339), .A2(n14888), .ZN(n10340) );
  OR2_X1 U12926 ( .A1(n10340), .A2(n10849), .ZN(n10859) );
  OAI211_X1 U12927 ( .C1(n10863), .C2(n14946), .A(n10856), .B(n10859), .ZN(
        n10347) );
  INV_X1 U12928 ( .A(n10347), .ZN(n10342) );
  AOI22_X1 U12929 ( .A1(n14900), .A2(n12312), .B1(n15265), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n10341) );
  OAI21_X1 U12930 ( .B1(n10342), .B2(n15265), .A(n10341), .ZN(P1_U3530) );
  AOI22_X1 U12931 ( .A1(n14900), .A2(n12324), .B1(n15265), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n10343) );
  OAI21_X1 U12932 ( .B1(n10344), .B2(n15265), .A(n10343), .ZN(P1_U3532) );
  INV_X1 U12933 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10345) );
  OAI22_X1 U12934 ( .A1(n15011), .A2(n12314), .B1(n15259), .B2(n10345), .ZN(
        n10346) );
  AOI21_X1 U12935 ( .B1(n10347), .B2(n15259), .A(n10346), .ZN(n10348) );
  INV_X1 U12936 ( .A(n10348), .ZN(P1_U3465) );
  INV_X1 U12937 ( .A(n10349), .ZN(n10351) );
  OAI222_X1 U12938 ( .A1(n13756), .A2(n10351), .B1(n12609), .B2(n10350), .C1(
        n13054), .C2(P3_U3151), .ZN(P3_U3277) );
  INV_X1 U12939 ( .A(n10532), .ZN(n10367) );
  INV_X1 U12940 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15526) );
  NAND2_X1 U12941 ( .A1(n10784), .A2(n10352), .ZN(n10353) );
  OAI21_X1 U12942 ( .B1(n10357), .B2(n12734), .A(n10356), .ZN(n10358) );
  INV_X1 U12943 ( .A(n15520), .ZN(n12061) );
  NAND3_X1 U12944 ( .A1(n12061), .A2(n10359), .A3(n6801), .ZN(n10360) );
  OAI211_X1 U12945 ( .C1(n10361), .C2(n15512), .A(n10531), .B(n10360), .ZN(
        n10362) );
  NAND2_X1 U12946 ( .A1(n10362), .A2(n12874), .ZN(n10366) );
  INV_X1 U12947 ( .A(n12880), .ZN(n12864) );
  OAI22_X1 U12948 ( .A1(n10629), .A2(n12867), .B1(n8254), .B2(n12885), .ZN(
        n10364) );
  AOI21_X1 U12949 ( .B1(n12864), .B2(n15516), .A(n10364), .ZN(n10365) );
  OAI211_X1 U12950 ( .C1(n10367), .C2(n15526), .A(n10366), .B(n10365), .ZN(
        P3_U3162) );
  INV_X1 U12951 ( .A(n10368), .ZN(n12010) );
  NAND2_X1 U12952 ( .A1(n12010), .A2(n10369), .ZN(n10370) );
  XNOR2_X1 U12953 ( .A(n10372), .B(n12592), .ZN(n10374) );
  NAND2_X1 U12954 ( .A1(n13912), .A2(n13997), .ZN(n10375) );
  XNOR2_X1 U12955 ( .A(n10374), .B(n10375), .ZN(n12012) );
  INV_X1 U12956 ( .A(n10374), .ZN(n10376) );
  NAND2_X1 U12957 ( .A1(n10376), .A2(n10375), .ZN(n10377) );
  XNOR2_X1 U12958 ( .A(n10655), .B(n12592), .ZN(n10378) );
  AND2_X1 U12959 ( .A1(n13911), .A2(n13997), .ZN(n10379) );
  NAND2_X1 U12960 ( .A1(n10378), .A2(n10379), .ZN(n10385) );
  INV_X1 U12961 ( .A(n10378), .ZN(n10384) );
  INV_X1 U12962 ( .A(n10379), .ZN(n10380) );
  NAND2_X1 U12963 ( .A1(n10384), .A2(n10380), .ZN(n10381) );
  NAND2_X1 U12964 ( .A1(n10385), .A2(n10381), .ZN(n10565) );
  NAND2_X1 U12965 ( .A1(n13910), .A2(n13997), .ZN(n10638) );
  INV_X1 U12966 ( .A(n10387), .ZN(n10383) );
  AOI21_X1 U12967 ( .B1(n10386), .B2(n10383), .A(n13872), .ZN(n10390) );
  INV_X1 U12968 ( .A(n13875), .ZN(n13817) );
  NOR3_X1 U12969 ( .A1(n13817), .A2(n12006), .A3(n10384), .ZN(n10389) );
  NAND2_X1 U12970 ( .A1(n10386), .A2(n10385), .ZN(n10388) );
  OAI21_X1 U12971 ( .B1(n10390), .B2(n10389), .A(n10641), .ZN(n10399) );
  NOR2_X1 U12972 ( .A1(n15111), .A2(n10391), .ZN(n10397) );
  NAND2_X1 U12973 ( .A1(n13911), .A2(n14025), .ZN(n10393) );
  NAND2_X1 U12974 ( .A1(n13909), .A2(n14027), .ZN(n10392) );
  NAND2_X1 U12975 ( .A1(n10393), .A2(n10392), .ZN(n10612) );
  INV_X1 U12976 ( .A(n10612), .ZN(n10395) );
  OAI21_X1 U12977 ( .B1(n13853), .B2(n10395), .A(n10394), .ZN(n10396) );
  AOI211_X1 U12978 ( .C1(n15326), .C2(n15107), .A(n10397), .B(n10396), .ZN(
        n10398) );
  NAND2_X1 U12979 ( .A1(n10399), .A2(n10398), .ZN(P2_U3185) );
  INV_X1 U12980 ( .A(n14946), .ZN(n15248) );
  XNOR2_X1 U12981 ( .A(n12330), .B(n14472), .ZN(n12492) );
  INV_X1 U12982 ( .A(n12492), .ZN(n11062) );
  NAND2_X1 U12983 ( .A1(n15243), .A2(n10417), .ZN(n10401) );
  OR2_X1 U12984 ( .A1(n10402), .A2(n11448), .ZN(n10405) );
  AOI22_X1 U12985 ( .A1(n11845), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11844), 
        .B2(n10403), .ZN(n10404) );
  NAND2_X1 U12986 ( .A1(n10405), .A2(n10404), .ZN(n14429) );
  XNOR2_X1 U12987 ( .A(n14429), .B(n14471), .ZN(n12495) );
  INV_X1 U12988 ( .A(n12495), .ZN(n10410) );
  OAI21_X1 U12989 ( .B1(n10406), .B2(n10410), .A(n10461), .ZN(n10816) );
  NAND2_X1 U12990 ( .A1(n15243), .A2(n11070), .ZN(n11069) );
  AOI21_X1 U12991 ( .B1(n11069), .B2(n14429), .A(n14828), .ZN(n10407) );
  AND2_X1 U12992 ( .A1(n10474), .A2(n10407), .ZN(n10825) );
  INV_X1 U12993 ( .A(n12326), .ZN(n14473) );
  OR2_X1 U12994 ( .A1(n12325), .A2(n14473), .ZN(n11061) );
  NAND2_X1 U12995 ( .A1(n11063), .A2(n11061), .ZN(n10408) );
  NAND2_X1 U12996 ( .A1(n10408), .A2(n12492), .ZN(n11065) );
  NAND2_X1 U12997 ( .A1(n12330), .A2(n10417), .ZN(n10409) );
  XNOR2_X1 U12998 ( .A(n10457), .B(n10410), .ZN(n10420) );
  NAND2_X1 U12999 ( .A1(n11985), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10416) );
  INV_X1 U13000 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10411) );
  OR2_X1 U13001 ( .A1(n11944), .A2(n10411), .ZN(n10415) );
  NAND2_X1 U13002 ( .A1(n10412), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10466) );
  OAI21_X1 U13003 ( .B1(n10412), .B2(P1_REG3_REG_7__SCAN_IN), .A(n10466), .ZN(
        n10953) );
  OR2_X1 U13004 ( .A1(n11986), .A2(n10953), .ZN(n10414) );
  OR2_X1 U13005 ( .A1(n12454), .A2(n9631), .ZN(n10413) );
  NAND4_X1 U13006 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n14470) );
  INV_X1 U13007 ( .A(n14470), .ZN(n10513) );
  OAI22_X1 U13008 ( .A1(n10417), .A2(n14824), .B1(n10513), .B2(n14826), .ZN(
        n10418) );
  AOI21_X1 U13009 ( .B1(n10816), .B2(n14629), .A(n10418), .ZN(n10419) );
  OAI21_X1 U13010 ( .B1(n15228), .B2(n10420), .A(n10419), .ZN(n10820) );
  AOI211_X1 U13011 ( .C1(n15248), .C2(n10816), .A(n10825), .B(n10820), .ZN(
        n10424) );
  OAI22_X1 U13012 ( .A1(n15011), .A2(n12341), .B1(n15259), .B2(n10113), .ZN(
        n10421) );
  INV_X1 U13013 ( .A(n10421), .ZN(n10422) );
  OAI21_X1 U13014 ( .B1(n10424), .B2(n15257), .A(n10422), .ZN(P1_U3477) );
  AOI22_X1 U13015 ( .A1(n14900), .A2(n14429), .B1(n15265), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n10423) );
  OAI21_X1 U13016 ( .B1(n10424), .B2(n15265), .A(n10423), .ZN(P1_U3534) );
  OAI222_X1 U13017 ( .A1(n13060), .A2(P3_U3151), .B1(n13756), .B2(n10426), 
        .C1(n10425), .C2(n12609), .ZN(P3_U3276) );
  OR2_X1 U13018 ( .A1(n6587), .A2(n11076), .ZN(n10431) );
  NAND2_X1 U13019 ( .A1(n6587), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10430) );
  AND2_X1 U13020 ( .A1(n10431), .A2(n10430), .ZN(n10433) );
  AND2_X1 U13021 ( .A1(n10433), .A2(n10451), .ZN(n11086) );
  INV_X1 U13022 ( .A(n11086), .ZN(n10432) );
  OAI21_X1 U13023 ( .B1(n10451), .B2(n10433), .A(n10432), .ZN(n10434) );
  AOI21_X1 U13024 ( .B1(n10435), .B2(n10434), .A(n11085), .ZN(n10453) );
  NAND2_X1 U13025 ( .A1(n10436), .A2(n10443), .ZN(n10437) );
  INV_X1 U13026 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15592) );
  AOI22_X1 U13027 ( .A1(n10451), .A2(P3_REG1_REG_6__SCAN_IN), .B1(n15592), 
        .B2(n11093), .ZN(n10439) );
  AOI21_X1 U13028 ( .B1(n10440), .B2(n10439), .A(n11092), .ZN(n10442) );
  AND2_X1 U13029 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n11037) );
  AOI21_X1 U13030 ( .B1(n15417), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n11037), .ZN(
        n10441) );
  OAI21_X1 U13031 ( .B1(n15407), .B2(n10442), .A(n10441), .ZN(n10450) );
  AOI22_X1 U13032 ( .A1(n10451), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n11076), 
        .B2(n11093), .ZN(n10446) );
  AOI21_X1 U13033 ( .B1(n10447), .B2(n10446), .A(n11078), .ZN(n10448) );
  NOR2_X1 U13034 ( .A1(n15408), .A2(n10448), .ZN(n10449) );
  AOI211_X1 U13035 ( .C1(n15421), .C2(n10451), .A(n10450), .B(n10449), .ZN(
        n10452) );
  OAI21_X1 U13036 ( .B1(n10453), .B2(n15406), .A(n10452), .ZN(P3_U3188) );
  OR2_X1 U13037 ( .A1(n10454), .A2(n11448), .ZN(n10456) );
  AOI22_X1 U13038 ( .A1(n11845), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11844), 
        .B2(n14552), .ZN(n10455) );
  NAND2_X1 U13039 ( .A1(n10456), .A2(n10455), .ZN(n12345) );
  XNOR2_X1 U13040 ( .A(n12345), .B(n10513), .ZN(n12497) );
  INV_X1 U13041 ( .A(n14471), .ZN(n12340) );
  NAND2_X1 U13042 ( .A1(n10457), .A2(n14429), .ZN(n10458) );
  XOR2_X1 U13043 ( .A(n10569), .B(n12497), .Z(n10948) );
  OR2_X1 U13044 ( .A1(n14429), .A2(n14471), .ZN(n10460) );
  NAND2_X1 U13045 ( .A1(n10462), .A2(n12497), .ZN(n10575) );
  OAI21_X1 U13046 ( .B1(n10462), .B2(n12497), .A(n10575), .ZN(n10463) );
  INV_X1 U13047 ( .A(n10463), .ZN(n10958) );
  NAND2_X1 U13048 ( .A1(n14471), .A2(n14791), .ZN(n10473) );
  NAND2_X1 U13049 ( .A1(n11985), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10471) );
  INV_X1 U13050 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10464) );
  OR2_X1 U13051 ( .A1(n11944), .A2(n10464), .ZN(n10470) );
  INV_X1 U13052 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10465) );
  AND2_X1 U13053 ( .A1(n10466), .A2(n10465), .ZN(n10467) );
  NOR2_X1 U13054 ( .A1(n10466), .A2(n10465), .ZN(n10579) );
  OR2_X1 U13055 ( .A1(n10467), .A2(n10579), .ZN(n10969) );
  OR2_X1 U13056 ( .A1(n11986), .A2(n10969), .ZN(n10469) );
  OR2_X1 U13057 ( .A1(n12454), .A2(n9632), .ZN(n10468) );
  NAND4_X1 U13058 ( .A1(n10471), .A2(n10470), .A3(n10469), .A4(n10468), .ZN(
        n14469) );
  NAND2_X1 U13059 ( .A1(n14469), .A2(n14850), .ZN(n10472) );
  NAND2_X1 U13060 ( .A1(n10473), .A2(n10472), .ZN(n10517) );
  INV_X1 U13061 ( .A(n10517), .ZN(n10951) );
  INV_X1 U13062 ( .A(n12345), .ZN(n10522) );
  NAND2_X1 U13063 ( .A1(n10522), .A2(n10475), .ZN(n10587) );
  OAI211_X1 U13064 ( .C1(n10522), .C2(n10475), .A(n14888), .B(n10587), .ZN(
        n10949) );
  OAI211_X1 U13065 ( .C1(n10958), .C2(n15229), .A(n10951), .B(n10949), .ZN(
        n10476) );
  AOI21_X1 U13066 ( .B1(n14939), .B2(n10948), .A(n10476), .ZN(n10480) );
  OAI22_X1 U13067 ( .A1(n15011), .A2(n10522), .B1(n15259), .B2(n10411), .ZN(
        n10477) );
  INV_X1 U13068 ( .A(n10477), .ZN(n10478) );
  OAI21_X1 U13069 ( .B1(n10480), .B2(n15257), .A(n10478), .ZN(P1_U3480) );
  AOI22_X1 U13070 ( .A1(n14900), .A2(n12345), .B1(n15265), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n10479) );
  OAI21_X1 U13071 ( .B1(n10480), .B2(n15265), .A(n10479), .ZN(P1_U3535) );
  NAND2_X1 U13072 ( .A1(n10482), .A2(n10481), .ZN(n10485) );
  NAND2_X1 U13073 ( .A1(n13743), .A2(n10483), .ZN(n10484) );
  AND2_X1 U13074 ( .A1(n10485), .A2(n10484), .ZN(n10486) );
  MUX2_X1 U13075 ( .A(n10526), .B(P3_REG2_REG_0__SCAN_IN), .S(n15489), .Z(
        n10492) );
  INV_X1 U13076 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10490) );
  OAI22_X1 U13077 ( .A1(n13587), .A2(n10524), .B1(n15525), .B2(n10490), .ZN(
        n10491) );
  OR2_X1 U13078 ( .A1(n10492), .A2(n10491), .ZN(P3_U3233) );
  NAND2_X1 U13079 ( .A1(n10494), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10493) );
  MUX2_X1 U13080 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10493), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n10495) );
  NAND2_X1 U13081 ( .A1(n10495), .A2(n11021), .ZN(n11393) );
  INV_X1 U13082 ( .A(n11814), .ZN(n10528) );
  OAI222_X1 U13083 ( .A1(P1_U3086), .A2(n11393), .B1(n15030), .B2(n10528), 
        .C1(n10496), .C2(n15024), .ZN(P1_U3339) );
  NAND2_X1 U13084 ( .A1(n14429), .A2(n12708), .ZN(n10501) );
  NAND2_X1 U13085 ( .A1(n10103), .A2(n14471), .ZN(n10500) );
  NAND2_X1 U13086 ( .A1(n10501), .A2(n10500), .ZN(n10502) );
  XNOR2_X1 U13087 ( .A(n10502), .B(n11728), .ZN(n10506) );
  NAND2_X1 U13088 ( .A1(n14429), .A2(n10103), .ZN(n10505) );
  NAND2_X1 U13089 ( .A1(n12709), .A2(n14471), .ZN(n10504) );
  NAND2_X1 U13090 ( .A1(n10505), .A2(n10504), .ZN(n10507) );
  XNOR2_X1 U13091 ( .A(n10506), .B(n10507), .ZN(n14427) );
  NAND2_X1 U13092 ( .A1(n14428), .A2(n14427), .ZN(n14426) );
  INV_X1 U13093 ( .A(n10506), .ZN(n10508) );
  NAND2_X1 U13094 ( .A1(n10508), .A2(n10507), .ZN(n10509) );
  NAND2_X1 U13095 ( .A1(n12345), .A2(n12708), .ZN(n10511) );
  NAND2_X1 U13096 ( .A1(n10103), .A2(n14470), .ZN(n10510) );
  NAND2_X1 U13097 ( .A1(n10511), .A2(n10510), .ZN(n10512) );
  XNOR2_X1 U13098 ( .A(n10512), .B(n12710), .ZN(n10758) );
  NOR2_X1 U13099 ( .A1(n6812), .A2(n10513), .ZN(n10514) );
  AOI21_X1 U13100 ( .B1(n12345), .B2(n10103), .A(n10514), .ZN(n10756) );
  XNOR2_X1 U13101 ( .A(n10758), .B(n10756), .ZN(n10515) );
  OAI211_X1 U13102 ( .C1(n10516), .C2(n10515), .A(n10760), .B(n14425), .ZN(
        n10521) );
  INV_X1 U13103 ( .A(n14410), .ZN(n14362) );
  AND2_X1 U13104 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14545) );
  AOI21_X1 U13105 ( .B1(n14362), .B2(n10517), .A(n14545), .ZN(n10518) );
  OAI21_X1 U13106 ( .B1(n14441), .B2(n10953), .A(n10518), .ZN(n10519) );
  INV_X1 U13107 ( .A(n10519), .ZN(n10520) );
  OAI211_X1 U13108 ( .C1(n10522), .C2(n14450), .A(n10521), .B(n10520), .ZN(
        P1_U3213) );
  INV_X1 U13109 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10523) );
  OAI22_X1 U13110 ( .A1(n13741), .A2(n10524), .B1(n15582), .B2(n10523), .ZN(
        n10525) );
  AOI21_X1 U13111 ( .B1(n10526), .B2(n15582), .A(n10525), .ZN(n10527) );
  INV_X1 U13112 ( .A(n10527), .ZN(P3_U3390) );
  OAI222_X1 U13113 ( .A1(n14312), .A2(n10529), .B1(n11776), .B2(P2_U3088), 
        .C1(n10596), .C2(n10528), .ZN(P2_U3311) );
  MUX2_X1 U13114 ( .A(n15496), .B(n12068), .S(n12734), .Z(n10530) );
  XNOR2_X1 U13115 ( .A(n7799), .B(n6604), .ZN(n10623) );
  XNOR2_X1 U13116 ( .A(n10623), .B(n7798), .ZN(n10621) );
  XNOR2_X1 U13117 ( .A(n10622), .B(n10621), .ZN(n10537) );
  NAND2_X1 U13118 ( .A1(n10532), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13119 ( .A1(n12896), .A2(n12878), .B1(n12869), .B2(n10533), .ZN(
        n10534) );
  OAI211_X1 U13120 ( .C1(n15493), .C2(n12880), .A(n10535), .B(n10534), .ZN(
        n10536) );
  AOI21_X1 U13121 ( .B1(n10537), .B2(n12874), .A(n10536), .ZN(n10538) );
  INV_X1 U13122 ( .A(n10538), .ZN(P3_U3177) );
  NAND2_X1 U13123 ( .A1(n11021), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10539) );
  XNOR2_X1 U13124 ( .A(n10539), .B(P1_IR_REG_17__SCAN_IN), .ZN(n11820) );
  INV_X1 U13125 ( .A(n11820), .ZN(n11527) );
  INV_X1 U13126 ( .A(n11819), .ZN(n10595) );
  OAI222_X1 U13127 ( .A1(P1_U3086), .A2(n11527), .B1(n15030), .B2(n10595), 
        .C1(n10540), .C2(n15024), .ZN(P1_U3338) );
  OAI21_X1 U13128 ( .B1(n10542), .B2(n10546), .A(n10541), .ZN(n10659) );
  OAI211_X1 U13129 ( .C1(n10562), .C2(n10543), .A(n10037), .B(n10609), .ZN(
        n10657) );
  INV_X1 U13130 ( .A(n10657), .ZN(n10553) );
  OAI22_X1 U13131 ( .A1(n10645), .A2(n15098), .B1(n10544), .B2(n15096), .ZN(
        n10559) );
  NAND3_X1 U13132 ( .A1(n10547), .A2(n10546), .A3(n10545), .ZN(n10548) );
  AOI21_X1 U13133 ( .B1(n10549), .B2(n10548), .A(n15125), .ZN(n10550) );
  AOI211_X1 U13134 ( .C1(n10551), .C2(n10659), .A(n10559), .B(n10550), .ZN(
        n10652) );
  INV_X1 U13135 ( .A(n10652), .ZN(n10552) );
  AOI211_X1 U13136 ( .C1(n15390), .C2(n10659), .A(n10553), .B(n10552), .ZN(
        n10558) );
  INV_X1 U13137 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10554) );
  OAI22_X1 U13138 ( .A1(n14287), .A2(n10562), .B1(n15393), .B2(n10554), .ZN(
        n10555) );
  INV_X1 U13139 ( .A(n10555), .ZN(n10556) );
  OAI21_X1 U13140 ( .B1(n10558), .B2(n15391), .A(n10556), .ZN(P2_U3448) );
  AOI22_X1 U13141 ( .A1(n14248), .A2(n10655), .B1(n6794), .B2(
        P2_REG1_REG_6__SCAN_IN), .ZN(n10557) );
  OAI21_X1 U13142 ( .B1(n10558), .B2(n6794), .A(n10557), .ZN(P2_U3505) );
  NAND2_X1 U13143 ( .A1(n15106), .A2(n10559), .ZN(n10561) );
  OAI211_X1 U13144 ( .C1(n13888), .C2(n10562), .A(n10561), .B(n10560), .ZN(
        n10567) );
  INV_X1 U13145 ( .A(n10386), .ZN(n10564) );
  AOI211_X1 U13146 ( .C1(n10565), .C2(n10563), .A(n13872), .B(n10564), .ZN(
        n10566) );
  AOI211_X1 U13147 ( .C1(n13855), .C2(n10654), .A(n10567), .B(n10566), .ZN(
        n10568) );
  INV_X1 U13148 ( .A(n10568), .ZN(P2_U3211) );
  OR2_X1 U13149 ( .A1(n10570), .A2(n11448), .ZN(n10573) );
  AOI22_X1 U13150 ( .A1(n11845), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11844), 
        .B2(n10571), .ZN(n10572) );
  INV_X1 U13151 ( .A(n14469), .ZN(n10754) );
  XNOR2_X1 U13152 ( .A(n12351), .B(n10754), .ZN(n12498) );
  XNOR2_X1 U13153 ( .A(n10723), .B(n12498), .ZN(n10976) );
  OR2_X1 U13154 ( .A1(n12345), .A2(n14470), .ZN(n10574) );
  OAI21_X1 U13155 ( .B1(n10576), .B2(n12498), .A(n10733), .ZN(n10577) );
  INV_X1 U13156 ( .A(n10577), .ZN(n10979) );
  NAND2_X1 U13157 ( .A1(n14470), .A2(n14791), .ZN(n10586) );
  NAND2_X1 U13158 ( .A1(n11985), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10584) );
  INV_X1 U13159 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10578) );
  OR2_X1 U13160 ( .A1(n11944), .A2(n10578), .ZN(n10583) );
  NAND2_X1 U13161 ( .A1(n10579), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10736) );
  OR2_X1 U13162 ( .A1(n10579), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10580) );
  NAND2_X1 U13163 ( .A1(n10736), .A2(n10580), .ZN(n11053) );
  OR2_X1 U13164 ( .A1(n11986), .A2(n11053), .ZN(n10582) );
  OR2_X1 U13165 ( .A1(n12454), .A2(n13354), .ZN(n10581) );
  NAND4_X1 U13166 ( .A1(n10584), .A2(n10583), .A3(n10582), .A4(n10581), .ZN(
        n14468) );
  NAND2_X1 U13167 ( .A1(n14468), .A2(n14850), .ZN(n10585) );
  NAND2_X1 U13168 ( .A1(n10586), .A2(n10585), .ZN(n10971) );
  INV_X1 U13169 ( .A(n10971), .ZN(n10589) );
  AOI21_X1 U13170 ( .B1(n12351), .B2(n10587), .A(n14828), .ZN(n10588) );
  NAND2_X1 U13171 ( .A1(n10588), .A2(n10744), .ZN(n10973) );
  OAI211_X1 U13172 ( .C1(n10979), .C2(n15229), .A(n10589), .B(n10973), .ZN(
        n10590) );
  AOI21_X1 U13173 ( .B1(n10976), .B2(n14939), .A(n10590), .ZN(n10594) );
  AOI22_X1 U13174 ( .A1(n14900), .A2(n12351), .B1(n15265), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n10591) );
  OAI21_X1 U13175 ( .B1(n10594), .B2(n15265), .A(n10591), .ZN(P1_U3536) );
  INV_X1 U13176 ( .A(n15011), .ZN(n14988) );
  NOR2_X1 U13177 ( .A1(n15259), .A2(n10464), .ZN(n10592) );
  AOI21_X1 U13178 ( .B1(n14988), .B2(n12351), .A(n10592), .ZN(n10593) );
  OAI21_X1 U13179 ( .B1(n10594), .B2(n15257), .A(n10593), .ZN(P1_U3483) );
  INV_X1 U13180 ( .A(n11784), .ZN(n15310) );
  OAI222_X1 U13181 ( .A1(n14312), .A2(n13533), .B1(n15310), .B2(P2_U3088), 
        .C1(n10596), .C2(n10595), .ZN(P2_U3310) );
  NAND2_X1 U13182 ( .A1(n6581), .A2(n10597), .ZN(n10599) );
  NAND2_X1 U13183 ( .A1(n15329), .A2(n12004), .ZN(n10598) );
  OAI211_X1 U13184 ( .C1(n12003), .C2(n15334), .A(n10599), .B(n10598), .ZN(
        n10602) );
  MUX2_X1 U13185 ( .A(n10600), .B(P2_REG2_REG_5__SCAN_IN), .S(n8990), .Z(
        n10601) );
  AOI211_X1 U13186 ( .C1(n14168), .C2(n10603), .A(n10602), .B(n10601), .ZN(
        n10604) );
  INV_X1 U13187 ( .A(n10604), .ZN(P2_U3260) );
  OAI21_X1 U13188 ( .B1(n10607), .B2(n10610), .A(n10606), .ZN(n15336) );
  INV_X1 U13189 ( .A(n10608), .ZN(n10702) );
  AOI211_X1 U13190 ( .C1(n15326), .C2(n10609), .A(n13997), .B(n10702), .ZN(
        n15328) );
  XOR2_X1 U13191 ( .A(n10611), .B(n10610), .Z(n10613) );
  AOI21_X1 U13192 ( .B1(n10613), .B2(n6580), .A(n10612), .ZN(n15339) );
  INV_X1 U13193 ( .A(n15339), .ZN(n10614) );
  AOI211_X1 U13194 ( .C1(n15372), .C2(n15336), .A(n15328), .B(n10614), .ZN(
        n10619) );
  INV_X1 U13195 ( .A(n14287), .ZN(n14294) );
  INV_X1 U13196 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10615) );
  NOR2_X1 U13197 ( .A1(n15393), .A2(n10615), .ZN(n10616) );
  AOI21_X1 U13198 ( .B1(n14294), .B2(n15326), .A(n10616), .ZN(n10617) );
  OAI21_X1 U13199 ( .B1(n10619), .B2(n15391), .A(n10617), .ZN(P2_U3451) );
  AOI22_X1 U13200 ( .A1(n14248), .A2(n15326), .B1(n6794), .B2(
        P2_REG1_REG_7__SCAN_IN), .ZN(n10618) );
  OAI21_X1 U13201 ( .B1(n10619), .B2(n6794), .A(n10618), .ZN(P2_U3506) );
  NAND2_X1 U13202 ( .A1(n10622), .A2(n10621), .ZN(n10627) );
  NAND2_X1 U13203 ( .A1(n10629), .A2(n10623), .ZN(n10626) );
  NAND2_X1 U13204 ( .A1(n10627), .A2(n10626), .ZN(n10624) );
  XNOR2_X1 U13205 ( .A(n15483), .B(n12734), .ZN(n10787) );
  AOI21_X1 U13206 ( .B1(n10624), .B2(n10625), .A(n12872), .ZN(n10628) );
  NAND2_X1 U13207 ( .A1(n10628), .A2(n10789), .ZN(n10633) );
  INV_X1 U13208 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15484) );
  NOR2_X1 U13209 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15484), .ZN(n15416) );
  OAI22_X1 U13210 ( .A1(n10912), .A2(n12867), .B1(n10629), .B2(n12880), .ZN(
        n10630) );
  AOI211_X1 U13211 ( .C1(n12869), .C2(n10631), .A(n15416), .B(n10630), .ZN(
        n10632) );
  OAI211_X1 U13212 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11604), .A(n10633), .B(
        n10632), .ZN(P3_U3158) );
  XNOR2_X1 U13213 ( .A(n10704), .B(n13792), .ZN(n10634) );
  NAND2_X1 U13214 ( .A1(n13909), .A2(n13997), .ZN(n10635) );
  NAND2_X1 U13215 ( .A1(n10634), .A2(n10635), .ZN(n10872) );
  INV_X1 U13216 ( .A(n10634), .ZN(n10637) );
  INV_X1 U13217 ( .A(n10635), .ZN(n10636) );
  NAND2_X1 U13218 ( .A1(n10637), .A2(n10636), .ZN(n10874) );
  NAND2_X1 U13219 ( .A1(n10872), .A2(n10874), .ZN(n10642) );
  INV_X1 U13220 ( .A(n10638), .ZN(n10639) );
  XOR2_X1 U13221 ( .A(n10642), .B(n10873), .Z(n10649) );
  INV_X1 U13222 ( .A(n10703), .ZN(n10644) );
  OAI21_X1 U13223 ( .B1(n15111), .B2(n10644), .A(n10643), .ZN(n10647) );
  OAI22_X1 U13224 ( .A1(n13883), .A2(n10902), .B1(n13881), .B2(n10645), .ZN(
        n10646) );
  AOI211_X1 U13225 ( .C1(n10704), .C2(n15107), .A(n10647), .B(n10646), .ZN(
        n10648) );
  OAI21_X1 U13226 ( .B1(n10649), .B2(n13872), .A(n10648), .ZN(P2_U3193) );
  INV_X1 U13227 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n10651) );
  NAND2_X1 U13228 ( .A1(n13133), .A2(P3_U3897), .ZN(n10650) );
  OAI21_X1 U13229 ( .B1(P3_U3897), .B2(n10651), .A(n10650), .ZN(P3_U3517) );
  MUX2_X1 U13230 ( .A(n10653), .B(n10652), .S(n14163), .Z(n10661) );
  AOI22_X1 U13231 ( .A1(n15132), .A2(n10655), .B1(n15329), .B2(n10654), .ZN(
        n10656) );
  OAI21_X1 U13232 ( .B1(n14152), .B2(n10657), .A(n10656), .ZN(n10658) );
  AOI21_X1 U13233 ( .B1(n10659), .B2(n14168), .A(n10658), .ZN(n10660) );
  NAND2_X1 U13234 ( .A1(n10661), .A2(n10660), .ZN(P2_U3259) );
  OAI21_X1 U13235 ( .B1(n10664), .B2(n10663), .A(n10662), .ZN(n15364) );
  OAI21_X1 U13236 ( .B1(n10667), .B2(n10666), .A(n10665), .ZN(n10668) );
  NAND2_X1 U13237 ( .A1(n10668), .A2(n6580), .ZN(n10670) );
  AOI22_X1 U13238 ( .A1(n14025), .A2(n13915), .B1(n13913), .B2(n14027), .ZN(
        n10669) );
  AND2_X1 U13239 ( .A1(n10670), .A2(n10669), .ZN(n15361) );
  OAI21_X1 U13240 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n14147), .A(n15361), .ZN(
        n10671) );
  MUX2_X1 U13241 ( .A(n10671), .B(P2_REG2_REG_3__SCAN_IN), .S(n8990), .Z(
        n10674) );
  OAI211_X1 U13242 ( .C1(n10672), .C2(n15360), .A(n10037), .B(n10683), .ZN(
        n15359) );
  OAI22_X1 U13243 ( .A1(n14152), .A2(n15359), .B1(n15360), .B2(n15334), .ZN(
        n10673) );
  AOI211_X1 U13244 ( .C1(n15337), .C2(n15364), .A(n10674), .B(n10673), .ZN(
        n10675) );
  INV_X1 U13245 ( .A(n10675), .ZN(P2_U3262) );
  OAI21_X1 U13246 ( .B1(n10678), .B2(n10677), .A(n10676), .ZN(n10679) );
  AOI222_X1 U13247 ( .A1(n6580), .A2(n10679), .B1(n13912), .B2(n14027), .C1(
        n13914), .C2(n14025), .ZN(n15368) );
  MUX2_X1 U13248 ( .A(n9472), .B(n15368), .S(n14163), .Z(n10691) );
  OAI21_X1 U13249 ( .B1(n10682), .B2(n10681), .A(n10680), .ZN(n15371) );
  AOI21_X1 U13250 ( .B1(n10683), .B2(n10687), .A(n13997), .ZN(n10685) );
  NAND2_X1 U13251 ( .A1(n10685), .A2(n10684), .ZN(n15366) );
  AOI22_X1 U13252 ( .A1(n15132), .A2(n10687), .B1(n15329), .B2(n10686), .ZN(
        n10688) );
  OAI21_X1 U13253 ( .B1(n14152), .B2(n15366), .A(n10688), .ZN(n10689) );
  AOI21_X1 U13254 ( .B1(n15337), .B2(n15371), .A(n10689), .ZN(n10690) );
  NAND2_X1 U13255 ( .A1(n10691), .A2(n10690), .ZN(P2_U3261) );
  NAND2_X1 U13256 ( .A1(n10692), .A2(n10695), .ZN(n10693) );
  NAND2_X1 U13257 ( .A1(n10694), .A2(n10693), .ZN(n10700) );
  AOI22_X1 U13258 ( .A1(n14025), .A2(n13910), .B1(n13908), .B2(n14027), .ZN(
        n10699) );
  XNOR2_X1 U13259 ( .A(n10696), .B(n10695), .ZN(n10697) );
  NAND2_X1 U13260 ( .A1(n10697), .A2(n6580), .ZN(n10698) );
  OAI211_X1 U13261 ( .C1(n10700), .C2(n9899), .A(n10699), .B(n10698), .ZN(
        n15375) );
  INV_X1 U13262 ( .A(n15375), .ZN(n10709) );
  INV_X1 U13263 ( .A(n10700), .ZN(n15377) );
  INV_X1 U13264 ( .A(n10701), .ZN(n10776) );
  OAI211_X1 U13265 ( .C1(n7500), .C2(n10702), .A(n10776), .B(n10037), .ZN(
        n15374) );
  AOI22_X1 U13266 ( .A1(n15331), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10703), 
        .B2(n15329), .ZN(n10706) );
  NAND2_X1 U13267 ( .A1(n15132), .A2(n10704), .ZN(n10705) );
  OAI211_X1 U13268 ( .C1(n15374), .C2(n14152), .A(n10706), .B(n10705), .ZN(
        n10707) );
  AOI21_X1 U13269 ( .B1(n15377), .B2(n14168), .A(n10707), .ZN(n10708) );
  OAI21_X1 U13270 ( .B1(n10709), .B2(n15331), .A(n10708), .ZN(P2_U3257) );
  XNOR2_X1 U13271 ( .A(n10710), .B(n12204), .ZN(n15548) );
  NAND2_X1 U13272 ( .A1(n15548), .A2(n15502), .ZN(n10718) );
  NAND2_X1 U13273 ( .A1(n15476), .A2(n10711), .ZN(n10712) );
  XNOR2_X1 U13274 ( .A(n10712), .B(n12204), .ZN(n10716) );
  NAND2_X1 U13275 ( .A1(n12896), .A2(n15515), .ZN(n10714) );
  NAND2_X1 U13276 ( .A1(n15459), .A2(n15517), .ZN(n10713) );
  NAND2_X1 U13277 ( .A1(n10714), .A2(n10713), .ZN(n10715) );
  AOI21_X1 U13278 ( .B1(n10716), .B2(n15513), .A(n10715), .ZN(n10717) );
  NOR2_X1 U13279 ( .A1(n15504), .A2(n12060), .ZN(n15505) );
  NOR2_X1 U13280 ( .A1(n10786), .A2(n15559), .ZN(n15547) );
  AOI22_X1 U13281 ( .A1(n15547), .A2(n15485), .B1(n15508), .B2(n10785), .ZN(
        n10719) );
  OAI21_X1 U13282 ( .B1(n10297), .B2(n15530), .A(n10719), .ZN(n10720) );
  AOI21_X1 U13283 ( .B1(n15548), .B2(n15444), .A(n10720), .ZN(n10721) );
  OAI21_X1 U13284 ( .B1(n15550), .B2(n15489), .A(n10721), .ZN(P3_U3229) );
  INV_X1 U13285 ( .A(n12498), .ZN(n10722) );
  OR2_X1 U13286 ( .A1(n12351), .A2(n10754), .ZN(n10724) );
  NAND2_X1 U13287 ( .A1(n10725), .A2(n10724), .ZN(n10729) );
  INV_X1 U13288 ( .A(n10729), .ZN(n10731) );
  OR2_X1 U13289 ( .A1(n10726), .A2(n11448), .ZN(n10728) );
  AOI22_X1 U13290 ( .A1(n11845), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11844), 
        .B2(n14572), .ZN(n10727) );
  INV_X1 U13291 ( .A(n14468), .ZN(n11201) );
  INV_X1 U13292 ( .A(n12499), .ZN(n10730) );
  OR2_X2 U13293 ( .A1(n10729), .A2(n12499), .ZN(n11106) );
  OAI21_X1 U13294 ( .B1(n10731), .B2(n10730), .A(n11106), .ZN(n10959) );
  OR2_X1 U13295 ( .A1(n12351), .A2(n14469), .ZN(n10732) );
  OAI21_X1 U13296 ( .B1(n10734), .B2(n12499), .A(n11115), .ZN(n10735) );
  INV_X1 U13297 ( .A(n10735), .ZN(n10968) );
  NAND2_X1 U13298 ( .A1(n12450), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10742) );
  OR2_X1 U13299 ( .A1(n12289), .A2(n9625), .ZN(n10741) );
  NAND2_X1 U13300 ( .A1(n10736), .A2(n13417), .ZN(n10737) );
  NAND2_X1 U13301 ( .A1(n11121), .A2(n10737), .ZN(n11204) );
  OR2_X1 U13302 ( .A1(n11986), .A2(n11204), .ZN(n10740) );
  OR2_X1 U13303 ( .A1(n12454), .A2(n10738), .ZN(n10739) );
  NAND4_X1 U13304 ( .A1(n10742), .A2(n10741), .A3(n10740), .A4(n10739), .ZN(
        n14467) );
  AOI22_X1 U13305 ( .A1(n14791), .A2(n14469), .B1(n14467), .B2(n14850), .ZN(
        n10961) );
  INV_X1 U13306 ( .A(n12356), .ZN(n11058) );
  AOI21_X1 U13307 ( .B1(n12356), .B2(n10744), .A(n14828), .ZN(n10745) );
  NAND2_X1 U13308 ( .A1(n11157), .A2(n10745), .ZN(n10963) );
  OAI211_X1 U13309 ( .C1(n10968), .C2(n15229), .A(n10961), .B(n10963), .ZN(
        n10746) );
  AOI21_X1 U13310 ( .B1(n14939), .B2(n10959), .A(n10746), .ZN(n10750) );
  AOI22_X1 U13311 ( .A1(n12356), .A2(n14900), .B1(n15265), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n10747) );
  OAI21_X1 U13312 ( .B1(n10750), .B2(n15265), .A(n10747), .ZN(P1_U3537) );
  OAI22_X1 U13313 ( .A1(n11058), .A2(n15011), .B1(n15259), .B2(n10578), .ZN(
        n10748) );
  INV_X1 U13314 ( .A(n10748), .ZN(n10749) );
  OAI21_X1 U13315 ( .B1(n10750), .B2(n15257), .A(n10749), .ZN(P1_U3486) );
  NAND2_X1 U13316 ( .A1(n12351), .A2(n12708), .ZN(n10752) );
  NAND2_X1 U13317 ( .A1(n10103), .A2(n14469), .ZN(n10751) );
  NAND2_X1 U13318 ( .A1(n10752), .A2(n10751), .ZN(n10753) );
  XNOR2_X1 U13319 ( .A(n10753), .B(n11728), .ZN(n11046) );
  NOR2_X1 U13320 ( .A1(n6812), .A2(n10754), .ZN(n10755) );
  AOI21_X1 U13321 ( .B1(n12351), .B2(n10103), .A(n10755), .ZN(n11045) );
  XNOR2_X1 U13322 ( .A(n11046), .B(n11045), .ZN(n10764) );
  INV_X1 U13323 ( .A(n10756), .ZN(n10757) );
  NAND2_X1 U13324 ( .A1(n10758), .A2(n10757), .ZN(n10759) );
  INV_X1 U13325 ( .A(n10764), .ZN(n10761) );
  INV_X1 U13326 ( .A(n11048), .ZN(n10762) );
  AOI21_X1 U13327 ( .B1(n10764), .B2(n10763), .A(n10762), .ZN(n10768) );
  AOI22_X1 U13328 ( .A1(n14362), .A2(n10971), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10765) );
  OAI21_X1 U13329 ( .B1(n14441), .B2(n10969), .A(n10765), .ZN(n10766) );
  AOI21_X1 U13330 ( .B1(n12351), .B2(n9832), .A(n10766), .ZN(n10767) );
  OAI21_X1 U13331 ( .B1(n10768), .B2(n14456), .A(n10767), .ZN(P1_U3221) );
  XNOR2_X1 U13332 ( .A(n10769), .B(n10770), .ZN(n10886) );
  INV_X1 U13333 ( .A(n14168), .ZN(n10781) );
  XNOR2_X1 U13334 ( .A(n10771), .B(n10770), .ZN(n10773) );
  OAI22_X1 U13335 ( .A1(n10881), .A2(n15096), .B1(n11226), .B2(n15098), .ZN(
        n10772) );
  AOI21_X1 U13336 ( .B1(n10773), .B2(n6580), .A(n10772), .ZN(n10774) );
  OAI21_X1 U13337 ( .B1(n10886), .B2(n9899), .A(n10774), .ZN(n10887) );
  NAND2_X1 U13338 ( .A1(n10887), .A2(n14163), .ZN(n10780) );
  INV_X1 U13339 ( .A(n10775), .ZN(n10810) );
  AOI211_X1 U13340 ( .C1(n10890), .C2(n10776), .A(n13997), .B(n10810), .ZN(
        n10888) );
  AOI22_X1 U13341 ( .A1(n15331), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10879), 
        .B2(n15329), .ZN(n10777) );
  OAI21_X1 U13342 ( .B1(n10893), .B2(n15334), .A(n10777), .ZN(n10778) );
  AOI21_X1 U13343 ( .B1(n10888), .B2(n6581), .A(n10778), .ZN(n10779) );
  OAI211_X1 U13344 ( .C1(n10886), .C2(n10781), .A(n10780), .B(n10779), .ZN(
        P2_U3256) );
  INV_X1 U13345 ( .A(n10785), .ZN(n10798) );
  XNOR2_X1 U13346 ( .A(n10786), .B(n12771), .ZN(n10909) );
  XNOR2_X1 U13347 ( .A(n10909), .B(n15474), .ZN(n10791) );
  NAND2_X1 U13348 ( .A1(n10787), .A2(n12896), .ZN(n10788) );
  AND2_X2 U13349 ( .A1(n10789), .A2(n10788), .ZN(n10790) );
  OAI21_X1 U13350 ( .B1(n10791), .B2(n10790), .A(n10911), .ZN(n10792) );
  NAND2_X1 U13351 ( .A1(n10792), .A2(n12874), .ZN(n10797) );
  OAI22_X1 U13352 ( .A1(n11035), .A2(n12867), .B1(n15495), .B2(n12880), .ZN(
        n10793) );
  AOI211_X1 U13353 ( .C1(n12869), .C2(n10795), .A(n10794), .B(n10793), .ZN(
        n10796) );
  OAI211_X1 U13354 ( .C1(n10798), .C2(n11604), .A(n10797), .B(n10796), .ZN(
        P3_U3170) );
  INV_X1 U13355 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n10801) );
  NAND2_X1 U13356 ( .A1(n10799), .A2(P3_U3897), .ZN(n10800) );
  OAI21_X1 U13357 ( .B1(P3_U3897), .B2(n10801), .A(n10800), .ZN(P3_U3519) );
  XNOR2_X1 U13358 ( .A(n10802), .B(n10803), .ZN(n10808) );
  XNOR2_X1 U13359 ( .A(n10804), .B(n10803), .ZN(n10806) );
  OAI22_X1 U13360 ( .A1(n10902), .A2(n15096), .B1(n10903), .B2(n15098), .ZN(
        n10805) );
  AOI21_X1 U13361 ( .B1(n10806), .B2(n6580), .A(n10805), .ZN(n10807) );
  OAI21_X1 U13362 ( .B1(n10808), .B2(n9899), .A(n10807), .ZN(n15381) );
  INV_X1 U13363 ( .A(n15381), .ZN(n10815) );
  INV_X1 U13364 ( .A(n10808), .ZN(n15383) );
  INV_X1 U13365 ( .A(n10906), .ZN(n15380) );
  OAI211_X1 U13366 ( .C1(n15380), .C2(n10810), .A(n10037), .B(n10987), .ZN(
        n15379) );
  AOI22_X1 U13367 ( .A1(n8990), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10899), 
        .B2(n15329), .ZN(n10812) );
  NAND2_X1 U13368 ( .A1(n10906), .A2(n15132), .ZN(n10811) );
  OAI211_X1 U13369 ( .C1(n15379), .C2(n14152), .A(n10812), .B(n10811), .ZN(
        n10813) );
  AOI21_X1 U13370 ( .B1(n15383), .B2(n14168), .A(n10813), .ZN(n10814) );
  OAI21_X1 U13371 ( .B1(n10815), .B2(n15331), .A(n10814), .ZN(P2_U3255) );
  INV_X1 U13372 ( .A(n10816), .ZN(n10828) );
  NOR2_X1 U13373 ( .A1(n10817), .A2(n12528), .ZN(n10819) );
  NAND2_X1 U13374 ( .A1(n10819), .A2(n10818), .ZN(n14607) );
  OR2_X1 U13375 ( .A1(n12300), .A2(n11695), .ZN(n12294) );
  NOR2_X1 U13376 ( .A1(n14855), .A2(n12294), .ZN(n14846) );
  INV_X1 U13377 ( .A(n14846), .ZN(n14798) );
  INV_X1 U13378 ( .A(n10820), .ZN(n10821) );
  MUX2_X1 U13379 ( .A(n9622), .B(n10821), .S(n14840), .Z(n10827) );
  INV_X1 U13380 ( .A(n10822), .ZN(n10823) );
  OAI22_X1 U13381 ( .A1(n14831), .A2(n12341), .B1(n14852), .B2(n14431), .ZN(
        n10824) );
  AOI21_X1 U13382 ( .B1(n14835), .B2(n10825), .A(n10824), .ZN(n10826) );
  OAI211_X1 U13383 ( .C1(n10828), .C2(n14798), .A(n10827), .B(n10826), .ZN(
        P1_U3287) );
  INV_X1 U13384 ( .A(n10829), .ZN(n10838) );
  INV_X1 U13385 ( .A(n10831), .ZN(n10832) );
  MUX2_X1 U13386 ( .A(n9570), .B(n10832), .S(n14840), .Z(n10837) );
  OAI22_X1 U13387 ( .A1(n14831), .A2(n12325), .B1(n14852), .B2(n10833), .ZN(
        n10834) );
  AOI21_X1 U13388 ( .B1(n14835), .B2(n10835), .A(n10834), .ZN(n10836) );
  OAI211_X1 U13389 ( .C1(n10838), .C2(n14838), .A(n10837), .B(n10836), .ZN(
        P1_U3289) );
  OR2_X1 U13390 ( .A1(n10839), .A2(n12491), .ZN(n10840) );
  NAND2_X1 U13391 ( .A1(n10841), .A2(n10840), .ZN(n15238) );
  INV_X1 U13392 ( .A(n15238), .ZN(n10855) );
  OAI21_X1 U13393 ( .B1(n10843), .B2(n12317), .A(n10842), .ZN(n10845) );
  OAI22_X1 U13394 ( .A1(n12315), .A2(n14824), .B1(n12326), .B2(n14826), .ZN(
        n10844) );
  AOI21_X1 U13395 ( .B1(n10845), .B2(n14939), .A(n10844), .ZN(n10847) );
  NAND2_X1 U13396 ( .A1(n15238), .A2(n14629), .ZN(n10846) );
  AND2_X1 U13397 ( .A1(n10847), .A2(n10846), .ZN(n15240) );
  MUX2_X1 U13398 ( .A(n15240), .B(n10848), .S(n14855), .Z(n10854) );
  INV_X1 U13399 ( .A(n15236), .ZN(n14332) );
  OAI21_X1 U13400 ( .B1(n10849), .B2(n15236), .A(n14888), .ZN(n10851) );
  OR2_X1 U13401 ( .A1(n10851), .A2(n10850), .ZN(n15235) );
  OAI22_X1 U13402 ( .A1(n14783), .A2(n15235), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14852), .ZN(n10852) );
  AOI21_X1 U13403 ( .B1(n14858), .B2(n14332), .A(n10852), .ZN(n10853) );
  OAI211_X1 U13404 ( .C1(n14798), .C2(n10855), .A(n10854), .B(n10853), .ZN(
        P1_U3290) );
  MUX2_X1 U13405 ( .A(n10857), .B(n10856), .S(n14840), .Z(n10862) );
  OAI22_X1 U13406 ( .A1(n14783), .A2(n10859), .B1(n10858), .B2(n14852), .ZN(
        n10860) );
  AOI21_X1 U13407 ( .B1(n14858), .B2(n12312), .A(n10860), .ZN(n10861) );
  OAI211_X1 U13408 ( .C1(n14798), .C2(n10863), .A(n10862), .B(n10861), .ZN(
        P1_U3291) );
  INV_X1 U13409 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n10866) );
  INV_X1 U13410 ( .A(n13094), .ZN(n10864) );
  NAND2_X1 U13411 ( .A1(n10864), .A2(P3_U3897), .ZN(n10865) );
  OAI21_X1 U13412 ( .B1(P3_U3897), .B2(n10866), .A(n10865), .ZN(P3_U3520) );
  XNOR2_X1 U13413 ( .A(n10890), .B(n13792), .ZN(n10867) );
  NAND2_X1 U13414 ( .A1(n13908), .A2(n13997), .ZN(n10868) );
  NAND2_X1 U13415 ( .A1(n10867), .A2(n10868), .ZN(n10897) );
  INV_X1 U13416 ( .A(n10867), .ZN(n10870) );
  INV_X1 U13417 ( .A(n10868), .ZN(n10869) );
  NAND2_X1 U13418 ( .A1(n10870), .A2(n10869), .ZN(n10871) );
  NAND2_X1 U13419 ( .A1(n10897), .A2(n10871), .ZN(n10878) );
  INV_X1 U13420 ( .A(n10898), .ZN(n10876) );
  AOI21_X1 U13421 ( .B1(n10878), .B2(n10877), .A(n10876), .ZN(n10885) );
  INV_X1 U13422 ( .A(n10879), .ZN(n10880) );
  NAND2_X1 U13423 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n13932) );
  OAI21_X1 U13424 ( .B1(n15111), .B2(n10880), .A(n13932), .ZN(n10883) );
  OAI22_X1 U13425 ( .A1(n13883), .A2(n11226), .B1(n13881), .B2(n10881), .ZN(
        n10882) );
  AOI211_X1 U13426 ( .C1(n10890), .C2(n15107), .A(n10883), .B(n10882), .ZN(
        n10884) );
  OAI21_X1 U13427 ( .B1(n10885), .B2(n13872), .A(n10884), .ZN(P2_U3203) );
  INV_X1 U13428 ( .A(n10886), .ZN(n10889) );
  AOI211_X1 U13429 ( .C1(n15390), .C2(n10889), .A(n10888), .B(n10887), .ZN(
        n10896) );
  AOI22_X1 U13430 ( .A1(n10890), .A2(n14248), .B1(n6794), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n10891) );
  OAI21_X1 U13431 ( .B1(n10896), .B2(n6794), .A(n10891), .ZN(P2_U3508) );
  INV_X1 U13432 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10892) );
  OAI22_X1 U13433 ( .A1(n10893), .A2(n14287), .B1(n15393), .B2(n10892), .ZN(
        n10894) );
  INV_X1 U13434 ( .A(n10894), .ZN(n10895) );
  OAI21_X1 U13435 ( .B1(n10896), .B2(n15391), .A(n10895), .ZN(P2_U3457) );
  XNOR2_X1 U13436 ( .A(n10906), .B(n13792), .ZN(n11212) );
  NAND2_X1 U13437 ( .A1(n13907), .A2(n13997), .ZN(n11211) );
  XNOR2_X1 U13438 ( .A(n11212), .B(n11211), .ZN(n11214) );
  XNOR2_X1 U13439 ( .A(n11215), .B(n11214), .ZN(n10908) );
  INV_X1 U13440 ( .A(n10899), .ZN(n10901) );
  OAI21_X1 U13441 ( .B1(n15111), .B2(n10901), .A(n10900), .ZN(n10905) );
  OAI22_X1 U13442 ( .A1(n13883), .A2(n10903), .B1(n13881), .B2(n10902), .ZN(
        n10904) );
  AOI211_X1 U13443 ( .C1(n10906), .C2(n15107), .A(n10905), .B(n10904), .ZN(
        n10907) );
  OAI21_X1 U13444 ( .B1(n10908), .B2(n13872), .A(n10907), .ZN(P2_U3189) );
  NAND2_X1 U13445 ( .A1(n10912), .A2(n10909), .ZN(n10910) );
  XNOR2_X1 U13446 ( .A(n10925), .B(n12771), .ZN(n11029) );
  XNOR2_X1 U13447 ( .A(n11029), .B(n15459), .ZN(n11031) );
  XOR2_X1 U13448 ( .A(n11032), .B(n11031), .Z(n10918) );
  OAI22_X1 U13449 ( .A1(n11173), .A2(n12867), .B1(n10912), .B2(n12880), .ZN(
        n10913) );
  AOI211_X1 U13450 ( .C1(n12869), .C2(n10915), .A(n10914), .B(n10913), .ZN(
        n10917) );
  NAND2_X1 U13451 ( .A1(n12882), .A2(n10926), .ZN(n10916) );
  OAI211_X1 U13452 ( .C1(n10918), .C2(n12872), .A(n10917), .B(n10916), .ZN(
        P3_U3167) );
  INV_X1 U13453 ( .A(n15462), .ZN(n10919) );
  AOI21_X1 U13454 ( .B1(n12202), .B2(n10920), .A(n10919), .ZN(n10924) );
  AOI22_X1 U13455 ( .A1(n15515), .A2(n15474), .B1(n12895), .B2(n15517), .ZN(
        n10923) );
  XNOR2_X1 U13456 ( .A(n10921), .B(n12202), .ZN(n15553) );
  NAND2_X1 U13457 ( .A1(n15553), .A2(n15502), .ZN(n10922) );
  OAI211_X1 U13458 ( .C1(n10924), .C2(n15497), .A(n10923), .B(n10922), .ZN(
        n15551) );
  INV_X1 U13459 ( .A(n15551), .ZN(n10931) );
  INV_X1 U13460 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10928) );
  NOR2_X1 U13461 ( .A1(n10925), .A2(n15559), .ZN(n15552) );
  AOI22_X1 U13462 ( .A1(n15552), .A2(n15485), .B1(n15508), .B2(n10926), .ZN(
        n10927) );
  OAI21_X1 U13463 ( .B1(n10928), .B2(n15530), .A(n10927), .ZN(n10929) );
  AOI21_X1 U13464 ( .B1(n15553), .B2(n15444), .A(n10929), .ZN(n10930) );
  OAI21_X1 U13465 ( .B1(n10931), .B2(n15489), .A(n10930), .ZN(P3_U3228) );
  OAI21_X1 U13466 ( .B1(n10939), .B2(n11461), .A(n10932), .ZN(n10933) );
  INV_X1 U13467 ( .A(n10933), .ZN(n10934) );
  XNOR2_X1 U13468 ( .A(n10933), .B(n11642), .ZN(n15204) );
  NOR2_X1 U13469 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15204), .ZN(n15203) );
  AOI21_X1 U13470 ( .B1(n10934), .B2(n15211), .A(n15203), .ZN(n10937) );
  INV_X1 U13471 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11392) );
  NOR2_X1 U13472 ( .A1(n11393), .A2(n11392), .ZN(n10935) );
  AOI21_X1 U13473 ( .B1(n11392), .B2(n11393), .A(n10935), .ZN(n10936) );
  NAND2_X1 U13474 ( .A1(n10936), .A2(n10937), .ZN(n11391) );
  OAI211_X1 U13475 ( .C1(n10937), .C2(n10936), .A(n14576), .B(n11391), .ZN(
        n10947) );
  NAND2_X1 U13476 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14371)
         );
  AOI21_X1 U13477 ( .B1(n11434), .B2(n10939), .A(n10938), .ZN(n10940) );
  INV_X1 U13478 ( .A(n10940), .ZN(n10941) );
  XNOR2_X1 U13479 ( .A(n10940), .B(n11642), .ZN(n15206) );
  NOR2_X1 U13480 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n15206), .ZN(n15205) );
  AOI21_X1 U13481 ( .B1(n15211), .B2(n10941), .A(n15205), .ZN(n10943) );
  XNOR2_X1 U13482 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n11393), .ZN(n10942) );
  NAND2_X1 U13483 ( .A1(n10942), .A2(n10943), .ZN(n11387) );
  OAI211_X1 U13484 ( .C1(n10943), .C2(n10942), .A(n14565), .B(n11387), .ZN(
        n10944) );
  NAND2_X1 U13485 ( .A1(n14371), .A2(n10944), .ZN(n10945) );
  AOI21_X1 U13486 ( .B1(n15199), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10945), 
        .ZN(n10946) );
  OAI211_X1 U13487 ( .C1(n15212), .C2(n11393), .A(n10947), .B(n10946), .ZN(
        P1_U3259) );
  NAND2_X1 U13488 ( .A1(n10948), .A2(n14856), .ZN(n10957) );
  NOR2_X1 U13489 ( .A1(n10949), .A2(n14783), .ZN(n10955) );
  MUX2_X1 U13490 ( .A(n10951), .B(n10950), .S(n14855), .Z(n10952) );
  OAI21_X1 U13491 ( .B1(n14852), .B2(n10953), .A(n10952), .ZN(n10954) );
  AOI211_X1 U13492 ( .C1(n14858), .C2(n12345), .A(n10955), .B(n10954), .ZN(
        n10956) );
  OAI211_X1 U13493 ( .C1(n10958), .C2(n14838), .A(n10957), .B(n10956), .ZN(
        P1_U3286) );
  NAND2_X1 U13494 ( .A1(n10959), .A2(n14856), .ZN(n10967) );
  MUX2_X1 U13495 ( .A(n10961), .B(n10960), .S(n14855), .Z(n10962) );
  OAI21_X1 U13496 ( .B1(n14852), .B2(n11053), .A(n10962), .ZN(n10965) );
  NOR2_X1 U13497 ( .A1(n10963), .A2(n14783), .ZN(n10964) );
  AOI211_X1 U13498 ( .C1(n14858), .C2(n12356), .A(n10965), .B(n10964), .ZN(
        n10966) );
  OAI211_X1 U13499 ( .C1(n10968), .C2(n14838), .A(n10967), .B(n10966), .ZN(
        P1_U3284) );
  INV_X1 U13500 ( .A(n10969), .ZN(n10970) );
  INV_X1 U13501 ( .A(n14852), .ZN(n14842) );
  AOI22_X1 U13502 ( .A1(n14840), .A2(n10971), .B1(n10970), .B2(n14842), .ZN(
        n10972) );
  OAI21_X1 U13503 ( .B1(n13476), .B2(n14840), .A(n10972), .ZN(n10975) );
  NOR2_X1 U13504 ( .A1(n10973), .A2(n14783), .ZN(n10974) );
  AOI211_X1 U13505 ( .C1(n14858), .C2(n12351), .A(n10975), .B(n10974), .ZN(
        n10978) );
  NAND2_X1 U13506 ( .A1(n10976), .A2(n14856), .ZN(n10977) );
  OAI211_X1 U13507 ( .C1(n10979), .C2(n14838), .A(n10978), .B(n10977), .ZN(
        P1_U3285) );
  XNOR2_X1 U13508 ( .A(n10980), .B(n10981), .ZN(n10986) );
  XNOR2_X1 U13509 ( .A(n10982), .B(n10981), .ZN(n10984) );
  OAI22_X1 U13510 ( .A1(n11417), .A2(n15098), .B1(n11226), .B2(n15096), .ZN(
        n10983) );
  AOI21_X1 U13511 ( .B1(n10984), .B2(n6580), .A(n10983), .ZN(n10985) );
  OAI21_X1 U13512 ( .B1(n10986), .B2(n9899), .A(n10985), .ZN(n15387) );
  INV_X1 U13513 ( .A(n15387), .ZN(n10992) );
  INV_X1 U13514 ( .A(n10986), .ZN(n15389) );
  OAI211_X1 U13515 ( .C1(n8991), .C2(n10809), .A(n10037), .B(n15136), .ZN(
        n15385) );
  AOI22_X1 U13516 ( .A1(n8990), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11224), 
        .B2(n15329), .ZN(n10989) );
  NAND2_X1 U13517 ( .A1(n11229), .A2(n15132), .ZN(n10988) );
  OAI211_X1 U13518 ( .C1(n15385), .C2(n14152), .A(n10989), .B(n10988), .ZN(
        n10990) );
  AOI21_X1 U13519 ( .B1(n15389), .B2(n14168), .A(n10990), .ZN(n10991) );
  OAI21_X1 U13520 ( .B1(n10992), .B2(n15331), .A(n10991), .ZN(P2_U3254) );
  INV_X1 U13521 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10995) );
  NOR2_X1 U13522 ( .A1(n11002), .A2(n10995), .ZN(n10994) );
  AOI21_X1 U13523 ( .B1(n10995), .B2(n11002), .A(n10994), .ZN(n15290) );
  NAND2_X1 U13524 ( .A1(n15291), .A2(n15290), .ZN(n15289) );
  OAI21_X1 U13525 ( .B1(n10995), .B2(n11002), .A(n15289), .ZN(n11267) );
  XNOR2_X1 U13526 ( .A(n11278), .B(n11267), .ZN(n10996) );
  OAI211_X1 U13527 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n10996), .A(n15319), 
        .B(n11269), .ZN(n11006) );
  NAND2_X1 U13528 ( .A1(n11268), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10997) );
  OAI21_X1 U13529 ( .B1(n11268), .B2(P2_REG1_REG_14__SCAN_IN), .A(n10997), 
        .ZN(n10998) );
  INV_X1 U13530 ( .A(n10998), .ZN(n11004) );
  INV_X1 U13531 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n15154) );
  AOI21_X1 U13532 ( .B1(n15160), .B2(n11000), .A(n10999), .ZN(n15295) );
  NOR2_X1 U13533 ( .A1(n11002), .A2(n15154), .ZN(n11001) );
  AOI21_X1 U13534 ( .B1(n15154), .B2(n11002), .A(n11001), .ZN(n15294) );
  NAND2_X1 U13535 ( .A1(n15295), .A2(n15294), .ZN(n15293) );
  OAI21_X1 U13536 ( .B1(n15154), .B2(n11002), .A(n15293), .ZN(n11003) );
  NAND2_X1 U13537 ( .A1(n11003), .A2(n11004), .ZN(n11277) );
  OAI211_X1 U13538 ( .C1(n11004), .C2(n11003), .A(n15317), .B(n11277), .ZN(
        n11005) );
  NAND2_X1 U13539 ( .A1(n11006), .A2(n11005), .ZN(n11008) );
  NAND2_X1 U13540 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n15108)
         );
  INV_X1 U13541 ( .A(n15108), .ZN(n11007) );
  AOI211_X1 U13542 ( .C1(n15314), .C2(P2_ADDR_REG_14__SCAN_IN), .A(n11008), 
        .B(n11007), .ZN(n11009) );
  OAI21_X1 U13543 ( .B1(n11278), .B2(n15311), .A(n11009), .ZN(P2_U3228) );
  XNOR2_X1 U13544 ( .A(n11010), .B(n12207), .ZN(n11014) );
  NAND2_X1 U13545 ( .A1(n12894), .A2(n15517), .ZN(n11012) );
  NAND2_X1 U13546 ( .A1(n12895), .A2(n15515), .ZN(n11011) );
  NAND2_X1 U13547 ( .A1(n11012), .A2(n11011), .ZN(n11013) );
  AOI21_X1 U13548 ( .B1(n11014), .B2(n15513), .A(n11013), .ZN(n15564) );
  OR2_X1 U13549 ( .A1(n11015), .A2(n12207), .ZN(n11016) );
  NAND2_X1 U13550 ( .A1(n11017), .A2(n11016), .ZN(n15562) );
  OR2_X1 U13551 ( .A1(n15502), .A2(n15505), .ZN(n15521) );
  AOI22_X1 U13552 ( .A1(n15489), .A2(P3_REG2_REG_7__SCAN_IN), .B1(n15508), 
        .B2(n11166), .ZN(n11018) );
  OAI21_X1 U13553 ( .B1(n13587), .B2(n15560), .A(n11018), .ZN(n11019) );
  AOI21_X1 U13554 ( .B1(n15562), .B2(n15071), .A(n11019), .ZN(n11020) );
  OAI21_X1 U13555 ( .B1(n15564), .B2(n15489), .A(n11020), .ZN(P3_U3226) );
  INV_X1 U13556 ( .A(n11830), .ZN(n11024) );
  OAI21_X1 U13557 ( .B1(n11021), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n11022) );
  XNOR2_X1 U13558 ( .A(n11022), .B(P1_IR_REG_18__SCAN_IN), .ZN(n11831) );
  INV_X1 U13559 ( .A(n11831), .ZN(n11535) );
  OAI222_X1 U13560 ( .A1(n15024), .A2(n13404), .B1(n15030), .B2(n11024), .C1(
        n11535), .C2(P1_U3086), .ZN(P1_U3337) );
  INV_X1 U13561 ( .A(n13952), .ZN(n11023) );
  OAI222_X1 U13562 ( .A1(n14312), .A2(n11025), .B1(n10596), .B2(n11024), .C1(
        P2_U3088), .C2(n11023), .ZN(P2_U3309) );
  INV_X1 U13563 ( .A(n11026), .ZN(n11028) );
  OAI222_X1 U13564 ( .A1(n12060), .A2(P3_U3151), .B1(n13756), .B2(n11028), 
        .C1(n11027), .C2(n12609), .ZN(P3_U3274) );
  INV_X1 U13565 ( .A(n15470), .ZN(n11041) );
  INV_X1 U13566 ( .A(n11029), .ZN(n11030) );
  XNOR2_X1 U13567 ( .A(n11038), .B(n6801), .ZN(n11167) );
  XNOR2_X1 U13568 ( .A(n11167), .B(n12895), .ZN(n11033) );
  OAI211_X1 U13569 ( .C1(n11034), .C2(n11033), .A(n11170), .B(n12874), .ZN(
        n11040) );
  OAI22_X1 U13570 ( .A1(n15451), .A2(n12867), .B1(n11035), .B2(n12880), .ZN(
        n11036) );
  AOI211_X1 U13571 ( .C1(n12869), .C2(n11038), .A(n11037), .B(n11036), .ZN(
        n11039) );
  OAI211_X1 U13572 ( .C1(n11041), .C2(n11604), .A(n11040), .B(n11039), .ZN(
        P3_U3179) );
  INV_X1 U13573 ( .A(n11042), .ZN(n11044) );
  OAI22_X1 U13574 ( .A1(n12236), .A2(P3_U3151), .B1(SI_22_), .B2(n12609), .ZN(
        n11043) );
  AOI21_X1 U13575 ( .B1(n11044), .B2(n13749), .A(n11043), .ZN(P3_U3273) );
  NAND2_X1 U13576 ( .A1(n11046), .A2(n11045), .ZN(n11047) );
  AOI22_X1 U13577 ( .A1(n12356), .A2(n10103), .B1(n12709), .B2(n14468), .ZN(
        n11191) );
  INV_X1 U13578 ( .A(n11191), .ZN(n11049) );
  AOI22_X1 U13579 ( .A1(n12356), .A2(n12708), .B1(n10103), .B2(n14468), .ZN(
        n11050) );
  XOR2_X1 U13580 ( .A(n12710), .B(n11050), .Z(n11051) );
  NAND2_X1 U13581 ( .A1(n11052), .A2(n11051), .ZN(n11193) );
  OAI211_X1 U13582 ( .C1(n11052), .C2(n11051), .A(n11193), .B(n14425), .ZN(
        n11057) );
  NOR2_X1 U13583 ( .A1(n14441), .A2(n11053), .ZN(n11055) );
  INV_X1 U13584 ( .A(n14467), .ZN(n11135) );
  NAND2_X1 U13585 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n14568) );
  OAI21_X1 U13586 ( .B1(n14449), .B2(n11135), .A(n14568), .ZN(n11054) );
  AOI211_X1 U13587 ( .C1(n14447), .C2(n14469), .A(n11055), .B(n11054), .ZN(
        n11056) );
  OAI211_X1 U13588 ( .C1(n11058), .C2(n14450), .A(n11057), .B(n11056), .ZN(
        P1_U3231) );
  OAI21_X1 U13589 ( .B1(n11060), .B2(n11062), .A(n11059), .ZN(n15247) );
  OAI22_X1 U13590 ( .A1(n12340), .A2(n14826), .B1(n12326), .B2(n14824), .ZN(
        n11067) );
  NAND3_X1 U13591 ( .A1(n11063), .A2(n11062), .A3(n11061), .ZN(n11064) );
  AOI21_X1 U13592 ( .B1(n11065), .B2(n11064), .A(n15228), .ZN(n11066) );
  AOI211_X1 U13593 ( .C1(n14629), .C2(n15247), .A(n11067), .B(n11066), .ZN(
        n15244) );
  MUX2_X1 U13594 ( .A(n11068), .B(n15244), .S(n14840), .Z(n11075) );
  OAI211_X1 U13595 ( .C1(n15243), .C2(n11070), .A(n14888), .B(n11069), .ZN(
        n15242) );
  AOI22_X1 U13596 ( .A1(n14858), .A2(n12330), .B1(n11071), .B2(n14842), .ZN(
        n11072) );
  OAI21_X1 U13597 ( .B1(n14783), .B2(n15242), .A(n11072), .ZN(n11073) );
  AOI21_X1 U13598 ( .B1(n14846), .B2(n15247), .A(n11073), .ZN(n11074) );
  NAND2_X1 U13599 ( .A1(n11075), .A2(n11074), .ZN(P1_U3288) );
  NOR2_X1 U13600 ( .A1(n10451), .A2(n11076), .ZN(n11077) );
  INV_X1 U13601 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11079) );
  AOI21_X1 U13602 ( .B1(n11080), .B2(n11079), .A(n11233), .ZN(n11099) );
  OR2_X1 U13603 ( .A1(n6587), .A2(n11079), .ZN(n11082) );
  NAND2_X1 U13604 ( .A1(n6587), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n11081) );
  AND2_X1 U13605 ( .A1(n11082), .A2(n11081), .ZN(n11084) );
  AND2_X1 U13606 ( .A1(n11084), .A2(n11251), .ZN(n11241) );
  INV_X1 U13607 ( .A(n11241), .ZN(n11083) );
  OAI21_X1 U13608 ( .B1(n11251), .B2(n11084), .A(n11083), .ZN(n11088) );
  NOR2_X1 U13609 ( .A1(n11087), .A2(n11088), .ZN(n11240) );
  AOI21_X1 U13610 ( .B1(n11088), .B2(n11087), .A(n11240), .ZN(n11091) );
  INV_X1 U13611 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n11089) );
  NOR2_X1 U13612 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11089), .ZN(n11175) );
  AOI21_X1 U13613 ( .B1(n15417), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11175), .ZN(
        n11090) );
  OAI21_X1 U13614 ( .B1(n11091), .B2(n15406), .A(n11090), .ZN(n11097) );
  INV_X1 U13615 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15594) );
  XNOR2_X1 U13616 ( .A(n11251), .B(n11250), .ZN(n11094) );
  AOI21_X1 U13617 ( .B1(n15594), .B2(n11094), .A(n11252), .ZN(n11095) );
  NOR2_X1 U13618 ( .A1(n11095), .A2(n15407), .ZN(n11096) );
  AOI211_X1 U13619 ( .C1(n15421), .C2(n11251), .A(n11097), .B(n11096), .ZN(
        n11098) );
  OAI21_X1 U13620 ( .B1(n11099), .B2(n15408), .A(n11098), .ZN(P3_U3189) );
  INV_X1 U13621 ( .A(n11843), .ZN(n11101) );
  OAI222_X1 U13622 ( .A1(P1_U3086), .A2(n11695), .B1(n15030), .B2(n11101), 
        .C1(n11100), .C2(n15024), .ZN(P1_U3336) );
  OAI222_X1 U13623 ( .A1(n14312), .A2(n11102), .B1(n10596), .B2(n11101), .C1(
        P2_U3088), .C2(n11795), .ZN(P2_U3308) );
  INV_X1 U13624 ( .A(n11858), .ZN(n11164) );
  OAI222_X1 U13625 ( .A1(n10596), .A2(n11164), .B1(n11104), .B2(P2_U3088), 
        .C1(n11103), .C2(n14312), .ZN(P2_U3307) );
  NAND2_X1 U13626 ( .A1(n12356), .A2(n11201), .ZN(n11105) );
  NAND2_X1 U13627 ( .A1(n11107), .A2(n12456), .ZN(n11110) );
  AOI22_X1 U13628 ( .A1(n11845), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11108), 
        .B2(n11844), .ZN(n11109) );
  XNOR2_X1 U13629 ( .A(n15249), .B(n14467), .ZN(n12500) );
  NAND2_X1 U13630 ( .A1(n11111), .A2(n11116), .ZN(n11112) );
  NAND3_X1 U13631 ( .A1(n11137), .A2(n14939), .A3(n11112), .ZN(n11114) );
  NAND2_X1 U13632 ( .A1(n14468), .A2(n14791), .ZN(n11113) );
  NAND2_X1 U13633 ( .A1(n11114), .A2(n11113), .ZN(n15253) );
  INV_X1 U13634 ( .A(n15253), .ZN(n11134) );
  NAND2_X1 U13635 ( .A1(n11117), .A2(n11116), .ZN(n11154) );
  OAI21_X1 U13636 ( .B1(n11117), .B2(n11116), .A(n11154), .ZN(n15255) );
  INV_X1 U13637 ( .A(n11157), .ZN(n11118) );
  XNOR2_X1 U13638 ( .A(n11118), .B(n15249), .ZN(n11129) );
  NAND2_X1 U13639 ( .A1(n11985), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11127) );
  INV_X1 U13640 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11119) );
  OR2_X1 U13641 ( .A1(n11944), .A2(n11119), .ZN(n11126) );
  NAND2_X1 U13642 ( .A1(n11121), .A2(n11120), .ZN(n11122) );
  NAND2_X1 U13643 ( .A1(n11144), .A2(n11122), .ZN(n11483) );
  OR2_X1 U13644 ( .A1(n11986), .A2(n11483), .ZN(n11125) );
  OR2_X1 U13645 ( .A1(n12454), .A2(n11123), .ZN(n11124) );
  NAND4_X1 U13646 ( .A1(n11127), .A2(n11126), .A3(n11125), .A4(n11124), .ZN(
        n14466) );
  AND2_X1 U13647 ( .A1(n14466), .A2(n14850), .ZN(n11128) );
  AOI21_X1 U13648 ( .B1(n11129), .B2(n14888), .A(n11128), .ZN(n15250) );
  OAI22_X1 U13649 ( .A1(n14840), .A2(n9625), .B1(n11204), .B2(n14852), .ZN(
        n11130) );
  AOI21_X1 U13650 ( .B1(n15249), .B2(n14858), .A(n11130), .ZN(n11131) );
  OAI21_X1 U13651 ( .B1(n15250), .B2(n14783), .A(n11131), .ZN(n11132) );
  AOI21_X1 U13652 ( .B1(n15255), .B2(n14857), .A(n11132), .ZN(n11133) );
  OAI21_X1 U13653 ( .B1(n11134), .B2(n14855), .A(n11133), .ZN(P1_U3283) );
  OR2_X1 U13654 ( .A1(n15249), .A2(n11135), .ZN(n11136) );
  NAND2_X1 U13655 ( .A1(n11138), .A2(n12456), .ZN(n11141) );
  AOI22_X1 U13656 ( .A1(n11845), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11844), 
        .B2(n11139), .ZN(n11140) );
  XNOR2_X1 U13657 ( .A(n12369), .B(n14466), .ZN(n12501) );
  XNOR2_X1 U13658 ( .A(n11294), .B(n11155), .ZN(n11142) );
  NAND2_X1 U13659 ( .A1(n11142), .A2(n14939), .ZN(n11152) );
  AND2_X1 U13660 ( .A1(n11144), .A2(n11143), .ZN(n11145) );
  NOR2_X1 U13661 ( .A1(n11287), .A2(n11145), .ZN(n11570) );
  NAND2_X1 U13662 ( .A1(n11878), .A2(n11570), .ZN(n11150) );
  INV_X1 U13663 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11146) );
  OR2_X1 U13664 ( .A1(n11944), .A2(n11146), .ZN(n11149) );
  OR2_X1 U13665 ( .A1(n12454), .A2(n9695), .ZN(n11148) );
  OR2_X1 U13666 ( .A1(n12289), .A2(n9688), .ZN(n11147) );
  NAND4_X1 U13667 ( .A1(n11150), .A2(n11149), .A3(n11148), .A4(n11147), .ZN(
        n14465) );
  AOI22_X1 U13668 ( .A1(n14791), .A2(n14467), .B1(n14465), .B2(n14850), .ZN(
        n11151) );
  NAND2_X1 U13669 ( .A1(n11152), .A2(n11151), .ZN(n15169) );
  INV_X1 U13670 ( .A(n15169), .ZN(n11163) );
  OR2_X1 U13671 ( .A1(n15249), .A2(n14467), .ZN(n11153) );
  OAI21_X1 U13672 ( .B1(n11156), .B2(n11155), .A(n11302), .ZN(n15171) );
  INV_X1 U13673 ( .A(n12369), .ZN(n15168) );
  NAND2_X1 U13674 ( .A1(n15168), .A2(n11158), .ZN(n11306) );
  OAI211_X1 U13675 ( .C1(n15168), .C2(n11158), .A(n14888), .B(n11306), .ZN(
        n15167) );
  OAI22_X1 U13676 ( .A1(n14840), .A2(n9691), .B1(n11483), .B2(n14852), .ZN(
        n11159) );
  AOI21_X1 U13677 ( .B1(n12369), .B2(n14858), .A(n11159), .ZN(n11160) );
  OAI21_X1 U13678 ( .B1(n15167), .B2(n14783), .A(n11160), .ZN(n11161) );
  AOI21_X1 U13679 ( .B1(n15171), .B2(n14857), .A(n11161), .ZN(n11162) );
  OAI21_X1 U13680 ( .B1(n11163), .B2(n14855), .A(n11162), .ZN(P1_U3282) );
  OAI222_X1 U13681 ( .A1(n11165), .A2(P1_U3086), .B1(n15030), .B2(n11164), 
        .C1(n13338), .C2(n15024), .ZN(P1_U3335) );
  INV_X1 U13682 ( .A(n11166), .ZN(n11179) );
  INV_X1 U13683 ( .A(n11167), .ZN(n11168) );
  NAND2_X1 U13684 ( .A1(n11168), .A2(n12895), .ZN(n11169) );
  NAND2_X1 U13685 ( .A1(n11170), .A2(n11169), .ZN(n11172) );
  XNOR2_X1 U13686 ( .A(n11171), .B(n12771), .ZN(n11328) );
  NAND2_X1 U13687 ( .A1(n11172), .A2(n11328), .ZN(n11331) );
  OAI211_X1 U13688 ( .C1(n11172), .C2(n11328), .A(n11331), .B(n12874), .ZN(
        n11178) );
  OAI22_X1 U13689 ( .A1(n11544), .A2(n12867), .B1(n11173), .B2(n12880), .ZN(
        n11174) );
  AOI211_X1 U13690 ( .C1(n12869), .C2(n11176), .A(n11175), .B(n11174), .ZN(
        n11177) );
  OAI211_X1 U13691 ( .C1(n11179), .C2(n11604), .A(n11178), .B(n11177), .ZN(
        P3_U3153) );
  XNOR2_X1 U13692 ( .A(n11181), .B(n11180), .ZN(n11182) );
  OAI222_X1 U13693 ( .A1(n15098), .A2(n13880), .B1(n11182), .B2(n15125), .C1(
        n15096), .C2(n11417), .ZN(n15151) );
  INV_X1 U13694 ( .A(n15151), .ZN(n11190) );
  XNOR2_X1 U13695 ( .A(n11184), .B(n11183), .ZN(n15153) );
  AOI21_X1 U13696 ( .B1(n15148), .B2(n15137), .A(n13997), .ZN(n11185) );
  NAND2_X1 U13697 ( .A1(n11185), .A2(n15120), .ZN(n15149) );
  AOI22_X1 U13698 ( .A1(n8990), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11415), 
        .B2(n15329), .ZN(n11187) );
  NAND2_X1 U13699 ( .A1(n15148), .A2(n15132), .ZN(n11186) );
  OAI211_X1 U13700 ( .C1(n15149), .C2(n14152), .A(n11187), .B(n11186), .ZN(
        n11188) );
  AOI21_X1 U13701 ( .B1(n15153), .B2(n15337), .A(n11188), .ZN(n11189) );
  OAI21_X1 U13702 ( .B1(n11190), .B2(n15331), .A(n11189), .ZN(P2_U3252) );
  NAND2_X1 U13703 ( .A1(n15249), .A2(n12708), .ZN(n11195) );
  NAND2_X1 U13704 ( .A1(n10103), .A2(n14467), .ZN(n11194) );
  NAND2_X1 U13705 ( .A1(n11195), .A2(n11194), .ZN(n11196) );
  XNOR2_X1 U13706 ( .A(n11196), .B(n12710), .ZN(n11474) );
  NAND2_X1 U13707 ( .A1(n15249), .A2(n10103), .ZN(n11198) );
  NAND2_X1 U13708 ( .A1(n12709), .A2(n14467), .ZN(n11197) );
  NAND2_X1 U13709 ( .A1(n11198), .A2(n11197), .ZN(n11471) );
  INV_X1 U13710 ( .A(n11471), .ZN(n11475) );
  XNOR2_X1 U13711 ( .A(n11474), .B(n11475), .ZN(n11199) );
  XNOR2_X1 U13712 ( .A(n11473), .B(n11199), .ZN(n11207) );
  OAI21_X1 U13713 ( .B1(n11567), .B2(n11201), .A(n11200), .ZN(n11202) );
  AOI21_X1 U13714 ( .B1(n14438), .B2(n14466), .A(n11202), .ZN(n11203) );
  OAI21_X1 U13715 ( .B1(n11204), .B2(n14441), .A(n11203), .ZN(n11205) );
  AOI21_X1 U13716 ( .B1(n15249), .B2(n9832), .A(n11205), .ZN(n11206) );
  OAI21_X1 U13717 ( .B1(n11207), .B2(n14456), .A(n11206), .ZN(P1_U3217) );
  NAND2_X1 U13718 ( .A1(n11208), .A2(n13749), .ZN(n11209) );
  OAI211_X1 U13719 ( .C1(n11210), .C2(n12609), .A(n11209), .B(n12235), .ZN(
        P3_U3272) );
  XNOR2_X1 U13720 ( .A(n11229), .B(n13792), .ZN(n11216) );
  NAND2_X1 U13721 ( .A1(n13906), .A2(n13997), .ZN(n11217) );
  NAND2_X1 U13722 ( .A1(n11216), .A2(n11217), .ZN(n11312) );
  INV_X1 U13723 ( .A(n11216), .ZN(n11219) );
  INV_X1 U13724 ( .A(n11217), .ZN(n11218) );
  NAND2_X1 U13725 ( .A1(n11219), .A2(n11218), .ZN(n11220) );
  NAND2_X1 U13726 ( .A1(n11312), .A2(n11220), .ZN(n11222) );
  INV_X1 U13727 ( .A(n11313), .ZN(n11221) );
  AOI21_X1 U13728 ( .B1(n11223), .B2(n11222), .A(n11221), .ZN(n11231) );
  INV_X1 U13729 ( .A(n11224), .ZN(n11225) );
  NAND2_X1 U13730 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n13938)
         );
  OAI21_X1 U13731 ( .B1(n15111), .B2(n11225), .A(n13938), .ZN(n11228) );
  OAI22_X1 U13732 ( .A1(n13883), .A2(n11417), .B1(n13881), .B2(n11226), .ZN(
        n11227) );
  AOI211_X1 U13733 ( .C1(n11229), .C2(n15107), .A(n11228), .B(n11227), .ZN(
        n11230) );
  OAI21_X1 U13734 ( .B1(n11231), .B2(n13872), .A(n11230), .ZN(P2_U3208) );
  NOR2_X1 U13735 ( .A1(n11251), .A2(n11232), .ZN(n11234) );
  NAND2_X1 U13736 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n11254), .ZN(n11235) );
  OAI21_X1 U13737 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11254), .A(n11235), .ZN(
        n11339) );
  INV_X1 U13738 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11236) );
  AOI21_X1 U13739 ( .B1(n11237), .B2(n11236), .A(n11357), .ZN(n11263) );
  OR2_X1 U13740 ( .A1(n6587), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11239) );
  INV_X1 U13741 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15596) );
  NAND2_X1 U13742 ( .A1(n6587), .A2(n15596), .ZN(n11238) );
  NAND2_X1 U13743 ( .A1(n11239), .A2(n11238), .ZN(n11243) );
  INV_X1 U13744 ( .A(n11254), .ZN(n11352) );
  AND2_X1 U13745 ( .A1(n11243), .A2(n11352), .ZN(n11244) );
  NOR2_X1 U13746 ( .A1(n11241), .A2(n11240), .ZN(n11341) );
  INV_X1 U13747 ( .A(n11244), .ZN(n11242) );
  OAI21_X1 U13748 ( .B1(n11352), .B2(n11243), .A(n11242), .ZN(n11342) );
  OR2_X1 U13749 ( .A1(n6587), .A2(n11236), .ZN(n11246) );
  NAND2_X1 U13750 ( .A1(n6587), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n11245) );
  AND2_X1 U13751 ( .A1(n11246), .A2(n11245), .ZN(n11247) );
  AND2_X1 U13752 ( .A1(n11247), .A2(n11374), .ZN(n11360) );
  NOR2_X1 U13753 ( .A1(n11247), .A2(n11374), .ZN(n11363) );
  NOR2_X1 U13754 ( .A1(n11360), .A2(n11363), .ZN(n11248) );
  XNOR2_X1 U13755 ( .A(n11362), .B(n11248), .ZN(n11249) );
  OR2_X1 U13756 ( .A1(n11249), .A2(n15406), .ZN(n11262) );
  INV_X1 U13757 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15598) );
  NAND2_X1 U13758 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n11254), .ZN(n11253) );
  OAI21_X1 U13759 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n11254), .A(n11253), .ZN(
        n11347) );
  NOR2_X1 U13760 ( .A1(n15598), .A2(n11255), .ZN(n11375) );
  AOI21_X1 U13761 ( .B1(n15598), .B2(n11255), .A(n11375), .ZN(n11256) );
  OR2_X1 U13762 ( .A1(n11256), .A2(n15407), .ZN(n11258) );
  AND2_X1 U13763 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11547) );
  AOI21_X1 U13764 ( .B1(n15417), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11547), .ZN(
        n11257) );
  OAI211_X1 U13765 ( .C1(n12916), .C2(n11259), .A(n11258), .B(n11257), .ZN(
        n11260) );
  INV_X1 U13766 ( .A(n11260), .ZN(n11261) );
  OAI211_X1 U13767 ( .C1(n11263), .C2(n15408), .A(n11262), .B(n11261), .ZN(
        P3_U3191) );
  INV_X1 U13768 ( .A(n11868), .ZN(n11265) );
  OAI222_X1 U13769 ( .A1(P1_U3086), .A2(n12298), .B1(n15030), .B2(n11265), 
        .C1(n11869), .C2(n15024), .ZN(P1_U3334) );
  OAI222_X1 U13770 ( .A1(n14312), .A2(n11266), .B1(n10596), .B2(n11265), .C1(
        P2_U3088), .C2(n11264), .ZN(P2_U3306) );
  NAND2_X1 U13771 ( .A1(n11268), .A2(n11267), .ZN(n11270) );
  NAND2_X1 U13772 ( .A1(n15301), .A2(n11271), .ZN(n11272) );
  XNOR2_X1 U13773 ( .A(n11279), .B(n11271), .ZN(n15303) );
  NAND2_X1 U13774 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15303), .ZN(n15302) );
  NAND2_X1 U13775 ( .A1(n11272), .A2(n15302), .ZN(n11276) );
  NAND2_X1 U13776 ( .A1(n11776), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n11273) );
  OAI21_X1 U13777 ( .B1(n11776), .B2(P2_REG2_REG_16__SCAN_IN), .A(n11273), 
        .ZN(n11275) );
  INV_X1 U13778 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11625) );
  NAND2_X1 U13779 ( .A1(n11776), .A2(n11625), .ZN(n11274) );
  OAI211_X1 U13780 ( .C1(n11276), .C2(n11275), .A(n11775), .B(n15319), .ZN(
        n11286) );
  NAND2_X1 U13781 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n13832)
         );
  XNOR2_X1 U13782 ( .A(n11776), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n11782) );
  INV_X1 U13783 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n15147) );
  OAI21_X1 U13784 ( .B1(n15147), .B2(n11278), .A(n11277), .ZN(n11280) );
  NAND2_X1 U13785 ( .A1(n15301), .A2(n11280), .ZN(n11281) );
  XNOR2_X1 U13786 ( .A(n11280), .B(n11279), .ZN(n15305) );
  NAND2_X1 U13787 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n15305), .ZN(n15304) );
  NAND2_X1 U13788 ( .A1(n11281), .A2(n15304), .ZN(n11783) );
  XOR2_X1 U13789 ( .A(n11782), .B(n11783), .Z(n11282) );
  NAND2_X1 U13790 ( .A1(n15317), .A2(n11282), .ZN(n11283) );
  NAND2_X1 U13791 ( .A1(n13832), .A2(n11283), .ZN(n11284) );
  AOI21_X1 U13792 ( .B1(n15314), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11284), 
        .ZN(n11285) );
  OAI211_X1 U13793 ( .C1(n15311), .C2(n11776), .A(n11286), .B(n11285), .ZN(
        P2_U3230) );
  OR2_X1 U13794 ( .A1(n11287), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11288) );
  NAND2_X1 U13795 ( .A1(n11287), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n11432) );
  AND2_X1 U13796 ( .A1(n11288), .A2(n11432), .ZN(n11613) );
  NAND2_X1 U13797 ( .A1(n11878), .A2(n11613), .ZN(n11293) );
  OR2_X1 U13798 ( .A1(n12289), .A2(n9873), .ZN(n11292) );
  INV_X1 U13799 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11289) );
  OR2_X1 U13800 ( .A1(n11944), .A2(n11289), .ZN(n11291) );
  OR2_X1 U13801 ( .A1(n12454), .A2(n11501), .ZN(n11290) );
  NAND4_X1 U13802 ( .A1(n11293), .A2(n11292), .A3(n11291), .A4(n11290), .ZN(
        n14464) );
  INV_X1 U13803 ( .A(n14466), .ZN(n11568) );
  OR2_X1 U13804 ( .A1(n12369), .A2(n11568), .ZN(n11295) );
  AOI22_X1 U13805 ( .A1(n11845), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n11298), 
        .B2(n11844), .ZN(n11299) );
  XNOR2_X1 U13806 ( .A(n11429), .B(n7309), .ZN(n11300) );
  OAI222_X1 U13807 ( .A1(n14826), .A2(n11611), .B1(n11300), .B2(n15228), .C1(
        n14824), .C2(n11568), .ZN(n11504) );
  INV_X1 U13808 ( .A(n11504), .ZN(n11311) );
  OR2_X1 U13809 ( .A1(n12369), .A2(n14466), .ZN(n11301) );
  OAI21_X1 U13810 ( .B1(n11304), .B2(n11303), .A(n11422), .ZN(n11506) );
  INV_X1 U13811 ( .A(n12375), .ZN(n11573) );
  INV_X1 U13812 ( .A(n11440), .ZN(n11305) );
  AOI211_X1 U13813 ( .C1(n12375), .C2(n11306), .A(n14828), .B(n11305), .ZN(
        n11505) );
  NAND2_X1 U13814 ( .A1(n11505), .A2(n14835), .ZN(n11308) );
  AOI22_X1 U13815 ( .A1(n14855), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11570), 
        .B2(n14842), .ZN(n11307) );
  OAI211_X1 U13816 ( .C1(n11573), .C2(n14831), .A(n11308), .B(n11307), .ZN(
        n11309) );
  AOI21_X1 U13817 ( .B1(n14857), .B2(n11506), .A(n11309), .ZN(n11310) );
  OAI21_X1 U13818 ( .B1(n11311), .B2(n14855), .A(n11310), .ZN(P1_U3281) );
  XNOR2_X1 U13819 ( .A(n15135), .B(n13792), .ZN(n11315) );
  NAND2_X1 U13820 ( .A1(n13905), .A2(n13997), .ZN(n11316) );
  NAND2_X1 U13821 ( .A1(n11315), .A2(n11316), .ZN(n11320) );
  NOR3_X1 U13822 ( .A1(n11315), .A2(n11417), .A3(n13817), .ZN(n11314) );
  AOI21_X1 U13823 ( .B1(n11413), .B2(n15104), .A(n11314), .ZN(n11327) );
  INV_X1 U13824 ( .A(n11315), .ZN(n11318) );
  INV_X1 U13825 ( .A(n11316), .ZN(n11317) );
  NAND2_X1 U13826 ( .A1(n11318), .A2(n11317), .ZN(n11412) );
  AOI21_X1 U13827 ( .B1(n11412), .B2(n11320), .A(n11319), .ZN(n11326) );
  NAND2_X1 U13828 ( .A1(n13906), .A2(n14025), .ZN(n11322) );
  NAND2_X1 U13829 ( .A1(n11414), .A2(n14027), .ZN(n11321) );
  AND2_X1 U13830 ( .A1(n11322), .A2(n11321), .ZN(n15127) );
  OAI22_X1 U13831 ( .A1(n13853), .A2(n15127), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13485), .ZN(n11323) );
  AOI21_X1 U13832 ( .B1(n15131), .B2(n13855), .A(n11323), .ZN(n11325) );
  NAND2_X1 U13833 ( .A1(n15135), .A2(n15107), .ZN(n11324) );
  OAI211_X1 U13834 ( .C1(n11327), .C2(n11326), .A(n11325), .B(n11324), .ZN(
        P2_U3196) );
  INV_X1 U13835 ( .A(n15454), .ZN(n11337) );
  INV_X1 U13836 ( .A(n11328), .ZN(n11329) );
  NAND2_X1 U13837 ( .A1(n11329), .A2(n15460), .ZN(n11330) );
  NAND2_X1 U13838 ( .A1(n11331), .A2(n11330), .ZN(n11332) );
  XNOR2_X1 U13839 ( .A(n15453), .B(n6801), .ZN(n11537) );
  XNOR2_X1 U13840 ( .A(n11537), .B(n12894), .ZN(n11333) );
  NAND2_X1 U13841 ( .A1(n11332), .A2(n11333), .ZN(n11540) );
  OAI211_X1 U13842 ( .C1(n11332), .C2(n11333), .A(n11540), .B(n12874), .ZN(
        n11336) );
  AND2_X1 U13843 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n11343) );
  OAI22_X1 U13844 ( .A1(n15452), .A2(n12867), .B1(n15451), .B2(n12880), .ZN(
        n11334) );
  AOI211_X1 U13845 ( .C1(n12869), .C2(n15453), .A(n11343), .B(n11334), .ZN(
        n11335) );
  OAI211_X1 U13846 ( .C1(n11337), .C2(n11604), .A(n11336), .B(n11335), .ZN(
        P3_U3161) );
  AOI21_X1 U13847 ( .B1(n6738), .B2(n11339), .A(n11338), .ZN(n11354) );
  AOI21_X1 U13848 ( .B1(n11342), .B2(n11341), .A(n11340), .ZN(n11345) );
  AOI21_X1 U13849 ( .B1(n15417), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n11343), .ZN(
        n11344) );
  OAI21_X1 U13850 ( .B1(n11345), .B2(n15406), .A(n11344), .ZN(n11351) );
  AOI21_X1 U13851 ( .B1(n11348), .B2(n11347), .A(n11346), .ZN(n11349) );
  NOR2_X1 U13852 ( .A1(n11349), .A2(n15407), .ZN(n11350) );
  AOI211_X1 U13853 ( .C1(n15421), .C2(n11352), .A(n11351), .B(n11350), .ZN(
        n11353) );
  OAI21_X1 U13854 ( .B1(n11354), .B2(n15408), .A(n11353), .ZN(P3_U3190) );
  NOR2_X1 U13855 ( .A1(n11374), .A2(n11355), .ZN(n11356) );
  NAND2_X1 U13856 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11670), .ZN(n11358) );
  OAI21_X1 U13857 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11670), .A(n11358), 
        .ZN(n11359) );
  AOI21_X1 U13858 ( .B1(n6734), .B2(n11359), .A(n11663), .ZN(n11386) );
  INV_X1 U13859 ( .A(n11360), .ZN(n11361) );
  OAI21_X1 U13860 ( .B1(n11363), .B2(n11362), .A(n11361), .ZN(n11368) );
  INV_X1 U13861 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11364) );
  OR2_X1 U13862 ( .A1(n6587), .A2(n11364), .ZN(n11366) );
  NAND2_X1 U13863 ( .A1(n6587), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n11365) );
  NAND2_X1 U13864 ( .A1(n11366), .A2(n11365), .ZN(n11669) );
  XNOR2_X1 U13865 ( .A(n11669), .B(n11383), .ZN(n11367) );
  OAI21_X1 U13866 ( .B1(n11368), .B2(n11367), .A(n11671), .ZN(n11369) );
  NAND2_X1 U13867 ( .A1(n11369), .A2(n15422), .ZN(n11385) );
  INV_X1 U13868 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11372) );
  INV_X1 U13869 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11370) );
  NOR2_X1 U13870 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11370), .ZN(n11600) );
  INV_X1 U13871 ( .A(n11600), .ZN(n11371) );
  OAI21_X1 U13872 ( .B1(n15414), .B2(n11372), .A(n11371), .ZN(n11382) );
  NOR2_X1 U13873 ( .A1(n11374), .A2(n11373), .ZN(n11376) );
  NAND2_X1 U13874 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11670), .ZN(n11377) );
  OAI21_X1 U13875 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n11670), .A(n11377), 
        .ZN(n11378) );
  AOI21_X1 U13876 ( .B1(n11379), .B2(n11378), .A(n6735), .ZN(n11380) );
  NOR2_X1 U13877 ( .A1(n11380), .A2(n15407), .ZN(n11381) );
  AOI211_X1 U13878 ( .C1(n15421), .C2(n11383), .A(n11382), .B(n11381), .ZN(
        n11384) );
  OAI211_X1 U13879 ( .C1(n11386), .C2(n15408), .A(n11385), .B(n11384), .ZN(
        P3_U3192) );
  NAND2_X1 U13880 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14382)
         );
  INV_X1 U13881 ( .A(n11393), .ZN(n11815) );
  INV_X1 U13882 ( .A(n11387), .ZN(n11388) );
  AOI21_X1 U13883 ( .B1(n11815), .B2(P1_REG1_REG_16__SCAN_IN), .A(n11388), 
        .ZN(n11528) );
  XNOR2_X1 U13884 ( .A(n11820), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n11529) );
  XOR2_X1 U13885 ( .A(n11528), .B(n11529), .Z(n11389) );
  NAND2_X1 U13886 ( .A1(n14565), .A2(n11389), .ZN(n11390) );
  NAND2_X1 U13887 ( .A1(n14382), .A2(n11390), .ZN(n11398) );
  OAI21_X1 U13888 ( .B1(n11393), .B2(n11392), .A(n11391), .ZN(n11394) );
  INV_X1 U13889 ( .A(n11394), .ZN(n11396) );
  INV_X1 U13890 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11525) );
  MUX2_X1 U13891 ( .A(n11525), .B(P1_REG2_REG_17__SCAN_IN), .S(n11820), .Z(
        n11395) );
  NOR2_X1 U13892 ( .A1(n11395), .A2(n11396), .ZN(n11523) );
  AOI211_X1 U13893 ( .C1(n11396), .C2(n11395), .A(n11523), .B(n15210), .ZN(
        n11397) );
  AOI211_X1 U13894 ( .C1(n15199), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n11398), 
        .B(n11397), .ZN(n11399) );
  OAI21_X1 U13895 ( .B1(n11527), .B2(n15212), .A(n11399), .ZN(P1_U3260) );
  XNOR2_X1 U13896 ( .A(n11400), .B(n12203), .ZN(n15572) );
  NAND2_X1 U13897 ( .A1(n15572), .A2(n15502), .ZN(n11408) );
  XNOR2_X1 U13898 ( .A(n11401), .B(n11402), .ZN(n11406) );
  NAND2_X1 U13899 ( .A1(n12894), .A2(n15515), .ZN(n11404) );
  NAND2_X1 U13900 ( .A1(n12892), .A2(n15517), .ZN(n11403) );
  NAND2_X1 U13901 ( .A1(n11404), .A2(n11403), .ZN(n11405) );
  AOI21_X1 U13902 ( .B1(n11406), .B2(n15513), .A(n11405), .ZN(n11407) );
  NOR2_X1 U13903 ( .A1(n11536), .A2(n15559), .ZN(n15571) );
  AOI22_X1 U13904 ( .A1(n15571), .A2(n15485), .B1(n15508), .B2(n11549), .ZN(
        n11409) );
  OAI21_X1 U13905 ( .B1(n11236), .B2(n15530), .A(n11409), .ZN(n11410) );
  AOI21_X1 U13906 ( .B1(n15572), .B2(n15444), .A(n11410), .ZN(n11411) );
  OAI21_X1 U13907 ( .B1(n15574), .B2(n15489), .A(n11411), .ZN(P3_U3224) );
  NAND2_X1 U13908 ( .A1(n11413), .A2(n11412), .ZN(n12537) );
  XNOR2_X1 U13909 ( .A(n15148), .B(n12592), .ZN(n12540) );
  NAND2_X1 U13910 ( .A1(n11414), .A2(n13997), .ZN(n12538) );
  XNOR2_X1 U13911 ( .A(n12540), .B(n12538), .ZN(n12536) );
  XNOR2_X1 U13912 ( .A(n12537), .B(n12536), .ZN(n11421) );
  INV_X1 U13913 ( .A(n11415), .ZN(n11416) );
  OAI22_X1 U13914 ( .A1(n15111), .A2(n11416), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8684), .ZN(n11419) );
  OAI22_X1 U13915 ( .A1(n13883), .A2(n13880), .B1(n13881), .B2(n11417), .ZN(
        n11418) );
  AOI211_X1 U13916 ( .C1(n15148), .C2(n15107), .A(n11419), .B(n11418), .ZN(
        n11420) );
  OAI21_X1 U13917 ( .B1(n11421), .B2(n13872), .A(n11420), .ZN(P2_U3206) );
  NAND2_X1 U13918 ( .A1(n11423), .A2(n12456), .ZN(n11426) );
  AOI22_X1 U13919 ( .A1(n11424), .A2(n11844), .B1(n11845), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n11425) );
  XNOR2_X1 U13920 ( .A(n12380), .B(n11611), .ZN(n12505) );
  OAI21_X1 U13921 ( .B1(n11427), .B2(n12505), .A(n11447), .ZN(n11428) );
  INV_X1 U13922 ( .A(n11428), .ZN(n11499) );
  OR2_X1 U13923 ( .A1(n12375), .A2(n7113), .ZN(n11430) );
  XNOR2_X1 U13924 ( .A(n11467), .B(n12505), .ZN(n11439) );
  NAND2_X1 U13925 ( .A1(n11432), .A2(n11431), .ZN(n11433) );
  NAND2_X1 U13926 ( .A1(n11647), .A2(n11433), .ZN(n11744) );
  OAI22_X1 U13927 ( .A1(n11744), .A2(n11986), .B1(n12454), .B2(n11434), .ZN(
        n11437) );
  NAND2_X1 U13928 ( .A1(n12450), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11435) );
  OAI21_X1 U13929 ( .B1(n11461), .B2(n12289), .A(n11435), .ZN(n11436) );
  AOI22_X1 U13930 ( .A1(n14463), .A2(n14850), .B1(n14465), .B2(n14791), .ZN(
        n11616) );
  INV_X1 U13931 ( .A(n11616), .ZN(n11438) );
  AOI21_X1 U13932 ( .B1(n11439), .B2(n14939), .A(n11438), .ZN(n11498) );
  AOI21_X1 U13933 ( .B1(n12380), .B2(n11440), .A(n7151), .ZN(n11496) );
  INV_X1 U13934 ( .A(n14659), .ZN(n11441) );
  AOI22_X1 U13935 ( .A1(n11496), .A2(n11441), .B1(n11613), .B2(n14842), .ZN(
        n11442) );
  AOI21_X1 U13936 ( .B1(n11498), .B2(n11442), .A(n14855), .ZN(n11443) );
  INV_X1 U13937 ( .A(n11443), .ZN(n11445) );
  AOI22_X1 U13938 ( .A1(n12380), .A2(n14858), .B1(n14855), .B2(
        P1_REG2_REG_13__SCAN_IN), .ZN(n11444) );
  OAI211_X1 U13939 ( .C1(n11499), .C2(n14838), .A(n11445), .B(n11444), .ZN(
        P1_U3280) );
  OR2_X1 U13940 ( .A1(n12380), .A2(n14464), .ZN(n11446) );
  AOI22_X1 U13941 ( .A1(n11450), .A2(n11844), .B1(n11845), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11451) );
  INV_X1 U13942 ( .A(n14463), .ZN(n11730) );
  NAND2_X1 U13943 ( .A1(n11746), .A2(n11730), .ZN(n12385) );
  NAND2_X1 U13944 ( .A1(n12387), .A2(n12385), .ZN(n12504) );
  INV_X1 U13945 ( .A(n12504), .ZN(n11652) );
  OAI21_X1 U13946 ( .B1(n6718), .B2(n12504), .A(n11640), .ZN(n11490) );
  XNOR2_X1 U13947 ( .A(n11647), .B(P1_REG3_REG_15__SCAN_IN), .ZN(n14453) );
  NAND2_X1 U13948 ( .A1(n14453), .A2(n11878), .ZN(n11458) );
  INV_X1 U13949 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11455) );
  NAND2_X1 U13950 ( .A1(n12450), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11454) );
  NAND2_X1 U13951 ( .A1(n11985), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11453) );
  OAI211_X1 U13952 ( .C1(n11455), .C2(n12454), .A(n11454), .B(n11453), .ZN(
        n11456) );
  INV_X1 U13953 ( .A(n11456), .ZN(n11457) );
  NAND2_X1 U13954 ( .A1(n11458), .A2(n11457), .ZN(n14462) );
  INV_X1 U13955 ( .A(n14462), .ZN(n14823) );
  OAI22_X1 U13956 ( .A1(n14823), .A2(n14826), .B1(n11611), .B2(n14824), .ZN(
        n11487) );
  INV_X1 U13957 ( .A(n11744), .ZN(n11459) );
  AOI22_X1 U13958 ( .A1(n14840), .A2(n11487), .B1(n11459), .B2(n14842), .ZN(
        n11460) );
  OAI21_X1 U13959 ( .B1(n11461), .B2(n14840), .A(n11460), .ZN(n11465) );
  AOI21_X1 U13960 ( .B1(n11746), .B2(n11462), .A(n14828), .ZN(n11463) );
  NAND2_X1 U13961 ( .A1(n11463), .A2(n11657), .ZN(n11488) );
  NOR2_X1 U13962 ( .A1(n11488), .A2(n14783), .ZN(n11464) );
  AOI211_X1 U13963 ( .C1(n14858), .C2(n11746), .A(n11465), .B(n11464), .ZN(
        n11469) );
  INV_X1 U13964 ( .A(n12505), .ZN(n11466) );
  XNOR2_X1 U13965 ( .A(n11653), .B(n12504), .ZN(n11492) );
  NAND2_X1 U13966 ( .A1(n11492), .A2(n14856), .ZN(n11468) );
  OAI211_X1 U13967 ( .C1(n11490), .C2(n14838), .A(n11469), .B(n11468), .ZN(
        P1_U3279) );
  AOI22_X1 U13968 ( .A1(n12369), .A2(n12708), .B1(n10103), .B2(n14466), .ZN(
        n11470) );
  XNOR2_X1 U13969 ( .A(n11470), .B(n12710), .ZN(n11557) );
  AOI22_X1 U13970 ( .A1(n12369), .A2(n10103), .B1(n12709), .B2(n14466), .ZN(
        n11558) );
  XNOR2_X1 U13971 ( .A(n11557), .B(n11558), .ZN(n11479) );
  OR2_X1 U13972 ( .A1(n11474), .A2(n11471), .ZN(n11472) );
  NAND2_X1 U13973 ( .A1(n11474), .A2(n11471), .ZN(n11476) );
  AOI21_X1 U13974 ( .B1(n11479), .B2(n6839), .A(n11564), .ZN(n11486) );
  OAI21_X1 U13975 ( .B1(n14449), .B2(n7113), .A(n11480), .ZN(n11481) );
  AOI21_X1 U13976 ( .B1(n14447), .B2(n14467), .A(n11481), .ZN(n11482) );
  OAI21_X1 U13977 ( .B1(n11483), .B2(n14441), .A(n11482), .ZN(n11484) );
  AOI21_X1 U13978 ( .B1(n12369), .B2(n9832), .A(n11484), .ZN(n11485) );
  OAI21_X1 U13979 ( .B1(n11486), .B2(n14456), .A(n11485), .ZN(P1_U3236) );
  AOI21_X1 U13980 ( .B1(n11746), .B2(n14966), .A(n11487), .ZN(n11489) );
  OAI211_X1 U13981 ( .C1(n11490), .C2(n15229), .A(n11489), .B(n11488), .ZN(
        n11491) );
  AOI21_X1 U13982 ( .B1(n14939), .B2(n11492), .A(n11491), .ZN(n11495) );
  NAND2_X1 U13983 ( .A1(n15257), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11493) );
  OAI21_X1 U13984 ( .B1(n11495), .B2(n15257), .A(n11493), .ZN(P1_U3501) );
  NAND2_X1 U13985 ( .A1(n15265), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11494) );
  OAI21_X1 U13986 ( .B1(n11495), .B2(n15265), .A(n11494), .ZN(P1_U3542) );
  AOI22_X1 U13987 ( .A1(n11496), .A2(n14888), .B1(n12380), .B2(n14966), .ZN(
        n11497) );
  OAI211_X1 U13988 ( .C1(n11499), .C2(n15229), .A(n11498), .B(n11497), .ZN(
        n11502) );
  NAND2_X1 U13989 ( .A1(n11502), .A2(n15267), .ZN(n11500) );
  OAI21_X1 U13990 ( .B1(n15267), .B2(n11501), .A(n11500), .ZN(P1_U3541) );
  NAND2_X1 U13991 ( .A1(n11502), .A2(n15259), .ZN(n11503) );
  OAI21_X1 U13992 ( .B1(n15259), .B2(n11289), .A(n11503), .ZN(P1_U3498) );
  AOI211_X1 U13993 ( .C1(n15256), .C2(n11506), .A(n11505), .B(n11504), .ZN(
        n11510) );
  OAI22_X1 U13994 ( .A1(n11573), .A2(n15011), .B1(n15259), .B2(n11146), .ZN(
        n11507) );
  INV_X1 U13995 ( .A(n11507), .ZN(n11508) );
  OAI21_X1 U13996 ( .B1(n11510), .B2(n15257), .A(n11508), .ZN(P1_U3495) );
  AOI22_X1 U13997 ( .A1(n12375), .A2(n14900), .B1(n15265), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n11509) );
  OAI21_X1 U13998 ( .B1(n11510), .B2(n15265), .A(n11509), .ZN(P1_U3540) );
  XNOR2_X1 U13999 ( .A(n11511), .B(n11513), .ZN(n14260) );
  OAI211_X1 U14000 ( .C1(n11514), .C2(n11513), .A(n11512), .B(n6580), .ZN(
        n11516) );
  AOI22_X1 U14001 ( .A1(n13902), .A2(n14027), .B1(n14025), .B2(n13904), .ZN(
        n11515) );
  NAND2_X1 U14002 ( .A1(n11516), .A2(n11515), .ZN(n14255) );
  NOR2_X1 U14003 ( .A1(n14147), .A2(n13879), .ZN(n11517) );
  OAI21_X1 U14004 ( .B1(n14255), .B2(n11517), .A(n14163), .ZN(n11522) );
  XNOR2_X1 U14005 ( .A(n15121), .B(n14257), .ZN(n11518) );
  NOR2_X1 U14006 ( .A1(n11518), .A2(n13997), .ZN(n14256) );
  INV_X1 U14007 ( .A(n14257), .ZN(n13889) );
  OAI22_X1 U14008 ( .A1(n13889), .A2(n15334), .B1(n11519), .B2(n14163), .ZN(
        n11520) );
  AOI21_X1 U14009 ( .B1(n14256), .B2(n6581), .A(n11520), .ZN(n11521) );
  OAI211_X1 U14010 ( .C1(n14260), .C2(n14137), .A(n11522), .B(n11521), .ZN(
        P2_U3250) );
  INV_X1 U14011 ( .A(n11523), .ZN(n11524) );
  OAI21_X1 U14012 ( .B1(n11525), .B2(n11527), .A(n11524), .ZN(n11686) );
  XNOR2_X1 U14013 ( .A(n11686), .B(n11535), .ZN(n11526) );
  NAND2_X1 U14014 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n11526), .ZN(n11688) );
  OAI211_X1 U14015 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n11526), .A(n14576), 
        .B(n11688), .ZN(n11534) );
  NAND2_X1 U14016 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14420)
         );
  INV_X1 U14017 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13374) );
  OAI22_X1 U14018 ( .A1(n11529), .A2(n11528), .B1(n13374), .B2(n11527), .ZN(
        n11682) );
  XNOR2_X1 U14019 ( .A(n11535), .B(n11682), .ZN(n11530) );
  NAND2_X1 U14020 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n11530), .ZN(n11684) );
  OAI211_X1 U14021 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n11530), .A(n14565), 
        .B(n11684), .ZN(n11531) );
  NAND2_X1 U14022 ( .A1(n14420), .A2(n11531), .ZN(n11532) );
  AOI21_X1 U14023 ( .B1(n15199), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n11532), 
        .ZN(n11533) );
  OAI211_X1 U14024 ( .C1(n15212), .C2(n11535), .A(n11534), .B(n11533), .ZN(
        P1_U3261) );
  XNOR2_X1 U14025 ( .A(n11536), .B(n6801), .ZN(n11592) );
  XNOR2_X1 U14026 ( .A(n11592), .B(n12893), .ZN(n11543) );
  INV_X1 U14027 ( .A(n11537), .ZN(n11538) );
  NAND2_X1 U14028 ( .A1(n11538), .A2(n12894), .ZN(n11539) );
  INV_X1 U14029 ( .A(n11595), .ZN(n11541) );
  AOI21_X1 U14030 ( .B1(n11543), .B2(n11542), .A(n11541), .ZN(n11552) );
  OAI22_X1 U14031 ( .A1(n11545), .A2(n12867), .B1(n11544), .B2(n12880), .ZN(
        n11546) );
  AOI211_X1 U14032 ( .C1(n12869), .C2(n11548), .A(n11547), .B(n11546), .ZN(
        n11551) );
  NAND2_X1 U14033 ( .A1(n12882), .A2(n11549), .ZN(n11550) );
  OAI211_X1 U14034 ( .C1(n11552), .C2(n12872), .A(n11551), .B(n11550), .ZN(
        P3_U3171) );
  NAND2_X1 U14035 ( .A1(n12375), .A2(n12708), .ZN(n11554) );
  NAND2_X1 U14036 ( .A1(n10103), .A2(n14465), .ZN(n11553) );
  NAND2_X1 U14037 ( .A1(n11554), .A2(n11553), .ZN(n11555) );
  XNOR2_X1 U14038 ( .A(n11555), .B(n11728), .ZN(n11606) );
  NOR2_X1 U14039 ( .A1(n6812), .A2(n7113), .ZN(n11556) );
  AOI21_X1 U14040 ( .B1(n12375), .B2(n10103), .A(n11556), .ZN(n11607) );
  XNOR2_X1 U14041 ( .A(n11606), .B(n11607), .ZN(n11562) );
  INV_X1 U14042 ( .A(n11557), .ZN(n11560) );
  INV_X1 U14043 ( .A(n11558), .ZN(n11559) );
  NOR2_X1 U14044 ( .A1(n11560), .A2(n11559), .ZN(n11563) );
  OAI21_X1 U14045 ( .B1(n11564), .B2(n11563), .A(n11562), .ZN(n11565) );
  NAND3_X1 U14046 ( .A1(n6723), .A2(n14425), .A3(n11565), .ZN(n11572) );
  AOI22_X1 U14047 ( .A1(n14438), .A2(n14464), .B1(P1_REG3_REG_12__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11566) );
  OAI21_X1 U14048 ( .B1(n11568), .B2(n11567), .A(n11566), .ZN(n11569) );
  AOI21_X1 U14049 ( .B1(n11570), .B2(n14454), .A(n11569), .ZN(n11571) );
  OAI211_X1 U14050 ( .C1(n11573), .C2(n14450), .A(n11572), .B(n11571), .ZN(
        P1_U3224) );
  NAND2_X1 U14051 ( .A1(n11889), .A2(n11574), .ZN(n11575) );
  OAI211_X1 U14052 ( .C1(n11890), .C2(n15024), .A(n11575), .B(n12531), .ZN(
        P1_U3332) );
  NAND2_X1 U14053 ( .A1(n11889), .A2(n14306), .ZN(n11577) );
  OAI211_X1 U14054 ( .C1(n11578), .C2(n14312), .A(n11577), .B(n11576), .ZN(
        P2_U3304) );
  XNOR2_X1 U14055 ( .A(n13569), .B(n12208), .ZN(n11579) );
  NAND2_X1 U14056 ( .A1(n11579), .A2(n15513), .ZN(n11581) );
  AOI22_X1 U14057 ( .A1(n15517), .A2(n12891), .B1(n12892), .B2(n15515), .ZN(
        n11580) );
  NAND2_X1 U14058 ( .A1(n11581), .A2(n11580), .ZN(n15088) );
  INV_X1 U14059 ( .A(n15088), .ZN(n11587) );
  XNOR2_X1 U14060 ( .A(n11582), .B(n12208), .ZN(n15084) );
  AOI22_X1 U14061 ( .A1(n15489), .A2(P3_REG2_REG_11__SCAN_IN), .B1(n15508), 
        .B2(n12846), .ZN(n11583) );
  OAI21_X1 U14062 ( .B1(n13587), .B2(n11584), .A(n11583), .ZN(n11585) );
  AOI21_X1 U14063 ( .B1(n15084), .B2(n15071), .A(n11585), .ZN(n11586) );
  OAI21_X1 U14064 ( .B1(n11587), .B2(n15489), .A(n11586), .ZN(P3_U3222) );
  INV_X1 U14065 ( .A(n11588), .ZN(n11589) );
  OAI222_X1 U14066 ( .A1(n11591), .A2(P3_U3151), .B1(n12609), .B2(n11590), 
        .C1(n13756), .C2(n11589), .ZN(P3_U3271) );
  INV_X1 U14067 ( .A(n15442), .ZN(n11605) );
  INV_X1 U14068 ( .A(n11592), .ZN(n11593) );
  NAND2_X1 U14069 ( .A1(n15452), .A2(n11593), .ZN(n11594) );
  XNOR2_X1 U14070 ( .A(n15443), .B(n6801), .ZN(n12238) );
  XNOR2_X1 U14071 ( .A(n12238), .B(n12892), .ZN(n11596) );
  AOI21_X1 U14072 ( .B1(n11597), .B2(n11596), .A(n12872), .ZN(n11598) );
  NAND2_X1 U14073 ( .A1(n11598), .A2(n12240), .ZN(n11603) );
  OAI22_X1 U14074 ( .A1(n15435), .A2(n12867), .B1(n15452), .B2(n12880), .ZN(
        n11599) );
  AOI211_X1 U14075 ( .C1(n12869), .C2(n11601), .A(n11600), .B(n11599), .ZN(
        n11602) );
  OAI211_X1 U14076 ( .C1(n11605), .C2(n11604), .A(n11603), .B(n11602), .ZN(
        P3_U3157) );
  INV_X1 U14077 ( .A(n11606), .ZN(n11609) );
  INV_X1 U14078 ( .A(n11607), .ZN(n11608) );
  AOI22_X1 U14079 ( .A1(n12380), .A2(n12708), .B1(n10103), .B2(n14464), .ZN(
        n11610) );
  XNOR2_X1 U14080 ( .A(n11610), .B(n12710), .ZN(n11734) );
  NOR2_X1 U14081 ( .A1(n6812), .A2(n11611), .ZN(n11612) );
  AOI21_X1 U14082 ( .B1(n12380), .B2(n10103), .A(n11612), .ZN(n11735) );
  XNOR2_X1 U14083 ( .A(n11734), .B(n11735), .ZN(n11736) );
  XNOR2_X1 U14084 ( .A(n11737), .B(n11736), .ZN(n11619) );
  NAND2_X1 U14085 ( .A1(n14454), .A2(n11613), .ZN(n11615) );
  OAI211_X1 U14086 ( .C1(n11616), .C2(n14410), .A(n11615), .B(n11614), .ZN(
        n11617) );
  AOI21_X1 U14087 ( .B1(n12380), .B2(n9832), .A(n11617), .ZN(n11618) );
  OAI21_X1 U14088 ( .B1(n11619), .B2(n14456), .A(n11618), .ZN(P1_U3234) );
  OAI21_X1 U14089 ( .B1(n11621), .B2(n8725), .A(n11620), .ZN(n14254) );
  INV_X1 U14090 ( .A(n11622), .ZN(n11624) );
  INV_X1 U14091 ( .A(n11708), .ZN(n11623) );
  AOI211_X1 U14092 ( .C1(n14251), .C2(n11624), .A(n13997), .B(n11623), .ZN(
        n14250) );
  OAI22_X1 U14093 ( .A1(n11626), .A2(n15334), .B1(n14163), .B2(n11625), .ZN(
        n11627) );
  AOI21_X1 U14094 ( .B1(n14250), .B2(n6581), .A(n11627), .ZN(n11635) );
  OAI211_X1 U14095 ( .C1(n11630), .C2(n11629), .A(n11628), .B(n6580), .ZN(
        n11632) );
  AOI22_X1 U14096 ( .A1(n13901), .A2(n14027), .B1(n14025), .B2(n13903), .ZN(
        n11631) );
  AND2_X1 U14097 ( .A1(n11632), .A2(n11631), .ZN(n14252) );
  OAI21_X1 U14098 ( .B1(n13833), .B2(n14147), .A(n14252), .ZN(n11633) );
  NAND2_X1 U14099 ( .A1(n11633), .A2(n14163), .ZN(n11634) );
  OAI211_X1 U14100 ( .C1(n14254), .C2(n14137), .A(n11635), .B(n11634), .ZN(
        P2_U3249) );
  INV_X1 U14101 ( .A(n11636), .ZN(n11637) );
  OAI222_X1 U14102 ( .A1(n11638), .A2(P3_U3151), .B1(n12609), .B2(n13365), 
        .C1(n13756), .C2(n11637), .ZN(P3_U3270) );
  NAND2_X1 U14103 ( .A1(n11746), .A2(n14463), .ZN(n11639) );
  NAND2_X1 U14104 ( .A1(n11641), .A2(n12456), .ZN(n11644) );
  AOI22_X1 U14105 ( .A1(n11845), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11844), 
        .B2(n11642), .ZN(n11643) );
  NAND2_X1 U14106 ( .A1(n14967), .A2(n14823), .ZN(n12396) );
  NAND2_X1 U14107 ( .A1(n12388), .A2(n12396), .ZN(n12506) );
  XNOR2_X1 U14108 ( .A(n11812), .B(n12506), .ZN(n14969) );
  INV_X1 U14109 ( .A(n11647), .ZN(n11645) );
  AOI21_X1 U14110 ( .B1(n11645), .B2(P1_REG3_REG_15__SCAN_IN), .A(
        P1_REG3_REG_16__SCAN_IN), .ZN(n11648) );
  NAND2_X1 U14111 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n11646) );
  OR2_X1 U14112 ( .A1(n11648), .A2(n11823), .ZN(n14832) );
  AOI22_X1 U14113 ( .A1(n11985), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n12450), 
        .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n11651) );
  INV_X1 U14114 ( .A(n12454), .ZN(n11874) );
  NAND2_X1 U14115 ( .A1(n11874), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11650) );
  OAI211_X1 U14116 ( .C1(n14832), .C2(n11986), .A(n11651), .B(n11650), .ZN(
        n14461) );
  INV_X1 U14117 ( .A(n14461), .ZN(n14805) );
  NAND2_X1 U14118 ( .A1(n11653), .A2(n11652), .ZN(n11654) );
  NAND2_X1 U14119 ( .A1(n11654), .A2(n12387), .ZN(n11964) );
  INV_X1 U14120 ( .A(n12506), .ZN(n11963) );
  XNOR2_X1 U14121 ( .A(n11964), .B(n11963), .ZN(n11655) );
  OAI222_X1 U14122 ( .A1(n14826), .A2(n14805), .B1(n14824), .B2(n11730), .C1(
        n15228), .C2(n11655), .ZN(n14964) );
  NAND2_X1 U14123 ( .A1(n14964), .A2(n14840), .ZN(n11661) );
  INV_X1 U14124 ( .A(n14829), .ZN(n11656) );
  AOI211_X1 U14125 ( .C1(n14967), .C2(n11657), .A(n14828), .B(n11656), .ZN(
        n14965) );
  AOI22_X1 U14126 ( .A1(n14855), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n14453), 
        .B2(n14842), .ZN(n11658) );
  OAI21_X1 U14127 ( .B1(n7152), .B2(n14831), .A(n11658), .ZN(n11659) );
  AOI21_X1 U14128 ( .B1(n14965), .B2(n14835), .A(n11659), .ZN(n11660) );
  OAI211_X1 U14129 ( .C1(n14969), .C2(n14838), .A(n11661), .B(n11660), .ZN(
        P1_U3278) );
  INV_X1 U14130 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n15089) );
  NOR2_X1 U14131 ( .A1(n15089), .A2(n11662), .ZN(n11749) );
  AOI21_X1 U14132 ( .B1(n11662), .B2(n15089), .A(n11749), .ZN(n11681) );
  INV_X1 U14133 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11667) );
  AOI21_X1 U14134 ( .B1(n11668), .B2(n11667), .A(n11753), .ZN(n11678) );
  MUX2_X1 U14135 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6587), .Z(n11765) );
  XOR2_X1 U14136 ( .A(n11764), .B(n11765), .Z(n11674) );
  OR2_X1 U14137 ( .A1(n11670), .A2(n11669), .ZN(n11672) );
  OAI21_X1 U14138 ( .B1(n11674), .B2(n11673), .A(n11763), .ZN(n11675) );
  NAND2_X1 U14139 ( .A1(n11675), .A2(n15422), .ZN(n11677) );
  AND2_X1 U14140 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12847) );
  AOI21_X1 U14141 ( .B1(n15417), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12847), 
        .ZN(n11676) );
  OAI211_X1 U14142 ( .C1(n11678), .C2(n15408), .A(n11677), .B(n11676), .ZN(
        n11679) );
  AOI21_X1 U14143 ( .B1(n7041), .B2(n15421), .A(n11679), .ZN(n11680) );
  OAI21_X1 U14144 ( .B1(n11681), .B2(n15407), .A(n11680), .ZN(P3_U3193) );
  INV_X1 U14145 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n11699) );
  NAND2_X1 U14146 ( .A1(n11831), .A2(n11682), .ZN(n11683) );
  NAND2_X1 U14147 ( .A1(n11684), .A2(n11683), .ZN(n11685) );
  INV_X1 U14148 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14943) );
  XNOR2_X1 U14149 ( .A(n11685), .B(n14943), .ZN(n11693) );
  NAND2_X1 U14150 ( .A1(n11831), .A2(n11686), .ZN(n11687) );
  NAND2_X1 U14151 ( .A1(n11688), .A2(n11687), .ZN(n11689) );
  XOR2_X1 U14152 ( .A(n11689), .B(P1_REG2_REG_19__SCAN_IN), .Z(n11694) );
  INV_X1 U14153 ( .A(n11694), .ZN(n11690) );
  NAND2_X1 U14154 ( .A1(n11690), .A2(n14576), .ZN(n11691) );
  OAI211_X1 U14155 ( .C1(n11693), .C2(n15208), .A(n11691), .B(n15212), .ZN(
        n11692) );
  INV_X1 U14156 ( .A(n11692), .ZN(n11697) );
  AOI22_X1 U14157 ( .A1(n11694), .A2(n14576), .B1(n11693), .B2(n14565), .ZN(
        n11696) );
  MUX2_X1 U14158 ( .A(n11697), .B(n11696), .S(n11695), .Z(n11698) );
  NAND2_X1 U14159 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14343)
         );
  OAI211_X1 U14160 ( .C1(n11699), .C2(n15216), .A(n11698), .B(n14343), .ZN(
        P1_U3262) );
  OR2_X1 U14161 ( .A1(n11700), .A2(n11703), .ZN(n11701) );
  NAND2_X1 U14162 ( .A1(n11702), .A2(n11701), .ZN(n14243) );
  XNOR2_X1 U14163 ( .A(n11704), .B(n11703), .ZN(n11705) );
  NAND2_X1 U14164 ( .A1(n11705), .A2(n6580), .ZN(n11707) );
  AOI22_X1 U14165 ( .A1(n13900), .A2(n14027), .B1(n14025), .B2(n13902), .ZN(
        n11706) );
  NAND2_X1 U14166 ( .A1(n11707), .A2(n11706), .ZN(n14244) );
  NAND2_X1 U14167 ( .A1(n14244), .A2(n14163), .ZN(n11715) );
  AOI21_X1 U14168 ( .B1(n11708), .B2(n14293), .A(n13997), .ZN(n11709) );
  AND2_X1 U14169 ( .A1(n11709), .A2(n6631), .ZN(n14245) );
  NAND2_X1 U14170 ( .A1(n14293), .A2(n15132), .ZN(n11712) );
  INV_X1 U14171 ( .A(n11710), .ZN(n13844) );
  AOI22_X1 U14172 ( .A1(n8990), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13844), 
        .B2(n15329), .ZN(n11711) );
  NAND2_X1 U14173 ( .A1(n11712), .A2(n11711), .ZN(n11713) );
  AOI21_X1 U14174 ( .B1(n14245), .B2(n6581), .A(n11713), .ZN(n11714) );
  OAI211_X1 U14175 ( .C1(n14243), .C2(n14137), .A(n11715), .B(n11714), .ZN(
        P2_U3248) );
  INV_X1 U14176 ( .A(n11716), .ZN(n11717) );
  OAI222_X1 U14177 ( .A1(n11718), .A2(P3_U3151), .B1(n12609), .B2(n13511), 
        .C1(n13756), .C2(n11717), .ZN(P3_U3269) );
  INV_X1 U14178 ( .A(n11902), .ZN(n11720) );
  OAI222_X1 U14179 ( .A1(P1_U3086), .A2(n9397), .B1(n15030), .B2(n11720), .C1(
        n11903), .C2(n15024), .ZN(P1_U3331) );
  OAI222_X1 U14180 ( .A1(n14312), .A2(n11721), .B1(n10596), .B2(n11720), .C1(
        n11719), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U14181 ( .A(n11915), .ZN(n11724) );
  OAI222_X1 U14182 ( .A1(n14312), .A2(n11723), .B1(n10596), .B2(n11724), .C1(
        n11722), .C2(P2_U3088), .ZN(P2_U3302) );
  OAI222_X1 U14183 ( .A1(P1_U3086), .A2(n11725), .B1(n15030), .B2(n11724), 
        .C1(n13373), .C2(n15024), .ZN(P1_U3330) );
  NAND2_X1 U14184 ( .A1(n11746), .A2(n12708), .ZN(n11727) );
  NAND2_X1 U14185 ( .A1(n10103), .A2(n14463), .ZN(n11726) );
  NAND2_X1 U14186 ( .A1(n11727), .A2(n11726), .ZN(n11729) );
  XNOR2_X1 U14187 ( .A(n11729), .B(n11728), .ZN(n11733) );
  NOR2_X1 U14188 ( .A1(n6812), .A2(n11730), .ZN(n11731) );
  AOI21_X1 U14189 ( .B1(n11746), .B2(n10103), .A(n11731), .ZN(n11732) );
  NAND2_X1 U14190 ( .A1(n11733), .A2(n11732), .ZN(n12617) );
  OAI21_X1 U14191 ( .B1(n11733), .B2(n11732), .A(n12617), .ZN(n11740) );
  AOI21_X1 U14192 ( .B1(n11740), .B2(n11739), .A(n11738), .ZN(n11748) );
  OAI21_X1 U14193 ( .B1(n14449), .B2(n14823), .A(n11741), .ZN(n11742) );
  AOI21_X1 U14194 ( .B1(n14447), .B2(n14464), .A(n11742), .ZN(n11743) );
  OAI21_X1 U14195 ( .B1(n11744), .B2(n14441), .A(n11743), .ZN(n11745) );
  AOI21_X1 U14196 ( .B1(n11746), .B2(n9832), .A(n11745), .ZN(n11747) );
  OAI21_X1 U14197 ( .B1(n11748), .B2(n14456), .A(n11747), .ZN(P1_U3215) );
  NOR2_X1 U14198 ( .A1(n6653), .A2(n11749), .ZN(n11752) );
  NAND2_X1 U14199 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n12898), .ZN(n11750) );
  OAI21_X1 U14200 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n12898), .A(n11750), 
        .ZN(n11751) );
  AOI21_X1 U14201 ( .B1(n11752), .B2(n11751), .A(n12900), .ZN(n11772) );
  NAND2_X1 U14202 ( .A1(n12898), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12910) );
  OAI21_X1 U14203 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n12898), .A(n12910), 
        .ZN(n11756) );
  AOI21_X1 U14204 ( .B1(n11756), .B2(n11755), .A(n12909), .ZN(n11758) );
  NOR2_X1 U14205 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13347), .ZN(n12790) );
  AOI21_X1 U14206 ( .B1(n15417), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12790), 
        .ZN(n11757) );
  OAI21_X1 U14207 ( .B1(n15408), .B2(n11758), .A(n11757), .ZN(n11769) );
  INV_X1 U14208 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11759) );
  NOR2_X1 U14209 ( .A1(n6587), .A2(n11759), .ZN(n11760) );
  AOI21_X1 U14210 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n6587), .A(n11760), .ZN(
        n11761) );
  NOR2_X1 U14211 ( .A1(n11761), .A2(n11770), .ZN(n12906) );
  AOI21_X1 U14212 ( .B1(n11761), .B2(n11770), .A(n12906), .ZN(n11762) );
  INV_X1 U14213 ( .A(n11762), .ZN(n11767) );
  AOI211_X1 U14214 ( .C1(n11767), .C2(n11766), .A(n15406), .B(n12905), .ZN(
        n11768) );
  AOI211_X1 U14215 ( .C1(n15421), .C2(n11770), .A(n11769), .B(n11768), .ZN(
        n11771) );
  OAI21_X1 U14216 ( .B1(n11772), .B2(n15407), .A(n11771), .ZN(P3_U3194) );
  INV_X1 U14217 ( .A(n12447), .ZN(n15022) );
  OAI222_X1 U14218 ( .A1(n10596), .A2(n15022), .B1(n11773), .B2(P2_U3088), 
        .C1(n12020), .C2(n14312), .ZN(P2_U3298) );
  INV_X1 U14219 ( .A(n11941), .ZN(n15026) );
  OAI222_X1 U14220 ( .A1(n10596), .A2(n15026), .B1(n8980), .B2(P2_U3088), .C1(
        n11774), .C2(n14312), .ZN(P2_U3300) );
  NOR2_X1 U14221 ( .A1(n15310), .A2(n11777), .ZN(n11778) );
  AOI21_X1 U14222 ( .B1(n11777), .B2(n15310), .A(n11778), .ZN(n15321) );
  NAND2_X1 U14223 ( .A1(n15322), .A2(n15321), .ZN(n15320) );
  OAI21_X1 U14224 ( .B1(n11777), .B2(n15310), .A(n15320), .ZN(n11779) );
  NOR2_X1 U14225 ( .A1(n11779), .A2(n13952), .ZN(n11780) );
  INV_X1 U14226 ( .A(n11794), .ZN(n11792) );
  AOI22_X1 U14227 ( .A1(n11783), .A2(n11782), .B1(n11781), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n15315) );
  XNOR2_X1 U14228 ( .A(n11784), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15316) );
  INV_X1 U14229 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11785) );
  OAI22_X1 U14230 ( .A1(n15315), .A2(n15316), .B1(n11785), .B2(n15310), .ZN(
        n11787) );
  XNOR2_X1 U14231 ( .A(n11787), .B(n13952), .ZN(n13951) );
  OR2_X1 U14232 ( .A1(n13951), .A2(n11786), .ZN(n11789) );
  NAND2_X1 U14233 ( .A1(n11787), .A2(n13952), .ZN(n11788) );
  NAND2_X1 U14234 ( .A1(n11789), .A2(n11788), .ZN(n11790) );
  XNOR2_X1 U14235 ( .A(n11790), .B(n13336), .ZN(n11793) );
  NOR2_X1 U14236 ( .A1(n11793), .A2(n15269), .ZN(n11791) );
  AOI22_X1 U14237 ( .A1(n11794), .A2(n15319), .B1(n15317), .B2(n11793), .ZN(
        n11796) );
  NAND2_X1 U14238 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13785)
         );
  OAI211_X1 U14239 ( .C1(n11799), .C2(n11798), .A(n11797), .B(n13785), .ZN(
        P2_U3233) );
  OAI22_X1 U14240 ( .A1(n13817), .A2(n11801), .B1(n9906), .B2(n13872), .ZN(
        n11804) );
  INV_X1 U14241 ( .A(n11802), .ZN(n11803) );
  NAND3_X1 U14242 ( .A1(n11804), .A2(n11803), .A3(n10131), .ZN(n11809) );
  INV_X1 U14243 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n13514) );
  OAI22_X1 U14244 ( .A1(n11806), .A2(n13514), .B1(n13853), .B2(n11805), .ZN(
        n11807) );
  AOI21_X1 U14245 ( .B1(n14158), .B2(n15107), .A(n11807), .ZN(n11808) );
  OAI211_X1 U14246 ( .C1(n11800), .C2(n13872), .A(n11809), .B(n11808), .ZN(
        P2_U3209) );
  NAND2_X1 U14247 ( .A1(n14307), .A2(n12456), .ZN(n11811) );
  OR2_X1 U14248 ( .A1(n12458), .A2(n11999), .ZN(n11810) );
  OR2_X1 U14249 ( .A1(n14967), .A2(n14462), .ZN(n11813) );
  AOI22_X1 U14250 ( .A1(n11845), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11844), 
        .B2(n11815), .ZN(n11816) );
  XNOR2_X1 U14251 ( .A(n14830), .B(n14461), .ZN(n12507) );
  OR2_X1 U14252 ( .A1(n14830), .A2(n14461), .ZN(n11818) );
  NAND2_X1 U14253 ( .A1(n11819), .A2(n12456), .ZN(n11822) );
  AOI22_X1 U14254 ( .A1(n11845), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11844), 
        .B2(n11820), .ZN(n11821) );
  NAND2_X2 U14255 ( .A1(n11822), .A2(n11821), .ZN(n14954) );
  NOR2_X1 U14256 ( .A1(n11823), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11824) );
  OR2_X1 U14257 ( .A1(n11834), .A2(n11824), .ZN(n14811) );
  AOI22_X1 U14258 ( .A1(n11985), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n12450), 
        .B2(P1_REG0_REG_17__SCAN_IN), .ZN(n11826) );
  OR2_X1 U14259 ( .A1(n12454), .A2(n13374), .ZN(n11825) );
  OAI211_X1 U14260 ( .C1(n14811), .C2(n11986), .A(n11826), .B(n11825), .ZN(
        n14790) );
  NAND2_X1 U14261 ( .A1(n14954), .A2(n14790), .ZN(n11827) );
  OR2_X1 U14262 ( .A1(n14954), .A2(n14790), .ZN(n11828) );
  NAND2_X1 U14263 ( .A1(n11830), .A2(n12456), .ZN(n11833) );
  AOI22_X1 U14264 ( .A1(n11845), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11844), 
        .B2(n11831), .ZN(n11832) );
  NAND2_X2 U14265 ( .A1(n11833), .A2(n11832), .ZN(n14786) );
  NAND2_X1 U14266 ( .A1(n11834), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11849) );
  OR2_X1 U14267 ( .A1(n11834), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11835) );
  AND2_X1 U14268 ( .A1(n11849), .A2(n11835), .ZN(n14778) );
  NAND2_X1 U14269 ( .A1(n14778), .A2(n11878), .ZN(n11840) );
  INV_X1 U14270 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14950) );
  NAND2_X1 U14271 ( .A1(n12450), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11837) );
  INV_X1 U14272 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14780) );
  OR2_X1 U14273 ( .A1(n12289), .A2(n14780), .ZN(n11836) );
  OAI211_X1 U14274 ( .C1(n12454), .C2(n14950), .A(n11837), .B(n11836), .ZN(
        n11838) );
  INV_X1 U14275 ( .A(n11838), .ZN(n11839) );
  NAND2_X1 U14276 ( .A1(n11840), .A2(n11839), .ZN(n14802) );
  NOR2_X1 U14277 ( .A1(n14786), .A2(n14802), .ZN(n11842) );
  NAND2_X1 U14278 ( .A1(n14786), .A2(n14802), .ZN(n11841) );
  NAND2_X1 U14279 ( .A1(n11843), .A2(n12456), .ZN(n11847) );
  AOI22_X1 U14280 ( .A1(n11845), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14768), 
        .B2(n11844), .ZN(n11846) );
  INV_X1 U14281 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n11848) );
  NAND2_X1 U14282 ( .A1(n11849), .A2(n11848), .ZN(n11850) );
  AND2_X1 U14283 ( .A1(n11861), .A2(n11850), .ZN(n14770) );
  NAND2_X1 U14284 ( .A1(n14770), .A2(n11878), .ZN(n11855) );
  NAND2_X1 U14285 ( .A1(n11985), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n11852) );
  NAND2_X1 U14286 ( .A1(n12450), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11851) );
  OAI211_X1 U14287 ( .C1(n14943), .C2(n12454), .A(n11852), .B(n11851), .ZN(
        n11853) );
  INV_X1 U14288 ( .A(n11853), .ZN(n11854) );
  NAND2_X1 U14289 ( .A1(n11855), .A2(n11854), .ZN(n14792) );
  OR2_X1 U14290 ( .A1(n14765), .A2(n14792), .ZN(n11856) );
  NAND2_X1 U14291 ( .A1(n11858), .A2(n12456), .ZN(n11860) );
  OR2_X1 U14292 ( .A1(n12458), .A2(n13338), .ZN(n11859) );
  INV_X1 U14293 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14401) );
  AND2_X1 U14294 ( .A1(n11861), .A2(n14401), .ZN(n11862) );
  NOR2_X1 U14295 ( .A1(n11862), .A2(n11872), .ZN(n14755) );
  INV_X1 U14296 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14933) );
  NAND2_X1 U14297 ( .A1(n11985), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11864) );
  NAND2_X1 U14298 ( .A1(n12450), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11863) );
  OAI211_X1 U14299 ( .C1(n14933), .C2(n12454), .A(n11864), .B(n11863), .ZN(
        n11865) );
  AOI21_X1 U14300 ( .B1(n14755), .B2(n11878), .A(n11865), .ZN(n14352) );
  INV_X1 U14301 ( .A(n14352), .ZN(n14460) );
  NAND2_X1 U14302 ( .A1(n14999), .A2(n14460), .ZN(n11970) );
  OR2_X1 U14303 ( .A1(n14999), .A2(n14460), .ZN(n11866) );
  NAND2_X1 U14304 ( .A1(n11970), .A2(n11866), .ZN(n12511) );
  INV_X1 U14305 ( .A(n12511), .ZN(n14752) );
  OR2_X1 U14306 ( .A1(n14999), .A2(n14352), .ZN(n11867) );
  NAND2_X1 U14307 ( .A1(n11868), .A2(n12456), .ZN(n11871) );
  OR2_X1 U14308 ( .A1(n12458), .A2(n11869), .ZN(n11870) );
  OR2_X1 U14309 ( .A1(n11872), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11873) );
  NAND2_X1 U14310 ( .A1(n11872), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11882) );
  AND2_X1 U14311 ( .A1(n11873), .A2(n11882), .ZN(n14738) );
  INV_X1 U14312 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n14740) );
  NAND2_X1 U14313 ( .A1(n11874), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n11876) );
  NAND2_X1 U14314 ( .A1(n12450), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11875) );
  OAI211_X1 U14315 ( .C1(n12289), .C2(n14740), .A(n11876), .B(n11875), .ZN(
        n11877) );
  AOI21_X1 U14316 ( .B1(n14738), .B2(n11878), .A(n11877), .ZN(n14398) );
  XNOR2_X1 U14317 ( .A(n14925), .B(n14398), .ZN(n14734) );
  NAND2_X1 U14318 ( .A1(n14925), .A2(n14398), .ZN(n11879) );
  NAND2_X1 U14319 ( .A1(n11880), .A2(n11879), .ZN(n14722) );
  OR2_X1 U14320 ( .A1(n8804), .A2(n7274), .ZN(n11881) );
  XNOR2_X1 U14321 ( .A(n11881), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15033) );
  NAND2_X1 U14322 ( .A1(n12450), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11887) );
  INV_X1 U14323 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14725) );
  OR2_X1 U14324 ( .A1(n12289), .A2(n14725), .ZN(n11886) );
  NAND2_X1 U14325 ( .A1(n11883), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11894) );
  OAI21_X1 U14326 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n11883), .A(n11894), 
        .ZN(n14726) );
  OR2_X1 U14327 ( .A1(n11986), .A2(n14726), .ZN(n11885) );
  INV_X1 U14328 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n13352) );
  OR2_X1 U14329 ( .A1(n12454), .A2(n13352), .ZN(n11884) );
  XNOR2_X1 U14330 ( .A(n14917), .B(n14351), .ZN(n14718) );
  INV_X1 U14331 ( .A(n14718), .ZN(n14723) );
  NAND2_X1 U14332 ( .A1(n14722), .A2(n14723), .ZN(n14721) );
  NAND2_X1 U14333 ( .A1(n14917), .A2(n14351), .ZN(n11888) );
  NAND2_X1 U14334 ( .A1(n11889), .A2(n12456), .ZN(n11892) );
  OR2_X1 U14335 ( .A1(n12458), .A2(n11890), .ZN(n11891) );
  NAND2_X1 U14336 ( .A1(n11985), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11900) );
  INV_X1 U14337 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n11893) );
  OR2_X1 U14338 ( .A1(n11944), .A2(n11893), .ZN(n11899) );
  INV_X1 U14339 ( .A(n11906), .ZN(n11908) );
  OAI21_X1 U14340 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n11895), .A(n11908), 
        .ZN(n14701) );
  OR2_X1 U14341 ( .A1(n11986), .A2(n14701), .ZN(n11898) );
  INV_X1 U14342 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n11896) );
  OR2_X1 U14343 ( .A1(n12454), .A2(n11896), .ZN(n11897) );
  NAND4_X1 U14344 ( .A1(n11900), .A2(n11899), .A3(n11898), .A4(n11897), .ZN(
        n14685) );
  XNOR2_X1 U14345 ( .A(n14909), .B(n14685), .ZN(n14708) );
  OR2_X2 U14346 ( .A1(n14698), .A2(n14708), .ZN(n14700) );
  NAND2_X1 U14347 ( .A1(n14909), .A2(n14685), .ZN(n11901) );
  NAND2_X1 U14348 ( .A1(n11902), .A2(n12456), .ZN(n11905) );
  OR2_X1 U14349 ( .A1(n12458), .A2(n11903), .ZN(n11904) );
  NAND2_X1 U14350 ( .A1(n11985), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11913) );
  INV_X1 U14351 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14991) );
  OR2_X1 U14352 ( .A1(n11944), .A2(n14991), .ZN(n11912) );
  INV_X1 U14353 ( .A(n11919), .ZN(n11921) );
  INV_X1 U14354 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n11907) );
  NAND2_X1 U14355 ( .A1(n11908), .A2(n11907), .ZN(n11909) );
  NAND2_X1 U14356 ( .A1(n11921), .A2(n11909), .ZN(n14692) );
  OR2_X1 U14357 ( .A1(n11986), .A2(n14692), .ZN(n11911) );
  INV_X1 U14358 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14906) );
  OR2_X1 U14359 ( .A1(n12454), .A2(n14906), .ZN(n11910) );
  NAND4_X1 U14360 ( .A1(n11913), .A2(n11912), .A3(n11911), .A4(n11910), .ZN(
        n14711) );
  INV_X1 U14361 ( .A(n14711), .ZN(n11974) );
  XNOR2_X1 U14362 ( .A(n14691), .B(n11974), .ZN(n12514) );
  OR2_X1 U14363 ( .A1(n14691), .A2(n14711), .ZN(n11914) );
  NAND2_X1 U14364 ( .A1(n11915), .A2(n12456), .ZN(n11917) );
  OR2_X1 U14365 ( .A1(n12458), .A2(n13373), .ZN(n11916) );
  NAND2_X1 U14366 ( .A1(n11985), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11928) );
  INV_X1 U14367 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n11918) );
  OR2_X1 U14368 ( .A1(n11944), .A2(n11918), .ZN(n11927) );
  INV_X1 U14369 ( .A(n11932), .ZN(n11923) );
  INV_X1 U14370 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n11920) );
  NAND2_X1 U14371 ( .A1(n11921), .A2(n11920), .ZN(n11922) );
  NAND2_X1 U14372 ( .A1(n11923), .A2(n11922), .ZN(n14671) );
  OR2_X1 U14373 ( .A1(n11986), .A2(n14671), .ZN(n11926) );
  INV_X1 U14374 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n11924) );
  OR2_X1 U14375 ( .A1(n12454), .A2(n11924), .ZN(n11925) );
  NAND4_X1 U14376 ( .A1(n11928), .A2(n11927), .A3(n11926), .A4(n11925), .ZN(
        n14684) );
  XNOR2_X1 U14377 ( .A(n14987), .B(n14684), .ZN(n12515) );
  NAND2_X1 U14378 ( .A1(n14987), .A2(n14684), .ZN(n11929) );
  NAND2_X1 U14379 ( .A1(n14666), .A2(n11929), .ZN(n14650) );
  NAND2_X1 U14380 ( .A1(n14311), .A2(n12456), .ZN(n11931) );
  OR2_X1 U14381 ( .A1(n12458), .A2(n15028), .ZN(n11930) );
  NAND2_X1 U14382 ( .A1(n11985), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11937) );
  INV_X1 U14383 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n13457) );
  OR2_X1 U14384 ( .A1(n11944), .A2(n13457), .ZN(n11936) );
  NAND2_X1 U14385 ( .A1(n11932), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11945) );
  OAI21_X1 U14386 ( .B1(n11932), .B2(P1_REG3_REG_26__SCAN_IN), .A(n11945), 
        .ZN(n14661) );
  OR2_X1 U14387 ( .A1(n11986), .A2(n14661), .ZN(n11935) );
  INV_X1 U14388 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n11933) );
  OR2_X1 U14389 ( .A1(n12454), .A2(n11933), .ZN(n11934) );
  NAND4_X1 U14390 ( .A1(n11937), .A2(n11936), .A3(n11935), .A4(n11934), .ZN(
        n14633) );
  INV_X1 U14391 ( .A(n14633), .ZN(n11938) );
  NAND2_X1 U14392 ( .A1(n14887), .A2(n11938), .ZN(n11979) );
  OR2_X1 U14393 ( .A1(n14887), .A2(n11938), .ZN(n11939) );
  NAND2_X1 U14394 ( .A1(n11979), .A2(n11939), .ZN(n14649) );
  AND2_X1 U14395 ( .A1(n14887), .A2(n14633), .ZN(n11940) );
  NAND2_X1 U14396 ( .A1(n11941), .A2(n12456), .ZN(n11943) );
  OR2_X1 U14397 ( .A1(n12458), .A2(n15025), .ZN(n11942) );
  NAND2_X1 U14398 ( .A1(n11985), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n11950) );
  INV_X1 U14399 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14982) );
  OR2_X1 U14400 ( .A1(n11944), .A2(n14982), .ZN(n11949) );
  INV_X1 U14401 ( .A(n11945), .ZN(n11946) );
  NAND2_X1 U14402 ( .A1(n11946), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11953) );
  OAI21_X1 U14403 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n11946), .A(n11953), 
        .ZN(n14642) );
  OR2_X1 U14404 ( .A1(n11986), .A2(n14642), .ZN(n11948) );
  INV_X1 U14405 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n14885) );
  OR2_X1 U14406 ( .A1(n12454), .A2(n14885), .ZN(n11947) );
  NAND4_X1 U14407 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n14656) );
  XNOR2_X1 U14408 ( .A(n14878), .B(n14656), .ZN(n14631) );
  INV_X1 U14409 ( .A(n14631), .ZN(n14625) );
  OR2_X1 U14410 ( .A1(n14878), .A2(n14656), .ZN(n11951) );
  NAND2_X1 U14411 ( .A1(n12450), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11959) );
  INV_X1 U14412 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n11952) );
  OR2_X1 U14413 ( .A1(n12454), .A2(n11952), .ZN(n11958) );
  INV_X1 U14414 ( .A(n11953), .ZN(n11954) );
  NAND2_X1 U14415 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n11954), .ZN(n14606) );
  OAI21_X1 U14416 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(n11954), .A(n14606), 
        .ZN(n14617) );
  OR2_X1 U14417 ( .A1(n11986), .A2(n14617), .ZN(n11957) );
  INV_X1 U14418 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n11955) );
  OR2_X1 U14419 ( .A1(n12289), .A2(n11955), .ZN(n11956) );
  NAND4_X1 U14420 ( .A1(n11959), .A2(n11958), .A3(n11957), .A4(n11956), .ZN(
        n14634) );
  INV_X1 U14421 ( .A(n14634), .ZN(n11960) );
  NAND2_X1 U14422 ( .A1(n14980), .A2(n11960), .ZN(n14598) );
  OR2_X1 U14423 ( .A1(n14980), .A2(n11960), .ZN(n11961) );
  OR2_X1 U14424 ( .A1(n14596), .A2(n11962), .ZN(n14615) );
  NAND2_X1 U14425 ( .A1(n11964), .A2(n11963), .ZN(n11965) );
  NAND2_X1 U14426 ( .A1(n14830), .A2(n14805), .ZN(n11966) );
  INV_X1 U14427 ( .A(n14790), .ZN(n14825) );
  XNOR2_X1 U14428 ( .A(n14954), .B(n14825), .ZN(n12394) );
  INV_X1 U14429 ( .A(n12394), .ZN(n14799) );
  OR2_X1 U14430 ( .A1(n14954), .A2(n14825), .ZN(n12393) );
  INV_X1 U14431 ( .A(n14802), .ZN(n14383) );
  NOR2_X1 U14432 ( .A1(n14786), .A2(n14383), .ZN(n11967) );
  INV_X1 U14433 ( .A(n14792), .ZN(n14421) );
  NAND2_X1 U14434 ( .A1(n14765), .A2(n14421), .ZN(n11968) );
  INV_X1 U14435 ( .A(n14398), .ZN(n14459) );
  NAND2_X1 U14436 ( .A1(n14719), .A2(n14718), .ZN(n14717) );
  INV_X1 U14437 ( .A(n14351), .ZN(n14712) );
  OR2_X1 U14438 ( .A1(n14917), .A2(n14712), .ZN(n11971) );
  NAND2_X1 U14439 ( .A1(n14717), .A2(n11971), .ZN(n14709) );
  INV_X1 U14440 ( .A(n14685), .ZN(n11972) );
  NAND2_X1 U14441 ( .A1(n14909), .A2(n11972), .ZN(n11973) );
  OR2_X1 U14442 ( .A1(n14691), .A2(n11974), .ZN(n11975) );
  INV_X1 U14443 ( .A(n14684), .ZN(n11976) );
  NAND2_X1 U14444 ( .A1(n14987), .A2(n11976), .ZN(n11977) );
  INV_X1 U14445 ( .A(n14649), .ZN(n14655) );
  NAND2_X1 U14446 ( .A1(n14654), .A2(n14655), .ZN(n14653) );
  NAND2_X1 U14447 ( .A1(n14653), .A2(n11979), .ZN(n14632) );
  INV_X1 U14448 ( .A(n14656), .ZN(n11980) );
  NAND2_X1 U14449 ( .A1(n14878), .A2(n11980), .ZN(n11982) );
  NAND2_X1 U14450 ( .A1(n14630), .A2(n11982), .ZN(n11981) );
  NAND2_X1 U14451 ( .A1(n11981), .A2(n12517), .ZN(n14599) );
  INV_X1 U14452 ( .A(n12517), .ZN(n11983) );
  NAND3_X1 U14453 ( .A1(n14630), .A2(n11983), .A3(n11982), .ZN(n11984) );
  NAND2_X1 U14454 ( .A1(n14599), .A2(n11984), .ZN(n11994) );
  NAND2_X1 U14455 ( .A1(n12450), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11991) );
  NAND2_X1 U14456 ( .A1(n11985), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11990) );
  OR2_X1 U14457 ( .A1(n11986), .A2(n14606), .ZN(n11989) );
  INV_X1 U14458 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n11987) );
  OR2_X1 U14459 ( .A1(n12454), .A2(n11987), .ZN(n11988) );
  NAND4_X1 U14460 ( .A1(n11991), .A2(n11990), .A3(n11989), .A4(n11988), .ZN(
        n14458) );
  AOI22_X1 U14461 ( .A1(n14850), .A2(n14458), .B1(n14656), .B2(n14791), .ZN(
        n11992) );
  INV_X1 U14462 ( .A(n11992), .ZN(n11993) );
  INV_X1 U14463 ( .A(n14954), .ZN(n14810) );
  NAND2_X1 U14464 ( .A1(n14810), .A2(n14827), .ZN(n14807) );
  AND2_X2 U14465 ( .A1(n14753), .A2(n14925), .ZN(n14737) );
  NAND2_X1 U14466 ( .A1(n14917), .A2(n14737), .ZN(n14724) );
  NAND2_X1 U14467 ( .A1(n14980), .A2(n6633), .ZN(n11995) );
  NAND2_X1 U14468 ( .A1(n11995), .A2(n14888), .ZN(n11996) );
  OR2_X1 U14469 ( .A1(n14603), .A2(n11996), .ZN(n14620) );
  AOI21_X1 U14470 ( .B1(n14900), .B2(n14980), .A(n11997), .ZN(n11998) );
  INV_X1 U14471 ( .A(n11998), .ZN(P1_U3556) );
  INV_X1 U14472 ( .A(n14307), .ZN(n12000) );
  OAI222_X1 U14473 ( .A1(n14490), .A2(P1_U3086), .B1(n15030), .B2(n12000), 
        .C1(n11999), .C2(n15024), .ZN(P1_U3327) );
  INV_X1 U14474 ( .A(n12457), .ZN(n15019) );
  OAI222_X1 U14475 ( .A1(n10596), .A2(n15019), .B1(n12001), .B2(P2_U3088), 
        .C1(n12036), .C2(n14312), .ZN(P2_U3297) );
  OAI21_X1 U14476 ( .B1(n13888), .B2(n12003), .A(n12002), .ZN(n12008) );
  INV_X1 U14477 ( .A(n12004), .ZN(n12005) );
  OAI22_X1 U14478 ( .A1(n13883), .A2(n12006), .B1(n15111), .B2(n12005), .ZN(
        n12007) );
  AOI211_X1 U14479 ( .C1(n12009), .C2(n13913), .A(n12008), .B(n12007), .ZN(
        n12017) );
  OAI22_X1 U14480 ( .A1(n13817), .A2(n12011), .B1(n12010), .B2(n13872), .ZN(
        n12015) );
  INV_X1 U14481 ( .A(n12012), .ZN(n12014) );
  NAND3_X1 U14482 ( .A1(n12015), .A2(n12014), .A3(n12013), .ZN(n12016) );
  OAI211_X1 U14483 ( .C1(n12018), .C2(n13872), .A(n12017), .B(n12016), .ZN(
        P2_U3199) );
  NAND2_X1 U14484 ( .A1(n12020), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12021) );
  NAND2_X1 U14485 ( .A1(n12022), .A2(n12021), .ZN(n12024) );
  NAND2_X1 U14486 ( .A1(n15021), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12023) );
  NOR2_X1 U14487 ( .A1(n12036), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12025) );
  INV_X1 U14488 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n15018) );
  OAI22_X1 U14489 ( .A1(n12038), .A2(n12025), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n15018), .ZN(n12027) );
  XNOR2_X1 U14490 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n12026) );
  XNOR2_X1 U14491 ( .A(n12027), .B(n12026), .ZN(n13750) );
  INV_X1 U14492 ( .A(SI_31_), .ZN(n13745) );
  NOR2_X1 U14493 ( .A1(n12040), .A2(n13745), .ZN(n12028) );
  NAND2_X1 U14494 ( .A1(n12029), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12033) );
  NAND2_X1 U14495 ( .A1(n12030), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12032) );
  NAND2_X1 U14496 ( .A1(n7830), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12031) );
  AND3_X1 U14497 ( .A1(n12033), .A2(n12032), .A3(n12031), .ZN(n12034) );
  NAND2_X1 U14498 ( .A1(n12035), .A2(n12034), .ZN(n12886) );
  NAND2_X1 U14499 ( .A1(n13079), .A2(n12886), .ZN(n12224) );
  XNOR2_X1 U14500 ( .A(n12036), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n12037) );
  XNOR2_X1 U14501 ( .A(n12038), .B(n12037), .ZN(n12606) );
  NAND2_X1 U14502 ( .A1(n12606), .A2(n12039), .ZN(n12042) );
  INV_X1 U14503 ( .A(SI_30_), .ZN(n12608) );
  OR2_X1 U14504 ( .A1(n12040), .A2(n12608), .ZN(n12041) );
  NAND2_X1 U14505 ( .A1(n12042), .A2(n12041), .ZN(n12044) );
  NAND2_X1 U14506 ( .A1(n12044), .A2(n12047), .ZN(n12195) );
  AND3_X1 U14507 ( .A1(n12224), .A2(n12043), .A3(n12195), .ZN(n12190) );
  NAND2_X1 U14508 ( .A1(n12046), .A2(n12045), .ZN(n12050) );
  INV_X1 U14509 ( .A(n12886), .ZN(n13075) );
  NAND2_X1 U14510 ( .A1(n12048), .A2(n13075), .ZN(n12223) );
  INV_X1 U14511 ( .A(n12047), .ZN(n12887) );
  NAND2_X1 U14512 ( .A1(n12050), .A2(n7624), .ZN(n12051) );
  XNOR2_X1 U14513 ( .A(n12053), .B(n12165), .ZN(n12168) );
  INV_X1 U14514 ( .A(n13175), .ZN(n13643) );
  NAND2_X1 U14515 ( .A1(n12071), .A2(n12054), .ZN(n12057) );
  NAND2_X1 U14516 ( .A1(n12070), .A2(n12055), .ZN(n12056) );
  MUX2_X1 U14517 ( .A(n12057), .B(n12056), .S(n12165), .Z(n12080) );
  NAND2_X1 U14518 ( .A1(n12059), .A2(n12058), .ZN(n12062) );
  MUX2_X1 U14519 ( .A(n12062), .B(n12061), .S(n12060), .Z(n12066) );
  OAI21_X1 U14520 ( .B1(n12064), .B2(n12063), .A(n12183), .ZN(n12065) );
  NAND4_X1 U14521 ( .A1(n12066), .A2(n12204), .A3(n12068), .A4(n12065), .ZN(
        n12079) );
  AOI21_X1 U14522 ( .B1(n12067), .B2(n12069), .A(n12080), .ZN(n12077) );
  MUX2_X1 U14523 ( .A(n12071), .B(n12070), .S(n12183), .Z(n12072) );
  NAND2_X1 U14524 ( .A1(n12204), .A2(n12072), .ZN(n12076) );
  MUX2_X1 U14525 ( .A(n12074), .B(n12073), .S(n12165), .Z(n12075) );
  OAI21_X1 U14526 ( .B1(n12077), .B2(n12076), .A(n12075), .ZN(n12078) );
  OAI21_X1 U14527 ( .B1(n12080), .B2(n12079), .A(n12078), .ZN(n12086) );
  NAND2_X1 U14528 ( .A1(n12088), .A2(n12081), .ZN(n12084) );
  NAND2_X1 U14529 ( .A1(n12087), .A2(n12082), .ZN(n12083) );
  MUX2_X1 U14530 ( .A(n12084), .B(n12083), .S(n12183), .Z(n12085) );
  AOI21_X1 U14531 ( .B1(n12086), .B2(n12202), .A(n12085), .ZN(n12094) );
  MUX2_X1 U14532 ( .A(n12088), .B(n12087), .S(n12165), .Z(n12089) );
  NAND2_X1 U14533 ( .A1(n12089), .A2(n12207), .ZN(n12093) );
  XNOR2_X1 U14534 ( .A(n12894), .B(n15453), .ZN(n15449) );
  NAND2_X1 U14535 ( .A1(n15460), .A2(n15560), .ZN(n12091) );
  MUX2_X1 U14536 ( .A(n12091), .B(n12090), .S(n12183), .Z(n12092) );
  OAI211_X1 U14537 ( .C1(n12094), .C2(n12093), .A(n15449), .B(n12092), .ZN(
        n12098) );
  MUX2_X1 U14538 ( .A(n12096), .B(n12095), .S(n12165), .Z(n12097) );
  NAND3_X1 U14539 ( .A1(n12098), .A2(n12203), .A3(n12097), .ZN(n12102) );
  MUX2_X1 U14540 ( .A(n12100), .B(n12099), .S(n12183), .Z(n12101) );
  NAND3_X1 U14541 ( .A1(n12102), .A2(n15439), .A3(n12101), .ZN(n12106) );
  NAND2_X1 U14542 ( .A1(n12892), .A2(n15443), .ZN(n12104) );
  MUX2_X1 U14543 ( .A(n12104), .B(n12103), .S(n12165), .Z(n12105) );
  AOI21_X1 U14544 ( .B1(n12106), .B2(n12105), .A(n7011), .ZN(n12109) );
  AOI21_X1 U14545 ( .B1(n12112), .B2(n12107), .A(n12183), .ZN(n12108) );
  OAI21_X1 U14546 ( .B1(n12109), .B2(n12108), .A(n12110), .ZN(n12115) );
  OAI21_X1 U14547 ( .B1(n15435), .B2(n15085), .A(n12110), .ZN(n12111) );
  NAND2_X1 U14548 ( .A1(n12111), .A2(n12183), .ZN(n12114) );
  INV_X1 U14549 ( .A(n12112), .ZN(n12113) );
  AOI22_X1 U14550 ( .A1(n12115), .A2(n12114), .B1(n12183), .B2(n12113), .ZN(
        n12120) );
  MUX2_X1 U14551 ( .A(n12118), .B(n12117), .S(n12183), .Z(n12119) );
  OAI211_X1 U14552 ( .C1(n12120), .C2(n8272), .A(n8005), .B(n12119), .ZN(
        n12124) );
  INV_X1 U14553 ( .A(n6828), .ZN(n15074) );
  NAND2_X1 U14554 ( .A1(n15074), .A2(n12833), .ZN(n12121) );
  MUX2_X1 U14555 ( .A(n12122), .B(n12121), .S(n12183), .Z(n12123) );
  NAND3_X1 U14556 ( .A1(n12124), .A2(n13558), .A3(n12123), .ZN(n12129) );
  OAI21_X1 U14557 ( .B1(n13676), .B2(n13560), .A(n12125), .ZN(n12126) );
  NAND2_X1 U14558 ( .A1(n12126), .A2(n12165), .ZN(n12128) );
  INV_X1 U14559 ( .A(n12131), .ZN(n12127) );
  AOI21_X1 U14560 ( .B1(n12129), .B2(n12128), .A(n12127), .ZN(n12134) );
  AOI21_X1 U14561 ( .B1(n12131), .B2(n12130), .A(n12165), .ZN(n12133) );
  NAND2_X1 U14562 ( .A1(n13246), .A2(n12183), .ZN(n12132) );
  OAI22_X1 U14563 ( .A1(n12134), .A2(n12133), .B1(n13676), .B2(n12132), .ZN(
        n12141) );
  INV_X1 U14564 ( .A(n12135), .ZN(n12140) );
  NAND2_X1 U14565 ( .A1(n13729), .A2(n13212), .ZN(n12148) );
  INV_X1 U14566 ( .A(n12136), .ZN(n12137) );
  NAND2_X1 U14567 ( .A1(n12142), .A2(n12137), .ZN(n12138) );
  NAND4_X1 U14568 ( .A1(n12148), .A2(n12183), .A3(n12139), .A4(n12138), .ZN(
        n12143) );
  AOI22_X1 U14569 ( .A1(n12141), .A2(n13254), .B1(n12140), .B2(n12143), .ZN(
        n12146) );
  AND3_X1 U14570 ( .A1(n12147), .A2(n12165), .A3(n12142), .ZN(n12145) );
  INV_X1 U14571 ( .A(n12143), .ZN(n12144) );
  OAI22_X1 U14572 ( .A1(n12146), .A2(n8282), .B1(n12145), .B2(n12144), .ZN(
        n12150) );
  MUX2_X1 U14573 ( .A(n12148), .B(n12147), .S(n12183), .Z(n12149) );
  NAND3_X1 U14574 ( .A1(n12150), .A2(n13207), .A3(n12149), .ZN(n12154) );
  XNOR2_X1 U14575 ( .A(n13198), .B(n13211), .ZN(n12197) );
  INV_X1 U14576 ( .A(n12889), .ZN(n13223) );
  NAND2_X1 U14577 ( .A1(n12271), .A2(n13223), .ZN(n12152) );
  MUX2_X1 U14578 ( .A(n12152), .B(n12151), .S(n12183), .Z(n12153) );
  NAND3_X1 U14579 ( .A1(n12154), .A2(n12197), .A3(n12153), .ZN(n12158) );
  AND2_X1 U14580 ( .A1(n12160), .A2(n12159), .ZN(n12196) );
  MUX2_X1 U14581 ( .A(n12156), .B(n12155), .S(n12165), .Z(n12157) );
  AND3_X1 U14582 ( .A1(n12158), .A2(n12196), .A3(n12157), .ZN(n12164) );
  INV_X1 U14583 ( .A(n12159), .ZN(n12162) );
  INV_X1 U14584 ( .A(n12160), .ZN(n12161) );
  MUX2_X1 U14585 ( .A(n12162), .B(n12161), .S(n12183), .Z(n12163) );
  OAI33_X1 U14586 ( .A1(n13151), .A2(n13643), .A3(n12165), .B1(n13168), .B2(
        n12164), .B3(n12163), .ZN(n12166) );
  AOI21_X1 U14587 ( .B1(n12166), .B2(n13147), .A(n13135), .ZN(n12167) );
  OAI21_X1 U14588 ( .B1(n13146), .B2(n12168), .A(n12167), .ZN(n12173) );
  INV_X1 U14589 ( .A(n13127), .ZN(n12172) );
  NAND3_X1 U14590 ( .A1(n12173), .A2(n12172), .A3(n12169), .ZN(n12170) );
  NAND2_X1 U14591 ( .A1(n12170), .A2(n13103), .ZN(n12177) );
  NAND3_X1 U14592 ( .A1(n12173), .A2(n12172), .A3(n12171), .ZN(n12175) );
  NAND2_X1 U14593 ( .A1(n12175), .A2(n12174), .ZN(n12176) );
  NAND2_X1 U14594 ( .A1(n12178), .A2(n13102), .ZN(n12182) );
  AOI21_X1 U14595 ( .B1(n12182), .B2(n12179), .A(n13090), .ZN(n12185) );
  AND3_X1 U14596 ( .A1(n12182), .A2(n12181), .A3(n12180), .ZN(n12184) );
  INV_X1 U14597 ( .A(n12186), .ZN(n12188) );
  INV_X1 U14598 ( .A(n12190), .ZN(n12193) );
  INV_X1 U14599 ( .A(n12223), .ZN(n12191) );
  OAI21_X1 U14600 ( .B1(n12191), .B2(n7637), .A(n12224), .ZN(n12192) );
  OAI21_X1 U14601 ( .B1(n12194), .B2(n12193), .A(n12192), .ZN(n12229) );
  INV_X1 U14602 ( .A(n12195), .ZN(n12222) );
  INV_X1 U14603 ( .A(n13259), .ZN(n13258) );
  INV_X1 U14604 ( .A(n10359), .ZN(n12198) );
  NAND4_X1 U14605 ( .A1(n12201), .A2(n12200), .A3(n12199), .A4(n12198), .ZN(
        n12206) );
  NAND4_X1 U14606 ( .A1(n12067), .A2(n12204), .A3(n12203), .A4(n12202), .ZN(
        n12205) );
  NOR2_X1 U14607 ( .A1(n12206), .A2(n12205), .ZN(n12210) );
  AND3_X1 U14608 ( .A1(n15068), .A2(n12207), .A3(n15439), .ZN(n12209) );
  NAND4_X1 U14609 ( .A1(n12210), .A2(n12209), .A3(n12208), .A4(n15449), .ZN(
        n12211) );
  NOR2_X1 U14610 ( .A1(n12211), .A2(n8272), .ZN(n12212) );
  NAND3_X1 U14611 ( .A1(n13558), .A2(n12212), .A3(n8005), .ZN(n12213) );
  NOR3_X1 U14612 ( .A1(n12214), .A2(n13258), .A3(n12213), .ZN(n12215) );
  NAND4_X1 U14613 ( .A1(n13207), .A2(n6618), .A3(n13233), .A4(n12215), .ZN(
        n12216) );
  NOR3_X1 U14614 ( .A1(n13182), .A2(n13194), .A3(n12216), .ZN(n12217) );
  NAND2_X1 U14615 ( .A1(n13164), .A2(n12217), .ZN(n12218) );
  NOR4_X1 U14616 ( .A1(n13127), .A2(n13135), .A3(n13154), .A4(n12218), .ZN(
        n12219) );
  NAND3_X1 U14617 ( .A1(n13093), .A2(n13102), .A3(n12219), .ZN(n12220) );
  NAND3_X1 U14618 ( .A1(n12225), .A2(n12224), .A3(n12223), .ZN(n12226) );
  XNOR2_X1 U14619 ( .A(n12226), .B(n13073), .ZN(n12227) );
  INV_X1 U14620 ( .A(n12235), .ZN(n12231) );
  NAND3_X1 U14621 ( .A1(n12233), .A2(n12232), .A3(n6587), .ZN(n12234) );
  OAI211_X1 U14622 ( .C1(n12236), .C2(n12235), .A(n12234), .B(P3_B_REG_SCAN_IN), .ZN(n12237) );
  NAND2_X1 U14623 ( .A1(n12238), .A2(n12892), .ZN(n12239) );
  XNOR2_X1 U14624 ( .A(n15085), .B(n6801), .ZN(n12241) );
  NAND2_X1 U14625 ( .A1(n12845), .A2(n15435), .ZN(n12245) );
  INV_X1 U14626 ( .A(n12241), .ZN(n12242) );
  OR2_X1 U14627 ( .A1(n12243), .A2(n12242), .ZN(n12244) );
  NAND2_X1 U14628 ( .A1(n12245), .A2(n12244), .ZN(n12788) );
  XNOR2_X1 U14629 ( .A(n12791), .B(n6801), .ZN(n12246) );
  XNOR2_X1 U14630 ( .A(n12246), .B(n12891), .ZN(n12789) );
  NAND2_X1 U14631 ( .A1(n12246), .A2(n13600), .ZN(n12247) );
  XNOR2_X1 U14632 ( .A(n13740), .B(n12771), .ZN(n12831) );
  AND2_X1 U14633 ( .A1(n12831), .A2(n12830), .ZN(n12248) );
  INV_X1 U14634 ( .A(n12831), .ZN(n12249) );
  NAND2_X1 U14635 ( .A1(n12249), .A2(n15065), .ZN(n12250) );
  XNOR2_X1 U14636 ( .A(n6828), .B(n12771), .ZN(n12253) );
  XNOR2_X1 U14637 ( .A(n12253), .B(n12833), .ZN(n12747) );
  INV_X1 U14638 ( .A(n12747), .ZN(n12251) );
  INV_X1 U14639 ( .A(n12253), .ZN(n12254) );
  NAND2_X1 U14640 ( .A1(n12254), .A2(n13601), .ZN(n12255) );
  AND2_X2 U14641 ( .A1(n12744), .A2(n12255), .ZN(n12877) );
  XNOR2_X1 U14642 ( .A(n13680), .B(n6801), .ZN(n12256) );
  XNOR2_X1 U14643 ( .A(n12256), .B(n13582), .ZN(n12876) );
  INV_X1 U14644 ( .A(n12256), .ZN(n12257) );
  NAND2_X1 U14645 ( .A1(n12257), .A2(n13582), .ZN(n12258) );
  NAND2_X1 U14646 ( .A1(n12875), .A2(n12258), .ZN(n12807) );
  XNOR2_X1 U14647 ( .A(n13676), .B(n6801), .ZN(n12259) );
  XNOR2_X1 U14648 ( .A(n12259), .B(n13246), .ZN(n12808) );
  NAND2_X1 U14649 ( .A1(n12807), .A2(n12808), .ZN(n12262) );
  INV_X1 U14650 ( .A(n12259), .ZN(n12260) );
  NAND2_X1 U14651 ( .A1(n12260), .A2(n13246), .ZN(n12261) );
  XNOR2_X1 U14652 ( .A(n13674), .B(n6801), .ZN(n12815) );
  AND2_X1 U14653 ( .A1(n12815), .A2(n12890), .ZN(n12265) );
  INV_X1 U14654 ( .A(n12815), .ZN(n12263) );
  NAND2_X1 U14655 ( .A1(n12263), .A2(n13263), .ZN(n12264) );
  XNOR2_X1 U14656 ( .A(n13242), .B(n6801), .ZN(n12266) );
  XNOR2_X1 U14657 ( .A(n12266), .B(n13247), .ZN(n12856) );
  INV_X1 U14658 ( .A(n12266), .ZN(n12267) );
  XNOR2_X1 U14659 ( .A(n13729), .B(n12771), .ZN(n12268) );
  XNOR2_X1 U14660 ( .A(n12268), .B(n13212), .ZN(n12762) );
  INV_X1 U14661 ( .A(n12268), .ZN(n12269) );
  NAND2_X1 U14662 ( .A1(n12269), .A2(n13212), .ZN(n12270) );
  NAND2_X1 U14663 ( .A1(n12761), .A2(n12270), .ZN(n12824) );
  XNOR2_X1 U14664 ( .A(n12271), .B(n6801), .ZN(n12272) );
  XNOR2_X1 U14665 ( .A(n12272), .B(n12889), .ZN(n12823) );
  NAND2_X1 U14666 ( .A1(n12824), .A2(n12823), .ZN(n12822) );
  INV_X1 U14667 ( .A(n12272), .ZN(n12273) );
  NAND2_X1 U14668 ( .A1(n12273), .A2(n12889), .ZN(n12274) );
  NAND2_X1 U14669 ( .A1(n12822), .A2(n12274), .ZN(n12781) );
  XNOR2_X1 U14670 ( .A(n13198), .B(n12771), .ZN(n12275) );
  XNOR2_X1 U14671 ( .A(n12275), .B(n13211), .ZN(n12782) );
  OR2_X2 U14672 ( .A1(n12781), .A2(n12782), .ZN(n12779) );
  INV_X1 U14673 ( .A(n12275), .ZN(n12276) );
  NAND2_X1 U14674 ( .A1(n12276), .A2(n13185), .ZN(n12277) );
  NAND2_X2 U14675 ( .A1(n12779), .A2(n12277), .ZN(n12733) );
  XNOR2_X1 U14676 ( .A(n13187), .B(n12771), .ZN(n12721) );
  XNOR2_X1 U14677 ( .A(n12733), .B(n12721), .ZN(n12839) );
  INV_X1 U14678 ( .A(n12721), .ZN(n12723) );
  AND2_X1 U14679 ( .A1(n12733), .A2(n12723), .ZN(n12278) );
  XNOR2_X1 U14680 ( .A(n13175), .B(n6801), .ZN(n12726) );
  XNOR2_X1 U14681 ( .A(n13640), .B(n6801), .ZN(n12730) );
  AOI22_X1 U14682 ( .A1(n13152), .A2(n12878), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12281) );
  OAI21_X1 U14683 ( .B1(n13186), .B2(n12880), .A(n12281), .ZN(n12283) );
  NOR2_X1 U14684 ( .A1(n13640), .A2(n12885), .ZN(n12282) );
  AOI211_X1 U14685 ( .C1(n13159), .C2(n12882), .A(n12283), .B(n12282), .ZN(
        n12284) );
  NAND2_X1 U14686 ( .A1(n14298), .A2(n12456), .ZN(n12287) );
  INV_X1 U14687 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12285) );
  OR2_X1 U14688 ( .A1(n12458), .A2(n12285), .ZN(n12286) );
  INV_X1 U14689 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14864) );
  NAND2_X1 U14690 ( .A1(n12450), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12291) );
  INV_X1 U14691 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n12288) );
  OR2_X1 U14692 ( .A1(n12289), .A2(n12288), .ZN(n12290) );
  OAI211_X1 U14693 ( .C1(n12454), .C2(n14864), .A(n12291), .B(n12290), .ZN(
        n14587) );
  INV_X1 U14694 ( .A(n14587), .ZN(n12480) );
  XNOR2_X1 U14695 ( .A(n14583), .B(n12480), .ZN(n12520) );
  NOR2_X1 U14696 ( .A1(n15034), .A2(n12296), .ZN(n12292) );
  OR2_X1 U14697 ( .A1(n12293), .A2(n12292), .ZN(n12295) );
  NAND2_X1 U14698 ( .A1(n12295), .A2(n12294), .ZN(n12477) );
  NOR2_X1 U14699 ( .A1(n12520), .A2(n12477), .ZN(n12527) );
  MUX2_X1 U14700 ( .A(n14470), .B(n12345), .S(n12413), .Z(n12350) );
  NAND2_X1 U14701 ( .A1(n12299), .A2(n12455), .ZN(n12297) );
  OAI21_X1 U14702 ( .B1(n12299), .B2(n12298), .A(n12297), .ZN(n12301) );
  OAI21_X1 U14703 ( .B1(n15232), .B2(n12300), .A(n12301), .ZN(n12304) );
  INV_X1 U14704 ( .A(n12301), .ZN(n12302) );
  AOI22_X1 U14705 ( .A1(n14476), .A2(n12304), .B1(n12303), .B2(n12302), .ZN(
        n12306) );
  NAND2_X1 U14706 ( .A1(n12487), .A2(n12339), .ZN(n12305) );
  AOI21_X1 U14707 ( .B1(n12306), .B2(n12305), .A(n12490), .ZN(n12311) );
  OAI21_X1 U14708 ( .B1(n12311), .B2(n12310), .A(n12309), .ZN(n12318) );
  OAI21_X1 U14709 ( .B1(n12315), .B2(n12314), .A(n12313), .ZN(n12316) );
  NAND3_X1 U14710 ( .A1(n12318), .A2(n12317), .A3(n12316), .ZN(n12323) );
  AND2_X1 U14711 ( .A1(n15236), .A2(n14474), .ZN(n12320) );
  MUX2_X1 U14712 ( .A(n12320), .B(n12319), .S(n6588), .Z(n12321) );
  INV_X1 U14713 ( .A(n12321), .ZN(n12322) );
  MUX2_X1 U14714 ( .A(n14473), .B(n12324), .S(n6588), .Z(n12328) );
  MUX2_X1 U14715 ( .A(n12326), .B(n12325), .S(n12339), .Z(n12327) );
  MUX2_X1 U14716 ( .A(n12330), .B(n14472), .S(n6588), .Z(n12334) );
  NAND2_X1 U14717 ( .A1(n12333), .A2(n12334), .ZN(n12332) );
  MUX2_X1 U14718 ( .A(n12330), .B(n14472), .S(n12339), .Z(n12331) );
  NAND2_X1 U14719 ( .A1(n12332), .A2(n12331), .ZN(n12338) );
  INV_X1 U14720 ( .A(n12333), .ZN(n12336) );
  NAND2_X1 U14721 ( .A1(n12336), .A2(n12335), .ZN(n12337) );
  NAND2_X1 U14722 ( .A1(n12338), .A2(n12337), .ZN(n12344) );
  MUX2_X1 U14723 ( .A(n14429), .B(n14471), .S(n12339), .Z(n12343) );
  MUX2_X1 U14724 ( .A(n12341), .B(n12340), .S(n6588), .Z(n12342) );
  MUX2_X1 U14725 ( .A(n12345), .B(n14470), .S(n12413), .Z(n12346) );
  NAND2_X1 U14726 ( .A1(n12347), .A2(n12346), .ZN(n12348) );
  OAI21_X1 U14727 ( .B1(n12350), .B2(n12349), .A(n12348), .ZN(n12353) );
  MUX2_X1 U14728 ( .A(n14469), .B(n12351), .S(n6588), .Z(n12354) );
  INV_X1 U14729 ( .A(n6588), .ZN(n12413) );
  MUX2_X1 U14730 ( .A(n14469), .B(n12351), .S(n12413), .Z(n12352) );
  INV_X1 U14731 ( .A(n12354), .ZN(n12355) );
  MUX2_X1 U14732 ( .A(n14468), .B(n12356), .S(n12413), .Z(n12360) );
  MUX2_X1 U14733 ( .A(n14468), .B(n12356), .S(n12439), .Z(n12357) );
  NAND2_X1 U14734 ( .A1(n12358), .A2(n12357), .ZN(n12364) );
  INV_X1 U14735 ( .A(n12360), .ZN(n12361) );
  NAND2_X1 U14736 ( .A1(n12362), .A2(n12361), .ZN(n12363) );
  NAND2_X1 U14737 ( .A1(n12364), .A2(n12363), .ZN(n12366) );
  MUX2_X1 U14738 ( .A(n14467), .B(n15249), .S(n12439), .Z(n12367) );
  MUX2_X1 U14739 ( .A(n14467), .B(n15249), .S(n12413), .Z(n12365) );
  INV_X1 U14740 ( .A(n12367), .ZN(n12368) );
  MUX2_X1 U14741 ( .A(n14466), .B(n12369), .S(n12413), .Z(n12372) );
  MUX2_X1 U14742 ( .A(n14466), .B(n12369), .S(n6588), .Z(n12370) );
  NAND2_X1 U14743 ( .A1(n12371), .A2(n12370), .ZN(n12374) );
  NAND2_X1 U14744 ( .A1(n12374), .A2(n12373), .ZN(n12377) );
  MUX2_X1 U14745 ( .A(n14465), .B(n12375), .S(n12417), .Z(n12378) );
  MUX2_X1 U14746 ( .A(n14465), .B(n12375), .S(n12467), .Z(n12376) );
  INV_X1 U14747 ( .A(n12378), .ZN(n12379) );
  MUX2_X1 U14748 ( .A(n14464), .B(n12380), .S(n12467), .Z(n12383) );
  MUX2_X1 U14749 ( .A(n14464), .B(n12380), .S(n12417), .Z(n12381) );
  INV_X1 U14750 ( .A(n12381), .ZN(n12382) );
  AOI21_X1 U14751 ( .B1(n12396), .B2(n12385), .A(n12439), .ZN(n12386) );
  NAND2_X1 U14752 ( .A1(n12388), .A2(n12387), .ZN(n12389) );
  NAND2_X1 U14753 ( .A1(n12389), .A2(n12439), .ZN(n12398) );
  MUX2_X1 U14754 ( .A(n14805), .B(n15012), .S(n12467), .Z(n12402) );
  AND2_X1 U14755 ( .A1(n14461), .A2(n12467), .ZN(n12390) );
  AOI21_X1 U14756 ( .B1(n14830), .B2(n12439), .A(n12390), .ZN(n12392) );
  NAND2_X1 U14757 ( .A1(n14954), .A2(n14825), .ZN(n12391) );
  NAND3_X1 U14758 ( .A1(n12393), .A2(n12392), .A3(n12391), .ZN(n12403) );
  OAI21_X1 U14759 ( .B1(n12394), .B2(n12402), .A(n12403), .ZN(n12395) );
  OAI21_X1 U14760 ( .B1(n12467), .B2(n12396), .A(n12395), .ZN(n12397) );
  AND2_X1 U14761 ( .A1(n14790), .A2(n12417), .ZN(n12400) );
  OAI21_X1 U14762 ( .B1(n14790), .B2(n12439), .A(n14954), .ZN(n12399) );
  OAI21_X1 U14763 ( .B1(n12400), .B2(n14954), .A(n12399), .ZN(n12401) );
  OAI21_X1 U14764 ( .B1(n12403), .B2(n12402), .A(n12401), .ZN(n12404) );
  NAND2_X1 U14765 ( .A1(n14786), .A2(n12467), .ZN(n12406) );
  OR2_X1 U14766 ( .A1(n14786), .A2(n12467), .ZN(n12405) );
  MUX2_X1 U14767 ( .A(n12406), .B(n12405), .S(n14802), .Z(n12407) );
  NAND2_X1 U14768 ( .A1(n12408), .A2(n14763), .ZN(n12412) );
  NAND2_X1 U14769 ( .A1(n14792), .A2(n12439), .ZN(n12410) );
  OR2_X1 U14770 ( .A1(n14792), .A2(n12439), .ZN(n12409) );
  MUX2_X1 U14771 ( .A(n12410), .B(n12409), .S(n14765), .Z(n12411) );
  NAND2_X1 U14772 ( .A1(n12412), .A2(n12411), .ZN(n12416) );
  INV_X1 U14773 ( .A(n14999), .ZN(n14754) );
  MUX2_X1 U14774 ( .A(n14460), .B(n14754), .S(n12467), .Z(n12415) );
  INV_X1 U14775 ( .A(n12413), .ZN(n12417) );
  MUX2_X1 U14776 ( .A(n14352), .B(n14999), .S(n12417), .Z(n12414) );
  INV_X1 U14777 ( .A(n14925), .ZN(n14742) );
  MUX2_X1 U14778 ( .A(n14459), .B(n14742), .S(n12417), .Z(n12419) );
  MUX2_X1 U14779 ( .A(n14398), .B(n14925), .S(n12467), .Z(n12418) );
  INV_X1 U14780 ( .A(n14917), .ZN(n14729) );
  MUX2_X1 U14781 ( .A(n14712), .B(n14729), .S(n12467), .Z(n12422) );
  MUX2_X1 U14782 ( .A(n14351), .B(n14917), .S(n12439), .Z(n12420) );
  NOR2_X1 U14783 ( .A1(n12423), .A2(n12422), .ZN(n12424) );
  MUX2_X1 U14784 ( .A(n14685), .B(n14909), .S(n12439), .Z(n12425) );
  MUX2_X1 U14785 ( .A(n14685), .B(n14909), .S(n12467), .Z(n12427) );
  NAND2_X1 U14786 ( .A1(n12429), .A2(n12428), .ZN(n12431) );
  MUX2_X1 U14787 ( .A(n14711), .B(n14691), .S(n12467), .Z(n12432) );
  MUX2_X1 U14788 ( .A(n14711), .B(n14691), .S(n12439), .Z(n12430) );
  INV_X1 U14789 ( .A(n12413), .ZN(n12439) );
  MUX2_X1 U14790 ( .A(n14684), .B(n14987), .S(n12439), .Z(n12435) );
  MUX2_X1 U14791 ( .A(n14684), .B(n14987), .S(n12467), .Z(n12433) );
  MUX2_X1 U14792 ( .A(n14633), .B(n14887), .S(n12467), .Z(n12438) );
  MUX2_X1 U14793 ( .A(n14633), .B(n14887), .S(n12439), .Z(n12437) );
  MUX2_X1 U14794 ( .A(n14656), .B(n14878), .S(n12439), .Z(n12442) );
  MUX2_X1 U14795 ( .A(n14656), .B(n14878), .S(n12467), .Z(n12440) );
  INV_X1 U14796 ( .A(n12442), .ZN(n12443) );
  MUX2_X1 U14797 ( .A(n14634), .B(n14980), .S(n12413), .Z(n12446) );
  MUX2_X1 U14798 ( .A(n14634), .B(n14980), .S(n12439), .Z(n12444) );
  NAND2_X1 U14799 ( .A1(n12447), .A2(n12456), .ZN(n12449) );
  OR2_X1 U14800 ( .A1(n12458), .A2(n15021), .ZN(n12448) );
  MUX2_X1 U14801 ( .A(n14458), .B(n14870), .S(n12439), .Z(n12470) );
  INV_X1 U14802 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14868) );
  NAND2_X1 U14803 ( .A1(n12450), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12453) );
  INV_X1 U14804 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n12451) );
  OR2_X1 U14805 ( .A1(n12289), .A2(n12451), .ZN(n12452) );
  OAI211_X1 U14806 ( .C1(n12454), .C2(n14868), .A(n12453), .B(n12452), .ZN(
        n14604) );
  OAI21_X1 U14807 ( .B1(n14587), .B2(n12455), .A(n14604), .ZN(n12461) );
  NAND2_X1 U14808 ( .A1(n12457), .A2(n12456), .ZN(n12460) );
  OR2_X1 U14809 ( .A1(n12458), .A2(n15018), .ZN(n12459) );
  MUX2_X1 U14810 ( .A(n12461), .B(n14977), .S(n12467), .Z(n12471) );
  NAND2_X1 U14811 ( .A1(n14591), .A2(n12439), .ZN(n12466) );
  NAND2_X1 U14812 ( .A1(n12467), .A2(n14587), .ZN(n12463) );
  NAND2_X1 U14813 ( .A1(n12463), .A2(n12462), .ZN(n12464) );
  NAND2_X1 U14814 ( .A1(n12464), .A2(n14604), .ZN(n12465) );
  NAND2_X1 U14815 ( .A1(n12466), .A2(n12465), .ZN(n12472) );
  INV_X1 U14816 ( .A(n14458), .ZN(n12468) );
  MUX2_X1 U14817 ( .A(n12468), .B(n14611), .S(n12467), .Z(n12469) );
  INV_X1 U14818 ( .A(n12471), .ZN(n12474) );
  INV_X1 U14819 ( .A(n12472), .ZN(n12473) );
  NAND2_X1 U14820 ( .A1(n12476), .A2(n12475), .ZN(n12526) );
  INV_X1 U14821 ( .A(n12477), .ZN(n12483) );
  INV_X1 U14822 ( .A(n12520), .ZN(n12479) );
  AND2_X1 U14823 ( .A1(n12477), .A2(n12522), .ZN(n12484) );
  INV_X1 U14824 ( .A(n12484), .ZN(n12478) );
  NOR2_X1 U14825 ( .A1(n12479), .A2(n12478), .ZN(n12482) );
  MUX2_X1 U14826 ( .A(n12480), .B(n14973), .S(n12439), .Z(n12481) );
  OAI21_X1 U14827 ( .B1(n14587), .B2(n14583), .A(n12481), .ZN(n12485) );
  MUX2_X1 U14828 ( .A(n12483), .B(n12482), .S(n12485), .Z(n12525) );
  NAND2_X1 U14829 ( .A1(n12485), .A2(n12484), .ZN(n12524) );
  INV_X1 U14830 ( .A(n14604), .ZN(n12486) );
  XOR2_X1 U14831 ( .A(n14458), .B(n14870), .Z(n14600) );
  INV_X1 U14832 ( .A(n14763), .ZN(n12510) );
  INV_X1 U14833 ( .A(n12487), .ZN(n12488) );
  OAI21_X1 U14834 ( .B1(n15232), .B2(n12489), .A(n12488), .ZN(n15226) );
  NOR4_X1 U14835 ( .A1(n12491), .A2(n10328), .A3(n12490), .A4(n15226), .ZN(
        n12494) );
  NAND4_X1 U14836 ( .A1(n12495), .A2(n12494), .A3(n12493), .A4(n12492), .ZN(
        n12496) );
  NOR4_X1 U14837 ( .A1(n12499), .A2(n12498), .A3(n12497), .A4(n12496), .ZN(
        n12502) );
  NAND4_X1 U14838 ( .A1(n7309), .A2(n12502), .A3(n12501), .A4(n12500), .ZN(
        n12503) );
  NOR4_X1 U14839 ( .A1(n12506), .A2(n12505), .A3(n12504), .A4(n12503), .ZN(
        n12508) );
  NAND3_X1 U14840 ( .A1(n14799), .A2(n12508), .A3(n12507), .ZN(n12509) );
  NOR4_X1 U14841 ( .A1(n12511), .A2(n12510), .A3(n7426), .A4(n12509), .ZN(
        n12512) );
  NAND4_X1 U14842 ( .A1(n14708), .A2(n14718), .A3(n12512), .A4(n14734), .ZN(
        n12513) );
  NOR3_X1 U14843 ( .A1(n14649), .A2(n12514), .A3(n12513), .ZN(n12516) );
  NAND4_X1 U14844 ( .A1(n12517), .A2(n12516), .A3(n12515), .A4(n14631), .ZN(
        n12518) );
  XNOR2_X1 U14845 ( .A(n12521), .B(n14768), .ZN(n12523) );
  NOR3_X1 U14846 ( .A1(n12528), .A2(n6584), .A3(n14824), .ZN(n12530) );
  OAI21_X1 U14847 ( .B1(n12531), .B2(n15034), .A(P1_B_REG_SCAN_IN), .ZN(n12529) );
  OAI22_X1 U14848 ( .A1(n12532), .A2(n12531), .B1(n12530), .B2(n12529), .ZN(
        P1_U3242) );
  INV_X1 U14849 ( .A(n12533), .ZN(n12534) );
  OAI222_X1 U14850 ( .A1(n12609), .A2(n12535), .B1(n13756), .B2(n12534), .C1(
        P3_U3151), .C2(n8297), .ZN(P3_U3267) );
  XNOR2_X1 U14851 ( .A(n14222), .B(n12592), .ZN(n12568) );
  NAND2_X1 U14852 ( .A1(n13897), .A2(n13997), .ZN(n12569) );
  NAND2_X1 U14853 ( .A1(n12537), .A2(n12536), .ZN(n12542) );
  INV_X1 U14854 ( .A(n12538), .ZN(n12539) );
  NAND2_X1 U14855 ( .A1(n12540), .A2(n12539), .ZN(n12541) );
  XNOR2_X1 U14856 ( .A(n15119), .B(n13792), .ZN(n12543) );
  NAND2_X1 U14857 ( .A1(n13904), .A2(n13997), .ZN(n12544) );
  NAND2_X1 U14858 ( .A1(n12543), .A2(n12544), .ZN(n12549) );
  INV_X1 U14859 ( .A(n12543), .ZN(n12546) );
  INV_X1 U14860 ( .A(n12544), .ZN(n12545) );
  NAND2_X1 U14861 ( .A1(n12546), .A2(n12545), .ZN(n12547) );
  NAND2_X1 U14862 ( .A1(n12549), .A2(n12547), .ZN(n15100) );
  XOR2_X1 U14863 ( .A(n12592), .B(n14257), .Z(n12551) );
  NAND2_X1 U14864 ( .A1(n13903), .A2(n13997), .ZN(n13874) );
  XNOR2_X1 U14865 ( .A(n14251), .B(n13792), .ZN(n12553) );
  NAND2_X1 U14866 ( .A1(n13902), .A2(n13997), .ZN(n12552) );
  NAND2_X1 U14867 ( .A1(n12553), .A2(n12552), .ZN(n12554) );
  OAI21_X1 U14868 ( .B1(n12553), .B2(n12552), .A(n12554), .ZN(n13831) );
  INV_X1 U14869 ( .A(n12554), .ZN(n12555) );
  XNOR2_X1 U14870 ( .A(n14293), .B(n13792), .ZN(n12557) );
  NAND2_X1 U14871 ( .A1(n13901), .A2(n13997), .ZN(n12556) );
  NAND2_X1 U14872 ( .A1(n12557), .A2(n12556), .ZN(n12558) );
  OAI21_X1 U14873 ( .B1(n12557), .B2(n12556), .A(n12558), .ZN(n13840) );
  INV_X1 U14874 ( .A(n12558), .ZN(n12559) );
  XNOR2_X1 U14875 ( .A(n14237), .B(n12592), .ZN(n12561) );
  NAND2_X1 U14876 ( .A1(n13900), .A2(n13997), .ZN(n12560) );
  XNOR2_X1 U14877 ( .A(n12561), .B(n12560), .ZN(n13865) );
  INV_X1 U14878 ( .A(n12560), .ZN(n12562) );
  XNOR2_X1 U14879 ( .A(n14233), .B(n12592), .ZN(n13777) );
  AND2_X1 U14880 ( .A1(n13899), .A2(n13997), .ZN(n12563) );
  NOR2_X1 U14881 ( .A1(n13777), .A2(n12563), .ZN(n13781) );
  INV_X1 U14882 ( .A(n13777), .ZN(n12565) );
  INV_X1 U14883 ( .A(n12563), .ZN(n12564) );
  NOR2_X1 U14884 ( .A1(n12565), .A2(n12564), .ZN(n13782) );
  XNOR2_X1 U14885 ( .A(n14116), .B(n12592), .ZN(n12567) );
  AND2_X1 U14886 ( .A1(n13898), .A2(n13997), .ZN(n12566) );
  NAND2_X1 U14887 ( .A1(n12567), .A2(n12566), .ZN(n13858) );
  XNOR2_X1 U14888 ( .A(n12568), .B(n12569), .ZN(n13808) );
  XNOR2_X1 U14889 ( .A(n14087), .B(n12592), .ZN(n12578) );
  INV_X1 U14890 ( .A(n12571), .ZN(n12572) );
  AOI22_X1 U14891 ( .A1(n12572), .A2(n15104), .B1(n13875), .B2(n13896), .ZN(
        n12577) );
  AOI22_X1 U14892 ( .A1(n13895), .A2(n14027), .B1(n14025), .B2(n13897), .ZN(
        n14083) );
  OAI22_X1 U14893 ( .A1(n14083), .A2(n13853), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12573), .ZN(n12574) );
  AOI21_X1 U14894 ( .B1(n14088), .B2(n13855), .A(n12574), .ZN(n12576) );
  NAND2_X1 U14895 ( .A1(n14087), .A2(n15107), .ZN(n12575) );
  OAI211_X1 U14896 ( .C1(n12581), .C2(n12577), .A(n12576), .B(n12575), .ZN(
        P2_U3207) );
  AND2_X1 U14897 ( .A1(n12579), .A2(n12578), .ZN(n12580) );
  XNOR2_X1 U14898 ( .A(n14210), .B(n12592), .ZN(n12583) );
  XNOR2_X1 U14899 ( .A(n12585), .B(n12583), .ZN(n13770) );
  AND2_X1 U14900 ( .A1(n13895), .A2(n13997), .ZN(n12582) );
  NAND2_X1 U14901 ( .A1(n13770), .A2(n12582), .ZN(n13769) );
  INV_X1 U14902 ( .A(n12583), .ZN(n12584) );
  XNOR2_X1 U14903 ( .A(n14205), .B(n13792), .ZN(n13818) );
  NAND2_X1 U14904 ( .A1(n14026), .A2(n13997), .ZN(n12586) );
  NOR2_X1 U14905 ( .A1(n13818), .A2(n12586), .ZN(n12591) );
  AOI21_X1 U14906 ( .B1(n13818), .B2(n12586), .A(n12591), .ZN(n13850) );
  XNOR2_X1 U14907 ( .A(n14031), .B(n12592), .ZN(n12594) );
  AND2_X1 U14908 ( .A1(n13894), .A2(n13997), .ZN(n12587) );
  NAND2_X1 U14909 ( .A1(n12594), .A2(n12587), .ZN(n12593) );
  INV_X1 U14910 ( .A(n12594), .ZN(n12589) );
  INV_X1 U14911 ( .A(n12587), .ZN(n12588) );
  NAND2_X1 U14912 ( .A1(n12589), .A2(n12588), .ZN(n12590) );
  AND2_X1 U14913 ( .A1(n12593), .A2(n12590), .ZN(n13816) );
  XNOR2_X1 U14914 ( .A(n14196), .B(n12592), .ZN(n13759) );
  NAND2_X1 U14915 ( .A1(n14028), .A2(n13997), .ZN(n13757) );
  XNOR2_X1 U14916 ( .A(n13759), .B(n13757), .ZN(n12596) );
  NAND3_X1 U14917 ( .A1(n12594), .A2(n13875), .A3(n13894), .ZN(n12595) );
  OAI21_X1 U14918 ( .B1(n13814), .B2(n13872), .A(n12595), .ZN(n12598) );
  INV_X1 U14919 ( .A(n12596), .ZN(n12597) );
  NAND2_X1 U14920 ( .A1(n12598), .A2(n12597), .ZN(n12602) );
  AOI22_X1 U14921 ( .A1(n13893), .A2(n14027), .B1(n14025), .B2(n13894), .ZN(
        n14017) );
  AOI22_X1 U14922 ( .A1(n14011), .A2(n13855), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12599) );
  OAI21_X1 U14923 ( .B1(n14017), .B2(n13853), .A(n12599), .ZN(n12600) );
  AOI21_X1 U14924 ( .B1(n14196), .B2(n15107), .A(n12600), .ZN(n12601) );
  OAI211_X1 U14925 ( .C1(n13761), .C2(n13872), .A(n12602), .B(n12601), .ZN(
        P2_U3212) );
  INV_X1 U14926 ( .A(n12603), .ZN(n12604) );
  OAI222_X1 U14927 ( .A1(n14312), .A2(n12605), .B1(n10596), .B2(n12604), .C1(
        P2_U3088), .C2(n9019), .ZN(P2_U3305) );
  INV_X1 U14928 ( .A(n12606), .ZN(n12607) );
  OAI222_X1 U14929 ( .A1(P3_U3151), .A2(n6587), .B1(n12609), .B2(n12612), .C1(
        n13756), .C2(n12611), .ZN(P3_U3268) );
  AND2_X1 U14930 ( .A1(n12709), .A2(n14792), .ZN(n12613) );
  AOI21_X1 U14931 ( .B1(n14765), .B2(n10103), .A(n12613), .ZN(n12650) );
  NAND2_X1 U14932 ( .A1(n14765), .A2(n12708), .ZN(n12615) );
  NAND2_X1 U14933 ( .A1(n14792), .A2(n10103), .ZN(n12614) );
  NAND2_X1 U14934 ( .A1(n12615), .A2(n12614), .ZN(n12616) );
  XNOR2_X1 U14935 ( .A(n12616), .B(n12710), .ZN(n12649) );
  NAND2_X1 U14936 ( .A1(n14967), .A2(n12708), .ZN(n12620) );
  NAND2_X1 U14937 ( .A1(n10103), .A2(n14462), .ZN(n12619) );
  NAND2_X1 U14938 ( .A1(n12620), .A2(n12619), .ZN(n12621) );
  XNOR2_X1 U14939 ( .A(n12621), .B(n12710), .ZN(n12623) );
  XNOR2_X2 U14940 ( .A(n12622), .B(n12623), .ZN(n14446) );
  OAI22_X1 U14941 ( .A1(n7152), .A2(n6749), .B1(n14823), .B2(n6812), .ZN(
        n14445) );
  NAND2_X1 U14942 ( .A1(n14830), .A2(n12708), .ZN(n12625) );
  NAND2_X1 U14943 ( .A1(n10103), .A2(n14461), .ZN(n12624) );
  NAND2_X1 U14944 ( .A1(n12625), .A2(n12624), .ZN(n12626) );
  XNOR2_X1 U14945 ( .A(n12626), .B(n12710), .ZN(n12630) );
  NAND2_X1 U14946 ( .A1(n14830), .A2(n10103), .ZN(n12628) );
  NAND2_X1 U14947 ( .A1(n12709), .A2(n14461), .ZN(n12627) );
  NAND2_X1 U14948 ( .A1(n12628), .A2(n12627), .ZN(n12629) );
  NOR2_X1 U14949 ( .A1(n12630), .A2(n12629), .ZN(n12631) );
  AOI21_X1 U14950 ( .B1(n12630), .B2(n12629), .A(n12631), .ZN(n14369) );
  INV_X1 U14951 ( .A(n12631), .ZN(n12632) );
  NAND2_X1 U14952 ( .A1(n14954), .A2(n12708), .ZN(n12634) );
  NAND2_X1 U14953 ( .A1(n10103), .A2(n14790), .ZN(n12633) );
  NAND2_X1 U14954 ( .A1(n12634), .A2(n12633), .ZN(n12635) );
  XNOR2_X1 U14955 ( .A(n12635), .B(n12710), .ZN(n12638) );
  NAND2_X1 U14956 ( .A1(n14954), .A2(n10103), .ZN(n12637) );
  NAND2_X1 U14957 ( .A1(n12709), .A2(n14790), .ZN(n12636) );
  NAND2_X1 U14958 ( .A1(n12637), .A2(n12636), .ZN(n12639) );
  NAND2_X1 U14959 ( .A1(n12638), .A2(n12639), .ZN(n14379) );
  INV_X1 U14960 ( .A(n12638), .ZN(n12641) );
  INV_X1 U14961 ( .A(n12639), .ZN(n12640) );
  NAND2_X1 U14962 ( .A1(n12641), .A2(n12640), .ZN(n14378) );
  NAND2_X1 U14963 ( .A1(n14786), .A2(n12708), .ZN(n12643) );
  NAND2_X1 U14964 ( .A1(n14802), .A2(n10103), .ZN(n12642) );
  NAND2_X1 U14965 ( .A1(n12643), .A2(n12642), .ZN(n12644) );
  XNOR2_X1 U14966 ( .A(n12644), .B(n12710), .ZN(n12647) );
  AOI22_X1 U14967 ( .A1(n14786), .A2(n10103), .B1(n12709), .B2(n14802), .ZN(
        n12645) );
  XNOR2_X1 U14968 ( .A(n12647), .B(n12645), .ZN(n14417) );
  INV_X1 U14969 ( .A(n12645), .ZN(n12646) );
  XOR2_X1 U14970 ( .A(n12650), .B(n12649), .Z(n14337) );
  OAI22_X1 U14971 ( .A1(n14999), .A2(n12666), .B1(n14352), .B2(n6749), .ZN(
        n12651) );
  XNOR2_X1 U14972 ( .A(n12651), .B(n12710), .ZN(n12655) );
  AND2_X1 U14973 ( .A1(n14460), .A2(n12709), .ZN(n12652) );
  AOI21_X1 U14974 ( .B1(n14754), .B2(n10103), .A(n12652), .ZN(n12653) );
  XNOR2_X1 U14975 ( .A(n12655), .B(n12653), .ZN(n14396) );
  INV_X1 U14976 ( .A(n12653), .ZN(n12654) );
  NAND2_X1 U14977 ( .A1(n12655), .A2(n12654), .ZN(n12656) );
  OAI22_X1 U14978 ( .A1(n14925), .A2(n12666), .B1(n14398), .B2(n6749), .ZN(
        n12657) );
  XNOR2_X1 U14979 ( .A(n12657), .B(n12710), .ZN(n12659) );
  OAI22_X1 U14980 ( .A1(n14925), .A2(n6749), .B1(n14398), .B2(n6812), .ZN(
        n12660) );
  XNOR2_X1 U14981 ( .A(n12659), .B(n12660), .ZN(n14350) );
  INV_X1 U14982 ( .A(n14350), .ZN(n12658) );
  INV_X1 U14983 ( .A(n12659), .ZN(n12662) );
  INV_X1 U14984 ( .A(n12660), .ZN(n12661) );
  NAND2_X1 U14985 ( .A1(n12662), .A2(n12661), .ZN(n12663) );
  OAI22_X1 U14986 ( .A1(n14917), .A2(n6749), .B1(n14351), .B2(n6812), .ZN(
        n12669) );
  OAI22_X1 U14987 ( .A1(n14917), .A2(n12666), .B1(n14351), .B2(n6749), .ZN(
        n12667) );
  XNOR2_X1 U14988 ( .A(n12667), .B(n12710), .ZN(n12668) );
  XOR2_X1 U14989 ( .A(n12669), .B(n12668), .Z(n14407) );
  INV_X1 U14990 ( .A(n12668), .ZN(n12671) );
  INV_X1 U14991 ( .A(n12669), .ZN(n12670) );
  NAND2_X1 U14992 ( .A1(n12671), .A2(n12670), .ZN(n12672) );
  NAND2_X1 U14993 ( .A1(n14909), .A2(n12708), .ZN(n12674) );
  NAND2_X1 U14994 ( .A1(n10103), .A2(n14685), .ZN(n12673) );
  NAND2_X1 U14995 ( .A1(n12674), .A2(n12673), .ZN(n12675) );
  XNOR2_X1 U14996 ( .A(n12675), .B(n12710), .ZN(n12676) );
  AOI22_X1 U14997 ( .A1(n14909), .A2(n10103), .B1(n12709), .B2(n14685), .ZN(
        n12677) );
  XNOR2_X1 U14998 ( .A(n12676), .B(n12677), .ZN(n14323) );
  INV_X1 U14999 ( .A(n12676), .ZN(n12678) );
  NAND2_X1 U15000 ( .A1(n14691), .A2(n12708), .ZN(n12680) );
  NAND2_X1 U15001 ( .A1(n10103), .A2(n14711), .ZN(n12679) );
  NAND2_X1 U15002 ( .A1(n12680), .A2(n12679), .ZN(n12681) );
  XNOR2_X1 U15003 ( .A(n12681), .B(n12710), .ZN(n12682) );
  AOI22_X1 U15004 ( .A1(n14691), .A2(n10103), .B1(n12709), .B2(n14711), .ZN(
        n12683) );
  XNOR2_X1 U15005 ( .A(n12682), .B(n12683), .ZN(n14389) );
  NAND2_X1 U15006 ( .A1(n14388), .A2(n14389), .ZN(n12686) );
  INV_X1 U15007 ( .A(n12682), .ZN(n12684) );
  NAND2_X1 U15008 ( .A1(n12684), .A2(n12683), .ZN(n12685) );
  NAND2_X1 U15009 ( .A1(n14987), .A2(n12708), .ZN(n12688) );
  NAND2_X1 U15010 ( .A1(n10103), .A2(n14684), .ZN(n12687) );
  NAND2_X1 U15011 ( .A1(n12688), .A2(n12687), .ZN(n12689) );
  XNOR2_X1 U15012 ( .A(n12689), .B(n12710), .ZN(n12690) );
  AOI22_X1 U15013 ( .A1(n14987), .A2(n10103), .B1(n12709), .B2(n14684), .ZN(
        n12691) );
  XNOR2_X1 U15014 ( .A(n12690), .B(n12691), .ZN(n14359) );
  NAND2_X1 U15015 ( .A1(n14358), .A2(n14359), .ZN(n12694) );
  INV_X1 U15016 ( .A(n12690), .ZN(n12692) );
  NAND2_X1 U15017 ( .A1(n12692), .A2(n12691), .ZN(n12693) );
  NAND2_X1 U15018 ( .A1(n14887), .A2(n12708), .ZN(n12696) );
  NAND2_X1 U15019 ( .A1(n10103), .A2(n14633), .ZN(n12695) );
  NAND2_X1 U15020 ( .A1(n12696), .A2(n12695), .ZN(n12697) );
  XNOR2_X1 U15021 ( .A(n12697), .B(n12710), .ZN(n12698) );
  AOI22_X1 U15022 ( .A1(n14887), .A2(n10103), .B1(n12709), .B2(n14633), .ZN(
        n12699) );
  XNOR2_X1 U15023 ( .A(n12698), .B(n12699), .ZN(n14437) );
  INV_X1 U15024 ( .A(n12698), .ZN(n12700) );
  NAND2_X1 U15025 ( .A1(n12700), .A2(n12699), .ZN(n12701) );
  NAND2_X1 U15026 ( .A1(n14878), .A2(n12708), .ZN(n12703) );
  NAND2_X1 U15027 ( .A1(n10103), .A2(n14656), .ZN(n12702) );
  NAND2_X1 U15028 ( .A1(n12703), .A2(n12702), .ZN(n12704) );
  XNOR2_X1 U15029 ( .A(n12704), .B(n12710), .ZN(n12705) );
  AOI22_X1 U15030 ( .A1(n14878), .A2(n10103), .B1(n12709), .B2(n14656), .ZN(
        n12706) );
  XNOR2_X1 U15031 ( .A(n12705), .B(n12706), .ZN(n14316) );
  INV_X1 U15032 ( .A(n12705), .ZN(n12707) );
  AOI22_X1 U15033 ( .A1(n14980), .A2(n12708), .B1(n10103), .B2(n14634), .ZN(
        n12713) );
  AOI22_X1 U15034 ( .A1(n14980), .A2(n10103), .B1(n12709), .B2(n14634), .ZN(
        n12711) );
  XNOR2_X1 U15035 ( .A(n12711), .B(n12710), .ZN(n12712) );
  XOR2_X1 U15036 ( .A(n12713), .B(n12712), .Z(n12714) );
  AOI22_X1 U15037 ( .A1(n14447), .A2(n14656), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12716) );
  NAND2_X1 U15038 ( .A1(n14438), .A2(n14458), .ZN(n12715) );
  OAI211_X1 U15039 ( .C1(n14441), .C2(n14617), .A(n12716), .B(n12715), .ZN(
        n12717) );
  AOI21_X1 U15040 ( .B1(n14980), .B2(n9832), .A(n12717), .ZN(n12718) );
  OAI21_X1 U15041 ( .B1(n12719), .B2(n14456), .A(n12718), .ZN(P1_U3220) );
  XNOR2_X1 U15042 ( .A(n13703), .B(n6801), .ZN(n12768) );
  XNOR2_X1 U15043 ( .A(n12768), .B(n12888), .ZN(n12769) );
  INV_X1 U15044 ( .A(n12730), .ZN(n12720) );
  OAI22_X1 U15045 ( .A1(n12720), .A2(n12725), .B1(n13186), .B2(n12726), .ZN(
        n12722) );
  AOI21_X1 U15046 ( .B1(n12721), .B2(n13170), .A(n12722), .ZN(n12732) );
  AOI21_X1 U15047 ( .B1(n12726), .B2(n13186), .A(n12725), .ZN(n12729) );
  INV_X1 U15048 ( .A(n12722), .ZN(n12724) );
  NAND3_X1 U15049 ( .A1(n12724), .A2(n13197), .A3(n12723), .ZN(n12728) );
  NAND3_X1 U15050 ( .A1(n12726), .A2(n13186), .A3(n12725), .ZN(n12727) );
  OAI211_X1 U15051 ( .C1(n12730), .C2(n12729), .A(n12728), .B(n12727), .ZN(
        n12731) );
  XNOR2_X1 U15052 ( .A(n13711), .B(n6801), .ZN(n12735) );
  XNOR2_X1 U15053 ( .A(n12735), .B(n13152), .ZN(n12800) );
  XNOR2_X1 U15054 ( .A(n13707), .B(n6801), .ZN(n12736) );
  XNOR2_X1 U15055 ( .A(n12736), .B(n13110), .ZN(n12863) );
  INV_X1 U15056 ( .A(n12736), .ZN(n12737) );
  XOR2_X1 U15057 ( .A(n12769), .B(n12770), .Z(n12743) );
  AOI22_X1 U15058 ( .A1(n13133), .A2(n12864), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12739) );
  NAND2_X1 U15059 ( .A1(n13116), .A2(n12882), .ZN(n12738) );
  OAI211_X1 U15060 ( .C1(n13111), .C2(n12867), .A(n12739), .B(n12738), .ZN(
        n12740) );
  AOI21_X1 U15061 ( .B1(n12741), .B2(n12869), .A(n12740), .ZN(n12742) );
  OAI21_X1 U15062 ( .B1(n12743), .B2(n12872), .A(n12742), .ZN(P3_U3154) );
  INV_X1 U15063 ( .A(n12744), .ZN(n12745) );
  AOI21_X1 U15064 ( .B1(n12747), .B2(n12746), .A(n12745), .ZN(n12754) );
  NAND2_X1 U15065 ( .A1(n12882), .A2(n13588), .ZN(n12750) );
  INV_X1 U15066 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n12748) );
  NOR2_X1 U15067 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12748), .ZN(n12926) );
  AOI21_X1 U15068 ( .B1(n13582), .B2(n12878), .A(n12926), .ZN(n12749) );
  OAI211_X1 U15069 ( .C1(n12830), .C2(n12880), .A(n12750), .B(n12749), .ZN(
        n12751) );
  AOI21_X1 U15070 ( .B1(n6828), .B2(n12869), .A(n12751), .ZN(n12753) );
  OAI21_X1 U15071 ( .B1(n12754), .B2(n12872), .A(n12753), .ZN(P3_U3155) );
  XNOR2_X1 U15072 ( .A(n12755), .B(n13186), .ZN(n12760) );
  AOI22_X1 U15073 ( .A1(n13171), .A2(n12878), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12757) );
  NAND2_X1 U15074 ( .A1(n12882), .A2(n13174), .ZN(n12756) );
  OAI211_X1 U15075 ( .C1(n13197), .C2(n12880), .A(n12757), .B(n12756), .ZN(
        n12758) );
  AOI21_X1 U15076 ( .B1(n13175), .B2(n12869), .A(n12758), .ZN(n12759) );
  OAI21_X1 U15077 ( .B1(n12760), .B2(n12872), .A(n12759), .ZN(P3_U3156) );
  OAI211_X1 U15078 ( .C1(n12763), .C2(n12762), .A(n12761), .B(n12874), .ZN(
        n12767) );
  NAND2_X1 U15079 ( .A1(n12889), .A2(n12878), .ZN(n12764) );
  NAND2_X1 U15080 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n13069)
         );
  OAI211_X1 U15081 ( .C1(n13222), .C2(n12880), .A(n12764), .B(n13069), .ZN(
        n12765) );
  AOI21_X1 U15082 ( .B1(n13225), .B2(n12882), .A(n12765), .ZN(n12766) );
  OAI211_X1 U15083 ( .C1(n12885), .C2(n13729), .A(n12767), .B(n12766), .ZN(
        P3_U3159) );
  XNOR2_X1 U15084 ( .A(n13093), .B(n12771), .ZN(n12772) );
  XNOR2_X1 U15085 ( .A(n12773), .B(n12772), .ZN(n12778) );
  AOI22_X1 U15086 ( .A1(n12888), .A2(n12864), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12775) );
  NAND2_X1 U15087 ( .A1(n13097), .A2(n12882), .ZN(n12774) );
  OAI211_X1 U15088 ( .C1(n13094), .C2(n12867), .A(n12775), .B(n12774), .ZN(
        n12776) );
  AOI21_X1 U15089 ( .B1(n13096), .B2(n12869), .A(n12776), .ZN(n12777) );
  OAI21_X1 U15090 ( .B1(n12778), .B2(n12872), .A(n12777), .ZN(P3_U3160) );
  INV_X1 U15091 ( .A(n12779), .ZN(n12780) );
  AOI21_X1 U15092 ( .B1(n12782), .B2(n12781), .A(n12780), .ZN(n12787) );
  AOI22_X1 U15093 ( .A1(n12864), .A2(n12889), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12784) );
  NAND2_X1 U15094 ( .A1(n12882), .A2(n13199), .ZN(n12783) );
  OAI211_X1 U15095 ( .C1(n13197), .C2(n12867), .A(n12784), .B(n12783), .ZN(
        n12785) );
  AOI21_X1 U15096 ( .B1(n13198), .B2(n12869), .A(n12785), .ZN(n12786) );
  OAI21_X1 U15097 ( .B1(n12787), .B2(n12872), .A(n12786), .ZN(P3_U3163) );
  XNOR2_X1 U15098 ( .A(n12788), .B(n12789), .ZN(n12797) );
  AOI21_X1 U15099 ( .B1(n15065), .B2(n12878), .A(n12790), .ZN(n12795) );
  NAND2_X1 U15100 ( .A1(n12882), .A2(n15067), .ZN(n12794) );
  NAND2_X1 U15101 ( .A1(n12791), .A2(n12869), .ZN(n12793) );
  OR2_X1 U15102 ( .A1(n15435), .A2(n12880), .ZN(n12792) );
  NAND4_X1 U15103 ( .A1(n12795), .A2(n12794), .A3(n12793), .A4(n12792), .ZN(
        n12796) );
  AOI21_X1 U15104 ( .B1(n12797), .B2(n12874), .A(n12796), .ZN(n12798) );
  INV_X1 U15105 ( .A(n12798), .ZN(P3_U3164) );
  XOR2_X1 U15106 ( .A(n12800), .B(n12799), .Z(n12806) );
  AOI22_X1 U15107 ( .A1(n13171), .A2(n12864), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12802) );
  NAND2_X1 U15108 ( .A1(n13140), .A2(n12882), .ZN(n12801) );
  OAI211_X1 U15109 ( .C1(n13110), .C2(n12867), .A(n12802), .B(n12801), .ZN(
        n12803) );
  AOI21_X1 U15110 ( .B1(n12804), .B2(n12869), .A(n12803), .ZN(n12805) );
  OAI21_X1 U15111 ( .B1(n12806), .B2(n12872), .A(n12805), .ZN(P3_U3165) );
  XNOR2_X1 U15112 ( .A(n12807), .B(n12808), .ZN(n12813) );
  NAND2_X1 U15113 ( .A1(n12890), .A2(n12878), .ZN(n12809) );
  NAND2_X1 U15114 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12988)
         );
  OAI211_X1 U15115 ( .C1(n13262), .C2(n12880), .A(n12809), .B(n12988), .ZN(
        n12810) );
  AOI21_X1 U15116 ( .B1(n13264), .B2(n12882), .A(n12810), .ZN(n12812) );
  NAND2_X1 U15117 ( .A1(n13676), .A2(n12869), .ZN(n12811) );
  OAI211_X1 U15118 ( .C1(n12813), .C2(n12872), .A(n12812), .B(n12811), .ZN(
        P3_U3166) );
  XNOR2_X1 U15119 ( .A(n12815), .B(n13263), .ZN(n12816) );
  XNOR2_X1 U15120 ( .A(n12814), .B(n12816), .ZN(n12821) );
  AND2_X1 U15121 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13015) );
  AOI21_X1 U15122 ( .B1(n13247), .B2(n12878), .A(n13015), .ZN(n12817) );
  OAI21_X1 U15123 ( .B1(n13560), .B2(n12880), .A(n12817), .ZN(n12819) );
  NOR2_X1 U15124 ( .A1(n13674), .A2(n12885), .ZN(n12818) );
  AOI211_X1 U15125 ( .C1(n13249), .C2(n12882), .A(n12819), .B(n12818), .ZN(
        n12820) );
  OAI21_X1 U15126 ( .B1(n12821), .B2(n12872), .A(n12820), .ZN(P3_U3168) );
  OAI211_X1 U15127 ( .C1(n12824), .C2(n12823), .A(n12822), .B(n12874), .ZN(
        n12828) );
  AOI22_X1 U15128 ( .A1(n13211), .A2(n12878), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12825) );
  OAI21_X1 U15129 ( .B1(n13235), .B2(n12880), .A(n12825), .ZN(n12826) );
  AOI21_X1 U15130 ( .B1(n13215), .B2(n12882), .A(n12826), .ZN(n12827) );
  OAI211_X1 U15131 ( .C1(n13725), .C2(n12885), .A(n12828), .B(n12827), .ZN(
        P3_U3173) );
  XNOR2_X1 U15132 ( .A(n12831), .B(n12830), .ZN(n12832) );
  XNOR2_X1 U15133 ( .A(n12829), .B(n12832), .ZN(n12838) );
  AND2_X1 U15134 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12913) );
  AOI21_X1 U15135 ( .B1(n12833), .B2(n12878), .A(n12913), .ZN(n12834) );
  OAI21_X1 U15136 ( .B1(n13600), .B2(n12880), .A(n12834), .ZN(n12836) );
  NOR2_X1 U15137 ( .A1(n13740), .A2(n12885), .ZN(n12835) );
  AOI211_X1 U15138 ( .C1(n13602), .C2(n12882), .A(n12836), .B(n12835), .ZN(
        n12837) );
  OAI21_X1 U15139 ( .B1(n12838), .B2(n12872), .A(n12837), .ZN(P3_U3174) );
  XNOR2_X1 U15140 ( .A(n12839), .B(n13170), .ZN(n12844) );
  AOI22_X1 U15141 ( .A1(n12864), .A2(n13211), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12841) );
  NAND2_X1 U15142 ( .A1(n12882), .A2(n13188), .ZN(n12840) );
  OAI211_X1 U15143 ( .C1(n13186), .C2(n12867), .A(n12841), .B(n12840), .ZN(
        n12842) );
  AOI21_X1 U15144 ( .B1(n13187), .B2(n12869), .A(n12842), .ZN(n12843) );
  OAI21_X1 U15145 ( .B1(n12844), .B2(n12872), .A(n12843), .ZN(P3_U3175) );
  XNOR2_X1 U15146 ( .A(n12845), .B(n15435), .ZN(n12853) );
  NAND2_X1 U15147 ( .A1(n12882), .A2(n12846), .ZN(n12851) );
  AOI21_X1 U15148 ( .B1(n12891), .B2(n12878), .A(n12847), .ZN(n12850) );
  NAND2_X1 U15149 ( .A1(n12869), .A2(n15085), .ZN(n12849) );
  NAND2_X1 U15150 ( .A1(n12864), .A2(n12892), .ZN(n12848) );
  NAND4_X1 U15151 ( .A1(n12851), .A2(n12850), .A3(n12849), .A4(n12848), .ZN(
        n12852) );
  AOI21_X1 U15152 ( .B1(n12853), .B2(n12874), .A(n12852), .ZN(n12854) );
  INV_X1 U15153 ( .A(n12854), .ZN(P3_U3176) );
  INV_X1 U15154 ( .A(n13242), .ZN(n13733) );
  OAI211_X1 U15155 ( .C1(n12857), .C2(n12856), .A(n12855), .B(n12874), .ZN(
        n12861) );
  AND2_X1 U15156 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n13045) );
  AOI21_X1 U15157 ( .B1(n13212), .B2(n12878), .A(n13045), .ZN(n12858) );
  OAI21_X1 U15158 ( .B1(n13263), .B2(n12880), .A(n12858), .ZN(n12859) );
  AOI21_X1 U15159 ( .B1(n13236), .B2(n12882), .A(n12859), .ZN(n12860) );
  OAI211_X1 U15160 ( .C1(n13733), .C2(n12885), .A(n12861), .B(n12860), .ZN(
        P3_U3178) );
  XOR2_X1 U15161 ( .A(n12863), .B(n12862), .Z(n12873) );
  AOI22_X1 U15162 ( .A1(n13152), .A2(n12864), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12866) );
  NAND2_X1 U15163 ( .A1(n13125), .A2(n12882), .ZN(n12865) );
  OAI211_X1 U15164 ( .C1(n13123), .C2(n12867), .A(n12866), .B(n12865), .ZN(
        n12868) );
  AOI21_X1 U15165 ( .B1(n12870), .B2(n12869), .A(n12868), .ZN(n12871) );
  OAI21_X1 U15166 ( .B1(n12873), .B2(n12872), .A(n12871), .ZN(P3_U3180) );
  INV_X1 U15167 ( .A(n13680), .ZN(n13563) );
  OAI211_X1 U15168 ( .C1(n12877), .C2(n12876), .A(n6601), .B(n12874), .ZN(
        n12884) );
  NAND2_X1 U15169 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12968)
         );
  NAND2_X1 U15170 ( .A1(n13246), .A2(n12878), .ZN(n12879) );
  OAI211_X1 U15171 ( .C1(n13601), .C2(n12880), .A(n12968), .B(n12879), .ZN(
        n12881) );
  AOI21_X1 U15172 ( .B1(n13561), .B2(n12882), .A(n12881), .ZN(n12883) );
  OAI211_X1 U15173 ( .C1(n13563), .C2(n12885), .A(n12884), .B(n12883), .ZN(
        P3_U3181) );
  MUX2_X1 U15174 ( .A(n12886), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12897), .Z(
        P3_U3522) );
  MUX2_X1 U15175 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12887), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U15176 ( .A(n12888), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12897), .Z(
        P3_U3518) );
  MUX2_X1 U15177 ( .A(n13152), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12897), .Z(
        P3_U3516) );
  MUX2_X1 U15178 ( .A(n13171), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12897), .Z(
        P3_U3515) );
  MUX2_X1 U15179 ( .A(n13151), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12897), .Z(
        P3_U3514) );
  MUX2_X1 U15180 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n13170), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U15181 ( .A(n13211), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12897), .Z(
        P3_U3512) );
  MUX2_X1 U15182 ( .A(n12889), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12897), .Z(
        P3_U3511) );
  MUX2_X1 U15183 ( .A(n13212), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12897), .Z(
        P3_U3510) );
  MUX2_X1 U15184 ( .A(n13247), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12897), .Z(
        P3_U3509) );
  MUX2_X1 U15185 ( .A(n12890), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12897), .Z(
        P3_U3508) );
  MUX2_X1 U15186 ( .A(n13246), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12897), .Z(
        P3_U3507) );
  MUX2_X1 U15187 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n15065), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15188 ( .A(n12891), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12897), .Z(
        P3_U3503) );
  MUX2_X1 U15189 ( .A(n12892), .B(P3_DATAO_REG_10__SCAN_IN), .S(n12897), .Z(
        P3_U3501) );
  MUX2_X1 U15190 ( .A(n12893), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12897), .Z(
        P3_U3500) );
  MUX2_X1 U15191 ( .A(n12894), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12897), .Z(
        P3_U3499) );
  MUX2_X1 U15192 ( .A(n15460), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12897), .Z(
        P3_U3498) );
  MUX2_X1 U15193 ( .A(n12895), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12897), .Z(
        P3_U3497) );
  MUX2_X1 U15194 ( .A(n15459), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12897), .Z(
        P3_U3496) );
  MUX2_X1 U15195 ( .A(n15474), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12897), .Z(
        P3_U3495) );
  MUX2_X1 U15196 ( .A(n12896), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12897), .Z(
        P3_U3494) );
  MUX2_X1 U15197 ( .A(n6592), .B(P3_DATAO_REG_2__SCAN_IN), .S(n12897), .Z(
        P3_U3493) );
  MUX2_X1 U15198 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n9975), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15199 ( .A(n15516), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12897), .Z(
        P3_U3491) );
  AND2_X1 U15200 ( .A1(n12898), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12899) );
  INV_X1 U15201 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n13687) );
  AOI21_X1 U15202 ( .B1(n12902), .B2(n13687), .A(n12941), .ZN(n12921) );
  INV_X1 U15203 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13604) );
  OR2_X1 U15204 ( .A1(n6587), .A2(n13604), .ZN(n12904) );
  NAND2_X1 U15205 ( .A1(n6587), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n12903) );
  NAND2_X1 U15206 ( .A1(n12904), .A2(n12903), .ZN(n12933) );
  XOR2_X1 U15207 ( .A(n12932), .B(n12933), .Z(n12908) );
  OAI21_X1 U15208 ( .B1(n12908), .B2(n12907), .A(n12931), .ZN(n12919) );
  AOI21_X1 U15209 ( .B1(n12912), .B2(n13604), .A(n12923), .ZN(n12915) );
  AOI21_X1 U15210 ( .B1(n15417), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12913), 
        .ZN(n12914) );
  OAI21_X1 U15211 ( .B1(n15408), .B2(n12915), .A(n12914), .ZN(n12918) );
  NOR2_X1 U15212 ( .A1(n12916), .A2(n12932), .ZN(n12917) );
  AOI211_X1 U15213 ( .C1(n15422), .C2(n12919), .A(n12918), .B(n12917), .ZN(
        n12920) );
  OAI21_X1 U15214 ( .B1(n12921), .B2(n15407), .A(n12920), .ZN(P3_U3195) );
  INV_X1 U15215 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n13590) );
  MUX2_X1 U15216 ( .A(n13590), .B(P3_REG2_REG_14__SCAN_IN), .S(n12955), .Z(
        n12927) );
  AND2_X1 U15217 ( .A1(n12927), .A2(n12924), .ZN(n12925) );
  OAI21_X1 U15218 ( .B1(n12949), .B2(n12925), .A(n15425), .ZN(n12939) );
  AOI21_X1 U15219 ( .B1(n15417), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12926), 
        .ZN(n12938) );
  OR2_X1 U15220 ( .A1(n6587), .A2(n12927), .ZN(n12930) );
  INV_X1 U15221 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n15078) );
  MUX2_X1 U15222 ( .A(n15078), .B(P3_REG1_REG_14__SCAN_IN), .S(n12955), .Z(
        n12942) );
  INV_X1 U15223 ( .A(n12942), .ZN(n12928) );
  NAND2_X1 U15224 ( .A1(n6587), .A2(n12928), .ZN(n12929) );
  AND2_X1 U15225 ( .A1(n12930), .A2(n12929), .ZN(n12934) );
  NAND2_X1 U15226 ( .A1(n12935), .A2(n12934), .ZN(n12936) );
  NAND3_X1 U15227 ( .A1(n12958), .A2(n15422), .A3(n12936), .ZN(n12937) );
  NAND3_X1 U15228 ( .A1(n12939), .A2(n12938), .A3(n12937), .ZN(n12946) );
  NOR2_X1 U15229 ( .A1(n12943), .A2(n12942), .ZN(n12951) );
  AOI21_X1 U15230 ( .B1(n12943), .B2(n12942), .A(n12951), .ZN(n12944) );
  NOR2_X1 U15231 ( .A1(n12944), .A2(n15407), .ZN(n12945) );
  AOI211_X1 U15232 ( .C1(n15421), .C2(n12947), .A(n12946), .B(n12945), .ZN(
        n12948) );
  INV_X1 U15233 ( .A(n12948), .ZN(P3_U3196) );
  INV_X1 U15234 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12962) );
  AOI21_X1 U15235 ( .B1(n12950), .B2(n12962), .A(n12977), .ZN(n12975) );
  INV_X1 U15236 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12953) );
  AOI21_X1 U15237 ( .B1(n12953), .B2(n12952), .A(n12993), .ZN(n12954) );
  NOR2_X1 U15238 ( .A1(n12954), .A2(n15407), .ZN(n12973) );
  NAND2_X1 U15239 ( .A1(n6587), .A2(n15078), .ZN(n12956) );
  OAI211_X1 U15240 ( .C1(n6587), .C2(P3_REG2_REG_14__SCAN_IN), .A(n12956), .B(
        n12955), .ZN(n12957) );
  NAND2_X1 U15241 ( .A1(n12958), .A2(n12957), .ZN(n12960) );
  NOR2_X1 U15242 ( .A1(n12960), .A2(n12959), .ZN(n12961) );
  OR2_X1 U15243 ( .A1(n6587), .A2(n12962), .ZN(n12964) );
  NAND2_X1 U15244 ( .A1(n6587), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12963) );
  NAND2_X1 U15245 ( .A1(n12964), .A2(n12963), .ZN(n12965) );
  OAI21_X1 U15246 ( .B1(n12966), .B2(n12965), .A(n15422), .ZN(n12967) );
  NOR2_X1 U15247 ( .A1(n12967), .A2(n12983), .ZN(n12972) );
  NAND2_X1 U15248 ( .A1(n15421), .A2(n12992), .ZN(n12969) );
  OAI211_X1 U15249 ( .C1(n12970), .C2(n15414), .A(n12969), .B(n12968), .ZN(
        n12971) );
  NOR3_X1 U15250 ( .A1(n12973), .A2(n12972), .A3(n12971), .ZN(n12974) );
  OAI21_X1 U15251 ( .B1(n12975), .B2(n15408), .A(n12974), .ZN(P3_U3197) );
  NOR2_X1 U15252 ( .A1(n12992), .A2(n12976), .ZN(n12978) );
  INV_X1 U15253 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n13415) );
  AOI22_X1 U15254 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13011), .B1(n13019), 
        .B2(n13415), .ZN(n12979) );
  AOI21_X1 U15255 ( .B1(n12980), .B2(n12979), .A(n13002), .ZN(n13001) );
  INV_X1 U15256 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n12990) );
  OR2_X1 U15257 ( .A1(n6587), .A2(n13415), .ZN(n12982) );
  NAND2_X1 U15258 ( .A1(n6587), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12981) );
  AND2_X1 U15259 ( .A1(n12982), .A2(n12981), .ZN(n13012) );
  XNOR2_X1 U15260 ( .A(n13012), .B(n13019), .ZN(n12986) );
  OAI21_X1 U15261 ( .B1(n12986), .B2(n12985), .A(n13009), .ZN(n12987) );
  NAND2_X1 U15262 ( .A1(n12987), .A2(n15422), .ZN(n12989) );
  OAI211_X1 U15263 ( .C1(n15414), .C2(n12990), .A(n12989), .B(n12988), .ZN(
        n12999) );
  INV_X1 U15264 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12994) );
  AOI22_X1 U15265 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n13011), .B1(n13019), 
        .B2(n12994), .ZN(n12995) );
  AOI21_X1 U15266 ( .B1(n12996), .B2(n12995), .A(n13018), .ZN(n12997) );
  NOR2_X1 U15267 ( .A1(n12997), .A2(n15407), .ZN(n12998) );
  AOI211_X1 U15268 ( .C1(n15421), .C2(n13011), .A(n12999), .B(n12998), .ZN(
        n13000) );
  OAI21_X1 U15269 ( .B1(n13001), .B2(n15408), .A(n13000), .ZN(P3_U3198) );
  XOR2_X1 U15270 ( .A(n13028), .B(n13020), .Z(n13004) );
  INV_X1 U15271 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n13003) );
  AOI21_X1 U15272 ( .B1(n13004), .B2(n13003), .A(n13029), .ZN(n13027) );
  OR2_X1 U15273 ( .A1(n6587), .A2(n13003), .ZN(n13006) );
  NAND2_X1 U15274 ( .A1(n6587), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n13005) );
  NAND2_X1 U15275 ( .A1(n13006), .A2(n13005), .ZN(n13007) );
  AND2_X1 U15276 ( .A1(n13007), .A2(n13020), .ZN(n13042) );
  NOR2_X1 U15277 ( .A1(n13007), .A2(n13020), .ZN(n13008) );
  NOR2_X1 U15278 ( .A1(n13042), .A2(n13008), .ZN(n13014) );
  OAI21_X1 U15279 ( .B1(n13014), .B2(n13013), .A(n15422), .ZN(n13017) );
  AND2_X1 U15280 ( .A1(n13014), .A2(n13013), .ZN(n13041) );
  AOI21_X1 U15281 ( .B1(n15417), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n13015), 
        .ZN(n13016) );
  OAI21_X1 U15282 ( .B1(n13017), .B2(n13041), .A(n13016), .ZN(n13025) );
  INV_X1 U15283 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13022) );
  AOI21_X1 U15284 ( .B1(n13022), .B2(n13021), .A(n13033), .ZN(n13023) );
  NOR2_X1 U15285 ( .A1(n13023), .A2(n15407), .ZN(n13024) );
  AOI211_X1 U15286 ( .C1(n15421), .C2(n7265), .A(n13025), .B(n13024), .ZN(
        n13026) );
  OAI21_X1 U15287 ( .B1(n13027), .B2(n15408), .A(n13026), .ZN(P3_U3199) );
  NOR2_X1 U15288 ( .A1(n7265), .A2(n13028), .ZN(n13030) );
  NAND2_X1 U15289 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n13054), .ZN(n13065) );
  OAI21_X1 U15290 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n13054), .A(n13065), 
        .ZN(n13031) );
  AOI21_X1 U15291 ( .B1(n6704), .B2(n13031), .A(n13066), .ZN(n13052) );
  NOR2_X1 U15292 ( .A1(n7265), .A2(n13032), .ZN(n13034) );
  INV_X1 U15293 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n13669) );
  AOI22_X1 U15294 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n13057), .B1(n13054), 
        .B2(n13669), .ZN(n13035) );
  NOR2_X1 U15295 ( .A1(n13036), .A2(n13035), .ZN(n13053) );
  AOI21_X1 U15296 ( .B1(n13036), .B2(n13035), .A(n13053), .ZN(n13037) );
  NOR2_X1 U15297 ( .A1(n13037), .A2(n15407), .ZN(n13050) );
  NAND2_X1 U15298 ( .A1(n15421), .A2(n13057), .ZN(n13048) );
  INV_X1 U15299 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13238) );
  OR2_X1 U15300 ( .A1(n6587), .A2(n13238), .ZN(n13040) );
  NAND2_X1 U15301 ( .A1(n6587), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n13039) );
  AND2_X1 U15302 ( .A1(n13040), .A2(n13039), .ZN(n13044) );
  XNOR2_X1 U15303 ( .A(n13054), .B(n13056), .ZN(n13043) );
  NAND2_X1 U15304 ( .A1(n13044), .A2(n13043), .ZN(n13059) );
  OAI21_X1 U15305 ( .B1(n13044), .B2(n13043), .A(n13059), .ZN(n13046) );
  AOI21_X1 U15306 ( .B1(n13046), .B2(n15422), .A(n13045), .ZN(n13047) );
  OAI21_X1 U15307 ( .B1(n13052), .B2(n15408), .A(n13051), .ZN(P3_U3200) );
  XNOR2_X1 U15308 ( .A(n13060), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n13062) );
  AOI21_X1 U15309 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(n13054), .A(n13053), 
        .ZN(n13055) );
  NAND2_X1 U15310 ( .A1(n13057), .A2(n13056), .ZN(n13058) );
  NAND2_X1 U15311 ( .A1(n13059), .A2(n13058), .ZN(n13064) );
  INV_X1 U15312 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n13061) );
  MUX2_X1 U15313 ( .A(n13061), .B(P3_REG2_REG_19__SCAN_IN), .S(n13060), .Z(
        n13067) );
  MUX2_X1 U15314 ( .A(n13067), .B(n13062), .S(n6587), .Z(n13063) );
  XNOR2_X1 U15315 ( .A(n13064), .B(n13063), .ZN(n13072) );
  OAI21_X1 U15316 ( .B1(n15414), .B2(n13070), .A(n13069), .ZN(n13071) );
  INV_X1 U15317 ( .A(n13076), .ZN(n13077) );
  NAND2_X1 U15318 ( .A1(n13077), .A2(n15508), .ZN(n13084) );
  OAI21_X1 U15319 ( .B1(n15489), .B2(n13615), .A(n13084), .ZN(n13080) );
  AOI21_X1 U15320 ( .B1(n15489), .B2(P3_REG2_REG_31__SCAN_IN), .A(n13080), 
        .ZN(n13078) );
  OAI21_X1 U15321 ( .B1(n13079), .B2(n13587), .A(n13078), .ZN(P3_U3202) );
  AOI21_X1 U15322 ( .B1(n15489), .B2(P3_REG2_REG_30__SCAN_IN), .A(n13080), 
        .ZN(n13081) );
  OAI21_X1 U15323 ( .B1(n13695), .B2(n13587), .A(n13081), .ZN(P3_U3203) );
  INV_X1 U15324 ( .A(n13082), .ZN(n13089) );
  NAND2_X1 U15325 ( .A1(n15489), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n13083) );
  OAI211_X1 U15326 ( .C1(n13085), .C2(n13587), .A(n13084), .B(n13083), .ZN(
        n13086) );
  AOI21_X1 U15327 ( .B1(n13087), .B2(n15071), .A(n13086), .ZN(n13088) );
  OAI21_X1 U15328 ( .B1(n13089), .B2(n15489), .A(n13088), .ZN(P3_U3204) );
  INV_X1 U15329 ( .A(n13621), .ZN(n13101) );
  OAI22_X1 U15330 ( .A1(n13094), .A2(n15494), .B1(n13123), .B2(n15492), .ZN(
        n13095) );
  AOI22_X1 U15331 ( .A1(n13097), .A2(n15508), .B1(n15489), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n13098) );
  OAI21_X1 U15332 ( .B1(n13699), .B2(n13587), .A(n13098), .ZN(n13099) );
  AOI21_X1 U15333 ( .B1(n13620), .B2(n15530), .A(n13099), .ZN(n13100) );
  OAI21_X1 U15334 ( .B1(n13101), .B2(n13606), .A(n13100), .ZN(P3_U3205) );
  INV_X1 U15335 ( .A(n13629), .ZN(n13104) );
  AOI21_X1 U15336 ( .B1(n13104), .B2(n13103), .A(n13102), .ZN(n13105) );
  NOR2_X1 U15337 ( .A1(n13106), .A2(n13105), .ZN(n13115) );
  INV_X1 U15338 ( .A(n15502), .ZN(n15481) );
  OAI21_X1 U15339 ( .B1(n13109), .B2(n13108), .A(n13107), .ZN(n13113) );
  OAI22_X1 U15340 ( .A1(n13111), .A2(n15494), .B1(n13110), .B2(n15492), .ZN(
        n13112) );
  AOI21_X1 U15341 ( .B1(n13113), .B2(n15513), .A(n13112), .ZN(n13114) );
  OAI21_X1 U15342 ( .B1(n13115), .B2(n15481), .A(n13114), .ZN(n13624) );
  INV_X1 U15343 ( .A(n13624), .ZN(n13120) );
  INV_X1 U15344 ( .A(n13115), .ZN(n13625) );
  AOI22_X1 U15345 ( .A1(n13116), .A2(n15508), .B1(n15489), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n13117) );
  OAI21_X1 U15346 ( .B1(n13703), .B2(n13587), .A(n13117), .ZN(n13118) );
  AOI21_X1 U15347 ( .B1(n13625), .B2(n15444), .A(n13118), .ZN(n13119) );
  OAI21_X1 U15348 ( .B1(n13120), .B2(n15489), .A(n13119), .ZN(P3_U3206) );
  XNOR2_X1 U15349 ( .A(n13121), .B(n13127), .ZN(n13124) );
  OAI222_X1 U15350 ( .A1(n13124), .A2(n15497), .B1(n15494), .B2(n13123), .C1(
        n15492), .C2(n13122), .ZN(n13630) );
  AOI22_X1 U15351 ( .A1(n13125), .A2(n15508), .B1(n15489), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n13126) );
  OAI21_X1 U15352 ( .B1(n13707), .B2(n13587), .A(n13126), .ZN(n13130) );
  AND2_X1 U15353 ( .A1(n6591), .A2(n13127), .ZN(n13628) );
  NOR3_X1 U15354 ( .A1(n13629), .A2(n13628), .A3(n13606), .ZN(n13129) );
  AOI211_X1 U15355 ( .C1(n15530), .C2(n13630), .A(n13130), .B(n13129), .ZN(
        n13131) );
  INV_X1 U15356 ( .A(n13131), .ZN(P3_U3207) );
  XOR2_X1 U15357 ( .A(n13135), .B(n13132), .Z(n13139) );
  AOI22_X1 U15358 ( .A1(n13133), .A2(n15517), .B1(n15515), .B2(n13171), .ZN(
        n13138) );
  OAI211_X1 U15359 ( .C1(n13136), .C2(n13135), .A(n13134), .B(n15513), .ZN(
        n13137) );
  OAI211_X1 U15360 ( .C1(n13139), .C2(n15481), .A(n13138), .B(n13137), .ZN(
        n13634) );
  INV_X1 U15361 ( .A(n13634), .ZN(n13144) );
  INV_X1 U15362 ( .A(n13139), .ZN(n13635) );
  AOI22_X1 U15363 ( .A1(n13140), .A2(n15508), .B1(n15489), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n13141) );
  OAI21_X1 U15364 ( .B1(n13711), .B2(n13587), .A(n13141), .ZN(n13142) );
  AOI21_X1 U15365 ( .B1(n13635), .B2(n15444), .A(n13142), .ZN(n13143) );
  OAI21_X1 U15366 ( .B1(n13144), .B2(n15489), .A(n13143), .ZN(P3_U3208) );
  NAND2_X1 U15367 ( .A1(n13145), .A2(n13164), .ZN(n13166) );
  AND2_X1 U15368 ( .A1(n13166), .A2(n13146), .ZN(n13150) );
  AOI21_X1 U15369 ( .B1(n13166), .B2(n13148), .A(n13147), .ZN(n13149) );
  NAND2_X1 U15370 ( .A1(n13638), .A2(n15502), .ZN(n13158) );
  AOI22_X1 U15371 ( .A1(n13152), .A2(n15517), .B1(n15515), .B2(n13151), .ZN(
        n13157) );
  OAI211_X1 U15372 ( .C1(n13155), .C2(n13154), .A(n13153), .B(n15513), .ZN(
        n13156) );
  NAND3_X1 U15373 ( .A1(n13158), .A2(n13157), .A3(n13156), .ZN(n13642) );
  INV_X1 U15374 ( .A(n13642), .ZN(n13163) );
  AOI22_X1 U15375 ( .A1(n13159), .A2(n15508), .B1(P3_REG2_REG_24__SCAN_IN), 
        .B2(n15489), .ZN(n13160) );
  OAI21_X1 U15376 ( .B1(n13640), .B2(n13587), .A(n13160), .ZN(n13161) );
  AOI21_X1 U15377 ( .B1(n13638), .B2(n15444), .A(n13161), .ZN(n13162) );
  OAI21_X1 U15378 ( .B1(n13163), .B2(n15489), .A(n13162), .ZN(P3_U3209) );
  OR2_X1 U15379 ( .A1(n13145), .A2(n13164), .ZN(n13165) );
  NAND2_X1 U15380 ( .A1(n13166), .A2(n13165), .ZN(n13645) );
  OAI211_X1 U15381 ( .C1(n13169), .C2(n13168), .A(n13167), .B(n15513), .ZN(
        n13173) );
  AOI22_X1 U15382 ( .A1(n13171), .A2(n15517), .B1(n15515), .B2(n13170), .ZN(
        n13172) );
  OAI211_X1 U15383 ( .C1(n15481), .C2(n13645), .A(n13173), .B(n13172), .ZN(
        n13647) );
  INV_X1 U15384 ( .A(n15444), .ZN(n13178) );
  AOI22_X1 U15385 ( .A1(n15489), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n13174), 
        .B2(n15508), .ZN(n13177) );
  INV_X1 U15386 ( .A(n13587), .ZN(n13611) );
  NAND2_X1 U15387 ( .A1(n13175), .A2(n13611), .ZN(n13176) );
  OAI211_X1 U15388 ( .C1(n13645), .C2(n13178), .A(n13177), .B(n13176), .ZN(
        n13179) );
  AOI21_X1 U15389 ( .B1(n13647), .B2(n15530), .A(n13179), .ZN(n13180) );
  INV_X1 U15390 ( .A(n13180), .ZN(P3_U3210) );
  XNOR2_X1 U15391 ( .A(n13181), .B(n13182), .ZN(n13649) );
  INV_X1 U15392 ( .A(n13649), .ZN(n13192) );
  XNOR2_X1 U15393 ( .A(n13183), .B(n13182), .ZN(n13184) );
  OAI222_X1 U15394 ( .A1(n15494), .A2(n13186), .B1(n15492), .B2(n13185), .C1(
        n13184), .C2(n15497), .ZN(n13648) );
  INV_X1 U15395 ( .A(n13187), .ZN(n13717) );
  AOI22_X1 U15396 ( .A1(n15489), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15508), 
        .B2(n13188), .ZN(n13189) );
  OAI21_X1 U15397 ( .B1(n13717), .B2(n13587), .A(n13189), .ZN(n13190) );
  AOI21_X1 U15398 ( .B1(n13648), .B2(n15530), .A(n13190), .ZN(n13191) );
  OAI21_X1 U15399 ( .B1(n13192), .B2(n13606), .A(n13191), .ZN(P3_U3211) );
  XNOR2_X1 U15400 ( .A(n13193), .B(n13194), .ZN(n13653) );
  INV_X1 U15401 ( .A(n13653), .ZN(n13203) );
  XNOR2_X1 U15402 ( .A(n13195), .B(n13194), .ZN(n13196) );
  OAI222_X1 U15403 ( .A1(n15494), .A2(n13197), .B1(n15492), .B2(n13223), .C1(
        n15497), .C2(n13196), .ZN(n13652) );
  INV_X1 U15404 ( .A(n13198), .ZN(n13721) );
  AOI22_X1 U15405 ( .A1(n15489), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15508), 
        .B2(n13199), .ZN(n13200) );
  OAI21_X1 U15406 ( .B1(n13721), .B2(n13587), .A(n13200), .ZN(n13201) );
  AOI21_X1 U15407 ( .B1(n13652), .B2(n15530), .A(n13201), .ZN(n13202) );
  OAI21_X1 U15408 ( .B1(n13606), .B2(n13203), .A(n13202), .ZN(P3_U3212) );
  NAND2_X1 U15409 ( .A1(n13204), .A2(n8287), .ZN(n13205) );
  NAND2_X1 U15410 ( .A1(n13206), .A2(n13205), .ZN(n13656) );
  NAND2_X1 U15411 ( .A1(n13208), .A2(n13207), .ZN(n13209) );
  NAND3_X1 U15412 ( .A1(n13210), .A2(n15513), .A3(n13209), .ZN(n13214) );
  AOI22_X1 U15413 ( .A1(n15515), .A2(n13212), .B1(n13211), .B2(n15517), .ZN(
        n13213) );
  INV_X1 U15414 ( .A(n13657), .ZN(n13218) );
  AOI22_X1 U15415 ( .A1(n15489), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15508), 
        .B2(n13215), .ZN(n13216) );
  OAI21_X1 U15416 ( .B1(n13725), .B2(n13587), .A(n13216), .ZN(n13217) );
  AOI21_X1 U15417 ( .B1(n13218), .B2(n15530), .A(n13217), .ZN(n13219) );
  OAI21_X1 U15418 ( .B1(n13606), .B2(n13656), .A(n13219), .ZN(P3_U3213) );
  XNOR2_X1 U15419 ( .A(n13220), .B(n6618), .ZN(n13221) );
  OAI222_X1 U15420 ( .A1(n15494), .A2(n13223), .B1(n15492), .B2(n13222), .C1(
        n15497), .C2(n13221), .ZN(n13661) );
  INV_X1 U15421 ( .A(n13661), .ZN(n13229) );
  OAI21_X1 U15422 ( .B1(n6717), .B2(n6618), .A(n13224), .ZN(n13662) );
  AOI22_X1 U15423 ( .A1(n15489), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15508), 
        .B2(n13225), .ZN(n13226) );
  OAI21_X1 U15424 ( .B1(n13729), .B2(n13587), .A(n13226), .ZN(n13227) );
  AOI21_X1 U15425 ( .B1(n13662), .B2(n15071), .A(n13227), .ZN(n13228) );
  OAI21_X1 U15426 ( .B1(n13229), .B2(n15489), .A(n13228), .ZN(P3_U3214) );
  INV_X1 U15427 ( .A(n13230), .ZN(n13231) );
  AOI21_X1 U15428 ( .B1(n13233), .B2(n13232), .A(n13231), .ZN(n13234) );
  OAI222_X1 U15429 ( .A1(n15494), .A2(n13235), .B1(n15492), .B2(n13263), .C1(
        n15497), .C2(n13234), .ZN(n13666) );
  INV_X1 U15430 ( .A(n13666), .ZN(n13244) );
  INV_X1 U15431 ( .A(n13236), .ZN(n13237) );
  OAI22_X1 U15432 ( .A1(n15530), .A2(n13238), .B1(n13237), .B2(n15525), .ZN(
        n13241) );
  AND2_X1 U15433 ( .A1(n13239), .A2(n8282), .ZN(n13665) );
  NOR3_X1 U15434 ( .A1(n8075), .A2(n13665), .A3(n13606), .ZN(n13240) );
  AOI211_X1 U15435 ( .C1(n13611), .C2(n13242), .A(n13241), .B(n13240), .ZN(
        n13243) );
  OAI21_X1 U15436 ( .B1(n13244), .B2(n15489), .A(n13243), .ZN(P3_U3215) );
  XNOR2_X1 U15437 ( .A(n13245), .B(n13254), .ZN(n13248) );
  AOI222_X1 U15438 ( .A1(n15513), .A2(n13248), .B1(n13247), .B2(n15517), .C1(
        n13246), .C2(n15515), .ZN(n13673) );
  INV_X1 U15439 ( .A(n13674), .ZN(n13252) );
  INV_X1 U15440 ( .A(n13249), .ZN(n13250) );
  OAI22_X1 U15441 ( .A1(n15530), .A2(n13003), .B1(n13250), .B2(n15525), .ZN(
        n13251) );
  AOI21_X1 U15442 ( .B1(n13252), .B2(n13611), .A(n13251), .ZN(n13256) );
  XNOR2_X1 U15443 ( .A(n13253), .B(n13254), .ZN(n13671) );
  NAND2_X1 U15444 ( .A1(n13671), .A2(n15071), .ZN(n13255) );
  OAI211_X1 U15445 ( .C1(n13673), .C2(n15489), .A(n13256), .B(n13255), .ZN(
        P3_U3216) );
  XNOR2_X1 U15446 ( .A(n13257), .B(n13258), .ZN(n13678) );
  XNOR2_X1 U15447 ( .A(n13260), .B(n13259), .ZN(n13261) );
  OAI222_X1 U15448 ( .A1(n15494), .A2(n13263), .B1(n15492), .B2(n13262), .C1(
        n13261), .C2(n15497), .ZN(n13675) );
  INV_X1 U15449 ( .A(n13676), .ZN(n13266) );
  AOI22_X1 U15450 ( .A1(n15489), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15508), 
        .B2(n13264), .ZN(n13265) );
  OAI21_X1 U15451 ( .B1(n13266), .B2(n13587), .A(n13265), .ZN(n13267) );
  AOI21_X1 U15452 ( .B1(n13675), .B2(n15530), .A(n13267), .ZN(n13268) );
  OAI21_X1 U15453 ( .B1(n13678), .B2(n13606), .A(n13268), .ZN(P3_U3217) );
  NAND2_X1 U15454 ( .A1(keyinput54), .A2(keyinput91), .ZN(n13269) );
  NOR3_X1 U15455 ( .A1(keyinput82), .A2(keyinput68), .A3(n13269), .ZN(n13270)
         );
  NAND3_X1 U15456 ( .A1(keyinput107), .A2(keyinput5), .A3(n13270), .ZN(n13281)
         );
  NAND4_X1 U15457 ( .A1(keyinput62), .A2(keyinput94), .A3(keyinput98), .A4(
        keyinput78), .ZN(n13271) );
  NOR3_X1 U15458 ( .A1(keyinput31), .A2(keyinput52), .A3(n13271), .ZN(n13279)
         );
  NOR4_X1 U15459 ( .A1(keyinput83), .A2(keyinput108), .A3(keyinput25), .A4(
        keyinput41), .ZN(n13272) );
  NAND3_X1 U15460 ( .A1(keyinput23), .A2(keyinput56), .A3(n13272), .ZN(n13277)
         );
  INV_X1 U15461 ( .A(keyinput27), .ZN(n13273) );
  NAND4_X1 U15462 ( .A1(keyinput26), .A2(keyinput30), .A3(keyinput86), .A4(
        n13273), .ZN(n13276) );
  NOR3_X1 U15463 ( .A1(keyinput42), .A2(keyinput69), .A3(keyinput118), .ZN(
        n13274) );
  NAND2_X1 U15464 ( .A1(keyinput3), .A2(n13274), .ZN(n13275) );
  NOR4_X1 U15465 ( .A1(keyinput71), .A2(n13277), .A3(n13276), .A4(n13275), 
        .ZN(n13278) );
  NAND4_X1 U15466 ( .A1(keyinput33), .A2(keyinput43), .A3(n13279), .A4(n13278), 
        .ZN(n13280) );
  NOR4_X1 U15467 ( .A1(keyinput121), .A2(keyinput39), .A3(n13281), .A4(n13280), 
        .ZN(n13332) );
  INV_X1 U15468 ( .A(keyinput125), .ZN(n13282) );
  NAND4_X1 U15469 ( .A1(keyinput6), .A2(keyinput65), .A3(keyinput110), .A4(
        n13282), .ZN(n13289) );
  NOR2_X1 U15470 ( .A1(keyinput99), .A2(keyinput17), .ZN(n13283) );
  NAND3_X1 U15471 ( .A1(keyinput88), .A2(keyinput77), .A3(n13283), .ZN(n13288)
         );
  NOR2_X1 U15472 ( .A1(keyinput21), .A2(keyinput81), .ZN(n13284) );
  NAND3_X1 U15473 ( .A1(keyinput57), .A2(keyinput36), .A3(n13284), .ZN(n13287)
         );
  INV_X1 U15474 ( .A(keyinput120), .ZN(n13285) );
  NAND4_X1 U15475 ( .A1(keyinput9), .A2(keyinput19), .A3(keyinput7), .A4(
        n13285), .ZN(n13286) );
  NOR4_X1 U15476 ( .A1(n13289), .A2(n13288), .A3(n13287), .A4(n13286), .ZN(
        n13331) );
  NOR2_X1 U15477 ( .A1(keyinput67), .A2(keyinput37), .ZN(n13290) );
  NAND3_X1 U15478 ( .A1(keyinput29), .A2(keyinput116), .A3(n13290), .ZN(n13296) );
  INV_X1 U15479 ( .A(keyinput44), .ZN(n13291) );
  NAND4_X1 U15480 ( .A1(keyinput92), .A2(keyinput127), .A3(keyinput106), .A4(
        n13291), .ZN(n13295) );
  INV_X1 U15481 ( .A(keyinput115), .ZN(n13292) );
  NAND4_X1 U15482 ( .A1(keyinput97), .A2(keyinput113), .A3(keyinput74), .A4(
        n13292), .ZN(n13294) );
  OR4_X1 U15483 ( .A1(keyinput105), .A2(keyinput18), .A3(keyinput73), .A4(
        keyinput72), .ZN(n13293) );
  NOR4_X1 U15484 ( .A1(n13296), .A2(n13295), .A3(n13294), .A4(n13293), .ZN(
        n13330) );
  NOR2_X1 U15485 ( .A1(keyinput85), .A2(keyinput45), .ZN(n13297) );
  NAND3_X1 U15486 ( .A1(keyinput93), .A2(keyinput109), .A3(n13297), .ZN(n13328) );
  NOR2_X1 U15487 ( .A1(keyinput58), .A2(keyinput87), .ZN(n13298) );
  NAND3_X1 U15488 ( .A1(keyinput95), .A2(keyinput89), .A3(n13298), .ZN(n13327)
         );
  NAND2_X1 U15489 ( .A1(keyinput15), .A2(keyinput24), .ZN(n13299) );
  NOR3_X1 U15490 ( .A1(keyinput4), .A2(keyinput34), .A3(n13299), .ZN(n13309)
         );
  NOR4_X1 U15491 ( .A1(keyinput96), .A2(keyinput104), .A3(keyinput53), .A4(
        keyinput40), .ZN(n13308) );
  NOR2_X1 U15492 ( .A1(keyinput63), .A2(keyinput84), .ZN(n13300) );
  NAND3_X1 U15493 ( .A1(keyinput66), .A2(keyinput101), .A3(n13300), .ZN(n13306) );
  INV_X1 U15494 ( .A(keyinput111), .ZN(n13301) );
  NAND4_X1 U15495 ( .A1(keyinput51), .A2(keyinput123), .A3(keyinput20), .A4(
        n13301), .ZN(n13305) );
  NAND4_X1 U15496 ( .A1(keyinput49), .A2(keyinput80), .A3(keyinput11), .A4(
        keyinput50), .ZN(n13304) );
  NOR2_X1 U15497 ( .A1(keyinput8), .A2(keyinput119), .ZN(n13302) );
  NAND3_X1 U15498 ( .A1(keyinput100), .A2(keyinput117), .A3(n13302), .ZN(
        n13303) );
  NOR4_X1 U15499 ( .A1(n13306), .A2(n13305), .A3(n13304), .A4(n13303), .ZN(
        n13307) );
  NAND3_X1 U15500 ( .A1(n13309), .A2(n13308), .A3(n13307), .ZN(n13326) );
  NOR2_X1 U15501 ( .A1(keyinput114), .A2(keyinput46), .ZN(n13310) );
  NAND3_X1 U15502 ( .A1(keyinput47), .A2(keyinput14), .A3(n13310), .ZN(n13311)
         );
  NOR3_X1 U15503 ( .A1(keyinput126), .A2(keyinput0), .A3(n13311), .ZN(n13324)
         );
  NAND2_X1 U15504 ( .A1(keyinput12), .A2(keyinput70), .ZN(n13312) );
  NOR3_X1 U15505 ( .A1(keyinput16), .A2(keyinput1), .A3(n13312), .ZN(n13313)
         );
  NAND3_X1 U15506 ( .A1(keyinput90), .A2(keyinput13), .A3(n13313), .ZN(n13322)
         );
  NAND2_X1 U15507 ( .A1(keyinput32), .A2(keyinput64), .ZN(n13314) );
  NOR3_X1 U15508 ( .A1(keyinput122), .A2(keyinput102), .A3(n13314), .ZN(n13320) );
  NAND2_X1 U15509 ( .A1(keyinput124), .A2(keyinput103), .ZN(n13315) );
  NOR3_X1 U15510 ( .A1(keyinput75), .A2(keyinput59), .A3(n13315), .ZN(n13319)
         );
  NOR4_X1 U15511 ( .A1(keyinput76), .A2(keyinput28), .A3(keyinput38), .A4(
        keyinput48), .ZN(n13318) );
  INV_X1 U15512 ( .A(keyinput10), .ZN(n13316) );
  NOR4_X1 U15513 ( .A1(keyinput2), .A2(keyinput55), .A3(keyinput61), .A4(
        n13316), .ZN(n13317) );
  NAND4_X1 U15514 ( .A1(n13320), .A2(n13319), .A3(n13318), .A4(n13317), .ZN(
        n13321) );
  NOR4_X1 U15515 ( .A1(keyinput79), .A2(keyinput35), .A3(n13322), .A4(n13321), 
        .ZN(n13323) );
  NAND4_X1 U15516 ( .A1(keyinput112), .A2(keyinput22), .A3(n13324), .A4(n13323), .ZN(n13325) );
  NOR4_X1 U15517 ( .A1(n13328), .A2(n13327), .A3(n13326), .A4(n13325), .ZN(
        n13329) );
  NAND4_X1 U15518 ( .A1(n13332), .A2(n13331), .A3(n13330), .A4(n13329), .ZN(
        n13333) );
  NAND2_X1 U15519 ( .A1(n13333), .A2(keyinput60), .ZN(n13334) );
  MUX2_X1 U15520 ( .A(keyinput60), .B(n13334), .S(P1_IR_REG_27__SCAN_IN), .Z(
        n13555) );
  AOI22_X1 U15521 ( .A1(n13336), .A2(keyinput18), .B1(n15028), .B2(keyinput73), 
        .ZN(n13335) );
  OAI221_X1 U15522 ( .B1(n13336), .B2(keyinput18), .C1(n15028), .C2(keyinput73), .A(n13335), .ZN(n13345) );
  AOI22_X1 U15523 ( .A1(n13339), .A2(keyinput72), .B1(n13338), .B2(keyinput115), .ZN(n13337) );
  OAI221_X1 U15524 ( .B1(n13339), .B2(keyinput72), .C1(n13338), .C2(
        keyinput115), .A(n13337), .ZN(n13344) );
  AOI22_X1 U15525 ( .A1(n15487), .A2(keyinput97), .B1(keyinput113), .B2(n13821), .ZN(n13340) );
  OAI221_X1 U15526 ( .B1(n15487), .B2(keyinput97), .C1(n13821), .C2(
        keyinput113), .A(n13340), .ZN(n13343) );
  INV_X1 U15527 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15341) );
  AOI22_X1 U15528 ( .A1(n15025), .A2(keyinput74), .B1(keyinput99), .B2(n15341), 
        .ZN(n13341) );
  OAI221_X1 U15529 ( .B1(n15025), .B2(keyinput74), .C1(n15341), .C2(keyinput99), .A(n13341), .ZN(n13342) );
  NOR4_X1 U15530 ( .A1(n13345), .A2(n13344), .A3(n13343), .A4(n13342), .ZN(
        n13360) );
  INV_X1 U15531 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U15532 ( .A1(n13663), .A2(keyinput75), .B1(n13347), .B2(keyinput124), .ZN(n13346) );
  OAI221_X1 U15533 ( .B1(n13663), .B2(keyinput75), .C1(n13347), .C2(
        keyinput124), .A(n13346), .ZN(n13358) );
  AOI22_X1 U15534 ( .A1(n10848), .A2(keyinput59), .B1(n13349), .B2(keyinput64), 
        .ZN(n13348) );
  OAI221_X1 U15535 ( .B1(n10848), .B2(keyinput59), .C1(n13349), .C2(keyinput64), .A(n13348), .ZN(n13357) );
  AOI22_X1 U15536 ( .A1(n13352), .A2(keyinput122), .B1(n13351), .B2(keyinput32), .ZN(n13350) );
  OAI221_X1 U15537 ( .B1(n13352), .B2(keyinput122), .C1(n13351), .C2(
        keyinput32), .A(n13350), .ZN(n13356) );
  AOI22_X1 U15538 ( .A1(n13354), .A2(keyinput102), .B1(n15220), .B2(
        keyinput114), .ZN(n13353) );
  OAI221_X1 U15539 ( .B1(n13354), .B2(keyinput102), .C1(n15220), .C2(
        keyinput114), .A(n13353), .ZN(n13355) );
  NOR4_X1 U15540 ( .A1(n13358), .A2(n13357), .A3(n13356), .A4(n13355), .ZN(
        n13359) );
  NAND2_X1 U15541 ( .A1(n13360), .A2(n13359), .ZN(n13554) );
  INV_X1 U15542 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n13363) );
  INV_X1 U15543 ( .A(keyinput37), .ZN(n13362) );
  AOI22_X1 U15544 ( .A1(n13363), .A2(keyinput67), .B1(P3_DATAO_REG_29__SCAN_IN), .B2(n13362), .ZN(n13361) );
  OAI221_X1 U15545 ( .B1(n13363), .B2(keyinput67), .C1(n13362), .C2(
        P3_DATAO_REG_29__SCAN_IN), .A(n13361), .ZN(n13395) );
  AOI22_X1 U15546 ( .A1(n13366), .A2(keyinput9), .B1(n13365), .B2(keyinput7), 
        .ZN(n13364) );
  OAI221_X1 U15547 ( .B1(n13366), .B2(keyinput9), .C1(n13365), .C2(keyinput7), 
        .A(n13364), .ZN(n13368) );
  XOR2_X1 U15548 ( .A(keyinput108), .B(P3_DATAO_REG_28__SCAN_IN), .Z(n13367)
         );
  NOR2_X1 U15549 ( .A1(n13368), .A2(n13367), .ZN(n13378) );
  XNOR2_X1 U15550 ( .A(keyinput77), .B(n15598), .ZN(n13371) );
  INV_X1 U15551 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n13369) );
  XNOR2_X1 U15552 ( .A(keyinput26), .B(n13369), .ZN(n13370) );
  NOR2_X1 U15553 ( .A1(n13371), .A2(n13370), .ZN(n13377) );
  AOI22_X1 U15554 ( .A1(n13374), .A2(keyinput39), .B1(n13373), .B2(keyinput107), .ZN(n13372) );
  OAI221_X1 U15555 ( .B1(n13374), .B2(keyinput39), .C1(n13373), .C2(
        keyinput107), .A(n13372), .ZN(n13375) );
  INV_X1 U15556 ( .A(n13375), .ZN(n13376) );
  NAND3_X1 U15557 ( .A1(n13378), .A2(n13377), .A3(n13376), .ZN(n13394) );
  INV_X1 U15558 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15575) );
  AOI22_X1 U15559 ( .A1(n9461), .A2(keyinput71), .B1(n15575), .B2(keyinput81), 
        .ZN(n13379) );
  OAI221_X1 U15560 ( .B1(n9461), .B2(keyinput71), .C1(n15575), .C2(keyinput81), 
        .A(n13379), .ZN(n13389) );
  INV_X1 U15561 ( .A(keyinput65), .ZN(n13381) );
  AOI22_X1 U15562 ( .A1(n15218), .A2(keyinput17), .B1(P3_DATAO_REG_11__SCAN_IN), .B2(n13381), .ZN(n13380) );
  OAI221_X1 U15563 ( .B1(n15218), .B2(keyinput17), .C1(n13381), .C2(
        P3_DATAO_REG_11__SCAN_IN), .A(n13380), .ZN(n13388) );
  INV_X1 U15564 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15241) );
  INV_X1 U15565 ( .A(keyinput105), .ZN(n13383) );
  AOI22_X1 U15566 ( .A1(n15241), .A2(keyinput116), .B1(P3_ADDR_REG_15__SCAN_IN), .B2(n13383), .ZN(n13382) );
  OAI221_X1 U15567 ( .B1(n15241), .B2(keyinput116), .C1(n13383), .C2(
        P3_ADDR_REG_15__SCAN_IN), .A(n13382), .ZN(n13387) );
  INV_X1 U15568 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n13385) );
  INV_X1 U15569 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15538) );
  AOI22_X1 U15570 ( .A1(n13385), .A2(keyinput120), .B1(n15538), .B2(keyinput57), .ZN(n13384) );
  OAI221_X1 U15571 ( .B1(n13385), .B2(keyinput120), .C1(n15538), .C2(
        keyinput57), .A(n13384), .ZN(n13386) );
  OR4_X1 U15572 ( .A1(n13389), .A2(n13388), .A3(n13387), .A4(n13386), .ZN(
        n13393) );
  AOI22_X1 U15573 ( .A1(n15587), .A2(keyinput83), .B1(n13391), .B2(keyinput25), 
        .ZN(n13390) );
  OAI221_X1 U15574 ( .B1(n15587), .B2(keyinput83), .C1(n13391), .C2(keyinput25), .A(n13390), .ZN(n13392) );
  NOR4_X1 U15575 ( .A1(n13395), .A2(n13394), .A3(n13393), .A4(n13392), .ZN(
        n13471) );
  INV_X1 U15576 ( .A(keyinput55), .ZN(n13397) );
  AOI22_X1 U15577 ( .A1(n13398), .A2(keyinput10), .B1(P3_ADDR_REG_1__SCAN_IN), 
        .B2(n13397), .ZN(n13396) );
  OAI221_X1 U15578 ( .B1(n13398), .B2(keyinput10), .C1(n13397), .C2(
        P3_ADDR_REG_1__SCAN_IN), .A(n13396), .ZN(n13409) );
  INV_X1 U15579 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15165) );
  INV_X1 U15580 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15342) );
  AOI22_X1 U15581 ( .A1(n15165), .A2(keyinput61), .B1(n15342), .B2(keyinput76), 
        .ZN(n13399) );
  OAI221_X1 U15582 ( .B1(n15165), .B2(keyinput61), .C1(n15342), .C2(keyinput76), .A(n13399), .ZN(n13408) );
  AOI22_X1 U15583 ( .A1(n13402), .A2(keyinput28), .B1(keyinput38), .B2(n13401), 
        .ZN(n13400) );
  OAI221_X1 U15584 ( .B1(n13402), .B2(keyinput28), .C1(n13401), .C2(keyinput38), .A(n13400), .ZN(n13407) );
  AOI22_X1 U15585 ( .A1(n13405), .A2(keyinput48), .B1(n13404), .B2(keyinput16), 
        .ZN(n13403) );
  OAI221_X1 U15586 ( .B1(n13405), .B2(keyinput48), .C1(n13404), .C2(keyinput16), .A(n13403), .ZN(n13406) );
  NOR4_X1 U15587 ( .A1(n13409), .A2(n13408), .A3(n13407), .A4(n13406), .ZN(
        n13470) );
  INV_X1 U15588 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n15163) );
  OAI22_X1 U15589 ( .A1(n15163), .A2(keyinput118), .B1(n14263), .B2(keyinput42), .ZN(n13410) );
  AOI221_X1 U15590 ( .B1(n15163), .B2(keyinput118), .C1(keyinput42), .C2(
        n14263), .A(n13410), .ZN(n13469) );
  INV_X1 U15591 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13413) );
  INV_X1 U15592 ( .A(keyinput45), .ZN(n13412) );
  AOI22_X1 U15593 ( .A1(n13413), .A2(keyinput93), .B1(P2_ADDR_REG_7__SCAN_IN), 
        .B2(n13412), .ZN(n13411) );
  OAI221_X1 U15594 ( .B1(n13413), .B2(keyinput93), .C1(n13412), .C2(
        P2_ADDR_REG_7__SCAN_IN), .A(n13411), .ZN(n13423) );
  AOI22_X1 U15595 ( .A1(n10738), .A2(keyinput87), .B1(n13415), .B2(keyinput58), 
        .ZN(n13414) );
  OAI221_X1 U15596 ( .B1(n10738), .B2(keyinput87), .C1(n13415), .C2(keyinput58), .A(n13414), .ZN(n13422) );
  AOI22_X1 U15597 ( .A1(n7756), .A2(keyinput109), .B1(keyinput123), .B2(n13417), .ZN(n13416) );
  OAI221_X1 U15598 ( .B1(n7756), .B2(keyinput109), .C1(n13417), .C2(
        keyinput123), .A(n13416), .ZN(n13421) );
  XNOR2_X1 U15599 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput89), .ZN(n13419)
         );
  XNOR2_X1 U15600 ( .A(P1_REG0_REG_31__SCAN_IN), .B(keyinput85), .ZN(n13418)
         );
  NAND2_X1 U15601 ( .A1(n13419), .A2(n13418), .ZN(n13420) );
  NOR4_X1 U15602 ( .A1(n13423), .A2(n13422), .A3(n13421), .A4(n13420), .ZN(
        n13467) );
  INV_X1 U15603 ( .A(keyinput40), .ZN(n13425) );
  AOI22_X1 U15604 ( .A1(n13426), .A2(keyinput34), .B1(P1_ADDR_REG_12__SCAN_IN), 
        .B2(n13425), .ZN(n13424) );
  OAI221_X1 U15605 ( .B1(n13426), .B2(keyinput34), .C1(n13425), .C2(
        P1_ADDR_REG_12__SCAN_IN), .A(n13424), .ZN(n13437) );
  INV_X1 U15606 ( .A(keyinput95), .ZN(n13428) );
  AOI22_X1 U15607 ( .A1(n12451), .A2(keyinput15), .B1(P3_DATAO_REG_15__SCAN_IN), .B2(n13428), .ZN(n13427) );
  OAI221_X1 U15608 ( .B1(n12451), .B2(keyinput15), .C1(n13428), .C2(
        P3_DATAO_REG_15__SCAN_IN), .A(n13427), .ZN(n13436) );
  INV_X1 U15609 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15343) );
  AOI22_X1 U15610 ( .A1(n13430), .A2(keyinput24), .B1(n15343), .B2(keyinput53), 
        .ZN(n13429) );
  OAI221_X1 U15611 ( .B1(n13430), .B2(keyinput24), .C1(n15343), .C2(keyinput53), .A(n13429), .ZN(n13435) );
  INV_X1 U15612 ( .A(keyinput4), .ZN(n13431) );
  XOR2_X1 U15613 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n13431), .Z(n13433) );
  XNOR2_X1 U15614 ( .A(P3_IR_REG_27__SCAN_IN), .B(keyinput104), .ZN(n13432) );
  NAND2_X1 U15615 ( .A1(n13433), .A2(n13432), .ZN(n13434) );
  NOR4_X1 U15616 ( .A1(n13437), .A2(n13436), .A3(n13435), .A4(n13434), .ZN(
        n13466) );
  INV_X1 U15617 ( .A(keyinput80), .ZN(n13439) );
  AOI22_X1 U15618 ( .A1(n13440), .A2(keyinput11), .B1(P3_DATAO_REG_30__SCAN_IN), .B2(n13439), .ZN(n13438) );
  OAI221_X1 U15619 ( .B1(n13440), .B2(keyinput11), .C1(n13439), .C2(
        P3_DATAO_REG_30__SCAN_IN), .A(n13438), .ZN(n13451) );
  INV_X1 U15620 ( .A(keyinput100), .ZN(n13442) );
  AOI22_X1 U15621 ( .A1(n13443), .A2(keyinput49), .B1(P2_ADDR_REG_13__SCAN_IN), 
        .B2(n13442), .ZN(n13441) );
  OAI221_X1 U15622 ( .B1(n13443), .B2(keyinput49), .C1(n13442), .C2(
        P2_ADDR_REG_13__SCAN_IN), .A(n13441), .ZN(n13450) );
  INV_X1 U15623 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n13445) );
  AOI22_X1 U15624 ( .A1(n14165), .A2(keyinput119), .B1(keyinput103), .B2(
        n13445), .ZN(n13444) );
  OAI221_X1 U15625 ( .B1(n14165), .B2(keyinput119), .C1(n13445), .C2(
        keyinput103), .A(n13444), .ZN(n13449) );
  INV_X1 U15626 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15373) );
  INV_X1 U15627 ( .A(keyinput50), .ZN(n13447) );
  AOI22_X1 U15628 ( .A1(n15373), .A2(keyinput117), .B1(
        P3_DATAO_REG_14__SCAN_IN), .B2(n13447), .ZN(n13446) );
  OAI221_X1 U15629 ( .B1(n15373), .B2(keyinput117), .C1(n13447), .C2(
        P3_DATAO_REG_14__SCAN_IN), .A(n13446), .ZN(n13448) );
  NOR4_X1 U15630 ( .A1(n13451), .A2(n13450), .A3(n13449), .A4(n13448), .ZN(
        n13465) );
  INV_X1 U15631 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13453) );
  INV_X1 U15632 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n15009) );
  AOI22_X1 U15633 ( .A1(n13453), .A2(keyinput66), .B1(keyinput101), .B2(n15009), .ZN(n13452) );
  OAI221_X1 U15634 ( .B1(n13453), .B2(keyinput66), .C1(n15009), .C2(
        keyinput101), .A(n13452), .ZN(n13463) );
  AOI22_X1 U15635 ( .A1(n13455), .A2(keyinput51), .B1(n9419), .B2(keyinput111), 
        .ZN(n13454) );
  OAI221_X1 U15636 ( .B1(n13455), .B2(keyinput51), .C1(n9419), .C2(keyinput111), .A(n13454), .ZN(n13462) );
  AOI22_X1 U15637 ( .A1(n14906), .A2(keyinput84), .B1(n13457), .B2(keyinput8), 
        .ZN(n13456) );
  OAI221_X1 U15638 ( .B1(n14906), .B2(keyinput84), .C1(n13457), .C2(keyinput8), 
        .A(n13456), .ZN(n13461) );
  XNOR2_X1 U15639 ( .A(P3_IR_REG_15__SCAN_IN), .B(keyinput20), .ZN(n13459) );
  XNOR2_X1 U15640 ( .A(P3_IR_REG_3__SCAN_IN), .B(keyinput63), .ZN(n13458) );
  NAND2_X1 U15641 ( .A1(n13459), .A2(n13458), .ZN(n13460) );
  NOR4_X1 U15642 ( .A1(n13463), .A2(n13462), .A3(n13461), .A4(n13460), .ZN(
        n13464) );
  AND4_X1 U15643 ( .A1(n13467), .A2(n13466), .A3(n13465), .A4(n13464), .ZN(
        n13468) );
  NAND4_X1 U15644 ( .A1(n13471), .A2(n13470), .A3(n13469), .A4(n13468), .ZN(
        n13553) );
  AOI22_X1 U15645 ( .A1(n13474), .A2(keyinput56), .B1(keyinput121), .B2(n13473), .ZN(n13472) );
  OAI221_X1 U15646 ( .B1(n13474), .B2(keyinput56), .C1(n13473), .C2(
        keyinput121), .A(n13472), .ZN(n13482) );
  INV_X1 U15647 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15219) );
  AOI22_X1 U15648 ( .A1(n15219), .A2(keyinput125), .B1(keyinput19), .B2(n13476), .ZN(n13475) );
  OAI221_X1 U15649 ( .B1(n15219), .B2(keyinput125), .C1(n13476), .C2(
        keyinput19), .A(n13475), .ZN(n13481) );
  AOI22_X1 U15650 ( .A1(n8684), .A2(keyinput92), .B1(keyinput127), .B2(n15221), 
        .ZN(n13477) );
  OAI221_X1 U15651 ( .B1(n8684), .B2(keyinput92), .C1(n15221), .C2(keyinput127), .A(n13477), .ZN(n13480) );
  XNOR2_X1 U15652 ( .A(n13478), .B(keyinput70), .ZN(n13479) );
  OR4_X1 U15653 ( .A1(n13482), .A2(n13481), .A3(n13480), .A4(n13479), .ZN(
        n13497) );
  INV_X1 U15654 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13484) );
  OAI22_X1 U15655 ( .A1(n13485), .A2(keyinput62), .B1(n13484), .B2(keyinput94), 
        .ZN(n13483) );
  AOI221_X1 U15656 ( .B1(n13485), .B2(keyinput62), .C1(keyinput94), .C2(n13484), .A(n13483), .ZN(n13495) );
  INV_X1 U15657 ( .A(keyinput43), .ZN(n13487) );
  OAI22_X1 U15658 ( .A1(n13488), .A2(keyinput31), .B1(n13487), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n13486) );
  AOI221_X1 U15659 ( .B1(n13488), .B2(keyinput31), .C1(P1_REG2_REG_21__SCAN_IN), .C2(n13487), .A(n13486), .ZN(n13494) );
  INV_X1 U15660 ( .A(keyinput96), .ZN(n13490) );
  OAI22_X1 U15661 ( .A1(keyinput78), .A2(n7123), .B1(n13490), .B2(
        P2_ADDR_REG_1__SCAN_IN), .ZN(n13489) );
  AOI221_X1 U15662 ( .B1(n7123), .B2(keyinput78), .C1(n13490), .C2(
        P2_ADDR_REG_1__SCAN_IN), .A(n13489), .ZN(n13493) );
  OAI22_X1 U15663 ( .A1(n15350), .A2(keyinput52), .B1(n10950), .B2(keyinput98), 
        .ZN(n13491) );
  AOI221_X1 U15664 ( .B1(n15350), .B2(keyinput52), .C1(keyinput98), .C2(n10950), .A(n13491), .ZN(n13492) );
  NAND4_X1 U15665 ( .A1(n13495), .A2(n13494), .A3(n13493), .A4(n13492), .ZN(
        n13496) );
  NOR2_X1 U15666 ( .A1(n13497), .A2(n13496), .ZN(n13551) );
  AOI22_X1 U15667 ( .A1(n13590), .A2(keyinput47), .B1(n7774), .B2(keyinput14), 
        .ZN(n13498) );
  OAI221_X1 U15668 ( .B1(n13590), .B2(keyinput47), .C1(n7774), .C2(keyinput14), 
        .A(n13498), .ZN(n13509) );
  INV_X1 U15669 ( .A(keyinput126), .ZN(n13500) );
  AOI22_X1 U15670 ( .A1(n13501), .A2(keyinput46), .B1(P3_ADDR_REG_7__SCAN_IN), 
        .B2(n13500), .ZN(n13499) );
  OAI221_X1 U15671 ( .B1(n13501), .B2(keyinput46), .C1(n13500), .C2(
        P3_ADDR_REG_7__SCAN_IN), .A(n13499), .ZN(n13508) );
  AOI22_X1 U15672 ( .A1(n13503), .A2(keyinput0), .B1(keyinput112), .B2(n7248), 
        .ZN(n13502) );
  OAI221_X1 U15673 ( .B1(n13503), .B2(keyinput0), .C1(n7248), .C2(keyinput112), 
        .A(n13502), .ZN(n13507) );
  AOI22_X1 U15674 ( .A1(n15484), .A2(keyinput22), .B1(keyinput2), .B2(n13505), 
        .ZN(n13504) );
  OAI221_X1 U15675 ( .B1(n15484), .B2(keyinput22), .C1(n13505), .C2(keyinput2), 
        .A(n13504), .ZN(n13506) );
  NOR4_X1 U15676 ( .A1(n13509), .A2(n13508), .A3(n13507), .A4(n13506), .ZN(
        n13550) );
  OAI22_X1 U15677 ( .A1(n13512), .A2(keyinput86), .B1(n13511), .B2(keyinput33), 
        .ZN(n13510) );
  AOI221_X1 U15678 ( .B1(n13512), .B2(keyinput86), .C1(keyinput33), .C2(n13511), .A(n13510), .ZN(n13549) );
  AOI22_X1 U15679 ( .A1(n13514), .A2(keyinput1), .B1(keyinput79), .B2(n14991), 
        .ZN(n13513) );
  OAI221_X1 U15680 ( .B1(n13514), .B2(keyinput1), .C1(n14991), .C2(keyinput79), 
        .A(n13513), .ZN(n13530) );
  XNOR2_X1 U15681 ( .A(SI_24_), .B(keyinput68), .ZN(n13518) );
  XNOR2_X1 U15682 ( .A(P1_REG3_REG_19__SCAN_IN), .B(keyinput5), .ZN(n13517) );
  XNOR2_X1 U15683 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput27), .ZN(n13516) );
  XNOR2_X1 U15684 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput3), .ZN(n13515) );
  NAND4_X1 U15685 ( .A1(n13518), .A2(n13517), .A3(n13516), .A4(n13515), .ZN(
        n13529) );
  XNOR2_X1 U15686 ( .A(P3_IR_REG_7__SCAN_IN), .B(keyinput90), .ZN(n13522) );
  XNOR2_X1 U15687 ( .A(P3_IR_REG_28__SCAN_IN), .B(keyinput91), .ZN(n13521) );
  XNOR2_X1 U15688 ( .A(P1_REG3_REG_17__SCAN_IN), .B(keyinput12), .ZN(n13520)
         );
  XNOR2_X1 U15689 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput13), .ZN(n13519)
         );
  NAND4_X1 U15690 ( .A1(n13522), .A2(n13521), .A3(n13520), .A4(n13519), .ZN(
        n13528) );
  XNOR2_X1 U15691 ( .A(P2_REG1_REG_22__SCAN_IN), .B(keyinput35), .ZN(n13526)
         );
  XNOR2_X1 U15692 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput106), .ZN(n13525)
         );
  XNOR2_X1 U15693 ( .A(P3_IR_REG_22__SCAN_IN), .B(keyinput44), .ZN(n13524) );
  XNOR2_X1 U15694 ( .A(P3_IR_REG_17__SCAN_IN), .B(keyinput29), .ZN(n13523) );
  NAND4_X1 U15695 ( .A1(n13526), .A2(n13525), .A3(n13524), .A4(n13523), .ZN(
        n13527) );
  NOR4_X1 U15696 ( .A1(n13530), .A2(n13529), .A3(n13528), .A4(n13527), .ZN(
        n13547) );
  INV_X1 U15697 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15344) );
  INV_X1 U15698 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15358) );
  OAI22_X1 U15699 ( .A1(n15344), .A2(keyinput82), .B1(n15358), .B2(keyinput54), 
        .ZN(n13531) );
  AOI221_X1 U15700 ( .B1(n15344), .B2(keyinput82), .C1(keyinput54), .C2(n15358), .A(n13531), .ZN(n13546) );
  INV_X1 U15701 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n13534) );
  OAI22_X1 U15702 ( .A1(n13534), .A2(keyinput69), .B1(n13533), .B2(keyinput30), 
        .ZN(n13532) );
  AOI221_X1 U15703 ( .B1(n13534), .B2(keyinput69), .C1(keyinput30), .C2(n13533), .A(n13532), .ZN(n13545) );
  INV_X1 U15704 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15558) );
  AOI22_X1 U15705 ( .A1(n15558), .A2(keyinput41), .B1(n7775), .B2(keyinput23), 
        .ZN(n13535) );
  OAI221_X1 U15706 ( .B1(n15558), .B2(keyinput41), .C1(n7775), .C2(keyinput23), 
        .A(n13535), .ZN(n13543) );
  XNOR2_X1 U15707 ( .A(n15222), .B(keyinput6), .ZN(n13542) );
  INV_X1 U15708 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n13536) );
  XOR2_X1 U15709 ( .A(n13536), .B(keyinput36), .Z(n13540) );
  XNOR2_X1 U15710 ( .A(P3_IR_REG_9__SCAN_IN), .B(keyinput110), .ZN(n13539) );
  XNOR2_X1 U15711 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput88), .ZN(n13538) );
  XNOR2_X1 U15712 ( .A(P3_IR_REG_24__SCAN_IN), .B(keyinput21), .ZN(n13537) );
  NAND4_X1 U15713 ( .A1(n13540), .A2(n13539), .A3(n13538), .A4(n13537), .ZN(
        n13541) );
  NOR3_X1 U15714 ( .A1(n13543), .A2(n13542), .A3(n13541), .ZN(n13544) );
  AND4_X1 U15715 ( .A1(n13547), .A2(n13546), .A3(n13545), .A4(n13544), .ZN(
        n13548) );
  NAND4_X1 U15716 ( .A1(n13551), .A2(n13550), .A3(n13549), .A4(n13548), .ZN(
        n13552) );
  NOR4_X1 U15717 ( .A1(n13555), .A2(n13554), .A3(n13553), .A4(n13552), .ZN(
        n13567) );
  XOR2_X1 U15718 ( .A(n13556), .B(n13558), .Z(n13682) );
  XOR2_X1 U15719 ( .A(n13558), .B(n13557), .Z(n13559) );
  OAI222_X1 U15720 ( .A1(n15492), .A2(n13601), .B1(n15494), .B2(n13560), .C1(
        n13559), .C2(n15497), .ZN(n13679) );
  AOI22_X1 U15721 ( .A1(n15489), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15508), 
        .B2(n13561), .ZN(n13562) );
  OAI21_X1 U15722 ( .B1(n13563), .B2(n13587), .A(n13562), .ZN(n13564) );
  AOI21_X1 U15723 ( .B1(n13679), .B2(n15530), .A(n13564), .ZN(n13565) );
  OAI21_X1 U15724 ( .B1(n13606), .B2(n13682), .A(n13565), .ZN(n13566) );
  XOR2_X1 U15725 ( .A(n13567), .B(n13566), .Z(P3_U3218) );
  NAND2_X1 U15726 ( .A1(n13569), .A2(n13568), .ZN(n13577) );
  NAND2_X1 U15727 ( .A1(n13577), .A2(n13570), .ZN(n15063) );
  NAND2_X1 U15728 ( .A1(n15063), .A2(n13571), .ZN(n13573) );
  NAND2_X1 U15729 ( .A1(n13573), .A2(n13572), .ZN(n13597) );
  NAND2_X1 U15730 ( .A1(n13595), .A2(n13574), .ZN(n13575) );
  NAND2_X1 U15731 ( .A1(n13575), .A2(n8005), .ZN(n13581) );
  NAND2_X1 U15732 ( .A1(n13577), .A2(n13576), .ZN(n13579) );
  NAND2_X1 U15733 ( .A1(n13579), .A2(n13578), .ZN(n13580) );
  NAND3_X1 U15734 ( .A1(n13581), .A2(n15513), .A3(n13580), .ZN(n13584) );
  AOI22_X1 U15735 ( .A1(n15065), .A2(n15515), .B1(n15517), .B2(n13582), .ZN(
        n13583) );
  NAND2_X1 U15736 ( .A1(n13584), .A2(n13583), .ZN(n15075) );
  INV_X1 U15737 ( .A(n15075), .ZN(n13594) );
  OAI21_X1 U15738 ( .B1(n13586), .B2(n8005), .A(n13585), .ZN(n15077) );
  NOR2_X1 U15739 ( .A1(n15074), .A2(n13587), .ZN(n13592) );
  INV_X1 U15740 ( .A(n13588), .ZN(n13589) );
  OAI22_X1 U15741 ( .A1(n15530), .A2(n13590), .B1(n13589), .B2(n15525), .ZN(
        n13591) );
  AOI211_X1 U15742 ( .C1(n15077), .C2(n15071), .A(n13592), .B(n13591), .ZN(
        n13593) );
  OAI21_X1 U15743 ( .B1(n15489), .B2(n13594), .A(n13593), .ZN(P3_U3219) );
  INV_X1 U15744 ( .A(n13595), .ZN(n13596) );
  AOI21_X1 U15745 ( .B1(n13598), .B2(n13597), .A(n13596), .ZN(n13599) );
  OAI222_X1 U15746 ( .A1(n15494), .A2(n13601), .B1(n15492), .B2(n13600), .C1(
        n15497), .C2(n13599), .ZN(n13684) );
  INV_X1 U15747 ( .A(n13684), .ZN(n13613) );
  INV_X1 U15748 ( .A(n13740), .ZN(n13610) );
  INV_X1 U15749 ( .A(n13602), .ZN(n13603) );
  OAI22_X1 U15750 ( .A1(n15530), .A2(n13604), .B1(n13603), .B2(n15525), .ZN(
        n13609) );
  INV_X1 U15751 ( .A(n13685), .ZN(n13607) );
  AND2_X1 U15752 ( .A1(n13605), .A2(n8272), .ZN(n13683) );
  NOR3_X1 U15753 ( .A1(n13607), .A2(n13683), .A3(n13606), .ZN(n13608) );
  AOI211_X1 U15754 ( .C1(n13611), .C2(n13610), .A(n13609), .B(n13608), .ZN(
        n13612) );
  OAI21_X1 U15755 ( .B1(n13613), .B2(n15489), .A(n13612), .ZN(P3_U3220) );
  INV_X1 U15756 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n13617) );
  INV_X1 U15757 ( .A(n13689), .ZN(n13614) );
  NAND2_X1 U15758 ( .A1(n12048), .A2(n13614), .ZN(n13616) );
  INV_X1 U15759 ( .A(n13615), .ZN(n13690) );
  NAND2_X1 U15760 ( .A1(n13690), .A2(n15603), .ZN(n13619) );
  OAI211_X1 U15761 ( .C1(n15603), .C2(n13617), .A(n13616), .B(n13619), .ZN(
        P3_U3490) );
  NAND2_X1 U15762 ( .A1(n15600), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n13618) );
  OAI211_X1 U15763 ( .C1(n13695), .C2(n13689), .A(n13619), .B(n13618), .ZN(
        P3_U3489) );
  INV_X1 U15764 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n13622) );
  MUX2_X1 U15765 ( .A(n13622), .B(n13696), .S(n15603), .Z(n13623) );
  OAI21_X1 U15766 ( .B1(n13699), .B2(n13689), .A(n13623), .ZN(P3_U3487) );
  INV_X1 U15767 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13626) );
  AOI21_X1 U15768 ( .B1(n15579), .B2(n13625), .A(n13624), .ZN(n13700) );
  MUX2_X1 U15769 ( .A(n13626), .B(n13700), .S(n15603), .Z(n13627) );
  OAI21_X1 U15770 ( .B1(n13703), .B2(n13689), .A(n13627), .ZN(P3_U3486) );
  INV_X1 U15771 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13632) );
  NOR3_X1 U15772 ( .A1(n13629), .A2(n13628), .A3(n15532), .ZN(n13631) );
  NOR2_X1 U15773 ( .A1(n13631), .A2(n13630), .ZN(n13704) );
  MUX2_X1 U15774 ( .A(n13632), .B(n13704), .S(n15603), .Z(n13633) );
  OAI21_X1 U15775 ( .B1(n13707), .B2(n13689), .A(n13633), .ZN(P3_U3485) );
  INV_X1 U15776 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13636) );
  AOI21_X1 U15777 ( .B1(n15579), .B2(n13635), .A(n13634), .ZN(n13708) );
  MUX2_X1 U15778 ( .A(n13636), .B(n13708), .S(n15603), .Z(n13637) );
  OAI21_X1 U15779 ( .B1(n13711), .B2(n13689), .A(n13637), .ZN(P3_U3484) );
  NAND2_X1 U15780 ( .A1(n13638), .A2(n15579), .ZN(n13639) );
  OAI21_X1 U15781 ( .B1(n13640), .B2(n15559), .A(n13639), .ZN(n13641) );
  MUX2_X1 U15782 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13712), .S(n15603), .Z(
        P3_U3483) );
  OAI22_X1 U15783 ( .A1(n13645), .A2(n13644), .B1(n13643), .B2(n15559), .ZN(
        n13646) );
  OR2_X1 U15784 ( .A1(n13647), .A2(n13646), .ZN(n13713) );
  MUX2_X1 U15785 ( .A(n13713), .B(P3_REG1_REG_23__SCAN_IN), .S(n15600), .Z(
        P3_U3482) );
  INV_X1 U15786 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13650) );
  AOI21_X1 U15787 ( .B1(n15569), .B2(n13649), .A(n13648), .ZN(n13714) );
  MUX2_X1 U15788 ( .A(n13650), .B(n13714), .S(n15603), .Z(n13651) );
  OAI21_X1 U15789 ( .B1(n13717), .B2(n13689), .A(n13651), .ZN(P3_U3481) );
  INV_X1 U15790 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13654) );
  AOI21_X1 U15791 ( .B1(n13653), .B2(n15569), .A(n13652), .ZN(n13718) );
  MUX2_X1 U15792 ( .A(n13654), .B(n13718), .S(n15603), .Z(n13655) );
  OAI21_X1 U15793 ( .B1(n13721), .B2(n13689), .A(n13655), .ZN(P3_U3480) );
  OR2_X1 U15794 ( .A1(n13656), .A2(n15532), .ZN(n13658) );
  NAND2_X1 U15795 ( .A1(n13658), .A2(n13657), .ZN(n13722) );
  MUX2_X1 U15796 ( .A(n13722), .B(P3_REG1_REG_20__SCAN_IN), .S(n15600), .Z(
        n13659) );
  INV_X1 U15797 ( .A(n13659), .ZN(n13660) );
  OAI21_X1 U15798 ( .B1(n13725), .B2(n13689), .A(n13660), .ZN(P3_U3479) );
  AOI21_X1 U15799 ( .B1(n15569), .B2(n13662), .A(n13661), .ZN(n13726) );
  MUX2_X1 U15800 ( .A(n13663), .B(n13726), .S(n15603), .Z(n13664) );
  OAI21_X1 U15801 ( .B1(n13689), .B2(n13729), .A(n13664), .ZN(P3_U3478) );
  NOR2_X1 U15802 ( .A1(n13665), .A2(n15532), .ZN(n13668) );
  AOI21_X1 U15803 ( .B1(n13668), .B2(n13667), .A(n13666), .ZN(n13730) );
  MUX2_X1 U15804 ( .A(n13669), .B(n13730), .S(n15603), .Z(n13670) );
  OAI21_X1 U15805 ( .B1(n13733), .B2(n13689), .A(n13670), .ZN(P3_U3477) );
  NAND2_X1 U15806 ( .A1(n13671), .A2(n15569), .ZN(n13672) );
  OAI211_X1 U15807 ( .C1(n13674), .C2(n15559), .A(n13673), .B(n13672), .ZN(
        n13734) );
  MUX2_X1 U15808 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n13734), .S(n15603), .Z(
        P3_U3476) );
  AOI21_X1 U15809 ( .B1(n15523), .B2(n13676), .A(n13675), .ZN(n13677) );
  OAI21_X1 U15810 ( .B1(n15532), .B2(n13678), .A(n13677), .ZN(n13735) );
  MUX2_X1 U15811 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n13735), .S(n15603), .Z(
        P3_U3475) );
  AOI21_X1 U15812 ( .B1(n15523), .B2(n13680), .A(n13679), .ZN(n13681) );
  OAI21_X1 U15813 ( .B1(n15532), .B2(n13682), .A(n13681), .ZN(n13736) );
  MUX2_X1 U15814 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n13736), .S(n15603), .Z(
        P3_U3474) );
  NOR2_X1 U15815 ( .A1(n13683), .A2(n15532), .ZN(n13686) );
  AOI21_X1 U15816 ( .B1(n13686), .B2(n13685), .A(n13684), .ZN(n13737) );
  MUX2_X1 U15817 ( .A(n13687), .B(n13737), .S(n15603), .Z(n13688) );
  OAI21_X1 U15818 ( .B1(n13689), .B2(n13740), .A(n13688), .ZN(P3_U3472) );
  INV_X1 U15819 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n13692) );
  NAND2_X1 U15820 ( .A1(n12048), .A2(n8344), .ZN(n13691) );
  NAND2_X1 U15821 ( .A1(n13690), .A2(n15582), .ZN(n13694) );
  OAI211_X1 U15822 ( .C1(n15582), .C2(n13692), .A(n13691), .B(n13694), .ZN(
        P3_U3458) );
  NAND2_X1 U15823 ( .A1(n8348), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n13693) );
  OAI211_X1 U15824 ( .C1(n13695), .C2(n13741), .A(n13694), .B(n13693), .ZN(
        P3_U3457) );
  INV_X1 U15825 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13697) );
  MUX2_X1 U15826 ( .A(n13697), .B(n13696), .S(n15582), .Z(n13698) );
  OAI21_X1 U15827 ( .B1(n13699), .B2(n13741), .A(n13698), .ZN(P3_U3455) );
  INV_X1 U15828 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13701) );
  MUX2_X1 U15829 ( .A(n13701), .B(n13700), .S(n15582), .Z(n13702) );
  OAI21_X1 U15830 ( .B1(n13703), .B2(n13741), .A(n13702), .ZN(P3_U3454) );
  INV_X1 U15831 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13705) );
  MUX2_X1 U15832 ( .A(n13705), .B(n13704), .S(n15582), .Z(n13706) );
  OAI21_X1 U15833 ( .B1(n13707), .B2(n13741), .A(n13706), .ZN(P3_U3453) );
  INV_X1 U15834 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13709) );
  MUX2_X1 U15835 ( .A(n13709), .B(n13708), .S(n15582), .Z(n13710) );
  OAI21_X1 U15836 ( .B1(n13711), .B2(n13741), .A(n13710), .ZN(P3_U3452) );
  MUX2_X1 U15837 ( .A(n13712), .B(P3_REG0_REG_24__SCAN_IN), .S(n8348), .Z(
        P3_U3451) );
  MUX2_X1 U15838 ( .A(n13713), .B(P3_REG0_REG_23__SCAN_IN), .S(n8348), .Z(
        P3_U3450) );
  INV_X1 U15839 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13715) );
  MUX2_X1 U15840 ( .A(n13715), .B(n13714), .S(n15582), .Z(n13716) );
  OAI21_X1 U15841 ( .B1(n13717), .B2(n13741), .A(n13716), .ZN(P3_U3449) );
  INV_X1 U15842 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13719) );
  MUX2_X1 U15843 ( .A(n13719), .B(n13718), .S(n15582), .Z(n13720) );
  OAI21_X1 U15844 ( .B1(n13721), .B2(n13741), .A(n13720), .ZN(P3_U3448) );
  MUX2_X1 U15845 ( .A(n13722), .B(P3_REG0_REG_20__SCAN_IN), .S(n8348), .Z(
        n13723) );
  INV_X1 U15846 ( .A(n13723), .ZN(n13724) );
  OAI21_X1 U15847 ( .B1(n13725), .B2(n13741), .A(n13724), .ZN(P3_U3447) );
  INV_X1 U15848 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13727) );
  MUX2_X1 U15849 ( .A(n13727), .B(n13726), .S(n15582), .Z(n13728) );
  OAI21_X1 U15850 ( .B1(n13741), .B2(n13729), .A(n13728), .ZN(P3_U3446) );
  INV_X1 U15851 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13731) );
  MUX2_X1 U15852 ( .A(n13731), .B(n13730), .S(n15582), .Z(n13732) );
  OAI21_X1 U15853 ( .B1(n13733), .B2(n13741), .A(n13732), .ZN(P3_U3444) );
  MUX2_X1 U15854 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n13734), .S(n15582), .Z(
        P3_U3441) );
  MUX2_X1 U15855 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n13735), .S(n15582), .Z(
        P3_U3438) );
  MUX2_X1 U15856 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n13736), .S(n15582), .Z(
        P3_U3435) );
  INV_X1 U15857 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n13738) );
  MUX2_X1 U15858 ( .A(n13738), .B(n13737), .S(n15582), .Z(n13739) );
  OAI21_X1 U15859 ( .B1(n13741), .B2(n13740), .A(n13739), .ZN(P3_U3429) );
  MUX2_X1 U15860 ( .A(n13743), .B(P3_D_REG_0__SCAN_IN), .S(n13742), .Z(
        P3_U3376) );
  INV_X1 U15861 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13744) );
  NAND3_X1 U15862 ( .A1(n13744), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n13746) );
  OAI22_X1 U15863 ( .A1(n13747), .A2(n13746), .B1(n13745), .B2(n12609), .ZN(
        n13748) );
  AOI21_X1 U15864 ( .B1(n13750), .B2(n13749), .A(n13748), .ZN(n13751) );
  INV_X1 U15865 ( .A(n13751), .ZN(P3_U3264) );
  INV_X1 U15866 ( .A(n13752), .ZN(n13755) );
  OAI222_X1 U15867 ( .A1(n13756), .A2(n13755), .B1(n13754), .B2(P3_U3151), 
        .C1(n13753), .C2(n12609), .ZN(P3_U3266) );
  INV_X1 U15868 ( .A(n13757), .ZN(n13758) );
  XNOR2_X1 U15869 ( .A(n14189), .B(n13792), .ZN(n13789) );
  NAND2_X1 U15870 ( .A1(n13893), .A2(n13997), .ZN(n13762) );
  NOR2_X1 U15871 ( .A1(n13789), .A2(n13762), .ZN(n13799) );
  AOI21_X1 U15872 ( .B1(n13789), .B2(n13762), .A(n13799), .ZN(n13763) );
  OAI211_X1 U15873 ( .C1(n13764), .C2(n13763), .A(n13803), .B(n15104), .ZN(
        n13768) );
  AOI22_X1 U15874 ( .A1(n13892), .A2(n14027), .B1(n14025), .B2(n14028), .ZN(
        n13994) );
  AOI22_X1 U15875 ( .A1(n13999), .A2(n13855), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13765) );
  OAI21_X1 U15876 ( .B1(n13994), .B2(n13853), .A(n13765), .ZN(n13766) );
  AOI21_X1 U15877 ( .B1(n14189), .B2(n15107), .A(n13766), .ZN(n13767) );
  NAND2_X1 U15878 ( .A1(n13768), .A2(n13767), .ZN(P2_U3186) );
  INV_X1 U15879 ( .A(n13769), .ZN(n13776) );
  AOI22_X1 U15880 ( .A1(n13770), .A2(n15104), .B1(n13875), .B2(n13895), .ZN(
        n13775) );
  NOR2_X1 U15881 ( .A1(n15111), .A2(n14073), .ZN(n13773) );
  AOI22_X1 U15882 ( .A1(n14026), .A2(n14027), .B1(n14025), .B2(n13896), .ZN(
        n14070) );
  OAI22_X1 U15883 ( .A1(n14070), .A2(n13853), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13771), .ZN(n13772) );
  AOI211_X1 U15884 ( .C1(n14210), .C2(n15107), .A(n13773), .B(n13772), .ZN(
        n13774) );
  OAI21_X1 U15885 ( .B1(n13776), .B2(n13775), .A(n13774), .ZN(P2_U3188) );
  NAND3_X1 U15886 ( .A1(n13777), .A2(n13875), .A3(n13899), .ZN(n13778) );
  OAI21_X1 U15887 ( .B1(n13779), .B2(n13872), .A(n13778), .ZN(n13784) );
  OAI21_X1 U15888 ( .B1(n13782), .B2(n13781), .A(n13780), .ZN(n13783) );
  NAND2_X1 U15889 ( .A1(n13784), .A2(n13783), .ZN(n13788) );
  AOI22_X1 U15890 ( .A1(n13898), .A2(n14027), .B1(n14025), .B2(n13900), .ZN(
        n14133) );
  OAI21_X1 U15891 ( .B1(n14133), .B2(n13853), .A(n13785), .ZN(n13786) );
  AOI21_X1 U15892 ( .B1(n14128), .B2(n13855), .A(n13786), .ZN(n13787) );
  OAI211_X1 U15893 ( .C1(n8992), .C2(n13888), .A(n13788), .B(n13787), .ZN(
        P2_U3191) );
  INV_X1 U15894 ( .A(n13789), .ZN(n13790) );
  NAND3_X1 U15895 ( .A1(n13790), .A2(n13875), .A3(n13893), .ZN(n13791) );
  NAND2_X1 U15896 ( .A1(n13892), .A2(n13997), .ZN(n13793) );
  XNOR2_X1 U15897 ( .A(n13793), .B(n13792), .ZN(n13794) );
  XNOR2_X1 U15898 ( .A(n14270), .B(n13794), .ZN(n13800) );
  NAND2_X1 U15899 ( .A1(n13795), .A2(n13800), .ZN(n13806) );
  AOI22_X1 U15900 ( .A1(n13893), .A2(n14025), .B1(n13891), .B2(n14027), .ZN(
        n13981) );
  INV_X1 U15901 ( .A(n13983), .ZN(n13796) );
  AOI22_X1 U15902 ( .A1(n13796), .A2(n13855), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13797) );
  OAI21_X1 U15903 ( .B1(n13981), .B2(n13853), .A(n13797), .ZN(n13798) );
  AOI21_X1 U15904 ( .B1(n14270), .B2(n15107), .A(n13798), .ZN(n13805) );
  INV_X1 U15905 ( .A(n13799), .ZN(n13802) );
  INV_X1 U15906 ( .A(n13800), .ZN(n13801) );
  NAND4_X1 U15907 ( .A1(n13803), .A2(n15104), .A3(n13802), .A4(n13801), .ZN(
        n13804) );
  NAND3_X1 U15908 ( .A1(n13806), .A2(n13805), .A3(n13804), .ZN(P2_U3192) );
  OAI211_X1 U15909 ( .C1(n13809), .C2(n13808), .A(n13807), .B(n15104), .ZN(
        n13813) );
  AOI22_X1 U15910 ( .A1(n13896), .A2(n14027), .B1(n14025), .B2(n13898), .ZN(
        n14097) );
  OAI22_X1 U15911 ( .A1(n14097), .A2(n13853), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13810), .ZN(n13811) );
  AOI21_X1 U15912 ( .B1(n14102), .B2(n13855), .A(n13811), .ZN(n13812) );
  OAI211_X1 U15913 ( .C1(n14105), .C2(n13888), .A(n13813), .B(n13812), .ZN(
        P2_U3195) );
  INV_X1 U15914 ( .A(n13814), .ZN(n13828) );
  OR2_X1 U15915 ( .A1(n13815), .A2(n13816), .ZN(n13820) );
  NOR3_X1 U15916 ( .A1(n13818), .A2(n13822), .A3(n13817), .ZN(n13819) );
  AOI21_X1 U15917 ( .B1(n13820), .B2(n15104), .A(n13819), .ZN(n13827) );
  OAI22_X1 U15918 ( .A1(n14035), .A2(n15111), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13821), .ZN(n13825) );
  OAI22_X1 U15919 ( .A1(n13823), .A2(n13883), .B1(n13822), .B2(n13881), .ZN(
        n13824) );
  AOI211_X1 U15920 ( .C1(n14031), .C2(n15107), .A(n13825), .B(n13824), .ZN(
        n13826) );
  OAI21_X1 U15921 ( .B1(n13828), .B2(n13827), .A(n13826), .ZN(P2_U3197) );
  AOI21_X1 U15922 ( .B1(n13831), .B2(n13830), .A(n13829), .ZN(n13838) );
  OAI21_X1 U15923 ( .B1(n15111), .B2(n13833), .A(n13832), .ZN(n13836) );
  OAI22_X1 U15924 ( .A1(n13883), .A2(n13834), .B1(n13881), .B2(n15099), .ZN(
        n13835) );
  AOI211_X1 U15925 ( .C1(n14251), .C2(n15107), .A(n13836), .B(n13835), .ZN(
        n13837) );
  OAI21_X1 U15926 ( .B1(n13838), .B2(n13872), .A(n13837), .ZN(P2_U3198) );
  AOI21_X1 U15927 ( .B1(n13841), .B2(n13840), .A(n13839), .ZN(n13847) );
  AND2_X1 U15928 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n15313) );
  OAI22_X1 U15929 ( .A1(n13883), .A2(n13842), .B1(n13881), .B2(n13882), .ZN(
        n13843) );
  AOI211_X1 U15930 ( .C1(n13855), .C2(n13844), .A(n15313), .B(n13843), .ZN(
        n13846) );
  NAND2_X1 U15931 ( .A1(n14293), .A2(n15107), .ZN(n13845) );
  OAI211_X1 U15932 ( .C1(n13847), .C2(n13872), .A(n13846), .B(n13845), .ZN(
        P2_U3200) );
  INV_X1 U15933 ( .A(n13815), .ZN(n13848) );
  OAI211_X1 U15934 ( .C1(n13850), .C2(n13849), .A(n13848), .B(n15104), .ZN(
        n13857) );
  INV_X1 U15935 ( .A(n13851), .ZN(n14055) );
  AOI22_X1 U15936 ( .A1(n13894), .A2(n14027), .B1(n14025), .B2(n13895), .ZN(
        n14045) );
  OAI22_X1 U15937 ( .A1(n14045), .A2(n13853), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13852), .ZN(n13854) );
  AOI21_X1 U15938 ( .B1(n14055), .B2(n13855), .A(n13854), .ZN(n13856) );
  OAI211_X1 U15939 ( .C1(n8993), .C2(n13888), .A(n13857), .B(n13856), .ZN(
        P2_U3201) );
  NAND2_X1 U15940 ( .A1(n6730), .A2(n13858), .ZN(n13859) );
  XNOR2_X1 U15941 ( .A(n6714), .B(n13859), .ZN(n13864) );
  OAI22_X1 U15942 ( .A1(n15111), .A2(n14117), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13860), .ZN(n13862) );
  OAI22_X1 U15943 ( .A1(n13883), .A2(n14114), .B1(n13881), .B2(n14113), .ZN(
        n13861) );
  AOI211_X1 U15944 ( .C1(n14116), .C2(n15107), .A(n13862), .B(n13861), .ZN(
        n13863) );
  OAI21_X1 U15945 ( .B1(n13864), .B2(n13872), .A(n13863), .ZN(P2_U3205) );
  XNOR2_X1 U15946 ( .A(n13866), .B(n13865), .ZN(n13873) );
  AND2_X1 U15947 ( .A1(n13901), .A2(n14025), .ZN(n13867) );
  AOI21_X1 U15948 ( .B1(n13899), .B2(n14027), .A(n13867), .ZN(n14139) );
  INV_X1 U15949 ( .A(n14139), .ZN(n13868) );
  AOI22_X1 U15950 ( .A1(n15106), .A2(n13868), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13869) );
  OAI21_X1 U15951 ( .B1(n14148), .B2(n15111), .A(n13869), .ZN(n13870) );
  AOI21_X1 U15952 ( .B1(n14237), .B2(n15107), .A(n13870), .ZN(n13871) );
  OAI21_X1 U15953 ( .B1(n13873), .B2(n13872), .A(n13871), .ZN(P2_U3210) );
  NAND2_X1 U15954 ( .A1(n15104), .A2(n13874), .ZN(n13878) );
  NAND2_X1 U15955 ( .A1(n13875), .A2(n13903), .ZN(n13877) );
  MUX2_X1 U15956 ( .A(n13878), .B(n13877), .S(n13876), .Z(n13887) );
  NOR2_X1 U15957 ( .A1(n15111), .A2(n13879), .ZN(n13885) );
  OAI22_X1 U15958 ( .A1(n13883), .A2(n13882), .B1(n13881), .B2(n13880), .ZN(
        n13884) );
  AOI211_X1 U15959 ( .C1(P2_REG3_REG_15__SCAN_IN), .C2(P2_U3088), .A(n13885), 
        .B(n13884), .ZN(n13886) );
  OAI211_X1 U15960 ( .C1(n13889), .C2(n13888), .A(n13887), .B(n13886), .ZN(
        P2_U3213) );
  MUX2_X1 U15961 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13963), .S(n6589), .Z(
        P2_U3562) );
  MUX2_X1 U15962 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13890), .S(n6589), .Z(
        P2_U3561) );
  MUX2_X1 U15963 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13891), .S(n6589), .Z(
        P2_U3560) );
  MUX2_X1 U15964 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13892), .S(n6589), .Z(
        P2_U3559) );
  MUX2_X1 U15965 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13893), .S(n6589), .Z(
        P2_U3558) );
  MUX2_X1 U15966 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n14028), .S(n6589), .Z(
        P2_U3557) );
  MUX2_X1 U15967 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13894), .S(n6589), .Z(
        P2_U3556) );
  MUX2_X1 U15968 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n14026), .S(n6589), .Z(
        P2_U3555) );
  MUX2_X1 U15969 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13895), .S(n6589), .Z(
        P2_U3554) );
  MUX2_X1 U15970 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13896), .S(n6589), .Z(
        P2_U3553) );
  MUX2_X1 U15971 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13897), .S(n6589), .Z(
        P2_U3552) );
  MUX2_X1 U15972 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13898), .S(n6589), .Z(
        P2_U3551) );
  MUX2_X1 U15973 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13899), .S(n6589), .Z(
        P2_U3550) );
  MUX2_X1 U15974 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13900), .S(n6589), .Z(
        P2_U3549) );
  MUX2_X1 U15975 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13901), .S(n6589), .Z(
        P2_U3548) );
  MUX2_X1 U15976 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13902), .S(n6589), .Z(
        P2_U3547) );
  MUX2_X1 U15977 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13903), .S(n6589), .Z(
        P2_U3546) );
  MUX2_X1 U15978 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13904), .S(n6589), .Z(
        P2_U3545) );
  MUX2_X1 U15979 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13905), .S(n6589), .Z(
        P2_U3543) );
  MUX2_X1 U15980 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13906), .S(n6589), .Z(
        P2_U3542) );
  MUX2_X1 U15981 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13907), .S(n6589), .Z(
        P2_U3541) );
  MUX2_X1 U15982 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13908), .S(n6589), .Z(
        P2_U3540) );
  MUX2_X1 U15983 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13909), .S(n6589), .Z(
        P2_U3539) );
  MUX2_X1 U15984 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13910), .S(n6589), .Z(
        P2_U3538) );
  MUX2_X1 U15985 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13911), .S(n6589), .Z(
        P2_U3537) );
  MUX2_X1 U15986 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13912), .S(n6589), .Z(
        P2_U3536) );
  MUX2_X1 U15987 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13913), .S(n6589), .Z(
        P2_U3535) );
  MUX2_X1 U15988 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13914), .S(n6589), .Z(
        P2_U3534) );
  MUX2_X1 U15989 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13915), .S(n6589), .Z(
        P2_U3533) );
  MUX2_X1 U15990 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9901), .S(n6589), .Z(
        P2_U3532) );
  MUX2_X1 U15991 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n9026), .S(n6589), .Z(
        P2_U3531) );
  NOR3_X1 U15992 ( .A1(n13922), .A2(n13916), .A3(n15281), .ZN(n13919) );
  NOR3_X1 U15993 ( .A1(n13926), .A2(n13917), .A3(n15269), .ZN(n13918) );
  OR3_X1 U15994 ( .A1(n13919), .A2(n15300), .A3(n13918), .ZN(n13924) );
  OAI21_X1 U15995 ( .B1(n13922), .B2(n13921), .A(n13920), .ZN(n13923) );
  AOI22_X1 U15996 ( .A1(n13924), .A2(n13925), .B1(n15319), .B2(n13923), .ZN(
        n13933) );
  NAND2_X1 U15997 ( .A1(n15314), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n13931) );
  NOR3_X1 U15998 ( .A1(n13926), .A2(P2_REG1_REG_9__SCAN_IN), .A3(n13925), .ZN(
        n13929) );
  INV_X1 U15999 ( .A(n13927), .ZN(n13928) );
  OAI21_X1 U16000 ( .B1(n13929), .B2(n13928), .A(n15317), .ZN(n13930) );
  NAND4_X1 U16001 ( .A1(n13933), .A2(n13932), .A3(n13931), .A4(n13930), .ZN(
        P2_U3223) );
  OAI21_X1 U16002 ( .B1(n13936), .B2(n13935), .A(n13934), .ZN(n13937) );
  NAND2_X1 U16003 ( .A1(n13937), .A2(n15319), .ZN(n13950) );
  OAI21_X1 U16004 ( .B1(n15311), .B2(n13939), .A(n13938), .ZN(n13940) );
  AOI21_X1 U16005 ( .B1(n15314), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n13940), 
        .ZN(n13949) );
  INV_X1 U16006 ( .A(n13941), .ZN(n13944) );
  MUX2_X1 U16007 ( .A(n15402), .B(P2_REG1_REG_11__SCAN_IN), .S(n13942), .Z(
        n13943) );
  NAND2_X1 U16008 ( .A1(n13944), .A2(n13943), .ZN(n13946) );
  OAI211_X1 U16009 ( .C1(n13947), .C2(n13946), .A(n13945), .B(n15317), .ZN(
        n13948) );
  NAND3_X1 U16010 ( .A1(n13950), .A2(n13949), .A3(n13948), .ZN(P2_U3225) );
  XOR2_X1 U16011 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13951), .Z(n13961) );
  NAND2_X1 U16012 ( .A1(n15300), .A2(n13952), .ZN(n13954) );
  NAND2_X1 U16013 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3088), .ZN(n13953)
         );
  NAND2_X1 U16014 ( .A1(n13954), .A2(n13953), .ZN(n13959) );
  AOI21_X1 U16015 ( .B1(n13956), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13955), 
        .ZN(n13957) );
  NOR2_X1 U16016 ( .A1(n13957), .A2(n15281), .ZN(n13958) );
  AOI211_X1 U16017 ( .C1(n15314), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13959), 
        .B(n13958), .ZN(n13960) );
  OAI21_X1 U16018 ( .B1(n13961), .B2(n15269), .A(n13960), .ZN(P2_U3232) );
  XNOR2_X1 U16019 ( .A(n14264), .B(n13970), .ZN(n13962) );
  NAND2_X1 U16020 ( .A1(n14174), .A2(n6581), .ZN(n13966) );
  AND2_X1 U16021 ( .A1(n13964), .A2(n13963), .ZN(n14173) );
  INV_X1 U16022 ( .A(n14173), .ZN(n14176) );
  NOR2_X1 U16023 ( .A1(n15331), .A2(n14176), .ZN(n13971) );
  AOI21_X1 U16024 ( .B1(n8990), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13971), .ZN(
        n13965) );
  OAI211_X1 U16025 ( .C1(n14264), .C2(n15334), .A(n13966), .B(n13965), .ZN(
        P2_U3234) );
  NAND2_X1 U16026 ( .A1(n14266), .A2(n13967), .ZN(n13968) );
  NAND2_X1 U16027 ( .A1(n13968), .A2(n10037), .ZN(n13969) );
  AOI21_X1 U16028 ( .B1(n8990), .B2(P2_REG2_REG_30__SCAN_IN), .A(n13971), .ZN(
        n13973) );
  NAND2_X1 U16029 ( .A1(n14266), .A2(n15132), .ZN(n13972) );
  OAI211_X1 U16030 ( .C1(n6699), .C2(n14152), .A(n13973), .B(n13972), .ZN(
        P2_U3235) );
  NAND2_X1 U16031 ( .A1(n13976), .A2(n13975), .ZN(n14185) );
  NOR2_X1 U16032 ( .A1(n13978), .A2(n13977), .ZN(n13980) );
  OAI21_X1 U16033 ( .B1(n13983), .B2(n14147), .A(n14184), .ZN(n13984) );
  NAND2_X1 U16034 ( .A1(n13984), .A2(n14163), .ZN(n13992) );
  AOI21_X1 U16035 ( .B1(n14270), .B2(n6629), .A(n13997), .ZN(n13986) );
  NAND2_X1 U16036 ( .A1(n13986), .A2(n13985), .ZN(n14183) );
  INV_X1 U16037 ( .A(n14183), .ZN(n13990) );
  INV_X1 U16038 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13987) );
  OAI22_X1 U16039 ( .A1(n13988), .A2(n15334), .B1(n14163), .B2(n13987), .ZN(
        n13989) );
  AOI21_X1 U16040 ( .B1(n13990), .B2(n6581), .A(n13989), .ZN(n13991) );
  OAI211_X1 U16041 ( .C1(n14137), .C2(n14185), .A(n13992), .B(n13991), .ZN(
        P2_U3237) );
  XNOR2_X1 U16042 ( .A(n14003), .B(n13993), .ZN(n13996) );
  INV_X1 U16043 ( .A(n13994), .ZN(n13995) );
  AOI21_X1 U16044 ( .B1(n13996), .B2(n6580), .A(n13995), .ZN(n14192) );
  AOI21_X1 U16045 ( .B1(n14189), .B2(n14008), .A(n13997), .ZN(n13998) );
  NAND2_X1 U16046 ( .A1(n13998), .A2(n6629), .ZN(n14191) );
  AOI22_X1 U16047 ( .A1(n13999), .A2(n15329), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15331), .ZN(n14001) );
  NAND2_X1 U16048 ( .A1(n14189), .A2(n15132), .ZN(n14000) );
  OAI211_X1 U16049 ( .C1(n14191), .C2(n14152), .A(n14001), .B(n14000), .ZN(
        n14002) );
  INV_X1 U16050 ( .A(n14002), .ZN(n14006) );
  NAND2_X1 U16051 ( .A1(n14004), .A2(n14003), .ZN(n14187) );
  NAND3_X1 U16052 ( .A1(n14188), .A2(n14187), .A3(n15337), .ZN(n14005) );
  OAI211_X1 U16053 ( .C1(n14192), .C2(n15331), .A(n14006), .B(n14005), .ZN(
        P2_U3238) );
  XNOR2_X1 U16054 ( .A(n14007), .B(n14015), .ZN(n14198) );
  INV_X1 U16055 ( .A(n14034), .ZN(n14010) );
  INV_X1 U16056 ( .A(n14008), .ZN(n14009) );
  AOI211_X1 U16057 ( .C1(n14196), .C2(n14010), .A(n13997), .B(n14009), .ZN(
        n14194) );
  AOI22_X1 U16058 ( .A1(n14011), .A2(n15329), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15331), .ZN(n14012) );
  OAI21_X1 U16059 ( .B1(n14013), .B2(n15334), .A(n14012), .ZN(n14014) );
  AOI21_X1 U16060 ( .B1(n14194), .B2(n6581), .A(n14014), .ZN(n14020) );
  XNOR2_X1 U16061 ( .A(n14016), .B(n14015), .ZN(n14018) );
  OAI21_X1 U16062 ( .B1(n14018), .B2(n15125), .A(n14017), .ZN(n14195) );
  NAND2_X1 U16063 ( .A1(n14195), .A2(n14163), .ZN(n14019) );
  OAI211_X1 U16064 ( .C1(n14198), .C2(n14137), .A(n14020), .B(n14019), .ZN(
        P2_U3239) );
  XNOR2_X1 U16065 ( .A(n14021), .B(n14023), .ZN(n14201) );
  INV_X1 U16066 ( .A(n14201), .ZN(n14041) );
  OAI21_X1 U16067 ( .B1(n14024), .B2(n14023), .A(n14022), .ZN(n14029) );
  AOI222_X1 U16068 ( .A1(n6580), .A2(n14029), .B1(n14028), .B2(n14027), .C1(
        n14026), .C2(n14025), .ZN(n14030) );
  INV_X1 U16069 ( .A(n14030), .ZN(n14199) );
  INV_X1 U16070 ( .A(n14031), .ZN(n14276) );
  NAND2_X1 U16071 ( .A1(n14031), .A2(n14053), .ZN(n14032) );
  NAND2_X1 U16072 ( .A1(n14032), .A2(n10037), .ZN(n14033) );
  NOR2_X1 U16073 ( .A1(n14034), .A2(n14033), .ZN(n14200) );
  NAND2_X1 U16074 ( .A1(n14200), .A2(n6581), .ZN(n14038) );
  INV_X1 U16075 ( .A(n14035), .ZN(n14036) );
  AOI22_X1 U16076 ( .A1(n14036), .A2(n15329), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n15331), .ZN(n14037) );
  OAI211_X1 U16077 ( .C1(n14276), .C2(n15334), .A(n14038), .B(n14037), .ZN(
        n14039) );
  AOI21_X1 U16078 ( .B1(n14199), .B2(n14163), .A(n14039), .ZN(n14040) );
  OAI21_X1 U16079 ( .B1(n14041), .B2(n14137), .A(n14040), .ZN(P2_U3240) );
  INV_X1 U16080 ( .A(n14042), .ZN(n14044) );
  OAI21_X1 U16081 ( .B1(n14044), .B2(n14048), .A(n14043), .ZN(n14047) );
  INV_X1 U16082 ( .A(n14045), .ZN(n14046) );
  AOI21_X1 U16083 ( .B1(n14047), .B2(n6580), .A(n14046), .ZN(n14207) );
  NAND2_X1 U16084 ( .A1(n14049), .A2(n14048), .ZN(n14050) );
  NAND2_X1 U16085 ( .A1(n14051), .A2(n14050), .ZN(n14208) );
  INV_X1 U16086 ( .A(n14208), .ZN(n14059) );
  AOI21_X1 U16087 ( .B1(n14205), .B2(n14064), .A(n13997), .ZN(n14054) );
  AND2_X1 U16088 ( .A1(n14054), .A2(n14053), .ZN(n14204) );
  NAND2_X1 U16089 ( .A1(n14204), .A2(n6581), .ZN(n14057) );
  AOI22_X1 U16090 ( .A1(n14055), .A2(n15329), .B1(n8990), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n14056) );
  OAI211_X1 U16091 ( .C1(n8993), .C2(n15334), .A(n14057), .B(n14056), .ZN(
        n14058) );
  AOI21_X1 U16092 ( .B1(n14059), .B2(n15337), .A(n14058), .ZN(n14060) );
  OAI21_X1 U16093 ( .B1(n14207), .B2(n15331), .A(n14060), .ZN(P2_U3241) );
  OAI21_X1 U16094 ( .B1(n14062), .B2(n14068), .A(n14061), .ZN(n14063) );
  INV_X1 U16095 ( .A(n14063), .ZN(n14213) );
  AOI211_X1 U16096 ( .C1(n14210), .C2(n14085), .A(n13997), .B(n14052), .ZN(
        n14209) );
  INV_X1 U16097 ( .A(n14210), .ZN(n14066) );
  INV_X1 U16098 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14065) );
  OAI22_X1 U16099 ( .A1(n14066), .A2(n15334), .B1(n14065), .B2(n14163), .ZN(
        n14067) );
  AOI21_X1 U16100 ( .B1(n14209), .B2(n6581), .A(n14067), .ZN(n14076) );
  XNOR2_X1 U16101 ( .A(n14069), .B(n14068), .ZN(n14072) );
  INV_X1 U16102 ( .A(n14070), .ZN(n14071) );
  AOI21_X1 U16103 ( .B1(n14072), .B2(n6580), .A(n14071), .ZN(n14211) );
  OAI21_X1 U16104 ( .B1(n14073), .B2(n14147), .A(n14211), .ZN(n14074) );
  NAND2_X1 U16105 ( .A1(n14074), .A2(n14163), .ZN(n14075) );
  OAI211_X1 U16106 ( .C1(n14213), .C2(n14137), .A(n14076), .B(n14075), .ZN(
        P2_U3242) );
  NAND2_X1 U16107 ( .A1(n14082), .A2(n14077), .ZN(n14078) );
  NAND2_X1 U16108 ( .A1(n14079), .A2(n14078), .ZN(n14214) );
  OAI211_X1 U16109 ( .C1(n14082), .C2(n14081), .A(n14080), .B(n6580), .ZN(
        n14084) );
  NAND2_X1 U16110 ( .A1(n14084), .A2(n14083), .ZN(n14215) );
  NAND2_X1 U16111 ( .A1(n14215), .A2(n14163), .ZN(n14092) );
  AOI21_X1 U16112 ( .B1(n14087), .B2(n14099), .A(n13997), .ZN(n14086) );
  AND2_X1 U16113 ( .A1(n14086), .A2(n14085), .ZN(n14216) );
  INV_X1 U16114 ( .A(n14087), .ZN(n14282) );
  AOI22_X1 U16115 ( .A1(n8990), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n14088), 
        .B2(n15329), .ZN(n14089) );
  OAI21_X1 U16116 ( .B1(n14282), .B2(n15334), .A(n14089), .ZN(n14090) );
  AOI21_X1 U16117 ( .B1(n6581), .B2(n14216), .A(n14090), .ZN(n14091) );
  OAI211_X1 U16118 ( .C1(n14214), .C2(n14137), .A(n14092), .B(n14091), .ZN(
        P2_U3243) );
  XNOR2_X1 U16119 ( .A(n14093), .B(n14094), .ZN(n14224) );
  XNOR2_X1 U16120 ( .A(n14096), .B(n14095), .ZN(n14098) );
  OAI21_X1 U16121 ( .B1(n14098), .B2(n15125), .A(n14097), .ZN(n14221) );
  INV_X1 U16122 ( .A(n14115), .ZN(n14101) );
  INV_X1 U16123 ( .A(n14099), .ZN(n14100) );
  AOI211_X1 U16124 ( .C1(n14222), .C2(n14101), .A(n13997), .B(n14100), .ZN(
        n14220) );
  NAND2_X1 U16125 ( .A1(n14220), .A2(n6581), .ZN(n14104) );
  AOI22_X1 U16126 ( .A1(n8990), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14102), 
        .B2(n15329), .ZN(n14103) );
  OAI211_X1 U16127 ( .C1(n14105), .C2(n15334), .A(n14104), .B(n14103), .ZN(
        n14106) );
  AOI21_X1 U16128 ( .B1(n14163), .B2(n14221), .A(n14106), .ZN(n14107) );
  OAI21_X1 U16129 ( .B1(n14137), .B2(n14224), .A(n14107), .ZN(P2_U3244) );
  XOR2_X1 U16130 ( .A(n14111), .B(n14108), .Z(n14227) );
  INV_X1 U16131 ( .A(n14227), .ZN(n14123) );
  AOI21_X1 U16132 ( .B1(n14111), .B2(n14110), .A(n6964), .ZN(n14112) );
  OAI222_X1 U16133 ( .A1(n15098), .A2(n14114), .B1(n15096), .B2(n14113), .C1(
        n15125), .C2(n14112), .ZN(n14225) );
  INV_X1 U16134 ( .A(n14116), .ZN(n14288) );
  AOI211_X1 U16135 ( .C1(n14116), .C2(n14126), .A(n13997), .B(n14115), .ZN(
        n14226) );
  NAND2_X1 U16136 ( .A1(n14226), .A2(n6581), .ZN(n14120) );
  INV_X1 U16137 ( .A(n14117), .ZN(n14118) );
  AOI22_X1 U16138 ( .A1(n8990), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n14118), 
        .B2(n15329), .ZN(n14119) );
  OAI211_X1 U16139 ( .C1(n14288), .C2(n15334), .A(n14120), .B(n14119), .ZN(
        n14121) );
  AOI21_X1 U16140 ( .B1(n14225), .B2(n14163), .A(n14121), .ZN(n14122) );
  OAI21_X1 U16141 ( .B1(n14137), .B2(n14123), .A(n14122), .ZN(P2_U3245) );
  XNOR2_X1 U16142 ( .A(n14124), .B(n14131), .ZN(n14235) );
  INV_X1 U16143 ( .A(n14126), .ZN(n14127) );
  AOI211_X1 U16144 ( .C1(n14233), .C2(n14145), .A(n13997), .B(n14127), .ZN(
        n14232) );
  AOI22_X1 U16145 ( .A1(n8990), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14128), 
        .B2(n15329), .ZN(n14129) );
  OAI21_X1 U16146 ( .B1(n8992), .B2(n15334), .A(n14129), .ZN(n14130) );
  AOI21_X1 U16147 ( .B1(n14232), .B2(n6581), .A(n14130), .ZN(n14136) );
  XOR2_X1 U16148 ( .A(n14132), .B(n14131), .Z(n14134) );
  OAI21_X1 U16149 ( .B1(n14134), .B2(n15125), .A(n14133), .ZN(n14231) );
  NAND2_X1 U16150 ( .A1(n14231), .A2(n14163), .ZN(n14135) );
  OAI211_X1 U16151 ( .C1(n14137), .C2(n14235), .A(n14136), .B(n14135), .ZN(
        P2_U3246) );
  XNOR2_X1 U16152 ( .A(n14142), .B(n6713), .ZN(n14138) );
  NAND2_X1 U16153 ( .A1(n14138), .A2(n6580), .ZN(n14140) );
  NAND2_X1 U16154 ( .A1(n14140), .A2(n14139), .ZN(n14241) );
  INV_X1 U16155 ( .A(n14241), .ZN(n14155) );
  OR2_X1 U16156 ( .A1(n14142), .A2(n14141), .ZN(n14143) );
  NAND2_X1 U16157 ( .A1(n14144), .A2(n14143), .ZN(n14236) );
  AOI21_X1 U16158 ( .B1(n14237), .B2(n6631), .A(n13997), .ZN(n14146) );
  NAND2_X1 U16159 ( .A1(n14146), .A2(n14145), .ZN(n14238) );
  INV_X1 U16160 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n14149) );
  OAI22_X1 U16161 ( .A1(n14163), .A2(n14149), .B1(n14148), .B2(n14147), .ZN(
        n14150) );
  AOI21_X1 U16162 ( .B1(n14237), .B2(n15132), .A(n14150), .ZN(n14151) );
  OAI21_X1 U16163 ( .B1(n14238), .B2(n14152), .A(n14151), .ZN(n14153) );
  AOI21_X1 U16164 ( .B1(n15337), .B2(n14236), .A(n14153), .ZN(n14154) );
  OAI21_X1 U16165 ( .B1(n14155), .B2(n15331), .A(n14154), .ZN(P2_U3247) );
  AOI22_X1 U16166 ( .A1(n6581), .A2(n14157), .B1(n14168), .B2(n14156), .ZN(
        n14162) );
  AOI22_X1 U16167 ( .A1(n15132), .A2(n14158), .B1(n15329), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n14161) );
  MUX2_X1 U16168 ( .A(n13398), .B(n14159), .S(n14163), .Z(n14160) );
  NAND3_X1 U16169 ( .A1(n14162), .A2(n14161), .A3(n14160), .ZN(P2_U3263) );
  MUX2_X1 U16170 ( .A(n14165), .B(n14164), .S(n14163), .Z(n14172) );
  AOI22_X1 U16171 ( .A1(n15132), .A2(n14166), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n15329), .ZN(n14171) );
  AOI22_X1 U16172 ( .A1(n6581), .A2(n14169), .B1(n14168), .B2(n14167), .ZN(
        n14170) );
  NAND3_X1 U16173 ( .A1(n14172), .A2(n14171), .A3(n14170), .ZN(P2_U3264) );
  INV_X1 U16174 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n14175) );
  NOR2_X1 U16175 ( .A1(n14174), .A2(n14173), .ZN(n14262) );
  AOI21_X1 U16176 ( .B1(n14258), .B2(n14179), .A(n14178), .ZN(n14180) );
  OAI211_X1 U16177 ( .C1(n14261), .C2(n14182), .A(n14181), .B(n14180), .ZN(
        n14268) );
  MUX2_X1 U16178 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n14268), .S(n15404), .Z(
        P2_U3528) );
  MUX2_X1 U16179 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14269), .S(n15404), .Z(
        n14186) );
  NAND3_X1 U16180 ( .A1(n14188), .A2(n15372), .A3(n14187), .ZN(n14193) );
  NAND2_X1 U16181 ( .A1(n14189), .A2(n14258), .ZN(n14190) );
  NAND4_X1 U16182 ( .A1(n14193), .A2(n14192), .A3(n14191), .A4(n14190), .ZN(
        n14271) );
  MUX2_X1 U16183 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14271), .S(n15404), .Z(
        P2_U3526) );
  AOI211_X1 U16184 ( .C1(n14258), .C2(n14196), .A(n14195), .B(n14194), .ZN(
        n14197) );
  OAI21_X1 U16185 ( .B1(n14261), .B2(n14198), .A(n14197), .ZN(n14272) );
  MUX2_X1 U16186 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14272), .S(n15404), .Z(
        P2_U3525) );
  AOI211_X1 U16187 ( .C1(n15372), .C2(n14201), .A(n14200), .B(n14199), .ZN(
        n14273) );
  MUX2_X1 U16188 ( .A(n14202), .B(n14273), .S(n15404), .Z(n14203) );
  OAI21_X1 U16189 ( .B1(n14276), .B2(n14230), .A(n14203), .ZN(P2_U3524) );
  AOI21_X1 U16190 ( .B1(n14258), .B2(n14205), .A(n14204), .ZN(n14206) );
  OAI211_X1 U16191 ( .C1(n14261), .C2(n14208), .A(n14207), .B(n14206), .ZN(
        n14277) );
  MUX2_X1 U16192 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14277), .S(n15404), .Z(
        P2_U3523) );
  AOI21_X1 U16193 ( .B1(n14258), .B2(n14210), .A(n14209), .ZN(n14212) );
  OAI211_X1 U16194 ( .C1(n14261), .C2(n14213), .A(n14212), .B(n14211), .ZN(
        n14278) );
  MUX2_X1 U16195 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14278), .S(n15404), .Z(
        P2_U3522) );
  NOR2_X1 U16196 ( .A1(n14214), .A2(n14261), .ZN(n14217) );
  NOR3_X1 U16197 ( .A1(n14217), .A2(n14216), .A3(n14215), .ZN(n14280) );
  MUX2_X1 U16198 ( .A(n14280), .B(n14218), .S(n6794), .Z(n14219) );
  OAI21_X1 U16199 ( .B1(n14282), .B2(n14230), .A(n14219), .ZN(P2_U3521) );
  AOI211_X1 U16200 ( .C1(n14258), .C2(n14222), .A(n14221), .B(n14220), .ZN(
        n14223) );
  OAI21_X1 U16201 ( .B1(n14261), .B2(n14224), .A(n14223), .ZN(n14283) );
  MUX2_X1 U16202 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14283), .S(n15404), .Z(
        P2_U3520) );
  AOI211_X1 U16203 ( .C1(n14227), .C2(n15372), .A(n14226), .B(n14225), .ZN(
        n14284) );
  MUX2_X1 U16204 ( .A(n14228), .B(n14284), .S(n15404), .Z(n14229) );
  OAI21_X1 U16205 ( .B1(n14288), .B2(n14230), .A(n14229), .ZN(P2_U3519) );
  AOI211_X1 U16206 ( .C1(n14258), .C2(n14233), .A(n14232), .B(n14231), .ZN(
        n14234) );
  OAI21_X1 U16207 ( .B1(n14261), .B2(n14235), .A(n14234), .ZN(n14289) );
  MUX2_X1 U16208 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14289), .S(n15404), .Z(
        P2_U3518) );
  AND2_X1 U16209 ( .A1(n14236), .A2(n15372), .ZN(n14242) );
  INV_X1 U16210 ( .A(n14237), .ZN(n14239) );
  OAI21_X1 U16211 ( .B1(n14239), .B2(n15386), .A(n14238), .ZN(n14240) );
  MUX2_X1 U16212 ( .A(n14290), .B(P2_REG1_REG_18__SCAN_IN), .S(n6794), .Z(
        P2_U3517) );
  NOR2_X1 U16213 ( .A1(n14243), .A2(n14261), .ZN(n14246) );
  MUX2_X1 U16214 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14291), .S(n15404), .Z(
        n14247) );
  AOI21_X1 U16215 ( .B1(n14248), .B2(n14293), .A(n14247), .ZN(n14249) );
  INV_X1 U16216 ( .A(n14249), .ZN(P2_U3516) );
  AOI21_X1 U16217 ( .B1(n14258), .B2(n14251), .A(n14250), .ZN(n14253) );
  OAI211_X1 U16218 ( .C1(n14261), .C2(n14254), .A(n14253), .B(n14252), .ZN(
        n14296) );
  MUX2_X1 U16219 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14296), .S(n15404), .Z(
        P2_U3515) );
  AOI211_X1 U16220 ( .C1(n14258), .C2(n14257), .A(n14256), .B(n14255), .ZN(
        n14259) );
  OAI21_X1 U16221 ( .B1(n14261), .B2(n14260), .A(n14259), .ZN(n14297) );
  MUX2_X1 U16222 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n14297), .S(n15404), .Z(
        P2_U3514) );
  AOI21_X1 U16223 ( .B1(n14294), .B2(n14266), .A(n14265), .ZN(n14267) );
  INV_X1 U16224 ( .A(n14267), .ZN(P2_U3497) );
  MUX2_X1 U16225 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n14268), .S(n15393), .Z(
        P2_U3496) );
  MUX2_X1 U16226 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14271), .S(n15393), .Z(
        P2_U3494) );
  MUX2_X1 U16227 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14272), .S(n15393), .Z(
        P2_U3493) );
  INV_X1 U16228 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14274) );
  MUX2_X1 U16229 ( .A(n14274), .B(n14273), .S(n15393), .Z(n14275) );
  OAI21_X1 U16230 ( .B1(n14276), .B2(n14287), .A(n14275), .ZN(P2_U3492) );
  MUX2_X1 U16231 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14277), .S(n15393), .Z(
        P2_U3491) );
  MUX2_X1 U16232 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14278), .S(n15393), .Z(
        P2_U3490) );
  INV_X1 U16233 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n14279) );
  MUX2_X1 U16234 ( .A(n14280), .B(n14279), .S(n15391), .Z(n14281) );
  OAI21_X1 U16235 ( .B1(n14282), .B2(n14287), .A(n14281), .ZN(P2_U3489) );
  MUX2_X1 U16236 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14283), .S(n15393), .Z(
        P2_U3488) );
  INV_X1 U16237 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n14285) );
  MUX2_X1 U16238 ( .A(n14285), .B(n14284), .S(n15393), .Z(n14286) );
  OAI21_X1 U16239 ( .B1(n14288), .B2(n14287), .A(n14286), .ZN(P2_U3487) );
  MUX2_X1 U16240 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14289), .S(n15393), .Z(
        P2_U3486) );
  MUX2_X1 U16241 ( .A(n14290), .B(P2_REG0_REG_18__SCAN_IN), .S(n15391), .Z(
        P2_U3484) );
  MUX2_X1 U16242 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14291), .S(n15393), .Z(
        n14292) );
  AOI21_X1 U16243 ( .B1(n14294), .B2(n14293), .A(n14292), .ZN(n14295) );
  INV_X1 U16244 ( .A(n14295), .ZN(P2_U3481) );
  MUX2_X1 U16245 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14296), .S(n15393), .Z(
        P2_U3478) );
  MUX2_X1 U16246 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n14297), .S(n15393), .Z(
        P2_U3475) );
  INV_X1 U16247 ( .A(n14298), .ZN(n15017) );
  INV_X1 U16248 ( .A(n14299), .ZN(n14302) );
  NOR4_X1 U16249 ( .A1(n14302), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3088), 
        .A4(n14300), .ZN(n14303) );
  AOI21_X1 U16250 ( .B1(n14304), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14303), 
        .ZN(n14305) );
  OAI21_X1 U16251 ( .B1(n15017), .B2(n10596), .A(n14305), .ZN(P2_U3296) );
  NAND2_X1 U16252 ( .A1(n14307), .A2(n14306), .ZN(n14309) );
  OAI211_X1 U16253 ( .C1(n14312), .C2(n14310), .A(n14309), .B(n14308), .ZN(
        P2_U3299) );
  INV_X1 U16254 ( .A(n14311), .ZN(n15029) );
  OAI222_X1 U16255 ( .A1(n10596), .A2(n15029), .B1(P2_U3088), .B2(n14314), 
        .C1(n14313), .C2(n14312), .ZN(P2_U3301) );
  MUX2_X1 U16256 ( .A(n14315), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  AOI22_X1 U16257 ( .A1(n14447), .A2(n14633), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14318) );
  NAND2_X1 U16258 ( .A1(n14438), .A2(n14634), .ZN(n14317) );
  OAI211_X1 U16259 ( .C1(n14441), .C2(n14642), .A(n14318), .B(n14317), .ZN(
        n14319) );
  AOI21_X1 U16260 ( .B1(n14878), .B2(n9832), .A(n14319), .ZN(n14320) );
  OAI21_X1 U16261 ( .B1(n14321), .B2(n14456), .A(n14320), .ZN(P1_U3214) );
  XOR2_X1 U16262 ( .A(n14323), .B(n14322), .Z(n14328) );
  AOI22_X1 U16263 ( .A1(n14447), .A2(n14712), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14325) );
  NAND2_X1 U16264 ( .A1(n14438), .A2(n14711), .ZN(n14324) );
  OAI211_X1 U16265 ( .C1(n14441), .C2(n14701), .A(n14325), .B(n14324), .ZN(
        n14326) );
  AOI21_X1 U16266 ( .B1(n14909), .B2(n9832), .A(n14326), .ZN(n14327) );
  OAI21_X1 U16267 ( .B1(n14328), .B2(n14456), .A(n14327), .ZN(P1_U3216) );
  AOI21_X1 U16268 ( .B1(n14330), .B2(n14329), .A(n14456), .ZN(n14331) );
  NAND2_X1 U16269 ( .A1(n14331), .A2(n10094), .ZN(n14336) );
  AOI22_X1 U16270 ( .A1(n14332), .A2(n9832), .B1(n14447), .B2(n14475), .ZN(
        n14335) );
  AOI22_X1 U16271 ( .A1(n14438), .A2(n14473), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14334) );
  INV_X1 U16272 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14508) );
  NAND2_X1 U16273 ( .A1(n14454), .A2(n14508), .ZN(n14333) );
  NAND4_X1 U16274 ( .A1(n14336), .A2(n14335), .A3(n14334), .A4(n14333), .ZN(
        P1_U3218) );
  AOI21_X1 U16275 ( .B1(n14338), .B2(n14337), .A(n14456), .ZN(n14340) );
  NAND2_X1 U16276 ( .A1(n14340), .A2(n14339), .ZN(n14346) );
  OR2_X1 U16277 ( .A1(n14352), .A2(n14826), .ZN(n14342) );
  NAND2_X1 U16278 ( .A1(n14802), .A2(n14791), .ZN(n14341) );
  AND2_X1 U16279 ( .A1(n14342), .A2(n14341), .ZN(n14935) );
  OAI21_X1 U16280 ( .B1(n14935), .B2(n14410), .A(n14343), .ZN(n14344) );
  AOI21_X1 U16281 ( .B1(n14770), .B2(n14454), .A(n14344), .ZN(n14345) );
  OAI211_X1 U16282 ( .C1(n7153), .C2(n14450), .A(n14346), .B(n14345), .ZN(
        P1_U3219) );
  INV_X1 U16283 ( .A(n14347), .ZN(n14348) );
  AOI21_X1 U16284 ( .B1(n14350), .B2(n14349), .A(n14348), .ZN(n14357) );
  INV_X1 U16285 ( .A(n14738), .ZN(n14354) );
  OAI22_X1 U16286 ( .A1(n14352), .A2(n14824), .B1(n14351), .B2(n14826), .ZN(
        n14922) );
  AOI22_X1 U16287 ( .A1(n14922), .A2(n14362), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14353) );
  OAI21_X1 U16288 ( .B1(n14354), .B2(n14441), .A(n14353), .ZN(n14355) );
  AOI21_X1 U16289 ( .B1(n14742), .B2(n9832), .A(n14355), .ZN(n14356) );
  OAI21_X1 U16290 ( .B1(n14357), .B2(n14456), .A(n14356), .ZN(P1_U3223) );
  XOR2_X1 U16291 ( .A(n14359), .B(n14358), .Z(n14366) );
  NAND2_X1 U16292 ( .A1(n14711), .A2(n14791), .ZN(n14361) );
  NAND2_X1 U16293 ( .A1(n14633), .A2(n14850), .ZN(n14360) );
  NAND2_X1 U16294 ( .A1(n14361), .A2(n14360), .ZN(n14670) );
  AOI22_X1 U16295 ( .A1(n14362), .A2(n14670), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14363) );
  OAI21_X1 U16296 ( .B1(n14441), .B2(n14671), .A(n14363), .ZN(n14364) );
  AOI21_X1 U16297 ( .B1(n14987), .B2(n9832), .A(n14364), .ZN(n14365) );
  OAI21_X1 U16298 ( .B1(n14366), .B2(n14456), .A(n14365), .ZN(P1_U3225) );
  OAI21_X1 U16299 ( .B1(n14369), .B2(n14368), .A(n14367), .ZN(n14370) );
  NAND2_X1 U16300 ( .A1(n14370), .A2(n14425), .ZN(n14375) );
  NOR2_X1 U16301 ( .A1(n14441), .A2(n14832), .ZN(n14373) );
  OAI21_X1 U16302 ( .B1(n14449), .B2(n14825), .A(n14371), .ZN(n14372) );
  AOI211_X1 U16303 ( .C1(n14447), .C2(n14462), .A(n14373), .B(n14372), .ZN(
        n14374) );
  OAI211_X1 U16304 ( .C1(n15012), .C2(n14450), .A(n14375), .B(n14374), .ZN(
        P1_U3226) );
  NOR2_X1 U16305 ( .A1(n14376), .A2(n7339), .ZN(n14381) );
  AOI21_X1 U16306 ( .B1(n14379), .B2(n14378), .A(n14377), .ZN(n14380) );
  OAI21_X1 U16307 ( .B1(n14381), .B2(n14380), .A(n14425), .ZN(n14387) );
  NOR2_X1 U16308 ( .A1(n14441), .A2(n14811), .ZN(n14385) );
  OAI21_X1 U16309 ( .B1(n14449), .B2(n14383), .A(n14382), .ZN(n14384) );
  AOI211_X1 U16310 ( .C1(n14447), .C2(n14461), .A(n14385), .B(n14384), .ZN(
        n14386) );
  OAI211_X1 U16311 ( .C1(n14810), .C2(n14450), .A(n14387), .B(n14386), .ZN(
        P1_U3228) );
  XOR2_X1 U16312 ( .A(n14389), .B(n14388), .Z(n14394) );
  AOI22_X1 U16313 ( .A1(n14447), .A2(n14685), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14391) );
  NAND2_X1 U16314 ( .A1(n14438), .A2(n14684), .ZN(n14390) );
  OAI211_X1 U16315 ( .C1(n14441), .C2(n14692), .A(n14391), .B(n14390), .ZN(
        n14392) );
  AOI21_X1 U16316 ( .B1(n14691), .B2(n9832), .A(n14392), .ZN(n14393) );
  OAI21_X1 U16317 ( .B1(n14394), .B2(n14456), .A(n14393), .ZN(P1_U3229) );
  OAI211_X1 U16318 ( .C1(n14397), .C2(n14396), .A(n14395), .B(n14425), .ZN(
        n14404) );
  OR2_X1 U16319 ( .A1(n14398), .A2(n14826), .ZN(n14400) );
  NAND2_X1 U16320 ( .A1(n14792), .A2(n14791), .ZN(n14399) );
  AND2_X1 U16321 ( .A1(n14400), .A2(n14399), .ZN(n14747) );
  OAI22_X1 U16322 ( .A1(n14747), .A2(n14410), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14401), .ZN(n14402) );
  AOI21_X1 U16323 ( .B1(n14755), .B2(n14454), .A(n14402), .ZN(n14403) );
  OAI211_X1 U16324 ( .C1(n14999), .C2(n14450), .A(n14404), .B(n14403), .ZN(
        P1_U3233) );
  OAI21_X1 U16325 ( .B1(n14407), .B2(n14406), .A(n14405), .ZN(n14408) );
  NAND2_X1 U16326 ( .A1(n14408), .A2(n14425), .ZN(n14414) );
  INV_X1 U16327 ( .A(n14726), .ZN(n14412) );
  AOI22_X1 U16328 ( .A1(n14459), .A2(n14791), .B1(n14850), .B2(n14685), .ZN(
        n14915) );
  INV_X1 U16329 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14409) );
  OAI22_X1 U16330 ( .A1(n14915), .A2(n14410), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14409), .ZN(n14411) );
  AOI21_X1 U16331 ( .B1(n14412), .B2(n14454), .A(n14411), .ZN(n14413) );
  OAI211_X1 U16332 ( .C1(n14450), .C2(n14917), .A(n14414), .B(n14413), .ZN(
        P1_U3235) );
  INV_X1 U16333 ( .A(n14786), .ZN(n15006) );
  OAI21_X1 U16334 ( .B1(n14417), .B2(n14416), .A(n14415), .ZN(n14418) );
  NAND2_X1 U16335 ( .A1(n14418), .A2(n14425), .ZN(n14424) );
  NAND2_X1 U16336 ( .A1(n14447), .A2(n14790), .ZN(n14419) );
  OAI211_X1 U16337 ( .C1(n14449), .C2(n14421), .A(n14420), .B(n14419), .ZN(
        n14422) );
  AOI21_X1 U16338 ( .B1(n14778), .B2(n14454), .A(n14422), .ZN(n14423) );
  OAI211_X1 U16339 ( .C1(n15006), .C2(n14450), .A(n14424), .B(n14423), .ZN(
        P1_U3238) );
  OAI211_X1 U16340 ( .C1(n14428), .C2(n14427), .A(n14426), .B(n14425), .ZN(
        n14435) );
  AOI22_X1 U16341 ( .A1(n14429), .A2(n9832), .B1(n14447), .B2(n14472), .ZN(
        n14434) );
  AOI21_X1 U16342 ( .B1(n14438), .B2(n14470), .A(n14430), .ZN(n14433) );
  OR2_X1 U16343 ( .A1(n14441), .A2(n14431), .ZN(n14432) );
  NAND4_X1 U16344 ( .A1(n14435), .A2(n14434), .A3(n14433), .A4(n14432), .ZN(
        P1_U3239) );
  XOR2_X1 U16345 ( .A(n14437), .B(n14436), .Z(n14444) );
  AOI22_X1 U16346 ( .A1(n14447), .A2(n14684), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14440) );
  NAND2_X1 U16347 ( .A1(n14438), .A2(n14656), .ZN(n14439) );
  OAI211_X1 U16348 ( .C1(n14441), .C2(n14661), .A(n14440), .B(n14439), .ZN(
        n14442) );
  AOI21_X1 U16349 ( .B1(n14887), .B2(n9832), .A(n14442), .ZN(n14443) );
  OAI21_X1 U16350 ( .B1(n14444), .B2(n14456), .A(n14443), .ZN(P1_U3240) );
  XNOR2_X1 U16351 ( .A(n14446), .B(n14445), .ZN(n14457) );
  NAND2_X1 U16352 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15214)
         );
  NAND2_X1 U16353 ( .A1(n14447), .A2(n14463), .ZN(n14448) );
  OAI211_X1 U16354 ( .C1(n14449), .C2(n14805), .A(n15214), .B(n14448), .ZN(
        n14452) );
  NOR2_X1 U16355 ( .A1(n7152), .A2(n14450), .ZN(n14451) );
  AOI211_X1 U16356 ( .C1(n14454), .C2(n14453), .A(n14452), .B(n14451), .ZN(
        n14455) );
  OAI21_X1 U16357 ( .B1(n14457), .B2(n14456), .A(n14455), .ZN(P1_U3241) );
  MUX2_X1 U16358 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14587), .S(n14496), .Z(
        P1_U3591) );
  MUX2_X1 U16359 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14604), .S(n14496), .Z(
        P1_U3590) );
  MUX2_X1 U16360 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14458), .S(n14496), .Z(
        P1_U3589) );
  MUX2_X1 U16361 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14634), .S(n14496), .Z(
        P1_U3588) );
  MUX2_X1 U16362 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14656), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16363 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14633), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16364 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14684), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16365 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14711), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16366 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14685), .S(n14496), .Z(
        P1_U3583) );
  MUX2_X1 U16367 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14712), .S(n14496), .Z(
        P1_U3582) );
  MUX2_X1 U16368 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14459), .S(n14496), .Z(
        P1_U3581) );
  MUX2_X1 U16369 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14460), .S(n14496), .Z(
        P1_U3580) );
  MUX2_X1 U16370 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14792), .S(n14496), .Z(
        P1_U3579) );
  MUX2_X1 U16371 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14802), .S(n14496), .Z(
        P1_U3578) );
  MUX2_X1 U16372 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14790), .S(n14496), .Z(
        P1_U3577) );
  MUX2_X1 U16373 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14461), .S(n14496), .Z(
        P1_U3576) );
  MUX2_X1 U16374 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14462), .S(n14496), .Z(
        P1_U3575) );
  MUX2_X1 U16375 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14463), .S(n14496), .Z(
        P1_U3574) );
  MUX2_X1 U16376 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14464), .S(n14496), .Z(
        P1_U3573) );
  MUX2_X1 U16377 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14465), .S(n14496), .Z(
        P1_U3572) );
  MUX2_X1 U16378 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14466), .S(n14496), .Z(
        P1_U3571) );
  MUX2_X1 U16379 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14467), .S(n14496), .Z(
        P1_U3570) );
  MUX2_X1 U16380 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14468), .S(n14496), .Z(
        P1_U3569) );
  MUX2_X1 U16381 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14469), .S(n14496), .Z(
        P1_U3568) );
  MUX2_X1 U16382 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14470), .S(n14496), .Z(
        P1_U3567) );
  MUX2_X1 U16383 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14471), .S(n14496), .Z(
        P1_U3566) );
  MUX2_X1 U16384 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14472), .S(n14496), .Z(
        P1_U3565) );
  MUX2_X1 U16385 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14473), .S(n14496), .Z(
        P1_U3564) );
  MUX2_X1 U16386 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14474), .S(n14496), .Z(
        P1_U3563) );
  MUX2_X1 U16387 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14475), .S(n14496), .Z(
        P1_U3562) );
  MUX2_X1 U16388 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14851), .S(n14496), .Z(
        P1_U3561) );
  MUX2_X1 U16389 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14476), .S(n14496), .Z(
        P1_U3560) );
  OAI211_X1 U16390 ( .C1(n14492), .C2(n14478), .A(n14576), .B(n14477), .ZN(
        n14489) );
  INV_X1 U16391 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14481) );
  MUX2_X1 U16392 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n14479), .S(n14484), .Z(
        n14480) );
  OAI21_X1 U16393 ( .B1(n9754), .B2(n14481), .A(n14480), .ZN(n14482) );
  NAND3_X1 U16394 ( .A1(n14565), .A2(n14483), .A3(n14482), .ZN(n14488) );
  INV_X1 U16395 ( .A(n14484), .ZN(n14485) );
  NAND2_X1 U16396 ( .A1(n14571), .A2(n14485), .ZN(n14487) );
  AOI22_X1 U16397 ( .A1(n15199), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14486) );
  NAND4_X1 U16398 ( .A1(n14489), .A2(n14488), .A3(n14487), .A4(n14486), .ZN(
        P1_U3244) );
  NOR2_X1 U16399 ( .A1(n6584), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14491) );
  NOR2_X1 U16400 ( .A1(n14491), .A2(n14490), .ZN(n15196) );
  MUX2_X1 U16401 ( .A(n14493), .B(n14492), .S(n15197), .Z(n14495) );
  NAND2_X1 U16402 ( .A1(n14495), .A2(n14494), .ZN(n14497) );
  OAI211_X1 U16403 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n15196), .A(n14497), .B(
        n14496), .ZN(n14542) );
  AOI22_X1 U16404 ( .A1(n15199), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14507) );
  OAI211_X1 U16405 ( .C1(n14499), .C2(n14498), .A(n14565), .B(n14513), .ZN(
        n14503) );
  OAI211_X1 U16406 ( .C1(n14501), .C2(n14500), .A(n14576), .B(n14518), .ZN(
        n14502) );
  OAI211_X1 U16407 ( .C1(n15212), .C2(n14504), .A(n14503), .B(n14502), .ZN(
        n14505) );
  INV_X1 U16408 ( .A(n14505), .ZN(n14506) );
  NAND3_X1 U16409 ( .A1(n14542), .A2(n14507), .A3(n14506), .ZN(P1_U3245) );
  OAI22_X1 U16410 ( .A1(n15216), .A2(n14509), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14508), .ZN(n14510) );
  AOI21_X1 U16411 ( .B1(n14515), .B2(n14571), .A(n14510), .ZN(n14522) );
  MUX2_X1 U16412 ( .A(n9824), .B(P1_REG1_REG_3__SCAN_IN), .S(n14515), .Z(
        n14511) );
  NAND3_X1 U16413 ( .A1(n14513), .A2(n14512), .A3(n14511), .ZN(n14514) );
  NAND3_X1 U16414 ( .A1(n14565), .A2(n14530), .A3(n14514), .ZN(n14521) );
  MUX2_X1 U16415 ( .A(n10848), .B(P1_REG2_REG_3__SCAN_IN), .S(n14515), .Z(
        n14516) );
  NAND3_X1 U16416 ( .A1(n14518), .A2(n14517), .A3(n14516), .ZN(n14519) );
  NAND3_X1 U16417 ( .A1(n14576), .A2(n14536), .A3(n14519), .ZN(n14520) );
  NAND3_X1 U16418 ( .A1(n14522), .A2(n14521), .A3(n14520), .ZN(P1_U3246) );
  AOI21_X1 U16419 ( .B1(n15199), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14523), .ZN(
        n14524) );
  OAI21_X1 U16420 ( .B1(n15212), .B2(n14525), .A(n14524), .ZN(n14526) );
  INV_X1 U16421 ( .A(n14526), .ZN(n14541) );
  INV_X1 U16422 ( .A(n14527), .ZN(n14532) );
  NAND3_X1 U16423 ( .A1(n14530), .A2(n14529), .A3(n14528), .ZN(n14531) );
  NAND3_X1 U16424 ( .A1(n14565), .A2(n14532), .A3(n14531), .ZN(n14540) );
  INV_X1 U16425 ( .A(n14533), .ZN(n14538) );
  NAND3_X1 U16426 ( .A1(n14536), .A2(n14535), .A3(n14534), .ZN(n14537) );
  NAND3_X1 U16427 ( .A1(n14576), .A2(n14538), .A3(n14537), .ZN(n14539) );
  NAND4_X1 U16428 ( .A1(n14542), .A2(n14541), .A3(n14540), .A4(n14539), .ZN(
        P1_U3247) );
  NOR2_X1 U16429 ( .A1(n15212), .A2(n14543), .ZN(n14544) );
  AOI211_X1 U16430 ( .C1(n15199), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n14545), .B(
        n14544), .ZN(n14560) );
  OR3_X1 U16431 ( .A1(n14548), .A2(n14547), .A3(n14546), .ZN(n14549) );
  NAND3_X1 U16432 ( .A1(n14565), .A2(n14550), .A3(n14549), .ZN(n14559) );
  INV_X1 U16433 ( .A(n14551), .ZN(n14554) );
  MUX2_X1 U16434 ( .A(n10950), .B(P1_REG2_REG_7__SCAN_IN), .S(n14552), .Z(
        n14553) );
  NAND2_X1 U16435 ( .A1(n14554), .A2(n14553), .ZN(n14556) );
  OAI211_X1 U16436 ( .C1(n14557), .C2(n14556), .A(n14576), .B(n14555), .ZN(
        n14558) );
  NAND3_X1 U16437 ( .A1(n14560), .A2(n14559), .A3(n14558), .ZN(P1_U3250) );
  INV_X1 U16438 ( .A(n14561), .ZN(n14567) );
  NOR3_X1 U16439 ( .A1(n14564), .A2(n14563), .A3(n14562), .ZN(n14566) );
  OAI21_X1 U16440 ( .B1(n14567), .B2(n14566), .A(n14565), .ZN(n14582) );
  INV_X1 U16441 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14569) );
  OAI21_X1 U16442 ( .B1(n15216), .B2(n14569), .A(n14568), .ZN(n14570) );
  AOI21_X1 U16443 ( .B1(n14572), .B2(n14571), .A(n14570), .ZN(n14581) );
  MUX2_X1 U16444 ( .A(n10960), .B(P1_REG2_REG_9__SCAN_IN), .S(n14572), .Z(
        n14575) );
  INV_X1 U16445 ( .A(n14573), .ZN(n14574) );
  NAND2_X1 U16446 ( .A1(n14575), .A2(n14574), .ZN(n14578) );
  OAI211_X1 U16447 ( .C1(n14579), .C2(n14578), .A(n14577), .B(n14576), .ZN(
        n14580) );
  NAND3_X1 U16448 ( .A1(n14582), .A2(n14581), .A3(n14580), .ZN(P1_U3252) );
  NAND2_X1 U16449 ( .A1(n14611), .A2(n14603), .ZN(n14602) );
  XNOR2_X1 U16450 ( .A(n14584), .B(n14583), .ZN(n14863) );
  NOR2_X1 U16451 ( .A1(n14783), .A2(n14828), .ZN(n14859) );
  NAND2_X1 U16452 ( .A1(n14863), .A2(n14859), .ZN(n14590) );
  INV_X1 U16453 ( .A(P1_B_REG_SCAN_IN), .ZN(n14585) );
  NOR2_X1 U16454 ( .A1(n6584), .A2(n14585), .ZN(n14586) );
  NOR2_X1 U16455 ( .A1(n14826), .A2(n14586), .ZN(n14605) );
  AND2_X1 U16456 ( .A1(n14605), .A2(n14587), .ZN(n14866) );
  INV_X1 U16457 ( .A(n14866), .ZN(n14588) );
  NOR2_X1 U16458 ( .A1(n14855), .A2(n14588), .ZN(n14593) );
  AOI21_X1 U16459 ( .B1(n14855), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14593), 
        .ZN(n14589) );
  OAI211_X1 U16460 ( .C1(n14973), .C2(n14831), .A(n14590), .B(n14589), .ZN(
        P1_U3263) );
  XNOR2_X1 U16461 ( .A(n14591), .B(n14602), .ZN(n14592) );
  NOR2_X1 U16462 ( .A1(n14592), .A2(n14828), .ZN(n14867) );
  NAND2_X1 U16463 ( .A1(n14867), .A2(n14835), .ZN(n14595) );
  AOI21_X1 U16464 ( .B1(n14855), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14593), 
        .ZN(n14594) );
  OAI211_X1 U16465 ( .C1(n14977), .C2(n14831), .A(n14595), .B(n14594), .ZN(
        P1_U3264) );
  NAND2_X1 U16466 ( .A1(n14599), .A2(n14598), .ZN(n14601) );
  XOR2_X1 U16467 ( .A(n14601), .B(n14600), .Z(n14875) );
  OAI211_X1 U16468 ( .C1(n14611), .C2(n14603), .A(n14888), .B(n14602), .ZN(
        n14874) );
  NOR2_X1 U16469 ( .A1(n14874), .A2(n14783), .ZN(n14613) );
  NAND2_X1 U16470 ( .A1(n14605), .A2(n14604), .ZN(n14871) );
  OAI22_X1 U16471 ( .A1(n14607), .A2(n14871), .B1(n14606), .B2(n14852), .ZN(
        n14609) );
  NAND2_X1 U16472 ( .A1(n14634), .A2(n14791), .ZN(n14872) );
  NOR2_X1 U16473 ( .A1(n14855), .A2(n14872), .ZN(n14608) );
  AOI211_X1 U16474 ( .C1(n14855), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14609), 
        .B(n14608), .ZN(n14610) );
  OAI21_X1 U16475 ( .B1(n14611), .B2(n14831), .A(n14610), .ZN(n14612) );
  AOI211_X1 U16476 ( .C1(n14875), .C2(n14856), .A(n14613), .B(n14612), .ZN(
        n14614) );
  OAI21_X1 U16477 ( .B1(n14876), .B2(n14838), .A(n14614), .ZN(P1_U3356) );
  INV_X1 U16478 ( .A(n14615), .ZN(n14622) );
  NAND2_X1 U16479 ( .A1(n14855), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n14616) );
  OAI21_X1 U16480 ( .B1(n14852), .B2(n14617), .A(n14616), .ZN(n14618) );
  AOI21_X1 U16481 ( .B1(n14980), .B2(n14858), .A(n14618), .ZN(n14619) );
  OAI21_X1 U16482 ( .B1(n14620), .B2(n14783), .A(n14619), .ZN(n14621) );
  AOI21_X1 U16483 ( .B1(n14622), .B2(n14857), .A(n14621), .ZN(n14623) );
  OAI21_X1 U16484 ( .B1(n14624), .B2(n14855), .A(n14623), .ZN(P1_U3265) );
  OR2_X1 U16485 ( .A1(n14626), .A2(n14625), .ZN(n14627) );
  NAND2_X1 U16486 ( .A1(n14628), .A2(n14627), .ZN(n14877) );
  NAND2_X1 U16487 ( .A1(n14877), .A2(n14629), .ZN(n14640) );
  OAI21_X1 U16488 ( .B1(n14632), .B2(n14631), .A(n14630), .ZN(n14638) );
  NAND2_X1 U16489 ( .A1(n14633), .A2(n14791), .ZN(n14636) );
  NAND2_X1 U16490 ( .A1(n14634), .A2(n14850), .ZN(n14635) );
  NAND2_X1 U16491 ( .A1(n14636), .A2(n14635), .ZN(n14637) );
  AOI21_X1 U16492 ( .B1(n14638), .B2(n14939), .A(n14637), .ZN(n14639) );
  NAND2_X1 U16493 ( .A1(n14640), .A2(n14639), .ZN(n14884) );
  INV_X1 U16494 ( .A(n14884), .ZN(n14648) );
  AOI21_X1 U16495 ( .B1(n14878), .B2(n14651), .A(n14828), .ZN(n14641) );
  NAND2_X1 U16496 ( .A1(n14641), .A2(n6633), .ZN(n14880) );
  INV_X1 U16497 ( .A(n14642), .ZN(n14643) );
  AOI22_X1 U16498 ( .A1(n14855), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14643), 
        .B2(n14842), .ZN(n14645) );
  NAND2_X1 U16499 ( .A1(n14878), .A2(n14858), .ZN(n14644) );
  OAI211_X1 U16500 ( .C1(n14880), .C2(n14783), .A(n14645), .B(n14644), .ZN(
        n14646) );
  AOI21_X1 U16501 ( .B1(n14877), .B2(n14846), .A(n14646), .ZN(n14647) );
  OAI21_X1 U16502 ( .B1(n14648), .B2(n14855), .A(n14647), .ZN(P1_U3266) );
  XNOR2_X1 U16503 ( .A(n14650), .B(n14649), .ZN(n14892) );
  INV_X1 U16504 ( .A(n14651), .ZN(n14652) );
  AOI21_X1 U16505 ( .B1(n14887), .B2(n14668), .A(n14652), .ZN(n14889) );
  INV_X1 U16506 ( .A(n14889), .ZN(n14658) );
  OAI21_X1 U16507 ( .B1(n14655), .B2(n14654), .A(n14653), .ZN(n14657) );
  AOI222_X1 U16508 ( .A1(n14939), .A2(n14657), .B1(n14656), .B2(n14850), .C1(
        n14684), .C2(n14791), .ZN(n14891) );
  OAI21_X1 U16509 ( .B1(n14659), .B2(n14658), .A(n14891), .ZN(n14660) );
  NAND2_X1 U16510 ( .A1(n14660), .A2(n14840), .ZN(n14665) );
  INV_X1 U16511 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n14662) );
  OAI22_X1 U16512 ( .A1(n14840), .A2(n14662), .B1(n14661), .B2(n14852), .ZN(
        n14663) );
  AOI21_X1 U16513 ( .B1(n14887), .B2(n14858), .A(n14663), .ZN(n14664) );
  OAI211_X1 U16514 ( .C1(n14892), .C2(n14838), .A(n14665), .B(n14664), .ZN(
        P1_U3267) );
  OAI21_X1 U16515 ( .B1(n14667), .B2(n14677), .A(n14666), .ZN(n14898) );
  AOI21_X1 U16516 ( .B1(n14987), .B2(n14689), .A(n14828), .ZN(n14669) );
  NAND2_X1 U16517 ( .A1(n14669), .A2(n14668), .ZN(n14894) );
  INV_X1 U16518 ( .A(n14894), .ZN(n14676) );
  INV_X1 U16519 ( .A(n14987), .ZN(n14674) );
  INV_X1 U16520 ( .A(n14670), .ZN(n14893) );
  OAI22_X1 U16521 ( .A1(n14855), .A2(n14893), .B1(n14671), .B2(n14852), .ZN(
        n14672) );
  AOI21_X1 U16522 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n14855), .A(n14672), 
        .ZN(n14673) );
  OAI21_X1 U16523 ( .B1(n14674), .B2(n14831), .A(n14673), .ZN(n14675) );
  AOI21_X1 U16524 ( .B1(n14676), .B2(n14835), .A(n14675), .ZN(n14680) );
  XNOR2_X1 U16525 ( .A(n14678), .B(n14677), .ZN(n14895) );
  NAND2_X1 U16526 ( .A1(n14895), .A2(n14856), .ZN(n14679) );
  OAI211_X1 U16527 ( .C1(n14898), .C2(n14838), .A(n14680), .B(n14679), .ZN(
        P1_U3268) );
  INV_X1 U16528 ( .A(n14681), .ZN(n14682) );
  AOI21_X1 U16529 ( .B1(n7297), .B2(n14683), .A(n14682), .ZN(n14902) );
  AOI22_X1 U16530 ( .A1(n14791), .A2(n14685), .B1(n14684), .B2(n14850), .ZN(
        n14688) );
  OAI211_X1 U16531 ( .C1(n6676), .C2(n7297), .A(n14939), .B(n6802), .ZN(n14687) );
  OAI211_X1 U16532 ( .C1(n14902), .C2(n14789), .A(n14688), .B(n14687), .ZN(
        n14903) );
  NAND2_X1 U16533 ( .A1(n14903), .A2(n14840), .ZN(n14697) );
  INV_X1 U16534 ( .A(n14689), .ZN(n14690) );
  AOI211_X1 U16535 ( .C1(n14691), .C2(n14703), .A(n14828), .B(n14690), .ZN(
        n14904) );
  INV_X1 U16536 ( .A(n14692), .ZN(n14693) );
  AOI22_X1 U16537 ( .A1(n14855), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14693), 
        .B2(n14842), .ZN(n14694) );
  OAI21_X1 U16538 ( .B1(n7157), .B2(n14831), .A(n14694), .ZN(n14695) );
  AOI21_X1 U16539 ( .B1(n14904), .B2(n14835), .A(n14695), .ZN(n14696) );
  OAI211_X1 U16540 ( .C1(n14902), .C2(n14798), .A(n14697), .B(n14696), .ZN(
        P1_U3269) );
  NAND2_X1 U16541 ( .A1(n14698), .A2(n14708), .ZN(n14699) );
  NAND2_X1 U16542 ( .A1(n14700), .A2(n14699), .ZN(n14908) );
  INV_X1 U16543 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n14702) );
  OAI22_X1 U16544 ( .A1(n14840), .A2(n14702), .B1(n14701), .B2(n14852), .ZN(
        n14706) );
  AOI21_X1 U16545 ( .B1(n14909), .B2(n14724), .A(n14828), .ZN(n14704) );
  NAND2_X1 U16546 ( .A1(n14704), .A2(n14703), .ZN(n14911) );
  NOR2_X1 U16547 ( .A1(n14911), .A2(n14783), .ZN(n14705) );
  AOI211_X1 U16548 ( .C1(n14858), .C2(n14909), .A(n14706), .B(n14705), .ZN(
        n14716) );
  OAI21_X1 U16549 ( .B1(n14709), .B2(n14708), .A(n14707), .ZN(n14710) );
  NAND2_X1 U16550 ( .A1(n14710), .A2(n14939), .ZN(n14714) );
  AOI22_X1 U16551 ( .A1(n14712), .A2(n14791), .B1(n14850), .B2(n14711), .ZN(
        n14713) );
  NAND2_X1 U16552 ( .A1(n14714), .A2(n14713), .ZN(n14913) );
  NAND2_X1 U16553 ( .A1(n14913), .A2(n14840), .ZN(n14715) );
  OAI211_X1 U16554 ( .C1(n14908), .C2(n14838), .A(n14716), .B(n14715), .ZN(
        P1_U3270) );
  OAI21_X1 U16555 ( .B1(n14719), .B2(n14718), .A(n14717), .ZN(n14720) );
  INV_X1 U16556 ( .A(n14720), .ZN(n14921) );
  INV_X1 U16557 ( .A(n14856), .ZN(n14776) );
  OAI21_X1 U16558 ( .B1(n14723), .B2(n14722), .A(n14721), .ZN(n14919) );
  OAI211_X1 U16559 ( .C1(n14917), .C2(n14737), .A(n14888), .B(n14724), .ZN(
        n14916) );
  NOR2_X1 U16560 ( .A1(n14840), .A2(n14725), .ZN(n14728) );
  OAI22_X1 U16561 ( .A1(n14915), .A2(n14855), .B1(n14726), .B2(n14852), .ZN(
        n14727) );
  AOI211_X1 U16562 ( .C1(n14729), .C2(n14858), .A(n14728), .B(n14727), .ZN(
        n14730) );
  OAI21_X1 U16563 ( .B1(n14916), .B2(n14783), .A(n14730), .ZN(n14731) );
  AOI21_X1 U16564 ( .B1(n14919), .B2(n14857), .A(n14731), .ZN(n14732) );
  OAI21_X1 U16565 ( .B1(n14921), .B2(n14776), .A(n14732), .ZN(P1_U3271) );
  XNOR2_X1 U16566 ( .A(n14733), .B(n14734), .ZN(n14929) );
  XNOR2_X1 U16567 ( .A(n14735), .B(n14734), .ZN(n14927) );
  NOR2_X1 U16568 ( .A1(n14753), .A2(n14925), .ZN(n14736) );
  OR3_X1 U16569 ( .A1(n14737), .A2(n14736), .A3(n14828), .ZN(n14924) );
  AOI22_X1 U16570 ( .A1(n14922), .A2(n14840), .B1(n14738), .B2(n14842), .ZN(
        n14739) );
  OAI21_X1 U16571 ( .B1(n14740), .B2(n14840), .A(n14739), .ZN(n14741) );
  AOI21_X1 U16572 ( .B1(n14742), .B2(n14858), .A(n14741), .ZN(n14743) );
  OAI21_X1 U16573 ( .B1(n14924), .B2(n14783), .A(n14743), .ZN(n14744) );
  AOI21_X1 U16574 ( .B1(n14927), .B2(n14857), .A(n14744), .ZN(n14745) );
  OAI21_X1 U16575 ( .B1(n14776), .B2(n14929), .A(n14745), .ZN(P1_U3272) );
  OAI211_X1 U16576 ( .C1(n6677), .C2(n14752), .A(n14746), .B(n14939), .ZN(
        n14748) );
  NAND2_X1 U16577 ( .A1(n14748), .A2(n14747), .ZN(n14931) );
  INV_X1 U16578 ( .A(n14931), .ZN(n14760) );
  INV_X1 U16579 ( .A(n14749), .ZN(n14750) );
  AOI21_X1 U16580 ( .B1(n14752), .B2(n14751), .A(n14750), .ZN(n14932) );
  AOI211_X1 U16581 ( .C1(n14754), .C2(n14767), .A(n14828), .B(n14753), .ZN(
        n14930) );
  NAND2_X1 U16582 ( .A1(n14930), .A2(n14835), .ZN(n14757) );
  AOI22_X1 U16583 ( .A1(n14855), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14755), 
        .B2(n14842), .ZN(n14756) );
  OAI211_X1 U16584 ( .C1(n14999), .C2(n14831), .A(n14757), .B(n14756), .ZN(
        n14758) );
  AOI21_X1 U16585 ( .B1(n14857), .B2(n14932), .A(n14758), .ZN(n14759) );
  OAI21_X1 U16586 ( .B1(n14855), .B2(n14760), .A(n14759), .ZN(P1_U3273) );
  XNOR2_X1 U16587 ( .A(n14762), .B(n14763), .ZN(n14940) );
  INV_X1 U16588 ( .A(n14940), .ZN(n14775) );
  XNOR2_X1 U16589 ( .A(n14764), .B(n14763), .ZN(n14938) );
  NAND2_X1 U16590 ( .A1(n14765), .A2(n14781), .ZN(n14766) );
  NAND3_X1 U16591 ( .A1(n14767), .A2(n14888), .A3(n14766), .ZN(n14936) );
  OAI21_X1 U16592 ( .B1(n14936), .B2(n14768), .A(n14935), .ZN(n14769) );
  NAND2_X1 U16593 ( .A1(n14769), .A2(n14840), .ZN(n14772) );
  AOI22_X1 U16594 ( .A1(n14855), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n14770), 
        .B2(n14842), .ZN(n14771) );
  OAI211_X1 U16595 ( .C1(n7153), .C2(n14831), .A(n14772), .B(n14771), .ZN(
        n14773) );
  AOI21_X1 U16596 ( .B1(n14857), .B2(n14938), .A(n14773), .ZN(n14774) );
  OAI21_X1 U16597 ( .B1(n14776), .B2(n14775), .A(n14774), .ZN(P1_U3274) );
  XNOR2_X1 U16598 ( .A(n14788), .B(n14777), .ZN(n14947) );
  INV_X1 U16599 ( .A(n14778), .ZN(n14779) );
  OAI22_X1 U16600 ( .A1(n14840), .A2(n14780), .B1(n14779), .B2(n14852), .ZN(
        n14785) );
  AOI21_X1 U16601 ( .B1(n14786), .B2(n14807), .A(n14828), .ZN(n14782) );
  NAND2_X1 U16602 ( .A1(n14782), .A2(n14781), .ZN(n14945) );
  NOR2_X1 U16603 ( .A1(n14945), .A2(n14783), .ZN(n14784) );
  AOI211_X1 U16604 ( .C1(n14858), .C2(n14786), .A(n14785), .B(n14784), .ZN(
        n14797) );
  XNOR2_X1 U16605 ( .A(n14788), .B(n14787), .ZN(n14795) );
  OR2_X1 U16606 ( .A1(n14947), .A2(n14789), .ZN(n14794) );
  AOI22_X1 U16607 ( .A1(n14792), .A2(n14850), .B1(n14791), .B2(n14790), .ZN(
        n14793) );
  OAI211_X1 U16608 ( .C1(n15228), .C2(n14795), .A(n14794), .B(n14793), .ZN(
        n14949) );
  NAND2_X1 U16609 ( .A1(n14949), .A2(n14840), .ZN(n14796) );
  OAI211_X1 U16610 ( .C1(n14947), .C2(n14798), .A(n14797), .B(n14796), .ZN(
        P1_U3275) );
  XNOR2_X1 U16611 ( .A(n14800), .B(n14799), .ZN(n14957) );
  AOI21_X1 U16612 ( .B1(n14801), .B2(n12394), .A(n15228), .ZN(n14804) );
  AOI22_X1 U16613 ( .A1(n14804), .A2(n14803), .B1(n14850), .B2(n14802), .ZN(
        n14955) );
  INV_X1 U16614 ( .A(n14955), .ZN(n14806) );
  NOR2_X1 U16615 ( .A1(n14805), .A2(n14824), .ZN(n14953) );
  OAI21_X1 U16616 ( .B1(n14806), .B2(n14953), .A(n14840), .ZN(n14815) );
  INV_X1 U16617 ( .A(n14827), .ZN(n14809) );
  INV_X1 U16618 ( .A(n14807), .ZN(n14808) );
  AOI211_X1 U16619 ( .C1(n14954), .C2(n14809), .A(n14828), .B(n14808), .ZN(
        n14952) );
  NOR2_X1 U16620 ( .A1(n14810), .A2(n14831), .ZN(n14813) );
  OAI22_X1 U16621 ( .A1(n14840), .A2(n11525), .B1(n14811), .B2(n14852), .ZN(
        n14812) );
  AOI211_X1 U16622 ( .C1(n14952), .C2(n14835), .A(n14813), .B(n14812), .ZN(
        n14814) );
  OAI211_X1 U16623 ( .C1(n14957), .C2(n14838), .A(n14815), .B(n14814), .ZN(
        P1_U3276) );
  OAI21_X1 U16624 ( .B1(n14817), .B2(n14821), .A(n14816), .ZN(n14960) );
  INV_X1 U16625 ( .A(n14960), .ZN(n14839) );
  INV_X1 U16626 ( .A(n14818), .ZN(n14819) );
  AOI21_X1 U16627 ( .B1(n14821), .B2(n14820), .A(n14819), .ZN(n14822) );
  OAI222_X1 U16628 ( .A1(n14826), .A2(n14825), .B1(n14824), .B2(n14823), .C1(
        n15228), .C2(n14822), .ZN(n14958) );
  NAND2_X1 U16629 ( .A1(n14958), .A2(n14840), .ZN(n14837) );
  AOI211_X1 U16630 ( .C1(n14830), .C2(n14829), .A(n14828), .B(n14827), .ZN(
        n14959) );
  NOR2_X1 U16631 ( .A1(n15012), .A2(n14831), .ZN(n14834) );
  OAI22_X1 U16632 ( .A1(n14840), .A2(n11392), .B1(n14832), .B2(n14852), .ZN(
        n14833) );
  AOI211_X1 U16633 ( .C1(n14959), .C2(n14835), .A(n14834), .B(n14833), .ZN(
        n14836) );
  OAI211_X1 U16634 ( .C1(n14839), .C2(n14838), .A(n14837), .B(n14836), .ZN(
        P1_U3277) );
  MUX2_X1 U16635 ( .A(n9567), .B(n14841), .S(n14840), .Z(n14849) );
  AOI22_X1 U16636 ( .A1(n14859), .A2(n14843), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n14842), .ZN(n14848) );
  AOI22_X1 U16637 ( .A1(n14846), .A2(n14845), .B1(n14858), .B2(n14844), .ZN(
        n14847) );
  NAND3_X1 U16638 ( .A1(n14849), .A2(n14848), .A3(n14847), .ZN(P1_U3292) );
  NAND2_X1 U16639 ( .A1(n14851), .A2(n14850), .ZN(n15225) );
  OAI22_X1 U16640 ( .A1(n14855), .A2(n15225), .B1(n14853), .B2(n14852), .ZN(
        n14854) );
  AOI21_X1 U16641 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n14855), .A(n14854), .ZN(
        n14862) );
  OAI21_X1 U16642 ( .B1(n14857), .B2(n14856), .A(n15226), .ZN(n14861) );
  OAI21_X1 U16643 ( .B1(n14859), .B2(n14858), .A(n15232), .ZN(n14860) );
  NAND3_X1 U16644 ( .A1(n14862), .A2(n14861), .A3(n14860), .ZN(P1_U3293) );
  AOI21_X1 U16645 ( .B1(n14863), .B2(n14888), .A(n14866), .ZN(n14970) );
  MUX2_X1 U16646 ( .A(n14864), .B(n14970), .S(n15267), .Z(n14865) );
  OAI21_X1 U16647 ( .B1(n14973), .B2(n14963), .A(n14865), .ZN(P1_U3559) );
  NOR2_X1 U16648 ( .A1(n14867), .A2(n14866), .ZN(n14974) );
  MUX2_X1 U16649 ( .A(n14868), .B(n14974), .S(n15267), .Z(n14869) );
  OAI21_X1 U16650 ( .B1(n14977), .B2(n14963), .A(n14869), .ZN(P1_U3558) );
  NAND2_X1 U16651 ( .A1(n14870), .A2(n14966), .ZN(n14873) );
  NAND2_X1 U16652 ( .A1(n14877), .A2(n15248), .ZN(n14882) );
  NAND2_X1 U16653 ( .A1(n14878), .A2(n14966), .ZN(n14879) );
  AND2_X1 U16654 ( .A1(n14880), .A2(n14879), .ZN(n14881) );
  NAND2_X1 U16655 ( .A1(n14882), .A2(n14881), .ZN(n14883) );
  NOR2_X1 U16656 ( .A1(n14884), .A2(n14883), .ZN(n14981) );
  MUX2_X1 U16657 ( .A(n14885), .B(n14981), .S(n15267), .Z(n14886) );
  INV_X1 U16658 ( .A(n14886), .ZN(P1_U3555) );
  AOI22_X1 U16659 ( .A1(n14889), .A2(n14888), .B1(n14887), .B2(n14966), .ZN(
        n14890) );
  OAI211_X1 U16660 ( .C1(n15229), .C2(n14892), .A(n14891), .B(n14890), .ZN(
        n14984) );
  MUX2_X1 U16661 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14984), .S(n15267), .Z(
        P1_U3554) );
  AND2_X1 U16662 ( .A1(n14894), .A2(n14893), .ZN(n14897) );
  NAND2_X1 U16663 ( .A1(n14895), .A2(n14939), .ZN(n14896) );
  OAI211_X1 U16664 ( .C1(n14898), .C2(n15229), .A(n14897), .B(n14896), .ZN(
        n14985) );
  MUX2_X1 U16665 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14985), .S(n15264), .Z(
        n14899) );
  AOI21_X1 U16666 ( .B1(n14900), .B2(n14987), .A(n14899), .ZN(n14901) );
  INV_X1 U16667 ( .A(n14901), .ZN(P1_U3553) );
  INV_X1 U16668 ( .A(n14902), .ZN(n14905) );
  AOI211_X1 U16669 ( .C1(n15248), .C2(n14905), .A(n14904), .B(n14903), .ZN(
        n14990) );
  MUX2_X1 U16670 ( .A(n14906), .B(n14990), .S(n15264), .Z(n14907) );
  OAI21_X1 U16671 ( .B1(n7157), .B2(n14963), .A(n14907), .ZN(P1_U3552) );
  NOR2_X1 U16672 ( .A1(n14908), .A2(n15229), .ZN(n14914) );
  NAND2_X1 U16673 ( .A1(n14909), .A2(n14966), .ZN(n14910) );
  NAND2_X1 U16674 ( .A1(n14911), .A2(n14910), .ZN(n14912) );
  MUX2_X1 U16675 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14993), .S(n15264), .Z(
        P1_U3551) );
  INV_X1 U16676 ( .A(n14966), .ZN(n15251) );
  OAI211_X1 U16677 ( .C1(n15251), .C2(n14917), .A(n14916), .B(n14915), .ZN(
        n14918) );
  AOI21_X1 U16678 ( .B1(n14919), .B2(n15256), .A(n14918), .ZN(n14920) );
  OAI21_X1 U16679 ( .B1(n14921), .B2(n15228), .A(n14920), .ZN(n14994) );
  MUX2_X1 U16680 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14994), .S(n15264), .Z(
        P1_U3550) );
  INV_X1 U16681 ( .A(n14922), .ZN(n14923) );
  OAI211_X1 U16682 ( .C1(n14925), .C2(n15251), .A(n14924), .B(n14923), .ZN(
        n14926) );
  AOI21_X1 U16683 ( .B1(n14927), .B2(n15256), .A(n14926), .ZN(n14928) );
  OAI21_X1 U16684 ( .B1(n14929), .B2(n15228), .A(n14928), .ZN(n14995) );
  MUX2_X1 U16685 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14995), .S(n15264), .Z(
        P1_U3549) );
  AOI211_X1 U16686 ( .C1(n14932), .C2(n15256), .A(n14931), .B(n14930), .ZN(
        n14996) );
  MUX2_X1 U16687 ( .A(n14933), .B(n14996), .S(n15264), .Z(n14934) );
  OAI21_X1 U16688 ( .B1(n14999), .B2(n14963), .A(n14934), .ZN(P1_U3548) );
  NAND2_X1 U16689 ( .A1(n14936), .A2(n14935), .ZN(n14937) );
  AOI21_X1 U16690 ( .B1(n14938), .B2(n15256), .A(n14937), .ZN(n14942) );
  NAND2_X1 U16691 ( .A1(n14940), .A2(n14939), .ZN(n14941) );
  AND2_X1 U16692 ( .A1(n14942), .A2(n14941), .ZN(n15000) );
  MUX2_X1 U16693 ( .A(n14943), .B(n15000), .S(n15264), .Z(n14944) );
  OAI21_X1 U16694 ( .B1(n7153), .B2(n14963), .A(n14944), .ZN(P1_U3547) );
  OAI21_X1 U16695 ( .B1(n14947), .B2(n14946), .A(n14945), .ZN(n14948) );
  NOR2_X1 U16696 ( .A1(n14949), .A2(n14948), .ZN(n15003) );
  MUX2_X1 U16697 ( .A(n14950), .B(n15003), .S(n15264), .Z(n14951) );
  OAI21_X1 U16698 ( .B1(n15006), .B2(n14963), .A(n14951), .ZN(P1_U3546) );
  AOI211_X1 U16699 ( .C1(n14954), .C2(n14966), .A(n14953), .B(n14952), .ZN(
        n14956) );
  OAI211_X1 U16700 ( .C1(n15229), .C2(n14957), .A(n14956), .B(n14955), .ZN(
        n15007) );
  MUX2_X1 U16701 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15007), .S(n15264), .Z(
        P1_U3545) );
  INV_X1 U16702 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14961) );
  AOI211_X1 U16703 ( .C1(n15256), .C2(n14960), .A(n14959), .B(n14958), .ZN(
        n15008) );
  MUX2_X1 U16704 ( .A(n14961), .B(n15008), .S(n15267), .Z(n14962) );
  OAI21_X1 U16705 ( .B1(n15012), .B2(n14963), .A(n14962), .ZN(P1_U3544) );
  AOI211_X1 U16706 ( .C1(n14967), .C2(n14966), .A(n14965), .B(n14964), .ZN(
        n14968) );
  OAI21_X1 U16707 ( .B1(n15229), .B2(n14969), .A(n14968), .ZN(n15013) );
  MUX2_X1 U16708 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15013), .S(n15267), .Z(
        P1_U3543) );
  INV_X1 U16709 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14971) );
  MUX2_X1 U16710 ( .A(n14971), .B(n14970), .S(n15259), .Z(n14972) );
  OAI21_X1 U16711 ( .B1(n14973), .B2(n15011), .A(n14972), .ZN(P1_U3527) );
  INV_X1 U16712 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14975) );
  MUX2_X1 U16713 ( .A(n14975), .B(n14974), .S(n15259), .Z(n14976) );
  OAI21_X1 U16714 ( .B1(n14977), .B2(n15011), .A(n14976), .ZN(P1_U3526) );
  MUX2_X1 U16715 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14978), .S(n15259), .Z(
        P1_U3525) );
  MUX2_X1 U16716 ( .A(n14982), .B(n14981), .S(n15259), .Z(n14983) );
  INV_X1 U16717 ( .A(n14983), .ZN(P1_U3523) );
  MUX2_X1 U16718 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14984), .S(n15259), .Z(
        P1_U3522) );
  MUX2_X1 U16719 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14985), .S(n15259), .Z(
        n14986) );
  AOI21_X1 U16720 ( .B1(n14988), .B2(n14987), .A(n14986), .ZN(n14989) );
  INV_X1 U16721 ( .A(n14989), .ZN(P1_U3521) );
  MUX2_X1 U16722 ( .A(n14991), .B(n14990), .S(n15259), .Z(n14992) );
  OAI21_X1 U16723 ( .B1(n7157), .B2(n15011), .A(n14992), .ZN(P1_U3520) );
  MUX2_X1 U16724 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14993), .S(n15259), .Z(
        P1_U3519) );
  MUX2_X1 U16725 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14994), .S(n15259), .Z(
        P1_U3518) );
  MUX2_X1 U16726 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14995), .S(n15259), .Z(
        P1_U3517) );
  INV_X1 U16727 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n14997) );
  MUX2_X1 U16728 ( .A(n14997), .B(n14996), .S(n15259), .Z(n14998) );
  OAI21_X1 U16729 ( .B1(n14999), .B2(n15011), .A(n14998), .ZN(P1_U3516) );
  INV_X1 U16730 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n15001) );
  MUX2_X1 U16731 ( .A(n15001), .B(n15000), .S(n15259), .Z(n15002) );
  OAI21_X1 U16732 ( .B1(n7153), .B2(n15011), .A(n15002), .ZN(P1_U3515) );
  INV_X1 U16733 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n15004) );
  MUX2_X1 U16734 ( .A(n15004), .B(n15003), .S(n15259), .Z(n15005) );
  OAI21_X1 U16735 ( .B1(n15006), .B2(n15011), .A(n15005), .ZN(P1_U3513) );
  MUX2_X1 U16736 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15007), .S(n15259), .Z(
        P1_U3510) );
  MUX2_X1 U16737 ( .A(n15009), .B(n15008), .S(n15259), .Z(n15010) );
  OAI21_X1 U16738 ( .B1(n15012), .B2(n15011), .A(n15010), .ZN(P1_U3507) );
  MUX2_X1 U16739 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15013), .S(n15259), .Z(
        P1_U3504) );
  NOR4_X1 U16740 ( .A1(n7629), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9318), .ZN(n15014) );
  AOI21_X1 U16741 ( .B1(n15015), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15014), 
        .ZN(n15016) );
  OAI21_X1 U16742 ( .B1(n15017), .B2(n15030), .A(n15016), .ZN(P1_U3324) );
  OAI222_X1 U16743 ( .A1(P1_U3086), .A2(n15020), .B1(n15030), .B2(n15019), 
        .C1(n15018), .C2(n15024), .ZN(P1_U3325) );
  OAI222_X1 U16744 ( .A1(P1_U3086), .A2(n15023), .B1(n15030), .B2(n15022), 
        .C1(n15021), .C2(n15024), .ZN(P1_U3326) );
  OAI222_X1 U16745 ( .A1(P1_U3086), .A2(n6584), .B1(n15030), .B2(n15026), .C1(
        n15025), .C2(n15024), .ZN(P1_U3328) );
  OAI222_X1 U16746 ( .A1(n15032), .A2(P1_U3086), .B1(n15030), .B2(n15029), 
        .C1(n15028), .C2(n15024), .ZN(P1_U3329) );
  MUX2_X1 U16747 ( .A(n15034), .B(n15033), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16748 ( .A(n15035), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U16749 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15038) );
  OAI21_X1 U16750 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15038), 
        .ZN(U28) );
  AOI21_X1 U16751 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15039) );
  OAI21_X1 U16752 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15039), 
        .ZN(U29) );
  OAI21_X1 U16753 ( .B1(n15042), .B2(n15041), .A(n15040), .ZN(n15043) );
  XNOR2_X1 U16754 ( .A(n15043), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16755 ( .B1(n15046), .B2(n15045), .A(n15044), .ZN(SUB_1596_U57) );
  OAI21_X1 U16756 ( .B1(n15049), .B2(n15048), .A(n15047), .ZN(n15050) );
  XNOR2_X1 U16757 ( .A(n15050), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  OAI21_X1 U16758 ( .B1(n15053), .B2(n15052), .A(n15051), .ZN(SUB_1596_U54) );
  OAI21_X1 U16759 ( .B1(n15056), .B2(n15055), .A(n15054), .ZN(n15057) );
  XNOR2_X1 U16760 ( .A(n15057), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OAI222_X1 U16761 ( .A1(n15062), .A2(n15061), .B1(n15062), .B2(n15060), .C1(
        n15059), .C2(n15058), .ZN(SUB_1596_U63) );
  XNOR2_X1 U16762 ( .A(n15063), .B(n15068), .ZN(n15066) );
  AOI222_X1 U16763 ( .A1(n15513), .A2(n15066), .B1(n15065), .B2(n15517), .C1(
        n15064), .C2(n15515), .ZN(n15079) );
  AOI22_X1 U16764 ( .A1(n15508), .A2(n15067), .B1(n15489), .B2(
        P3_REG2_REG_12__SCAN_IN), .ZN(n15073) );
  XNOR2_X1 U16765 ( .A(n15069), .B(n15068), .ZN(n15082) );
  NOR2_X1 U16766 ( .A1(n15070), .A2(n15559), .ZN(n15081) );
  AOI22_X1 U16767 ( .A1(n15082), .A2(n15071), .B1(n15485), .B2(n15081), .ZN(
        n15072) );
  OAI211_X1 U16768 ( .C1(n15489), .C2(n15079), .A(n15073), .B(n15072), .ZN(
        P3_U3221) );
  NOR2_X1 U16769 ( .A1(n15074), .A2(n15559), .ZN(n15076) );
  AOI211_X1 U16770 ( .C1(n15569), .C2(n15077), .A(n15076), .B(n15075), .ZN(
        n15091) );
  AOI22_X1 U16771 ( .A1(n15603), .A2(n15091), .B1(n15078), .B2(n15600), .ZN(
        P3_U3473) );
  INV_X1 U16772 ( .A(n15079), .ZN(n15080) );
  AOI211_X1 U16773 ( .C1(n15082), .C2(n15569), .A(n15081), .B(n15080), .ZN(
        n15093) );
  INV_X1 U16774 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n15083) );
  AOI22_X1 U16775 ( .A1(n15603), .A2(n15093), .B1(n15083), .B2(n15600), .ZN(
        P3_U3471) );
  AND2_X1 U16776 ( .A1(n15084), .A2(n15569), .ZN(n15087) );
  AND2_X1 U16777 ( .A1(n15085), .A2(n15523), .ZN(n15086) );
  NOR3_X1 U16778 ( .A1(n15088), .A2(n15087), .A3(n15086), .ZN(n15095) );
  AOI22_X1 U16779 ( .A1(n15603), .A2(n15095), .B1(n15089), .B2(n15600), .ZN(
        P3_U3470) );
  INV_X1 U16780 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n15090) );
  AOI22_X1 U16781 ( .A1(n15582), .A2(n15091), .B1(n15090), .B2(n8348), .ZN(
        P3_U3432) );
  INV_X1 U16782 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n15092) );
  AOI22_X1 U16783 ( .A1(n15582), .A2(n15093), .B1(n15092), .B2(n8348), .ZN(
        P3_U3426) );
  INV_X1 U16784 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n15094) );
  AOI22_X1 U16785 ( .A1(n15582), .A2(n15095), .B1(n15094), .B2(n8348), .ZN(
        P3_U3423) );
  OAI22_X1 U16786 ( .A1(n15099), .A2(n15098), .B1(n15097), .B2(n15096), .ZN(
        n15113) );
  NAND2_X1 U16787 ( .A1(n15101), .A2(n15100), .ZN(n15102) );
  NAND2_X1 U16788 ( .A1(n15103), .A2(n15102), .ZN(n15105) );
  AOI222_X1 U16789 ( .A1(n15107), .A2(n15119), .B1(n15113), .B2(n15106), .C1(
        n15105), .C2(n15104), .ZN(n15109) );
  OAI211_X1 U16790 ( .C1(n15111), .C2(n15110), .A(n15109), .B(n15108), .ZN(
        P2_U3187) );
  XOR2_X1 U16791 ( .A(n15117), .B(n15112), .Z(n15115) );
  AOI21_X1 U16792 ( .B1(n15115), .B2(n6580), .A(n15113), .ZN(n15143) );
  AOI222_X1 U16793 ( .A1(n15119), .A2(n15132), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n15331), .C1(n15329), .C2(n15116), .ZN(n15124) );
  XNOR2_X1 U16794 ( .A(n15118), .B(n15117), .ZN(n15146) );
  OAI211_X1 U16795 ( .C1(n7138), .C2(n7139), .A(n10037), .B(n15121), .ZN(
        n15142) );
  INV_X1 U16796 ( .A(n15142), .ZN(n15122) );
  AOI22_X1 U16797 ( .A1(n15146), .A2(n15337), .B1(n6581), .B2(n15122), .ZN(
        n15123) );
  OAI211_X1 U16798 ( .C1(n15331), .C2(n15143), .A(n15124), .B(n15123), .ZN(
        P2_U3251) );
  AOI21_X1 U16799 ( .B1(n15126), .B2(n15134), .A(n15125), .ZN(n15130) );
  INV_X1 U16800 ( .A(n15127), .ZN(n15128) );
  AOI21_X1 U16801 ( .B1(n15130), .B2(n15129), .A(n15128), .ZN(n15156) );
  AOI222_X1 U16802 ( .A1(n15135), .A2(n15132), .B1(P2_REG2_REG_12__SCAN_IN), 
        .B2(n15331), .C1(n15329), .C2(n15131), .ZN(n15141) );
  XNOR2_X1 U16803 ( .A(n15133), .B(n15134), .ZN(n15159) );
  INV_X1 U16804 ( .A(n15135), .ZN(n15157) );
  INV_X1 U16805 ( .A(n15136), .ZN(n15138) );
  OAI211_X1 U16806 ( .C1(n15157), .C2(n15138), .A(n10037), .B(n15137), .ZN(
        n15155) );
  INV_X1 U16807 ( .A(n15155), .ZN(n15139) );
  AOI22_X1 U16808 ( .A1(n15159), .A2(n15337), .B1(n6581), .B2(n15139), .ZN(
        n15140) );
  OAI211_X1 U16809 ( .C1(n8990), .C2(n15156), .A(n15141), .B(n15140), .ZN(
        P2_U3253) );
  OAI21_X1 U16810 ( .B1(n7138), .B2(n15386), .A(n15142), .ZN(n15145) );
  INV_X1 U16811 ( .A(n15143), .ZN(n15144) );
  AOI211_X1 U16812 ( .C1(n15372), .C2(n15146), .A(n15145), .B(n15144), .ZN(
        n15162) );
  AOI22_X1 U16813 ( .A1(n15404), .A2(n15162), .B1(n15147), .B2(n6794), .ZN(
        P2_U3513) );
  INV_X1 U16814 ( .A(n15148), .ZN(n15150) );
  OAI21_X1 U16815 ( .B1(n15150), .B2(n15386), .A(n15149), .ZN(n15152) );
  AOI211_X1 U16816 ( .C1(n15153), .C2(n15372), .A(n15152), .B(n15151), .ZN(
        n15164) );
  AOI22_X1 U16817 ( .A1(n15404), .A2(n15164), .B1(n15154), .B2(n6794), .ZN(
        P2_U3512) );
  OAI211_X1 U16818 ( .C1(n15157), .C2(n15386), .A(n15156), .B(n15155), .ZN(
        n15158) );
  AOI21_X1 U16819 ( .B1(n15372), .B2(n15159), .A(n15158), .ZN(n15166) );
  AOI22_X1 U16820 ( .A1(n15404), .A2(n15166), .B1(n15160), .B2(n6794), .ZN(
        P2_U3511) );
  INV_X1 U16821 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n15161) );
  AOI22_X1 U16822 ( .A1(n15393), .A2(n15162), .B1(n15161), .B2(n15391), .ZN(
        P2_U3472) );
  AOI22_X1 U16823 ( .A1(n15393), .A2(n15164), .B1(n15163), .B2(n15391), .ZN(
        P2_U3469) );
  AOI22_X1 U16824 ( .A1(n15393), .A2(n15166), .B1(n15165), .B2(n15391), .ZN(
        P2_U3466) );
  OAI21_X1 U16825 ( .B1(n15168), .B2(n15251), .A(n15167), .ZN(n15170) );
  AOI211_X1 U16826 ( .C1(n15256), .C2(n15171), .A(n15170), .B(n15169), .ZN(
        n15172) );
  AOI22_X1 U16827 ( .A1(n15267), .A2(n15172), .B1(n11123), .B2(n15265), .ZN(
        P1_U3539) );
  AOI22_X1 U16828 ( .A1(n15259), .A2(n15172), .B1(n11119), .B2(n15257), .ZN(
        P1_U3492) );
  OAI21_X1 U16829 ( .B1(n15175), .B2(n15174), .A(n15173), .ZN(n15176) );
  XNOR2_X1 U16830 ( .A(n15176), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16831 ( .B1(n15179), .B2(n15178), .A(n15177), .ZN(SUB_1596_U68) );
  OAI21_X1 U16832 ( .B1(n15182), .B2(n15181), .A(n15180), .ZN(n15183) );
  XNOR2_X1 U16833 ( .A(n15183), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U16834 ( .B1(n15186), .B2(n15185), .A(n15184), .ZN(n15187) );
  XNOR2_X1 U16835 ( .A(n15187), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AOI21_X1 U16836 ( .B1(n15190), .B2(n15189), .A(n15188), .ZN(n15191) );
  XOR2_X1 U16837 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15191), .Z(SUB_1596_U65)
         );
  OAI21_X1 U16838 ( .B1(n15194), .B2(n15193), .A(n15192), .ZN(n15195) );
  XNOR2_X1 U16839 ( .A(n15195), .B(P2_ADDR_REG_16__SCAN_IN), .ZN(SUB_1596_U64)
         );
  OAI21_X1 U16840 ( .B1(n15197), .B2(P1_REG1_REG_0__SCAN_IN), .A(n15196), .ZN(
        n15198) );
  XOR2_X1 U16841 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15198), .Z(n15202) );
  AOI22_X1 U16842 ( .A1(n15199), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15200) );
  OAI21_X1 U16843 ( .B1(n15202), .B2(n15201), .A(n15200), .ZN(P1_U3243) );
  AOI21_X1 U16844 ( .B1(n15204), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15203), 
        .ZN(n15209) );
  AOI21_X1 U16845 ( .B1(n15206), .B2(P1_REG1_REG_15__SCAN_IN), .A(n15205), 
        .ZN(n15207) );
  OAI222_X1 U16846 ( .A1(n15212), .A2(n15211), .B1(n15210), .B2(n15209), .C1(
        n15208), .C2(n15207), .ZN(n15213) );
  INV_X1 U16847 ( .A(n15213), .ZN(n15215) );
  OAI211_X1 U16848 ( .C1(n15217), .C2(n15216), .A(n15215), .B(n15214), .ZN(
        P1_U3258) );
  AND2_X1 U16849 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15224), .ZN(P1_U3294) );
  AND2_X1 U16850 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15224), .ZN(P1_U3295) );
  AND2_X1 U16851 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15224), .ZN(P1_U3296) );
  INV_X1 U16852 ( .A(n15224), .ZN(n15223) );
  NOR2_X1 U16853 ( .A1(n15223), .A2(n15218), .ZN(P1_U3297) );
  AND2_X1 U16854 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15224), .ZN(P1_U3298) );
  AND2_X1 U16855 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15224), .ZN(P1_U3299) );
  AND2_X1 U16856 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15224), .ZN(P1_U3300) );
  NOR2_X1 U16857 ( .A1(n15223), .A2(n15219), .ZN(P1_U3301) );
  AND2_X1 U16858 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15224), .ZN(P1_U3302) );
  AND2_X1 U16859 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15224), .ZN(P1_U3303) );
  AND2_X1 U16860 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15224), .ZN(P1_U3304) );
  AND2_X1 U16861 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15224), .ZN(P1_U3305) );
  AND2_X1 U16862 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15224), .ZN(P1_U3306) );
  AND2_X1 U16863 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15224), .ZN(P1_U3307) );
  AND2_X1 U16864 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15224), .ZN(P1_U3308) );
  AND2_X1 U16865 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15224), .ZN(P1_U3309) );
  AND2_X1 U16866 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15224), .ZN(P1_U3310) );
  AND2_X1 U16867 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15224), .ZN(P1_U3311) );
  AND2_X1 U16868 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15224), .ZN(P1_U3312) );
  AND2_X1 U16869 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15224), .ZN(P1_U3313) );
  AND2_X1 U16870 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15224), .ZN(P1_U3314) );
  AND2_X1 U16871 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15224), .ZN(P1_U3315) );
  NOR2_X1 U16872 ( .A1(n15223), .A2(n15220), .ZN(P1_U3316) );
  AND2_X1 U16873 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15224), .ZN(P1_U3317) );
  NOR2_X1 U16874 ( .A1(n15223), .A2(n15221), .ZN(P1_U3318) );
  AND2_X1 U16875 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15224), .ZN(P1_U3319) );
  AND2_X1 U16876 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15224), .ZN(P1_U3320) );
  AND2_X1 U16877 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15224), .ZN(P1_U3321) );
  NOR2_X1 U16878 ( .A1(n15223), .A2(n15222), .ZN(P1_U3322) );
  AND2_X1 U16879 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15224), .ZN(P1_U3323) );
  INV_X1 U16880 ( .A(n15225), .ZN(n15231) );
  INV_X1 U16881 ( .A(n15226), .ZN(n15227) );
  AOI21_X1 U16882 ( .B1(n15229), .B2(n15228), .A(n15227), .ZN(n15230) );
  AOI211_X1 U16883 ( .C1(n15233), .C2(n15232), .A(n15231), .B(n15230), .ZN(
        n15260) );
  INV_X1 U16884 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U16885 ( .A1(n15259), .A2(n15260), .B1(n15234), .B2(n15257), .ZN(
        P1_U3459) );
  OAI21_X1 U16886 ( .B1(n15236), .B2(n15251), .A(n15235), .ZN(n15237) );
  AOI21_X1 U16887 ( .B1(n15238), .B2(n15248), .A(n15237), .ZN(n15239) );
  AND2_X1 U16888 ( .A1(n15240), .A2(n15239), .ZN(n15261) );
  AOI22_X1 U16889 ( .A1(n15259), .A2(n15261), .B1(n15241), .B2(n15257), .ZN(
        P1_U3468) );
  OAI21_X1 U16890 ( .B1(n15243), .B2(n15251), .A(n15242), .ZN(n15246) );
  INV_X1 U16891 ( .A(n15244), .ZN(n15245) );
  AOI211_X1 U16892 ( .C1(n15248), .C2(n15247), .A(n15246), .B(n15245), .ZN(
        n15263) );
  AOI22_X1 U16893 ( .A1(n15259), .A2(n15263), .B1(n10023), .B2(n15257), .ZN(
        P1_U3474) );
  INV_X1 U16894 ( .A(n15249), .ZN(n15252) );
  OAI21_X1 U16895 ( .B1(n15252), .B2(n15251), .A(n15250), .ZN(n15254) );
  AOI211_X1 U16896 ( .C1(n15256), .C2(n15255), .A(n15254), .B(n15253), .ZN(
        n15266) );
  INV_X1 U16897 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n15258) );
  AOI22_X1 U16898 ( .A1(n15259), .A2(n15266), .B1(n15258), .B2(n15257), .ZN(
        P1_U3489) );
  AOI22_X1 U16899 ( .A1(n15267), .A2(n15260), .B1(n9754), .B2(n15265), .ZN(
        P1_U3528) );
  AOI22_X1 U16900 ( .A1(n15264), .A2(n15261), .B1(n9824), .B2(n15265), .ZN(
        P1_U3531) );
  AOI22_X1 U16901 ( .A1(n15264), .A2(n15263), .B1(n15262), .B2(n15265), .ZN(
        P1_U3533) );
  AOI22_X1 U16902 ( .A1(n15267), .A2(n15266), .B1(n10738), .B2(n15265), .ZN(
        P1_U3538) );
  NOR2_X1 U16903 ( .A1(n15314), .A2(n6589), .ZN(P2_U3087) );
  AOI21_X1 U16904 ( .B1(n15317), .B2(P2_REG1_REG_0__SCAN_IN), .A(n15268), .ZN(
        n15273) );
  AOI22_X1 U16905 ( .A1(n15314), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n15272) );
  OAI22_X1 U16906 ( .A1(n15281), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n15269), .ZN(n15270) );
  OAI21_X1 U16907 ( .B1(n15300), .B2(n15270), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n15271) );
  OAI211_X1 U16908 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n15273), .A(n15272), .B(
        n15271), .ZN(P2_U3214) );
  INV_X1 U16909 ( .A(n15274), .ZN(n15275) );
  OAI21_X1 U16910 ( .B1(n15311), .B2(n15276), .A(n15275), .ZN(n15277) );
  AOI21_X1 U16911 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n15314), .A(n15277), .ZN(
        n15288) );
  OAI211_X1 U16912 ( .C1(n15280), .C2(n15279), .A(n15317), .B(n15278), .ZN(
        n15287) );
  AOI211_X1 U16913 ( .C1(n15284), .C2(n15283), .A(n15282), .B(n15281), .ZN(
        n15285) );
  INV_X1 U16914 ( .A(n15285), .ZN(n15286) );
  NAND3_X1 U16915 ( .A1(n15288), .A2(n15287), .A3(n15286), .ZN(P2_U3217) );
  AOI22_X1 U16916 ( .A1(n15314), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n15299) );
  OAI211_X1 U16917 ( .C1(n15291), .C2(n15290), .A(n15289), .B(n15319), .ZN(
        n15298) );
  NAND2_X1 U16918 ( .A1(n15300), .A2(n15292), .ZN(n15297) );
  OAI211_X1 U16919 ( .C1(n15295), .C2(n15294), .A(n15293), .B(n15317), .ZN(
        n15296) );
  NAND4_X1 U16920 ( .A1(n15299), .A2(n15298), .A3(n15297), .A4(n15296), .ZN(
        P2_U3227) );
  AOI22_X1 U16921 ( .A1(n15314), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n15309) );
  NAND2_X1 U16922 ( .A1(n15301), .A2(n15300), .ZN(n15308) );
  OAI211_X1 U16923 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15303), .A(n15319), 
        .B(n15302), .ZN(n15307) );
  OAI211_X1 U16924 ( .C1(n15305), .C2(P2_REG1_REG_15__SCAN_IN), .A(n15317), 
        .B(n15304), .ZN(n15306) );
  NAND4_X1 U16925 ( .A1(n15309), .A2(n15308), .A3(n15307), .A4(n15306), .ZN(
        P2_U3229) );
  NOR2_X1 U16926 ( .A1(n15311), .A2(n15310), .ZN(n15312) );
  AOI211_X1 U16927 ( .C1(P2_ADDR_REG_17__SCAN_IN), .C2(n15314), .A(n15313), 
        .B(n15312), .ZN(n15325) );
  XOR2_X1 U16928 ( .A(n15316), .B(n15315), .Z(n15318) );
  NAND2_X1 U16929 ( .A1(n15318), .A2(n15317), .ZN(n15324) );
  OAI211_X1 U16930 ( .C1(n15322), .C2(n15321), .A(n15320), .B(n15319), .ZN(
        n15323) );
  NAND3_X1 U16931 ( .A1(n15325), .A2(n15324), .A3(n15323), .ZN(P2_U3231) );
  NAND2_X1 U16932 ( .A1(n15328), .A2(n6581), .ZN(n15333) );
  AOI22_X1 U16933 ( .A1(n15331), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n15330), 
        .B2(n15329), .ZN(n15332) );
  OAI211_X1 U16934 ( .C1(n7140), .C2(n15334), .A(n15333), .B(n15332), .ZN(
        n15335) );
  AOI21_X1 U16935 ( .B1(n15337), .B2(n15336), .A(n15335), .ZN(n15338) );
  OAI21_X1 U16936 ( .B1(n8990), .B2(n15339), .A(n15338), .ZN(P2_U3258) );
  AND2_X1 U16937 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15346), .ZN(P2_U3266) );
  AND2_X1 U16938 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15346), .ZN(P2_U3267) );
  AND2_X1 U16939 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15346), .ZN(P2_U3268) );
  NOR2_X1 U16940 ( .A1(n15345), .A2(n15341), .ZN(P2_U3269) );
  AND2_X1 U16941 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15346), .ZN(P2_U3270) );
  AND2_X1 U16942 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15346), .ZN(P2_U3271) );
  AND2_X1 U16943 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15346), .ZN(P2_U3272) );
  AND2_X1 U16944 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15346), .ZN(P2_U3273) );
  AND2_X1 U16945 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15346), .ZN(P2_U3274) );
  AND2_X1 U16946 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15346), .ZN(P2_U3275) );
  AND2_X1 U16947 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15346), .ZN(P2_U3276) );
  AND2_X1 U16948 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15346), .ZN(P2_U3277) );
  NOR2_X1 U16949 ( .A1(n15345), .A2(n15342), .ZN(P2_U3278) );
  AND2_X1 U16950 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15346), .ZN(P2_U3279) );
  NOR2_X1 U16951 ( .A1(n15345), .A2(n15343), .ZN(P2_U3280) );
  AND2_X1 U16952 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15346), .ZN(P2_U3281) );
  AND2_X1 U16953 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15346), .ZN(P2_U3282) );
  AND2_X1 U16954 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15346), .ZN(P2_U3283) );
  AND2_X1 U16955 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15346), .ZN(P2_U3284) );
  AND2_X1 U16956 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15346), .ZN(P2_U3285) );
  AND2_X1 U16957 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15346), .ZN(P2_U3286) );
  AND2_X1 U16958 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15346), .ZN(P2_U3287) );
  NOR2_X1 U16959 ( .A1(n15345), .A2(n15344), .ZN(P2_U3288) );
  AND2_X1 U16960 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15346), .ZN(P2_U3289) );
  AND2_X1 U16961 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15346), .ZN(P2_U3290) );
  AND2_X1 U16962 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15346), .ZN(P2_U3291) );
  AND2_X1 U16963 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15346), .ZN(P2_U3292) );
  AND2_X1 U16964 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15346), .ZN(P2_U3293) );
  AND2_X1 U16965 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15346), .ZN(P2_U3294) );
  AND2_X1 U16966 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15346), .ZN(P2_U3295) );
  AOI22_X1 U16967 ( .A1(n15352), .A2(n15348), .B1(n15347), .B2(n15349), .ZN(
        P2_U3416) );
  AOI22_X1 U16968 ( .A1(n15352), .A2(n15351), .B1(n15350), .B2(n15349), .ZN(
        P2_U3417) );
  INV_X1 U16969 ( .A(n15353), .ZN(n15356) );
  INV_X1 U16970 ( .A(n15354), .ZN(n15355) );
  AOI211_X1 U16971 ( .C1(n15390), .C2(n15357), .A(n15356), .B(n15355), .ZN(
        n15395) );
  AOI22_X1 U16972 ( .A1(n15393), .A2(n15395), .B1(n15358), .B2(n15391), .ZN(
        P2_U3430) );
  OAI21_X1 U16973 ( .B1(n15360), .B2(n15386), .A(n15359), .ZN(n15363) );
  INV_X1 U16974 ( .A(n15361), .ZN(n15362) );
  AOI211_X1 U16975 ( .C1(n15372), .C2(n15364), .A(n15363), .B(n15362), .ZN(
        n15396) );
  INV_X1 U16976 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15365) );
  AOI22_X1 U16977 ( .A1(n15393), .A2(n15396), .B1(n15365), .B2(n15391), .ZN(
        P2_U3439) );
  OAI21_X1 U16978 ( .B1(n15367), .B2(n15386), .A(n15366), .ZN(n15370) );
  INV_X1 U16979 ( .A(n15368), .ZN(n15369) );
  AOI211_X1 U16980 ( .C1(n15372), .C2(n15371), .A(n15370), .B(n15369), .ZN(
        n15397) );
  AOI22_X1 U16981 ( .A1(n15393), .A2(n15397), .B1(n15373), .B2(n15391), .ZN(
        P2_U3442) );
  OAI21_X1 U16982 ( .B1(n7500), .B2(n15386), .A(n15374), .ZN(n15376) );
  AOI211_X1 U16983 ( .C1(n15390), .C2(n15377), .A(n15376), .B(n15375), .ZN(
        n15399) );
  INV_X1 U16984 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15378) );
  AOI22_X1 U16985 ( .A1(n15393), .A2(n15399), .B1(n15378), .B2(n15391), .ZN(
        P2_U3454) );
  OAI21_X1 U16986 ( .B1(n15380), .B2(n15386), .A(n15379), .ZN(n15382) );
  AOI211_X1 U16987 ( .C1(n15390), .C2(n15383), .A(n15382), .B(n15381), .ZN(
        n15401) );
  INV_X1 U16988 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15384) );
  AOI22_X1 U16989 ( .A1(n15393), .A2(n15401), .B1(n15384), .B2(n15391), .ZN(
        P2_U3460) );
  OAI21_X1 U16990 ( .B1(n8991), .B2(n15386), .A(n15385), .ZN(n15388) );
  AOI211_X1 U16991 ( .C1(n15390), .C2(n15389), .A(n15388), .B(n15387), .ZN(
        n15403) );
  INV_X1 U16992 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15392) );
  AOI22_X1 U16993 ( .A1(n15393), .A2(n15403), .B1(n15392), .B2(n15391), .ZN(
        P2_U3463) );
  AOI22_X1 U16994 ( .A1(n15404), .A2(n15395), .B1(n15394), .B2(n6794), .ZN(
        P2_U3499) );
  AOI22_X1 U16995 ( .A1(n15404), .A2(n15396), .B1(n9483), .B2(n6794), .ZN(
        P2_U3502) );
  AOI22_X1 U16996 ( .A1(n15404), .A2(n15397), .B1(n9486), .B2(n6794), .ZN(
        P2_U3503) );
  AOI22_X1 U16997 ( .A1(n15404), .A2(n15399), .B1(n15398), .B2(n6794), .ZN(
        P2_U3507) );
  AOI22_X1 U16998 ( .A1(n15404), .A2(n15401), .B1(n15400), .B2(n6794), .ZN(
        P2_U3509) );
  AOI22_X1 U16999 ( .A1(n15404), .A2(n15403), .B1(n15402), .B2(n6794), .ZN(
        P2_U3510) );
  NOR2_X1 U17000 ( .A1(P3_U3897), .A2(n15417), .ZN(P3_U3150) );
  AOI22_X1 U17001 ( .A1(n15421), .A2(P3_IR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n15413) );
  NOR2_X1 U17002 ( .A1(n15405), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n15410) );
  NAND3_X1 U17003 ( .A1(n15408), .A2(n15407), .A3(n15406), .ZN(n15409) );
  OAI21_X1 U17004 ( .B1(n15411), .B2(n15410), .A(n15409), .ZN(n15412) );
  OAI211_X1 U17005 ( .C1(n15415), .C2(n15414), .A(n15413), .B(n15412), .ZN(
        P3_U3182) );
  AOI21_X1 U17006 ( .B1(P3_ADDR_REG_3__SCAN_IN), .B2(n15417), .A(n15416), .ZN(
        n15433) );
  OAI21_X1 U17007 ( .B1(n15420), .B2(n15419), .A(n15418), .ZN(n15423) );
  AOI22_X1 U17008 ( .A1(n15423), .A2(n15422), .B1(n7258), .B2(n15421), .ZN(
        n15432) );
  OAI221_X1 U17009 ( .B1(n15424), .B2(n15487), .C1(n15424), .C2(n15426), .A(
        n15425), .ZN(n15431) );
  XNOR2_X1 U17010 ( .A(n15427), .B(n15587), .ZN(n15428) );
  NAND2_X1 U17011 ( .A1(n15429), .A2(n15428), .ZN(n15430) );
  NAND4_X1 U17012 ( .A1(n15433), .A2(n15432), .A3(n15431), .A4(n15430), .ZN(
        P3_U3185) );
  XNOR2_X1 U17013 ( .A(n15434), .B(n15439), .ZN(n15580) );
  OAI22_X1 U17014 ( .A1(n15452), .A2(n15492), .B1(n15435), .B2(n15494), .ZN(
        n15441) );
  INV_X1 U17015 ( .A(n15436), .ZN(n15437) );
  AOI211_X1 U17016 ( .C1(n15439), .C2(n15438), .A(n15497), .B(n15437), .ZN(
        n15440) );
  AOI211_X1 U17017 ( .C1(n15580), .C2(n15502), .A(n15441), .B(n15440), .ZN(
        n15576) );
  AOI22_X1 U17018 ( .A1(n15508), .A2(n15442), .B1(n15489), .B2(
        P3_REG2_REG_10__SCAN_IN), .ZN(n15446) );
  NOR2_X1 U17019 ( .A1(n15443), .A2(n15559), .ZN(n15578) );
  AOI22_X1 U17020 ( .A1(n15580), .A2(n15444), .B1(n15485), .B2(n15578), .ZN(
        n15445) );
  OAI211_X1 U17021 ( .C1(n15489), .C2(n15576), .A(n15446), .B(n15445), .ZN(
        P3_U3223) );
  XNOR2_X1 U17022 ( .A(n15447), .B(n15449), .ZN(n15568) );
  XOR2_X1 U17023 ( .A(n15449), .B(n15448), .Z(n15450) );
  OAI222_X1 U17024 ( .A1(n15494), .A2(n15452), .B1(n15492), .B2(n15451), .C1(
        n15497), .C2(n15450), .ZN(n15566) );
  AOI21_X1 U17025 ( .B1(n15521), .B2(n15568), .A(n15566), .ZN(n15457) );
  INV_X1 U17026 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n15456) );
  AND2_X1 U17027 ( .A1(n15453), .A2(n15523), .ZN(n15567) );
  AOI22_X1 U17028 ( .A1(n15485), .A2(n15567), .B1(n15508), .B2(n15454), .ZN(
        n15455) );
  OAI221_X1 U17029 ( .B1(n15489), .B2(n15457), .C1(n15530), .C2(n15456), .A(
        n15455), .ZN(P3_U3225) );
  XNOR2_X1 U17030 ( .A(n15458), .B(n15464), .ZN(n15468) );
  INV_X1 U17031 ( .A(n15468), .ZN(n15557) );
  AOI22_X1 U17032 ( .A1(n15517), .A2(n15460), .B1(n15459), .B2(n15515), .ZN(
        n15467) );
  AND2_X1 U17033 ( .A1(n15462), .A2(n15461), .ZN(n15465) );
  OAI211_X1 U17034 ( .C1(n15465), .C2(n15464), .A(n15463), .B(n15513), .ZN(
        n15466) );
  OAI211_X1 U17035 ( .C1(n15468), .C2(n15481), .A(n15467), .B(n15466), .ZN(
        n15555) );
  AOI21_X1 U17036 ( .B1(n15505), .B2(n15557), .A(n15555), .ZN(n15472) );
  NOR2_X1 U17037 ( .A1(n15469), .A2(n15559), .ZN(n15556) );
  AOI22_X1 U17038 ( .A1(n15556), .A2(n15485), .B1(n15508), .B2(n15470), .ZN(
        n15471) );
  OAI221_X1 U17039 ( .B1(n15489), .B2(n15472), .C1(n15530), .C2(n11076), .A(
        n15471), .ZN(P3_U3227) );
  XNOR2_X1 U17040 ( .A(n15473), .B(n15477), .ZN(n15482) );
  INV_X1 U17041 ( .A(n15482), .ZN(n15545) );
  AOI22_X1 U17042 ( .A1(n15515), .A2(n6592), .B1(n15474), .B2(n15517), .ZN(
        n15480) );
  AND2_X1 U17043 ( .A1(n15499), .A2(n15475), .ZN(n15478) );
  OAI211_X1 U17044 ( .C1(n15478), .C2(n15477), .A(n15476), .B(n15513), .ZN(
        n15479) );
  OAI211_X1 U17045 ( .C1(n15482), .C2(n15481), .A(n15480), .B(n15479), .ZN(
        n15543) );
  AOI21_X1 U17046 ( .B1(n15505), .B2(n15545), .A(n15543), .ZN(n15488) );
  NOR2_X1 U17047 ( .A1(n15483), .A2(n15559), .ZN(n15544) );
  AOI22_X1 U17048 ( .A1(n15544), .A2(n15485), .B1(n15508), .B2(n15484), .ZN(
        n15486) );
  OAI221_X1 U17049 ( .B1(n15489), .B2(n15488), .C1(n15530), .C2(n15487), .A(
        n15486), .ZN(P3_U3230) );
  OAI21_X1 U17050 ( .B1(n15491), .B2(n12067), .A(n15490), .ZN(n15541) );
  OAI22_X1 U17051 ( .A1(n15495), .A2(n15494), .B1(n15493), .B2(n15492), .ZN(
        n15501) );
  NAND3_X1 U17052 ( .A1(n15511), .A2(n12067), .A3(n15496), .ZN(n15498) );
  AOI21_X1 U17053 ( .B1(n15499), .B2(n15498), .A(n15497), .ZN(n15500) );
  AOI211_X1 U17054 ( .C1(n15502), .C2(n15541), .A(n15501), .B(n15500), .ZN(
        n15503) );
  INV_X1 U17055 ( .A(n15503), .ZN(n15539) );
  NOR2_X1 U17056 ( .A1(n7799), .A2(n15559), .ZN(n15540) );
  AOI22_X1 U17057 ( .A1(n15541), .A2(n15505), .B1(n15540), .B2(n15504), .ZN(
        n15506) );
  INV_X1 U17058 ( .A(n15506), .ZN(n15507) );
  AOI211_X1 U17059 ( .C1(n15508), .C2(P3_REG3_REG_2__SCAN_IN), .A(n15539), .B(
        n15507), .ZN(n15509) );
  AOI22_X1 U17060 ( .A1(n15489), .A2(n15510), .B1(n15509), .B2(n15530), .ZN(
        P3_U3231) );
  OAI21_X1 U17061 ( .B1(n10359), .B2(n15512), .A(n15511), .ZN(n15514) );
  NAND2_X1 U17062 ( .A1(n15514), .A2(n15513), .ZN(n15519) );
  AOI22_X1 U17063 ( .A1(n15517), .A2(n6592), .B1(n15516), .B2(n15515), .ZN(
        n15518) );
  NAND2_X1 U17064 ( .A1(n15519), .A2(n15518), .ZN(n15537) );
  XNOR2_X1 U17065 ( .A(n15520), .B(n10359), .ZN(n15533) );
  INV_X1 U17066 ( .A(n15521), .ZN(n15522) );
  NOR2_X1 U17067 ( .A1(n15533), .A2(n15522), .ZN(n15529) );
  NAND2_X1 U17068 ( .A1(n15524), .A2(n15523), .ZN(n15534) );
  OAI22_X1 U17069 ( .A1(n15534), .A2(n15527), .B1(n15526), .B2(n15525), .ZN(
        n15528) );
  NOR3_X1 U17070 ( .A1(n15537), .A2(n15529), .A3(n15528), .ZN(n15531) );
  AOI22_X1 U17071 ( .A1(n15489), .A2(n10175), .B1(n15531), .B2(n15530), .ZN(
        P3_U3232) );
  NOR2_X1 U17072 ( .A1(n15533), .A2(n15532), .ZN(n15536) );
  INV_X1 U17073 ( .A(n15534), .ZN(n15535) );
  NOR3_X1 U17074 ( .A1(n15537), .A2(n15536), .A3(n15535), .ZN(n15584) );
  AOI22_X1 U17075 ( .A1(n15582), .A2(n15584), .B1(n15538), .B2(n8348), .ZN(
        P3_U3393) );
  AOI211_X1 U17076 ( .C1(n15579), .C2(n15541), .A(n15540), .B(n15539), .ZN(
        n15586) );
  INV_X1 U17077 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15542) );
  AOI22_X1 U17078 ( .A1(n15582), .A2(n15586), .B1(n15542), .B2(n8348), .ZN(
        P3_U3396) );
  AOI211_X1 U17079 ( .C1(n15545), .C2(n15579), .A(n15544), .B(n15543), .ZN(
        n15588) );
  INV_X1 U17080 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15546) );
  AOI22_X1 U17081 ( .A1(n15582), .A2(n15588), .B1(n15546), .B2(n8348), .ZN(
        P3_U3399) );
  AOI21_X1 U17082 ( .B1(n15548), .B2(n15579), .A(n15547), .ZN(n15549) );
  AOI22_X1 U17083 ( .A1(n15582), .A2(n15590), .B1(n7813), .B2(n8348), .ZN(
        P3_U3402) );
  AOI211_X1 U17084 ( .C1(n15553), .C2(n15579), .A(n15552), .B(n15551), .ZN(
        n15591) );
  INV_X1 U17085 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15554) );
  AOI22_X1 U17086 ( .A1(n15582), .A2(n15591), .B1(n15554), .B2(n8348), .ZN(
        P3_U3405) );
  AOI211_X1 U17087 ( .C1(n15557), .C2(n15579), .A(n15556), .B(n15555), .ZN(
        n15593) );
  AOI22_X1 U17088 ( .A1(n15582), .A2(n15593), .B1(n15558), .B2(n8348), .ZN(
        P3_U3408) );
  NOR2_X1 U17089 ( .A1(n15560), .A2(n15559), .ZN(n15561) );
  AOI21_X1 U17090 ( .B1(n15562), .B2(n15569), .A(n15561), .ZN(n15563) );
  AND2_X1 U17091 ( .A1(n15564), .A2(n15563), .ZN(n15595) );
  INV_X1 U17092 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15565) );
  AOI22_X1 U17093 ( .A1(n15582), .A2(n15595), .B1(n15565), .B2(n8348), .ZN(
        P3_U3411) );
  AOI211_X1 U17094 ( .C1(n15569), .C2(n15568), .A(n15567), .B(n15566), .ZN(
        n15597) );
  INV_X1 U17095 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15570) );
  AOI22_X1 U17096 ( .A1(n15582), .A2(n15597), .B1(n15570), .B2(n8348), .ZN(
        P3_U3414) );
  AOI21_X1 U17097 ( .B1(n15572), .B2(n15579), .A(n15571), .ZN(n15573) );
  AND2_X1 U17098 ( .A1(n15574), .A2(n15573), .ZN(n15599) );
  AOI22_X1 U17099 ( .A1(n15582), .A2(n15599), .B1(n15575), .B2(n8348), .ZN(
        P3_U3417) );
  INV_X1 U17100 ( .A(n15576), .ZN(n15577) );
  AOI211_X1 U17101 ( .C1(n15580), .C2(n15579), .A(n15578), .B(n15577), .ZN(
        n15602) );
  INV_X1 U17102 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15581) );
  AOI22_X1 U17103 ( .A1(n15582), .A2(n15602), .B1(n15581), .B2(n8348), .ZN(
        P3_U3420) );
  AOI22_X1 U17104 ( .A1(n15603), .A2(n15584), .B1(n15583), .B2(n15600), .ZN(
        P3_U3460) );
  AOI22_X1 U17105 ( .A1(n15603), .A2(n15586), .B1(n15585), .B2(n15600), .ZN(
        P3_U3461) );
  AOI22_X1 U17106 ( .A1(n15603), .A2(n15588), .B1(n15587), .B2(n15600), .ZN(
        P3_U3462) );
  AOI22_X1 U17107 ( .A1(n15603), .A2(n15590), .B1(n15589), .B2(n15600), .ZN(
        P3_U3463) );
  AOI22_X1 U17108 ( .A1(n15603), .A2(n15591), .B1(n7050), .B2(n15600), .ZN(
        P3_U3464) );
  AOI22_X1 U17109 ( .A1(n15603), .A2(n15593), .B1(n15592), .B2(n15600), .ZN(
        P3_U3465) );
  AOI22_X1 U17110 ( .A1(n15603), .A2(n15595), .B1(n15594), .B2(n15600), .ZN(
        P3_U3466) );
  AOI22_X1 U17111 ( .A1(n15603), .A2(n15597), .B1(n15596), .B2(n15600), .ZN(
        P3_U3467) );
  AOI22_X1 U17112 ( .A1(n15603), .A2(n15599), .B1(n15598), .B2(n15600), .ZN(
        P3_U3468) );
  INV_X1 U17113 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15601) );
  AOI22_X1 U17114 ( .A1(n15603), .A2(n15602), .B1(n15601), .B2(n15600), .ZN(
        P3_U3469) );
  AOI21_X1 U17115 ( .B1(n15606), .B2(n15605), .A(n15604), .ZN(SUB_1596_U59) );
  OAI21_X1 U17116 ( .B1(n15609), .B2(n15608), .A(n15607), .ZN(SUB_1596_U58) );
  XNOR2_X1 U17117 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15610), .ZN(SUB_1596_U53)
         );
  OAI21_X1 U17118 ( .B1(n15613), .B2(n15612), .A(n15611), .ZN(SUB_1596_U56) );
  AOI21_X1 U17119 ( .B1(n15616), .B2(n15615), .A(n15614), .ZN(n15617) );
  XOR2_X1 U17120 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15617), .Z(SUB_1596_U60) );
  AOI21_X1 U17121 ( .B1(n15620), .B2(n15619), .A(n15618), .ZN(SUB_1596_U5) );
  INV_X1 U7479 ( .A(n7274), .ZN(n7620) );
  BUF_X2 U7678 ( .A(n7831), .Z(n6607) );
  AND2_X1 U7473 ( .A1(n8364), .A2(n8363), .ZN(n8709) );
  CLKBUF_X1 U8573 ( .A(n9236), .Z(n6847) );
  CLKBUF_X2 U8625 ( .A(n8205), .Z(n12040) );
endmodule

