

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4254, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136;

  NAND2_X1 U4759 ( .A1(n8607), .A2(n8606), .ZN(n8895) );
  AOI21_X1 U4760 ( .B1(n7494), .B2(n7493), .A(n7492), .ZN(n7838) );
  CLKBUF_X1 U4761 ( .A(n6507), .Z(n4259) );
  NAND2_X1 U4762 ( .A1(n4422), .A2(n4421), .ZN(n8113) );
  INV_X1 U4763 ( .A(n4597), .ZN(n6761) );
  BUF_X2 U4764 ( .A(n6606), .Z(n6791) );
  CLKBUF_X3 U4765 ( .A(n5828), .Z(n4274) );
  INV_X2 U4766 ( .A(n5196), .ZN(n5578) );
  INV_X1 U4767 ( .A(n5530), .ZN(n5571) );
  AND2_X1 U4768 ( .A1(n6507), .A2(n6506), .ZN(n7517) );
  AND2_X1 U4769 ( .A1(n4273), .A2(n4256), .ZN(n5085) );
  BUF_X1 U4770 ( .A(n6944), .Z(n4257) );
  NAND2_X1 U4771 ( .A1(n5970), .A2(n5971), .ZN(n8231) );
  MUX2_X1 U4772 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4994), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n4996) );
  XNOR2_X1 U4774 ( .A(n5981), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6000) );
  NAND4_X1 U4775 ( .A1(n5956), .A2(n6244), .A3(n6291), .A4(n5955), .ZN(n6509)
         );
  INV_X1 U4776 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5327) );
  INV_X1 U4777 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5623) );
  OR3_X1 U4778 ( .A1(n5781), .A2(n7870), .A3(n8758), .ZN(n5776) );
  INV_X1 U4779 ( .A(n5776), .ZN(n5778) );
  INV_X1 U4780 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5955) );
  AND2_X1 U4781 ( .A1(n7517), .A2(n6868), .ZN(n6603) );
  AND3_X1 U4782 ( .A1(n5963), .A2(n5962), .A3(n5961), .ZN(n6510) );
  INV_X1 U4783 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6512) );
  INV_X1 U4784 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6291) );
  NAND2_X1 U4785 ( .A1(n4420), .A2(n4419), .ZN(n4967) );
  CLKBUF_X3 U4786 ( .A(n5085), .Z(n4275) );
  INV_X1 U4787 ( .A(n5047), .ZN(n6983) );
  NAND2_X1 U4788 ( .A1(n4845), .A2(n9886), .ZN(n8080) );
  NOR2_X2 U4789 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5363) );
  AND4_X1 U4790 ( .A1(n5363), .A2(n5362), .A3(n5361), .A4(n5327), .ZN(n5364)
         );
  INV_X1 U4791 ( .A(n6791), .ZN(n6744) );
  NOR2_X1 U4792 ( .A1(n6794), .A2(n6586), .ZN(n6614) );
  NAND2_X1 U4793 ( .A1(n9300), .A2(n8301), .ZN(n8296) );
  AOI21_X1 U4794 ( .B1(n9313), .B2(n8224), .A(n8223), .ZN(n9294) );
  AND2_X1 U4795 ( .A1(n4899), .A2(n4513), .ZN(n4361) );
  NAND2_X1 U4796 ( .A1(n5346), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5386) );
  OAI21_X1 U4797 ( .B1(n8726), .B2(n4302), .A(n4494), .ZN(n8626) );
  NOR2_X2 U4798 ( .A1(n8080), .A2(n8085), .ZN(n8079) );
  INV_X1 U4799 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9015) );
  OR2_X1 U4801 ( .A1(n6233), .A2(n6232), .ZN(n6235) );
  XNOR2_X1 U4802 ( .A(n5968), .B(n5967), .ZN(n6524) );
  OAI21_X1 U4803 ( .B1(n7178), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7175), .ZN(
        n7429) );
  NOR2_X1 U4804 ( .A1(n9232), .A2(n9231), .ZN(n9230) );
  NOR2_X2 U4805 ( .A1(n8296), .A2(n9527), .ZN(n9287) );
  BUF_X1 U4806 ( .A(n6612), .Z(n7526) );
  NAND3_X1 U4807 ( .A1(n4511), .A2(n4509), .A3(n4361), .ZN(n5980) );
  AND2_X1 U4808 ( .A1(n8609), .A2(n5549), .ZN(n8261) );
  BUF_X2 U4809 ( .A(n5088), .Z(n5530) );
  NAND3_X2 U4810 ( .A1(n5009), .A2(n5010), .A3(n5011), .ZN(n8289) );
  XNOR2_X1 U4811 ( .A(n4984), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9020) );
  NAND2_X2 U4812 ( .A1(n4727), .A2(n4726), .ZN(n9724) );
  AND4_X1 U4813 ( .A1(n6114), .A2(n6113), .A3(n6112), .A4(n6111), .ZN(n7543)
         );
  BUF_X1 U4814 ( .A(n6000), .Z(n9663) );
  INV_X1 U4815 ( .A(n6508), .ZN(n6530) );
  INV_X1 U4816 ( .A(n5812), .ZN(n7229) );
  INV_X1 U4817 ( .A(n6137), .ZN(n6096) );
  XNOR2_X2 U4818 ( .A(n9724), .B(n6587), .ZN(n7267) );
  INV_X1 U4819 ( .A(n5231), .ZN(n5034) );
  XNOR2_X2 U4820 ( .A(n4369), .B(P1_ADDR_REG_6__SCAN_IN), .ZN(n10116) );
  OAI21_X2 U4821 ( .B1(n8524), .B2(n8523), .A(n8522), .ZN(n8546) );
  NAND2_X1 U4822 ( .A1(n9030), .A2(n7004), .ZN(n4254) );
  NAND2_X2 U4823 ( .A1(n9030), .A2(n7004), .ZN(n5047) );
  OR2_X2 U4824 ( .A1(n7445), .A2(n7529), .ZN(n7648) );
  OAI211_X2 U4825 ( .C1(n6106), .C2(n6938), .A(n6105), .B(n6104), .ZN(n7529)
         );
  NAND2_X2 U4826 ( .A1(n9484), .A2(n9490), .ZN(n9460) );
  NAND2_X2 U4827 ( .A1(n9374), .A2(n4345), .ZN(n4717) );
  NAND2_X2 U4828 ( .A1(n9375), .A2(n9376), .ZN(n9374) );
  AND3_X2 U4829 ( .A1(n5363), .A2(n4978), .A3(n5076), .ZN(n5626) );
  OR2_X2 U4830 ( .A1(n6958), .A2(n5059), .ZN(n5009) );
  NAND2_X2 U4831 ( .A1(n9389), .A2(n8217), .ZN(n9375) );
  XNOR2_X2 U4832 ( .A(n6895), .B(n7126), .ZN(n9240) );
  OAI21_X2 U4833 ( .B1(n7214), .B2(n7212), .A(n7213), .ZN(n7487) );
  XNOR2_X2 U4834 ( .A(n5082), .B(SI_4_), .ZN(n5080) );
  AOI21_X2 U4835 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8572), .A(n8571), .ZN(
        n9820) );
  OAI21_X2 U4836 ( .B1(n7829), .B2(n5851), .A(n4695), .ZN(n4694) );
  INV_X1 U4839 ( .A(n5972), .ZN(n6944) );
  AND4_X4 U4840 ( .A1(n6068), .A2(n6067), .A3(n4962), .A4(n6066), .ZN(n6080)
         );
  XNOR2_X2 U4841 ( .A(n5954), .B(n5961), .ZN(n6508) );
  NAND2_X2 U4842 ( .A1(n6871), .A2(n6872), .ZN(n6870) );
  OAI21_X2 U4843 ( .B1(n7595), .B2(n7594), .A(n4385), .ZN(n6871) );
  OAI22_X2 U4844 ( .A1(n7413), .A2(n7414), .B1(n7423), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7291) );
  OAI21_X2 U4845 ( .B1(n7719), .B2(n7718), .A(n7717), .ZN(n7768) );
  NAND2_X1 U4846 ( .A1(n4738), .A2(n7501), .ZN(n7719) );
  NOR2_X2 U4847 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4813) );
  NOR2_X2 U4848 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4812) );
  XNOR2_X2 U4849 ( .A(n5297), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7491) );
  INV_X2 U4850 ( .A(n5047), .ZN(n4258) );
  NAND2_X1 U4851 ( .A1(n9030), .A2(n7004), .ZN(n4273) );
  OAI21_X2 U4852 ( .B1(n7335), .B2(n7334), .A(n5836), .ZN(n7566) );
  XNOR2_X2 U4853 ( .A(n5607), .B(P2_IR_REG_19__SCAN_IN), .ZN(n7627) );
  NAND2_X2 U4854 ( .A1(n4699), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5607) );
  XNOR2_X2 U4855 ( .A(n6103), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6937) );
  XNOR2_X1 U4856 ( .A(n8591), .B(n5774), .ZN(n8888) );
  NAND2_X1 U4857 ( .A1(n8721), .A2(n8253), .ZN(n8255) );
  NAND2_X1 U4858 ( .A1(n4262), .A2(n4731), .ZN(n8747) );
  NAND2_X1 U4859 ( .A1(n6221), .A2(n6220), .ZN(n9606) );
  OAI21_X1 U4860 ( .B1(n4524), .B2(n4260), .A(n4263), .ZN(n7467) );
  NAND2_X1 U4861 ( .A1(n5789), .A2(n5788), .ZN(n7198) );
  INV_X2 U4862 ( .A(n6612), .ZN(n6792) );
  INV_X1 U4863 ( .A(n7362), .ZN(n4260) );
  BUF_X1 U4864 ( .A(n5833), .Z(n5909) );
  NAND2_X1 U4865 ( .A1(n7135), .A2(n7134), .ZN(n9509) );
  INV_X1 U4866 ( .A(n6817), .ZN(n6406) );
  INV_X2 U4867 ( .A(n7667), .ZN(n4931) );
  AND4_X1 U4868 ( .A1(n6100), .A2(n6099), .A3(n6098), .A4(n6097), .ZN(n7670)
         );
  INV_X1 U4869 ( .A(n7529), .ZN(n7521) );
  INV_X1 U4870 ( .A(n5823), .ZN(n9861) );
  INV_X4 U4871 ( .A(n6080), .ZN(n6587) );
  INV_X1 U4872 ( .A(n6868), .ZN(n6591) );
  MUX2_X1 U4873 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5977), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5979) );
  INV_X2 U4874 ( .A(n5972), .ZN(n5103) );
  NAND2_X1 U4875 ( .A1(n5109), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5152) );
  AND2_X1 U4876 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4272) );
  INV_X1 U4877 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6244) );
  INV_X2 U4878 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  CLKBUF_X2 U4879 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n9813) );
  OAI21_X1 U4880 ( .B1(n9539), .B2(n9735), .A(n4443), .ZN(n4442) );
  NOR2_X1 U4881 ( .A1(n4445), .A2(n4301), .ZN(n4444) );
  AND3_X1 U4882 ( .A1(n4537), .A2(n4911), .A3(n4536), .ZN(n4850) );
  AND4_X1 U4883 ( .A1(n6529), .A2(n7133), .A3(n6528), .A4(n6577), .ZN(n4956)
         );
  NOR2_X1 U4884 ( .A1(n9542), .A2(n4410), .ZN(n9544) );
  OAI21_X1 U4885 ( .B1(n8304), .B2(n8228), .A(n8227), .ZN(n8229) );
  OR2_X1 U4886 ( .A1(n4830), .A2(n6763), .ZN(n9117) );
  AOI21_X1 U4887 ( .B1(n9320), .B2(n9509), .A(n9319), .ZN(n9548) );
  NAND2_X1 U4888 ( .A1(n4412), .A2(n4411), .ZN(n4410) );
  AOI21_X1 U4889 ( .B1(n9277), .B2(n9719), .A(n9711), .ZN(n4661) );
  NAND2_X1 U4890 ( .A1(n8747), .A2(n8252), .ZN(n8721) );
  NAND2_X1 U4891 ( .A1(n9543), .A2(n9626), .ZN(n4411) );
  NAND2_X1 U4892 ( .A1(n6042), .A2(n6041), .ZN(n9550) );
  XNOR2_X1 U4893 ( .A(n5557), .B(n5556), .ZN(n9025) );
  NAND2_X1 U4894 ( .A1(n8768), .A2(n4278), .ZN(n4262) );
  NAND2_X1 U4895 ( .A1(n5469), .A2(n5468), .ZN(n8923) );
  NAND2_X1 U4896 ( .A1(n6337), .A2(n6336), .ZN(n9570) );
  NAND2_X1 U4897 ( .A1(n5454), .A2(n5453), .ZN(n8926) );
  CLKBUF_X1 U4898 ( .A(n8138), .Z(n4364) );
  NAND2_X1 U4899 ( .A1(n8103), .A2(n4740), .ZN(n8849) );
  NAND2_X1 U4900 ( .A1(n8032), .A2(n8031), .ZN(n8103) );
  NAND2_X1 U4901 ( .A1(n5369), .A2(n5368), .ZN(n8952) );
  AND2_X1 U4902 ( .A1(n5477), .A2(n5476), .ZN(n8349) );
  NAND2_X1 U4903 ( .A1(n7154), .A2(n7153), .ZN(n7155) );
  NAND2_X1 U4904 ( .A1(n9904), .A2(n8029), .ZN(n8032) );
  NAND2_X1 U4905 ( .A1(n7994), .A2(n7993), .ZN(n9904) );
  OR2_X1 U4906 ( .A1(n7710), .A2(n7709), .ZN(n4645) );
  AOI21_X1 U4907 ( .B1(n7683), .B2(n7679), .A(n7680), .ZN(n7901) );
  NAND2_X1 U4908 ( .A1(n9226), .A2(n4383), .ZN(n6921) );
  NAND2_X1 U4909 ( .A1(n6266), .A2(n6265), .ZN(n9595) );
  NAND2_X1 U4910 ( .A1(n6017), .A2(n6016), .ZN(n9334) );
  NAND2_X1 U4911 ( .A1(n4714), .A2(n4712), .ZN(n7885) );
  INV_X1 U4912 ( .A(n7893), .ZN(n9620) );
  NAND2_X1 U4913 ( .A1(n5263), .A2(n5262), .ZN(n5859) );
  INV_X1 U4914 ( .A(n4969), .ZN(n4845) );
  NAND2_X1 U4915 ( .A1(n6180), .A2(n6179), .ZN(n9625) );
  AND2_X1 U4916 ( .A1(n6209), .A2(n6208), .ZN(n8057) );
  NAND2_X2 U4917 ( .A1(n5217), .A2(n5216), .ZN(n8987) );
  NAND2_X1 U4918 ( .A1(n6169), .A2(n6168), .ZN(n7936) );
  NAND2_X1 U4919 ( .A1(n7467), .A2(n7466), .ZN(n4739) );
  NAND2_X1 U4920 ( .A1(n5184), .A2(n5207), .ZN(n4453) );
  NAND2_X1 U4921 ( .A1(n4524), .A2(n7202), .ZN(n7361) );
  NAND2_X1 U4922 ( .A1(n9733), .A2(n9725), .ZN(n9502) );
  OAI21_X2 U4923 ( .B1(n7090), .B2(n7066), .A(n7067), .ZN(n7163) );
  NAND2_X1 U4924 ( .A1(n6156), .A2(n6155), .ZN(n7791) );
  INV_X1 U4925 ( .A(n5347), .ZN(n5346) );
  NAND2_X1 U4926 ( .A1(n5211), .A2(n4954), .ZN(n5213) );
  AND2_X1 U4927 ( .A1(n6145), .A2(n6144), .ZN(n9788) );
  NAND2_X1 U4928 ( .A1(n7198), .A2(n7197), .ZN(n4525) );
  INV_X1 U4929 ( .A(n7500), .ZN(n7631) );
  AND2_X1 U4930 ( .A1(n5087), .A2(n5086), .ZN(n7500) );
  AND2_X1 U4931 ( .A1(n6131), .A2(n6130), .ZN(n9781) );
  AOI21_X1 U4932 ( .B1(n7362), .B2(n4264), .A(n7204), .ZN(n4263) );
  NAND2_X1 U4933 ( .A1(n7229), .A2(n7199), .ZN(n5789) );
  INV_X1 U4934 ( .A(n7202), .ZN(n4264) );
  AND2_X1 U4935 ( .A1(n7203), .A2(n9861), .ZN(n7204) );
  AND2_X1 U4936 ( .A1(n9839), .A2(n4360), .ZN(n7102) );
  INV_X1 U4937 ( .A(n7670), .ZN(n7530) );
  OR2_X1 U4938 ( .A1(n8282), .A2(n7328), .ZN(n5818) );
  XNOR2_X1 U4939 ( .A(n9199), .B(n6093), .ZN(n7136) );
  NAND2_X1 U4940 ( .A1(n4336), .A2(n4399), .ZN(n9197) );
  INV_X1 U4941 ( .A(n7543), .ZN(n9198) );
  INV_X1 U4942 ( .A(n5828), .ZN(n5833) );
  AND4_X1 U4943 ( .A1(n6152), .A2(n6151), .A3(n6150), .A4(n6149), .ZN(n7758)
         );
  AND4_X1 U4944 ( .A1(n6164), .A2(n6163), .A3(n6162), .A4(n6161), .ZN(n7910)
         );
  AND2_X1 U4945 ( .A1(n5079), .A2(n5078), .ZN(n9868) );
  AND4_X1 U4946 ( .A1(n5046), .A2(n5045), .A3(n5044), .A4(n5043), .ZN(n7203)
         );
  NAND2_X1 U4947 ( .A1(n4668), .A2(n4309), .ZN(n4667) );
  AND4_X1 U4948 ( .A1(n5133), .A2(n5132), .A3(n5131), .A4(n5130), .ZN(n7771)
         );
  OR2_X1 U4949 ( .A1(n5237), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5259) );
  AND2_X1 U4950 ( .A1(n5163), .A2(n5138), .ZN(n4774) );
  CLKBUF_X1 U4951 ( .A(n6021), .Z(n6397) );
  INV_X2 U4952 ( .A(n5059), .ZN(n5564) );
  NOR2_X1 U4953 ( .A1(n5229), .A2(n4568), .ZN(n4567) );
  AND2_X1 U4954 ( .A1(n4959), .A2(n5210), .ZN(n4954) );
  NAND2_X1 U4955 ( .A1(n9675), .A2(n6518), .ZN(n6868) );
  NAND2_X1 U4956 ( .A1(n4438), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5242) );
  AND2_X2 U4957 ( .A1(n5637), .A2(n7870), .ZN(n9838) );
  XNOR2_X1 U4958 ( .A(n6410), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6507) );
  INV_X2 U4959 ( .A(n6071), .ZN(n6362) );
  INV_X1 U4960 ( .A(n5218), .ZN(n4438) );
  NAND2_X1 U4962 ( .A1(n5952), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6410) );
  XNOR2_X1 U4963 ( .A(n5007), .B(n5008), .ZN(n6958) );
  AND2_X2 U4964 ( .A1(n9663), .A2(n5982), .ZN(n6109) );
  NAND2_X2 U4965 ( .A1(n4987), .A2(n4989), .ZN(n5196) );
  INV_X1 U4966 ( .A(n5059), .ZN(n4261) );
  NAND2_X1 U4967 ( .A1(n6000), .A2(n9666), .ZN(n6071) );
  INV_X1 U4968 ( .A(n9020), .ZN(n4987) );
  INV_X1 U4969 ( .A(n4989), .ZN(n9023) );
  NAND2_X1 U4970 ( .A1(n5608), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5609) );
  XNOR2_X1 U4971 ( .A(n5100), .B(SI_5_), .ZN(n5097) );
  NAND2_X1 U4972 ( .A1(n5187), .A2(n5186), .ZN(n5212) );
  NAND2_X1 U4973 ( .A1(n9016), .A2(n4270), .ZN(n4989) );
  NAND2_X1 U4974 ( .A1(n5614), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5615) );
  XNOR2_X1 U4975 ( .A(n5073), .B(n4558), .ZN(n5072) );
  NAND2_X2 U4976 ( .A1(n4257), .A2(P1_U3084), .ZN(n10109) );
  MUX2_X1 U4977 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5969), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5971) );
  NAND2_X1 U4978 ( .A1(n5970), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5968) );
  OAI21_X1 U4979 ( .B1(n6516), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6515) );
  CLKBUF_X1 U4980 ( .A(n4985), .Z(n9016) );
  AOI21_X1 U4981 ( .B1(n4998), .B2(n4272), .A(n4271), .ZN(n4270) );
  NAND2_X2 U4982 ( .A1(n5972), .A2(P2_U3152), .ZN(n9038) );
  INV_X2 U4983 ( .A(n5034), .ZN(n5164) );
  XNOR2_X1 U4984 ( .A(n5049), .B(n5076), .ZN(n7058) );
  NAND2_X1 U4985 ( .A1(n5154), .A2(n5153), .ZN(n5175) );
  NOR2_X1 U4986 ( .A1(n4326), .A2(n4840), .ZN(n4839) );
  AND2_X1 U4987 ( .A1(n5626), .A2(n4555), .ZN(n4389) );
  INV_X1 U4988 ( .A(n5152), .ZN(n5154) );
  AND2_X1 U4989 ( .A1(n5627), .A2(n5076), .ZN(n5366) );
  NAND3_X1 U4990 ( .A1(n4651), .A2(n4649), .A3(n4648), .ZN(n6904) );
  AND2_X1 U4991 ( .A1(n5976), .A2(n4951), .ZN(n4899) );
  NOR2_X1 U4992 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5951) );
  CLKBUF_X1 U4993 ( .A(n5001), .Z(n5002) );
  INV_X1 U4994 ( .A(n5950), .ZN(n4840) );
  AND3_X2 U4995 ( .A1(n5949), .A2(n5948), .A3(n5947), .ZN(n5966) );
  NAND4_X1 U4996 ( .A1(n5959), .A2(n5958), .A3(n6512), .A4(n5957), .ZN(n5960)
         );
  INV_X1 U4997 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6521) );
  INV_X1 U4998 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5361) );
  NOR2_X1 U4999 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4271) );
  NOR2_X1 U5000 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4971) );
  NOR2_X1 U5001 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4972) );
  INV_X1 U5002 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4650) );
  NOR2_X1 U5003 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4814) );
  INV_X1 U5004 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4267) );
  INV_X1 U5005 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n4266) );
  NAND3_X1 U5006 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5111) );
  AND3_X1 U5007 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6133) );
  INV_X1 U5008 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5610) );
  AND2_X1 U5009 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n5153) );
  INV_X1 U5010 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4456) );
  NOR2_X2 U5011 ( .A1(n4268), .A2(n4265), .ZN(n5625) );
  NAND4_X1 U5012 ( .A1(n5606), .A2(n4701), .A3(n4267), .A4(n4266), .ZN(n4265)
         );
  INV_X2 U5013 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4701) );
  INV_X2 U5014 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5606) );
  NAND4_X1 U5015 ( .A1(n4269), .A2(n5612), .A3(n5327), .A4(n5623), .ZN(n4268)
         );
  INV_X2 U5016 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5612) );
  NOR2_X2 U5017 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4269) );
  XNOR2_X1 U5018 ( .A(n5850), .B(n4365), .ZN(n7829) );
  NAND2_X1 U5019 ( .A1(n4824), .A2(n6730), .ZN(n9130) );
  OAI211_X1 U5020 ( .C1(n4586), .C2(n4589), .A(n4816), .B(n4584), .ZN(n4824)
         );
  XNOR2_X1 U5021 ( .A(n5120), .B(SI_6_), .ZN(n5117) );
  NOR2_X1 U5022 ( .A1(n9163), .A2(n6781), .ZN(n9160) );
  NAND2_X1 U5023 ( .A1(n9454), .A2(n8206), .ZN(n8208) );
  NAND2_X2 U5024 ( .A1(n6870), .A2(n6874), .ZN(n7830) );
  AOI21_X2 U5025 ( .B1(n7838), .B2(n7837), .A(n7836), .ZN(n7839) );
  NOR2_X2 U5026 ( .A1(n5812), .A2(n7328), .ZN(n7316) );
  NOR2_X2 U5027 ( .A1(n6894), .A2(n9230), .ZN(n6895) );
  OAI21_X2 U5028 ( .B1(n8145), .B2(n4721), .A(n4328), .ZN(n9454) );
  AOI211_X2 U5029 ( .C1(n9555), .C2(n9494), .A(n9350), .B(n9349), .ZN(n9351)
         );
  OAI21_X2 U5030 ( .B1(n7566), .B2(n4684), .A(n4682), .ZN(n7595) );
  OAI21_X2 U5031 ( .B1(n7577), .B2(n7575), .A(n7573), .ZN(n7335) );
  NAND2_X1 U5032 ( .A1(n8278), .A2(n5827), .ZN(n7577) );
  OAI21_X2 U5033 ( .B1(n8045), .B2(n8044), .A(n8043), .ZN(n8135) );
  NOR2_X2 U5034 ( .A1(n7478), .A2(n7477), .ZN(n7479) );
  INV_X2 U5035 ( .A(n7322), .ZN(n9853) );
  XNOR2_X1 U5036 ( .A(n7199), .B(n5828), .ZN(n7318) );
  AND2_X2 U5037 ( .A1(n7889), .A2(n7893), .ZN(n7973) );
  NOR2_X2 U5038 ( .A1(n7823), .A2(n9625), .ZN(n7889) );
  XNOR2_X2 U5039 ( .A(n5900), .B(n5899), .ZN(n8320) );
  AOI211_X2 U5040 ( .C1(n9626), .C2(n9527), .A(n9526), .B(n9525), .ZN(n9528)
         );
  OR2_X1 U5041 ( .A1(n8911), .A2(n8631), .ZN(n5760) );
  OR2_X1 U5042 ( .A1(n9543), .A2(n8306), .ZN(n8225) );
  AOI21_X1 U5043 ( .B1(n4627), .B2(n5768), .A(n4626), .ZN(n4625) );
  AOI21_X1 U5044 ( .B1(n4563), .B2(n4296), .A(n4561), .ZN(n4560) );
  INV_X1 U5045 ( .A(n4957), .ZN(n4561) );
  AND2_X1 U5046 ( .A1(n4782), .A2(n4781), .ZN(n4780) );
  INV_X1 U5047 ( .A(n5594), .ZN(n4781) );
  AOI21_X1 U5048 ( .B1(n4782), .B2(n4778), .A(n4777), .ZN(n4776) );
  NOR2_X1 U5049 ( .A1(n5593), .A2(SI_30_), .ZN(n4777) );
  NOR2_X1 U5050 ( .A1(n4785), .A2(n5594), .ZN(n4778) );
  NAND2_X1 U5052 ( .A1(n8258), .A2(n8639), .ZN(n4548) );
  NOR2_X1 U5053 ( .A1(n8306), .A2(n4597), .ZN(n6788) );
  NOR2_X1 U5054 ( .A1(n9296), .A2(n4865), .ZN(n4864) );
  INV_X1 U5055 ( .A(n8196), .ZN(n4865) );
  INV_X1 U5056 ( .A(n5683), .ZN(n4638) );
  OR2_X1 U5057 ( .A1(n7783), .A2(n8458), .ZN(n7986) );
  NAND2_X1 U5058 ( .A1(n4915), .A2(n4460), .ZN(n4459) );
  NAND2_X1 U5059 ( .A1(n5320), .A2(n5319), .ZN(n5339) );
  INV_X1 U5060 ( .A(SI_16_), .ZN(n5319) );
  NAND2_X1 U5061 ( .A1(n5231), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4559) );
  NAND2_X1 U5062 ( .A1(n4382), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4370) );
  INV_X1 U5063 ( .A(n5231), .ZN(n4382) );
  AOI21_X1 U5064 ( .B1(n4622), .B2(n4624), .A(n4337), .ZN(n4621) );
  INV_X1 U5065 ( .A(n4625), .ZN(n4624) );
  NAND2_X1 U5066 ( .A1(n4316), .A2(n4757), .ZN(n5805) );
  OAI21_X1 U5067 ( .B1(n5774), .B2(n5775), .A(n5772), .ZN(n5804) );
  OR2_X1 U5068 ( .A1(n8611), .A2(n8268), .ZN(n5770) );
  NOR2_X1 U5069 ( .A1(n8911), .A2(n8916), .ZN(n4856) );
  NOR2_X1 U5070 ( .A1(n8712), .A2(n4751), .ZN(n4750) );
  NAND2_X1 U5071 ( .A1(n5717), .A2(n5718), .ZN(n8244) );
  OR2_X1 U5072 ( .A1(n8900), .A2(n8632), .ZN(n5763) );
  NAND2_X1 U5073 ( .A1(n4982), .A2(n4981), .ZN(n4983) );
  INV_X1 U5074 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4982) );
  INV_X1 U5075 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U5076 ( .A1(n9666), .A2(n5983), .ZN(n6064) );
  OR2_X1 U5077 ( .A1(n9046), .A2(n9089), .ZN(n6706) );
  OR2_X1 U5078 ( .A1(n4943), .A2(n9334), .ZN(n8195) );
  NOR2_X1 U5079 ( .A1(n4887), .A2(n4884), .ZN(n4883) );
  INV_X1 U5080 ( .A(n8189), .ZN(n4884) );
  INV_X1 U5081 ( .A(n4888), .ZN(n4887) );
  OR2_X1 U5082 ( .A1(n9550), .A2(n9169), .ZN(n9312) );
  NAND2_X1 U5083 ( .A1(n9431), .A2(n4937), .ZN(n4936) );
  NOR2_X1 U5084 ( .A1(n9589), .A2(n9595), .ZN(n4937) );
  AND2_X1 U5085 ( .A1(n8146), .A2(n8144), .ZN(n4723) );
  NAND2_X1 U5086 ( .A1(n6221), .A2(n4575), .ZN(n8203) );
  AND2_X1 U5087 ( .A1(n9511), .A2(n6220), .ZN(n4575) );
  NAND2_X1 U5088 ( .A1(n7605), .A2(n7758), .ZN(n6468) );
  OR2_X1 U5089 ( .A1(n7605), .A2(n7758), .ZN(n7611) );
  NAND2_X1 U5090 ( .A1(n5998), .A2(n5997), .ZN(n9527) );
  NAND2_X1 U5091 ( .A1(n6508), .A2(n9278), .ZN(n6817) );
  INV_X1 U5092 ( .A(n5560), .ZN(n4786) );
  NAND2_X1 U5093 ( .A1(n5543), .A2(n5542), .ZN(n5557) );
  AOI21_X1 U5094 ( .B1(n4761), .B2(n4295), .A(n4759), .ZN(n4758) );
  AND2_X1 U5095 ( .A1(n4769), .A2(n5394), .ZN(n4768) );
  AND2_X1 U5096 ( .A1(n5412), .A2(n5400), .ZN(n5410) );
  XNOR2_X1 U5097 ( .A(n8028), .B(n4274), .ZN(n5850) );
  NAND2_X1 U5098 ( .A1(n4629), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U5099 ( .A1(n4441), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5436) );
  INV_X1 U5100 ( .A(n5779), .ZN(n4617) );
  NAND2_X1 U5101 ( .A1(n4491), .A2(n4490), .ZN(n5590) );
  AOI21_X1 U5102 ( .B1(n8648), .B2(n5571), .A(n5502), .ZN(n8631) );
  NAND2_X1 U5103 ( .A1(n4542), .A2(n4541), .ZN(n8669) );
  AOI21_X1 U5104 ( .B1(n4283), .B2(n4547), .A(n4329), .ZN(n4541) );
  NAND2_X1 U5105 ( .A1(n4532), .A2(n4531), .ZN(n4526) );
  NAND2_X1 U5106 ( .A1(n4922), .A2(n4313), .ZN(n5337) );
  INV_X1 U5107 ( .A(n5085), .ZN(n5331) );
  OR2_X1 U5108 ( .A1(n8968), .A2(n8835), .ZN(n5714) );
  NAND2_X1 U5109 ( .A1(n8849), .A2(n8243), .ZN(n4535) );
  OR2_X1 U5110 ( .A1(n8987), .A2(n8101), .ZN(n8107) );
  OR2_X1 U5111 ( .A1(n4285), .A2(n4743), .ZN(n4539) );
  AND2_X1 U5112 ( .A1(n8424), .A2(n8625), .ZN(n4745) );
  NAND2_X1 U5113 ( .A1(n6999), .A2(n9837), .ZN(n9830) );
  INV_X1 U5114 ( .A(n5048), .ZN(n5627) );
  OAI22_X1 U5115 ( .A1(n6863), .A2(n4597), .B1(n6791), .B2(n8301), .ZN(n6793)
         );
  NAND2_X1 U5116 ( .A1(n7148), .A2(n9769), .ZN(n7454) );
  AND2_X1 U5117 ( .A1(n6506), .A2(n6576), .ZN(n7139) );
  CLKBUF_X1 U5118 ( .A(n6071), .Z(n6393) );
  NAND2_X1 U5119 ( .A1(n7293), .A2(n4435), .ZN(n7552) );
  OR2_X1 U5120 ( .A1(n7296), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4435) );
  AND2_X1 U5121 ( .A1(n6368), .A2(n6367), .ZN(n8306) );
  NAND2_X1 U5122 ( .A1(n9306), .A2(n8195), .ZN(n8197) );
  NAND2_X1 U5123 ( .A1(n8195), .A2(n8196), .ZN(n9315) );
  NOR2_X1 U5124 ( .A1(n4720), .A2(n4719), .ZN(n4718) );
  INV_X1 U5125 ( .A(n4966), .ZN(n4719) );
  NAND2_X1 U5126 ( .A1(n4877), .A2(n4321), .ZN(n9424) );
  OAI22_X1 U5127 ( .A1(n4299), .A2(n4875), .B1(n9476), .B2(n8174), .ZN(n4874)
         );
  OR2_X1 U5128 ( .A1(n7702), .A2(n7133), .ZN(n9789) );
  OAI21_X1 U5129 ( .B1(n5292), .B2(n5291), .A(n5290), .ZN(n5318) );
  OAI21_X1 U5130 ( .B1(n5807), .B2(n4358), .A(n4408), .ZN(n4407) );
  NAND2_X1 U5131 ( .A1(n5782), .A2(P2_B_REG_SCAN_IN), .ZN(n4408) );
  OR2_X1 U5132 ( .A1(n7118), .A2(n9838), .ZN(n4643) );
  INV_X1 U5133 ( .A(n6576), .ZN(n9278) );
  INV_X1 U5134 ( .A(n6468), .ZN(n4506) );
  INV_X1 U5135 ( .A(n5684), .ZN(n4637) );
  AOI21_X1 U5136 ( .B1(n5675), .B2(n5674), .A(n4641), .ZN(n4640) );
  NOR2_X1 U5137 ( .A1(n5647), .A2(n5646), .ZN(n5686) );
  AOI21_X1 U5138 ( .B1(n4507), .B2(n6461), .A(n4505), .ZN(n4504) );
  NOR2_X1 U5139 ( .A1(n7734), .A2(n6817), .ZN(n4505) );
  NAND2_X1 U5140 ( .A1(n4507), .A2(n6467), .ZN(n4501) );
  NAND2_X1 U5141 ( .A1(n4503), .A2(n6406), .ZN(n4502) );
  INV_X1 U5142 ( .A(n6466), .ZN(n4503) );
  AND2_X1 U5143 ( .A1(n4523), .A2(n4610), .ZN(n6262) );
  AND2_X1 U5144 ( .A1(n6218), .A2(n4395), .ZN(n4610) );
  NAND2_X1 U5145 ( .A1(n4611), .A2(n6817), .ZN(n4523) );
  AOI21_X1 U5146 ( .B1(n4705), .B2(n6406), .A(n4396), .ZN(n4395) );
  NOR2_X1 U5147 ( .A1(n4496), .A2(n5422), .ZN(n4493) );
  INV_X1 U5148 ( .A(n4497), .ZN(n4496) );
  INV_X1 U5149 ( .A(n4927), .ZN(n4926) );
  AND2_X1 U5150 ( .A1(n4912), .A2(n5679), .ZN(n4461) );
  INV_X1 U5151 ( .A(n5677), .ZN(n4916) );
  OAI21_X1 U5152 ( .B1(n4521), .B2(n6357), .A(n9358), .ZN(n4520) );
  AND2_X1 U5153 ( .A1(n9315), .A2(n4614), .ZN(n4613) );
  AND2_X1 U5154 ( .A1(n6358), .A2(n9312), .ZN(n4614) );
  NAND2_X1 U5155 ( .A1(n6385), .A2(n6359), .ZN(n4612) );
  INV_X1 U5157 ( .A(n5490), .ZN(n4796) );
  INV_X1 U5158 ( .A(n5519), .ZN(n4795) );
  AND2_X1 U5159 ( .A1(n5517), .A2(n4792), .ZN(n4791) );
  NAND2_X1 U5160 ( .A1(n5378), .A2(n5377), .ZN(n5394) );
  INV_X1 U5161 ( .A(SI_19_), .ZN(n5377) );
  OAI21_X1 U5162 ( .B1(n5103), .B2(P1_DATAO_REG_11__SCAN_IN), .A(n4418), .ZN(
        n5226) );
  OAI21_X1 U5163 ( .B1(n5103), .B2(n4363), .A(n4362), .ZN(n5120) );
  NAND2_X1 U5164 ( .A1(n5103), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4362) );
  OAI21_X1 U5165 ( .B1(n5164), .B2(n4452), .A(n4451), .ZN(n5100) );
  INV_X1 U5166 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n4452) );
  NAND2_X1 U5167 ( .A1(n5164), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4451) );
  AND2_X1 U5168 ( .A1(n4679), .A2(n4677), .ZN(n4676) );
  INV_X1 U5169 ( .A(n5897), .ZN(n4677) );
  INV_X1 U5170 ( .A(n5896), .ZN(n4674) );
  INV_X1 U5171 ( .A(n9838), .ZN(n4668) );
  NOR2_X1 U5172 ( .A1(n5509), .A2(n8425), .ZN(n4439) );
  AOI21_X1 U5173 ( .B1(n4625), .B2(n4628), .A(n4623), .ZN(n4622) );
  INV_X1 U5174 ( .A(n5773), .ZN(n4623) );
  OR2_X1 U5175 ( .A1(n4288), .A2(n5769), .ZN(n4489) );
  OR2_X1 U5176 ( .A1(n8905), .A2(n8424), .ZN(n5639) );
  AND2_X1 U5177 ( .A1(n8712), .A2(n5741), .ZN(n4497) );
  NOR2_X1 U5178 ( .A1(n8942), .A2(n8948), .ZN(n4858) );
  OR2_X1 U5179 ( .A1(n8942), .A2(n8339), .ZN(n5737) );
  OR2_X1 U5180 ( .A1(n8952), .A2(n8372), .ZN(n5727) );
  NAND2_X1 U5181 ( .A1(n4917), .A2(n5646), .ZN(n4466) );
  INV_X1 U5182 ( .A(n4917), .ZN(n4467) );
  NAND2_X1 U5183 ( .A1(n7500), .A2(n8461), .ZN(n5792) );
  AND2_X1 U5184 ( .A1(n4294), .A2(n7469), .ZN(n7193) );
  INV_X1 U5185 ( .A(n5810), .ZN(n7108) );
  NAND2_X1 U5186 ( .A1(n5791), .A2(n7988), .ZN(n4553) );
  OAI21_X1 U5187 ( .B1(n5259), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5274) );
  INV_X1 U5188 ( .A(n5426), .ZN(n4763) );
  INV_X1 U5189 ( .A(n4762), .ZN(n4761) );
  OAI21_X1 U5190 ( .B1(n4765), .B2(n4295), .A(n5444), .ZN(n4762) );
  OAI22_X1 U5191 ( .A1(n6605), .A2(n7670), .B1(n6791), .B2(n7521), .ZN(n6608)
         );
  NAND2_X1 U5192 ( .A1(n9149), .A2(n9148), .ZN(n4820) );
  CLKBUF_X1 U5193 ( .A(n9042), .Z(n9043) );
  INV_X1 U5194 ( .A(n9666), .ZN(n5982) );
  AND2_X1 U5195 ( .A1(n9404), .A2(n9420), .ZN(n8215) );
  OR2_X1 U5196 ( .A1(n9584), .A2(n6720), .ZN(n6414) );
  INV_X1 U5197 ( .A(n4880), .ZN(n4879) );
  OAI21_X1 U5198 ( .B1(n9467), .B2(n4881), .A(n8179), .ZN(n4880) );
  NOR2_X1 U5199 ( .A1(n4709), .A2(n4705), .ZN(n4704) );
  INV_X1 U5200 ( .A(n8141), .ZN(n4709) );
  INV_X1 U5201 ( .A(n8057), .ZN(n8042) );
  OR2_X1 U5202 ( .A1(n9615), .A2(n8136), .ZN(n6417) );
  OR2_X1 U5203 ( .A1(n7895), .A2(n4896), .ZN(n4895) );
  INV_X1 U5204 ( .A(n7817), .ZN(n4896) );
  OR2_X1 U5205 ( .A1(n9620), .A2(n7969), .ZN(n7966) );
  INV_X1 U5206 ( .A(n7804), .ZN(n7794) );
  INV_X1 U5207 ( .A(n4371), .ZN(n4722) );
  NAND2_X1 U5208 ( .A1(n4371), .A2(n4723), .ZN(n8204) );
  AOI21_X1 U5209 ( .B1(n5374), .B2(n4773), .A(n4334), .ZN(n4772) );
  INV_X1 U5210 ( .A(n5359), .ZN(n4773) );
  AOI21_X1 U5211 ( .B1(n4807), .B2(n4805), .A(n4804), .ZN(n4803) );
  NOR2_X1 U5212 ( .A1(n5317), .A2(n4810), .ZN(n4809) );
  INV_X1 U5213 ( .A(n5290), .ZN(n4810) );
  AOI21_X1 U5214 ( .B1(n4809), .B2(n5291), .A(n4808), .ZN(n4807) );
  INV_X1 U5215 ( .A(n5316), .ZN(n4808) );
  INV_X1 U5216 ( .A(n5287), .ZN(n5291) );
  OAI21_X1 U5217 ( .B1(n4567), .B2(n4296), .A(n5248), .ZN(n4564) );
  INV_X1 U5218 ( .A(SI_3_), .ZN(n4558) );
  NAND2_X1 U5219 ( .A1(n5231), .A2(n5055), .ZN(n5056) );
  OR2_X1 U5220 ( .A1(n5281), .A2(n5265), .ZN(n5307) );
  NOR2_X1 U5221 ( .A1(n4665), .A2(n8329), .ZN(n4664) );
  INV_X1 U5222 ( .A(n5881), .ZN(n4665) );
  NAND2_X1 U5223 ( .A1(n4439), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5548) );
  INV_X1 U5224 ( .A(n7567), .ZN(n4685) );
  NAND2_X1 U5225 ( .A1(n4440), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U5226 ( .A1(n5174), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5199) );
  INV_X1 U5227 ( .A(n5175), .ZN(n5174) );
  NAND2_X1 U5228 ( .A1(n4387), .A2(n4386), .ZN(n4385) );
  INV_X1 U5229 ( .A(n5843), .ZN(n4386) );
  INV_X1 U5230 ( .A(n5844), .ZN(n4387) );
  OR3_X1 U5231 ( .A1(n5436), .A2(n8337), .A3(n8404), .ZN(n5455) );
  AND2_X1 U5232 ( .A1(n8336), .A2(n4680), .ZN(n4679) );
  NAND2_X1 U5233 ( .A1(n8393), .A2(n5889), .ZN(n4680) );
  BUF_X1 U5234 ( .A(n5886), .Z(n4413) );
  OR2_X1 U5235 ( .A1(n8346), .A2(n8347), .ZN(n4671) );
  OR2_X1 U5236 ( .A1(n5507), .A2(n9991), .ZN(n5509) );
  INV_X1 U5237 ( .A(n4439), .ZN(n5528) );
  OR3_X1 U5238 ( .A1(n8121), .A2(n9036), .A3(n9034), .ZN(n6999) );
  NAND2_X1 U5239 ( .A1(n7487), .A2(n4455), .ZN(n7842) );
  OR2_X1 U5240 ( .A1(n7491), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4455) );
  AND2_X1 U5241 ( .A1(n4854), .A2(n8263), .ZN(n4853) );
  AOI21_X1 U5242 ( .B1(n8639), .B2(n4550), .A(n4331), .ZN(n4549) );
  INV_X1 U5243 ( .A(n8257), .ZN(n4550) );
  OR2_X1 U5244 ( .A1(n8916), .A2(n8451), .ZN(n8257) );
  AOI21_X1 U5245 ( .B1(n4546), .B2(n4746), .A(n4330), .ZN(n4545) );
  INV_X1 U5246 ( .A(n4750), .ZN(n4546) );
  INV_X1 U5247 ( .A(n4746), .ZN(n4547) );
  NOR2_X1 U5248 ( .A1(n8696), .A2(n4747), .ZN(n4746) );
  INV_X1 U5249 ( .A(n4749), .ZN(n4747) );
  OR2_X1 U5250 ( .A1(n8931), .A2(n8727), .ZN(n4749) );
  NAND2_X1 U5251 ( .A1(n8255), .A2(n4750), .ZN(n4748) );
  OR2_X1 U5252 ( .A1(n8931), .A2(n8340), .ZN(n5748) );
  AND2_X1 U5253 ( .A1(n5748), .A2(n5745), .ZN(n8712) );
  AND2_X1 U5254 ( .A1(n8734), .A2(n5737), .ZN(n8726) );
  NAND2_X1 U5255 ( .A1(n8726), .A2(n5422), .ZN(n8725) );
  NAND2_X1 U5256 ( .A1(n8250), .A2(n4734), .ZN(n4733) );
  INV_X1 U5257 ( .A(n8248), .ZN(n4734) );
  NOR2_X1 U5258 ( .A1(n4736), .A2(n8249), .ZN(n4735) );
  AOI21_X1 U5259 ( .B1(n4471), .B2(n4473), .A(n4469), .ZN(n4468) );
  AND2_X1 U5260 ( .A1(n4528), .A2(n4315), .ZN(n4531) );
  NAND2_X1 U5261 ( .A1(n4530), .A2(n4529), .ZN(n4528) );
  INV_X1 U5262 ( .A(n4534), .ZN(n4532) );
  INV_X1 U5263 ( .A(n8244), .ZN(n8809) );
  AND2_X1 U5264 ( .A1(n8825), .A2(n5313), .ZN(n5314) );
  OR2_X1 U5265 ( .A1(n5859), .A2(n8860), .ZN(n8815) );
  NAND2_X1 U5266 ( .A1(n4437), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5279) );
  INV_X1 U5267 ( .A(n5242), .ZN(n4437) );
  NOR2_X1 U5268 ( .A1(n8106), .A2(n4741), .ZN(n4740) );
  INV_X1 U5269 ( .A(n8102), .ZN(n4741) );
  NOR2_X1 U5270 ( .A1(n4919), .A2(n4918), .ZN(n4917) );
  INV_X1 U5271 ( .A(n4963), .ZN(n4919) );
  INV_X1 U5272 ( .A(n5785), .ZN(n4918) );
  NAND2_X1 U5273 ( .A1(n7982), .A2(n5786), .ZN(n4920) );
  NAND2_X1 U5274 ( .A1(n8028), .A2(n8021), .ZN(n5785) );
  NAND2_X1 U5275 ( .A1(n6964), .A2(n5564), .ZN(n4492) );
  NAND2_X1 U5276 ( .A1(n4462), .A2(n5793), .ZN(n7505) );
  NAND2_X1 U5277 ( .A1(n7470), .A2(n5669), .ZN(n4462) );
  NAND2_X1 U5278 ( .A1(n7505), .A2(n7504), .ZN(n7503) );
  NAND2_X1 U5279 ( .A1(n5062), .A2(n4260), .ZN(n7366) );
  INV_X1 U5280 ( .A(n8871), .ZN(n8831) );
  NAND2_X1 U5281 ( .A1(n4629), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5044) );
  INV_X1 U5282 ( .A(n7193), .ZN(n7466) );
  OR2_X1 U5283 ( .A1(n6985), .A2(n7004), .ZN(n8861) );
  INV_X1 U5284 ( .A(n7102), .ZN(n7197) );
  OR2_X1 U5285 ( .A1(n7106), .A2(n7623), .ZN(n7113) );
  INV_X1 U5286 ( .A(n8861), .ZN(n8819) );
  AND2_X1 U5287 ( .A1(n8647), .A2(n4298), .ZN(n8910) );
  INV_X1 U5288 ( .A(n7636), .ZN(n7626) );
  OR3_X1 U5289 ( .A1(n7625), .A2(n7624), .A3(n7623), .ZN(n7637) );
  AND2_X1 U5290 ( .A1(n5626), .A2(n4635), .ZN(n4634) );
  NOR2_X1 U5291 ( .A1(n4983), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4635) );
  NAND2_X1 U5292 ( .A1(n5617), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U5293 ( .A1(n5615), .A2(n5616), .ZN(n5617) );
  AND2_X1 U5294 ( .A1(n4950), .A2(n4701), .ZN(n4700) );
  OR2_X1 U5295 ( .A1(n5144), .A2(n5143), .ZN(n5325) );
  NAND2_X1 U5296 ( .A1(n6602), .A2(n6601), .ZN(n7309) );
  INV_X1 U5297 ( .A(n4820), .ZN(n4819) );
  AND2_X1 U5298 ( .A1(n4595), .A2(n8008), .ZN(n4594) );
  NAND2_X1 U5299 ( .A1(n4303), .A2(n6667), .ZN(n4595) );
  INV_X1 U5300 ( .A(n6667), .ZN(n4592) );
  NAND2_X1 U5301 ( .A1(n6661), .A2(n6660), .ZN(n7872) );
  OAI22_X1 U5302 ( .A1(n8128), .A2(n6606), .B1(n4597), .B2(n8136), .ZN(n6675)
         );
  NOR2_X1 U5303 ( .A1(n9169), .A2(n4597), .ZN(n6775) );
  INV_X1 U5304 ( .A(n9057), .ZN(n4829) );
  INV_X1 U5305 ( .A(n9116), .ZN(n4827) );
  NAND2_X1 U5306 ( .A1(n6157), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U5307 ( .A1(n4583), .A2(n4325), .ZN(n4587) );
  NAND2_X1 U5308 ( .A1(n6133), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6159) );
  AND2_X1 U5309 ( .A1(n6826), .A2(n9769), .ZN(n6820) );
  AND2_X1 U5310 ( .A1(n6508), .A2(n4259), .ZN(n4515) );
  OR2_X1 U5311 ( .A1(n9517), .A2(n5994), .ZN(n6572) );
  AOI21_X1 U5312 ( .B1(n4605), .B2(n9531), .A(n4606), .ZN(n4604) );
  NAND2_X1 U5313 ( .A1(n6408), .A2(n6409), .ZN(n4606) );
  NAND2_X1 U5314 ( .A1(n4607), .A2(n4609), .ZN(n4605) );
  NAND2_X1 U5315 ( .A1(n6403), .A2(n4518), .ZN(n4601) );
  NOR2_X1 U5316 ( .A1(n4607), .A2(n8228), .ZN(n4518) );
  NAND2_X1 U5317 ( .A1(n6405), .A2(n4397), .ZN(n4603) );
  AND2_X1 U5318 ( .A1(n8227), .A2(n4398), .ZN(n4397) );
  INV_X1 U5319 ( .A(n4609), .ZN(n4398) );
  AND2_X1 U5320 ( .A1(n6345), .A2(n6344), .ZN(n9142) );
  INV_X1 U5321 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n4898) );
  NOR2_X1 U5322 ( .A1(n7418), .A2(n4654), .ZN(n7294) );
  AND2_X1 U5323 ( .A1(n7423), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U5324 ( .A1(n4434), .A2(n4433), .ZN(n4647) );
  INV_X1 U5325 ( .A(n7553), .ZN(n4433) );
  AND2_X1 U5326 ( .A1(n4647), .A2(n4646), .ZN(n7710) );
  NAND2_X1 U5327 ( .A1(n7556), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4646) );
  NAND2_X1 U5328 ( .A1(n9228), .A2(n9227), .ZN(n9226) );
  NOR2_X1 U5329 ( .A1(n9252), .A2(n4409), .ZN(n6902) );
  AND2_X1 U5330 ( .A1(n7288), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4409) );
  NOR2_X1 U5331 ( .A1(n6902), .A2(n6901), .ZN(n9265) );
  OR2_X1 U5332 ( .A1(n9527), .A2(n8305), .ZN(n6498) );
  AND2_X1 U5333 ( .A1(n6389), .A2(n6388), .ZN(n8301) );
  INV_X1 U5334 ( .A(n9333), .ZN(n4449) );
  AOI21_X1 U5335 ( .B1(n4888), .B2(n4886), .A(n4324), .ZN(n4885) );
  NOR2_X1 U5336 ( .A1(n8187), .A2(n4906), .ZN(n4905) );
  INV_X1 U5337 ( .A(n8184), .ZN(n4906) );
  AND2_X1 U5338 ( .A1(n4907), .A2(n8186), .ZN(n4903) );
  OR2_X1 U5339 ( .A1(n8215), .A2(n8214), .ZN(n9405) );
  NAND2_X1 U5340 ( .A1(n9412), .A2(n8183), .ZN(n8185) );
  NAND2_X1 U5341 ( .A1(n4934), .A2(n4933), .ZN(n4932) );
  INV_X1 U5342 ( .A(n4936), .ZN(n4933) );
  AND2_X1 U5343 ( .A1(n6447), .A2(n8212), .ZN(n9418) );
  NAND2_X1 U5344 ( .A1(n6414), .A2(n8210), .ZN(n9434) );
  AND2_X1 U5345 ( .A1(n4966), .A2(n9432), .ZN(n9447) );
  INV_X1 U5346 ( .A(n8177), .ZN(n9468) );
  INV_X1 U5347 ( .A(n4868), .ZN(n4867) );
  AOI21_X1 U5348 ( .B1(n4868), .B2(n4875), .A(n4323), .ZN(n4866) );
  NAND2_X1 U5349 ( .A1(n9468), .A2(n9467), .ZN(n9466) );
  OR2_X1 U5350 ( .A1(n4723), .A2(n4721), .ZN(n4574) );
  INV_X1 U5351 ( .A(n8203), .ZN(n4721) );
  OR2_X1 U5352 ( .A1(n9599), .A2(n6688), .ZN(n9455) );
  INV_X1 U5353 ( .A(n8138), .ZN(n4871) );
  INV_X1 U5354 ( .A(n8137), .ZN(n4876) );
  AND2_X1 U5355 ( .A1(n6416), .A2(n8203), .ZN(n8146) );
  NAND2_X1 U5356 ( .A1(n4897), .A2(n7794), .ZN(n7818) );
  INV_X1 U5357 ( .A(n7795), .ZN(n4897) );
  NOR2_X1 U5358 ( .A1(n4715), .A2(n4713), .ZN(n4712) );
  INV_X1 U5359 ( .A(n7803), .ZN(n4713) );
  AOI21_X1 U5360 ( .B1(n7611), .B2(n6468), .A(n4863), .ZN(n4862) );
  INV_X1 U5361 ( .A(n7603), .ZN(n4863) );
  INV_X1 U5362 ( .A(n9197), .ZN(n7740) );
  INV_X1 U5363 ( .A(n7702), .ZN(n7455) );
  INV_X1 U5364 ( .A(n7139), .ZN(n7460) );
  OR2_X1 U5365 ( .A1(n7454), .A2(n7453), .ZN(n7618) );
  INV_X1 U5366 ( .A(n8128), .ZN(n9615) );
  INV_X1 U5367 ( .A(n9789), .ZN(n9627) );
  OR2_X1 U5368 ( .A1(n6817), .A2(n7133), .ZN(n9632) );
  AND2_X2 U5369 ( .A1(n7455), .A2(n7460), .ZN(n9626) );
  OR2_X1 U5370 ( .A1(n8099), .A2(n8230), .ZN(n6798) );
  AND2_X1 U5371 ( .A1(n8159), .A2(n8099), .ZN(n6518) );
  INV_X1 U5372 ( .A(n6509), .ZN(n4513) );
  NOR2_X1 U5373 ( .A1(n5960), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U5374 ( .A1(n4779), .A2(n4776), .ZN(n5600) );
  NAND2_X1 U5375 ( .A1(n5980), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5981) );
  XNOR2_X1 U5376 ( .A(n5595), .B(n5577), .ZN(n9019) );
  OAI21_X1 U5377 ( .B1(n5557), .B2(n4784), .A(n4782), .ZN(n5595) );
  NAND2_X1 U5378 ( .A1(n4797), .A2(n5490), .ZN(n5518) );
  NAND2_X1 U5379 ( .A1(n4798), .A2(n4792), .ZN(n4797) );
  NAND2_X1 U5380 ( .A1(n4764), .A2(n5426), .ZN(n5446) );
  NAND2_X1 U5381 ( .A1(n5413), .A2(n4765), .ZN(n4764) );
  XNOR2_X1 U5382 ( .A(n5375), .B(n5373), .ZN(n7514) );
  NAND2_X1 U5383 ( .A1(n4566), .A2(n5228), .ZN(n5250) );
  NAND2_X1 U5384 ( .A1(n5213), .A2(n4567), .ZN(n4566) );
  OR2_X1 U5385 ( .A1(n6177), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6206) );
  OR2_X1 U5386 ( .A1(n6119), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U5387 ( .A1(n4650), .A2(P1_IR_REG_1__SCAN_IN), .ZN(n4649) );
  NAND2_X1 U5388 ( .A1(n9659), .A2(P1_IR_REG_1__SCAN_IN), .ZN(n4648) );
  OR2_X1 U5389 ( .A1(n9689), .A2(n10118), .ZN(n4369) );
  NOR2_X1 U5390 ( .A1(n10127), .A2(n9695), .ZN(n9696) );
  AND2_X1 U5391 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9694), .ZN(n9695) );
  INV_X1 U5392 ( .A(n5849), .ZN(n4365) );
  AOI21_X2 U5393 ( .B1(n5571), .B2(P2_REG3_REG_2__SCAN_IN), .A(n4372), .ZN(
        n8282) );
  OR2_X1 U5394 ( .A1(n5065), .A2(n7231), .ZN(n5022) );
  OR2_X1 U5395 ( .A1(n5088), .A2(n7379), .ZN(n5012) );
  AND4_X1 U5396 ( .A1(n5224), .A2(n5223), .A3(n5222), .A4(n5221), .ZN(n8101)
         );
  AND4_X1 U5397 ( .A1(n5285), .A2(n5284), .A3(n5283), .A4(n5282), .ZN(n8834)
         );
  AND3_X1 U5398 ( .A1(n5353), .A2(n5352), .A3(n5351), .ZN(n8415) );
  AND2_X1 U5399 ( .A1(n5421), .A2(n5420), .ZN(n8736) );
  AND2_X1 U5400 ( .A1(n5393), .A2(n5392), .ZN(n8735) );
  AOI21_X1 U5401 ( .B1(n4689), .B2(n4691), .A(n4310), .ZN(n4686) );
  NAND2_X1 U5402 ( .A1(n5931), .A2(n8761), .ZN(n8445) );
  NAND2_X1 U5403 ( .A1(n5301), .A2(n5300), .ZN(n8968) );
  NAND2_X1 U5404 ( .A1(n5780), .A2(n7765), .ZN(n5807) );
  AOI21_X1 U5405 ( .B1(n4618), .B2(n4620), .A(n4617), .ZN(n4616) );
  XNOR2_X1 U5406 ( .A(n4392), .B(n7627), .ZN(n5806) );
  NOR2_X1 U5407 ( .A1(n5803), .A2(n4393), .ZN(n4392) );
  NAND2_X1 U5408 ( .A1(n8898), .A2(n4394), .ZN(n4393) );
  OR2_X1 U5409 ( .A1(n5605), .A2(n4482), .ZN(n4480) );
  NAND2_X1 U5410 ( .A1(n4484), .A2(n5619), .ZN(n4482) );
  NAND2_X1 U5411 ( .A1(n4485), .A2(n4487), .ZN(n4484) );
  NOR2_X1 U5412 ( .A1(n4483), .A2(n5618), .ZN(n4481) );
  AND2_X1 U5413 ( .A1(n4485), .A2(n4346), .ZN(n4483) );
  INV_X1 U5414 ( .A(n8680), .ZN(n8451) );
  INV_X1 U5415 ( .A(n8340), .ZN(n8727) );
  NAND2_X1 U5416 ( .A1(n4702), .A2(n5366), .ZN(n5381) );
  AND2_X1 U5417 ( .A1(n4698), .A2(n5364), .ZN(n4702) );
  XNOR2_X1 U5418 ( .A(n8569), .B(n9822), .ZN(n9815) );
  OR2_X1 U5419 ( .A1(n5932), .A2(n9830), .ZN(n8761) );
  OR2_X1 U5420 ( .A1(n4744), .A2(n4285), .ZN(n4536) );
  NAND2_X1 U5421 ( .A1(n4379), .A2(n9902), .ZN(n4378) );
  INV_X1 U5422 ( .A(n8925), .ZN(n4379) );
  AND2_X1 U5423 ( .A1(n5935), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8018) );
  NAND2_X1 U5424 ( .A1(n4579), .A2(n4582), .ZN(n4578) );
  AND2_X1 U5425 ( .A1(n6866), .A2(n4955), .ZN(n4582) );
  NAND2_X1 U5426 ( .A1(n4580), .A2(n6859), .ZN(n4579) );
  NAND2_X1 U5427 ( .A1(n6029), .A2(n6028), .ZN(n9559) );
  INV_X1 U5428 ( .A(n4815), .ZN(n9066) );
  AOI21_X1 U5429 ( .B1(n9151), .B2(n4821), .A(n4819), .ZN(n4815) );
  NAND2_X1 U5430 ( .A1(n4837), .A2(n6781), .ZN(n4833) );
  NAND2_X1 U5431 ( .A1(n4837), .A2(n4835), .ZN(n4834) );
  NOR2_X1 U5432 ( .A1(n6859), .A2(n6858), .ZN(n4837) );
  AND2_X1 U5433 ( .A1(n6816), .A2(n9165), .ZN(n4836) );
  INV_X1 U5434 ( .A(n8301), .ZN(n9536) );
  INV_X1 U5435 ( .A(n9404), .ZN(n9574) );
  INV_X1 U5436 ( .A(n9373), .ZN(n9564) );
  INV_X1 U5437 ( .A(n9431), .ZN(n9584) );
  INV_X1 U5438 ( .A(n9490), .ZN(n9599) );
  OAI21_X1 U5439 ( .B1(n4517), .B2(n4516), .A(n4514), .ZN(n6529) );
  AND2_X1 U5440 ( .A1(n6572), .A2(n4515), .ZN(n4514) );
  INV_X1 U5441 ( .A(n4603), .ZN(n4516) );
  NAND2_X1 U5442 ( .A1(n4601), .A2(n4604), .ZN(n4517) );
  OR2_X1 U5443 ( .A1(n6823), .A2(n6393), .ZN(n6401) );
  NAND2_X1 U5444 ( .A1(n6039), .A2(n6038), .ZN(n9377) );
  INV_X1 U5445 ( .A(n9142), .ZN(n9408) );
  NAND2_X1 U5446 ( .A1(n7390), .A2(n7391), .ZN(n7389) );
  AND2_X1 U5447 ( .A1(n6923), .A2(n8231), .ZN(n9719) );
  OAI21_X1 U5448 ( .B1(n9702), .B2(n9281), .A(n9280), .ZN(n4663) );
  INV_X1 U5449 ( .A(n9529), .ZN(n4416) );
  INV_X1 U5450 ( .A(n4415), .ZN(n4414) );
  AOI21_X1 U5451 ( .B1(n9525), .B2(n9514), .A(n8236), .ZN(n4415) );
  NAND2_X1 U5452 ( .A1(n4380), .A2(n8303), .ZN(n8295) );
  INV_X1 U5453 ( .A(n8308), .ZN(n9539) );
  INV_X1 U5454 ( .A(n9728), .ZN(n9499) );
  NAND2_X1 U5455 ( .A1(n9318), .A2(n9317), .ZN(n9319) );
  AND2_X1 U5456 ( .A1(n6058), .A2(n6057), .ZN(n7893) );
  CLKBUF_X1 U5457 ( .A(n9766), .Z(n9754) );
  INV_X1 U5458 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4598) );
  OAI21_X1 U5459 ( .B1(n6263), .B2(n4841), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4599) );
  NOR2_X1 U5460 ( .A1(n9950), .A2(n4359), .ZN(n9948) );
  INV_X2 U5461 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9702) );
  NOR2_X1 U5462 ( .A1(n6406), .A2(n4508), .ZN(n4507) );
  NAND2_X1 U5463 ( .A1(n4500), .A2(n4499), .ZN(n6176) );
  AOI21_X1 U5464 ( .B1(n4276), .B2(n4281), .A(n4339), .ZN(n4499) );
  NAND2_X1 U5465 ( .A1(n6141), .A2(n4276), .ZN(n4500) );
  NOR2_X1 U5466 ( .A1(n4638), .A2(n4637), .ZN(n4636) );
  NAND2_X1 U5467 ( .A1(n4912), .A2(n5680), .ZN(n4639) );
  NAND2_X1 U5468 ( .A1(n6417), .A2(n7963), .ZN(n4396) );
  OAI21_X1 U5469 ( .B1(n4281), .B2(n6141), .A(n4276), .ZN(n6203) );
  NAND2_X1 U5470 ( .A1(n5721), .A2(n4632), .ZN(n5734) );
  NOR2_X1 U5471 ( .A1(n5726), .A2(n4633), .ZN(n4632) );
  INV_X1 U5472 ( .A(n5727), .ZN(n4633) );
  AND2_X1 U5473 ( .A1(n5727), .A2(n5731), .ZN(n4631) );
  NOR4_X1 U5474 ( .A1(n5794), .A2(n4460), .A3(n7767), .A4(n7472), .ZN(n5795)
         );
  NAND2_X1 U5475 ( .A1(n5792), .A2(n7469), .ZN(n5657) );
  NAND2_X1 U5476 ( .A1(n8463), .A2(n9861), .ZN(n5668) );
  NAND2_X1 U5477 ( .A1(n7765), .A2(n5809), .ZN(n5810) );
  NOR2_X1 U5478 ( .A1(n8774), .A2(n5725), .ZN(n4474) );
  AND2_X1 U5479 ( .A1(n7986), .A2(n7985), .ZN(n7987) );
  INV_X1 U5480 ( .A(n8178), .ZN(n4881) );
  INV_X1 U5481 ( .A(n5463), .ZN(n4759) );
  INV_X1 U5482 ( .A(n5395), .ZN(n4771) );
  AND2_X1 U5483 ( .A1(n4772), .A2(n4771), .ZN(n4767) );
  NOR2_X1 U5484 ( .A1(n4806), .A2(n4801), .ZN(n4800) );
  INV_X1 U5485 ( .A(n5256), .ZN(n4801) );
  INV_X1 U5486 ( .A(n4809), .ZN(n4805) );
  INV_X1 U5487 ( .A(n4960), .ZN(n4804) );
  INV_X1 U5488 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5341) );
  INV_X1 U5489 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5251) );
  INV_X1 U5490 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5232) );
  AND2_X1 U5491 ( .A1(n5861), .A2(n5860), .ZN(n8355) );
  XNOR2_X1 U5492 ( .A(n5828), .B(n9853), .ZN(n5819) );
  NAND2_X1 U5493 ( .A1(n4488), .A2(n4322), .ZN(n4491) );
  NAND2_X1 U5494 ( .A1(n5775), .A2(n5809), .ZN(n4490) );
  NOR2_X1 U5495 ( .A1(n8905), .A2(n4855), .ZN(n4854) );
  INV_X1 U5496 ( .A(n4856), .ZN(n4855) );
  AND2_X1 U5497 ( .A1(n4495), .A2(n4923), .ZN(n4494) );
  NAND2_X1 U5498 ( .A1(n5478), .A2(n4493), .ZN(n4495) );
  AND2_X1 U5499 ( .A1(n8696), .A2(n5748), .ZN(n4927) );
  INV_X1 U5500 ( .A(n4297), .ZN(n4736) );
  NOR2_X1 U5501 ( .A1(n5859), .A2(n8977), .ZN(n4861) );
  OAI211_X1 U5502 ( .C1(n7505), .C2(n4913), .A(n4461), .B(n4459), .ZN(n4458)
         );
  INV_X1 U5503 ( .A(n5657), .ZN(n5669) );
  NAND2_X1 U5504 ( .A1(n7120), .A2(n9853), .ZN(n5664) );
  NAND2_X1 U5505 ( .A1(n8282), .A2(n7322), .ZN(n7363) );
  NOR2_X1 U5506 ( .A1(n4406), .A2(n9905), .ZN(n4852) );
  AOI21_X1 U5507 ( .B1(n4474), .B2(n4477), .A(n4472), .ZN(n4471) );
  INV_X1 U5508 ( .A(n5733), .ZN(n4472) );
  INV_X1 U5509 ( .A(n4474), .ZN(n4473) );
  NAND2_X1 U5510 ( .A1(n4914), .A2(n5679), .ZN(n7773) );
  NAND2_X1 U5511 ( .A1(n7503), .A2(n4915), .ZN(n4914) );
  AOI21_X1 U5512 ( .B1(n9829), .B2(n9835), .A(n9836), .ZN(n7625) );
  INV_X1 U5513 ( .A(n4983), .ZN(n4555) );
  NAND2_X1 U5514 ( .A1(n5076), .A2(n10062), .ZN(n4697) );
  OR2_X1 U5515 ( .A1(n5214), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U5516 ( .A1(n5001), .A2(n4974), .ZN(n5048) );
  INV_X1 U5517 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4974) );
  INV_X1 U5518 ( .A(n9297), .ZN(n6863) );
  CLKBUF_X1 U5519 ( .A(n7901), .Z(n7903) );
  INV_X1 U5520 ( .A(n6794), .ZN(n6784) );
  NOR2_X1 U5521 ( .A1(n4597), .A2(n9049), .ZN(n6683) );
  NAND2_X1 U5522 ( .A1(n6503), .A2(n4608), .ZN(n4607) );
  AND2_X1 U5523 ( .A1(n6498), .A2(n6817), .ZN(n4608) );
  NAND2_X1 U5524 ( .A1(n6567), .A2(n4308), .ZN(n4609) );
  NOR2_X1 U5525 ( .A1(n4317), .A2(n4612), .ZN(n4522) );
  NAND2_X1 U5526 ( .A1(n7713), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4644) );
  NOR2_X1 U5527 ( .A1(n4943), .A2(n4940), .ZN(n4939) );
  INV_X1 U5528 ( .A(n4941), .ZN(n4940) );
  NOR2_X1 U5529 ( .A1(n9550), .A2(n4942), .ZN(n4941) );
  NOR2_X1 U5530 ( .A1(n8193), .A2(n4889), .ZN(n4888) );
  INV_X1 U5531 ( .A(n8192), .ZN(n4889) );
  INV_X1 U5532 ( .A(n8191), .ZN(n4886) );
  OR2_X1 U5533 ( .A1(n9570), .A2(n9142), .ZN(n6448) );
  NAND2_X1 U5534 ( .A1(n4879), .A2(n4881), .ZN(n4878) );
  NOR2_X1 U5535 ( .A1(n4874), .A2(n8176), .ZN(n4868) );
  AND2_X1 U5536 ( .A1(n4948), .A2(n4282), .ZN(n4947) );
  INV_X1 U5537 ( .A(n4895), .ZN(n4892) );
  INV_X1 U5538 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U5539 ( .A1(n9781), .A2(n4931), .ZN(n4930) );
  AND2_X1 U5540 ( .A1(n6467), .A2(n6542), .ZN(n4729) );
  NAND2_X1 U5541 ( .A1(n6107), .A2(n6542), .ZN(n6125) );
  OR2_X1 U5542 ( .A1(n9736), .A2(n6811), .ZN(n7449) );
  AOI21_X1 U5543 ( .B1(n4785), .B2(n4783), .A(n4355), .ZN(n4782) );
  INV_X1 U5544 ( .A(n5556), .ZN(n4783) );
  NAND2_X1 U5545 ( .A1(n4710), .A2(n4280), .ZN(n5970) );
  AND2_X1 U5546 ( .A1(n5964), .A2(n6052), .ZN(n4710) );
  INV_X1 U5547 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4711) );
  NAND2_X1 U5548 ( .A1(n4790), .A2(n4788), .ZN(n5541) );
  AND2_X1 U5549 ( .A1(n4789), .A2(n4794), .ZN(n4788) );
  AOI21_X1 U5550 ( .B1(n5517), .B2(n4796), .A(n4795), .ZN(n4794) );
  AND2_X1 U5551 ( .A1(n5542), .A2(n5524), .ZN(n5540) );
  NOR2_X1 U5552 ( .A1(n5503), .A2(n4793), .ZN(n4792) );
  INV_X1 U5553 ( .A(n5482), .ZN(n4793) );
  AND2_X1 U5554 ( .A1(n6511), .A2(n6510), .ZN(n6519) );
  INV_X1 U5555 ( .A(SI_15_), .ZN(n9985) );
  NOR2_X1 U5556 ( .A1(n5427), .A2(n4766), .ZN(n4765) );
  INV_X1 U5557 ( .A(n5412), .ZN(n4766) );
  NAND2_X1 U5558 ( .A1(n5398), .A2(n5397), .ZN(n5412) );
  INV_X1 U5559 ( .A(SI_20_), .ZN(n5397) );
  NOR2_X1 U5560 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5950) );
  XNOR2_X1 U5561 ( .A(n5288), .B(SI_14_), .ZN(n5287) );
  INV_X1 U5562 ( .A(n5225), .ZN(n5229) );
  INV_X1 U5563 ( .A(n5212), .ZN(n4568) );
  XNOR2_X1 U5564 ( .A(n5226), .B(SI_11_), .ZN(n5225) );
  AND2_X1 U5565 ( .A1(n5207), .A2(n5206), .ZN(n5208) );
  NAND2_X1 U5566 ( .A1(n5075), .A2(n5074), .ZN(n4557) );
  INV_X1 U5567 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4753) );
  AND2_X1 U5568 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  NAND2_X1 U5569 ( .A1(n5264), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5281) );
  INV_X1 U5570 ( .A(n5279), .ZN(n5264) );
  AOI21_X1 U5571 ( .B1(n4679), .B2(n4675), .A(n4674), .ZN(n4673) );
  NOR2_X1 U5572 ( .A1(n5897), .A2(n5889), .ZN(n4675) );
  NAND2_X1 U5573 ( .A1(n4629), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U5574 ( .A1(n5875), .A2(n4968), .ZN(n4666) );
  INV_X1 U5575 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7847) );
  INV_X1 U5576 ( .A(n4440), .ZN(n5470) );
  AOI21_X1 U5577 ( .B1(n4692), .B2(n4694), .A(n4690), .ZN(n4689) );
  INV_X1 U5578 ( .A(n8002), .ZN(n4690) );
  INV_X1 U5579 ( .A(n4692), .ZN(n4691) );
  OR2_X1 U5580 ( .A1(n5940), .A2(n5939), .ZN(n8426) );
  OR2_X1 U5581 ( .A1(n5933), .A2(n9830), .ZN(n5940) );
  AOI21_X1 U5582 ( .B1(n4621), .B2(n4619), .A(n4327), .ZN(n4618) );
  INV_X1 U5583 ( .A(n4622), .ZN(n4619) );
  INV_X1 U5584 ( .A(n4621), .ZN(n4620) );
  NOR2_X1 U5585 ( .A1(n5805), .A2(n5804), .ZN(n4394) );
  NAND2_X1 U5586 ( .A1(n4757), .A2(n8758), .ZN(n4487) );
  INV_X1 U5587 ( .A(n4486), .ZN(n4485) );
  OAI22_X1 U5588 ( .A1(n5604), .A2(n4487), .B1(n4757), .B2(n8758), .ZN(n4486)
         );
  OR2_X1 U5589 ( .A1(n5196), .A2(n4988), .ZN(n4993) );
  NAND2_X1 U5590 ( .A1(n4629), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4556) );
  AOI21_X1 U5591 ( .B1(n7034), .B2(n7033), .A(n7032), .ZN(n8468) );
  OAI21_X1 U5592 ( .B1(n8468), .B2(n8466), .A(n8467), .ZN(n8481) );
  AOI21_X1 U5593 ( .B1(n8481), .B2(n8480), .A(n8479), .ZN(n8496) );
  AOI21_X1 U5594 ( .B1(n8509), .B2(n8508), .A(n8507), .ZN(n8524) );
  OR2_X1 U5595 ( .A1(n7055), .A2(n7056), .ZN(n7154) );
  AND2_X1 U5596 ( .A1(n7842), .A2(n4454), .ZN(n4425) );
  AND2_X1 U5597 ( .A1(n7496), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n7836) );
  INV_X1 U5598 ( .A(n8607), .ZN(n8592) );
  AND2_X1 U5599 ( .A1(n5535), .A2(n5534), .ZN(n8424) );
  OR2_X1 U5600 ( .A1(n8622), .A2(n5530), .ZN(n5535) );
  NAND2_X1 U5601 ( .A1(n8682), .A2(n4854), .ZN(n8620) );
  NAND2_X1 U5602 ( .A1(n8682), .A2(n8666), .ZN(n8660) );
  AND2_X1 U5603 ( .A1(n5515), .A2(n5514), .ZN(n8680) );
  NAND2_X1 U5604 ( .A1(n8770), .A2(n8259), .ZN(n8755) );
  NAND2_X1 U5605 ( .A1(n8770), .A2(n4858), .ZN(n4970) );
  INV_X1 U5606 ( .A(n4441), .ZN(n5403) );
  INV_X1 U5607 ( .A(n8787), .ZN(n4420) );
  NAND2_X1 U5608 ( .A1(n8872), .A2(n4861), .ZN(n8839) );
  AOI21_X1 U5609 ( .B1(n4305), .B2(n4467), .A(n4464), .ZN(n4463) );
  INV_X1 U5610 ( .A(n5783), .ZN(n4464) );
  INV_X1 U5611 ( .A(n8024), .ZN(n4422) );
  AND2_X1 U5612 ( .A1(n8107), .A2(n4963), .ZN(n8030) );
  NAND2_X1 U5613 ( .A1(n5171), .A2(n5170), .ZN(n8085) );
  OR2_X1 U5614 ( .A1(n8088), .A2(n7990), .ZN(n8074) );
  AND2_X1 U5615 ( .A1(n5644), .A2(n5684), .ZN(n8088) );
  NAND2_X1 U5616 ( .A1(n4847), .A2(n4846), .ZN(n4969) );
  INV_X1 U5617 ( .A(n7781), .ZN(n4847) );
  INV_X1 U5618 ( .A(n8761), .ZN(n8876) );
  NAND2_X1 U5619 ( .A1(n7366), .A2(n4312), .ZN(n7470) );
  NAND2_X1 U5620 ( .A1(n4843), .A2(n9861), .ZN(n7478) );
  INV_X1 U5621 ( .A(n4844), .ZN(n4843) );
  NAND2_X1 U5622 ( .A1(n7228), .A2(n7227), .ZN(n7364) );
  INV_X1 U5623 ( .A(n8293), .ZN(n4360) );
  AND2_X1 U5624 ( .A1(n8267), .A2(n5763), .ZN(n8598) );
  INV_X1 U5625 ( .A(n9905), .ZN(n8988) );
  NAND2_X1 U5626 ( .A1(n9838), .A2(n7765), .ZN(n9907) );
  NAND2_X1 U5627 ( .A1(n9838), .A2(n5939), .ZN(n9905) );
  INV_X1 U5628 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5616) );
  AND2_X1 U5629 ( .A1(n6858), .A2(n9165), .ZN(n4580) );
  OAI21_X1 U5630 ( .B1(n5413), .B2(n4295), .A(n4761), .ZN(n5464) );
  AND2_X1 U5631 ( .A1(n6664), .A2(n6663), .ZN(n7874) );
  NAND2_X1 U5632 ( .A1(n4823), .A2(n4822), .ZN(n4821) );
  INV_X1 U5633 ( .A(n9148), .ZN(n4822) );
  INV_X1 U5634 ( .A(n9149), .ZN(n4823) );
  NOR2_X1 U5635 ( .A1(n9142), .A2(n4597), .ZN(n6743) );
  AND2_X1 U5636 ( .A1(n6700), .A2(n6699), .ZN(n9106) );
  NAND2_X1 U5637 ( .A1(n9056), .A2(n9057), .ZN(n9118) );
  INV_X1 U5638 ( .A(n7674), .ZN(n4596) );
  INV_X1 U5639 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6181) );
  INV_X1 U5640 ( .A(n6592), .ZN(n6593) );
  NAND2_X1 U5641 ( .A1(n6603), .A2(n9201), .ZN(n6590) );
  OR2_X1 U5642 ( .A1(n4585), .A2(n4587), .ZN(n4584) );
  AND2_X1 U5643 ( .A1(n9065), .A2(n4817), .ZN(n4816) );
  NAND2_X1 U5644 ( .A1(n4818), .A2(n4820), .ZN(n4817) );
  INV_X1 U5645 ( .A(n4821), .ZN(n4818) );
  INV_X1 U5646 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6232) );
  INV_X1 U5647 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6210) );
  INV_X1 U5648 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6298) );
  AND2_X1 U5649 ( .A1(n6306), .A2(n6305), .ZN(n6720) );
  NOR2_X1 U5650 ( .A1(n6899), .A2(P1_U3084), .ZN(n7281) );
  OAI22_X1 U5651 ( .A1(n7343), .A2(n7344), .B1(n6946), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n9214) );
  AND2_X1 U5652 ( .A1(n7347), .A2(n6915), .ZN(n9220) );
  NAND2_X1 U5653 ( .A1(n7245), .A2(n4653), .ZN(n7176) );
  OR2_X1 U5654 ( .A1(n6916), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4653) );
  AND2_X1 U5655 ( .A1(n7433), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4655) );
  AND2_X1 U5656 ( .A1(n9272), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U5657 ( .A1(n5974), .A2(n5973), .ZN(n9288) );
  AND3_X2 U5658 ( .A1(n9353), .A2(n4938), .A3(n4939), .ZN(n9300) );
  AND2_X1 U5659 ( .A1(n6006), .A2(n6005), .ZN(n8305) );
  INV_X1 U5660 ( .A(n6009), .ZN(n6391) );
  NAND2_X1 U5661 ( .A1(n9316), .A2(n9510), .ZN(n9318) );
  NAND2_X1 U5662 ( .A1(n9353), .A2(n4939), .ZN(n9307) );
  OR2_X1 U5663 ( .A1(n9559), .A2(n9122), .ZN(n8219) );
  NAND2_X1 U5664 ( .A1(n9353), .A2(n9344), .ZN(n9339) );
  AOI21_X1 U5665 ( .B1(n4903), .B2(n4902), .A(n4320), .ZN(n4901) );
  INV_X1 U5666 ( .A(n4903), .ZN(n4900) );
  INV_X1 U5667 ( .A(n4905), .ZN(n4902) );
  NOR2_X1 U5668 ( .A1(n8214), .A2(n4725), .ZN(n4724) );
  NOR2_X1 U5669 ( .A1(n9460), .A2(n4935), .ZN(n9442) );
  INV_X1 U5670 ( .A(n4937), .ZN(n4935) );
  NAND2_X1 U5671 ( .A1(n8204), .A2(n8203), .ZN(n9473) );
  AND2_X1 U5672 ( .A1(n7973), .A2(n4945), .ZN(n9484) );
  NOR2_X1 U5673 ( .A1(n4946), .A2(n9606), .ZN(n4945) );
  INV_X1 U5674 ( .A(n4947), .ZN(n4946) );
  AOI21_X1 U5675 ( .B1(n8141), .B2(n4708), .A(n4707), .ZN(n4706) );
  INV_X1 U5676 ( .A(n8037), .ZN(n4708) );
  NAND2_X1 U5677 ( .A1(n7973), .A2(n4947), .ZN(n9497) );
  NAND2_X1 U5678 ( .A1(n8038), .A2(n8037), .ZN(n8142) );
  AND2_X1 U5679 ( .A1(n7973), .A2(n8057), .ZN(n8049) );
  NAND2_X1 U5680 ( .A1(n7967), .A2(n7966), .ZN(n8038) );
  AND4_X1 U5681 ( .A1(n6063), .A2(n6062), .A3(n6061), .A4(n6060), .ZN(n7969)
         );
  AND4_X1 U5682 ( .A1(n6201), .A2(n6200), .A3(n6199), .A4(n6198), .ZN(n8136)
         );
  NAND2_X1 U5683 ( .A1(n6108), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6198) );
  AND2_X1 U5684 ( .A1(n7815), .A2(n7803), .ZN(n7804) );
  OR2_X1 U5685 ( .A1(n7797), .A2(n7936), .ZN(n7823) );
  NAND2_X1 U5686 ( .A1(n4404), .A2(n4403), .ZN(n7797) );
  INV_X1 U5687 ( .A(n7616), .ZN(n4404) );
  NAND2_X1 U5688 ( .A1(n4929), .A2(n4928), .ZN(n7616) );
  NOR2_X1 U5689 ( .A1(n7605), .A2(n4930), .ZN(n4928) );
  NOR2_X1 U5690 ( .A1(n7648), .A2(n4930), .ZN(n7745) );
  NOR2_X1 U5691 ( .A1(n7648), .A2(n7667), .ZN(n7647) );
  NAND2_X1 U5692 ( .A1(n6108), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U5693 ( .A1(n6542), .A2(n6463), .ZN(n7533) );
  NOR2_X1 U5694 ( .A1(n9201), .A2(n7701), .ZN(n7268) );
  INV_X1 U5695 ( .A(n9541), .ZN(n4412) );
  NOR2_X1 U5696 ( .A1(n4722), .A2(n6240), .ZN(n4949) );
  INV_X1 U5697 ( .A(n9626), .ZN(n9787) );
  OR2_X1 U5698 ( .A1(n7149), .A2(n7454), .ZN(n7693) );
  AND2_X1 U5699 ( .A1(n6052), .A2(n5966), .ZN(n4512) );
  XNOR2_X1 U5700 ( .A(n5576), .B(n5563), .ZN(n9022) );
  NAND2_X1 U5701 ( .A1(n4787), .A2(n5560), .ZN(n5576) );
  CLKBUF_X1 U5702 ( .A(n6524), .Z(n7410) );
  XNOR2_X1 U5703 ( .A(n5541), .B(n5540), .ZN(n9029) );
  NAND2_X1 U5704 ( .A1(n4798), .A2(n5482), .ZN(n5504) );
  XNOR2_X1 U5705 ( .A(n5484), .B(n5479), .ZN(n8098) );
  NAND2_X1 U5706 ( .A1(n5953), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U5707 ( .A1(n5951), .A2(n4842), .ZN(n4841) );
  INV_X1 U5708 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4842) );
  OAI21_X1 U5709 ( .B1(n5360), .B2(n5373), .A(n4772), .ZN(n5396) );
  NAND2_X1 U5710 ( .A1(n4802), .A2(n4807), .ZN(n5338) );
  NAND2_X1 U5711 ( .A1(n5292), .A2(n4809), .ZN(n4802) );
  XNOR2_X1 U5712 ( .A(n5183), .B(n5182), .ZN(n6969) );
  OR2_X1 U5713 ( .A1(n6153), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n6165) );
  XNOR2_X1 U5714 ( .A(n5161), .B(n5162), .ZN(n6964) );
  CLKBUF_X1 U5715 ( .A(n5119), .Z(n5104) );
  INV_X1 U5716 ( .A(n5072), .ZN(n5070) );
  INV_X1 U5717 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10089) );
  AOI21_X1 U5718 ( .B1(n4368), .B2(n4367), .A(n4366), .ZN(n9688) );
  AND2_X1 U5719 ( .A1(n10089), .A2(n7399), .ZN(n4366) );
  INV_X1 U5720 ( .A(n10136), .ZN(n4367) );
  INV_X1 U5721 ( .A(n10135), .ZN(n4368) );
  INV_X1 U5722 ( .A(n4369), .ZN(n9690) );
  NAND2_X1 U5723 ( .A1(n4666), .A2(n5881), .ZN(n8330) );
  OR2_X1 U5724 ( .A1(n6847), .A2(n6846), .ZN(n6848) );
  NAND2_X1 U5725 ( .A1(n4306), .A2(n4685), .ZN(n4684) );
  AND4_X1 U5726 ( .A1(n5180), .A2(n5179), .A3(n5178), .A4(n5177), .ZN(n7984)
         );
  AND2_X1 U5727 ( .A1(n5443), .A2(n5442), .ZN(n8340) );
  AND2_X1 U5728 ( .A1(n5409), .A2(n5408), .ZN(n8339) );
  NAND2_X1 U5729 ( .A1(n4678), .A2(n5889), .ZN(n8335) );
  NAND2_X1 U5730 ( .A1(n4413), .A2(n5885), .ZN(n4678) );
  NAND2_X1 U5731 ( .A1(n7830), .A2(n4693), .ZN(n4688) );
  AND3_X1 U5732 ( .A1(n5311), .A2(n5310), .A3(n5309), .ZN(n8835) );
  NAND2_X1 U5733 ( .A1(n5402), .A2(n5401), .ZN(n8942) );
  OAI21_X1 U5734 ( .B1(n4413), .B2(n4681), .A(n4679), .ZN(n8399) );
  AND4_X1 U5735 ( .A1(n5247), .A2(n5246), .A3(n5245), .A4(n5244), .ZN(n8862)
         );
  AND4_X1 U5736 ( .A1(n5205), .A2(n5204), .A3(n5203), .A4(n5202), .ZN(n8021)
         );
  AOI21_X1 U5737 ( .B1(n7829), .B2(n7830), .A(n5851), .ZN(n7915) );
  CLKBUF_X1 U5738 ( .A(n7566), .Z(n4388) );
  NOR2_X1 U5739 ( .A1(n4388), .A2(n7567), .ZN(n7565) );
  AND2_X1 U5740 ( .A1(n5528), .A2(n5498), .ZN(n8648) );
  AND4_X1 U5741 ( .A1(n5272), .A2(n5271), .A3(n5270), .A4(n5269), .ZN(n8860)
         );
  OR2_X1 U5742 ( .A1(n8426), .A2(n8859), .ZN(n8441) );
  INV_X1 U5743 ( .A(n8349), .ZN(n8690) );
  NAND2_X1 U5744 ( .A1(n4629), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5068) );
  INV_X1 U5745 ( .A(n7203), .ZN(n8463) );
  OR2_X2 U5746 ( .A1(n6999), .A2(n6869), .ZN(n8464) );
  NAND2_X1 U5747 ( .A1(n4424), .A2(n4423), .ZN(n7016) );
  OR2_X1 U5748 ( .A1(n7020), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4424) );
  NAND2_X1 U5749 ( .A1(n7016), .A2(n7017), .ZN(n7034) );
  NAND2_X1 U5750 ( .A1(n8542), .A2(n8543), .ZN(n8541) );
  AOI21_X1 U5751 ( .B1(n8556), .B2(n7076), .A(n7075), .ZN(n7087) );
  AND2_X1 U5752 ( .A1(n7088), .A2(n7089), .ZN(n7090) );
  XNOR2_X1 U5753 ( .A(n7842), .B(n4454), .ZN(n7488) );
  AND2_X1 U5754 ( .A1(n6987), .A2(n6986), .ZN(n8585) );
  XNOR2_X1 U5755 ( .A(n4417), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8580) );
  OR2_X1 U5756 ( .A1(n9814), .A2(n8570), .ZN(n4417) );
  INV_X1 U5757 ( .A(n9807), .ZN(n9823) );
  NAND2_X1 U5758 ( .A1(n5602), .A2(n5601), .ZN(n5774) );
  AOI21_X1 U5759 ( .B1(n9019), .B2(n4261), .A(n4953), .ZN(n8593) );
  OR2_X1 U5760 ( .A1(n4406), .A2(n8605), .ZN(n8606) );
  NAND2_X1 U5761 ( .A1(n4911), .A2(n8602), .ZN(n8614) );
  NOR2_X1 U5762 ( .A1(n4744), .A2(n4743), .ZN(n4742) );
  OAI21_X1 U5763 ( .B1(n8667), .B2(n4551), .A(n4549), .ZN(n8617) );
  NAND2_X1 U5764 ( .A1(n5497), .A2(n5496), .ZN(n8911) );
  NAND2_X1 U5765 ( .A1(n8640), .A2(n8639), .ZN(n8638) );
  NAND2_X1 U5766 ( .A1(n8667), .A2(n8257), .ZN(n8640) );
  NAND2_X1 U5767 ( .A1(n4544), .A2(n4545), .ZN(n8674) );
  OR2_X1 U5768 ( .A1(n8255), .A2(n4547), .ZN(n4544) );
  NAND2_X1 U5769 ( .A1(n4375), .A2(n4373), .ZN(n8921) );
  INV_X1 U5770 ( .A(n4374), .ZN(n4373) );
  OAI211_X1 U5771 ( .C1(n8677), .C2(n8678), .A(n8653), .B(n8871), .ZN(n4375)
         );
  OAI21_X1 U5772 ( .B1(n8680), .B2(n8859), .A(n8679), .ZN(n4374) );
  NAND2_X1 U5773 ( .A1(n4748), .A2(n4746), .ZN(n8699) );
  NAND2_X1 U5774 ( .A1(n4748), .A2(n4749), .ZN(n8697) );
  AND2_X1 U5775 ( .A1(n8716), .A2(n8715), .ZN(n8934) );
  AND2_X1 U5776 ( .A1(n8725), .A2(n5741), .ZN(n8711) );
  AOI21_X1 U5777 ( .B1(n4278), .B2(n4733), .A(n4732), .ZN(n4731) );
  NAND2_X1 U5778 ( .A1(n4730), .A2(n4278), .ZN(n8746) );
  OR2_X1 U5779 ( .A1(n8768), .A2(n4733), .ZN(n4730) );
  NAND2_X1 U5780 ( .A1(n4921), .A2(n5735), .ZN(n8733) );
  NAND2_X1 U5781 ( .A1(n4737), .A2(n4297), .ZN(n8750) );
  OR2_X1 U5782 ( .A1(n8768), .A2(n8248), .ZN(n4737) );
  NAND2_X1 U5783 ( .A1(n4475), .A2(n5722), .ZN(n8775) );
  NAND2_X1 U5784 ( .A1(n5337), .A2(n4476), .ZN(n4475) );
  NAND2_X1 U5785 ( .A1(n8806), .A2(n8245), .ZN(n8793) );
  NAND2_X1 U5786 ( .A1(n4535), .A2(n4534), .ZN(n8808) );
  INV_X1 U5787 ( .A(n8242), .ZN(n4533) );
  NAND2_X1 U5788 ( .A1(n8103), .A2(n8102), .ZN(n8105) );
  NAND2_X1 U5789 ( .A1(n4920), .A2(n4917), .ZN(n8108) );
  NAND2_X1 U5790 ( .A1(n6971), .A2(n5564), .ZN(n5195) );
  NAND2_X1 U5791 ( .A1(n7503), .A2(n5677), .ZN(n7723) );
  NAND2_X1 U5792 ( .A1(n4739), .A2(n7468), .ZN(n7502) );
  NAND2_X1 U5793 ( .A1(n7366), .A2(n5654), .ZN(n7192) );
  OR2_X1 U5794 ( .A1(n7113), .A2(n7112), .ZN(n8687) );
  AND2_X1 U5795 ( .A1(n8772), .A2(n7111), .ZN(n8765) );
  INV_X1 U5796 ( .A(n8687), .ZN(n8884) );
  INV_X2 U5797 ( .A(n8772), .ZN(n8886) );
  NAND2_X1 U5798 ( .A1(n8772), .A2(n7109), .ZN(n8854) );
  AND2_X1 U5799 ( .A1(n5635), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9837) );
  NAND2_X1 U5800 ( .A1(n4985), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4984) );
  INV_X1 U5801 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9039) );
  INV_X1 U5802 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8119) );
  XNOR2_X1 U5803 ( .A(n5624), .B(n5623), .ZN(n8121) );
  NAND2_X1 U5804 ( .A1(n5622), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5624) );
  INV_X1 U5805 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8173) );
  INV_X1 U5806 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U5807 ( .A1(n5611), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5584) );
  INV_X1 U5808 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7766) );
  INV_X1 U5809 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7643) );
  INV_X1 U5810 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7437) );
  INV_X1 U5811 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7287) );
  OR2_X1 U5812 ( .A1(n5330), .A2(n5329), .ZN(n7921) );
  INV_X1 U5813 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7129) );
  INV_X1 U5814 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10071) );
  INV_X1 U5815 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6977) );
  INV_X1 U5816 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6965) );
  OR2_X1 U5817 ( .A1(n6868), .A2(n6880), .ZN(n6928) );
  AND4_X1 U5818 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n7688)
         );
  CLKBUF_X1 U5819 ( .A(n7872), .Z(n7873) );
  AOI21_X1 U5820 ( .B1(n4594), .B2(n4592), .A(n4335), .ZN(n4591) );
  INV_X1 U5821 ( .A(n4594), .ZN(n4593) );
  NAND2_X1 U5822 ( .A1(n6108), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U5823 ( .A1(n6278), .A2(n6277), .ZN(n9589) );
  OR2_X1 U5824 ( .A1(n6763), .A2(n4829), .ZN(n4828) );
  NAND2_X1 U5825 ( .A1(n4827), .A2(n4826), .ZN(n4825) );
  NAND2_X1 U5826 ( .A1(n6763), .A2(n4829), .ZN(n4826) );
  NAND2_X1 U5827 ( .A1(n4832), .A2(n6610), .ZN(n7673) );
  OAI21_X1 U5828 ( .B1(n7873), .B2(n4303), .A(n6667), .ZN(n8009) );
  INV_X1 U5829 ( .A(n9178), .ZN(n9155) );
  NAND2_X1 U5830 ( .A1(n4588), .A2(n4590), .ZN(n9151) );
  INV_X1 U5831 ( .A(n4587), .ZN(n4590) );
  NAND2_X1 U5832 ( .A1(n6829), .A2(n7188), .ZN(n9167) );
  AND2_X1 U5833 ( .A1(n6051), .A2(n6050), .ZN(n9169) );
  OR2_X1 U5834 ( .A1(n9326), .A2(n6393), .ZN(n6051) );
  INV_X1 U5835 ( .A(n9152), .ZN(n9180) );
  INV_X1 U5836 ( .A(n6506), .ZN(n7133) );
  AND2_X1 U5837 ( .A1(n4604), .A2(n7143), .ZN(n4602) );
  INV_X1 U5838 ( .A(n8306), .ZN(n9316) );
  INV_X1 U5839 ( .A(n9169), .ZN(n9348) );
  OR2_X1 U5840 ( .A1(n9370), .A2(n6393), .ZN(n6356) );
  INV_X1 U5841 ( .A(n6720), .ZN(n9450) );
  NAND2_X1 U5842 ( .A1(n6255), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6187) );
  INV_X1 U5843 ( .A(n4400), .ZN(n4399) );
  OAI21_X1 U5844 ( .B1(n6132), .B2(n4898), .A(n6139), .ZN(n4400) );
  CLKBUF_X2 U5845 ( .A(P1_U4006), .Z(n9200) );
  OAI21_X1 U5846 ( .B1(n6904), .B2(n6883), .A(n4652), .ZN(n7241) );
  NAND2_X1 U5847 ( .A1(n6904), .A2(n6883), .ZN(n4652) );
  NAND2_X1 U5848 ( .A1(n7241), .A2(n7240), .ZN(n7239) );
  OAI21_X1 U5849 ( .B1(n6937), .B2(n6909), .A(n4384), .ZN(n7391) );
  NAND2_X1 U5850 ( .A1(n6937), .A2(n6909), .ZN(n4384) );
  OR2_X1 U5851 ( .A1(n7395), .A2(n6912), .ZN(n7396) );
  AOI21_X1 U5852 ( .B1(n9218), .B2(n7251), .A(n7252), .ZN(n7254) );
  INV_X1 U5853 ( .A(n4647), .ZN(n7551) );
  OAI22_X1 U5854 ( .A1(n7549), .A2(n7550), .B1(n7556), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7706) );
  INV_X1 U5855 ( .A(n4645), .ZN(n7708) );
  NOR2_X1 U5856 ( .A1(n9240), .A2(n10016), .ZN(n9239) );
  NAND2_X1 U5857 ( .A1(n4658), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U5858 ( .A1(n6896), .A2(n4658), .ZN(n4656) );
  INV_X1 U5859 ( .A(n9253), .ZN(n4658) );
  NOR2_X1 U5860 ( .A1(n6922), .A2(n9241), .ZN(n9257) );
  AOI21_X1 U5861 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9272), .A(n9271), .ZN(
        n9716) );
  INV_X1 U5862 ( .A(n9281), .ZN(n9718) );
  NAND2_X1 U5863 ( .A1(n5993), .A2(n5992), .ZN(n9517) );
  INV_X1 U5864 ( .A(n9288), .ZN(n9524) );
  NAND2_X1 U5865 ( .A1(n9299), .A2(n9298), .ZN(n9542) );
  NAND2_X1 U5866 ( .A1(n8197), .A2(n8196), .ZN(n9293) );
  AOI21_X1 U5867 ( .B1(n4448), .B2(n9509), .A(n4446), .ZN(n9553) );
  OAI21_X1 U5868 ( .B1(n6862), .B2(n9474), .A(n4447), .ZN(n4446) );
  XNOR2_X1 U5869 ( .A(n9332), .B(n4449), .ZN(n4448) );
  NAND2_X1 U5870 ( .A1(n4890), .A2(n8192), .ZN(n9338) );
  NAND2_X1 U5871 ( .A1(n9352), .A2(n8191), .ZN(n4890) );
  AND2_X1 U5872 ( .A1(n6348), .A2(n6347), .ZN(n9373) );
  NAND2_X1 U5873 ( .A1(n4904), .A2(n4903), .ZN(n9382) );
  NAND2_X1 U5874 ( .A1(n8185), .A2(n4905), .ZN(n4904) );
  NAND2_X1 U5875 ( .A1(n8213), .A2(n8212), .ZN(n9406) );
  AND2_X1 U5876 ( .A1(n6321), .A2(n6320), .ZN(n9404) );
  AND2_X1 U5877 ( .A1(n6296), .A2(n6295), .ZN(n9431) );
  CLKBUF_X1 U5878 ( .A(n9424), .Z(n9425) );
  NAND2_X1 U5879 ( .A1(n9466), .A2(n8178), .ZN(n9441) );
  INV_X1 U5880 ( .A(n4874), .ZN(n4873) );
  NAND2_X1 U5881 ( .A1(n4871), .A2(n4870), .ZN(n4869) );
  AND2_X1 U5882 ( .A1(n6250), .A2(n6249), .ZN(n9490) );
  NAND2_X1 U5883 ( .A1(n4364), .A2(n4299), .ZN(n4872) );
  NAND2_X1 U5884 ( .A1(n4364), .A2(n8137), .ZN(n9496) );
  AND2_X1 U5885 ( .A1(n6194), .A2(n6193), .ZN(n8128) );
  NAND2_X1 U5886 ( .A1(n7818), .A2(n7817), .ZN(n7896) );
  OR2_X1 U5887 ( .A1(n6101), .A2(n6958), .ZN(n4727) );
  OR2_X1 U5888 ( .A1(n6124), .A2(n7244), .ZN(n4728) );
  INV_X1 U5889 ( .A(n9502), .ZN(n9462) );
  INV_X2 U5890 ( .A(n9799), .ZN(n9801) );
  INV_X1 U5891 ( .A(n4402), .ZN(n4401) );
  INV_X2 U5892 ( .A(n9795), .ZN(n9796) );
  NOR2_X1 U5893 ( .A1(n9738), .A2(n9737), .ZN(n9766) );
  AND2_X1 U5894 ( .A1(n6868), .A2(n6523), .ZN(n9769) );
  INV_X1 U5895 ( .A(n9769), .ZN(n9738) );
  AND2_X1 U5896 ( .A1(n5966), .A2(n4510), .ZN(n4509) );
  AND2_X1 U5897 ( .A1(n6510), .A2(n6052), .ZN(n4511) );
  XNOR2_X1 U5898 ( .A(n6514), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9675) );
  XNOR2_X1 U5899 ( .A(n6515), .B(P1_IR_REG_25__SCAN_IN), .ZN(n8159) );
  INV_X1 U5900 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10033) );
  INV_X1 U5901 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7731) );
  INV_X1 U5902 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7641) );
  INV_X1 U5903 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7290) );
  INV_X1 U5904 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7023) );
  INV_X1 U5905 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6982) );
  XNOR2_X1 U5906 ( .A(n6056), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7423) );
  INV_X1 U5907 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6968) );
  OR2_X1 U5908 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  AND2_X1 U5909 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9688), .ZN(n10117) );
  NOR2_X1 U5910 ( .A1(n9697), .A2(n10124), .ZN(n9955) );
  NOR2_X1 U5911 ( .A1(n4432), .A2(n4431), .ZN(n4430) );
  NOR2_X1 U5912 ( .A1(n9987), .A2(n9990), .ZN(n4431) );
  INV_X1 U5913 ( .A(n9967), .ZN(n4432) );
  AOI21_X1 U5914 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9943), .ZN(n9942) );
  NAND2_X1 U5915 ( .A1(n10053), .A2(n4429), .ZN(n4428) );
  INV_X1 U5916 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n4429) );
  OAI21_X1 U5917 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9931), .ZN(n10121) );
  OAI21_X1 U5918 ( .B1(n8625), .B2(n8432), .A(n5943), .ZN(n5944) );
  AND2_X1 U5919 ( .A1(n4480), .A2(n4479), .ZN(n4390) );
  INV_X1 U5920 ( .A(n4407), .ZN(n4642) );
  INV_X1 U5921 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n4909) );
  NAND2_X1 U5922 ( .A1(n4377), .A2(n4376), .ZN(P2_U3512) );
  NAND2_X1 U5923 ( .A1(n9912), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n4376) );
  AOI21_X1 U5924 ( .B1(n6860), .B2(n9165), .A(n4578), .ZN(n4576) );
  AND2_X1 U5925 ( .A1(n6859), .A2(n9165), .ZN(n4581) );
  NAND2_X1 U5926 ( .A1(n6860), .A2(n4836), .ZN(n6837) );
  INV_X1 U5927 ( .A(n4663), .ZN(n4662) );
  AOI21_X1 U5928 ( .B1(n4416), .B2(n9733), .A(n4414), .ZN(n8237) );
  INV_X1 U5929 ( .A(n4442), .ZN(n8310) );
  AOI21_X1 U5930 ( .B1(n9537), .B2(n9494), .A(n8309), .ZN(n4443) );
  NOR2_X1 U5931 ( .A1(n9548), .A2(n9735), .ZN(n9321) );
  NAND2_X1 U5932 ( .A1(n4573), .A2(n4571), .ZN(P1_U3519) );
  OR2_X1 U5933 ( .A1(n9796), .A2(n4572), .ZN(n4571) );
  NAND2_X1 U5934 ( .A1(n9637), .A2(n9796), .ZN(n4573) );
  INV_X1 U5935 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n4572) );
  AND2_X1 U5936 ( .A1(n4279), .A2(n4504), .ZN(n4276) );
  XNOR2_X1 U5937 ( .A(n4599), .B(n4598), .ZN(n6576) );
  AND2_X1 U5938 ( .A1(n4861), .A2(n4860), .ZN(n4277) );
  INV_X2 U5940 ( .A(n6021), .ZN(n6255) );
  NAND2_X1 U5941 ( .A1(n5774), .A2(n5775), .ZN(n4757) );
  NAND2_X1 U5942 ( .A1(n8675), .A2(n5478), .ZN(n8653) );
  OR2_X1 U5943 ( .A1(n4735), .A2(n8251), .ZN(n4278) );
  AND2_X1 U5944 ( .A1(n6468), .A2(n7611), .ZN(n4279) );
  AND4_X1 U5945 ( .A1(n6510), .A2(n5966), .A3(n4951), .A4(n4711), .ZN(n4280)
         );
  AND2_X1 U5946 ( .A1(n4501), .A2(n4502), .ZN(n4281) );
  INV_X1 U5947 ( .A(n8212), .ZN(n4725) );
  AND2_X1 U5948 ( .A1(n8128), .A2(n8057), .ZN(n4282) );
  AND2_X1 U5949 ( .A1(n4545), .A2(n4543), .ZN(n4283) );
  OR2_X1 U5950 ( .A1(n8896), .A2(n8993), .ZN(n4284) );
  OR2_X1 U5951 ( .A1(n4626), .A2(n4284), .ZN(n4285) );
  INV_X1 U5952 ( .A(n7966), .ZN(n4705) );
  AND2_X1 U5953 ( .A1(n6008), .A2(n6007), .ZN(n9311) );
  INV_X1 U5954 ( .A(n9311), .ZN(n4943) );
  AND2_X1 U5955 ( .A1(n5852), .A2(n5853), .ZN(n4286) );
  INV_X1 U5956 ( .A(n4875), .ZN(n4870) );
  NAND2_X1 U5957 ( .A1(n4300), .A2(n8139), .ZN(n4875) );
  AOI21_X1 U5958 ( .B1(n7286), .B2(n5564), .A(n5332), .ZN(n8804) );
  INV_X1 U5959 ( .A(n8804), .ZN(n8962) );
  AND2_X1 U5960 ( .A1(n8710), .A2(n5748), .ZN(n4287) );
  AND2_X1 U5961 ( .A1(n5763), .A2(n5770), .ZN(n4288) );
  AND2_X1 U5962 ( .A1(n4857), .A2(n4858), .ZN(n4289) );
  AND2_X1 U5963 ( .A1(n4961), .A2(n4958), .ZN(n4290) );
  AND2_X1 U5964 ( .A1(n8246), .A2(n8245), .ZN(n4291) );
  NAND2_X1 U5965 ( .A1(n7973), .A2(n4282), .ZN(n8150) );
  NAND2_X1 U5966 ( .A1(n4714), .A2(n7800), .ZN(n4292) );
  NOR2_X1 U5967 ( .A1(n9926), .A2(n5569), .ZN(n4293) );
  OR2_X1 U5968 ( .A1(n9626), .A2(n6814), .ZN(n9186) );
  XNOR2_X1 U5969 ( .A(n5584), .B(n5612), .ZN(n7870) );
  INV_X2 U5970 ( .A(n6096), .ZN(n6394) );
  OR2_X1 U5971 ( .A1(n8462), .A2(n9868), .ZN(n4294) );
  OR2_X1 U5972 ( .A1(n5445), .A2(n4763), .ZN(n4295) );
  OR2_X1 U5973 ( .A1(n4565), .A2(n5249), .ZN(n4296) );
  OR2_X1 U5974 ( .A1(n8773), .A2(n8372), .ZN(n4297) );
  NAND2_X1 U5975 ( .A1(n8682), .A2(n4856), .ZN(n4298) );
  NAND2_X1 U5976 ( .A1(n4465), .A2(n4463), .ZN(n8814) );
  NAND2_X1 U5977 ( .A1(n5760), .A2(n8627), .ZN(n8639) );
  INV_X1 U5978 ( .A(n8639), .ZN(n4551) );
  NOR2_X1 U5979 ( .A1(n8140), .A2(n4876), .ZN(n4299) );
  OR2_X1 U5980 ( .A1(n9606), .A2(n9511), .ZN(n4300) );
  NOR2_X1 U5981 ( .A1(n9534), .A2(n9533), .ZN(n4301) );
  OR2_X1 U5982 ( .A1(n4924), .A2(n4496), .ZN(n4302) );
  AND2_X1 U5983 ( .A1(n7875), .A2(n7874), .ZN(n4303) );
  AND2_X1 U5984 ( .A1(n5679), .A2(n5678), .ZN(n5791) );
  INV_X1 U5985 ( .A(n4915), .ZN(n4913) );
  NOR2_X1 U5986 ( .A1(n4916), .A2(n5676), .ZN(n4915) );
  AND2_X1 U5987 ( .A1(n5714), .A2(n5713), .ZN(n8825) );
  INV_X1 U5988 ( .A(n8825), .ZN(n4530) );
  INV_X1 U5989 ( .A(n5373), .ZN(n5374) );
  INV_X1 U5990 ( .A(n8207), .ZN(n4720) );
  OAI21_X1 U5991 ( .B1(n5213), .B2(n4296), .A(n4563), .ZN(n5273) );
  NAND2_X1 U5992 ( .A1(n8208), .A2(n8207), .ZN(n9446) );
  NAND2_X1 U5993 ( .A1(n4922), .A2(n5714), .ZN(n8798) );
  INV_X1 U5994 ( .A(n4413), .ZN(n8392) );
  NAND2_X1 U5995 ( .A1(n8190), .A2(n8189), .ZN(n9352) );
  NAND2_X1 U5996 ( .A1(n4838), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U5997 ( .A1(n8185), .A2(n8184), .ZN(n9397) );
  NAND2_X1 U5998 ( .A1(n4920), .A2(n5785), .ZN(n8020) );
  NAND2_X1 U5999 ( .A1(n4869), .A2(n4873), .ZN(n9478) );
  AND2_X1 U6000 ( .A1(n4535), .A2(n4533), .ZN(n4304) );
  AND2_X1 U6001 ( .A1(n4466), .A2(n5689), .ZN(n4305) );
  NAND2_X1 U6002 ( .A1(n5842), .A2(n5841), .ZN(n4306) );
  INV_X1 U6003 ( .A(n8143), .ZN(n4707) );
  NAND2_X1 U6004 ( .A1(n4492), .A2(n5149), .ZN(n7783) );
  AND2_X1 U6005 ( .A1(n9217), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4307) );
  INV_X1 U6006 ( .A(n9511), .ZN(n9476) );
  NAND2_X1 U6007 ( .A1(n4830), .A2(n6763), .ZN(n9056) );
  AND2_X1 U6008 ( .A1(n6500), .A2(n6406), .ZN(n4308) );
  AND2_X1 U6009 ( .A1(n6019), .A2(n6018), .ZN(n9344) );
  INV_X1 U6010 ( .A(n9344), .ZN(n4942) );
  XNOR2_X1 U6011 ( .A(n8926), .B(n8713), .ZN(n8696) );
  OR2_X1 U6012 ( .A1(n8028), .A2(n8021), .ZN(n5786) );
  INV_X1 U6013 ( .A(n8745), .ZN(n4732) );
  AND2_X1 U6014 ( .A1(n4669), .A2(n7870), .ZN(n4309) );
  NAND2_X1 U6015 ( .A1(n5277), .A2(n5276), .ZN(n8977) );
  AND2_X1 U6016 ( .A1(n5763), .A2(n5641), .ZN(n8265) );
  INV_X1 U6017 ( .A(n8265), .ZN(n4743) );
  AND2_X1 U6018 ( .A1(n5855), .A2(n5854), .ZN(n4310) );
  NAND2_X1 U6019 ( .A1(n6052), .A2(n5966), .ZN(n6191) );
  NOR2_X1 U6020 ( .A1(n9239), .A2(n6896), .ZN(n4311) );
  AND2_X1 U6021 ( .A1(n4294), .A2(n5654), .ZN(n4312) );
  INV_X1 U6022 ( .A(n8602), .ZN(n8603) );
  NAND2_X1 U6023 ( .A1(n5506), .A2(n5505), .ZN(n8916) );
  INV_X1 U6024 ( .A(n9531), .ZN(n9532) );
  NAND2_X1 U6025 ( .A1(n6498), .A2(n6567), .ZN(n9531) );
  AND2_X1 U6026 ( .A1(n5718), .A2(n5714), .ZN(n4313) );
  OR2_X1 U6027 ( .A1(n9536), .A2(n6863), .ZN(n8226) );
  NAND2_X1 U6028 ( .A1(n6420), .A2(n7800), .ZN(n7801) );
  NAND2_X1 U6029 ( .A1(n5383), .A2(n5382), .ZN(n8948) );
  AND2_X1 U6030 ( .A1(n7613), .A2(n4716), .ZN(n4314) );
  AND2_X1 U6031 ( .A1(n8654), .A2(n5750), .ZN(n8678) );
  INV_X1 U6032 ( .A(n8678), .ZN(n4543) );
  AND2_X1 U6033 ( .A1(n8244), .A2(n8807), .ZN(n4315) );
  NAND2_X1 U6034 ( .A1(n8593), .A2(n8599), .ZN(n4316) );
  INV_X1 U6035 ( .A(n8905), .ZN(n8625) );
  NAND2_X1 U6036 ( .A1(n5526), .A2(n5525), .ZN(n8905) );
  AND2_X1 U6037 ( .A1(n6383), .A2(n9315), .ZN(n4317) );
  AND2_X1 U6038 ( .A1(n4904), .A2(n8186), .ZN(n4318) );
  NAND2_X1 U6039 ( .A1(n9353), .A2(n4941), .ZN(n4944) );
  INV_X1 U6040 ( .A(n5889), .ZN(n4681) );
  AND2_X1 U6041 ( .A1(n6072), .A2(n6074), .ZN(n4319) );
  AND2_X1 U6042 ( .A1(n9570), .A2(n9408), .ZN(n4320) );
  INV_X1 U6043 ( .A(n4477), .ZN(n4476) );
  NAND2_X1 U6044 ( .A1(n4478), .A2(n5717), .ZN(n4477) );
  AND2_X1 U6045 ( .A1(n4878), .A2(n8180), .ZN(n4321) );
  AND2_X1 U6046 ( .A1(n4489), .A2(n4316), .ZN(n4322) );
  INV_X1 U6047 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n10062) );
  AND2_X1 U6048 ( .A1(n8225), .A2(n6412), .ZN(n9296) );
  NOR2_X1 U6049 ( .A1(n9599), .A2(n9458), .ZN(n4323) );
  AND2_X1 U6050 ( .A1(n6448), .A2(n8217), .ZN(n9390) );
  INV_X1 U6051 ( .A(n9390), .ZN(n4907) );
  NOR2_X1 U6052 ( .A1(n4942), .A2(n9362), .ZN(n4324) );
  NAND2_X1 U6053 ( .A1(n6718), .A2(n6717), .ZN(n4325) );
  OR2_X1 U6054 ( .A1(n4841), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n4326) );
  NAND2_X1 U6055 ( .A1(n4756), .A2(n4755), .ZN(n4327) );
  INV_X1 U6056 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7916) );
  AND2_X1 U6057 ( .A1(n9574), .A2(n6731), .ZN(n8214) );
  AND2_X1 U6058 ( .A1(n4574), .A2(n8205), .ZN(n4328) );
  NOR2_X1 U6059 ( .A1(n8923), .A2(n8690), .ZN(n4329) );
  NOR2_X1 U6060 ( .A1(n8695), .A2(n8405), .ZN(n4330) );
  NOR2_X1 U6061 ( .A1(n8911), .A2(n8450), .ZN(n4331) );
  OR2_X1 U6062 ( .A1(n6263), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4332) );
  NAND2_X1 U6063 ( .A1(n7578), .A2(n7500), .ZN(n4333) );
  AND2_X1 U6064 ( .A1(n5376), .A2(SI_18_), .ZN(n4334) );
  INV_X1 U6065 ( .A(n8898), .ZN(n4626) );
  AND2_X1 U6066 ( .A1(n6673), .A2(n6672), .ZN(n4335) );
  AND2_X1 U6067 ( .A1(n5731), .A2(n5735), .ZN(n8752) );
  INV_X1 U6068 ( .A(n8752), .ZN(n4469) );
  INV_X1 U6069 ( .A(n8289), .ZN(n7199) );
  INV_X1 U6070 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6979) );
  AND2_X1 U6071 ( .A1(n5770), .A2(n5771), .ZN(n8898) );
  INV_X1 U6072 ( .A(n5769), .ZN(n5771) );
  AND2_X1 U6073 ( .A1(n6140), .A2(n6138), .ZN(n4336) );
  NAND2_X1 U6074 ( .A1(n4316), .A2(n5772), .ZN(n4337) );
  NOR2_X1 U6075 ( .A1(n9543), .A2(n9316), .ZN(n4338) );
  OR2_X1 U6076 ( .A1(n4715), .A2(n4506), .ZN(n4339) );
  NAND2_X1 U6077 ( .A1(n5547), .A2(n5546), .ZN(n8900) );
  OR2_X1 U6078 ( .A1(n8958), .A2(n8415), .ZN(n5722) );
  OR2_X1 U6079 ( .A1(n5898), .A2(n8382), .ZN(n4340) );
  NAND2_X1 U6080 ( .A1(n5566), .A2(n5565), .ZN(n8611) );
  INV_X1 U6081 ( .A(n8611), .ZN(n4406) );
  NAND2_X1 U6082 ( .A1(n5435), .A2(n5434), .ZN(n8931) );
  NOR2_X1 U6083 ( .A1(n8899), .A2(n4852), .ZN(n4341) );
  AND2_X1 U6084 ( .A1(n4732), .A2(n5735), .ZN(n4342) );
  AND2_X1 U6085 ( .A1(n8265), .A2(n5771), .ZN(n4343) );
  AND2_X1 U6086 ( .A1(n7986), .A2(n8072), .ZN(n7774) );
  INV_X1 U6087 ( .A(n7774), .ZN(n4912) );
  AND2_X1 U6088 ( .A1(n6378), .A2(n8219), .ZN(n4344) );
  NAND2_X1 U6089 ( .A1(n8710), .A2(n4927), .ZN(n8675) );
  NOR2_X1 U6090 ( .A1(n9360), .A2(n8218), .ZN(n4345) );
  NAND2_X1 U6091 ( .A1(n5604), .A2(n7627), .ZN(n4346) );
  AND2_X1 U6092 ( .A1(n4729), .A2(n6406), .ZN(n4347) );
  AND2_X1 U6093 ( .A1(n5095), .A2(n5096), .ZN(n4348) );
  AND2_X1 U6094 ( .A1(n8611), .A2(n8268), .ZN(n5769) );
  AND2_X1 U6095 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4349) );
  NAND2_X1 U6096 ( .A1(n8346), .A2(n8347), .ZN(n4350) );
  NAND2_X1 U6097 ( .A1(n9106), .A2(n6706), .ZN(n4351) );
  OR2_X1 U6098 ( .A1(n9886), .A2(n8458), .ZN(n4352) );
  INV_X1 U6099 ( .A(n6109), .ZN(n6132) );
  INV_X1 U6100 ( .A(n7837), .ZN(n4454) );
  AND2_X1 U6101 ( .A1(n8872), .A2(n4277), .ZN(n4353) );
  NAND2_X1 U6102 ( .A1(n8872), .A2(n8880), .ZN(n8838) );
  OAI21_X1 U6103 ( .B1(n8849), .B2(n4532), .A(n4531), .ZN(n8806) );
  NAND2_X1 U6104 ( .A1(n6361), .A2(n6360), .ZN(n9543) );
  INV_X1 U6105 ( .A(n9543), .ZN(n4938) );
  OR2_X1 U6106 ( .A1(n9460), .A2(n9595), .ZN(n4354) );
  NAND2_X1 U6107 ( .A1(n4692), .A2(n4688), .ZN(n8001) );
  NAND2_X1 U6108 ( .A1(n4872), .A2(n8139), .ZN(n8175) );
  NAND2_X1 U6109 ( .A1(n7614), .A2(n7613), .ZN(n7802) );
  NAND2_X1 U6110 ( .A1(n5415), .A2(n5414), .ZN(n8936) );
  INV_X1 U6111 ( .A(n8936), .ZN(n4857) );
  NAND2_X1 U6112 ( .A1(n7604), .A2(n7603), .ZN(n7737) );
  OR2_X1 U6113 ( .A1(n8923), .A2(n8349), .ZN(n8654) );
  INV_X1 U6114 ( .A(n8654), .ZN(n4925) );
  INV_X1 U6115 ( .A(n4785), .ZN(n4784) );
  NOR2_X1 U6116 ( .A1(n4786), .A2(n5575), .ZN(n4785) );
  AND2_X1 U6117 ( .A1(n5519), .A2(n5495), .ZN(n5517) );
  AND2_X1 U6118 ( .A1(n5574), .A2(SI_29_), .ZN(n4355) );
  OR2_X1 U6119 ( .A1(n9460), .A2(n4936), .ZN(n4356) );
  INV_X2 U6120 ( .A(n9923), .ZN(n9926) );
  INV_X1 U6121 ( .A(n7780), .ZN(n4846) );
  INV_X1 U6122 ( .A(n9474), .ZN(n9510) );
  OR2_X1 U6123 ( .A1(n7142), .A2(n9669), .ZN(n9474) );
  OAI211_X1 U6124 ( .C1(n6124), .C2(n7403), .A(n6123), .B(n6122), .ZN(n7667)
         );
  INV_X2 U6125 ( .A(n9912), .ZN(n9913) );
  INV_X1 U6126 ( .A(n8282), .ZN(n7120) );
  INV_X4 U6127 ( .A(n9733), .ZN(n9735) );
  NAND2_X1 U6128 ( .A1(n7618), .A2(n9728), .ZN(n9733) );
  NAND2_X1 U6129 ( .A1(n6310), .A2(n6309), .ZN(n9580) );
  INV_X1 U6130 ( .A(n9580), .ZN(n4934) );
  NAND2_X1 U6131 ( .A1(n6231), .A2(n6230), .ZN(n9610) );
  INV_X1 U6132 ( .A(n9610), .ZN(n4948) );
  INV_X1 U6133 ( .A(n8968), .ZN(n4860) );
  NAND2_X1 U6134 ( .A1(n5345), .A2(n5344), .ZN(n8958) );
  INV_X1 U6135 ( .A(n8958), .ZN(n4419) );
  INV_X1 U6136 ( .A(n7791), .ZN(n4403) );
  INV_X1 U6137 ( .A(n8987), .ZN(n4421) );
  INV_X1 U6138 ( .A(n7648), .ZN(n4929) );
  INV_X1 U6139 ( .A(n9186), .ZN(n9165) );
  OAI21_X1 U6140 ( .B1(n7328), .B2(n7117), .A(n8018), .ZN(n5618) );
  AND2_X1 U6141 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n4357) );
  NAND2_X1 U6142 ( .A1(n7102), .A2(n7112), .ZN(n7326) );
  INV_X1 U6143 ( .A(n4669), .ZN(n7118) );
  NAND2_X1 U6144 ( .A1(n5781), .A2(n7627), .ZN(n4669) );
  OR2_X1 U6145 ( .A1(n7001), .A2(n4643), .ZN(n4358) );
  AND2_X1 U6146 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4359) );
  INV_X1 U6147 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4363) );
  NAND2_X1 U6148 ( .A1(n9362), .A2(n9506), .ZN(n4447) );
  NAND2_X1 U6149 ( .A1(n9348), .A2(n9506), .ZN(n9317) );
  AOI222_X1 U6150 ( .A1(n9348), .A2(n9510), .B1(n9509), .B2(n9347), .C1(n9377), 
        .C2(n9506), .ZN(n9557) );
  MUX2_X1 U6151 ( .A(n5744), .B(n5743), .S(n5776), .Z(n5749) );
  NAND4_X1 U6152 ( .A1(n4952), .A2(n5964), .A3(n6052), .A4(n6510), .ZN(n5975)
         );
  AND2_X2 U6153 ( .A1(n5966), .A2(n4951), .ZN(n4952) );
  INV_X1 U6154 ( .A(n9781), .ZN(n7602) );
  NAND2_X1 U6155 ( .A1(n9366), .A2(n8188), .ZN(n8190) );
  NAND2_X1 U6156 ( .A1(n8135), .A2(n8134), .ZN(n8138) );
  NAND4_X2 U6157 ( .A1(n4980), .A2(n4979), .A3(n5625), .A4(n5626), .ZN(n5633)
         );
  AOI21_X2 U6158 ( .B1(n8065), .B2(n8066), .A(n5858), .ZN(n8312) );
  NAND2_X1 U6159 ( .A1(n8182), .A2(n8181), .ZN(n9412) );
  NAND2_X1 U6160 ( .A1(n7607), .A2(n7801), .ZN(n7793) );
  NAND2_X1 U6161 ( .A1(n6465), .A2(n6422), .ZN(n6107) );
  NAND2_X1 U6162 ( .A1(n9417), .A2(n9418), .ZN(n8213) );
  AND3_X2 U6163 ( .A1(n6090), .A2(n6092), .A3(n6091), .ZN(n6093) );
  INV_X2 U6164 ( .A(n6124), .ZN(n7276) );
  NAND2_X2 U6165 ( .A1(n6524), .A2(n8231), .ZN(n6124) );
  NAND2_X1 U6166 ( .A1(n5356), .A2(n5355), .ZN(n5360) );
  NAND2_X1 U6167 ( .A1(n4760), .A2(n4758), .ZN(n5466) );
  INV_X1 U6168 ( .A(n4807), .ZN(n4806) );
  NAND2_X1 U6169 ( .A1(n5340), .A2(n5339), .ZN(n5354) );
  NAND2_X1 U6170 ( .A1(n4770), .A2(n4768), .ZN(n5411) );
  NAND2_X1 U6171 ( .A1(n5539), .A2(n5538), .ZN(n8628) );
  NAND2_X1 U6172 ( .A1(n5071), .A2(n5072), .ZN(n5075) );
  AND2_X1 U6173 ( .A1(n6073), .A2(n6075), .ZN(n4498) );
  NAND2_X1 U6174 ( .A1(n9935), .A2(n9936), .ZN(n9934) );
  NAND2_X1 U6175 ( .A1(n9948), .A2(n4430), .ZN(n9947) );
  NOR2_X1 U6176 ( .A1(n9952), .A2(n9951), .ZN(n9950) );
  NAND2_X1 U6177 ( .A1(n9934), .A2(n4428), .ZN(n9932) );
  NAND2_X1 U6178 ( .A1(n4427), .A2(n9693), .ZN(n9694) );
  NAND2_X1 U6179 ( .A1(n4426), .A2(n9691), .ZN(n9692) );
  OAI21_X1 U6180 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9937), .ZN(n9935) );
  OAI21_X1 U6181 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9940), .ZN(n9938) );
  OAI21_X1 U6182 ( .B1(n9927), .B2(n9683), .A(n9929), .ZN(n10131) );
  NOR2_X1 U6183 ( .A1(n9953), .A2(n4357), .ZN(n9952) );
  OAI21_X1 U6184 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9701), .A(n10120), .ZN(
        n9704) );
  NAND2_X1 U6185 ( .A1(n9503), .A2(n9504), .ZN(n8145) );
  NAND2_X1 U6186 ( .A1(n4370), .A2(n4559), .ZN(n5073) );
  NAND2_X1 U6187 ( .A1(n8211), .A2(n8210), .ZN(n9417) );
  NAND2_X1 U6188 ( .A1(n4458), .A2(n4352), .ZN(n8089) );
  NAND3_X1 U6189 ( .A1(n5021), .A2(n5022), .A3(n5023), .ZN(n4372) );
  NAND2_X1 U6190 ( .A1(n9001), .A2(n9913), .ZN(n4377) );
  NAND2_X1 U6191 ( .A1(n8924), .A2(n4378), .ZN(n9001) );
  INV_X1 U6192 ( .A(n8294), .ZN(n4380) );
  NAND2_X1 U6193 ( .A1(n5053), .A2(n5054), .ZN(n5058) );
  NAND2_X1 U6194 ( .A1(n5035), .A2(n5036), .ZN(n5053) );
  NAND2_X1 U6195 ( .A1(n5102), .A2(n5101), .ZN(n5119) );
  NAND2_X1 U6196 ( .A1(n4381), .A2(n5083), .ZN(n5099) );
  NAND2_X1 U6197 ( .A1(n4557), .A2(n5081), .ZN(n4381) );
  OR2_X1 U6198 ( .A1(n9234), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4383) );
  NAND2_X1 U6199 ( .A1(n6102), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6103) );
  NAND4_X1 U6200 ( .A1(n4389), .A2(n4979), .A3(n5625), .A4(n4980), .ZN(n4998)
         );
  NAND3_X1 U6201 ( .A1(n4391), .A2(n4642), .A3(n4390), .ZN(P2_U3244) );
  NAND3_X1 U6202 ( .A1(n5808), .A2(n5807), .A3(n8018), .ZN(n4391) );
  NAND2_X1 U6203 ( .A1(n4520), .A2(n4613), .ZN(n4519) );
  OAI21_X1 U6204 ( .B1(n6262), .B2(n6479), .A(n6480), .ZN(n6242) );
  AOI21_X1 U6205 ( .B1(n6370), .B2(n9387), .A(n6346), .ZN(n4521) );
  NAND2_X2 U6206 ( .A1(n7266), .A2(n6081), .ZN(n7137) );
  NAND2_X1 U6207 ( .A1(n4717), .A2(n8219), .ZN(n9345) );
  NAND2_X1 U6208 ( .A1(n4401), .A2(n9539), .ZN(n9637) );
  OAI21_X1 U6209 ( .B1(n9540), .B2(n9624), .A(n9538), .ZN(n4402) );
  NAND2_X1 U6210 ( .A1(n4775), .A2(n5138), .ZN(n5161) );
  NAND2_X1 U6211 ( .A1(n4999), .A2(n4998), .ZN(n7004) );
  NAND2_X1 U6212 ( .A1(n8277), .A2(n8279), .ZN(n8278) );
  NAND2_X1 U6213 ( .A1(n9535), .A2(n9528), .ZN(n4445) );
  NAND2_X1 U6214 ( .A1(n4405), .A2(n8809), .ZN(n5720) );
  NAND2_X1 U6215 ( .A1(n5716), .A2(n5715), .ZN(n4405) );
  NAND2_X1 U6216 ( .A1(n5209), .A2(n5206), .ZN(n5183) );
  NAND2_X1 U6217 ( .A1(n5136), .A2(n5135), .ZN(n4775) );
  NOR2_X1 U6218 ( .A1(n4538), .A2(n8603), .ZN(n4537) );
  NAND2_X1 U6219 ( .A1(n5734), .A2(n4631), .ZN(n4630) );
  NAND2_X1 U6220 ( .A1(n4630), .A2(n5735), .ZN(n5728) );
  INV_X1 U6221 ( .A(n4851), .ZN(n4540) );
  NAND2_X2 U6222 ( .A1(n5004), .A2(n5003), .ZN(n7020) );
  MUX2_X1 U6223 ( .A(n8582), .B(n8581), .S(n8758), .Z(n8584) );
  OR2_X2 U6224 ( .A1(n5633), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U6225 ( .A1(n7176), .A2(n7177), .ZN(n7175) );
  NAND2_X1 U6226 ( .A1(n7294), .A2(n7295), .ZN(n7293) );
  INV_X1 U6227 ( .A(n7552), .ZN(n4434) );
  NAND2_X1 U6228 ( .A1(n4660), .A2(n9278), .ZN(n4659) );
  NAND2_X1 U6229 ( .A1(n7247), .A2(n7246), .ZN(n7245) );
  XNOR2_X2 U6230 ( .A(n6893), .B(n7021), .ZN(n9232) );
  AND2_X2 U6231 ( .A1(n4645), .A2(n4644), .ZN(n6893) );
  NOR2_X1 U6232 ( .A1(n7420), .A2(n7419), .ZN(n7418) );
  NOR2_X1 U6233 ( .A1(n7386), .A2(n7385), .ZN(n7384) );
  NAND2_X1 U6234 ( .A1(n4703), .A2(n4706), .ZN(n9503) );
  NAND2_X1 U6235 ( .A1(n9331), .A2(n8221), .ZN(n9313) );
  NAND2_X1 U6236 ( .A1(n4717), .A2(n4344), .ZN(n9331) );
  NAND2_X1 U6237 ( .A1(n9388), .A2(n8216), .ZN(n9389) );
  OR2_X1 U6238 ( .A1(n6860), .A2(n6815), .ZN(n6838) );
  INV_X4 U6239 ( .A(n6603), .ZN(n6606) );
  NAND3_X1 U6240 ( .A1(n4832), .A2(n6610), .A3(n4596), .ZN(n7671) );
  INV_X1 U6241 ( .A(n4694), .ZN(n4693) );
  XNOR2_X2 U6242 ( .A(n5230), .B(n5225), .ZN(n6978) );
  XNOR2_X1 U6243 ( .A(n5038), .B(n5037), .ZN(n6956) );
  NAND2_X1 U6244 ( .A1(n8567), .A2(n8568), .ZN(n8569) );
  NAND2_X1 U6245 ( .A1(n5103), .A2(n6982), .ZN(n4418) );
  INV_X1 U6246 ( .A(n4564), .ZN(n4563) );
  INV_X1 U6247 ( .A(n5228), .ZN(n4565) );
  NAND2_X1 U6248 ( .A1(n4799), .A2(n4803), .ZN(n5340) );
  NAND2_X1 U6249 ( .A1(n4470), .A2(n4468), .ZN(n4921) );
  NAND2_X1 U6250 ( .A1(n4562), .A2(n4560), .ZN(n5257) );
  NOR2_X2 U6251 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5001) );
  NOR2_X1 U6252 ( .A1(n7841), .A2(n4425), .ZN(n7846) );
  NAND2_X1 U6253 ( .A1(n7846), .A2(n7845), .ZN(n7926) );
  AOI21_X1 U6254 ( .B1(n7163), .B2(n7161), .A(n7162), .ZN(n7214) );
  NOR2_X4 U6255 ( .A1(n4967), .A2(n8952), .ZN(n8770) );
  NOR2_X4 U6256 ( .A1(n8113), .A2(n8982), .ZN(n8872) );
  NAND2_X1 U6257 ( .A1(n4540), .A2(n4539), .ZN(n4538) );
  NAND2_X1 U6258 ( .A1(n5886), .A2(n4676), .ZN(n4672) );
  OAI21_X1 U6259 ( .B1(n8895), .B2(n9907), .A(n4341), .ZN(n4851) );
  NAND2_X1 U6260 ( .A1(n8894), .A2(n4850), .ZN(n8996) );
  NAND2_X1 U6261 ( .A1(n8996), .A2(n9913), .ZN(n4910) );
  NAND2_X1 U6262 ( .A1(n7960), .A2(n7959), .ZN(n7962) );
  NAND2_X1 U6263 ( .A1(n4891), .A2(n4893), .ZN(n7960) );
  AOI21_X2 U6264 ( .B1(n9324), .B2(n9333), .A(n8194), .ZN(n9306) );
  OAI21_X1 U6265 ( .B1(n4871), .B2(n4867), .A(n4866), .ZN(n8177) );
  AOI21_X1 U6266 ( .B1(n5633), .B2(n4349), .A(n4290), .ZN(n4999) );
  NAND2_X2 U6267 ( .A1(n6124), .A2(n4257), .ZN(n6101) );
  NAND2_X1 U6268 ( .A1(n7928), .A2(n7929), .ZN(n8567) );
  NAND2_X1 U6269 ( .A1(n7020), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4423) );
  AND2_X2 U6270 ( .A1(n8327), .A2(n5884), .ZN(n5886) );
  NAND2_X1 U6271 ( .A1(n4450), .A2(n5907), .ZN(n8422) );
  NAND2_X1 U6272 ( .A1(n10116), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U6273 ( .A1(n10130), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n4427) );
  NOR2_X1 U6274 ( .A1(n10126), .A2(n10125), .ZN(n10124) );
  NOR2_X1 U6275 ( .A1(n9945), .A2(n9944), .ZN(n9943) );
  NOR2_X1 U6276 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10117), .ZN(n9689) );
  NOR2_X1 U6277 ( .A1(n8381), .A2(n5901), .ZN(n5902) );
  NOR2_X2 U6278 ( .A1(n9265), .A2(n4436), .ZN(n9706) );
  OAI21_X1 U6279 ( .B1(n9276), .B2(n9275), .A(n4661), .ZN(n4660) );
  XNOR2_X1 U6280 ( .A(n9268), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9276) );
  OAI211_X1 U6281 ( .C1(n9279), .C2(n9278), .A(n4662), .B(n4659), .ZN(P1_U3260) );
  NOR2_X1 U6282 ( .A1(n9213), .A2(n4307), .ZN(n7247) );
  NOR2_X1 U6283 ( .A1(n7428), .A2(n4655), .ZN(n7420) );
  NAND2_X1 U6284 ( .A1(n5305), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5333) );
  INV_X1 U6285 ( .A(n4628), .ZN(n4627) );
  NOR2_X2 U6286 ( .A1(n5455), .A2(n8321), .ZN(n4440) );
  NOR2_X2 U6287 ( .A1(n5386), .A2(n5385), .ZN(n4441) );
  NAND2_X1 U6288 ( .A1(n6107), .A2(n4729), .ZN(n7654) );
  NAND2_X1 U6289 ( .A1(n6094), .A2(n6539), .ZN(n6465) );
  NAND2_X1 U6290 ( .A1(n7614), .A2(n4314), .ZN(n4714) );
  NAND2_X1 U6291 ( .A1(n7654), .A2(n7650), .ZN(n7610) );
  NAND2_X1 U6292 ( .A1(n9529), .A2(n4444), .ZN(n9636) );
  INV_X2 U6293 ( .A(n6101), .ZN(n6386) );
  INV_X1 U6294 ( .A(n8421), .ZN(n4450) );
  NAND2_X1 U6295 ( .A1(n4670), .A2(n4671), .ZN(n8421) );
  INV_X1 U6296 ( .A(n7914), .ZN(n4695) );
  NAND2_X1 U6297 ( .A1(n5870), .A2(n5869), .ZN(n8363) );
  NAND2_X1 U6298 ( .A1(n4686), .A2(n4687), .ZN(n8065) );
  XNOR2_X2 U6299 ( .A(n4453), .B(n4959), .ZN(n6971) );
  OR2_X2 U6300 ( .A1(n8320), .A2(n4340), .ZN(n5904) );
  NAND2_X1 U6301 ( .A1(n4775), .A2(n4774), .ZN(n5209) );
  NOR2_X2 U6302 ( .A1(n8704), .A2(n8926), .ZN(n8260) );
  NAND2_X1 U6303 ( .A1(n8079), .A2(n9906), .ZN(n8024) );
  NOR2_X4 U6304 ( .A1(n8692), .A2(n8923), .ZN(n8682) );
  NAND2_X1 U6305 ( .A1(n4910), .A2(n4908), .ZN(P2_U3517) );
  XNOR2_X2 U6306 ( .A(n5039), .B(P2_IR_REG_2__SCAN_IN), .ZN(n7039) );
  NAND3_X2 U6307 ( .A1(n9702), .A2(n4457), .A3(n4456), .ZN(n4754) );
  INV_X2 U6308 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4457) );
  INV_X1 U6309 ( .A(n7504), .ZN(n4460) );
  NAND2_X1 U6310 ( .A1(n7982), .A2(n4305), .ZN(n4465) );
  OAI21_X1 U6311 ( .B1(n5337), .B2(n4473), .A(n4471), .ZN(n8751) );
  NAND2_X1 U6312 ( .A1(n5337), .A2(n4471), .ZN(n4470) );
  NAND2_X1 U6313 ( .A1(n5337), .A2(n5717), .ZN(n8783) );
  INV_X1 U6314 ( .A(n8246), .ZN(n4478) );
  NAND2_X1 U6315 ( .A1(n5605), .A2(n4481), .ZN(n4479) );
  NAND2_X1 U6316 ( .A1(n8264), .A2(n4343), .ZN(n4488) );
  NAND2_X1 U6317 ( .A1(n4488), .A2(n4489), .ZN(n5588) );
  NAND2_X1 U6318 ( .A1(n8264), .A2(n8265), .ZN(n8267) );
  NAND2_X1 U6319 ( .A1(n8725), .A2(n4497), .ZN(n8710) );
  NAND2_X1 U6320 ( .A1(n7268), .A2(n7267), .ZN(n7266) );
  NAND2_X2 U6321 ( .A1(n4498), .A2(n4319), .ZN(n9201) );
  INV_X1 U6322 ( .A(n7734), .ZN(n4508) );
  NAND4_X1 U6323 ( .A1(n4512), .A2(n4899), .A3(n6510), .A4(n5964), .ZN(n5978)
         );
  NOR2_X2 U6324 ( .A1(n6509), .A2(n5960), .ZN(n5964) );
  NAND3_X1 U6325 ( .A1(n6384), .A2(n4522), .A3(n4519), .ZN(n6404) );
  NAND2_X1 U6326 ( .A1(n7222), .A2(n7201), .ZN(n4524) );
  NAND2_X1 U6327 ( .A1(n4525), .A2(n7200), .ZN(n7222) );
  NAND2_X1 U6328 ( .A1(n8849), .A2(n4531), .ZN(n4527) );
  NAND3_X1 U6329 ( .A1(n4527), .A2(n4526), .A3(n4291), .ZN(n8791) );
  NOR2_X1 U6330 ( .A1(n8825), .A2(n8242), .ZN(n4534) );
  NOR2_X1 U6331 ( .A1(n8242), .A2(n8243), .ZN(n4529) );
  AND2_X2 U6332 ( .A1(n4744), .A2(n4743), .ZN(n8893) );
  NAND2_X1 U6333 ( .A1(n8255), .A2(n4283), .ZN(n4542) );
  OAI22_X2 U6334 ( .A1(n8667), .A2(n4548), .B1(n4549), .B2(n4552), .ZN(n8618)
         );
  INV_X1 U6335 ( .A(n8258), .ZN(n4552) );
  OAI211_X1 U6336 ( .C1(n7768), .C2(n4554), .A(n7992), .B(n4553), .ZN(n7994)
         );
  NAND2_X1 U6337 ( .A1(n7768), .A2(n7767), .ZN(n7989) );
  INV_X1 U6338 ( .A(n7988), .ZN(n4554) );
  INV_X2 U6339 ( .A(n4629), .ZN(n5583) );
  AND4_X2 U6340 ( .A1(n4993), .A2(n4991), .A3(n4992), .A4(n4556), .ZN(n5812)
         );
  AND2_X2 U6341 ( .A1(n9023), .A2(n4987), .ZN(n4629) );
  XNOR2_X1 U6342 ( .A(n4557), .B(n5080), .ZN(n6941) );
  NAND2_X1 U6343 ( .A1(n5213), .A2(n4563), .ZN(n4562) );
  NAND2_X1 U6344 ( .A1(n5213), .A2(n5212), .ZN(n5230) );
  NAND2_X1 U6345 ( .A1(n5122), .A2(n5121), .ZN(n5136) );
  NAND3_X1 U6346 ( .A1(n4570), .A2(n4569), .A3(n5208), .ZN(n5211) );
  NAND2_X1 U6347 ( .A1(n5134), .A2(n4774), .ZN(n4569) );
  NAND3_X1 U6348 ( .A1(n5122), .A2(n4774), .A3(n5121), .ZN(n4570) );
  NAND2_X1 U6349 ( .A1(n9160), .A2(n4581), .ZN(n4577) );
  NAND2_X1 U6350 ( .A1(n4577), .A2(n4576), .ZN(P1_U3212) );
  NAND3_X1 U6351 ( .A1(n5965), .A2(n5966), .A3(n6052), .ZN(n6228) );
  AND4_X2 U6352 ( .A1(n5965), .A2(n5966), .A3(n6052), .A4(n5956), .ZN(n6219)
         );
  INV_X1 U6353 ( .A(n9042), .ZN(n4589) );
  NAND2_X1 U6354 ( .A1(n6715), .A2(n4351), .ZN(n4583) );
  OR2_X1 U6355 ( .A1(n6715), .A2(n4819), .ZN(n4585) );
  NAND2_X1 U6356 ( .A1(n9045), .A2(n6715), .ZN(n4588) );
  OR2_X1 U6357 ( .A1(n4587), .A2(n4819), .ZN(n4586) );
  OAI21_X2 U6358 ( .B1(n7872), .B2(n4593), .A(n4591), .ZN(n8124) );
  NOR2_X1 U6359 ( .A1(n8124), .A2(n8125), .ZN(n6678) );
  NAND2_X1 U6360 ( .A1(n7671), .A2(n6619), .ZN(n7857) );
  CLKBUF_X1 U6361 ( .A(n6605), .Z(n4597) );
  NOR2_X2 U6362 ( .A1(n9081), .A2(n9080), .ZN(n9163) );
  NOR2_X2 U6363 ( .A1(n9120), .A2(n6773), .ZN(n9081) );
  AOI21_X2 U6364 ( .B1(n4830), .B2(n4828), .A(n4825), .ZN(n9120) );
  NAND2_X2 U6365 ( .A1(n4831), .A2(n9138), .ZN(n4830) );
  NAND2_X1 U6366 ( .A1(n4600), .A2(n6531), .ZN(n6532) );
  NAND3_X1 U6367 ( .A1(n4603), .A2(n4602), .A3(n4601), .ZN(n4600) );
  NAND3_X1 U6368 ( .A1(n6202), .A2(n6418), .A3(n8143), .ZN(n4611) );
  NAND2_X1 U6369 ( .A1(n6107), .A2(n4347), .ZN(n6127) );
  NAND2_X1 U6370 ( .A1(n4615), .A2(n4616), .ZN(n5780) );
  NAND2_X1 U6371 ( .A1(n5767), .A2(n4618), .ZN(n4615) );
  NOR2_X1 U6372 ( .A1(n5765), .A2(n5766), .ZN(n4628) );
  NAND4_X1 U6373 ( .A1(n4634), .A2(n4979), .A3(n5625), .A4(n4980), .ZN(n4985)
         );
  OAI21_X1 U6374 ( .B1(n4640), .B2(n4639), .A(n4636), .ZN(n5685) );
  OAI21_X1 U6375 ( .B1(n5677), .B2(n5776), .A(n5791), .ZN(n4641) );
  NAND3_X1 U6376 ( .A1(n5093), .A2(n5094), .A3(n4348), .ZN(n8461) );
  NAND3_X1 U6377 ( .A1(n6086), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n4651) );
  OAI21_X1 U6378 ( .B1(n9240), .B2(n4657), .A(n4656), .ZN(n9252) );
  NAND2_X1 U6379 ( .A1(n4666), .A2(n4664), .ZN(n8327) );
  NAND2_X2 U6380 ( .A1(n5810), .A2(n4667), .ZN(n5828) );
  INV_X1 U6381 ( .A(n7870), .ZN(n5809) );
  NAND3_X1 U6382 ( .A1(n5904), .A2(n4350), .A3(n5903), .ZN(n4670) );
  NAND2_X1 U6383 ( .A1(n5904), .A2(n5903), .ZN(n8345) );
  NAND2_X1 U6384 ( .A1(n4672), .A2(n4673), .ZN(n5900) );
  NAND2_X1 U6385 ( .A1(n4683), .A2(n4306), .ZN(n4682) );
  NAND2_X1 U6386 ( .A1(n7560), .A2(n5839), .ZN(n4683) );
  NOR2_X1 U6387 ( .A1(n7565), .A2(n5840), .ZN(n7559) );
  NAND2_X1 U6388 ( .A1(n7830), .A2(n4689), .ZN(n4687) );
  AOI21_X2 U6389 ( .B1(n4693), .B2(n5851), .A(n4286), .ZN(n4692) );
  NOR2_X1 U6390 ( .A1(n5323), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5365) );
  NAND4_X1 U6391 ( .A1(n5364), .A2(n4700), .A3(n5627), .A4(n4696), .ZN(n5611)
         );
  NOR2_X1 U6392 ( .A1(n5323), .A2(n4697), .ZN(n4696) );
  CLKBUF_X1 U6393 ( .A(n5365), .Z(n4698) );
  NAND4_X1 U6394 ( .A1(n5366), .A2(n5365), .A3(n5364), .A4(n4701), .ZN(n4699)
         );
  XNOR2_X1 U6395 ( .A(n5824), .B(n5825), .ZN(n8279) );
  NAND2_X1 U6396 ( .A1(n7967), .A2(n4704), .ZN(n4703) );
  INV_X1 U6397 ( .A(n7801), .ZN(n4716) );
  INV_X1 U6398 ( .A(n7800), .ZN(n4715) );
  NAND2_X1 U6399 ( .A1(n8208), .A2(n4718), .ZN(n9433) );
  NAND2_X1 U6400 ( .A1(n9433), .A2(n8209), .ZN(n8211) );
  NAND2_X1 U6401 ( .A1(n8213), .A2(n4724), .ZN(n9388) );
  AND2_X2 U6402 ( .A1(n4728), .A2(n6069), .ZN(n4726) );
  NAND2_X2 U6403 ( .A1(n8669), .A2(n8668), .ZN(n8667) );
  NAND3_X1 U6404 ( .A1(n4739), .A2(n4333), .A3(n7468), .ZN(n4738) );
  NOR2_X2 U6405 ( .A1(n8893), .A2(n4742), .ZN(n8904) );
  OR2_X2 U6406 ( .A1(n8618), .A2(n4745), .ZN(n4744) );
  NAND2_X1 U6407 ( .A1(n8255), .A2(n8254), .ZN(n8703) );
  INV_X1 U6408 ( .A(n8254), .ZN(n4751) );
  NAND2_X4 U6409 ( .A1(n4754), .A2(n4752), .ZN(n5231) );
  NAND3_X1 U6410 ( .A1(n4753), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U6411 ( .A1(n5805), .A2(n5776), .ZN(n4756) );
  NAND2_X1 U6412 ( .A1(n5804), .A2(n5778), .ZN(n4755) );
  NAND2_X1 U6413 ( .A1(n5413), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U6414 ( .A1(n5413), .A2(n5412), .ZN(n5428) );
  NAND2_X1 U6415 ( .A1(n5360), .A2(n4767), .ZN(n4770) );
  NAND2_X1 U6416 ( .A1(n5360), .A2(n5359), .ZN(n5375) );
  NAND3_X1 U6417 ( .A1(n4772), .A2(n5373), .A3(n4771), .ZN(n4769) );
  NAND2_X1 U6418 ( .A1(n5557), .A2(n4780), .ZN(n4779) );
  NAND2_X1 U6419 ( .A1(n5557), .A2(n5556), .ZN(n4787) );
  NAND2_X1 U6420 ( .A1(n5484), .A2(n4791), .ZN(n4790) );
  NAND3_X1 U6421 ( .A1(n5517), .A2(n4792), .A3(n5483), .ZN(n4789) );
  OR2_X1 U6422 ( .A1(n5484), .A2(n5483), .ZN(n4798) );
  NAND2_X1 U6423 ( .A1(n5257), .A2(n5256), .ZN(n5292) );
  NAND2_X1 U6424 ( .A1(n5257), .A2(n4800), .ZN(n4799) );
  NAND2_X1 U6425 ( .A1(n4811), .A2(n6594), .ZN(n7354) );
  OAI21_X1 U6426 ( .B1(n7304), .B2(n7303), .A(n4811), .ZN(n7407) );
  NAND2_X1 U6427 ( .A1(n7304), .A2(n7303), .ZN(n4811) );
  AND3_X2 U6428 ( .A1(n4814), .A2(n4813), .A3(n4812), .ZN(n6052) );
  NAND2_X1 U6429 ( .A1(n9137), .A2(n9140), .ZN(n4831) );
  NAND2_X1 U6430 ( .A1(n6757), .A2(n6756), .ZN(n9138) );
  NAND2_X1 U6431 ( .A1(n7309), .A2(n7308), .ZN(n4832) );
  OAI21_X1 U6432 ( .B1(n9081), .B2(n4834), .A(n4833), .ZN(n6860) );
  INV_X1 U6433 ( .A(n9080), .ZN(n4835) );
  NAND2_X1 U6434 ( .A1(n6219), .A2(n5950), .ZN(n6263) );
  NAND2_X1 U6435 ( .A1(n6219), .A2(n4839), .ZN(n4838) );
  NAND2_X1 U6436 ( .A1(n7223), .A2(n9853), .ZN(n4844) );
  NAND2_X1 U6437 ( .A1(n5823), .A2(n4844), .ZN(n7372) );
  NAND2_X1 U6438 ( .A1(n7224), .A2(n4844), .ZN(n9854) );
  INV_X1 U6439 ( .A(n8894), .ZN(n4848) );
  AOI21_X1 U6440 ( .B1(n4848), .B2(n9926), .A(n4293), .ZN(n4849) );
  OAI21_X1 U6441 ( .B1(n4850), .B2(n9923), .A(n4849), .ZN(P2_U3549) );
  AND2_X2 U6442 ( .A1(n8682), .A2(n4853), .ZN(n8605) );
  NAND2_X1 U6443 ( .A1(n8770), .A2(n4289), .ZN(n4859) );
  OR2_X2 U6444 ( .A1(n4859), .A2(n8931), .ZN(n8704) );
  INV_X1 U6445 ( .A(n4859), .ZN(n8722) );
  NAND3_X1 U6446 ( .A1(n8872), .A2(n4277), .A3(n8804), .ZN(n8787) );
  NAND2_X1 U6447 ( .A1(n7604), .A2(n4862), .ZN(n7739) );
  NAND3_X1 U6448 ( .A1(n7538), .A2(n7537), .A3(n7540), .ZN(n7604) );
  AOI21_X2 U6449 ( .B1(n8197), .B2(n4864), .A(n4338), .ZN(n8294) );
  NAND2_X1 U6450 ( .A1(n8294), .A2(n8302), .ZN(n9534) );
  NAND2_X1 U6451 ( .A1(n9468), .A2(n4879), .ZN(n4877) );
  NAND2_X1 U6452 ( .A1(n8190), .A2(n4883), .ZN(n4882) );
  NAND2_X1 U6453 ( .A1(n4882), .A2(n4885), .ZN(n9324) );
  NAND2_X1 U6454 ( .A1(n7795), .A2(n4892), .ZN(n4891) );
  INV_X1 U6455 ( .A(n4894), .ZN(n4893) );
  OAI22_X1 U6456 ( .A1(n7794), .A2(n4895), .B1(n9193), .B2(n9625), .ZN(n4894)
         );
  OAI21_X2 U6457 ( .B1(n8185), .B2(n4900), .A(n4901), .ZN(n9366) );
  NAND2_X1 U6458 ( .A1(n5664), .A2(n7363), .ZN(n7201) );
  OAI211_X2 U6459 ( .C1(n5059), .C2(n6956), .A(n5040), .B(n5041), .ZN(n7322)
         );
  NAND2_X1 U6460 ( .A1(n8604), .A2(n8871), .ZN(n4911) );
  OR2_X1 U6461 ( .A1(n9913), .A2(n4909), .ZN(n4908) );
  NAND2_X1 U6462 ( .A1(n4921), .A2(n4342), .ZN(n8734) );
  NAND2_X1 U6463 ( .A1(n5315), .A2(n5314), .ZN(n4922) );
  AOI21_X1 U6464 ( .B1(n5478), .B2(n4926), .A(n4925), .ZN(n4923) );
  INV_X1 U6465 ( .A(n5478), .ZN(n4924) );
  NOR2_X2 U6466 ( .A1(n4932), .A2(n9460), .ZN(n9413) );
  INV_X1 U6467 ( .A(n4944), .ZN(n9325) );
  CLKBUF_X1 U6468 ( .A(n8311), .Z(n8354) );
  CLKBUF_X1 U6469 ( .A(n7317), .Z(n8284) );
  INV_X1 U6470 ( .A(n7317), .ZN(n5815) );
  INV_X1 U6471 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5620) );
  AND2_X2 U6472 ( .A1(n6089), .A2(n6102), .ZN(n9205) );
  NAND2_X1 U6473 ( .A1(n5946), .A2(n5945), .ZN(P2_U3216) );
  CLKBUF_X1 U6474 ( .A(n6465), .Z(n7441) );
  OAI211_X1 U6475 ( .C1(n6794), .C2(n7701), .A(n6590), .B(n6589), .ZN(n7303)
         );
  AOI21_X1 U6476 ( .B1(n6614), .B2(n9201), .A(n6593), .ZN(n7304) );
  CLKBUF_X1 U6477 ( .A(n7610), .Z(n7541) );
  INV_X1 U6478 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5146) );
  AND2_X2 U6479 ( .A1(n7479), .A2(n7500), .ZN(n7508) );
  INV_X1 U6480 ( .A(n5196), .ZN(n5172) );
  XNOR2_X1 U6481 ( .A(n5518), .B(n5517), .ZN(n9032) );
  CLKBUF_X1 U6482 ( .A(n9503), .Z(n9505) );
  INV_X1 U6483 ( .A(n9160), .ZN(n9166) );
  AND2_X1 U6484 ( .A1(n7818), .A2(n7796), .ZN(n7943) );
  INV_X1 U6485 ( .A(n7201), .ZN(n7227) );
  XNOR2_X1 U6486 ( .A(n5504), .B(n5503), .ZN(n8158) );
  XNOR2_X1 U6487 ( .A(n8598), .B(n8898), .ZN(n8604) );
  XNOR2_X1 U6488 ( .A(n6411), .B(n5959), .ZN(n6506) );
  NAND2_X1 U6489 ( .A1(n5588), .A2(n8593), .ZN(n5589) );
  NAND2_X1 U6490 ( .A1(n9020), .A2(n9023), .ZN(n5088) );
  NAND2_X1 U6491 ( .A1(n9020), .A2(n4989), .ZN(n5065) );
  AND2_X1 U6492 ( .A1(n5606), .A2(n5610), .ZN(n4950) );
  AND2_X1 U6493 ( .A1(n6521), .A2(n5965), .ZN(n4951) );
  AND2_X1 U6494 ( .A1(n4275), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n4953) );
  AND2_X1 U6495 ( .A1(n7143), .A2(n9669), .ZN(n9506) );
  OR2_X1 U6496 ( .A1(n4938), .A2(n9173), .ZN(n4955) );
  AND2_X1 U6497 ( .A1(n5256), .A2(n5255), .ZN(n4957) );
  NAND2_X1 U6498 ( .A1(n4997), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4958) );
  INV_X1 U6499 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5050) );
  AND2_X1 U6500 ( .A1(n5212), .A2(n5189), .ZN(n4959) );
  NAND2_X1 U6501 ( .A1(n8804), .A2(n8818), .ZN(n5718) );
  AND2_X1 U6502 ( .A1(n5339), .A2(n5322), .ZN(n4960) );
  NAND2_X1 U6503 ( .A1(n9015), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4961) );
  OR2_X1 U6504 ( .A1(n6071), .A2(n6065), .ZN(n4962) );
  NAND2_X1 U6505 ( .A1(n8987), .A2(n8101), .ZN(n4963) );
  AND2_X1 U6506 ( .A1(n8383), .A2(n8384), .ZN(n4964) );
  INV_X1 U6507 ( .A(n6614), .ZN(n6605) );
  INV_X1 U6508 ( .A(n8720), .ZN(n5422) );
  AND2_X1 U6509 ( .A1(n5760), .A2(n8642), .ZN(n4965) );
  NAND2_X1 U6510 ( .A1(n9589), .A2(n6288), .ZN(n4966) );
  NOR2_X1 U6511 ( .A1(n8410), .A2(n5880), .ZN(n4968) );
  NAND2_X1 U6512 ( .A1(n5466), .A2(n5465), .ZN(n5484) );
  INV_X1 U6513 ( .A(n8260), .ZN(n8692) );
  INV_X1 U6514 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5965) );
  INV_X1 U6515 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5956) );
  INV_X1 U6516 ( .A(n7316), .ZN(n5814) );
  INV_X1 U6517 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4981) );
  AND2_X1 U6518 ( .A1(n7991), .A2(n7987), .ZN(n7988) );
  INV_X1 U6519 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4975) );
  INV_X1 U6520 ( .A(n8222), .ZN(n8223) );
  INV_X1 U6521 ( .A(n8302), .ZN(n8303) );
  INV_X1 U6522 ( .A(SI_13_), .ZN(n5252) );
  INV_X1 U6523 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5198) );
  INV_X1 U6524 ( .A(n5865), .ZN(n5866) );
  NAND2_X1 U6525 ( .A1(n5668), .A2(n5654), .ZN(n7362) );
  AOI22_X1 U6526 ( .A1(n8601), .A2(n8819), .B1(n8600), .B2(n8599), .ZN(n8602)
         );
  INV_X1 U6527 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5084) );
  NOR2_X1 U6528 ( .A1(n6349), .A2(n9141), .ZN(n6030) );
  NOR2_X1 U6529 ( .A1(n6299), .A2(n6298), .ZN(n6297) );
  INV_X1 U6530 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7415) );
  OR2_X1 U6531 ( .A1(n6339), .A2(n6338), .ZN(n6349) );
  XNOR2_X1 U6532 ( .A(n8304), .B(n8303), .ZN(n8307) );
  OR2_X1 U6533 ( .A1(n6101), .A2(n6956), .ZN(n6092) );
  INV_X1 U6534 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10005) );
  INV_X1 U6535 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5961) );
  INV_X1 U6536 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n5258) );
  INV_X1 U6537 ( .A(n5162), .ZN(n5163) );
  INV_X1 U6538 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5265) );
  INV_X1 U6539 ( .A(n5825), .ZN(n5826) );
  INV_X1 U6540 ( .A(n5065), .ZN(n5302) );
  INV_X1 U6541 ( .A(n8018), .ZN(n7001) );
  AND2_X1 U6542 ( .A1(n5789), .A2(n5652), .ZN(n7228) );
  INV_X1 U6543 ( .A(n8696), .ZN(n8256) );
  AND2_X1 U6544 ( .A1(n6010), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6009) );
  AND2_X1 U6545 ( .A1(n6714), .A2(n9110), .ZN(n6715) );
  OR2_X1 U6546 ( .A1(n9161), .A2(n9162), .ZN(n6781) );
  OR2_X1 U6547 ( .A1(n6322), .A2(n9131), .ZN(n6339) );
  NAND2_X1 U6548 ( .A1(n6297), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6322) );
  INV_X1 U6549 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U6550 ( .A1(n6251), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6280) );
  INV_X1 U6551 ( .A(n8233), .ZN(n8234) );
  OR2_X1 U6552 ( .A1(n7142), .A2(n7139), .ZN(n7148) );
  NAND2_X1 U6553 ( .A1(n5293), .A2(n9985), .ZN(n5316) );
  XNOR2_X1 U6554 ( .A(n5828), .B(n5823), .ZN(n5824) );
  NAND2_X1 U6555 ( .A1(n5824), .A2(n5826), .ZN(n5827) );
  AND2_X1 U6556 ( .A1(n5850), .A2(n5849), .ZN(n5851) );
  OR2_X1 U6557 ( .A1(n5835), .A2(n5834), .ZN(n5836) );
  OR2_X1 U6558 ( .A1(n5940), .A2(n7110), .ZN(n5931) );
  OR2_X1 U6559 ( .A1(n5637), .A2(n7870), .ZN(n6985) );
  INV_X1 U6560 ( .A(n8593), .ZN(n8889) );
  INV_X1 U6561 ( .A(n5791), .ZN(n7767) );
  OR2_X1 U6562 ( .A1(n6985), .A2(n9027), .ZN(n8859) );
  NOR2_X1 U6563 ( .A1(n9907), .A2(n8758), .ZN(n7624) );
  AND2_X1 U6564 ( .A1(n5465), .A2(n5452), .ZN(n5463) );
  OR2_X1 U6565 ( .A1(n7142), .A2(n6880), .ZN(n6881) );
  AND2_X1 U6566 ( .A1(n6783), .A2(n6782), .ZN(n6858) );
  NAND2_X1 U6567 ( .A1(n6195), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6233) );
  OR2_X2 U6568 ( .A1(n6033), .A2(n9121), .ZN(n6043) );
  NAND2_X1 U6569 ( .A1(n6530), .A2(n4259), .ZN(n7142) );
  AND2_X1 U6570 ( .A1(n6391), .A2(n6012), .ZN(n9309) );
  AOI22_X1 U6571 ( .A1(n9202), .A2(n9203), .B1(n9205), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n7386) );
  NAND2_X1 U6572 ( .A1(n8226), .A2(n8227), .ZN(n8302) );
  INV_X1 U6573 ( .A(n9190), .ZN(n9049) );
  AND2_X1 U6574 ( .A1(n7141), .A2(n7140), .ZN(n9480) );
  OAI211_X1 U6575 ( .C1(n8159), .C2(n6798), .A(n9675), .B(n6797), .ZN(n9736)
         );
  XNOR2_X1 U6576 ( .A(n5376), .B(SI_18_), .ZN(n5373) );
  INV_X1 U6577 ( .A(n8429), .ZN(n8439) );
  AND2_X1 U6578 ( .A1(n7330), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8429) );
  INV_X1 U6579 ( .A(n5618), .ZN(n5619) );
  INV_X1 U6580 ( .A(n9827), .ZN(n8579) );
  INV_X1 U6581 ( .A(n9805), .ZN(n9821) );
  INV_X1 U6582 ( .A(n8859), .ZN(n8817) );
  OR2_X1 U6583 ( .A1(n7118), .A2(n7117), .ZN(n8871) );
  NAND2_X1 U6584 ( .A1(n7113), .A2(n8761), .ZN(n8772) );
  NAND2_X1 U6585 ( .A1(n5917), .A2(n5916), .ZN(n7636) );
  AND2_X1 U6586 ( .A1(n8853), .A2(n8852), .ZN(n8976) );
  AND2_X1 U6587 ( .A1(n8867), .A2(n9860), .ZN(n8993) );
  INV_X1 U6588 ( .A(n8993), .ZN(n9902) );
  AND2_X1 U6589 ( .A1(n5915), .A2(n5914), .ZN(n9829) );
  OR2_X1 U6590 ( .A1(n5629), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n5631) );
  INV_X1 U6591 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U6592 ( .A1(n8122), .A2(n6679), .ZN(n8165) );
  INV_X1 U6593 ( .A(n9173), .ZN(n9184) );
  OR2_X1 U6594 ( .A1(n9354), .A2(n6393), .ZN(n6039) );
  OR2_X1 U6595 ( .A1(n6071), .A2(n6070), .ZN(n6072) );
  AND2_X1 U6596 ( .A1(n6923), .A2(n9672), .ZN(n9709) );
  AND2_X1 U6597 ( .A1(n6926), .A2(n7410), .ZN(n9711) );
  INV_X1 U6598 ( .A(n9709), .ZN(n9251) );
  NAND2_X1 U6599 ( .A1(n9312), .A2(n6413), .ZN(n9333) );
  AND2_X1 U6600 ( .A1(n6449), .A2(n9358), .ZN(n9376) );
  AND2_X1 U6601 ( .A1(n6415), .A2(n8144), .ZN(n9504) );
  AND2_X1 U6602 ( .A1(n9733), .A2(n7461), .ZN(n9494) );
  OR2_X1 U6603 ( .A1(n9632), .A2(n6818), .ZN(n9728) );
  NAND2_X1 U6604 ( .A1(n6508), .A2(n7854), .ZN(n7702) );
  AND2_X1 U6605 ( .A1(n9480), .A2(n9632), .ZN(n9624) );
  XNOR2_X1 U6606 ( .A(n6517), .B(P1_IR_REG_24__SCAN_IN), .ZN(n8099) );
  INV_X1 U6607 ( .A(n8585), .ZN(n9817) );
  OR2_X1 U6608 ( .A1(n8426), .A2(n8861), .ZN(n8440) );
  INV_X1 U6609 ( .A(n8445), .ZN(n8432) );
  INV_X1 U6610 ( .A(n8632), .ZN(n8601) );
  INV_X1 U6611 ( .A(n8735), .ZN(n8776) );
  INV_X1 U6612 ( .A(n8834), .ZN(n8453) );
  INV_X1 U6613 ( .A(n8765), .ZN(n8879) );
  OR2_X1 U6614 ( .A1(n7637), .A2(n7636), .ZN(n9923) );
  OR2_X1 U6615 ( .A1(n7637), .A2(n7626), .ZN(n9912) );
  NOR2_X1 U6616 ( .A1(n9830), .A2(n9829), .ZN(n9831) );
  INV_X1 U6617 ( .A(n9831), .ZN(n9834) );
  INV_X1 U6618 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6995) );
  INV_X1 U6619 ( .A(n9167), .ZN(n9182) );
  AND2_X1 U6620 ( .A1(n6819), .A2(n9728), .ZN(n9173) );
  NAND2_X1 U6621 ( .A1(n6532), .A2(n9278), .ZN(n6583) );
  NAND2_X1 U6622 ( .A1(n6027), .A2(n6026), .ZN(n9362) );
  INV_X1 U6623 ( .A(n7688), .ZN(n9194) );
  INV_X1 U6624 ( .A(n9711), .ZN(n9261) );
  INV_X1 U6625 ( .A(n9719), .ZN(n9254) );
  NAND2_X1 U6626 ( .A1(n6929), .A2(n6928), .ZN(n9281) );
  NAND2_X1 U6627 ( .A1(n9733), .A2(n7528), .ZN(n9516) );
  OR2_X1 U6628 ( .A1(n7693), .A2(n7150), .ZN(n9799) );
  NOR2_X1 U6629 ( .A1(n7693), .A2(n7692), .ZN(n9655) );
  INV_X1 U6630 ( .A(n9655), .ZN(n9795) );
  INV_X1 U6631 ( .A(n4259), .ZN(n7854) );
  INV_X1 U6632 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7127) );
  INV_X1 U6633 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6975) );
  NOR2_X1 U6634 ( .A1(n10129), .A2(n10128), .ZN(n10127) );
  NOR2_X1 U6635 ( .A1(n9955), .A2(n9954), .ZN(n9953) );
  INV_X1 U6636 ( .A(n8464), .ZN(P2_U3966) );
  NOR2_X1 U6637 ( .A1(n6928), .A2(P1_U3084), .ZN(P1_U4006) );
  NOR2_X1 U6638 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4973) );
  NAND4_X1 U6639 ( .A1(n4973), .A2(n4972), .A3(n4971), .A4(n5146), .ZN(n5323)
         );
  INV_X1 U6640 ( .A(n5323), .ZN(n4980) );
  NAND3_X1 U6641 ( .A1(n10062), .A2(n4976), .A3(n4975), .ZN(n4977) );
  NOR2_X2 U6642 ( .A1(n5048), .A2(n4977), .ZN(n4979) );
  NOR2_X1 U6643 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4978) );
  INV_X1 U6644 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n4986) );
  INV_X1 U6645 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U6646 ( .A1(n5302), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4992) );
  INV_X1 U6647 ( .A(n5530), .ZN(n4990) );
  NAND2_X1 U6648 ( .A1(n4990), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U6649 ( .A1(n5633), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4994) );
  NAND2_X2 U6650 ( .A1(n4995), .A2(n4996), .ZN(n9030) );
  NAND2_X1 U6651 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n4997) );
  NAND2_X1 U6652 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n9813), .ZN(n5000) );
  MUX2_X1 U6653 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5000), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5004) );
  INV_X1 U6654 ( .A(n5002), .ZN(n5003) );
  INV_X1 U6655 ( .A(n7020), .ZN(n7031) );
  NAND2_X1 U6656 ( .A1(n6983), .A2(n7031), .ZN(n5011) );
  INV_X2 U6657 ( .A(n5231), .ZN(n5972) );
  NAND2_X1 U6658 ( .A1(n5085), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5010) );
  AND2_X1 U6659 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5024) );
  NAND2_X1 U6660 ( .A1(n5164), .A2(n5024), .ZN(n6078) );
  AND2_X1 U6661 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5029) );
  NAND2_X1 U6662 ( .A1(n5972), .A2(n5029), .ZN(n5018) );
  NAND2_X1 U6663 ( .A1(n6078), .A2(n5018), .ZN(n5006) );
  INV_X1 U6664 ( .A(SI_1_), .ZN(n5005) );
  XNOR2_X1 U6665 ( .A(n5006), .B(n5005), .ZN(n5008) );
  MUX2_X1 U6666 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5103), .Z(n5007) );
  NAND2_X2 U6667 ( .A1(n5047), .A2(n5972), .ZN(n5059) );
  NAND2_X1 U6668 ( .A1(n5812), .A2(n8289), .ZN(n5788) );
  NAND2_X1 U6669 ( .A1(n5172), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5015) );
  INV_X1 U6670 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9803) );
  OR2_X1 U6671 ( .A1(n5065), .A2(n9803), .ZN(n5014) );
  INV_X1 U6672 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9802) );
  INV_X1 U6673 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7379) );
  AND4_X2 U6674 ( .A1(n5015), .A2(n5014), .A3(n5013), .A4(n5012), .ZN(n8293)
         );
  NAND2_X1 U6675 ( .A1(n5972), .A2(SI_0_), .ZN(n5017) );
  INV_X1 U6676 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U6677 ( .A1(n5017), .A2(n5016), .ZN(n5019) );
  AND2_X1 U6678 ( .A1(n5019), .A2(n5018), .ZN(n9041) );
  MUX2_X1 U6679 ( .A(n9813), .B(n9041), .S(n4254), .Z(n9839) );
  NAND2_X1 U6680 ( .A1(n8293), .A2(n9839), .ZN(n7119) );
  NAND2_X1 U6681 ( .A1(n5788), .A2(n7119), .ZN(n5652) );
  NAND2_X1 U6682 ( .A1(n5172), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5023) );
  INV_X1 U6683 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7231) );
  INV_X1 U6684 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5020) );
  NOR2_X1 U6685 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5027) );
  INV_X1 U6686 ( .A(n5024), .ZN(n5026) );
  NAND2_X1 U6687 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(SI_1_), .ZN(n5025) );
  OAI21_X1 U6688 ( .B1(n5027), .B2(n5026), .A(n5025), .ZN(n5028) );
  NAND2_X1 U6689 ( .A1(n5231), .A2(n5028), .ZN(n5036) );
  NOR2_X1 U6690 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5032) );
  INV_X1 U6691 ( .A(n5029), .ZN(n5031) );
  NAND2_X1 U6692 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5030) );
  OAI21_X1 U6693 ( .B1(n5032), .B2(n5031), .A(n5030), .ZN(n5033) );
  NAND2_X1 U6694 ( .A1(n5034), .A2(n5033), .ZN(n5035) );
  INV_X1 U6695 ( .A(SI_2_), .ZN(n5051) );
  XNOR2_X1 U6696 ( .A(n5053), .B(n5051), .ZN(n5038) );
  MUX2_X1 U6697 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5103), .Z(n5037) );
  NAND2_X1 U6698 ( .A1(n5085), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5041) );
  OR2_X1 U6699 ( .A1(n5002), .A2(n9015), .ZN(n5039) );
  NAND2_X1 U6700 ( .A1(n4258), .A2(n7039), .ZN(n5040) );
  NAND2_X1 U6701 ( .A1(n7364), .A2(n7363), .ZN(n5062) );
  NAND2_X1 U6702 ( .A1(n5578), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5046) );
  INV_X1 U6703 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7059) );
  OR2_X1 U6704 ( .A1(n5350), .A2(n7059), .ZN(n5045) );
  INV_X1 U6705 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5042) );
  OR2_X1 U6706 ( .A1(n5088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5043) );
  OR2_X1 U6707 ( .A1(n5627), .A2(n9015), .ZN(n5049) );
  INV_X1 U6708 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6955) );
  NAND2_X1 U6709 ( .A1(n5231), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5052) );
  OAI211_X1 U6710 ( .C1(n5231), .C2(n6955), .A(n5052), .B(n5051), .ZN(n5054)
         );
  INV_X1 U6711 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5055) );
  OAI211_X1 U6712 ( .C1(n5231), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5056), .B(
        SI_2_), .ZN(n5057) );
  NAND2_X1 U6713 ( .A1(n5058), .A2(n5057), .ZN(n5071) );
  XNOR2_X1 U6714 ( .A(n5070), .B(n5071), .ZN(n6936) );
  NAND2_X1 U6715 ( .A1(n6936), .A2(n4261), .ZN(n5061) );
  NAND2_X1 U6716 ( .A1(n5085), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5060) );
  OAI211_X1 U6717 ( .C1(n5047), .C2(n7058), .A(n5061), .B(n5060), .ZN(n5823)
         );
  NAND2_X1 U6718 ( .A1(n7203), .A2(n5823), .ZN(n5654) );
  NAND2_X1 U6719 ( .A1(n5578), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5069) );
  INV_X1 U6720 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5063) );
  INV_X1 U6721 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5064) );
  OR2_X1 U6722 ( .A1(n5065), .A2(n5064), .ZN(n5067) );
  XNOR2_X1 U6723 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7579) );
  OR2_X1 U6724 ( .A1(n5088), .A2(n7579), .ZN(n5066) );
  NAND4_X1 U6725 ( .A1(n5069), .A2(n5068), .A3(n5067), .A4(n5066), .ZN(n8462)
         );
  NAND2_X1 U6726 ( .A1(n5073), .A2(SI_3_), .ZN(n5074) );
  MUX2_X1 U6727 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5231), .Z(n5082) );
  NAND2_X1 U6728 ( .A1(n6941), .A2(n4261), .ZN(n5079) );
  OR2_X1 U6729 ( .A1(n5366), .A2(n9015), .ZN(n5077) );
  XNOR2_X1 U6730 ( .A(n5077), .B(P2_IR_REG_4__SCAN_IN), .ZN(n8486) );
  AOI22_X1 U6731 ( .A1(n5085), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n4258), .B2(
        n8486), .ZN(n5078) );
  INV_X1 U6732 ( .A(n5080), .ZN(n5081) );
  NAND2_X1 U6733 ( .A1(n5082), .A2(SI_4_), .ZN(n5083) );
  XNOR2_X1 U6734 ( .A(n5099), .B(n5097), .ZN(n6943) );
  NAND2_X1 U6735 ( .A1(n6943), .A2(n5564), .ZN(n5087) );
  NAND2_X1 U6736 ( .A1(n5366), .A2(n5084), .ZN(n5144) );
  NAND2_X1 U6737 ( .A1(n5144), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5105) );
  XNOR2_X1 U6738 ( .A(n5105), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8499) );
  AOI22_X1 U6739 ( .A1(n5085), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n4258), .B2(
        n8499), .ZN(n5086) );
  NAND2_X1 U6740 ( .A1(n5578), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5096) );
  INV_X1 U6741 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7475) );
  OR2_X1 U6742 ( .A1(n5350), .A2(n7475), .ZN(n5095) );
  INV_X1 U6743 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5090) );
  NAND2_X1 U6744 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5089) );
  NAND2_X1 U6745 ( .A1(n5090), .A2(n5089), .ZN(n5091) );
  NAND2_X1 U6746 ( .A1(n5111), .A2(n5091), .ZN(n7481) );
  OR2_X1 U6747 ( .A1(n5530), .A2(n7481), .ZN(n5094) );
  INV_X1 U6748 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5092) );
  OR2_X1 U6749 ( .A1(n5583), .A2(n5092), .ZN(n5093) );
  NAND2_X1 U6750 ( .A1(n8462), .A2(n9868), .ZN(n7469) );
  INV_X1 U6751 ( .A(n8461), .ZN(n7578) );
  NAND2_X1 U6752 ( .A1(n7578), .A2(n7631), .ZN(n5793) );
  INV_X1 U6753 ( .A(n5097), .ZN(n5098) );
  NAND2_X1 U6754 ( .A1(n5099), .A2(n5098), .ZN(n5102) );
  NAND2_X1 U6755 ( .A1(n5100), .A2(SI_5_), .ZN(n5101) );
  XNOR2_X1 U6756 ( .A(n5104), .B(n5117), .ZN(n6949) );
  NAND2_X1 U6757 ( .A1(n6949), .A2(n5564), .ZN(n5108) );
  INV_X1 U6758 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9958) );
  NAND2_X1 U6759 ( .A1(n5105), .A2(n9958), .ZN(n5106) );
  NAND2_X1 U6760 ( .A1(n5106), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5124) );
  XNOR2_X1 U6761 ( .A(n5124), .B(P2_IR_REG_6__SCAN_IN), .ZN(n8514) );
  AOI22_X1 U6762 ( .A1(n4275), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8514), .B2(
        n4258), .ZN(n5107) );
  NAND2_X1 U6763 ( .A1(n5108), .A2(n5107), .ZN(n7716) );
  NAND2_X1 U6764 ( .A1(n5578), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5116) );
  INV_X1 U6765 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7507) );
  OR2_X1 U6766 ( .A1(n5350), .A2(n7507), .ZN(n5115) );
  INV_X1 U6767 ( .A(n5111), .ZN(n5109) );
  INV_X1 U6768 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6769 ( .A1(n5111), .A2(n5110), .ZN(n5112) );
  NAND2_X1 U6770 ( .A1(n5152), .A2(n5112), .ZN(n7568) );
  OR2_X1 U6771 ( .A1(n5530), .A2(n7568), .ZN(n5114) );
  INV_X1 U6772 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7045) );
  OR2_X1 U6773 ( .A1(n5583), .A2(n7045), .ZN(n5113) );
  NAND4_X1 U6774 ( .A1(n5116), .A2(n5115), .A3(n5114), .A4(n5113), .ZN(n8460)
         );
  XNOR2_X1 U6775 ( .A(n7716), .B(n8460), .ZN(n7504) );
  INV_X1 U6776 ( .A(n8460), .ZN(n7726) );
  NAND2_X1 U6777 ( .A1(n7716), .A2(n7726), .ZN(n5677) );
  INV_X1 U6778 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U6779 ( .A1(n5119), .A2(n5118), .ZN(n5122) );
  NAND2_X1 U6780 ( .A1(n5120), .A2(SI_6_), .ZN(n5121) );
  MUX2_X1 U6781 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5103), .Z(n5137) );
  XNOR2_X1 U6782 ( .A(n5137), .B(SI_7_), .ZN(n5134) );
  XNOR2_X1 U6783 ( .A(n5136), .B(n5134), .ZN(n6953) );
  NAND2_X1 U6784 ( .A1(n6953), .A2(n5564), .ZN(n5128) );
  INV_X1 U6785 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6786 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  NAND2_X1 U6787 ( .A1(n5125), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5126) );
  XNOR2_X1 U6788 ( .A(n5126), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8528) );
  AOI22_X1 U6789 ( .A1(n8528), .A2(n4258), .B1(n5085), .B2(
        P1_DATAO_REG_7__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6790 ( .A1(n5128), .A2(n5127), .ZN(n7780) );
  NAND2_X1 U6791 ( .A1(n5578), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5133) );
  INV_X1 U6792 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7062) );
  OR2_X1 U6793 ( .A1(n5350), .A2(n7062), .ZN(n5132) );
  XNOR2_X1 U6794 ( .A(n5152), .B(n8529), .ZN(n7720) );
  OR2_X1 U6795 ( .A1(n5530), .A2(n7720), .ZN(n5131) );
  INV_X1 U6796 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5129) );
  OR2_X1 U6797 ( .A1(n5583), .A2(n5129), .ZN(n5130) );
  AND2_X1 U6798 ( .A1(n7780), .A2(n7771), .ZN(n5676) );
  OR2_X1 U6799 ( .A1(n7780), .A2(n7771), .ZN(n5679) );
  INV_X1 U6800 ( .A(n5134), .ZN(n5135) );
  NAND2_X1 U6801 ( .A1(n5137), .A2(SI_7_), .ZN(n5138) );
  MUX2_X1 U6802 ( .A(n6965), .B(n6968), .S(n5164), .Z(n5140) );
  INV_X1 U6803 ( .A(SI_8_), .ZN(n5139) );
  NAND2_X1 U6804 ( .A1(n5140), .A2(n5139), .ZN(n5206) );
  INV_X1 U6805 ( .A(n5140), .ZN(n5141) );
  NAND2_X1 U6806 ( .A1(n5141), .A2(SI_8_), .ZN(n5142) );
  NAND2_X1 U6807 ( .A1(n5206), .A2(n5142), .ZN(n5162) );
  NAND2_X1 U6808 ( .A1(n5363), .A2(n5361), .ZN(n5143) );
  NAND2_X1 U6809 ( .A1(n5325), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5145) );
  MUX2_X1 U6810 ( .A(n5145), .B(P2_IR_REG_31__SCAN_IN), .S(n5146), .Z(n5148)
         );
  INV_X1 U6811 ( .A(n5325), .ZN(n5147) );
  NAND2_X1 U6812 ( .A1(n5147), .A2(n5146), .ZN(n5190) );
  NAND2_X1 U6813 ( .A1(n5148), .A2(n5190), .ZN(n8538) );
  INV_X1 U6814 ( .A(n8538), .ZN(n7048) );
  AOI22_X1 U6815 ( .A1(n4275), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7048), .B2(
        n4258), .ZN(n5149) );
  NAND2_X1 U6816 ( .A1(n5578), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5160) );
  INV_X1 U6817 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5150) );
  OR2_X1 U6818 ( .A1(n5350), .A2(n5150), .ZN(n5159) );
  INV_X1 U6819 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5151) );
  OAI21_X1 U6820 ( .B1(n5152), .B2(n8529), .A(n5151), .ZN(n5155) );
  NAND2_X1 U6821 ( .A1(n5155), .A2(n5175), .ZN(n7784) );
  OR2_X1 U6822 ( .A1(n5530), .A2(n7784), .ZN(n5158) );
  INV_X1 U6823 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5156) );
  OR2_X1 U6824 ( .A1(n5583), .A2(n5156), .ZN(n5157) );
  NAND4_X1 U6825 ( .A1(n5160), .A2(n5159), .A3(n5158), .A4(n5157), .ZN(n8458)
         );
  NAND2_X1 U6826 ( .A1(n7783), .A2(n8458), .ZN(n8072) );
  INV_X1 U6827 ( .A(n7783), .ZN(n9886) );
  INV_X1 U6828 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5165) );
  MUX2_X1 U6829 ( .A(n5165), .B(n6975), .S(n5164), .Z(n5167) );
  INV_X1 U6830 ( .A(SI_9_), .ZN(n5166) );
  NAND2_X1 U6831 ( .A1(n5167), .A2(n5166), .ZN(n5207) );
  INV_X1 U6832 ( .A(n5167), .ZN(n5168) );
  NAND2_X1 U6833 ( .A1(n5168), .A2(SI_9_), .ZN(n5210) );
  AND2_X1 U6834 ( .A1(n5207), .A2(n5210), .ZN(n5182) );
  NAND2_X1 U6835 ( .A1(n6969), .A2(n5564), .ZN(n5171) );
  NAND2_X1 U6836 ( .A1(n5190), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5169) );
  XNOR2_X1 U6837 ( .A(n5169), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8562) );
  AOI22_X1 U6838 ( .A1(n4258), .A2(n8562), .B1(n4275), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6839 ( .A1(n5578), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5180) );
  INV_X1 U6840 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5173) );
  OR2_X1 U6841 ( .A1(n5583), .A2(n5173), .ZN(n5179) );
  INV_X1 U6842 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U6843 ( .A1(n5175), .A2(n8557), .ZN(n5176) );
  NAND2_X1 U6844 ( .A1(n5199), .A2(n5176), .ZN(n8083) );
  OR2_X1 U6845 ( .A1(n5530), .A2(n8083), .ZN(n5178) );
  INV_X1 U6846 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7063) );
  OR2_X1 U6847 ( .A1(n5350), .A2(n7063), .ZN(n5177) );
  OR2_X1 U6848 ( .A1(n8085), .A2(n7984), .ZN(n5644) );
  NAND2_X1 U6849 ( .A1(n8085), .A2(n7984), .ZN(n5684) );
  NAND2_X1 U6850 ( .A1(n8089), .A2(n8088), .ZN(n5181) );
  NAND2_X1 U6851 ( .A1(n5181), .A2(n5684), .ZN(n7982) );
  NAND2_X1 U6852 ( .A1(n5183), .A2(n5182), .ZN(n5184) );
  INV_X1 U6853 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5185) );
  MUX2_X1 U6854 ( .A(n6977), .B(n5185), .S(n5103), .Z(n5187) );
  INV_X1 U6855 ( .A(SI_10_), .ZN(n5186) );
  INV_X1 U6856 ( .A(n5187), .ZN(n5188) );
  NAND2_X1 U6857 ( .A1(n5188), .A2(SI_10_), .ZN(n5189) );
  INV_X1 U6858 ( .A(n5190), .ZN(n5192) );
  INV_X1 U6859 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6860 ( .A1(n5192), .A2(n5191), .ZN(n5214) );
  NAND2_X1 U6861 ( .A1(n5214), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5193) );
  XNOR2_X1 U6862 ( .A(n5193), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7064) );
  AOI22_X1 U6863 ( .A1(n7064), .A2(n4258), .B1(n4275), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5194) );
  NAND2_X2 U6864 ( .A1(n5195), .A2(n5194), .ZN(n8028) );
  NAND2_X1 U6865 ( .A1(n4629), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5205) );
  INV_X1 U6866 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5197) );
  OR2_X1 U6867 ( .A1(n5196), .A2(n5197), .ZN(n5204) );
  OR2_X2 U6868 ( .A1(n5199), .A2(n5198), .ZN(n5218) );
  NAND2_X1 U6869 ( .A1(n5199), .A2(n5198), .ZN(n5200) );
  NAND2_X1 U6870 ( .A1(n5218), .A2(n5200), .ZN(n7995) );
  OR2_X1 U6871 ( .A1(n5530), .A2(n7995), .ZN(n5203) );
  INV_X1 U6872 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5201) );
  OR2_X1 U6873 ( .A1(n5350), .A2(n5201), .ZN(n5202) );
  NAND2_X1 U6874 ( .A1(n6978), .A2(n5564), .ZN(n5217) );
  NAND2_X1 U6875 ( .A1(n5237), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5215) );
  XNOR2_X1 U6876 ( .A(n5215), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7065) );
  AOI22_X1 U6877 ( .A1(n7065), .A2(n4258), .B1(n4275), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6878 ( .A1(n5578), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5224) );
  INV_X1 U6879 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7052) );
  OR2_X1 U6880 ( .A1(n5583), .A2(n7052), .ZN(n5223) );
  NAND2_X1 U6881 ( .A1(n5218), .A2(n7916), .ZN(n5219) );
  NAND2_X1 U6882 ( .A1(n5242), .A2(n5219), .ZN(n8025) );
  OR2_X1 U6883 ( .A1(n5530), .A2(n8025), .ZN(n5222) );
  INV_X1 U6884 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5220) );
  OR2_X1 U6885 ( .A1(n5350), .A2(n5220), .ZN(n5221) );
  INV_X1 U6886 ( .A(n5226), .ZN(n5227) );
  NAND2_X1 U6887 ( .A1(n5227), .A2(SI_11_), .ZN(n5228) );
  MUX2_X1 U6888 ( .A(n6995), .B(n5232), .S(n5164), .Z(n5234) );
  INV_X1 U6889 ( .A(SI_12_), .ZN(n5233) );
  NAND2_X1 U6890 ( .A1(n5234), .A2(n5233), .ZN(n5248) );
  INV_X1 U6891 ( .A(n5234), .ZN(n5235) );
  NAND2_X1 U6892 ( .A1(n5235), .A2(SI_12_), .ZN(n5236) );
  NAND2_X1 U6893 ( .A1(n5248), .A2(n5236), .ZN(n5249) );
  XNOR2_X1 U6894 ( .A(n5250), .B(n5249), .ZN(n6990) );
  NAND2_X1 U6895 ( .A1(n6990), .A2(n5564), .ZN(n5240) );
  NAND2_X1 U6896 ( .A1(n5259), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5238) );
  XNOR2_X1 U6897 ( .A(n5238), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7071) );
  AOI22_X1 U6898 ( .A1(n7071), .A2(n4258), .B1(n4275), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n5239) );
  NAND2_X2 U6899 ( .A1(n5240), .A2(n5239), .ZN(n8982) );
  NAND2_X1 U6900 ( .A1(n5578), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5247) );
  INV_X1 U6901 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8112) );
  OR2_X1 U6902 ( .A1(n5350), .A2(n8112), .ZN(n5246) );
  INV_X1 U6903 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U6904 ( .A1(n5242), .A2(n5241), .ZN(n5243) );
  NAND2_X1 U6905 ( .A1(n5279), .A2(n5243), .ZN(n8114) );
  OR2_X1 U6906 ( .A1(n5530), .A2(n8114), .ZN(n5245) );
  INV_X1 U6907 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7152) );
  OR2_X1 U6908 ( .A1(n5583), .A2(n7152), .ZN(n5244) );
  OR2_X1 U6909 ( .A1(n8982), .A2(n8862), .ZN(n5784) );
  AND2_X1 U6910 ( .A1(n5784), .A2(n8107), .ZN(n5689) );
  NAND2_X1 U6911 ( .A1(n8982), .A2(n8862), .ZN(n5783) );
  MUX2_X1 U6912 ( .A(n10071), .B(n5251), .S(n6944), .Z(n5253) );
  NAND2_X1 U6913 ( .A1(n5253), .A2(n5252), .ZN(n5256) );
  INV_X1 U6914 ( .A(n5253), .ZN(n5254) );
  NAND2_X1 U6915 ( .A1(n5254), .A2(SI_13_), .ZN(n5255) );
  MUX2_X1 U6916 ( .A(n5258), .B(n7023), .S(n5103), .Z(n5288) );
  XNOR2_X1 U6917 ( .A(n5292), .B(n5287), .ZN(n6997) );
  NAND2_X1 U6918 ( .A1(n6997), .A2(n5564), .ZN(n5263) );
  INV_X1 U6919 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5260) );
  NAND2_X1 U6920 ( .A1(n5274), .A2(n5260), .ZN(n5261) );
  NAND2_X1 U6921 ( .A1(n5261), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5297) );
  AOI22_X1 U6922 ( .A1(n7491), .A2(n6983), .B1(n4275), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6923 ( .A1(n5281), .A2(n5265), .ZN(n5266) );
  AND2_X1 U6924 ( .A1(n5307), .A2(n5266), .ZN(n8841) );
  NAND2_X1 U6925 ( .A1(n5571), .A2(n8841), .ZN(n5272) );
  INV_X1 U6926 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n5267) );
  OR2_X1 U6927 ( .A1(n5196), .A2(n5267), .ZN(n5271) );
  INV_X1 U6928 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n5268) );
  OR2_X1 U6929 ( .A1(n5350), .A2(n5268), .ZN(n5270) );
  INV_X1 U6930 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7208) );
  OR2_X1 U6931 ( .A1(n5583), .A2(n7208), .ZN(n5269) );
  XNOR2_X1 U6932 ( .A(n5273), .B(n4957), .ZN(n6992) );
  NAND2_X1 U6933 ( .A1(n6992), .A2(n5564), .ZN(n5277) );
  XNOR2_X1 U6934 ( .A(n5274), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7211) );
  NOR2_X1 U6935 ( .A1(n5331), .A2(n10071), .ZN(n5275) );
  AOI21_X1 U6936 ( .B1(n7211), .B2(n4258), .A(n5275), .ZN(n5276) );
  NAND2_X1 U6937 ( .A1(n5578), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5285) );
  INV_X1 U6938 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7160) );
  OR2_X1 U6939 ( .A1(n5350), .A2(n7160), .ZN(n5284) );
  INV_X1 U6940 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6941 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  NAND2_X1 U6942 ( .A1(n5281), .A2(n5280), .ZN(n8875) );
  OR2_X1 U6943 ( .A1(n5530), .A2(n8875), .ZN(n5283) );
  INV_X1 U6944 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9993) );
  OR2_X1 U6945 ( .A1(n5583), .A2(n9993), .ZN(n5282) );
  OR2_X1 U6946 ( .A1(n8977), .A2(n8834), .ZN(n5699) );
  AND2_X1 U6947 ( .A1(n8815), .A2(n5699), .ZN(n5286) );
  NAND2_X1 U6948 ( .A1(n8814), .A2(n5286), .ZN(n5315) );
  INV_X1 U6949 ( .A(n5288), .ZN(n5289) );
  NAND2_X1 U6950 ( .A1(n5289), .A2(SI_14_), .ZN(n5290) );
  MUX2_X1 U6951 ( .A(n7129), .B(n7127), .S(n5103), .Z(n5293) );
  INV_X1 U6952 ( .A(n5293), .ZN(n5294) );
  NAND2_X1 U6953 ( .A1(n5294), .A2(SI_15_), .ZN(n5295) );
  NAND2_X1 U6954 ( .A1(n5316), .A2(n5295), .ZN(n5317) );
  XNOR2_X1 U6955 ( .A(n5318), .B(n5317), .ZN(n7125) );
  NAND2_X1 U6956 ( .A1(n7125), .A2(n5564), .ZN(n5301) );
  INV_X1 U6957 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6958 ( .A1(n5297), .A2(n5296), .ZN(n5298) );
  NAND2_X1 U6959 ( .A1(n5298), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5299) );
  XNOR2_X1 U6960 ( .A(n5299), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7837) );
  AOI22_X1 U6961 ( .A1(n7837), .A2(n4258), .B1(n4275), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6962 ( .A1(n5579), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6963 ( .A1(n5578), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5303) );
  AND2_X1 U6964 ( .A1(n5304), .A2(n5303), .ZN(n5311) );
  INV_X1 U6965 ( .A(n5307), .ZN(n5305) );
  INV_X1 U6966 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6967 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  NAND2_X1 U6968 ( .A1(n5333), .A2(n5308), .ZN(n8822) );
  OR2_X1 U6969 ( .A1(n8822), .A2(n5530), .ZN(n5310) );
  NAND2_X1 U6970 ( .A1(n4629), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6971 ( .A1(n8968), .A2(n8835), .ZN(n5713) );
  NAND2_X1 U6972 ( .A1(n5859), .A2(n8860), .ZN(n5695) );
  NAND2_X1 U6973 ( .A1(n8977), .A2(n8834), .ZN(n8830) );
  NAND2_X1 U6974 ( .A1(n5695), .A2(n8830), .ZN(n5312) );
  NAND2_X1 U6975 ( .A1(n5312), .A2(n8815), .ZN(n5313) );
  MUX2_X1 U6976 ( .A(n7287), .B(n7290), .S(n4257), .Z(n5320) );
  INV_X1 U6977 ( .A(n5320), .ZN(n5321) );
  NAND2_X1 U6978 ( .A1(n5321), .A2(SI_16_), .ZN(n5322) );
  XNOR2_X1 U6979 ( .A(n5338), .B(n4960), .ZN(n7286) );
  INV_X1 U6980 ( .A(n4698), .ZN(n5324) );
  NOR2_X1 U6981 ( .A1(n5325), .A2(n5324), .ZN(n5328) );
  NOR2_X1 U6982 ( .A1(n5328), .A2(n9015), .ZN(n5326) );
  MUX2_X1 U6983 ( .A(n9015), .B(n5326), .S(P2_IR_REG_16__SCAN_IN), .Z(n5330)
         );
  NAND2_X1 U6984 ( .A1(n5328), .A2(n5327), .ZN(n5342) );
  INV_X1 U6985 ( .A(n5342), .ZN(n5329) );
  OAI22_X1 U6986 ( .A1(n7921), .A2(n5047), .B1(n5331), .B2(n7287), .ZN(n5332)
         );
  OR2_X2 U6987 ( .A1(n5333), .A2(n7847), .ZN(n5347) );
  NAND2_X1 U6988 ( .A1(n5333), .A2(n7847), .ZN(n5334) );
  NAND2_X1 U6989 ( .A1(n5347), .A2(n5334), .ZN(n8366) );
  AOI22_X1 U6990 ( .A1(n4629), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n5578), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n5336) );
  NAND2_X1 U6991 ( .A1(n5579), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5335) );
  OAI211_X1 U6992 ( .C1(n8366), .C2(n5530), .A(n5336), .B(n5335), .ZN(n8818)
         );
  INV_X1 U6993 ( .A(n8818), .ZN(n8442) );
  NAND2_X1 U6994 ( .A1(n8962), .A2(n8442), .ZN(n5717) );
  MUX2_X1 U6995 ( .A(n7437), .B(n5341), .S(n4256), .Z(n5357) );
  XNOR2_X1 U6996 ( .A(n5357), .B(SI_17_), .ZN(n5355) );
  XNOR2_X1 U6997 ( .A(n5354), .B(n5355), .ZN(n7341) );
  NAND2_X1 U6998 ( .A1(n7341), .A2(n5564), .ZN(n5345) );
  NAND2_X1 U6999 ( .A1(n5342), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5343) );
  XNOR2_X1 U7000 ( .A(n5343), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8572) );
  AOI22_X1 U7001 ( .A1(n8572), .A2(n6983), .B1(n4275), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n5344) );
  INV_X1 U7002 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9956) );
  NAND2_X1 U7003 ( .A1(n5347), .A2(n9956), .ZN(n5348) );
  NAND2_X1 U7004 ( .A1(n5386), .A2(n5348), .ZN(n8788) );
  OR2_X1 U7005 ( .A1(n8788), .A2(n5530), .ZN(n5353) );
  AOI22_X1 U7006 ( .A1(n4629), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n5578), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n5352) );
  INV_X1 U7007 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n5349) );
  OR2_X1 U7008 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  NAND2_X1 U7009 ( .A1(n8958), .A2(n8415), .ZN(n5723) );
  NAND2_X1 U7010 ( .A1(n5722), .A2(n5723), .ZN(n8246) );
  INV_X1 U7011 ( .A(n5354), .ZN(n5356) );
  INV_X1 U7012 ( .A(n5357), .ZN(n5358) );
  NAND2_X1 U7013 ( .A1(n5358), .A2(SI_17_), .ZN(n5359) );
  MUX2_X1 U7014 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4256), .Z(n5376) );
  NAND2_X1 U7015 ( .A1(n7514), .A2(n5564), .ZN(n5369) );
  NOR2_X1 U7016 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5362) );
  NAND2_X1 U7017 ( .A1(n5381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5367) );
  XNOR2_X1 U7018 ( .A(n5367), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U7019 ( .A1(n4275), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6983), .B2(
        n9822), .ZN(n5368) );
  XNOR2_X1 U7020 ( .A(n5386), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n8778) );
  INV_X1 U7021 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U7022 ( .A1(n5579), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U7023 ( .A1(n5578), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5370) );
  OAI211_X1 U7024 ( .C1(n8574), .C2(n5583), .A(n5371), .B(n5370), .ZN(n5372)
         );
  AOI21_X1 U7025 ( .B1(n8778), .B2(n5571), .A(n5372), .ZN(n8372) );
  NAND2_X1 U7026 ( .A1(n8952), .A2(n8372), .ZN(n5733) );
  NAND2_X1 U7027 ( .A1(n5727), .A2(n5733), .ZN(n8774) );
  MUX2_X1 U7028 ( .A(n7643), .B(n7641), .S(n4256), .Z(n5378) );
  INV_X1 U7029 ( .A(n5378), .ZN(n5379) );
  NAND2_X1 U7030 ( .A1(n5379), .A2(SI_19_), .ZN(n5380) );
  NAND2_X1 U7031 ( .A1(n5394), .A2(n5380), .ZN(n5395) );
  XNOR2_X1 U7032 ( .A(n5396), .B(n5395), .ZN(n7640) );
  NAND2_X1 U7033 ( .A1(n7640), .A2(n5564), .ZN(n5383) );
  AOI22_X1 U7034 ( .A1(n4275), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7627), .B2(
        n6983), .ZN(n5382) );
  INV_X1 U7035 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10037) );
  INV_X1 U7036 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5384) );
  OAI21_X1 U7037 ( .B1(n5386), .B2(n10037), .A(n5384), .ZN(n5387) );
  NAND2_X1 U7038 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n5385) );
  NAND2_X1 U7039 ( .A1(n5387), .A2(n5403), .ZN(n8762) );
  OR2_X1 U7040 ( .A1(n8762), .A2(n5530), .ZN(n5393) );
  INV_X1 U7041 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U7042 ( .A1(n5578), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U7043 ( .A1(n5579), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5388) );
  OAI211_X1 U7044 ( .C1(n5583), .C2(n5390), .A(n5389), .B(n5388), .ZN(n5391)
         );
  INV_X1 U7045 ( .A(n5391), .ZN(n5392) );
  OR2_X1 U7046 ( .A1(n8948), .A2(n8735), .ZN(n5731) );
  NAND2_X1 U7047 ( .A1(n8948), .A2(n8735), .ZN(n5735) );
  MUX2_X1 U7048 ( .A(n7766), .B(n7731), .S(n4256), .Z(n5398) );
  INV_X1 U7049 ( .A(n5398), .ZN(n5399) );
  NAND2_X1 U7050 ( .A1(n5399), .A2(SI_20_), .ZN(n5400) );
  XNOR2_X1 U7051 ( .A(n5411), .B(n5410), .ZN(n7730) );
  NAND2_X1 U7052 ( .A1(n7730), .A2(n5564), .ZN(n5402) );
  NAND2_X1 U7053 ( .A1(n4275), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5401) );
  INV_X1 U7054 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10018) );
  NAND2_X1 U7055 ( .A1(n5403), .A2(n10018), .ZN(n5404) );
  NAND2_X1 U7056 ( .A1(n5436), .A2(n5404), .ZN(n8740) );
  OR2_X1 U7057 ( .A1(n8740), .A2(n5530), .ZN(n5409) );
  INV_X1 U7058 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U7059 ( .A1(n5579), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U7060 ( .A1(n4629), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5405) );
  OAI211_X1 U7061 ( .C1(n5196), .C2(n10090), .A(n5406), .B(n5405), .ZN(n5407)
         );
  INV_X1 U7062 ( .A(n5407), .ZN(n5408) );
  NAND2_X1 U7063 ( .A1(n8942), .A2(n8339), .ZN(n5736) );
  NAND2_X1 U7064 ( .A1(n5737), .A2(n5736), .ZN(n8745) );
  NAND2_X1 U7065 ( .A1(n5411), .A2(n5410), .ZN(n5413) );
  MUX2_X1 U7066 ( .A(n7871), .B(n10033), .S(n4257), .Z(n5424) );
  XNOR2_X1 U7067 ( .A(n5424), .B(SI_21_), .ZN(n5423) );
  XNOR2_X1 U7068 ( .A(n5428), .B(n5423), .ZN(n7853) );
  NAND2_X1 U7069 ( .A1(n7853), .A2(n5564), .ZN(n5415) );
  NAND2_X1 U7070 ( .A1(n4275), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5414) );
  XNOR2_X1 U7071 ( .A(n5436), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U7072 ( .A1(n8723), .A2(n5571), .ZN(n5421) );
  INV_X1 U7073 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n5418) );
  NAND2_X1 U7074 ( .A1(n5578), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U7075 ( .A1(n5579), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5416) );
  OAI211_X1 U7076 ( .C1(n5418), .C2(n5583), .A(n5417), .B(n5416), .ZN(n5419)
         );
  INV_X1 U7077 ( .A(n5419), .ZN(n5420) );
  XNOR2_X1 U7078 ( .A(n8936), .B(n8736), .ZN(n8720) );
  NAND2_X1 U7079 ( .A1(n8936), .A2(n8736), .ZN(n5741) );
  INV_X1 U7080 ( .A(n5423), .ZN(n5427) );
  INV_X1 U7081 ( .A(n5424), .ZN(n5425) );
  NAND2_X1 U7082 ( .A1(n5425), .A2(SI_21_), .ZN(n5426) );
  INV_X1 U7083 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n5429) );
  MUX2_X1 U7084 ( .A(n8173), .B(n5429), .S(n4256), .Z(n5431) );
  INV_X1 U7085 ( .A(SI_22_), .ZN(n5430) );
  NAND2_X1 U7086 ( .A1(n5431), .A2(n5430), .ZN(n5444) );
  INV_X1 U7087 ( .A(n5431), .ZN(n5432) );
  NAND2_X1 U7088 ( .A1(n5432), .A2(SI_22_), .ZN(n5433) );
  NAND2_X1 U7089 ( .A1(n5444), .A2(n5433), .ZN(n5445) );
  XNOR2_X1 U7090 ( .A(n5446), .B(n5445), .ZN(n7980) );
  NAND2_X1 U7091 ( .A1(n7980), .A2(n5564), .ZN(n5435) );
  NAND2_X1 U7092 ( .A1(n4275), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5434) );
  INV_X1 U7093 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8337) );
  INV_X1 U7094 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8404) );
  OAI21_X1 U7095 ( .B1(n5436), .B2(n8337), .A(n8404), .ZN(n5437) );
  NAND2_X1 U7096 ( .A1(n5437), .A2(n5455), .ZN(n8706) );
  OR2_X1 U7097 ( .A1(n8706), .A2(n5530), .ZN(n5443) );
  INV_X1 U7098 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U7099 ( .A1(n5579), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U7100 ( .A1(n5578), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5438) );
  OAI211_X1 U7101 ( .C1(n5440), .C2(n5583), .A(n5439), .B(n5438), .ZN(n5441)
         );
  INV_X1 U7102 ( .A(n5441), .ZN(n5442) );
  NAND2_X1 U7103 ( .A1(n8931), .A2(n8340), .ZN(n5745) );
  INV_X1 U7104 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5448) );
  INV_X1 U7105 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5447) );
  MUX2_X1 U7106 ( .A(n5448), .B(n5447), .S(n4257), .Z(n5450) );
  INV_X1 U7107 ( .A(SI_23_), .ZN(n5449) );
  NAND2_X1 U7108 ( .A1(n5450), .A2(n5449), .ZN(n5465) );
  INV_X1 U7109 ( .A(n5450), .ZN(n5451) );
  NAND2_X1 U7110 ( .A1(n5451), .A2(SI_23_), .ZN(n5452) );
  XNOR2_X1 U7111 ( .A(n5464), .B(n5463), .ZN(n8017) );
  NAND2_X1 U7112 ( .A1(n8017), .A2(n5564), .ZN(n5454) );
  NAND2_X1 U7113 ( .A1(n4275), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5453) );
  INV_X1 U7114 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U7115 ( .A1(n5455), .A2(n8321), .ZN(n5456) );
  AND2_X1 U7116 ( .A1(n5470), .A2(n5456), .ZN(n8693) );
  NAND2_X1 U7117 ( .A1(n8693), .A2(n5571), .ZN(n5462) );
  INV_X1 U7118 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7119 ( .A1(n5578), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U7120 ( .A1(n5579), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5457) );
  OAI211_X1 U7121 ( .C1(n5459), .C2(n5583), .A(n5458), .B(n5457), .ZN(n5460)
         );
  INV_X1 U7122 ( .A(n5460), .ZN(n5461) );
  NAND2_X1 U7123 ( .A1(n5462), .A2(n5461), .ZN(n8713) );
  INV_X1 U7124 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n5467) );
  MUX2_X1 U7125 ( .A(n8119), .B(n5467), .S(n4257), .Z(n5480) );
  XNOR2_X1 U7126 ( .A(n5480), .B(SI_24_), .ZN(n5479) );
  NAND2_X1 U7127 ( .A1(n8098), .A2(n5564), .ZN(n5469) );
  NAND2_X1 U7128 ( .A1(n4275), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5468) );
  INV_X1 U7129 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U7130 ( .A1(n5470), .A2(n8387), .ZN(n5471) );
  NAND2_X1 U7131 ( .A1(n5507), .A2(n5471), .ZN(n8683) );
  OR2_X1 U7132 ( .A1(n8683), .A2(n5530), .ZN(n5477) );
  INV_X1 U7133 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U7134 ( .A1(n5579), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U7135 ( .A1(n5578), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5472) );
  OAI211_X1 U7136 ( .C1(n5474), .C2(n5583), .A(n5473), .B(n5472), .ZN(n5475)
         );
  INV_X1 U7137 ( .A(n5475), .ZN(n5476) );
  NAND2_X1 U7138 ( .A1(n8923), .A2(n8349), .ZN(n5750) );
  INV_X1 U7139 ( .A(n8713), .ZN(n8405) );
  NAND2_X1 U7140 ( .A1(n8926), .A2(n8405), .ZN(n8676) );
  AND2_X1 U7141 ( .A1(n8678), .A2(n8676), .ZN(n5478) );
  INV_X1 U7142 ( .A(n8626), .ZN(n5516) );
  INV_X1 U7143 ( .A(n5479), .ZN(n5483) );
  INV_X1 U7144 ( .A(n5480), .ZN(n5481) );
  NAND2_X1 U7145 ( .A1(n5481), .A2(SI_24_), .ZN(n5482) );
  INV_X1 U7146 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5485) );
  MUX2_X1 U7147 ( .A(n9039), .B(n5485), .S(n4256), .Z(n5487) );
  INV_X1 U7148 ( .A(SI_25_), .ZN(n5486) );
  NAND2_X1 U7149 ( .A1(n5487), .A2(n5486), .ZN(n5490) );
  INV_X1 U7150 ( .A(n5487), .ZN(n5488) );
  NAND2_X1 U7151 ( .A1(n5488), .A2(SI_25_), .ZN(n5489) );
  NAND2_X1 U7152 ( .A1(n5490), .A2(n5489), .ZN(n5503) );
  INV_X1 U7153 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9033) );
  INV_X1 U7154 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5491) );
  MUX2_X1 U7155 ( .A(n9033), .B(n5491), .S(n4256), .Z(n5493) );
  INV_X1 U7156 ( .A(SI_26_), .ZN(n5492) );
  NAND2_X1 U7157 ( .A1(n5493), .A2(n5492), .ZN(n5519) );
  INV_X1 U7158 ( .A(n5493), .ZN(n5494) );
  NAND2_X1 U7159 ( .A1(n5494), .A2(SI_26_), .ZN(n5495) );
  NAND2_X1 U7160 ( .A1(n9032), .A2(n5564), .ZN(n5497) );
  NAND2_X1 U7161 ( .A1(n4275), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5496) );
  INV_X1 U7162 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9991) );
  INV_X1 U7163 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U7164 ( .A1(n5509), .A2(n8425), .ZN(n5498) );
  INV_X1 U7165 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U7166 ( .A1(n5579), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U7167 ( .A1(n5578), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5499) );
  OAI211_X1 U7168 ( .C1(n5501), .C2(n5583), .A(n5500), .B(n5499), .ZN(n5502)
         );
  NAND2_X1 U7169 ( .A1(n8158), .A2(n5564), .ZN(n5506) );
  NAND2_X1 U7170 ( .A1(n4275), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7171 ( .A1(n5507), .A2(n9991), .ZN(n5508) );
  NAND2_X1 U7172 ( .A1(n5509), .A2(n5508), .ZN(n8663) );
  OR2_X1 U7173 ( .A1(n8663), .A2(n5530), .ZN(n5515) );
  INV_X1 U7174 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7175 ( .A1(n5579), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7176 ( .A1(n5578), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5510) );
  OAI211_X1 U7177 ( .C1(n5512), .C2(n5583), .A(n5511), .B(n5510), .ZN(n5513)
         );
  INV_X1 U7178 ( .A(n5513), .ZN(n5514) );
  OR2_X1 U7179 ( .A1(n8916), .A2(n8680), .ZN(n8642) );
  NAND2_X1 U7180 ( .A1(n5516), .A2(n4965), .ZN(n5539) );
  INV_X1 U7181 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9031) );
  INV_X1 U7182 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5520) );
  MUX2_X1 U7183 ( .A(n9031), .B(n5520), .S(n4257), .Z(n5522) );
  INV_X1 U7184 ( .A(SI_27_), .ZN(n5521) );
  NAND2_X1 U7185 ( .A1(n5522), .A2(n5521), .ZN(n5542) );
  INV_X1 U7186 ( .A(n5522), .ZN(n5523) );
  NAND2_X1 U7187 ( .A1(n5523), .A2(SI_27_), .ZN(n5524) );
  NAND2_X1 U7188 ( .A1(n9029), .A2(n5564), .ZN(n5526) );
  NAND2_X1 U7189 ( .A1(n4275), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5525) );
  INV_X1 U7190 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U7191 ( .A1(n5528), .A2(n5527), .ZN(n5529) );
  NAND2_X1 U7192 ( .A1(n5548), .A2(n5529), .ZN(n8622) );
  INV_X1 U7193 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10004) );
  NAND2_X1 U7194 ( .A1(n5578), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7195 ( .A1(n5579), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5531) );
  OAI211_X1 U7196 ( .C1(n5583), .C2(n10004), .A(n5532), .B(n5531), .ZN(n5533)
         );
  INV_X1 U7197 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U7198 ( .A1(n8905), .A2(n8424), .ZN(n5640) );
  NAND2_X1 U7199 ( .A1(n5639), .A2(n5640), .ZN(n8258) );
  AND2_X1 U7200 ( .A1(n8916), .A2(n8680), .ZN(n5755) );
  NAND2_X1 U7201 ( .A1(n5760), .A2(n5755), .ZN(n5536) );
  NAND2_X1 U7202 ( .A1(n8911), .A2(n8631), .ZN(n8627) );
  NAND2_X1 U7203 ( .A1(n5536), .A2(n8627), .ZN(n5537) );
  NOR2_X1 U7204 ( .A1(n8258), .A2(n5537), .ZN(n5538) );
  NAND2_X1 U7205 ( .A1(n8628), .A2(n5639), .ZN(n8264) );
  NAND2_X1 U7206 ( .A1(n5541), .A2(n5540), .ZN(n5543) );
  INV_X1 U7207 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5545) );
  INV_X1 U7208 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5544) );
  MUX2_X1 U7209 ( .A(n5545), .B(n5544), .S(n4256), .Z(n5559) );
  XNOR2_X1 U7210 ( .A(n5559), .B(SI_28_), .ZN(n5556) );
  NAND2_X1 U7211 ( .A1(n9025), .A2(n5564), .ZN(n5547) );
  NAND2_X1 U7212 ( .A1(n4275), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5546) );
  INV_X1 U7213 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6853) );
  OR2_X2 U7214 ( .A1(n5548), .A2(n6853), .ZN(n8609) );
  NAND2_X1 U7215 ( .A1(n5548), .A2(n6853), .ZN(n5549) );
  NAND2_X1 U7216 ( .A1(n8261), .A2(n5571), .ZN(n5555) );
  INV_X1 U7217 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U7218 ( .A1(n5579), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7219 ( .A1(n5578), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5550) );
  OAI211_X1 U7220 ( .C1(n5552), .C2(n5583), .A(n5551), .B(n5550), .ZN(n5553)
         );
  INV_X1 U7221 ( .A(n5553), .ZN(n5554) );
  AND2_X2 U7222 ( .A1(n5555), .A2(n5554), .ZN(n8632) );
  NAND2_X1 U7223 ( .A1(n8900), .A2(n8632), .ZN(n5641) );
  INV_X1 U7224 ( .A(SI_28_), .ZN(n5558) );
  NAND2_X1 U7225 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  INV_X1 U7226 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5562) );
  INV_X1 U7227 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n5561) );
  MUX2_X1 U7228 ( .A(n5562), .B(n5561), .S(n4257), .Z(n5573) );
  XNOR2_X1 U7229 ( .A(n5573), .B(SI_29_), .ZN(n5563) );
  NAND2_X1 U7230 ( .A1(n9022), .A2(n5564), .ZN(n5566) );
  NAND2_X1 U7231 ( .A1(n4275), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n5565) );
  INV_X1 U7232 ( .A(n8609), .ZN(n5572) );
  INV_X1 U7233 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U7234 ( .A1(n5578), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7235 ( .A1(n5579), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5567) );
  OAI211_X1 U7236 ( .C1(n5583), .C2(n5569), .A(n5568), .B(n5567), .ZN(n5570)
         );
  AOI21_X1 U7237 ( .B1(n5572), .B2(n5571), .A(n5570), .ZN(n8268) );
  INV_X1 U7238 ( .A(n5573), .ZN(n5574) );
  NOR2_X1 U7239 ( .A1(n5574), .A2(SI_29_), .ZN(n5575) );
  MUX2_X1 U7240 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4256), .Z(n5593) );
  XNOR2_X1 U7241 ( .A(n5593), .B(SI_30_), .ZN(n5577) );
  INV_X1 U7242 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7243 ( .A1(n5578), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7244 ( .A1(n5579), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5580) );
  OAI211_X1 U7245 ( .C1(n5583), .C2(n5582), .A(n5581), .B(n5580), .ZN(n8599)
         );
  INV_X1 U7246 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7247 ( .A1(n5579), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U7248 ( .A1(n5578), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n5585) );
  OAI211_X1 U7249 ( .C1(n5583), .C2(n5587), .A(n5586), .B(n5585), .ZN(n8588)
         );
  NAND2_X1 U7250 ( .A1(n5590), .A2(n5589), .ZN(n5605) );
  INV_X1 U7251 ( .A(n5593), .ZN(n5592) );
  INV_X1 U7252 ( .A(SI_30_), .ZN(n5591) );
  NOR2_X1 U7253 ( .A1(n5592), .A2(n5591), .ZN(n5594) );
  INV_X1 U7254 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5597) );
  INV_X1 U7255 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5596) );
  MUX2_X1 U7256 ( .A(n5597), .B(n5596), .S(n4256), .Z(n5598) );
  XNOR2_X1 U7257 ( .A(n5598), .B(SI_31_), .ZN(n5599) );
  XNOR2_X1 U7258 ( .A(n5600), .B(n5599), .ZN(n5991) );
  NAND2_X1 U7259 ( .A1(n5991), .A2(n5564), .ZN(n5602) );
  NAND2_X1 U7260 ( .A1(n4275), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n5601) );
  INV_X1 U7261 ( .A(n8588), .ZN(n5775) );
  INV_X1 U7262 ( .A(n8599), .ZN(n5603) );
  NAND2_X1 U7263 ( .A1(n8889), .A2(n5603), .ZN(n5772) );
  INV_X1 U7264 ( .A(n5804), .ZN(n5604) );
  INV_X2 U7265 ( .A(n7627), .ZN(n8758) );
  NAND2_X1 U7266 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  XNOR2_X2 U7267 ( .A(n5610), .B(n5609), .ZN(n7765) );
  AND2_X2 U7268 ( .A1(n7765), .A2(n8758), .ZN(n5934) );
  INV_X1 U7269 ( .A(n5611), .ZN(n5613) );
  NAND2_X1 U7270 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  XNOR2_X2 U7271 ( .A(n5615), .B(n5616), .ZN(n5637) );
  NAND2_X4 U7272 ( .A1(n5934), .A2(n9838), .ZN(n7112) );
  INV_X4 U7273 ( .A(n7112), .ZN(n7328) );
  INV_X1 U7274 ( .A(n7765), .ZN(n5930) );
  AND2_X1 U7275 ( .A1(n5809), .A2(n5930), .ZN(n7117) );
  XNOR2_X1 U7276 ( .A(n5621), .B(n5620), .ZN(n5635) );
  INV_X1 U7277 ( .A(n5635), .ZN(n5935) );
  NAND2_X1 U7278 ( .A1(n5621), .A2(n5620), .ZN(n5622) );
  NAND4_X1 U7279 ( .A1(n4698), .A2(n5627), .A3(n5626), .A4(n5625), .ZN(n5629)
         );
  NAND2_X1 U7280 ( .A1(n5629), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5628) );
  MUX2_X1 U7281 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5628), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5630) );
  NAND2_X1 U7282 ( .A1(n5630), .A2(n5631), .ZN(n9036) );
  NAND2_X1 U7283 ( .A1(n5631), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5632) );
  MUX2_X1 U7284 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5632), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5634) );
  NAND2_X1 U7285 ( .A1(n5634), .A2(n5633), .ZN(n9034) );
  INV_X1 U7286 ( .A(n9830), .ZN(n5636) );
  NOR2_X1 U7287 ( .A1(n9030), .A2(n7004), .ZN(n7014) );
  NAND4_X1 U7288 ( .A1(n5636), .A2(n7108), .A3(n7014), .A4(n8758), .ZN(n5638)
         );
  INV_X1 U7289 ( .A(n5637), .ZN(n5781) );
  MUX2_X1 U7290 ( .A(n7001), .B(n5638), .S(n5781), .Z(n5782) );
  INV_X1 U7291 ( .A(n5639), .ZN(n5643) );
  NAND2_X1 U7292 ( .A1(n5641), .A2(n5640), .ZN(n5642) );
  MUX2_X1 U7293 ( .A(n5643), .B(n5642), .S(n5776), .Z(n5768) );
  OR2_X1 U7294 ( .A1(n8936), .A2(n8736), .ZN(n5738) );
  AND2_X1 U7295 ( .A1(n4963), .A2(n5785), .ZN(n5651) );
  INV_X1 U7296 ( .A(n5644), .ZN(n5649) );
  NAND2_X1 U7297 ( .A1(n5785), .A2(n5684), .ZN(n5645) );
  MUX2_X1 U7298 ( .A(n5649), .B(n5645), .S(n5776), .Z(n5647) );
  INV_X1 U7299 ( .A(n5786), .ZN(n5646) );
  NAND2_X1 U7300 ( .A1(n8107), .A2(n5786), .ZN(n5648) );
  AOI21_X1 U7301 ( .B1(n5686), .B2(n5649), .A(n5648), .ZN(n5650) );
  MUX2_X1 U7302 ( .A(n5651), .B(n5650), .S(n5776), .Z(n5688) );
  INV_X1 U7303 ( .A(n8293), .ZN(n8465) );
  INV_X1 U7304 ( .A(n9839), .ZN(n7327) );
  NAND2_X1 U7305 ( .A1(n8465), .A2(n7327), .ZN(n5787) );
  AND2_X1 U7306 ( .A1(n5787), .A2(n5809), .ZN(n5661) );
  OAI211_X1 U7307 ( .C1(n5652), .C2(n5661), .A(n5664), .B(n5789), .ZN(n5653)
         );
  NAND3_X1 U7308 ( .A1(n5653), .A2(n5776), .A3(n7363), .ZN(n5656) );
  AOI21_X1 U7309 ( .B1(n4294), .B2(n5654), .A(n5778), .ZN(n5655) );
  AOI21_X1 U7310 ( .B1(n5656), .B2(n4260), .A(n5655), .ZN(n5660) );
  NAND2_X1 U7311 ( .A1(n5793), .A2(n4294), .ZN(n5658) );
  MUX2_X1 U7312 ( .A(n5658), .B(n5657), .S(n5776), .Z(n5670) );
  AND2_X1 U7313 ( .A1(n5677), .A2(n5793), .ZN(n5659) );
  OAI22_X1 U7314 ( .A1(n5660), .A2(n5670), .B1(n5778), .B2(n5659), .ZN(n5667)
         );
  OR2_X1 U7315 ( .A1(n7716), .A2(n7726), .ZN(n5671) );
  INV_X1 U7316 ( .A(n5661), .ZN(n5663) );
  INV_X1 U7317 ( .A(n5789), .ZN(n5662) );
  OAI211_X1 U7318 ( .C1(n5663), .C2(n5662), .A(n5788), .B(n7363), .ZN(n5665)
         );
  NAND3_X1 U7319 ( .A1(n5665), .A2(n5778), .A3(n5664), .ZN(n5666) );
  NAND3_X1 U7320 ( .A1(n5667), .A2(n5671), .A3(n5666), .ZN(n5675) );
  AOI22_X1 U7321 ( .A1(n5670), .A2(n5792), .B1(n5669), .B2(n5668), .ZN(n5673)
         );
  INV_X1 U7322 ( .A(n5671), .ZN(n5672) );
  OAI21_X1 U7323 ( .B1(n5673), .B2(n5672), .A(n5778), .ZN(n5674) );
  INV_X1 U7324 ( .A(n5676), .ZN(n5678) );
  MUX2_X1 U7325 ( .A(n5679), .B(n5678), .S(n5776), .Z(n5680) );
  NAND2_X1 U7326 ( .A1(n8458), .A2(n5776), .ZN(n5682) );
  INV_X1 U7327 ( .A(n8458), .ZN(n7725) );
  NAND2_X1 U7328 ( .A1(n7725), .A2(n5778), .ZN(n5681) );
  MUX2_X1 U7329 ( .A(n5682), .B(n5681), .S(n7783), .Z(n5683) );
  NAND2_X1 U7330 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  NAND2_X1 U7331 ( .A1(n5688), .A2(n5687), .ZN(n5694) );
  AND2_X2 U7332 ( .A1(n8815), .A2(n5695), .ZN(n8239) );
  INV_X1 U7333 ( .A(n5689), .ZN(n5691) );
  OAI21_X1 U7334 ( .B1(n5778), .B2(n4963), .A(n5783), .ZN(n5690) );
  AOI21_X1 U7335 ( .B1(n5778), .B2(n5691), .A(n5690), .ZN(n5693) );
  OR2_X1 U7336 ( .A1(n8977), .A2(n5776), .ZN(n5708) );
  NAND2_X1 U7337 ( .A1(n8977), .A2(n5776), .ZN(n5705) );
  MUX2_X1 U7338 ( .A(n5708), .B(n5705), .S(n8834), .Z(n5692) );
  NAND4_X1 U7339 ( .A1(n5694), .A2(n8239), .A3(n5693), .A4(n5692), .ZN(n5712)
         );
  MUX2_X1 U7340 ( .A(n5695), .B(n8815), .S(n5776), .Z(n5711) );
  INV_X1 U7341 ( .A(n8862), .ZN(n8454) );
  NAND2_X1 U7342 ( .A1(n8454), .A2(n5776), .ZN(n5700) );
  NOR2_X1 U7343 ( .A1(n5700), .A2(n8834), .ZN(n5697) );
  NAND2_X1 U7344 ( .A1(n8862), .A2(n5778), .ZN(n5701) );
  NAND2_X1 U7345 ( .A1(n8982), .A2(n5701), .ZN(n5696) );
  OAI21_X1 U7346 ( .B1(n8982), .B2(n5697), .A(n5696), .ZN(n5698) );
  NAND2_X1 U7347 ( .A1(n5699), .A2(n5698), .ZN(n5707) );
  INV_X1 U7348 ( .A(n5700), .ZN(n5703) );
  OAI21_X1 U7349 ( .B1(n8453), .B2(n5701), .A(n8982), .ZN(n5702) );
  OAI21_X1 U7350 ( .B1(n5703), .B2(n8982), .A(n5702), .ZN(n5704) );
  NAND2_X1 U7351 ( .A1(n8830), .A2(n5704), .ZN(n5706) );
  AOI22_X1 U7352 ( .A1(n5708), .A2(n5707), .B1(n5706), .B2(n5705), .ZN(n5709)
         );
  INV_X1 U7353 ( .A(n8239), .ZN(n5797) );
  OR2_X1 U7354 ( .A1(n5709), .A2(n5797), .ZN(n5710) );
  NAND4_X1 U7355 ( .A1(n8825), .A2(n5712), .A3(n5711), .A4(n5710), .ZN(n5716)
         );
  MUX2_X1 U7356 ( .A(n5714), .B(n5713), .S(n5776), .Z(n5715) );
  MUX2_X1 U7357 ( .A(n5718), .B(n5717), .S(n5776), .Z(n5719) );
  NAND3_X1 U7358 ( .A1(n4478), .A2(n5720), .A3(n5719), .ZN(n5721) );
  INV_X1 U7359 ( .A(n5722), .ZN(n5725) );
  NAND2_X1 U7360 ( .A1(n5733), .A2(n5723), .ZN(n5724) );
  MUX2_X1 U7361 ( .A(n5725), .B(n5724), .S(n5778), .Z(n5726) );
  NAND2_X1 U7362 ( .A1(n5728), .A2(n5737), .ZN(n5729) );
  NAND3_X1 U7363 ( .A1(n5729), .A2(n5736), .A3(n5741), .ZN(n5730) );
  NAND3_X1 U7364 ( .A1(n5748), .A2(n5738), .A3(n5730), .ZN(n5744) );
  INV_X1 U7365 ( .A(n5731), .ZN(n5732) );
  AOI21_X1 U7366 ( .B1(n5734), .B2(n5733), .A(n5732), .ZN(n5740) );
  NAND2_X1 U7367 ( .A1(n5736), .A2(n5735), .ZN(n5739) );
  OAI211_X1 U7368 ( .C1(n5740), .C2(n5739), .A(n5738), .B(n5737), .ZN(n5742)
         );
  NAND3_X1 U7369 ( .A1(n5745), .A2(n5742), .A3(n5741), .ZN(n5743) );
  NAND3_X1 U7370 ( .A1(n5749), .A2(n5745), .A3(n8696), .ZN(n5746) );
  OAI211_X1 U7371 ( .C1(n8405), .C2(n8926), .A(n8678), .B(n5746), .ZN(n5747)
         );
  NAND2_X1 U7372 ( .A1(n5747), .A2(n5750), .ZN(n5753) );
  NAND3_X1 U7373 ( .A1(n5749), .A2(n5748), .A3(n8696), .ZN(n5751) );
  AND3_X1 U7374 ( .A1(n5751), .A2(n8676), .A3(n5750), .ZN(n5752) );
  MUX2_X1 U7375 ( .A(n5753), .B(n5752), .S(n5776), .Z(n5759) );
  XNOR2_X1 U7376 ( .A(n8916), .B(n8451), .ZN(n8655) );
  OAI21_X1 U7377 ( .B1(n5778), .B2(n8654), .A(n8655), .ZN(n5758) );
  NAND2_X1 U7378 ( .A1(n5760), .A2(n5778), .ZN(n5754) );
  OAI21_X1 U7379 ( .B1(n8639), .B2(n5755), .A(n5754), .ZN(n5757) );
  OR3_X1 U7380 ( .A1(n8916), .A2(n8680), .A3(n5776), .ZN(n5756) );
  OAI211_X1 U7381 ( .C1(n5759), .C2(n5758), .A(n5757), .B(n5756), .ZN(n5762)
         );
  MUX2_X1 U7382 ( .A(n8627), .B(n5760), .S(n5776), .Z(n5761) );
  NAND3_X1 U7383 ( .A1(n5762), .A2(n5761), .A3(n4552), .ZN(n5764) );
  NAND2_X1 U7384 ( .A1(n5764), .A2(n5763), .ZN(n5767) );
  AND2_X1 U7385 ( .A1(n8601), .A2(n8900), .ZN(n5766) );
  INV_X1 U7386 ( .A(n8900), .ZN(n8263) );
  MUX2_X1 U7387 ( .A(n8632), .B(n8263), .S(n5778), .Z(n5765) );
  MUX2_X1 U7388 ( .A(n5771), .B(n5770), .S(n5776), .Z(n5773) );
  MUX2_X1 U7389 ( .A(n5776), .B(n5775), .S(n5774), .Z(n5777) );
  OAI21_X1 U7390 ( .B1(n5778), .B2(n8588), .A(n5777), .ZN(n5779) );
  NAND2_X1 U7391 ( .A1(n5784), .A2(n5783), .ZN(n8109) );
  NAND2_X1 U7392 ( .A1(n5786), .A2(n5785), .ZN(n7993) );
  NAND2_X1 U7393 ( .A1(n7119), .A2(n5787), .ZN(n9840) );
  NOR4_X1 U7394 ( .A1(n9840), .A2(n7201), .A3(n7198), .A4(n7765), .ZN(n5790)
         );
  NAND3_X1 U7395 ( .A1(n5790), .A2(n4260), .A3(n7193), .ZN(n5794) );
  NAND2_X1 U7396 ( .A1(n5793), .A2(n5792), .ZN(n7472) );
  NAND4_X1 U7397 ( .A1(n8030), .A2(n8088), .A3(n5795), .A4(n4912), .ZN(n5796)
         );
  NOR4_X1 U7398 ( .A1(n5797), .A2(n8109), .A3(n7993), .A4(n5796), .ZN(n5798)
         );
  XNOR2_X1 U7399 ( .A(n8977), .B(n8453), .ZN(n8863) );
  NAND4_X1 U7400 ( .A1(n8809), .A2(n8825), .A3(n5798), .A4(n8863), .ZN(n5799)
         );
  NOR4_X1 U7401 ( .A1(n4469), .A2(n8774), .A3(n8246), .A4(n5799), .ZN(n5800)
         );
  NAND4_X1 U7402 ( .A1(n8712), .A2(n4732), .A3(n5800), .A4(n5422), .ZN(n5801)
         );
  NOR4_X1 U7403 ( .A1(n8639), .A2(n8256), .A3(n4543), .A4(n5801), .ZN(n5802)
         );
  NAND4_X1 U7404 ( .A1(n8265), .A2(n4552), .A3(n5802), .A4(n8655), .ZN(n5803)
         );
  OAI22_X1 U7405 ( .A1(n5806), .A2(n5809), .B1(n5930), .B2(n4669), .ZN(n5808)
         );
  NAND2_X1 U7406 ( .A1(n5833), .A2(n7327), .ZN(n5811) );
  NAND2_X1 U7407 ( .A1(n7326), .A2(n5811), .ZN(n7317) );
  NAND2_X1 U7408 ( .A1(n7317), .A2(n7316), .ZN(n5813) );
  NAND2_X1 U7409 ( .A1(n5813), .A2(n7318), .ZN(n5817) );
  NAND2_X1 U7410 ( .A1(n5819), .A2(n5818), .ZN(n7315) );
  NAND2_X1 U7411 ( .A1(n5815), .A2(n5814), .ZN(n5816) );
  NAND3_X1 U7412 ( .A1(n5817), .A2(n7315), .A3(n5816), .ZN(n5822) );
  INV_X1 U7413 ( .A(n5818), .ZN(n5821) );
  INV_X1 U7414 ( .A(n5819), .ZN(n5820) );
  NAND2_X1 U7415 ( .A1(n5821), .A2(n5820), .ZN(n7314) );
  NAND2_X1 U7416 ( .A1(n5822), .A2(n7314), .ZN(n8277) );
  OR2_X1 U7417 ( .A1(n7203), .A2(n7328), .ZN(n5825) );
  INV_X1 U7418 ( .A(n9868), .ZN(n7477) );
  XNOR2_X1 U7419 ( .A(n7477), .B(n5828), .ZN(n5829) );
  AND2_X1 U7420 ( .A1(n7112), .A2(n8462), .ZN(n5830) );
  AND2_X1 U7421 ( .A1(n5829), .A2(n5830), .ZN(n7575) );
  INV_X1 U7422 ( .A(n5829), .ZN(n5832) );
  INV_X1 U7423 ( .A(n5830), .ZN(n5831) );
  NAND2_X1 U7424 ( .A1(n5832), .A2(n5831), .ZN(n7573) );
  XNOR2_X1 U7425 ( .A(n7500), .B(n4274), .ZN(n5835) );
  NAND2_X1 U7426 ( .A1(n7112), .A2(n8461), .ZN(n5834) );
  XNOR2_X1 U7427 ( .A(n5835), .B(n5834), .ZN(n7334) );
  XNOR2_X1 U7428 ( .A(n7716), .B(n5909), .ZN(n5838) );
  NAND2_X1 U7429 ( .A1(n7112), .A2(n8460), .ZN(n5837) );
  NAND2_X1 U7430 ( .A1(n5838), .A2(n5837), .ZN(n5839) );
  OAI21_X1 U7431 ( .B1(n5838), .B2(n5837), .A(n5839), .ZN(n7567) );
  INV_X1 U7432 ( .A(n5839), .ZN(n5840) );
  NOR2_X1 U7433 ( .A1(n7771), .A2(n7328), .ZN(n5841) );
  XNOR2_X1 U7434 ( .A(n7780), .B(n5828), .ZN(n5842) );
  XOR2_X1 U7435 ( .A(n5841), .B(n5842), .Z(n7560) );
  XNOR2_X1 U7436 ( .A(n9886), .B(n4274), .ZN(n5844) );
  NAND2_X1 U7437 ( .A1(n7112), .A2(n8458), .ZN(n5843) );
  XNOR2_X1 U7438 ( .A(n5844), .B(n5843), .ZN(n7594) );
  XNOR2_X1 U7439 ( .A(n8085), .B(n5909), .ZN(n5845) );
  OR2_X1 U7440 ( .A1(n7984), .A2(n7328), .ZN(n5846) );
  NAND2_X1 U7441 ( .A1(n5845), .A2(n5846), .ZN(n6872) );
  INV_X1 U7442 ( .A(n5845), .ZN(n5848) );
  INV_X1 U7443 ( .A(n5846), .ZN(n5847) );
  NAND2_X1 U7444 ( .A1(n5848), .A2(n5847), .ZN(n6874) );
  NOR2_X1 U7445 ( .A1(n8021), .A2(n7328), .ZN(n5849) );
  XNOR2_X1 U7446 ( .A(n8987), .B(n4274), .ZN(n5852) );
  NOR2_X1 U7447 ( .A1(n8101), .A2(n7328), .ZN(n5853) );
  XNOR2_X1 U7448 ( .A(n5852), .B(n5853), .ZN(n7914) );
  NOR2_X1 U7449 ( .A1(n8862), .A2(n7328), .ZN(n5854) );
  XNOR2_X1 U7450 ( .A(n8982), .B(n4274), .ZN(n5855) );
  XOR2_X1 U7451 ( .A(n5854), .B(n5855), .Z(n8002) );
  NOR2_X1 U7452 ( .A1(n8834), .A2(n7328), .ZN(n5856) );
  XNOR2_X1 U7453 ( .A(n8977), .B(n4274), .ZN(n5857) );
  XOR2_X1 U7454 ( .A(n5856), .B(n5857), .Z(n8066) );
  OR2_X1 U7455 ( .A1(n8860), .A2(n7328), .ZN(n5860) );
  INV_X1 U7456 ( .A(n5860), .ZN(n5863) );
  XNOR2_X1 U7457 ( .A(n5859), .B(n5909), .ZN(n5861) );
  INV_X1 U7458 ( .A(n5861), .ZN(n5862) );
  AOI21_X1 U7459 ( .B1(n5863), .B2(n5862), .A(n8355), .ZN(n8313) );
  NAND2_X1 U7460 ( .A1(n8312), .A2(n8313), .ZN(n8311) );
  XNOR2_X1 U7461 ( .A(n8968), .B(n4274), .ZN(n8358) );
  NOR2_X1 U7462 ( .A1(n8835), .A2(n7328), .ZN(n8437) );
  INV_X1 U7463 ( .A(n8355), .ZN(n5864) );
  OAI21_X1 U7464 ( .B1(n8358), .B2(n8437), .A(n5864), .ZN(n5865) );
  NAND2_X1 U7465 ( .A1(n8311), .A2(n5866), .ZN(n5870) );
  XNOR2_X1 U7466 ( .A(n8804), .B(n4274), .ZN(n5868) );
  NAND2_X1 U7467 ( .A1(n8818), .A2(n7112), .ZN(n5867) );
  NAND2_X1 U7468 ( .A1(n5868), .A2(n5867), .ZN(n5871) );
  OAI21_X1 U7469 ( .B1(n5868), .B2(n5867), .A(n5871), .ZN(n8361) );
  AOI21_X1 U7470 ( .B1(n8437), .B2(n8358), .A(n8361), .ZN(n5869) );
  NAND2_X1 U7471 ( .A1(n8363), .A2(n5871), .ZN(n8371) );
  INV_X1 U7472 ( .A(n8371), .ZN(n5875) );
  XNOR2_X1 U7473 ( .A(n8958), .B(n4274), .ZN(n5877) );
  NOR2_X1 U7474 ( .A1(n8415), .A2(n7328), .ZN(n5876) );
  XNOR2_X1 U7475 ( .A(n5877), .B(n5876), .ZN(n8410) );
  XNOR2_X1 U7476 ( .A(n8952), .B(n4274), .ZN(n5872) );
  NOR2_X1 U7477 ( .A1(n8372), .A2(n7328), .ZN(n5873) );
  NAND2_X1 U7478 ( .A1(n5872), .A2(n5873), .ZN(n5878) );
  INV_X1 U7479 ( .A(n5878), .ZN(n5874) );
  XOR2_X1 U7480 ( .A(n5873), .B(n5872), .Z(n8413) );
  NOR2_X1 U7481 ( .A1(n5874), .A2(n8413), .ZN(n5880) );
  NAND2_X1 U7482 ( .A1(n5877), .A2(n5876), .ZN(n8411) );
  AND2_X1 U7483 ( .A1(n8411), .A2(n5878), .ZN(n5879) );
  OR2_X1 U7484 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  XNOR2_X1 U7485 ( .A(n8948), .B(n5909), .ZN(n5883) );
  NAND2_X1 U7486 ( .A1(n8776), .A2(n7112), .ZN(n5882) );
  NAND2_X1 U7487 ( .A1(n5883), .A2(n5882), .ZN(n5884) );
  OAI21_X1 U7488 ( .B1(n5883), .B2(n5882), .A(n5884), .ZN(n8329) );
  XNOR2_X1 U7489 ( .A(n8942), .B(n4274), .ZN(n5888) );
  NOR2_X1 U7490 ( .A1(n8339), .A2(n7328), .ZN(n5887) );
  XNOR2_X1 U7491 ( .A(n5888), .B(n5887), .ZN(n8393) );
  INV_X1 U7492 ( .A(n8393), .ZN(n5885) );
  NAND2_X1 U7493 ( .A1(n5888), .A2(n5887), .ZN(n5889) );
  NOR2_X1 U7494 ( .A1(n8736), .A2(n7328), .ZN(n5891) );
  XNOR2_X1 U7495 ( .A(n8936), .B(n4274), .ZN(n5893) );
  XOR2_X1 U7496 ( .A(n5891), .B(n5893), .Z(n8336) );
  XNOR2_X1 U7497 ( .A(n8931), .B(n4274), .ZN(n8401) );
  NOR2_X1 U7498 ( .A1(n8340), .A2(n7328), .ZN(n5890) );
  NOR2_X1 U7499 ( .A1(n8401), .A2(n5890), .ZN(n5897) );
  NAND2_X1 U7500 ( .A1(n5893), .A2(n5891), .ZN(n8398) );
  INV_X1 U7501 ( .A(n5890), .ZN(n8400) );
  NAND2_X1 U7502 ( .A1(n8398), .A2(n8400), .ZN(n5895) );
  INV_X1 U7503 ( .A(n5891), .ZN(n5892) );
  NOR2_X1 U7504 ( .A1(n5892), .A2(n8340), .ZN(n5894) );
  AOI22_X1 U7505 ( .A1(n8401), .A2(n5895), .B1(n5894), .B2(n5893), .ZN(n5896)
         );
  XNOR2_X1 U7506 ( .A(n8926), .B(n4274), .ZN(n5899) );
  XNOR2_X1 U7507 ( .A(n8923), .B(n4274), .ZN(n8383) );
  NOR2_X1 U7508 ( .A1(n8383), .A2(n8690), .ZN(n5898) );
  NAND2_X1 U7509 ( .A1(n8713), .A2(n7112), .ZN(n8382) );
  NAND2_X1 U7510 ( .A1(n5900), .A2(n5899), .ZN(n8381) );
  NOR2_X1 U7511 ( .A1(n8349), .A2(n7328), .ZN(n8384) );
  NOR2_X1 U7512 ( .A1(n8383), .A2(n8384), .ZN(n5901) );
  NOR2_X1 U7513 ( .A1(n5902), .A2(n4964), .ZN(n5903) );
  XNOR2_X1 U7514 ( .A(n8916), .B(n4274), .ZN(n8346) );
  NOR2_X1 U7515 ( .A1(n8680), .A2(n7328), .ZN(n8347) );
  XNOR2_X1 U7516 ( .A(n8911), .B(n4274), .ZN(n5906) );
  NOR2_X1 U7517 ( .A1(n8631), .A2(n7328), .ZN(n5905) );
  NAND2_X1 U7518 ( .A1(n5906), .A2(n5905), .ZN(n5908) );
  OAI21_X1 U7519 ( .B1(n5906), .B2(n5905), .A(n5908), .ZN(n8420) );
  INV_X1 U7520 ( .A(n8420), .ZN(n5907) );
  NAND2_X1 U7521 ( .A1(n8422), .A2(n5908), .ZN(n5912) );
  XNOR2_X1 U7522 ( .A(n8905), .B(n5909), .ZN(n5911) );
  INV_X1 U7523 ( .A(n8424), .ZN(n8449) );
  NAND2_X1 U7524 ( .A1(n8449), .A2(n7112), .ZN(n5910) );
  NOR2_X1 U7525 ( .A1(n5911), .A2(n5910), .ZN(n6839) );
  AOI21_X1 U7526 ( .B1(n5911), .B2(n5910), .A(n6839), .ZN(n5929) );
  NAND2_X1 U7527 ( .A1(n5912), .A2(n5929), .ZN(n6841) );
  XNOR2_X1 U7529 ( .A(n8121), .B(P2_B_REG_SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7530 ( .A1(n5913), .A2(n9036), .ZN(n5915) );
  INV_X1 U7531 ( .A(n9034), .ZN(n5914) );
  INV_X1 U7532 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9832) );
  NAND2_X1 U7533 ( .A1(n9829), .A2(n9832), .ZN(n5917) );
  AND2_X1 U7534 ( .A1(n8121), .A2(n9034), .ZN(n9833) );
  INV_X1 U7535 ( .A(n9833), .ZN(n5916) );
  INV_X1 U7536 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9835) );
  AND2_X1 U7537 ( .A1(n9034), .A2(n9036), .ZN(n9836) );
  NOR2_X1 U7538 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .ZN(
        n9970) );
  NOR4_X1 U7539 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5920) );
  NOR4_X1 U7540 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5919) );
  NOR4_X1 U7541 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5918) );
  AND4_X1 U7542 ( .A1(n9970), .A2(n5920), .A3(n5919), .A4(n5918), .ZN(n5926)
         );
  NOR4_X1 U7543 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5924) );
  NOR4_X1 U7544 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5923) );
  NOR4_X1 U7545 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n5922) );
  NOR4_X1 U7546 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n5921) );
  AND4_X1 U7547 ( .A1(n5924), .A2(n5923), .A3(n5922), .A4(n5921), .ZN(n5925)
         );
  NAND2_X1 U7548 ( .A1(n5926), .A2(n5925), .ZN(n5927) );
  NAND2_X1 U7549 ( .A1(n9829), .A2(n5927), .ZN(n7105) );
  NAND3_X1 U7550 ( .A1(n7626), .A2(n7625), .A3(n7105), .ZN(n5933) );
  INV_X1 U7551 ( .A(n5934), .ZN(n5939) );
  INV_X1 U7552 ( .A(n6985), .ZN(n7002) );
  OR3_X2 U7553 ( .A1(n5940), .A2(n8988), .A3(n7002), .ZN(n8447) );
  INV_X1 U7554 ( .A(n8447), .ZN(n8314) );
  OAI211_X1 U7555 ( .C1(n5912), .C2(n5929), .A(n5928), .B(n8314), .ZN(n5946)
         );
  NAND2_X1 U7556 ( .A1(n9838), .A2(n5930), .ZN(n7110) );
  INV_X1 U7557 ( .A(n7624), .ZN(n5932) );
  NAND2_X1 U7558 ( .A1(n5933), .A2(n5932), .ZN(n5938) );
  NOR2_X1 U7559 ( .A1(n6985), .A2(n5934), .ZN(n7103) );
  NOR2_X1 U7560 ( .A1(n7103), .A2(n5935), .ZN(n5936) );
  AND2_X1 U7561 ( .A1(n5936), .A2(n6999), .ZN(n5937) );
  NAND2_X1 U7562 ( .A1(n5938), .A2(n5937), .ZN(n7330) );
  NOR2_X1 U7563 ( .A1(n8622), .A2(n8439), .ZN(n5942) );
  INV_X1 U7564 ( .A(n7004), .ZN(n9027) );
  OAI22_X1 U7565 ( .A1(n8632), .A2(n8441), .B1(n8631), .B2(n8440), .ZN(n5941)
         );
  AOI211_X1 U7566 ( .C1(P2_REG3_REG_27__SCAN_IN), .C2(P2_U3152), .A(n5942), 
        .B(n5941), .ZN(n5943) );
  INV_X1 U7567 ( .A(n5944), .ZN(n5945) );
  INV_X2 U7568 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X2 U7569 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5949) );
  NOR2_X2 U7570 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5948) );
  NOR2_X2 U7571 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5947) );
  INV_X2 U7572 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7573 ( .A1(n6411), .A2(n5959), .ZN(n5952) );
  NAND2_X1 U7574 ( .A1(n6410), .A2(n5955), .ZN(n5953) );
  INV_X1 U7575 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5958) );
  INV_X1 U7576 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5957) );
  NOR2_X1 U7577 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5963) );
  NOR2_X1 U7578 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5962) );
  NAND2_X1 U7579 ( .A1(n5975), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7580 ( .A1(n9019), .A2(n6386), .ZN(n5974) );
  AND2_X2 U7581 ( .A1(n6124), .A2(n5972), .ZN(n6143) );
  INV_X2 U7582 ( .A(n6143), .ZN(n6106) );
  NAND2_X1 U7583 ( .A1(n6387), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5973) );
  NOR2_X1 U7584 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n5976) );
  NAND2_X1 U7585 ( .A1(n5978), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5977) );
  AND2_X2 U7586 ( .A1(n5979), .A2(n5980), .ZN(n9666) );
  INV_X1 U7587 ( .A(n6000), .ZN(n5983) );
  INV_X1 U7588 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7589 ( .A1(n6301), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5985) );
  AND2_X2 U7590 ( .A1(n5983), .A2(n5982), .ZN(n6137) );
  NAND2_X1 U7591 ( .A1(n6394), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5984) );
  OAI211_X1 U7592 ( .C1(n6397), .C2(n5986), .A(n5985), .B(n5984), .ZN(n9282)
         );
  INV_X1 U7593 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5989) );
  INV_X2 U7594 ( .A(n6132), .ZN(n6301) );
  NAND2_X1 U7595 ( .A1(n6301), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7596 ( .A1(n6394), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5987) );
  OAI211_X1 U7597 ( .C1(n6397), .C2(n5989), .A(n5988), .B(n5987), .ZN(n9188)
         );
  NAND2_X1 U7598 ( .A1(n9282), .A2(n9188), .ZN(n5990) );
  NAND2_X1 U7599 ( .A1(n9288), .A2(n5990), .ZN(n6500) );
  NAND2_X1 U7600 ( .A1(n5991), .A2(n6386), .ZN(n5993) );
  INV_X4 U7601 ( .A(n6106), .ZN(n6387) );
  NAND2_X1 U7602 ( .A1(n6387), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5992) );
  INV_X1 U7603 ( .A(n9282), .ZN(n5994) );
  OAI21_X1 U7604 ( .B1(n6406), .B2(n6500), .A(n6572), .ZN(n5995) );
  NAND2_X1 U7605 ( .A1(n9517), .A2(n5994), .ZN(n6441) );
  NAND2_X1 U7606 ( .A1(n5995), .A2(n6441), .ZN(n6409) );
  INV_X1 U7607 ( .A(n9188), .ZN(n6438) );
  OR2_X1 U7608 ( .A1(n9288), .A2(n6438), .ZN(n6440) );
  NAND2_X1 U7609 ( .A1(n6440), .A2(n9282), .ZN(n5996) );
  AND2_X1 U7610 ( .A1(n5996), .A2(n9517), .ZN(n6407) );
  INV_X1 U7611 ( .A(n6407), .ZN(n6503) );
  NAND2_X1 U7612 ( .A1(n9022), .A2(n6386), .ZN(n5998) );
  NAND2_X1 U7613 ( .A1(n6387), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5997) );
  NOR2_X2 U7614 ( .A1(n6159), .A2(n6158), .ZN(n6157) );
  OR2_X2 U7615 ( .A1(n6182), .A2(n6181), .ZN(n6184) );
  OR2_X2 U7616 ( .A1(n6184), .A2(n7415), .ZN(n6211) );
  NOR2_X2 U7617 ( .A1(n6211), .A2(n6210), .ZN(n6195) );
  NOR2_X2 U7618 ( .A1(n6235), .A2(n10005), .ZN(n6224) );
  AND2_X2 U7619 ( .A1(n6224), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6251) );
  INV_X1 U7620 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6279) );
  OR2_X2 U7621 ( .A1(n6280), .A2(n6279), .ZN(n6299) );
  INV_X1 U7622 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9131) );
  INV_X1 U7623 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6338) );
  INV_X1 U7624 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9141) );
  NAND2_X1 U7625 ( .A1(n6030), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6033) );
  INV_X1 U7626 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9121) );
  INV_X1 U7627 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9082) );
  NOR2_X2 U7628 ( .A1(n6043), .A2(n9082), .ZN(n6010) );
  AND2_X1 U7629 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5999) );
  NAND2_X1 U7630 ( .A1(n6009), .A2(n5999), .ZN(n8199) );
  OR2_X1 U7631 ( .A1(n8199), .A2(n6393), .ZN(n6006) );
  INV_X1 U7632 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7633 ( .A1(n6394), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7634 ( .A1(n6301), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6001) );
  OAI211_X1 U7635 ( .C1(n6003), .C2(n6397), .A(n6002), .B(n6001), .ZN(n6004)
         );
  INV_X1 U7636 ( .A(n6004), .ZN(n6005) );
  NAND2_X1 U7637 ( .A1(n9527), .A2(n8305), .ZN(n6567) );
  NAND2_X1 U7638 ( .A1(n9032), .A2(n6386), .ZN(n6008) );
  NAND2_X1 U7639 ( .A1(n6387), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6007) );
  INV_X1 U7640 ( .A(n6010), .ZN(n6045) );
  INV_X1 U7641 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7642 ( .A1(n6045), .A2(n6011), .ZN(n6012) );
  NAND2_X1 U7643 ( .A1(n9309), .A2(n6362), .ZN(n6017) );
  INV_X1 U7644 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n10092) );
  NAND2_X1 U7645 ( .A1(n6301), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7646 ( .A1(n6394), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6013) );
  OAI211_X1 U7647 ( .C1(n6397), .C2(n10092), .A(n6014), .B(n6013), .ZN(n6015)
         );
  INV_X1 U7648 ( .A(n6015), .ZN(n6016) );
  NAND2_X1 U7649 ( .A1(n4943), .A2(n9334), .ZN(n8196) );
  NAND2_X1 U7650 ( .A1(n8098), .A2(n6386), .ZN(n6019) );
  NAND2_X1 U7651 ( .A1(n6387), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7652 ( .A1(n6033), .A2(n9121), .ZN(n6020) );
  AND2_X1 U7653 ( .A1(n6043), .A2(n6020), .ZN(n9342) );
  NAND2_X1 U7654 ( .A1(n9342), .A2(n6362), .ZN(n6027) );
  INV_X1 U7655 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7656 ( .A1(n6108), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7657 ( .A1(n6394), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6022) );
  OAI211_X1 U7658 ( .C1(n6132), .C2(n6024), .A(n6023), .B(n6022), .ZN(n6025)
         );
  INV_X1 U7659 ( .A(n6025), .ZN(n6026) );
  AND2_X1 U7660 ( .A1(n9344), .A2(n9362), .ZN(n8220) );
  NAND2_X1 U7661 ( .A1(n8017), .A2(n6386), .ZN(n6029) );
  NAND2_X1 U7662 ( .A1(n6387), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6028) );
  INV_X1 U7663 ( .A(n6030), .ZN(n6351) );
  INV_X1 U7664 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7665 ( .A1(n6351), .A2(n6031), .ZN(n6032) );
  NAND2_X1 U7666 ( .A1(n6033), .A2(n6032), .ZN(n9354) );
  INV_X1 U7667 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7668 ( .A1(n6394), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7669 ( .A1(n6301), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6034) );
  OAI211_X1 U7670 ( .C1(n6397), .C2(n6036), .A(n6035), .B(n6034), .ZN(n6037)
         );
  INV_X1 U7671 ( .A(n6037), .ZN(n6038) );
  INV_X1 U7672 ( .A(n9377), .ZN(n9122) );
  INV_X1 U7673 ( .A(n8219), .ZN(n6040) );
  OR2_X1 U7674 ( .A1(n8220), .A2(n6040), .ZN(n6490) );
  NOR2_X1 U7675 ( .A1(n6490), .A2(n6817), .ZN(n6358) );
  NAND2_X1 U7676 ( .A1(n8158), .A2(n6386), .ZN(n6042) );
  NAND2_X1 U7677 ( .A1(n6387), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7678 ( .A1(n6043), .A2(n9082), .ZN(n6044) );
  NAND2_X1 U7679 ( .A1(n6045), .A2(n6044), .ZN(n9326) );
  INV_X1 U7680 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7681 ( .A1(n6301), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7682 ( .A1(n6394), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6046) );
  OAI211_X1 U7683 ( .C1(n6397), .C2(n6048), .A(n6047), .B(n6046), .ZN(n6049)
         );
  INV_X1 U7684 ( .A(n6049), .ZN(n6050) );
  NAND2_X1 U7685 ( .A1(n6971), .A2(n6386), .ZN(n6058) );
  INV_X1 U7686 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7687 ( .A1(n6052), .A2(n6053), .ZN(n6153) );
  INV_X1 U7688 ( .A(n6165), .ZN(n6055) );
  INV_X1 U7689 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7690 ( .A1(n6055), .A2(n6054), .ZN(n6177) );
  NAND2_X1 U7691 ( .A1(n6206), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6056) );
  AOI22_X1 U7692 ( .A1(n6387), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7276), .B2(
        n7423), .ZN(n6057) );
  NAND2_X1 U7693 ( .A1(n6255), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7694 ( .A1(n6301), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7695 ( .A1(n6184), .A2(n7415), .ZN(n6059) );
  AND2_X1 U7696 ( .A1(n6211), .A2(n6059), .ZN(n7891) );
  NAND2_X1 U7697 ( .A1(n6362), .A2(n7891), .ZN(n6061) );
  NAND2_X1 U7698 ( .A1(n6394), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6060) );
  INV_X1 U7699 ( .A(n6064), .ZN(n6108) );
  NAND2_X1 U7700 ( .A1(n6108), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7701 ( .A1(n6109), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6067) );
  INV_X1 U7702 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7703 ( .A1(n6137), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7704 ( .A1(n6143), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7705 ( .A1(n6108), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7706 ( .A1(n6137), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7707 ( .A1(n6109), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6073) );
  INV_X1 U7708 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7709 ( .A1(n5103), .A2(SI_0_), .ZN(n6077) );
  INV_X1 U7710 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7711 ( .A1(n6077), .A2(n6076), .ZN(n6079) );
  AND2_X1 U7712 ( .A1(n6079), .A2(n6078), .ZN(n9678) );
  MUX2_X1 U7713 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9678), .S(n6124), .Z(n7462) );
  INV_X1 U7714 ( .A(n7462), .ZN(n7701) );
  NAND2_X1 U7715 ( .A1(n6080), .A2(n9724), .ZN(n6081) );
  NAND2_X1 U7716 ( .A1(n6362), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U7717 ( .A1(n6109), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7718 ( .A1(n6137), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7719 ( .A1(n6255), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6082) );
  NAND4_X2 U7720 ( .A1(n6085), .A2(n6084), .A3(n6083), .A4(n6082), .ZN(n9199)
         );
  NAND2_X1 U7721 ( .A1(n6143), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6091) );
  INV_X1 U7722 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7723 ( .A1(n4650), .A2(n6086), .ZN(n6115) );
  NAND2_X1 U7724 ( .A1(n6115), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6088) );
  INV_X1 U7725 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6087) );
  NAND2_X1 U7726 ( .A1(n6088), .A2(n6087), .ZN(n6102) );
  NAND2_X1 U7727 ( .A1(n7276), .A2(n9205), .ZN(n6090) );
  INV_X1 U7728 ( .A(n7136), .ZN(n6421) );
  NAND2_X1 U7729 ( .A1(n7137), .A2(n6421), .ZN(n6094) );
  INV_X1 U7730 ( .A(n9199), .ZN(n7440) );
  INV_X1 U7731 ( .A(n6093), .ZN(n7589) );
  NAND2_X1 U7732 ( .A1(n7440), .A2(n7589), .ZN(n6539) );
  NAND2_X1 U7733 ( .A1(n6109), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U7734 ( .A1(n6255), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6099) );
  INV_X1 U7735 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7736 ( .A1(n6362), .A2(n6095), .ZN(n6098) );
  NAND2_X1 U7737 ( .A1(n6137), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6097) );
  INV_X1 U7738 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6938) );
  INV_X1 U7739 ( .A(n6101), .ZN(n6121) );
  NAND2_X1 U7740 ( .A1(n6121), .A2(n6936), .ZN(n6105) );
  NAND2_X1 U7741 ( .A1(n7276), .A2(n6937), .ZN(n6104) );
  NAND2_X1 U7742 ( .A1(n7670), .A2(n7529), .ZN(n6542) );
  NAND2_X1 U7743 ( .A1(n7530), .A2(n7521), .ZN(n6463) );
  INV_X1 U7744 ( .A(n7533), .ZN(n6422) );
  NAND2_X1 U7745 ( .A1(n6109), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6113) );
  INV_X1 U7746 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6110) );
  XNOR2_X1 U7747 ( .A(n6110), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U7748 ( .A1(n6362), .A2(n7677), .ZN(n6112) );
  NAND2_X1 U7749 ( .A1(n6137), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6111) );
  INV_X1 U7750 ( .A(n6115), .ZN(n6117) );
  NOR2_X1 U7751 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6116) );
  NAND2_X1 U7752 ( .A1(n6117), .A2(n6116), .ZN(n6119) );
  NAND2_X1 U7753 ( .A1(n6119), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6118) );
  MUX2_X1 U7754 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6118), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n6120) );
  NAND2_X1 U7755 ( .A1(n6120), .A2(n6128), .ZN(n7403) );
  NAND2_X1 U7756 ( .A1(n6941), .A2(n6121), .ZN(n6123) );
  NAND2_X1 U7757 ( .A1(n6143), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7758 ( .A1(n7543), .A2(n7667), .ZN(n6467) );
  INV_X1 U7759 ( .A(n6467), .ZN(n6545) );
  NAND2_X2 U7760 ( .A1(n4931), .A2(n9198), .ZN(n7650) );
  NAND3_X1 U7761 ( .A1(n6125), .A2(n6817), .A3(n7650), .ZN(n6126) );
  NAND2_X1 U7762 ( .A1(n6127), .A2(n6126), .ZN(n6141) );
  NAND2_X1 U7763 ( .A1(n6943), .A2(n6121), .ZN(n6131) );
  NAND2_X1 U7764 ( .A1(n6128), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6129) );
  XNOR2_X1 U7765 ( .A(n6129), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6946) );
  AOI22_X1 U7766 ( .A1(n6143), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7276), .B2(
        n6946), .ZN(n6130) );
  NAND2_X1 U7767 ( .A1(n6255), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6140) );
  INV_X1 U7768 ( .A(n6133), .ZN(n6147) );
  INV_X1 U7769 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7770 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6134) );
  NAND2_X1 U7771 ( .A1(n6135), .A2(n6134), .ZN(n6136) );
  AND2_X1 U7772 ( .A1(n6147), .A2(n6136), .ZN(n7545) );
  NAND2_X1 U7773 ( .A1(n6362), .A2(n7545), .ZN(n6139) );
  NAND2_X1 U7774 ( .A1(n6137), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7775 ( .A1(n9781), .A2(n9197), .ZN(n6460) );
  NAND2_X1 U7776 ( .A1(n7740), .A2(n7602), .ZN(n7734) );
  NAND2_X1 U7777 ( .A1(n6460), .A2(n7650), .ZN(n6466) );
  NAND2_X1 U7778 ( .A1(n6949), .A2(n6386), .ZN(n6145) );
  OR2_X1 U7779 ( .A1(n6052), .A2(n9659), .ZN(n6142) );
  XNOR2_X1 U7780 ( .A(n6142), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9217) );
  AOI22_X1 U7781 ( .A1(n6387), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7276), .B2(
        n9217), .ZN(n6144) );
  INV_X1 U7782 ( .A(n9788), .ZN(n7605) );
  NAND2_X1 U7783 ( .A1(n6301), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6152) );
  INV_X1 U7784 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7785 ( .A1(n6147), .A2(n6146), .ZN(n6148) );
  AND2_X1 U7786 ( .A1(n6159), .A2(n6148), .ZN(n7866) );
  NAND2_X1 U7787 ( .A1(n6362), .A2(n7866), .ZN(n6150) );
  NAND2_X1 U7788 ( .A1(n6394), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7789 ( .A1(n6953), .A2(n6386), .ZN(n6156) );
  NAND2_X1 U7790 ( .A1(n6153), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6154) );
  XNOR2_X1 U7791 ( .A(n6154), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6916) );
  AOI22_X1 U7792 ( .A1(n6387), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7276), .B2(
        n6916), .ZN(n6155) );
  NAND2_X1 U7793 ( .A1(n6255), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7794 ( .A1(n6301), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6163) );
  INV_X1 U7795 ( .A(n6157), .ZN(n6170) );
  NAND2_X1 U7796 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  AND2_X1 U7797 ( .A1(n6170), .A2(n6160), .ZN(n7684) );
  NAND2_X1 U7798 ( .A1(n6362), .A2(n7684), .ZN(n6162) );
  NAND2_X1 U7799 ( .A1(n6394), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7800 ( .A1(n7791), .A2(n7910), .ZN(n7800) );
  OR2_X1 U7801 ( .A1(n7791), .A2(n7910), .ZN(n6420) );
  NAND2_X1 U7802 ( .A1(n6964), .A2(n6386), .ZN(n6169) );
  NAND2_X1 U7803 ( .A1(n6165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6166) );
  MUX2_X1 U7804 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6166), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n6167) );
  NAND2_X1 U7805 ( .A1(n6167), .A2(n6177), .ZN(n6966) );
  INV_X1 U7806 ( .A(n6966), .ZN(n7178) );
  AOI22_X1 U7807 ( .A1(n6387), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7276), .B2(
        n7178), .ZN(n6168) );
  NAND2_X1 U7808 ( .A1(n6255), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7809 ( .A1(n6301), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6174) );
  INV_X1 U7810 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7180) );
  NAND2_X1 U7811 ( .A1(n6170), .A2(n7180), .ZN(n6171) );
  AND2_X1 U7812 ( .A1(n6182), .A2(n6171), .ZN(n7935) );
  NAND2_X1 U7813 ( .A1(n6362), .A2(n7935), .ZN(n6173) );
  NAND2_X1 U7814 ( .A1(n6394), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6172) );
  OR2_X1 U7815 ( .A1(n7936), .A2(n7688), .ZN(n7815) );
  NAND3_X1 U7816 ( .A1(n6176), .A2(n6420), .A3(n7815), .ZN(n6189) );
  NAND2_X1 U7817 ( .A1(n7936), .A2(n7688), .ZN(n7803) );
  NAND2_X1 U7818 ( .A1(n6969), .A2(n6386), .ZN(n6180) );
  NAND2_X1 U7819 ( .A1(n6177), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6178) );
  XNOR2_X1 U7820 ( .A(n6178), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7433) );
  AOI22_X1 U7821 ( .A1(n6387), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7276), .B2(
        n7433), .ZN(n6179) );
  NAND2_X1 U7822 ( .A1(n6301), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7823 ( .A1(n6182), .A2(n6181), .ZN(n6183) );
  AND2_X1 U7824 ( .A1(n6184), .A2(n6183), .ZN(n7955) );
  NAND2_X1 U7825 ( .A1(n6362), .A2(n7955), .ZN(n6186) );
  NAND2_X1 U7826 ( .A1(n6394), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6185) );
  NAND4_X1 U7827 ( .A1(n6188), .A2(n6187), .A3(n6186), .A4(n6185), .ZN(n9193)
         );
  INV_X1 U7828 ( .A(n9193), .ZN(n7880) );
  NAND2_X1 U7829 ( .A1(n9625), .A2(n7880), .ZN(n7886) );
  NAND3_X1 U7830 ( .A1(n6189), .A2(n7803), .A3(n7886), .ZN(n6190) );
  OR2_X1 U7831 ( .A1(n9625), .A2(n7880), .ZN(n6419) );
  NAND3_X1 U7832 ( .A1(n6190), .A2(n7966), .A3(n6419), .ZN(n6202) );
  NAND2_X1 U7833 ( .A1(n6990), .A2(n6386), .ZN(n6194) );
  NAND2_X1 U7834 ( .A1(n6191), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6192) );
  XNOR2_X1 U7835 ( .A(n6192), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7556) );
  AOI22_X1 U7836 ( .A1(n6387), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7276), .B2(
        n7556), .ZN(n6193) );
  NAND2_X1 U7837 ( .A1(n6301), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7838 ( .A1(n6394), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6200) );
  INV_X1 U7839 ( .A(n6195), .ZN(n6213) );
  INV_X1 U7840 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7841 ( .A1(n6213), .A2(n6196), .ZN(n6197) );
  AND2_X1 U7842 ( .A1(n6233), .A2(n6197), .ZN(n8131) );
  NAND2_X1 U7843 ( .A1(n6362), .A2(n8131), .ZN(n6199) );
  NAND2_X1 U7844 ( .A1(n9615), .A2(n8136), .ZN(n8143) );
  NAND2_X1 U7845 ( .A1(n9620), .A2(n7969), .ZN(n6418) );
  AND2_X1 U7846 ( .A1(n6420), .A2(n7611), .ZN(n6469) );
  NAND2_X1 U7847 ( .A1(n7803), .A2(n7800), .ZN(n6454) );
  AOI21_X1 U7848 ( .B1(n6203), .B2(n6469), .A(n6454), .ZN(n6205) );
  AND2_X1 U7849 ( .A1(n6419), .A2(n7815), .ZN(n7884) );
  INV_X1 U7850 ( .A(n7884), .ZN(n6204) );
  AND2_X1 U7851 ( .A1(n6418), .A2(n7886), .ZN(n7964) );
  OAI211_X1 U7852 ( .C1(n6205), .C2(n6204), .A(n6406), .B(n7964), .ZN(n6218)
         );
  NAND2_X1 U7853 ( .A1(n6978), .A2(n6386), .ZN(n6209) );
  OAI21_X1 U7854 ( .B1(n6206), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6207) );
  XNOR2_X1 U7855 ( .A(n6207), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7296) );
  AOI22_X1 U7856 ( .A1(n6387), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7296), .B2(
        n7276), .ZN(n6208) );
  NAND2_X1 U7857 ( .A1(n6301), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7858 ( .A1(n6394), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7859 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  AND2_X1 U7860 ( .A1(n6213), .A2(n6212), .ZN(n8014) );
  NAND2_X1 U7861 ( .A1(n6362), .A2(n8014), .ZN(n6215) );
  NAND2_X1 U7862 ( .A1(n6255), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6214) );
  NAND4_X1 U7863 ( .A1(n6217), .A2(n6216), .A3(n6215), .A4(n6214), .ZN(n9191)
         );
  INV_X1 U7864 ( .A(n9191), .ZN(n8041) );
  XNOR2_X1 U7865 ( .A(n8057), .B(n8041), .ZN(n7963) );
  NAND2_X1 U7866 ( .A1(n8042), .A2(n8041), .ZN(n8037) );
  NAND2_X1 U7867 ( .A1(n8143), .A2(n8037), .ZN(n6456) );
  AND2_X1 U7868 ( .A1(n6456), .A2(n6417), .ZN(n6241) );
  NAND2_X1 U7869 ( .A1(n6997), .A2(n6386), .ZN(n6221) );
  OR2_X1 U7870 ( .A1(n6219), .A2(n9659), .ZN(n6245) );
  XNOR2_X1 U7871 ( .A(n6245), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9234) );
  AOI22_X1 U7872 ( .A1(n6387), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7276), .B2(
        n9234), .ZN(n6220) );
  INV_X1 U7873 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U7874 ( .A1(n6301), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7875 ( .A1(n6255), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6222) );
  AND2_X1 U7876 ( .A1(n6223), .A2(n6222), .ZN(n6227) );
  INV_X1 U7877 ( .A(n6224), .ZN(n6253) );
  NAND2_X1 U7878 ( .A1(n6235), .A2(n10005), .ZN(n6225) );
  NAND2_X1 U7879 ( .A1(n6253), .A2(n6225), .ZN(n9052) );
  OR2_X1 U7880 ( .A1(n9052), .A2(n6393), .ZN(n6226) );
  OAI211_X1 U7881 ( .C1(n6096), .C2(n10015), .A(n6227), .B(n6226), .ZN(n9511)
         );
  NAND2_X1 U7882 ( .A1(n9606), .A2(n9476), .ZN(n6416) );
  NAND2_X1 U7883 ( .A1(n6416), .A2(n6406), .ZN(n6243) );
  NAND2_X1 U7884 ( .A1(n6992), .A2(n6386), .ZN(n6231) );
  NAND2_X1 U7885 ( .A1(n6228), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6229) );
  XNOR2_X1 U7886 ( .A(n6229), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7713) );
  AOI22_X1 U7887 ( .A1(n6387), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7276), .B2(
        n7713), .ZN(n6230) );
  NAND2_X1 U7888 ( .A1(n6255), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7889 ( .A1(n6301), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7890 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  AND2_X1 U7891 ( .A1(n6235), .A2(n6234), .ZN(n9500) );
  NAND2_X1 U7892 ( .A1(n6362), .A2(n9500), .ZN(n6237) );
  NAND2_X1 U7893 ( .A1(n6394), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6236) );
  NAND4_X1 U7894 ( .A1(n6239), .A2(n6238), .A3(n6237), .A4(n6236), .ZN(n9190)
         );
  NAND2_X1 U7895 ( .A1(n9610), .A2(n9049), .ZN(n8144) );
  INV_X1 U7896 ( .A(n8144), .ZN(n6240) );
  OR3_X1 U7897 ( .A1(n6241), .A2(n6243), .A3(n6240), .ZN(n6261) );
  OR2_X1 U7898 ( .A1(n8042), .A2(n8041), .ZN(n8039) );
  AND2_X1 U7899 ( .A1(n6417), .A2(n8039), .ZN(n8141) );
  OR2_X1 U7900 ( .A1(n9610), .A2(n9049), .ZN(n6415) );
  OAI21_X1 U7901 ( .B1(n8141), .B2(n4707), .A(n6415), .ZN(n6479) );
  AND2_X1 U7902 ( .A1(n6416), .A2(n8144), .ZN(n6480) );
  NAND3_X1 U7903 ( .A1(n6242), .A2(n6817), .A3(n8203), .ZN(n6260) );
  AOI21_X1 U7904 ( .B1(n8203), .B2(n6415), .A(n6243), .ZN(n6258) );
  NAND2_X1 U7905 ( .A1(n7125), .A2(n6386), .ZN(n6250) );
  NAND2_X1 U7906 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  NAND2_X1 U7907 ( .A1(n6246), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6248) );
  INV_X1 U7908 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6247) );
  XNOR2_X1 U7909 ( .A(n6248), .B(n6247), .ZN(n7126) );
  INV_X1 U7910 ( .A(n7126), .ZN(n9245) );
  AOI22_X1 U7911 ( .A1(n9245), .A2(n7276), .B1(n6387), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n6249) );
  INV_X1 U7912 ( .A(n6251), .ZN(n6268) );
  INV_X1 U7913 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7914 ( .A1(n6253), .A2(n6252), .ZN(n6254) );
  NAND2_X1 U7915 ( .A1(n6268), .A2(n6254), .ZN(n9487) );
  AOI22_X1 U7916 ( .A1(n6255), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n6301), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7917 ( .A1(n6394), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6256) );
  OAI211_X1 U7918 ( .C1(n9487), .C2(n6393), .A(n6257), .B(n6256), .ZN(n9458)
         );
  INV_X1 U7919 ( .A(n9458), .ZN(n6688) );
  NAND2_X1 U7920 ( .A1(n9599), .A2(n6688), .ZN(n8205) );
  NAND2_X1 U7921 ( .A1(n9455), .A2(n8205), .ZN(n9479) );
  NOR2_X1 U7922 ( .A1(n6258), .A2(n9479), .ZN(n6259) );
  OAI211_X1 U7923 ( .C1(n6262), .C2(n6261), .A(n6260), .B(n6259), .ZN(n6276)
         );
  NAND2_X1 U7924 ( .A1(n7286), .A2(n6386), .ZN(n6266) );
  NAND2_X1 U7925 ( .A1(n6263), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6264) );
  XNOR2_X1 U7926 ( .A(n6264), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7288) );
  AOI22_X1 U7927 ( .A1(n6387), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7276), .B2(
        n7288), .ZN(n6265) );
  INV_X1 U7928 ( .A(n9595), .ZN(n6273) );
  INV_X1 U7929 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6272) );
  INV_X1 U7930 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U7931 ( .A1(n6268), .A2(n6267), .ZN(n6269) );
  NAND2_X1 U7932 ( .A1(n6280), .A2(n6269), .ZN(n9465) );
  OR2_X1 U7933 ( .A1(n9465), .A2(n6393), .ZN(n6271) );
  AOI22_X1 U7934 ( .A1(n6255), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n6301), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6270) );
  OAI211_X1 U7935 ( .C1(n6096), .C2(n6272), .A(n6271), .B(n6270), .ZN(n9448)
         );
  NAND2_X1 U7936 ( .A1(n6273), .A2(n9448), .ZN(n6474) );
  INV_X1 U7937 ( .A(n9448), .ZN(n9475) );
  NAND2_X1 U7938 ( .A1(n9595), .A2(n9475), .ZN(n8207) );
  NAND2_X1 U7939 ( .A1(n6474), .A2(n8207), .ZN(n9467) );
  INV_X1 U7940 ( .A(n9467), .ZN(n6275) );
  MUX2_X1 U7941 ( .A(n8205), .B(n9455), .S(n6817), .Z(n6274) );
  NAND3_X1 U7942 ( .A1(n6276), .A2(n6275), .A3(n6274), .ZN(n6290) );
  NAND2_X1 U7943 ( .A1(n7341), .A2(n6386), .ZN(n6278) );
  NAND2_X1 U7944 ( .A1(n4332), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6292) );
  XNOR2_X1 U7945 ( .A(n6292), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9272) );
  AOI22_X1 U7946 ( .A1(n7276), .A2(n9272), .B1(n6387), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7947 ( .A1(n6280), .A2(n6279), .ZN(n6281) );
  AND2_X1 U7948 ( .A1(n6299), .A2(n6281), .ZN(n9443) );
  NAND2_X1 U7949 ( .A1(n9443), .A2(n6362), .ZN(n6287) );
  INV_X1 U7950 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U7951 ( .A1(n6301), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U7952 ( .A1(n6394), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6282) );
  OAI211_X1 U7953 ( .C1(n6397), .C2(n6284), .A(n6283), .B(n6282), .ZN(n6285)
         );
  INV_X1 U7954 ( .A(n6285), .ZN(n6286) );
  NAND2_X1 U7955 ( .A1(n6287), .A2(n6286), .ZN(n9457) );
  INV_X1 U7956 ( .A(n9457), .ZN(n6288) );
  OR2_X1 U7957 ( .A1(n9589), .A2(n6288), .ZN(n9432) );
  MUX2_X1 U7958 ( .A(n6474), .B(n8207), .S(n6817), .Z(n6289) );
  NAND3_X1 U7959 ( .A1(n6290), .A2(n9447), .A3(n6289), .ZN(n6308) );
  NAND2_X1 U7960 ( .A1(n7514), .A2(n6386), .ZN(n6296) );
  NAND2_X1 U7961 ( .A1(n6292), .A2(n6291), .ZN(n6293) );
  NAND2_X1 U7962 ( .A1(n6293), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6294) );
  XNOR2_X1 U7963 ( .A(n6294), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9710) );
  AOI22_X1 U7964 ( .A1(n9710), .A2(n7276), .B1(n6387), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n6295) );
  INV_X1 U7965 ( .A(n6297), .ZN(n6312) );
  NAND2_X1 U7966 ( .A1(n6299), .A2(n6298), .ZN(n6300) );
  NAND2_X1 U7967 ( .A1(n6312), .A2(n6300), .ZN(n9428) );
  OR2_X1 U7968 ( .A1(n9428), .A2(n6393), .ZN(n6306) );
  INV_X1 U7969 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U7970 ( .A1(n6394), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7971 ( .A1(n6301), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6302) );
  OAI211_X1 U7972 ( .C1(n6397), .C2(n9270), .A(n6303), .B(n6302), .ZN(n6304)
         );
  INV_X1 U7973 ( .A(n6304), .ZN(n6305) );
  AND2_X1 U7974 ( .A1(n6414), .A2(n9432), .ZN(n8209) );
  NAND2_X1 U7975 ( .A1(n9584), .A2(n6720), .ZN(n8210) );
  AND2_X1 U7976 ( .A1(n8210), .A2(n4966), .ZN(n6453) );
  MUX2_X1 U7977 ( .A(n8209), .B(n6453), .S(n6406), .Z(n6307) );
  NAND2_X1 U7978 ( .A1(n6308), .A2(n6307), .ZN(n6332) );
  NAND2_X1 U7979 ( .A1(n7640), .A2(n6386), .ZN(n6310) );
  AOI22_X1 U7980 ( .A1(n9278), .A2(n7276), .B1(n6387), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n6309) );
  INV_X1 U7981 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7982 ( .A1(n6312), .A2(n6311), .ZN(n6313) );
  NAND2_X1 U7983 ( .A1(n6322), .A2(n6313), .ZN(n9414) );
  OR2_X1 U7984 ( .A1(n9414), .A2(n6393), .ZN(n6319) );
  INV_X1 U7985 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U7986 ( .A1(n6394), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6315) );
  NAND2_X1 U7987 ( .A1(n6301), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6314) );
  OAI211_X1 U7988 ( .C1(n6397), .C2(n6316), .A(n6315), .B(n6314), .ZN(n6317)
         );
  INV_X1 U7989 ( .A(n6317), .ZN(n6318) );
  NAND2_X1 U7990 ( .A1(n6319), .A2(n6318), .ZN(n9436) );
  INV_X1 U7991 ( .A(n9436), .ZN(n9153) );
  OR2_X1 U7992 ( .A1(n9580), .A2(n9153), .ZN(n6447) );
  NAND3_X1 U7993 ( .A1(n6332), .A2(n6414), .A3(n6447), .ZN(n6330) );
  NAND2_X1 U7994 ( .A1(n7730), .A2(n6386), .ZN(n6321) );
  NAND2_X1 U7995 ( .A1(n6387), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6320) );
  NAND2_X1 U7996 ( .A1(n6322), .A2(n9131), .ZN(n6323) );
  NAND2_X1 U7997 ( .A1(n6339), .A2(n6323), .ZN(n9401) );
  OR2_X1 U7998 ( .A1(n9401), .A2(n6393), .ZN(n6328) );
  INV_X1 U7999 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10050) );
  NAND2_X1 U8000 ( .A1(n6301), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U8001 ( .A1(n6394), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6324) );
  OAI211_X1 U8002 ( .C1(n6397), .C2(n10050), .A(n6325), .B(n6324), .ZN(n6326)
         );
  INV_X1 U8003 ( .A(n6326), .ZN(n6327) );
  NAND2_X1 U8004 ( .A1(n6328), .A2(n6327), .ZN(n9420) );
  INV_X1 U8005 ( .A(n9420), .ZN(n6731) );
  NOR2_X1 U8006 ( .A1(n8214), .A2(n6817), .ZN(n6329) );
  NAND2_X1 U8007 ( .A1(n6330), .A2(n6329), .ZN(n6333) );
  NAND2_X1 U8008 ( .A1(n9580), .A2(n9153), .ZN(n8212) );
  NAND2_X1 U8009 ( .A1(n6447), .A2(n6817), .ZN(n6331) );
  OAI22_X1 U8010 ( .A1(n6333), .A2(n4725), .B1(n8215), .B2(n6331), .ZN(n6335)
         );
  AND2_X1 U8011 ( .A1(n8212), .A2(n8210), .ZN(n6444) );
  NAND3_X1 U8012 ( .A1(n6333), .A2(n6444), .A3(n6332), .ZN(n6334) );
  NAND2_X1 U8013 ( .A1(n6335), .A2(n6334), .ZN(n6370) );
  INV_X1 U8014 ( .A(n8215), .ZN(n9387) );
  NAND2_X1 U8015 ( .A1(n7853), .A2(n6386), .ZN(n6337) );
  NAND2_X1 U8016 ( .A1(n6387), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U8017 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  AND2_X1 U8018 ( .A1(n6349), .A2(n6340), .ZN(n9384) );
  NAND2_X1 U8019 ( .A1(n9384), .A2(n6362), .ZN(n6345) );
  INV_X1 U8020 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9999) );
  NAND2_X1 U8021 ( .A1(n6394), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U8022 ( .A1(n6301), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6341) );
  OAI211_X1 U8023 ( .C1(n6397), .C2(n9999), .A(n6342), .B(n6341), .ZN(n6343)
         );
  INV_X1 U8024 ( .A(n6343), .ZN(n6344) );
  NAND2_X1 U8025 ( .A1(n9570), .A2(n9142), .ZN(n8217) );
  INV_X1 U8026 ( .A(n8217), .ZN(n6346) );
  NAND2_X1 U8027 ( .A1(n7980), .A2(n6386), .ZN(n6348) );
  NAND2_X1 U8028 ( .A1(n6387), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U8029 ( .A1(n6349), .A2(n9141), .ZN(n6350) );
  NAND2_X1 U8030 ( .A1(n6351), .A2(n6350), .ZN(n9370) );
  INV_X1 U8031 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n10076) );
  NAND2_X1 U8032 ( .A1(n6301), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U8033 ( .A1(n6394), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6352) );
  OAI211_X1 U8034 ( .C1(n10076), .C2(n6397), .A(n6353), .B(n6352), .ZN(n6354)
         );
  INV_X1 U8035 ( .A(n6354), .ZN(n6355) );
  NAND2_X1 U8036 ( .A1(n6356), .A2(n6355), .ZN(n9392) );
  INV_X1 U8037 ( .A(n9392), .ZN(n9076) );
  OR2_X1 U8038 ( .A1(n9564), .A2(n9076), .ZN(n6449) );
  NAND2_X1 U8039 ( .A1(n6449), .A2(n6448), .ZN(n6357) );
  NAND2_X1 U8040 ( .A1(n9564), .A2(n9076), .ZN(n9358) );
  NAND3_X1 U8041 ( .A1(n9311), .A2(n6817), .A3(n9334), .ZN(n6359) );
  NAND2_X1 U8042 ( .A1(n9029), .A2(n6386), .ZN(n6361) );
  NAND2_X1 U8043 ( .A1(n6387), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6360) );
  XNOR2_X1 U8044 ( .A(n6391), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9301) );
  NAND2_X1 U8045 ( .A1(n9301), .A2(n6362), .ZN(n6368) );
  INV_X1 U8046 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n6365) );
  NAND2_X1 U8047 ( .A1(n6394), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U8048 ( .A1(n6301), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6363) );
  OAI211_X1 U8049 ( .C1(n6397), .C2(n6365), .A(n6364), .B(n6363), .ZN(n6366)
         );
  INV_X1 U8050 ( .A(n6366), .ZN(n6367) );
  NAND2_X1 U8051 ( .A1(n9543), .A2(n8306), .ZN(n6412) );
  INV_X1 U8052 ( .A(n9334), .ZN(n6862) );
  NAND2_X1 U8053 ( .A1(n4943), .A2(n6862), .ZN(n8222) );
  NAND2_X1 U8054 ( .A1(n6412), .A2(n8222), .ZN(n6369) );
  NAND2_X1 U8055 ( .A1(n6369), .A2(n6406), .ZN(n6385) );
  INV_X1 U8056 ( .A(n6449), .ZN(n6376) );
  INV_X1 U8057 ( .A(n6370), .ZN(n6373) );
  NAND2_X1 U8058 ( .A1(n6448), .A2(n8214), .ZN(n6371) );
  AND2_X1 U8059 ( .A1(n6371), .A2(n8217), .ZN(n6372) );
  NAND2_X1 U8060 ( .A1(n6372), .A2(n9358), .ZN(n6452) );
  AOI21_X1 U8061 ( .B1(n6373), .B2(n6448), .A(n6452), .ZN(n6375) );
  NAND2_X1 U8062 ( .A1(n9550), .A2(n9169), .ZN(n6413) );
  NAND2_X1 U8063 ( .A1(n9559), .A2(n9122), .ZN(n6489) );
  INV_X1 U8064 ( .A(n9362), .ZN(n9083) );
  NAND2_X1 U8065 ( .A1(n4942), .A2(n9083), .ZN(n9330) );
  AND4_X1 U8066 ( .A1(n6413), .A2(n6817), .A3(n6489), .A4(n9330), .ZN(n6374)
         );
  OAI211_X1 U8067 ( .C1(n6376), .C2(n6375), .A(n9315), .B(n6374), .ZN(n6384)
         );
  AND2_X1 U8068 ( .A1(n6413), .A2(n9330), .ZN(n8221) );
  OAI21_X1 U8069 ( .B1(n8220), .B2(n6489), .A(n8221), .ZN(n6377) );
  NAND3_X1 U8070 ( .A1(n6377), .A2(n6406), .A3(n9312), .ZN(n6382) );
  INV_X1 U8071 ( .A(n9330), .ZN(n6379) );
  INV_X1 U8072 ( .A(n8220), .ZN(n6378) );
  OAI211_X1 U8073 ( .C1(n6379), .C2(n8219), .A(n6378), .B(n9312), .ZN(n6380)
         );
  NAND3_X1 U8074 ( .A1(n6380), .A2(n6817), .A3(n6413), .ZN(n6381) );
  NAND2_X1 U8075 ( .A1(n6382), .A2(n6381), .ZN(n6383) );
  INV_X1 U8076 ( .A(n8225), .ZN(n6402) );
  NAND2_X1 U8077 ( .A1(n9025), .A2(n6386), .ZN(n6389) );
  NAND2_X1 U8078 ( .A1(n6387), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6388) );
  INV_X1 U8079 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6861) );
  INV_X1 U8080 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6390) );
  OAI21_X1 U8081 ( .B1(n6391), .B2(n6861), .A(n6390), .ZN(n6392) );
  NAND2_X1 U8082 ( .A1(n6392), .A2(n8199), .ZN(n6823) );
  INV_X1 U8083 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U8084 ( .A1(n6301), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U8085 ( .A1(n6394), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6395) );
  OAI211_X1 U8086 ( .C1(n6398), .C2(n6397), .A(n6396), .B(n6395), .ZN(n6399)
         );
  INV_X1 U8087 ( .A(n6399), .ZN(n6400) );
  NAND2_X2 U8088 ( .A1(n6401), .A2(n6400), .ZN(n9297) );
  NAND2_X1 U8089 ( .A1(n9536), .A2(n6863), .ZN(n8227) );
  AND2_X1 U8090 ( .A1(n8227), .A2(n6412), .ZN(n6495) );
  OAI21_X1 U8091 ( .B1(n6404), .B2(n6402), .A(n6495), .ZN(n6403) );
  NAND3_X1 U8092 ( .A1(n6404), .A2(n8226), .A3(n8225), .ZN(n6405) );
  NAND2_X1 U8093 ( .A1(n6407), .A2(n6406), .ZN(n6408) );
  XNOR2_X1 U8094 ( .A(n9344), .B(n9362), .ZN(n9346) );
  INV_X1 U8095 ( .A(n9434), .ZN(n6431) );
  INV_X1 U8096 ( .A(n9479), .ZN(n6428) );
  NAND2_X1 U8097 ( .A1(n6417), .A2(n8143), .ZN(n8134) );
  INV_X1 U8098 ( .A(n7963), .ZN(n7968) );
  NAND2_X1 U8099 ( .A1(n7966), .A2(n6418), .ZN(n7959) );
  NAND2_X1 U8100 ( .A1(n6419), .A2(n7886), .ZN(n7819) );
  AND2_X1 U8101 ( .A1(n9201), .A2(n7701), .ZN(n6537) );
  NOR2_X1 U8102 ( .A1(n7268), .A2(n6537), .ZN(n7456) );
  NAND4_X1 U8103 ( .A1(n7456), .A2(n6422), .A3(n7267), .A4(n6421), .ZN(n6423)
         );
  NAND2_X1 U8104 ( .A1(n7734), .A2(n6460), .ZN(n7540) );
  NAND2_X2 U8105 ( .A1(n7650), .A2(n6467), .ZN(n7651) );
  NOR3_X1 U8106 ( .A1(n6423), .A2(n7540), .A3(n7651), .ZN(n6424) );
  NAND4_X1 U8107 ( .A1(n7804), .A2(n4716), .A3(n4279), .A4(n6424), .ZN(n6425)
         );
  OR3_X1 U8108 ( .A1(n7959), .A2(n7819), .A3(n6425), .ZN(n6426) );
  NOR3_X1 U8109 ( .A1(n8134), .A2(n7968), .A3(n6426), .ZN(n6427) );
  NAND4_X1 U8110 ( .A1(n6428), .A2(n9504), .A3(n8146), .A4(n6427), .ZN(n6429)
         );
  NOR2_X1 U8111 ( .A1(n9467), .A2(n6429), .ZN(n6430) );
  NAND4_X1 U8112 ( .A1(n9418), .A2(n6431), .A3(n9447), .A4(n6430), .ZN(n6432)
         );
  NOR2_X1 U8113 ( .A1(n9405), .A2(n6432), .ZN(n6433) );
  NAND3_X1 U8114 ( .A1(n9376), .A2(n9390), .A3(n6433), .ZN(n6434) );
  NAND2_X1 U8115 ( .A1(n8219), .A2(n6489), .ZN(n9360) );
  OR2_X1 U8116 ( .A1(n6434), .A2(n9360), .ZN(n6435) );
  NOR3_X1 U8117 ( .A1(n9333), .A2(n9346), .A3(n6435), .ZN(n6436) );
  NAND3_X1 U8118 ( .A1(n9296), .A2(n6436), .A3(n9315), .ZN(n6437) );
  NOR2_X1 U8119 ( .A1(n8302), .A2(n6437), .ZN(n6439) );
  NAND2_X1 U8120 ( .A1(n9288), .A2(n6438), .ZN(n6568) );
  NAND4_X1 U8121 ( .A1(n6572), .A2(n9532), .A3(n6439), .A4(n6568), .ZN(n6442)
         );
  NAND2_X1 U8122 ( .A1(n6441), .A2(n6440), .ZN(n6573) );
  OR2_X1 U8123 ( .A1(n6442), .A2(n6573), .ZN(n6443) );
  NAND2_X1 U8124 ( .A1(n6443), .A2(n7854), .ZN(n6531) );
  INV_X1 U8125 ( .A(n6444), .ZN(n6445) );
  OR2_X1 U8126 ( .A1(n6445), .A2(n8209), .ZN(n6446) );
  AND4_X1 U8127 ( .A1(n9387), .A2(n6448), .A3(n6447), .A4(n6446), .ZN(n6450)
         );
  OAI21_X1 U8128 ( .B1(n6452), .B2(n6450), .A(n6449), .ZN(n6451) );
  NOR2_X1 U8129 ( .A1(n6490), .A2(n6451), .ZN(n6558) );
  NOR2_X1 U8130 ( .A1(n6452), .A2(n4725), .ZN(n6534) );
  INV_X1 U8131 ( .A(n6453), .ZN(n6459) );
  INV_X1 U8132 ( .A(n6454), .ZN(n6457) );
  NOR2_X1 U8133 ( .A1(n7964), .A2(n4705), .ZN(n6455) );
  NOR2_X1 U8134 ( .A1(n6456), .A2(n6455), .ZN(n6475) );
  NAND4_X1 U8135 ( .A1(n8205), .A2(n6480), .A3(n6457), .A4(n6475), .ZN(n6458)
         );
  OR3_X1 U8136 ( .A1(n6459), .A2(n4720), .A3(n6458), .ZN(n6535) );
  INV_X1 U8137 ( .A(n6469), .ZN(n6546) );
  INV_X1 U8138 ( .A(n6460), .ZN(n6461) );
  NAND2_X1 U8139 ( .A1(n6468), .A2(n6461), .ZN(n7612) );
  INV_X1 U8140 ( .A(n7612), .ZN(n6462) );
  NOR2_X1 U8141 ( .A1(n6546), .A2(n6462), .ZN(n6544) );
  AND2_X1 U8142 ( .A1(n7650), .A2(n6463), .ZN(n6464) );
  NAND2_X1 U8143 ( .A1(n6544), .A2(n6464), .ZN(n6536) );
  INV_X1 U8144 ( .A(n7441), .ZN(n6473) );
  AOI21_X1 U8145 ( .B1(n6467), .B2(n6542), .A(n6466), .ZN(n6471) );
  AND2_X1 U8146 ( .A1(n6468), .A2(n7734), .ZN(n7609) );
  INV_X1 U8147 ( .A(n7609), .ZN(n6470) );
  OAI21_X1 U8148 ( .B1(n6471), .B2(n6470), .A(n6469), .ZN(n6472) );
  OAI21_X1 U8149 ( .B1(n6536), .B2(n6473), .A(n6472), .ZN(n6486) );
  AND2_X1 U8150 ( .A1(n6474), .A2(n9455), .ZN(n8206) );
  INV_X1 U8151 ( .A(n6475), .ZN(n6477) );
  AND2_X1 U8152 ( .A1(n7884), .A2(n7966), .ZN(n6476) );
  NOR2_X1 U8153 ( .A1(n6477), .A2(n6476), .ZN(n6478) );
  NOR2_X1 U8154 ( .A1(n6479), .A2(n6478), .ZN(n6482) );
  INV_X1 U8155 ( .A(n6480), .ZN(n6481) );
  OAI21_X1 U8156 ( .B1(n6482), .B2(n6481), .A(n8203), .ZN(n6483) );
  NAND2_X1 U8157 ( .A1(n6483), .A2(n8205), .ZN(n6484) );
  AOI21_X1 U8158 ( .B1(n8206), .B2(n6484), .A(n4720), .ZN(n6485) );
  NAND3_X1 U8159 ( .A1(n8210), .A2(n6485), .A3(n4966), .ZN(n6552) );
  OAI21_X1 U8160 ( .B1(n6535), .B2(n6486), .A(n6552), .ZN(n6487) );
  NAND2_X1 U8161 ( .A1(n6534), .A2(n6487), .ZN(n6488) );
  NAND2_X1 U8162 ( .A1(n6558), .A2(n6488), .ZN(n6492) );
  OR2_X1 U8163 ( .A1(n6490), .A2(n6489), .ZN(n6491) );
  AND2_X1 U8164 ( .A1(n8221), .A2(n6491), .ZN(n6559) );
  NAND2_X1 U8165 ( .A1(n6492), .A2(n6559), .ZN(n6494) );
  OR2_X1 U8166 ( .A1(n4943), .A2(n6862), .ZN(n6493) );
  AND2_X1 U8167 ( .A1(n6493), .A2(n9312), .ZN(n8224) );
  AND3_X1 U8168 ( .A1(n6494), .A2(n8224), .A3(n8225), .ZN(n6499) );
  AND2_X1 U8169 ( .A1(n8225), .A2(n8223), .ZN(n6497) );
  INV_X1 U8170 ( .A(n6495), .ZN(n6496) );
  OR2_X1 U8171 ( .A1(n6497), .A2(n6496), .ZN(n6533) );
  AND2_X1 U8172 ( .A1(n6498), .A2(n8226), .ZN(n6563) );
  OAI21_X1 U8173 ( .B1(n6499), .B2(n6533), .A(n6563), .ZN(n6501) );
  NAND3_X1 U8174 ( .A1(n6501), .A2(n6567), .A3(n6500), .ZN(n6502) );
  NAND2_X1 U8175 ( .A1(n6503), .A2(n6502), .ZN(n6504) );
  NAND3_X1 U8176 ( .A1(n6504), .A2(n4259), .A3(n6572), .ZN(n6505) );
  NAND3_X1 U8177 ( .A1(n6531), .A2(n6576), .A3(n6505), .ZN(n6528) );
  INV_X1 U8178 ( .A(n7517), .ZN(n6584) );
  NAND2_X1 U8179 ( .A1(n6530), .A2(n6576), .ZN(n7138) );
  OR2_X1 U8180 ( .A1(n6584), .A2(n7138), .ZN(n7527) );
  NOR2_X1 U8181 ( .A1(n6509), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n6511) );
  NAND3_X1 U8182 ( .A1(n6519), .A2(n6052), .A3(n4952), .ZN(n6516) );
  NAND2_X1 U8183 ( .A1(n6515), .A2(n6512), .ZN(n6513) );
  NAND2_X1 U8184 ( .A1(n6513), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8185 ( .A1(n6516), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6517) );
  INV_X1 U8186 ( .A(n6519), .ZN(n6520) );
  OAI21_X1 U8187 ( .B1(n6228), .B2(n6520), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6522) );
  XNOR2_X1 U8188 ( .A(n6522), .B(n6521), .ZN(n6867) );
  AND2_X1 U8189 ( .A1(n6867), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6523) );
  INV_X1 U8190 ( .A(n8231), .ZN(n9672) );
  INV_X1 U8191 ( .A(n7410), .ZN(n9669) );
  NAND3_X1 U8192 ( .A1(n9769), .A2(n9672), .A3(n9669), .ZN(n6525) );
  OR2_X1 U8193 ( .A1(n7527), .A2(n6525), .ZN(n6527) );
  NOR2_X1 U8194 ( .A1(n6867), .A2(P1_U3084), .ZN(n10112) );
  INV_X1 U8195 ( .A(P1_B_REG_SCAN_IN), .ZN(n8230) );
  AOI21_X1 U8196 ( .B1(n6508), .B2(n10112), .A(n8230), .ZN(n6526) );
  NAND2_X1 U8197 ( .A1(n6527), .A2(n6526), .ZN(n6577) );
  INV_X1 U8198 ( .A(n6577), .ZN(n6581) );
  INV_X1 U8199 ( .A(n6533), .ZN(n6566) );
  INV_X1 U8200 ( .A(n6534), .ZN(n6557) );
  INV_X1 U8201 ( .A(n6535), .ZN(n6555) );
  INV_X1 U8202 ( .A(n6536), .ZN(n6551) );
  INV_X1 U8203 ( .A(n6537), .ZN(n6538) );
  OAI211_X1 U8204 ( .C1(n6080), .C2(n9724), .A(n4259), .B(n6538), .ZN(n6540)
         );
  NAND2_X1 U8205 ( .A1(n6540), .A2(n6539), .ZN(n6541) );
  OAI22_X1 U8206 ( .A1(n7137), .A2(n6541), .B1(n7440), .B2(n7589), .ZN(n6543)
         );
  NAND2_X1 U8207 ( .A1(n6543), .A2(n6542), .ZN(n6550) );
  INV_X1 U8208 ( .A(n6544), .ZN(n6548) );
  NAND2_X1 U8209 ( .A1(n7612), .A2(n6545), .ZN(n6547) );
  OAI22_X1 U8210 ( .A1(n6548), .A2(n7609), .B1(n6547), .B2(n6546), .ZN(n6549)
         );
  AOI21_X1 U8211 ( .B1(n6551), .B2(n6550), .A(n6549), .ZN(n6554) );
  INV_X1 U8212 ( .A(n6552), .ZN(n6553) );
  AOI21_X1 U8213 ( .B1(n6555), .B2(n6554), .A(n6553), .ZN(n6556) );
  NOR2_X1 U8214 ( .A1(n6557), .A2(n6556), .ZN(n6561) );
  INV_X1 U8215 ( .A(n6558), .ZN(n6560) );
  OAI21_X1 U8216 ( .B1(n6561), .B2(n6560), .A(n6559), .ZN(n6562) );
  NAND3_X1 U8217 ( .A1(n9296), .A2(n8224), .A3(n6562), .ZN(n6565) );
  INV_X1 U8218 ( .A(n6563), .ZN(n6564) );
  AOI21_X1 U8219 ( .B1(n6566), .B2(n6565), .A(n6564), .ZN(n6571) );
  INV_X1 U8220 ( .A(n6567), .ZN(n6570) );
  INV_X1 U8221 ( .A(n6568), .ZN(n6569) );
  NOR3_X1 U8222 ( .A1(n6571), .A2(n6570), .A3(n6569), .ZN(n6574) );
  OAI21_X1 U8223 ( .B1(n6574), .B2(n6573), .A(n6572), .ZN(n6575) );
  NAND4_X1 U8224 ( .A1(n6575), .A2(n9278), .A3(n6506), .A4(n6577), .ZN(n6580)
         );
  INV_X1 U8225 ( .A(n6575), .ZN(n6578) );
  NAND3_X1 U8226 ( .A1(n6578), .A2(n7139), .A3(n6577), .ZN(n6579) );
  OAI211_X1 U8227 ( .C1(n10112), .C2(n6581), .A(n6580), .B(n6579), .ZN(n6582)
         );
  AOI21_X1 U8228 ( .B1(n4956), .B2(n6583), .A(n6582), .ZN(P1_U3240) );
  INV_X1 U8229 ( .A(n9724), .ZN(n7265) );
  OR2_X4 U8230 ( .A1(n7517), .A2(n6591), .ZN(n6794) );
  OAI22_X1 U8231 ( .A1(n7265), .A2(n6794), .B1(n6606), .B2(n6080), .ZN(n6585)
         );
  NAND2_X1 U8232 ( .A1(n6584), .A2(n7138), .ZN(n6612) );
  XNOR2_X1 U8233 ( .A(n6585), .B(n6792), .ZN(n7356) );
  AND2_X1 U8234 ( .A1(n6508), .A2(n7139), .ZN(n6586) );
  NOR2_X1 U8235 ( .A1(n6606), .A2(n7265), .ZN(n6588) );
  AOI21_X1 U8236 ( .B1(n6614), .B2(n6587), .A(n6588), .ZN(n7353) );
  NAND2_X1 U8237 ( .A1(n6591), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6589) );
  AOI22_X1 U8238 ( .A1(n6603), .A2(n7462), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6591), .ZN(n6592) );
  OR2_X1 U8239 ( .A1(n7303), .A2(n6792), .ZN(n6594) );
  OAI21_X1 U8240 ( .B1(n7356), .B2(n7353), .A(n7354), .ZN(n6596) );
  NAND2_X1 U8241 ( .A1(n7356), .A2(n7353), .ZN(n6595) );
  NAND2_X1 U8242 ( .A1(n6596), .A2(n6595), .ZN(n7185) );
  OAI22_X1 U8243 ( .A1(n6605), .A2(n7440), .B1(n6093), .B2(n6606), .ZN(n6599)
         );
  OAI22_X1 U8244 ( .A1(n6093), .A2(n6794), .B1(n6606), .B2(n7440), .ZN(n6597)
         );
  XNOR2_X1 U8245 ( .A(n6597), .B(n6792), .ZN(n6598) );
  XNOR2_X1 U8246 ( .A(n6599), .B(n6598), .ZN(n7184) );
  NAND2_X1 U8247 ( .A1(n7185), .A2(n7184), .ZN(n6602) );
  INV_X1 U8248 ( .A(n6598), .ZN(n6600) );
  OR2_X1 U8249 ( .A1(n6600), .A2(n6599), .ZN(n6601) );
  OAI22_X1 U8250 ( .A1(n7521), .A2(n6794), .B1(n6606), .B2(n7670), .ZN(n6604)
         );
  XNOR2_X1 U8251 ( .A(n6604), .B(n6792), .ZN(n6607) );
  XNOR2_X1 U8252 ( .A(n6607), .B(n6608), .ZN(n7308) );
  INV_X1 U8253 ( .A(n6607), .ZN(n6609) );
  OR2_X1 U8254 ( .A1(n6609), .A2(n6608), .ZN(n6610) );
  OR2_X1 U8255 ( .A1(n6606), .A2(n7543), .ZN(n6611) );
  OAI21_X1 U8256 ( .B1(n6794), .B2(n4931), .A(n6611), .ZN(n6613) );
  XNOR2_X1 U8257 ( .A(n6613), .B(n7526), .ZN(n6618) );
  NAND2_X1 U8258 ( .A1(n6750), .A2(n9198), .ZN(n6616) );
  OR2_X1 U8259 ( .A1(n6606), .A2(n4931), .ZN(n6615) );
  NAND2_X1 U8260 ( .A1(n6616), .A2(n6615), .ZN(n6617) );
  XNOR2_X1 U8261 ( .A(n6618), .B(n6617), .ZN(n7674) );
  NAND2_X1 U8262 ( .A1(n6617), .A2(n6618), .ZN(n6619) );
  OR2_X1 U8263 ( .A1(n6791), .A2(n7740), .ZN(n6620) );
  OAI21_X1 U8264 ( .B1(n6794), .B2(n9781), .A(n6620), .ZN(n6621) );
  XNOR2_X1 U8265 ( .A(n6792), .B(n6621), .ZN(n7754) );
  NOR2_X1 U8266 ( .A1(n6606), .A2(n9781), .ZN(n6622) );
  AOI21_X1 U8267 ( .B1(n6750), .B2(n9197), .A(n6622), .ZN(n7756) );
  OAI22_X1 U8268 ( .A1(n9788), .A2(n6794), .B1(n6606), .B2(n7758), .ZN(n6623)
         );
  XNOR2_X1 U8269 ( .A(n6623), .B(n6792), .ZN(n7860) );
  INV_X1 U8270 ( .A(n7758), .ZN(n9196) );
  NOR2_X1 U8271 ( .A1(n6791), .A2(n9788), .ZN(n6624) );
  AOI21_X1 U8272 ( .B1(n6750), .B2(n9196), .A(n6624), .ZN(n7859) );
  AOI22_X1 U8273 ( .A1(n7754), .A2(n7756), .B1(n7860), .B2(n7859), .ZN(n6625)
         );
  NAND2_X1 U8274 ( .A1(n7857), .A2(n6625), .ZN(n6633) );
  INV_X1 U8275 ( .A(n7754), .ZN(n7858) );
  INV_X1 U8276 ( .A(n7756), .ZN(n6628) );
  NAND2_X1 U8277 ( .A1(n7858), .A2(n6628), .ZN(n6626) );
  NAND2_X1 U8278 ( .A1(n6626), .A2(n7859), .ZN(n6631) );
  INV_X1 U8279 ( .A(n7860), .ZN(n6630) );
  INV_X1 U8280 ( .A(n7859), .ZN(n6627) );
  AND2_X1 U8281 ( .A1(n6628), .A2(n6627), .ZN(n6629) );
  AOI22_X1 U8282 ( .A1(n6631), .A2(n6630), .B1(n6629), .B2(n7858), .ZN(n6632)
         );
  NAND2_X1 U8283 ( .A1(n6633), .A2(n6632), .ZN(n7683) );
  INV_X1 U8284 ( .A(n7910), .ZN(n9195) );
  NAND2_X1 U8285 ( .A1(n6761), .A2(n9195), .ZN(n6635) );
  NAND2_X1 U8286 ( .A1(n7791), .A2(n6744), .ZN(n6634) );
  NAND2_X1 U8287 ( .A1(n6635), .A2(n6634), .ZN(n6641) );
  INV_X1 U8288 ( .A(n6641), .ZN(n6640) );
  NAND2_X1 U8289 ( .A1(n6784), .A2(n7791), .ZN(n6637) );
  OR2_X1 U8290 ( .A1(n6791), .A2(n7910), .ZN(n6636) );
  NAND2_X1 U8291 ( .A1(n6637), .A2(n6636), .ZN(n6638) );
  XNOR2_X1 U8292 ( .A(n6638), .B(n7526), .ZN(n6642) );
  INV_X1 U8293 ( .A(n6642), .ZN(n6639) );
  NAND2_X1 U8294 ( .A1(n6640), .A2(n6639), .ZN(n7679) );
  AND2_X1 U8295 ( .A1(n6642), .A2(n6641), .ZN(n7680) );
  NAND2_X1 U8296 ( .A1(n9625), .A2(n6784), .ZN(n6644) );
  OR2_X1 U8297 ( .A1(n6606), .A2(n7880), .ZN(n6643) );
  NAND2_X1 U8298 ( .A1(n6644), .A2(n6643), .ZN(n6645) );
  XNOR2_X1 U8299 ( .A(n6645), .B(n7526), .ZN(n7949) );
  NAND2_X1 U8300 ( .A1(n9625), .A2(n6744), .ZN(n6647) );
  NAND2_X1 U8301 ( .A1(n6761), .A2(n9193), .ZN(n6646) );
  NAND2_X1 U8302 ( .A1(n6647), .A2(n6646), .ZN(n7948) );
  NAND2_X1 U8303 ( .A1(n6761), .A2(n9194), .ZN(n6649) );
  NAND2_X1 U8304 ( .A1(n7936), .A2(n6744), .ZN(n6648) );
  NAND2_X1 U8305 ( .A1(n6649), .A2(n6648), .ZN(n6654) );
  NAND2_X1 U8306 ( .A1(n7936), .A2(n6784), .ZN(n6651) );
  OR2_X1 U8307 ( .A1(n6791), .A2(n7688), .ZN(n6650) );
  NAND2_X1 U8308 ( .A1(n6651), .A2(n6650), .ZN(n6652) );
  XNOR2_X1 U8309 ( .A(n6652), .B(n7526), .ZN(n7946) );
  AOI22_X1 U8310 ( .A1(n7949), .A2(n7948), .B1(n6654), .B2(n7946), .ZN(n6653)
         );
  NAND2_X1 U8311 ( .A1(n7901), .A2(n6653), .ZN(n6661) );
  INV_X1 U8312 ( .A(n7949), .ZN(n6659) );
  INV_X1 U8313 ( .A(n7946), .ZN(n7905) );
  INV_X1 U8314 ( .A(n6654), .ZN(n7902) );
  NAND2_X1 U8315 ( .A1(n7905), .A2(n7902), .ZN(n6655) );
  NAND2_X1 U8316 ( .A1(n6655), .A2(n7948), .ZN(n6658) );
  INV_X1 U8317 ( .A(n6655), .ZN(n6657) );
  INV_X1 U8318 ( .A(n7948), .ZN(n6656) );
  AOI22_X1 U8319 ( .A1(n6659), .A2(n6658), .B1(n6657), .B2(n6656), .ZN(n6660)
         );
  OAI22_X1 U8320 ( .A1(n7893), .A2(n6794), .B1(n7969), .B2(n6606), .ZN(n6662)
         );
  XNOR2_X1 U8321 ( .A(n6662), .B(n6792), .ZN(n7875) );
  OR2_X1 U8322 ( .A1(n7893), .A2(n6791), .ZN(n6664) );
  INV_X1 U8323 ( .A(n6605), .ZN(n6750) );
  INV_X1 U8324 ( .A(n7969), .ZN(n9192) );
  NAND2_X1 U8325 ( .A1(n6750), .A2(n9192), .ZN(n6663) );
  INV_X1 U8326 ( .A(n7875), .ZN(n6666) );
  INV_X1 U8327 ( .A(n7874), .ZN(n6665) );
  NAND2_X1 U8328 ( .A1(n6666), .A2(n6665), .ZN(n6667) );
  OAI22_X1 U8329 ( .A1(n8057), .A2(n6794), .B1(n8041), .B2(n6791), .ZN(n6668)
         );
  XNOR2_X1 U8330 ( .A(n6668), .B(n6792), .ZN(n6671) );
  OR2_X1 U8331 ( .A1(n8057), .A2(n6606), .ZN(n6670) );
  NAND2_X1 U8332 ( .A1(n6750), .A2(n9191), .ZN(n6669) );
  NAND2_X1 U8333 ( .A1(n6670), .A2(n6669), .ZN(n6672) );
  XNOR2_X1 U8334 ( .A(n6671), .B(n6672), .ZN(n8008) );
  INV_X1 U8335 ( .A(n6671), .ZN(n6673) );
  OAI22_X1 U8336 ( .A1(n8128), .A2(n6794), .B1(n8136), .B2(n6791), .ZN(n6674)
         );
  XNOR2_X1 U8337 ( .A(n6674), .B(n7526), .ZN(n6676) );
  OR2_X1 U8338 ( .A1(n6676), .A2(n6675), .ZN(n6679) );
  NAND2_X1 U8339 ( .A1(n6676), .A2(n6675), .ZN(n6677) );
  NAND2_X1 U8340 ( .A1(n6679), .A2(n6677), .ZN(n8125) );
  INV_X1 U8341 ( .A(n6678), .ZN(n8122) );
  NAND2_X1 U8342 ( .A1(n9610), .A2(n6784), .ZN(n6681) );
  OR2_X1 U8343 ( .A1(n6606), .A2(n9049), .ZN(n6680) );
  NAND2_X1 U8344 ( .A1(n6681), .A2(n6680), .ZN(n6682) );
  XNOR2_X1 U8345 ( .A(n6682), .B(n6792), .ZN(n6684) );
  AOI21_X1 U8346 ( .B1(n9610), .B2(n6744), .A(n6683), .ZN(n6685) );
  AND2_X1 U8347 ( .A1(n6684), .A2(n6685), .ZN(n8161) );
  INV_X1 U8348 ( .A(n6684), .ZN(n6687) );
  INV_X1 U8349 ( .A(n6685), .ZN(n6686) );
  NAND2_X1 U8350 ( .A1(n6687), .A2(n6686), .ZN(n8162) );
  OAI21_X1 U8351 ( .B1(n8165), .B2(n8161), .A(n8162), .ZN(n9042) );
  OAI22_X1 U8352 ( .A1(n9490), .A2(n6794), .B1(n6688), .B2(n6791), .ZN(n6689)
         );
  XNOR2_X1 U8353 ( .A(n6689), .B(n7526), .ZN(n9094) );
  OR2_X1 U8354 ( .A1(n9490), .A2(n6606), .ZN(n6691) );
  NAND2_X1 U8355 ( .A1(n6750), .A2(n9458), .ZN(n6690) );
  NAND2_X1 U8356 ( .A1(n6691), .A2(n6690), .ZN(n6707) );
  NAND2_X1 U8357 ( .A1(n9595), .A2(n6744), .ZN(n6693) );
  NAND2_X1 U8358 ( .A1(n6750), .A2(n9448), .ZN(n6692) );
  NAND2_X1 U8359 ( .A1(n6693), .A2(n6692), .ZN(n9096) );
  OAI21_X1 U8360 ( .B1(n9094), .B2(n6707), .A(n9096), .ZN(n6697) );
  NAND2_X1 U8361 ( .A1(n9595), .A2(n6784), .ZN(n6695) );
  NAND2_X1 U8362 ( .A1(n6744), .A2(n9448), .ZN(n6694) );
  NAND2_X1 U8363 ( .A1(n6695), .A2(n6694), .ZN(n6696) );
  XNOR2_X1 U8364 ( .A(n6696), .B(n6792), .ZN(n9097) );
  NAND2_X1 U8365 ( .A1(n6697), .A2(n9097), .ZN(n6700) );
  INV_X1 U8366 ( .A(n9094), .ZN(n9091) );
  INV_X1 U8367 ( .A(n9096), .ZN(n6698) );
  INV_X1 U8368 ( .A(n6707), .ZN(n9176) );
  NAND3_X1 U8369 ( .A1(n9091), .A2(n6698), .A3(n9176), .ZN(n6699) );
  NAND2_X1 U8370 ( .A1(n9606), .A2(n6784), .ZN(n6702) );
  OR2_X1 U8371 ( .A1(n6791), .A2(n9476), .ZN(n6701) );
  NAND2_X1 U8372 ( .A1(n6702), .A2(n6701), .ZN(n6703) );
  XNOR2_X1 U8373 ( .A(n6703), .B(n7526), .ZN(n9046) );
  NAND2_X1 U8374 ( .A1(n9606), .A2(n6744), .ZN(n6705) );
  NAND2_X1 U8375 ( .A1(n6761), .A2(n9511), .ZN(n6704) );
  NAND2_X1 U8376 ( .A1(n6705), .A2(n6704), .ZN(n9089) );
  INV_X1 U8377 ( .A(n9046), .ZN(n9044) );
  INV_X1 U8378 ( .A(n9089), .ZN(n9047) );
  INV_X1 U8379 ( .A(n9097), .ZN(n6708) );
  AOI22_X1 U8380 ( .A1(n6708), .A2(n9096), .B1(n9094), .B2(n6707), .ZN(n9105)
         );
  OAI21_X1 U8381 ( .B1(n9044), .B2(n9047), .A(n9105), .ZN(n6709) );
  NAND2_X1 U8382 ( .A1(n6709), .A2(n9106), .ZN(n6714) );
  NAND2_X1 U8383 ( .A1(n9589), .A2(n6784), .ZN(n6711) );
  NAND2_X1 U8384 ( .A1(n9457), .A2(n6744), .ZN(n6710) );
  NAND2_X1 U8385 ( .A1(n6711), .A2(n6710), .ZN(n6712) );
  XNOR2_X1 U8386 ( .A(n6712), .B(n7526), .ZN(n6716) );
  AND2_X1 U8387 ( .A1(n6761), .A2(n9457), .ZN(n6713) );
  AOI21_X1 U8388 ( .B1(n9589), .B2(n6744), .A(n6713), .ZN(n6717) );
  XNOR2_X1 U8389 ( .A(n6716), .B(n6717), .ZN(n9110) );
  INV_X1 U8390 ( .A(n6716), .ZN(n6718) );
  OAI22_X1 U8391 ( .A1(n9431), .A2(n6794), .B1(n6720), .B2(n6791), .ZN(n6719)
         );
  XNOR2_X1 U8392 ( .A(n6719), .B(n6792), .ZN(n9149) );
  OR2_X1 U8393 ( .A1(n9431), .A2(n6606), .ZN(n6722) );
  NAND2_X1 U8394 ( .A1(n9450), .A2(n6750), .ZN(n6721) );
  AND2_X1 U8395 ( .A1(n6722), .A2(n6721), .ZN(n9148) );
  NAND2_X1 U8396 ( .A1(n9580), .A2(n6784), .ZN(n6724) );
  NAND2_X1 U8397 ( .A1(n9436), .A2(n6744), .ZN(n6723) );
  NAND2_X1 U8398 ( .A1(n6724), .A2(n6723), .ZN(n6725) );
  XNOR2_X1 U8399 ( .A(n6725), .B(n7526), .ZN(n6727) );
  AND2_X1 U8400 ( .A1(n9436), .A2(n6761), .ZN(n6726) );
  AOI21_X1 U8401 ( .B1(n9580), .B2(n6744), .A(n6726), .ZN(n6728) );
  XNOR2_X1 U8402 ( .A(n6727), .B(n6728), .ZN(n9065) );
  INV_X1 U8403 ( .A(n6727), .ZN(n6729) );
  NAND2_X1 U8404 ( .A1(n6729), .A2(n6728), .ZN(n6730) );
  OAI22_X1 U8405 ( .A1(n9404), .A2(n6794), .B1(n6731), .B2(n6791), .ZN(n6732)
         );
  XNOR2_X1 U8406 ( .A(n6732), .B(n7526), .ZN(n6735) );
  OR2_X1 U8407 ( .A1(n9404), .A2(n6606), .ZN(n6734) );
  NAND2_X1 U8408 ( .A1(n9420), .A2(n6761), .ZN(n6733) );
  NAND2_X1 U8409 ( .A1(n6734), .A2(n6733), .ZN(n6736) );
  NAND2_X1 U8410 ( .A1(n6735), .A2(n6736), .ZN(n9127) );
  NAND2_X1 U8411 ( .A1(n9130), .A2(n9127), .ZN(n6739) );
  INV_X1 U8412 ( .A(n6735), .ZN(n6738) );
  INV_X1 U8413 ( .A(n6736), .ZN(n6737) );
  NAND2_X1 U8414 ( .A1(n6738), .A2(n6737), .ZN(n9128) );
  NAND2_X1 U8415 ( .A1(n6739), .A2(n9128), .ZN(n9072) );
  NAND2_X1 U8416 ( .A1(n9570), .A2(n6784), .ZN(n6741) );
  NAND2_X1 U8417 ( .A1(n9408), .A2(n6744), .ZN(n6740) );
  NAND2_X1 U8418 ( .A1(n6741), .A2(n6740), .ZN(n6742) );
  XNOR2_X1 U8419 ( .A(n6742), .B(n7526), .ZN(n6745) );
  AOI21_X1 U8420 ( .B1(n9570), .B2(n6744), .A(n6743), .ZN(n6746) );
  XNOR2_X1 U8421 ( .A(n6745), .B(n6746), .ZN(n9073) );
  NAND2_X1 U8422 ( .A1(n9072), .A2(n9073), .ZN(n6749) );
  INV_X1 U8423 ( .A(n6745), .ZN(n6747) );
  NAND2_X1 U8424 ( .A1(n6747), .A2(n6746), .ZN(n6748) );
  NAND2_X1 U8425 ( .A1(n6749), .A2(n6748), .ZN(n6754) );
  OR2_X1 U8426 ( .A1(n9373), .A2(n6791), .ZN(n6752) );
  NAND2_X1 U8427 ( .A1(n9392), .A2(n6750), .ZN(n6751) );
  AND2_X1 U8428 ( .A1(n6752), .A2(n6751), .ZN(n6755) );
  NAND2_X1 U8429 ( .A1(n6754), .A2(n6755), .ZN(n9137) );
  OAI22_X1 U8430 ( .A1(n9373), .A2(n6794), .B1(n9076), .B2(n6606), .ZN(n6753)
         );
  XNOR2_X1 U8431 ( .A(n6753), .B(n7526), .ZN(n9140) );
  INV_X1 U8432 ( .A(n6754), .ZN(n6757) );
  INV_X1 U8433 ( .A(n6755), .ZN(n6756) );
  NAND2_X1 U8434 ( .A1(n9559), .A2(n6784), .ZN(n6759) );
  NAND2_X1 U8435 ( .A1(n9377), .A2(n6744), .ZN(n6758) );
  NAND2_X1 U8436 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  XNOR2_X1 U8437 ( .A(n6760), .B(n7526), .ZN(n6763) );
  AND2_X1 U8438 ( .A1(n9377), .A2(n6761), .ZN(n6762) );
  AOI21_X1 U8439 ( .B1(n9559), .B2(n6744), .A(n6762), .ZN(n9057) );
  OAI22_X1 U8440 ( .A1(n9344), .A2(n6794), .B1(n9083), .B2(n6791), .ZN(n6764)
         );
  XNOR2_X1 U8441 ( .A(n6764), .B(n6792), .ZN(n6767) );
  OR2_X1 U8442 ( .A1(n9344), .A2(n6606), .ZN(n6766) );
  NAND2_X1 U8443 ( .A1(n9362), .A2(n6750), .ZN(n6765) );
  AND2_X1 U8444 ( .A1(n6766), .A2(n6765), .ZN(n6768) );
  NAND2_X1 U8445 ( .A1(n6767), .A2(n6768), .ZN(n6772) );
  INV_X1 U8446 ( .A(n6767), .ZN(n6770) );
  INV_X1 U8447 ( .A(n6768), .ZN(n6769) );
  NAND2_X1 U8448 ( .A1(n6770), .A2(n6769), .ZN(n6771) );
  NAND2_X1 U8449 ( .A1(n6772), .A2(n6771), .ZN(n9116) );
  INV_X1 U8450 ( .A(n6772), .ZN(n6773) );
  AOI22_X1 U8451 ( .A1(n9550), .A2(n6784), .B1(n6744), .B2(n9348), .ZN(n6774)
         );
  XNOR2_X1 U8452 ( .A(n6774), .B(n7526), .ZN(n6780) );
  AOI21_X1 U8453 ( .B1(n9550), .B2(n6744), .A(n6775), .ZN(n6779) );
  XNOR2_X1 U8454 ( .A(n6780), .B(n6779), .ZN(n9080) );
  OAI22_X1 U8455 ( .A1(n9311), .A2(n6794), .B1(n6862), .B2(n6791), .ZN(n6776)
         );
  XNOR2_X1 U8456 ( .A(n6776), .B(n7526), .ZN(n6783) );
  OR2_X1 U8457 ( .A1(n9311), .A2(n6606), .ZN(n6778) );
  NAND2_X1 U8458 ( .A1(n9334), .A2(n6761), .ZN(n6777) );
  NAND2_X1 U8459 ( .A1(n6778), .A2(n6777), .ZN(n6782) );
  XNOR2_X1 U8460 ( .A(n6783), .B(n6782), .ZN(n9161) );
  AND2_X1 U8461 ( .A1(n6780), .A2(n6779), .ZN(n9162) );
  NAND2_X1 U8462 ( .A1(n9543), .A2(n6784), .ZN(n6786) );
  NAND2_X1 U8463 ( .A1(n9316), .A2(n6744), .ZN(n6785) );
  NAND2_X1 U8464 ( .A1(n6786), .A2(n6785), .ZN(n6787) );
  XNOR2_X1 U8465 ( .A(n6787), .B(n6792), .ZN(n6790) );
  AOI21_X1 U8466 ( .B1(n9543), .B2(n6744), .A(n6788), .ZN(n6789) );
  NAND2_X1 U8467 ( .A1(n6790), .A2(n6789), .ZN(n6832) );
  OAI21_X1 U8468 ( .B1(n6790), .B2(n6789), .A(n6832), .ZN(n6859) );
  XNOR2_X1 U8469 ( .A(n6793), .B(n6792), .ZN(n6796) );
  OAI22_X1 U8470 ( .A1(n8301), .A2(n6794), .B1(n6863), .B2(n6606), .ZN(n6795)
         );
  XNOR2_X1 U8471 ( .A(n6796), .B(n6795), .ZN(n6816) );
  INV_X1 U8472 ( .A(n6816), .ZN(n6833) );
  NAND2_X1 U8473 ( .A1(n8099), .A2(n8230), .ZN(n6797) );
  OR2_X1 U8474 ( .A1(n9736), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6800) );
  OR2_X1 U8475 ( .A1(n9675), .A2(n8099), .ZN(n6799) );
  NAND2_X1 U8476 ( .A1(n6800), .A2(n6799), .ZN(n7450) );
  INV_X1 U8477 ( .A(n7450), .ZN(n9657) );
  NOR2_X1 U8478 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .ZN(
        n6804) );
  NOR4_X1 U8479 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6803) );
  NOR4_X1 U8480 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6802) );
  NOR4_X1 U8481 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6801) );
  NAND4_X1 U8482 ( .A1(n6804), .A2(n6803), .A3(n6802), .A4(n6801), .ZN(n6810)
         );
  NOR4_X1 U8483 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6808) );
  NOR4_X1 U8484 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6807) );
  NOR4_X1 U8485 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6806) );
  NOR4_X1 U8486 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6805) );
  NAND4_X1 U8487 ( .A1(n6808), .A2(n6807), .A3(n6806), .A4(n6805), .ZN(n6809)
         );
  NOR2_X1 U8488 ( .A1(n6810), .A2(n6809), .ZN(n6811) );
  NAND2_X1 U8489 ( .A1(n9657), .A2(n7449), .ZN(n7150) );
  OR2_X1 U8490 ( .A1(n9736), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6813) );
  OR2_X1 U8491 ( .A1(n9675), .A2(n8159), .ZN(n6812) );
  NAND2_X1 U8492 ( .A1(n6813), .A2(n6812), .ZN(n7451) );
  NOR2_X1 U8493 ( .A1(n7150), .A2(n7451), .ZN(n6826) );
  NAND2_X1 U8494 ( .A1(n6820), .A2(n7142), .ZN(n6814) );
  NAND3_X1 U8495 ( .A1(n6833), .A2(n9165), .A3(n6832), .ZN(n6815) );
  NOR2_X1 U8496 ( .A1(n7702), .A2(n6506), .ZN(n9725) );
  NAND2_X1 U8497 ( .A1(n9725), .A2(n6820), .ZN(n6819) );
  OR2_X1 U8498 ( .A1(n4259), .A2(n9738), .ZN(n6818) );
  INV_X1 U8499 ( .A(n6820), .ZN(n6821) );
  NOR2_X1 U8500 ( .A1(n7527), .A2(n6821), .ZN(n6822) );
  NAND2_X1 U8501 ( .A1(n6822), .A2(n9669), .ZN(n9178) );
  INV_X1 U8502 ( .A(n8305), .ZN(n9189) );
  NAND2_X1 U8503 ( .A1(n6822), .A2(n7410), .ZN(n9152) );
  NAND2_X1 U8504 ( .A1(n9189), .A2(n9180), .ZN(n6831) );
  INV_X1 U8505 ( .A(n6823), .ZN(n8299) );
  AND3_X1 U8506 ( .A1(n7148), .A2(n6868), .A3(n6867), .ZN(n6824) );
  OR2_X1 U8507 ( .A1(n9626), .A2(n6826), .ZN(n7186) );
  NAND2_X1 U8508 ( .A1(n6824), .A2(n7186), .ZN(n6825) );
  NAND2_X1 U8509 ( .A1(n6825), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6829) );
  INV_X1 U8510 ( .A(n6826), .ZN(n6827) );
  AND2_X1 U8511 ( .A1(n6827), .A2(n9769), .ZN(n6828) );
  NAND2_X1 U8512 ( .A1(n9725), .A2(n6828), .ZN(n7188) );
  AOI22_X1 U8513 ( .A1(n8299), .A2(n9167), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6830) );
  OAI211_X1 U8514 ( .C1(n8306), .C2(n9178), .A(n6831), .B(n6830), .ZN(n6835)
         );
  NOR3_X1 U8515 ( .A1(n6833), .A2(n6832), .A3(n9186), .ZN(n6834) );
  AOI211_X1 U8516 ( .C1(n9536), .C2(n9184), .A(n6835), .B(n6834), .ZN(n6836)
         );
  NAND3_X1 U8517 ( .A1(n6838), .A2(n6837), .A3(n6836), .ZN(P1_U3218) );
  INV_X1 U8518 ( .A(n6839), .ZN(n6840) );
  NAND2_X1 U8519 ( .A1(n6841), .A2(n6840), .ZN(n6852) );
  NOR2_X1 U8520 ( .A1(n8632), .A2(n7328), .ZN(n6842) );
  XNOR2_X1 U8521 ( .A(n6842), .B(n4274), .ZN(n6844) );
  INV_X1 U8522 ( .A(n6844), .ZN(n6845) );
  NOR3_X1 U8523 ( .A1(n8263), .A2(n8445), .A3(n6845), .ZN(n6843) );
  AOI21_X1 U8524 ( .B1(n8263), .B2(n6845), .A(n6843), .ZN(n6851) );
  NOR3_X1 U8525 ( .A1(n8263), .A2(n6844), .A3(n8445), .ZN(n6847) );
  NOR2_X1 U8526 ( .A1(n8900), .A2(n6845), .ZN(n6846) );
  NAND2_X1 U8527 ( .A1(n6852), .A2(n6848), .ZN(n6850) );
  OAI21_X1 U8528 ( .B1(n8263), .B2(n8432), .A(n8447), .ZN(n6849) );
  OAI211_X1 U8529 ( .C1(n6852), .C2(n6851), .A(n6850), .B(n6849), .ZN(n6857)
         );
  NOR2_X1 U8530 ( .A1(n6853), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6855) );
  OAI22_X1 U8531 ( .A1(n8268), .A2(n8441), .B1(n8424), .B2(n8440), .ZN(n6854)
         );
  AOI211_X1 U8532 ( .C1(n8261), .C2(n8429), .A(n6855), .B(n6854), .ZN(n6856)
         );
  NAND2_X1 U8533 ( .A1(n6857), .A2(n6856), .ZN(P2_U3222) );
  OAI22_X1 U8534 ( .A1(n6862), .A2(n9178), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6861), .ZN(n6865) );
  NOR2_X1 U8535 ( .A1(n6863), .A2(n9152), .ZN(n6864) );
  AOI211_X1 U8536 ( .C1(n9301), .C2(n9167), .A(n6865), .B(n6864), .ZN(n6866)
         );
  INV_X1 U8537 ( .A(n6867), .ZN(n6880) );
  INV_X1 U8538 ( .A(n9837), .ZN(n6869) );
  INV_X1 U8539 ( .A(n6870), .ZN(n6875) );
  AOI21_X1 U8540 ( .B1(n6874), .B2(n6872), .A(n6871), .ZN(n6873) );
  AOI211_X1 U8541 ( .C1(n6875), .C2(n6874), .A(n8447), .B(n6873), .ZN(n6879)
         );
  INV_X1 U8542 ( .A(n8085), .ZN(n9894) );
  NOR2_X1 U8543 ( .A1(n8432), .A2(n9894), .ZN(n6878) );
  OAI22_X1 U8544 ( .A1(n8439), .A2(n8083), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8557), .ZN(n6877) );
  OAI22_X1 U8545 ( .A1(n7725), .A2(n8440), .B1(n8441), .B2(n8021), .ZN(n6876)
         );
  OR4_X1 U8546 ( .A1(n6879), .A2(n6878), .A3(n6877), .A4(n6876), .ZN(P2_U3233)
         );
  NAND2_X1 U8547 ( .A1(n6881), .A2(n6928), .ZN(n6899) );
  OR2_X1 U8548 ( .A1(n6899), .A2(n7276), .ZN(n6882) );
  NAND2_X1 U8549 ( .A1(n6882), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8550 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6883) );
  INV_X1 U8551 ( .A(n6904), .ZN(n7244) );
  NAND2_X1 U8552 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n7408) );
  INV_X1 U8553 ( .A(n7408), .ZN(n7240) );
  OAI21_X1 U8554 ( .B1(n6883), .B2(n7244), .A(n7239), .ZN(n9202) );
  INV_X1 U8555 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6884) );
  XNOR2_X1 U8556 ( .A(n9205), .B(n6884), .ZN(n9203) );
  XNOR2_X1 U8557 ( .A(n6937), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n7385) );
  AOI21_X1 U8558 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6937), .A(n7384), .ZN(
        n7401) );
  INV_X1 U8559 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6885) );
  MUX2_X1 U8560 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6885), .S(n7403), .Z(n7400)
         );
  INV_X1 U8561 ( .A(n7400), .ZN(n6886) );
  AOI22_X1 U8562 ( .A1(n7401), .A2(n6886), .B1(n7403), .B2(n6885), .ZN(n7343)
         );
  XNOR2_X1 U8563 ( .A(n6946), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n7344) );
  XNOR2_X1 U8564 ( .A(n9217), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9215) );
  NOR2_X1 U8565 ( .A1(n9214), .A2(n9215), .ZN(n9213) );
  INV_X1 U8566 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6887) );
  MUX2_X1 U8567 ( .A(n6887), .B(P1_REG2_REG_7__SCAN_IN), .S(n6916), .Z(n6888)
         );
  INV_X1 U8568 ( .A(n6888), .ZN(n7246) );
  INV_X1 U8569 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6889) );
  MUX2_X1 U8570 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n6889), .S(n6966), .Z(n6890)
         );
  INV_X1 U8571 ( .A(n6890), .ZN(n7177) );
  XNOR2_X1 U8572 ( .A(n7433), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7430) );
  NOR2_X1 U8573 ( .A1(n7429), .A2(n7430), .ZN(n7428) );
  XNOR2_X1 U8574 ( .A(n7423), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7419) );
  XOR2_X1 U8575 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7296), .Z(n7295) );
  XNOR2_X1 U8576 ( .A(n7556), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7553) );
  INV_X1 U8577 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6891) );
  MUX2_X1 U8578 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n6891), .S(n7713), .Z(n6892)
         );
  INV_X1 U8579 ( .A(n6892), .ZN(n7709) );
  INV_X1 U8580 ( .A(n9234), .ZN(n7021) );
  NOR2_X1 U8581 ( .A1(n6893), .A2(n7021), .ZN(n6894) );
  INV_X1 U8582 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9231) );
  NOR2_X1 U8583 ( .A1(n6895), .A2(n7126), .ZN(n6896) );
  INV_X1 U8584 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10016) );
  NAND2_X1 U8585 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7288), .ZN(n6897) );
  OAI21_X1 U8586 ( .B1(n7288), .B2(P1_REG2_REG_16__SCAN_IN), .A(n6897), .ZN(
        n9253) );
  NAND2_X1 U8587 ( .A1(n9272), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6898) );
  OAI21_X1 U8588 ( .B1(n9272), .B2(P1_REG2_REG_17__SCAN_IN), .A(n6898), .ZN(
        n6901) );
  INV_X1 U8589 ( .A(n7281), .ZN(n6900) );
  NOR2_X1 U8590 ( .A1(n6900), .A2(n7410), .ZN(n6923) );
  AOI211_X1 U8591 ( .C1(n6902), .C2(n6901), .A(n9265), .B(n9251), .ZN(n6935)
         );
  XNOR2_X1 U8592 ( .A(n7021), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9227) );
  INV_X1 U8593 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7666) );
  INV_X1 U8594 ( .A(n6916), .ZN(n7257) );
  INV_X1 U8595 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6903) );
  MUX2_X1 U8596 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6903), .S(n6904), .Z(n7235)
         );
  AND2_X1 U8597 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n7236) );
  NAND2_X1 U8598 ( .A1(n7235), .A2(n7236), .ZN(n7234) );
  NAND2_X1 U8599 ( .A1(n6904), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U8600 ( .A1(n7234), .A2(n6905), .ZN(n9206) );
  INV_X1 U8601 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6906) );
  XNOR2_X1 U8602 ( .A(n9205), .B(n6906), .ZN(n9207) );
  NAND2_X1 U8603 ( .A1(n9206), .A2(n9207), .ZN(n6908) );
  NAND2_X1 U8604 ( .A1(n9205), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6907) );
  NAND2_X1 U8605 ( .A1(n6908), .A2(n6907), .ZN(n7390) );
  INV_X1 U8606 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U8607 ( .A1(n6937), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U8608 ( .A1(n7389), .A2(n6910), .ZN(n7395) );
  INV_X1 U8609 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6911) );
  MUX2_X1 U8610 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6911), .S(n7403), .Z(n6912)
         );
  NAND2_X1 U8611 ( .A1(n7403), .A2(n6911), .ZN(n6913) );
  AND2_X1 U8612 ( .A1(n7396), .A2(n6913), .ZN(n7349) );
  INV_X1 U8613 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6914) );
  MUX2_X1 U8614 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6914), .S(n6946), .Z(n7348)
         );
  NAND2_X1 U8615 ( .A1(n7349), .A2(n7348), .ZN(n7347) );
  NAND2_X1 U8616 ( .A1(n6946), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6915) );
  INV_X1 U8617 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9984) );
  MUX2_X1 U8618 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n9984), .S(n9217), .Z(n9219)
         );
  NAND2_X1 U8619 ( .A1(n9220), .A2(n9219), .ZN(n9218) );
  INV_X1 U8620 ( .A(n9217), .ZN(n6950) );
  NAND2_X1 U8621 ( .A1(n6950), .A2(n9984), .ZN(n7251) );
  MUX2_X1 U8622 ( .A(n7666), .B(P1_REG1_REG_7__SCAN_IN), .S(n6916), .Z(n7252)
         );
  AOI21_X1 U8623 ( .B1(n7666), .B2(n7257), .A(n7254), .ZN(n7174) );
  AND2_X1 U8624 ( .A1(n7178), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7172) );
  INV_X1 U8625 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U8626 ( .A1(n6966), .A2(n6917), .ZN(n7170) );
  OAI21_X1 U8627 ( .B1(n7174), .B2(n7172), .A(n7170), .ZN(n7426) );
  INV_X1 U8628 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6918) );
  XNOR2_X1 U8629 ( .A(n7433), .B(n6918), .ZN(n7427) );
  INV_X1 U8630 ( .A(n7433), .ZN(n6973) );
  AOI22_X1 U8631 ( .A1(n7426), .A2(n7427), .B1(n6973), .B2(n6918), .ZN(n7413)
         );
  XNOR2_X1 U8632 ( .A(n7423), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7414) );
  XOR2_X1 U8633 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n7296), .Z(n7292) );
  INV_X1 U8634 ( .A(n7296), .ZN(n6980) );
  INV_X1 U8635 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6919) );
  AOI22_X1 U8636 ( .A1(n7291), .A2(n7292), .B1(n6980), .B2(n6919), .ZN(n7549)
         );
  XNOR2_X1 U8637 ( .A(n7556), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7550) );
  INV_X1 U8638 ( .A(n7706), .ZN(n6920) );
  XNOR2_X1 U8639 ( .A(n7713), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7705) );
  OAI22_X1 U8640 ( .A1(n6920), .A2(n7705), .B1(n7713), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n9228) );
  NOR2_X1 U8641 ( .A1(n7126), .A2(n6921), .ZN(n6922) );
  INV_X1 U8642 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9242) );
  XNOR2_X1 U8643 ( .A(n7126), .B(n6921), .ZN(n9243) );
  NOR2_X1 U8644 ( .A1(n9242), .A2(n9243), .ZN(n9241) );
  XNOR2_X1 U8645 ( .A(n7288), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9256) );
  NOR2_X1 U8646 ( .A1(n9257), .A2(n9256), .ZN(n9255) );
  AOI21_X1 U8647 ( .B1(n7288), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9255), .ZN(
        n6925) );
  XNOR2_X1 U8648 ( .A(n9272), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n6924) );
  NOR2_X1 U8649 ( .A1(n6925), .A2(n6924), .ZN(n9271) );
  AOI211_X1 U8650 ( .C1(n6925), .C2(n6924), .A(n9271), .B(n9254), .ZN(n6934)
         );
  NAND2_X1 U8651 ( .A1(n7281), .A2(n9672), .ZN(n9275) );
  INV_X1 U8652 ( .A(n9275), .ZN(n6926) );
  INV_X1 U8653 ( .A(n9272), .ZN(n6927) );
  NOR2_X1 U8654 ( .A1(n9261), .A2(n6927), .ZN(n6933) );
  INV_X1 U8655 ( .A(P1_U3083), .ZN(n6929) );
  INV_X1 U8656 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U8657 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n6930) );
  OAI21_X1 U8658 ( .B1(n9281), .B2(n6931), .A(n6930), .ZN(n6932) );
  OR4_X1 U8659 ( .A1(n6935), .A2(n6934), .A3(n6933), .A4(n6932), .ZN(P1_U3258)
         );
  NOR2_X2 U8660 ( .A1(n4257), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10113) );
  INV_X1 U8661 ( .A(n10113), .ZN(n7855) );
  INV_X1 U8662 ( .A(n6936), .ZN(n6959) );
  INV_X1 U8663 ( .A(n6937), .ZN(n7394) );
  OAI222_X1 U8664 ( .A1(n7855), .A2(n6938), .B1(n10109), .B2(n6959), .C1(
        P1_U3084), .C2(n7394), .ZN(P1_U3350) );
  INV_X1 U8665 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6939) );
  OAI222_X1 U8666 ( .A1(n7244), .A2(P1_U3084), .B1(n10109), .B2(n6958), .C1(
        n6939), .C2(n7855), .ZN(P1_U3352) );
  INV_X1 U8667 ( .A(n9205), .ZN(n6940) );
  OAI222_X1 U8668 ( .A1(n6940), .A2(P1_U3084), .B1(n10109), .B2(n6956), .C1(
        n5055), .C2(n7855), .ZN(P1_U3351) );
  INV_X1 U8669 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6942) );
  INV_X1 U8670 ( .A(n6941), .ZN(n6960) );
  OAI222_X1 U8671 ( .A1(n7855), .A2(n6942), .B1(n10109), .B2(n6960), .C1(
        P1_U3084), .C2(n7403), .ZN(P1_U3349) );
  INV_X1 U8672 ( .A(n6943), .ZN(n6947) );
  AND2_X1 U8673 ( .A1(n4256), .A2(P2_U3152), .ZN(n9026) );
  AOI22_X1 U8674 ( .A1(n8499), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n9026), .ZN(n6945) );
  OAI21_X1 U8675 ( .B1(n6947), .B2(n9038), .A(n6945), .ZN(P2_U3353) );
  INV_X1 U8676 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6948) );
  INV_X1 U8677 ( .A(n6946), .ZN(n7352) );
  OAI222_X1 U8678 ( .A1(n7855), .A2(n6948), .B1(n10109), .B2(n6947), .C1(
        P1_U3084), .C2(n7352), .ZN(P1_U3348) );
  INV_X1 U8679 ( .A(n9026), .ZN(n9040) );
  INV_X1 U8680 ( .A(n6949), .ZN(n6951) );
  INV_X1 U8681 ( .A(n8514), .ZN(n7061) );
  OAI222_X1 U8682 ( .A1(n9040), .A2(n4363), .B1(n9038), .B2(n6951), .C1(
        P2_U3152), .C2(n7061), .ZN(P2_U3352) );
  INV_X1 U8683 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6952) );
  OAI222_X1 U8684 ( .A1(n7855), .A2(n6952), .B1(n10109), .B2(n6951), .C1(
        P1_U3084), .C2(n6950), .ZN(P1_U3347) );
  INV_X1 U8685 ( .A(n6953), .ZN(n6962) );
  AOI22_X1 U8686 ( .A1(n8528), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n9026), .ZN(n6954) );
  OAI21_X1 U8687 ( .B1(n6962), .B2(n9038), .A(n6954), .ZN(P2_U3351) );
  INV_X1 U8688 ( .A(n7039), .ZN(n7057) );
  OAI222_X1 U8689 ( .A1(n7057), .A2(P2_U3152), .B1(n9038), .B2(n6956), .C1(
        n6955), .C2(n9040), .ZN(P2_U3356) );
  INV_X1 U8690 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6957) );
  OAI222_X1 U8691 ( .A1(n7020), .A2(P2_U3152), .B1(n9038), .B2(n6958), .C1(
        n6957), .C2(n9040), .ZN(P2_U3357) );
  OAI222_X1 U8692 ( .A1(n9040), .A2(n5050), .B1(n9038), .B2(n6959), .C1(
        P2_U3152), .C2(n7058), .ZN(P2_U3355) );
  INV_X1 U8693 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6961) );
  INV_X1 U8694 ( .A(n8486), .ZN(n7060) );
  OAI222_X1 U8695 ( .A1(n9040), .A2(n6961), .B1(n9038), .B2(n6960), .C1(
        P2_U3152), .C2(n7060), .ZN(P2_U3354) );
  INV_X1 U8696 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6963) );
  OAI222_X1 U8697 ( .A1(n7855), .A2(n6963), .B1(n10109), .B2(n6962), .C1(
        P1_U3084), .C2(n7257), .ZN(P1_U3346) );
  INV_X1 U8698 ( .A(n6964), .ZN(n6967) );
  OAI222_X1 U8699 ( .A1(n9040), .A2(n6965), .B1(n9038), .B2(n6967), .C1(
        P2_U3152), .C2(n8538), .ZN(P2_U3350) );
  OAI222_X1 U8700 ( .A1(n7855), .A2(n6968), .B1(n10109), .B2(n6967), .C1(
        P1_U3084), .C2(n6966), .ZN(P1_U3345) );
  INV_X1 U8701 ( .A(n6969), .ZN(n6974) );
  AOI22_X1 U8702 ( .A1(n8562), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9026), .ZN(n6970) );
  OAI21_X1 U8703 ( .B1(n6974), .B2(n9038), .A(n6970), .ZN(P2_U3349) );
  INV_X1 U8704 ( .A(n6971), .ZN(n6976) );
  AOI22_X1 U8705 ( .A1(n7423), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10113), .ZN(n6972) );
  OAI21_X1 U8706 ( .B1(n6976), .B2(n10109), .A(n6972), .ZN(P1_U3343) );
  OAI222_X1 U8707 ( .A1(n7855), .A2(n6975), .B1(n10109), .B2(n6974), .C1(n6973), .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8708 ( .A(n7064), .ZN(n7078) );
  OAI222_X1 U8709 ( .A1(n9040), .A2(n6977), .B1(n9038), .B2(n6976), .C1(n7078), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8710 ( .A(n6978), .ZN(n6981) );
  INV_X1 U8711 ( .A(n7065), .ZN(n7093) );
  OAI222_X1 U8712 ( .A1(n9040), .A2(n6979), .B1(n9038), .B2(n6981), .C1(n7093), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  OAI222_X1 U8713 ( .A1(n7855), .A2(n6982), .B1(n10109), .B2(n6981), .C1(n6980), .C2(P1_U3084), .ZN(P1_U3342) );
  NAND2_X1 U8714 ( .A1(n9830), .A2(n7001), .ZN(n6984) );
  NAND2_X1 U8715 ( .A1(n6984), .A2(n4258), .ZN(n6987) );
  OR2_X1 U8716 ( .A1(n9830), .A2(n6985), .ZN(n6986) );
  NOR2_X1 U8717 ( .A1(n9817), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U8718 ( .A1(P2_U3966), .A2(n8588), .ZN(n6988) );
  OAI21_X1 U8719 ( .B1(P2_U3966), .B2(n5596), .A(n6988), .ZN(P2_U3583) );
  NAND2_X1 U8720 ( .A1(n9282), .A2(n9200), .ZN(n6989) );
  OAI21_X1 U8721 ( .B1(n9200), .B2(n5597), .A(n6989), .ZN(P1_U3586) );
  INV_X1 U8722 ( .A(n6990), .ZN(n6994) );
  AOI22_X1 U8723 ( .A1(n7556), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10113), .ZN(n6991) );
  OAI21_X1 U8724 ( .B1(n6994), .B2(n10109), .A(n6991), .ZN(P1_U3341) );
  INV_X1 U8725 ( .A(n6992), .ZN(n6996) );
  AOI22_X1 U8726 ( .A1(n7713), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10113), .ZN(n6993) );
  OAI21_X1 U8727 ( .B1(n6996), .B2(n10109), .A(n6993), .ZN(P1_U3340) );
  INV_X1 U8728 ( .A(n7071), .ZN(n7159) );
  OAI222_X1 U8729 ( .A1(n9040), .A2(n6995), .B1(n9038), .B2(n6994), .C1(
        P2_U3152), .C2(n7159), .ZN(P2_U3346) );
  INV_X1 U8730 ( .A(n7211), .ZN(n7158) );
  OAI222_X1 U8731 ( .A1(n9040), .A2(n10071), .B1(n9038), .B2(n6996), .C1(n7158), .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8732 ( .A(n6997), .ZN(n7022) );
  AOI22_X1 U8733 ( .A1(n7491), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n9026), .ZN(n6998) );
  OAI21_X1 U8734 ( .B1(n7022), .B2(n9038), .A(n6998), .ZN(P2_U3344) );
  OR2_X1 U8735 ( .A1(n6999), .A2(P2_U3152), .ZN(n7000) );
  OAI211_X1 U8736 ( .C1(n9830), .C2(n7002), .A(n7001), .B(n7000), .ZN(n7003)
         );
  NAND2_X1 U8737 ( .A1(n7003), .A2(n4254), .ZN(n7007) );
  NAND2_X1 U8738 ( .A1(n7007), .A2(n8464), .ZN(n7015) );
  NAND2_X1 U8739 ( .A1(n7015), .A2(n7004), .ZN(n9805) );
  INV_X1 U8740 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7114) );
  NOR2_X1 U8741 ( .A1(n7114), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7013) );
  NAND2_X1 U8742 ( .A1(n9813), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7011) );
  MUX2_X1 U8743 ( .A(n4986), .B(P2_REG1_REG_1__SCAN_IN), .S(n7020), .Z(n7006)
         );
  INV_X1 U8744 ( .A(n7006), .ZN(n7010) );
  INV_X1 U8745 ( .A(n7011), .ZN(n7005) );
  NAND2_X1 U8746 ( .A1(n7006), .A2(n7005), .ZN(n7025) );
  INV_X1 U8747 ( .A(n7025), .ZN(n7009) );
  INV_X1 U8748 ( .A(n7007), .ZN(n7008) );
  NAND2_X1 U8749 ( .A1(n7008), .A2(n9030), .ZN(n9807) );
  AOI211_X1 U8750 ( .C1(n7011), .C2(n7010), .A(n7009), .B(n9807), .ZN(n7012)
         );
  AOI211_X1 U8751 ( .C1(P2_ADDR_REG_1__SCAN_IN), .C2(n9817), .A(n7013), .B(
        n7012), .ZN(n7019) );
  AND2_X1 U8752 ( .A1(n9813), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7017) );
  INV_X1 U8753 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7122) );
  NAND2_X1 U8754 ( .A1(n7015), .A2(n7014), .ZN(n9827) );
  OAI211_X1 U8755 ( .C1(n7017), .C2(n7016), .A(n8579), .B(n7034), .ZN(n7018)
         );
  OAI211_X1 U8756 ( .C1(n9805), .C2(n7020), .A(n7019), .B(n7018), .ZN(P2_U3246) );
  OAI222_X1 U8757 ( .A1(n7855), .A2(n7023), .B1(n10109), .B2(n7022), .C1(n7021), .C2(P1_U3084), .ZN(P1_U3339) );
  INV_X1 U8758 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7225) );
  MUX2_X1 U8759 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5020), .S(n7039), .Z(n7027)
         );
  NAND2_X1 U8760 ( .A1(n7031), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7024) );
  NAND2_X1 U8761 ( .A1(n7025), .A2(n7024), .ZN(n7026) );
  NAND2_X1 U8762 ( .A1(n7026), .A2(n7027), .ZN(n7041) );
  OAI211_X1 U8763 ( .C1(n7027), .C2(n7026), .A(n9823), .B(n7041), .ZN(n7029)
         );
  NAND2_X1 U8764 ( .A1(n9817), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n7028) );
  OAI211_X1 U8765 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7225), .A(n7029), .B(n7028), .ZN(n7030) );
  AOI21_X1 U8766 ( .B1(n7039), .B2(n9821), .A(n7030), .ZN(n7038) );
  NAND2_X1 U8767 ( .A1(n7031), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7033) );
  MUX2_X1 U8768 ( .A(n7231), .B(P2_REG2_REG_2__SCAN_IN), .S(n7039), .Z(n7032)
         );
  INV_X1 U8769 ( .A(n8468), .ZN(n7036) );
  NAND3_X1 U8770 ( .A1(n7034), .A2(n7033), .A3(n7032), .ZN(n7035) );
  NAND3_X1 U8771 ( .A1(n8579), .A2(n7036), .A3(n7035), .ZN(n7037) );
  NAND2_X1 U8772 ( .A1(n7038), .A2(n7037), .ZN(P2_U3247) );
  XNOR2_X1 U8773 ( .A(n7071), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7056) );
  NAND2_X1 U8774 ( .A1(n7039), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7040) );
  NAND2_X1 U8775 ( .A1(n7041), .A2(n7040), .ZN(n8473) );
  XNOR2_X1 U8776 ( .A(n7058), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n8474) );
  NAND2_X1 U8777 ( .A1(n8473), .A2(n8474), .ZN(n8472) );
  INV_X1 U8778 ( .A(n7058), .ZN(n8471) );
  NAND2_X1 U8779 ( .A1(n8471), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7042) );
  NAND2_X1 U8780 ( .A1(n8472), .A2(n7042), .ZN(n8488) );
  MUX2_X1 U8781 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n5063), .S(n8486), .Z(n8489)
         );
  NAND2_X1 U8782 ( .A1(n8488), .A2(n8489), .ZN(n8487) );
  NAND2_X1 U8783 ( .A1(n8486), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7043) );
  NAND2_X1 U8784 ( .A1(n8487), .A2(n7043), .ZN(n8501) );
  MUX2_X1 U8785 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n5092), .S(n8499), .Z(n8502)
         );
  NAND2_X1 U8786 ( .A1(n8501), .A2(n8502), .ZN(n8500) );
  NAND2_X1 U8787 ( .A1(n8499), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7044) );
  NAND2_X1 U8788 ( .A1(n8500), .A2(n7044), .ZN(n8516) );
  XNOR2_X1 U8789 ( .A(n8514), .B(n7045), .ZN(n8517) );
  NAND2_X1 U8790 ( .A1(n8516), .A2(n8517), .ZN(n8515) );
  NAND2_X1 U8791 ( .A1(n8514), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7046) );
  NAND2_X1 U8792 ( .A1(n8515), .A2(n7046), .ZN(n8532) );
  MUX2_X1 U8793 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n5129), .S(n8528), .Z(n8533)
         );
  NAND2_X1 U8794 ( .A1(n8532), .A2(n8533), .ZN(n8531) );
  NAND2_X1 U8795 ( .A1(n8528), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U8796 ( .A1(n8531), .A2(n7047), .ZN(n8542) );
  MUX2_X1 U8797 ( .A(n5156), .B(P2_REG1_REG_8__SCAN_IN), .S(n8538), .Z(n8543)
         );
  NAND2_X1 U8798 ( .A1(n7048), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7049) );
  NAND2_X1 U8799 ( .A1(n8541), .A2(n7049), .ZN(n8560) );
  MUX2_X1 U8800 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n5173), .S(n8562), .Z(n8561)
         );
  NAND2_X1 U8801 ( .A1(n8560), .A2(n8561), .ZN(n8559) );
  NAND2_X1 U8802 ( .A1(n8562), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7050) );
  NAND2_X1 U8803 ( .A1(n8559), .A2(n7050), .ZN(n7083) );
  INV_X1 U8804 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9924) );
  MUX2_X1 U8805 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9924), .S(n7064), .Z(n7082)
         );
  NAND2_X1 U8806 ( .A1(n7083), .A2(n7082), .ZN(n7081) );
  NAND2_X1 U8807 ( .A1(n7064), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7051) );
  NAND2_X1 U8808 ( .A1(n7081), .A2(n7051), .ZN(n7098) );
  XNOR2_X1 U8809 ( .A(n7065), .B(n7052), .ZN(n7097) );
  NAND2_X1 U8810 ( .A1(n7098), .A2(n7097), .ZN(n7096) );
  NAND2_X1 U8811 ( .A1(n7065), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7053) );
  NAND2_X1 U8812 ( .A1(n7096), .A2(n7053), .ZN(n7055) );
  INV_X1 U8813 ( .A(n7154), .ZN(n7054) );
  AOI21_X1 U8814 ( .B1(n7056), .B2(n7055), .A(n7054), .ZN(n7074) );
  NOR2_X1 U8815 ( .A1(n7057), .A2(n7231), .ZN(n8466) );
  MUX2_X1 U8816 ( .A(n7059), .B(P2_REG2_REG_3__SCAN_IN), .S(n7058), .Z(n8467)
         );
  NAND2_X1 U8817 ( .A1(n8471), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8480) );
  MUX2_X1 U8818 ( .A(n5064), .B(P2_REG2_REG_4__SCAN_IN), .S(n8486), .Z(n8479)
         );
  NOR2_X1 U8819 ( .A1(n7060), .A2(n5064), .ZN(n8495) );
  MUX2_X1 U8820 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7475), .S(n8499), .Z(n8494)
         );
  OAI21_X1 U8821 ( .B1(n8496), .B2(n8495), .A(n8494), .ZN(n8509) );
  NAND2_X1 U8822 ( .A1(n8499), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8508) );
  MUX2_X1 U8823 ( .A(n7507), .B(P2_REG2_REG_6__SCAN_IN), .S(n8514), .Z(n8507)
         );
  NOR2_X1 U8824 ( .A1(n7061), .A2(n7507), .ZN(n8523) );
  MUX2_X1 U8825 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7062), .S(n8528), .Z(n8522)
         );
  NAND2_X1 U8826 ( .A1(n8528), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8545) );
  MUX2_X1 U8827 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n5150), .S(n8538), .Z(n8544)
         );
  AOI21_X1 U8828 ( .B1(n8546), .B2(n8545), .A(n8544), .ZN(n8554) );
  NOR2_X1 U8829 ( .A1(n8538), .A2(n5150), .ZN(n8553) );
  MUX2_X1 U8830 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7063), .S(n8562), .Z(n8552)
         );
  OAI21_X1 U8831 ( .B1(n8554), .B2(n8553), .A(n8552), .ZN(n8556) );
  NAND2_X1 U8832 ( .A1(n8562), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7076) );
  MUX2_X1 U8833 ( .A(n5201), .B(P2_REG2_REG_10__SCAN_IN), .S(n7064), .Z(n7075)
         );
  AOI21_X1 U8834 ( .B1(n7064), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7087), .ZN(
        n7088) );
  MUX2_X1 U8835 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n5220), .S(n7065), .Z(n7089)
         );
  NOR2_X1 U8836 ( .A1(n7065), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7066) );
  MUX2_X1 U8837 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8112), .S(n7071), .Z(n7067)
         );
  INV_X1 U8838 ( .A(n7163), .ZN(n7069) );
  NOR3_X1 U8839 ( .A1(n7090), .A2(n7067), .A3(n7066), .ZN(n7068) );
  OAI21_X1 U8840 ( .B1(n7069), .B2(n7068), .A(n8579), .ZN(n7073) );
  INV_X1 U8841 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U8842 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8003) );
  OAI21_X1 U8843 ( .B1(n8585), .B2(n9987), .A(n8003), .ZN(n7070) );
  AOI21_X1 U8844 ( .B1(n9821), .B2(n7071), .A(n7070), .ZN(n7072) );
  OAI211_X1 U8845 ( .C1(n7074), .C2(n9807), .A(n7073), .B(n7072), .ZN(P2_U3257) );
  NAND3_X1 U8846 ( .A1(n8556), .A2(n7076), .A3(n7075), .ZN(n7077) );
  NAND2_X1 U8847 ( .A1(n7077), .A2(n8579), .ZN(n7086) );
  NAND2_X1 U8848 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7831) );
  INV_X1 U8849 ( .A(n7831), .ZN(n7080) );
  NOR2_X1 U8850 ( .A1(n9805), .A2(n7078), .ZN(n7079) );
  AOI211_X1 U8851 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n9817), .A(n7080), .B(
        n7079), .ZN(n7085) );
  OAI211_X1 U8852 ( .C1(n7083), .C2(n7082), .A(n7081), .B(n9823), .ZN(n7084)
         );
  OAI211_X1 U8853 ( .C1(n7087), .C2(n7086), .A(n7085), .B(n7084), .ZN(P2_U3255) );
  INV_X1 U8854 ( .A(n7088), .ZN(n7092) );
  INV_X1 U8855 ( .A(n7089), .ZN(n7091) );
  AOI21_X1 U8856 ( .B1(n7092), .B2(n7091), .A(n7090), .ZN(n7101) );
  NOR2_X1 U8857 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7916), .ZN(n7095) );
  NOR2_X1 U8858 ( .A1(n9805), .A2(n7093), .ZN(n7094) );
  AOI211_X1 U8859 ( .C1(P2_ADDR_REG_11__SCAN_IN), .C2(n9817), .A(n7095), .B(
        n7094), .ZN(n7100) );
  OAI211_X1 U8860 ( .C1(n7098), .C2(n7097), .A(n7096), .B(n9823), .ZN(n7099)
         );
  OAI211_X1 U8861 ( .C1(n7101), .C2(n9827), .A(n7100), .B(n7099), .ZN(P2_U3256) );
  XNOR2_X1 U8862 ( .A(n7198), .B(n7102), .ZN(n9844) );
  NAND2_X1 U8863 ( .A1(n7625), .A2(n7636), .ZN(n7106) );
  NOR2_X1 U8864 ( .A1(n9830), .A2(n7103), .ZN(n7104) );
  NAND2_X1 U8865 ( .A1(n7105), .A2(n7104), .ZN(n7623) );
  XNOR2_X1 U8866 ( .A(n7108), .B(n5637), .ZN(n7107) );
  NAND2_X1 U8867 ( .A1(n7107), .A2(n8758), .ZN(n8867) );
  NAND2_X1 U8868 ( .A1(n7108), .A2(n7627), .ZN(n7373) );
  NAND2_X1 U8869 ( .A1(n8867), .A2(n7373), .ZN(n7109) );
  INV_X1 U8870 ( .A(n7110), .ZN(n7111) );
  NOR2_X2 U8871 ( .A1(n8289), .A2(n9839), .ZN(n7223) );
  INV_X1 U8872 ( .A(n7223), .ZN(n9847) );
  NAND2_X1 U8873 ( .A1(n8289), .A2(n9839), .ZN(n9845) );
  NAND2_X1 U8874 ( .A1(n9847), .A2(n9845), .ZN(n7115) );
  OAI22_X1 U8875 ( .A1(n8687), .A2(n7115), .B1(n7114), .B2(n8761), .ZN(n7116)
         );
  AOI21_X1 U8876 ( .B1(n8765), .B2(n8289), .A(n7116), .ZN(n7124) );
  XNOR2_X1 U8877 ( .A(n7198), .B(n7119), .ZN(n7121) );
  AOI222_X1 U8878 ( .A1(n8871), .A2(n7121), .B1(n8465), .B2(n8819), .C1(n7120), 
        .C2(n8817), .ZN(n9849) );
  MUX2_X1 U8879 ( .A(n7122), .B(n9849), .S(n8772), .Z(n7123) );
  OAI211_X1 U8880 ( .C1(n9844), .C2(n8854), .A(n7124), .B(n7123), .ZN(P2_U3295) );
  INV_X1 U8881 ( .A(n7125), .ZN(n7128) );
  OAI222_X1 U8882 ( .A1(n7855), .A2(n7127), .B1(n10109), .B2(n7128), .C1(
        P1_U3084), .C2(n7126), .ZN(P1_U3338) );
  OAI222_X1 U8883 ( .A1(n9040), .A2(n7129), .B1(n9038), .B2(n7128), .C1(
        P2_U3152), .C2(n4454), .ZN(P2_U3343) );
  INV_X1 U8884 ( .A(n9632), .ZN(n9794) );
  NAND2_X1 U8885 ( .A1(n9201), .A2(n7462), .ZN(n7258) );
  NOR2_X1 U8886 ( .A1(n7267), .A2(n7258), .ZN(n7259) );
  AOI21_X1 U8887 ( .B1(n9724), .B2(n6587), .A(n7259), .ZN(n7132) );
  NAND2_X1 U8888 ( .A1(n7258), .A2(n6080), .ZN(n7130) );
  NAND2_X1 U8889 ( .A1(n7130), .A2(n9724), .ZN(n7131) );
  OAI211_X1 U8890 ( .C1(n7258), .C2(n6080), .A(n7136), .B(n7131), .ZN(n7439)
         );
  OAI21_X1 U8891 ( .B1(n7132), .B2(n7136), .A(n7439), .ZN(n7590) );
  NOR2_X2 U8892 ( .A1(n9724), .A2(n7462), .ZN(n7263) );
  NAND2_X1 U8893 ( .A1(n7263), .A2(n6093), .ZN(n7445) );
  OAI21_X1 U8894 ( .B1(n7263), .B2(n6093), .A(n7445), .ZN(n7586) );
  OAI22_X1 U8895 ( .A1(n9787), .A2(n6093), .B1(n9789), .B2(n7586), .ZN(n7147)
         );
  NAND2_X1 U8896 ( .A1(n6530), .A2(n9278), .ZN(n7135) );
  NAND2_X1 U8897 ( .A1(n4259), .A2(n7133), .ZN(n7134) );
  INV_X1 U8898 ( .A(n9509), .ZN(n7743) );
  XNOR2_X1 U8899 ( .A(n7137), .B(n7136), .ZN(n7146) );
  OR2_X1 U8900 ( .A1(n7138), .A2(n7517), .ZN(n7141) );
  NAND3_X1 U8901 ( .A1(n6508), .A2(n4259), .A3(n7139), .ZN(n7140) );
  INV_X1 U8902 ( .A(n9480), .ZN(n7894) );
  NAND2_X1 U8903 ( .A1(n7590), .A2(n7894), .ZN(n7145) );
  INV_X1 U8904 ( .A(n7142), .ZN(n7143) );
  AOI22_X1 U8905 ( .A1(n9510), .A2(n7530), .B1(n9506), .B2(n6587), .ZN(n7144)
         );
  OAI211_X1 U8906 ( .C1(n7743), .C2(n7146), .A(n7145), .B(n7144), .ZN(n7584)
         );
  AOI211_X1 U8907 ( .C1(n9794), .C2(n7590), .A(n7147), .B(n7584), .ZN(n9772)
         );
  OAI21_X1 U8908 ( .B1(n9632), .B2(n4259), .A(n7451), .ZN(n7149) );
  NAND2_X1 U8909 ( .A1(n9799), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7151) );
  OAI21_X1 U8910 ( .B1(n9772), .B2(n9799), .A(n7151), .ZN(P1_U3525) );
  XNOR2_X1 U8911 ( .A(n7211), .B(n9993), .ZN(n7156) );
  NAND2_X1 U8912 ( .A1(n7159), .A2(n7152), .ZN(n7153) );
  NAND2_X1 U8913 ( .A1(n7155), .A2(n7156), .ZN(n7210) );
  OAI21_X1 U8914 ( .B1(n7156), .B2(n7155), .A(n7210), .ZN(n7168) );
  NAND2_X1 U8915 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8067) );
  NAND2_X1 U8916 ( .A1(n9817), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n7157) );
  OAI211_X1 U8917 ( .C1(n9805), .C2(n7158), .A(n8067), .B(n7157), .ZN(n7167)
         );
  NAND2_X1 U8918 ( .A1(n7159), .A2(n8112), .ZN(n7161) );
  MUX2_X1 U8919 ( .A(n7160), .B(P2_REG2_REG_13__SCAN_IN), .S(n7211), .Z(n7162)
         );
  INV_X1 U8920 ( .A(n7214), .ZN(n7165) );
  NAND3_X1 U8921 ( .A1(n7163), .A2(n7162), .A3(n7161), .ZN(n7164) );
  AOI21_X1 U8922 ( .B1(n7165), .B2(n7164), .A(n9827), .ZN(n7166) );
  AOI211_X1 U8923 ( .C1(n9823), .C2(n7168), .A(n7167), .B(n7166), .ZN(n7169)
         );
  INV_X1 U8924 ( .A(n7169), .ZN(P2_U3258) );
  INV_X1 U8925 ( .A(n7170), .ZN(n7171) );
  NOR2_X1 U8926 ( .A1(n7172), .A2(n7171), .ZN(n7173) );
  XNOR2_X1 U8927 ( .A(n7174), .B(n7173), .ZN(n7183) );
  OAI21_X1 U8928 ( .B1(n7177), .B2(n7176), .A(n7175), .ZN(n7179) );
  AOI22_X1 U8929 ( .A1(n7179), .A2(n9709), .B1(n7178), .B2(n9711), .ZN(n7182)
         );
  NOR2_X1 U8930 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7180), .ZN(n7907) );
  AOI21_X1 U8931 ( .B1(n9718), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7907), .ZN(
        n7181) );
  OAI211_X1 U8932 ( .C1(n9254), .C2(n7183), .A(n7182), .B(n7181), .ZN(P1_U3249) );
  XOR2_X1 U8933 ( .A(n7185), .B(n7184), .Z(n7191) );
  AOI22_X1 U8934 ( .A1(n9155), .A2(n6587), .B1(n9180), .B2(n7530), .ZN(n7190)
         );
  INV_X1 U8935 ( .A(n7454), .ZN(n7187) );
  NAND3_X1 U8936 ( .A1(n7188), .A2(n7187), .A3(n7186), .ZN(n7357) );
  AOI22_X1 U8937 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n7357), .B1(n9184), .B2(
        n7589), .ZN(n7189) );
  OAI211_X1 U8938 ( .C1(n7191), .C2(n9186), .A(n7190), .B(n7189), .ZN(P1_U3235) );
  XNOR2_X1 U8939 ( .A(n7192), .B(n7466), .ZN(n7194) );
  OAI222_X1 U8940 ( .A1(n8859), .A2(n7578), .B1(n8861), .B2(n7203), .C1(n7194), 
        .C2(n8831), .ZN(n9870) );
  INV_X1 U8941 ( .A(n9870), .ZN(n7207) );
  NOR2_X1 U8942 ( .A1(n8772), .A2(n5064), .ZN(n7196) );
  XNOR2_X1 U8943 ( .A(n7478), .B(n7477), .ZN(n9869) );
  OAI22_X1 U8944 ( .A1(n8687), .A2(n9869), .B1(n7579), .B2(n8761), .ZN(n7195)
         );
  AOI211_X1 U8945 ( .C1(n8765), .C2(n7477), .A(n7196), .B(n7195), .ZN(n7206)
         );
  INV_X1 U8946 ( .A(n8854), .ZN(n8811) );
  NAND2_X1 U8947 ( .A1(n5812), .A2(n7199), .ZN(n7200) );
  NAND2_X1 U8948 ( .A1(n8282), .A2(n9853), .ZN(n7202) );
  XNOR2_X1 U8949 ( .A(n7467), .B(n7466), .ZN(n9872) );
  NAND2_X1 U8950 ( .A1(n8811), .A2(n9872), .ZN(n7205) );
  OAI211_X1 U8951 ( .C1(n7207), .C2(n8886), .A(n7206), .B(n7205), .ZN(P2_U3292) );
  XNOR2_X1 U8952 ( .A(n7491), .B(n7208), .ZN(n7493) );
  OR2_X1 U8953 ( .A1(n7211), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7209) );
  XOR2_X1 U8954 ( .A(n7493), .B(n7494), .Z(n7221) );
  NOR2_X1 U8955 ( .A1(n7211), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7212) );
  MUX2_X1 U8956 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n5268), .S(n7491), .Z(n7213)
         );
  INV_X1 U8957 ( .A(n7487), .ZN(n7216) );
  NOR3_X1 U8958 ( .A1(n7214), .A2(n7213), .A3(n7212), .ZN(n7215) );
  OAI21_X1 U8959 ( .B1(n7216), .B2(n7215), .A(n8579), .ZN(n7220) );
  AND2_X1 U8960 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8317) );
  INV_X1 U8961 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7217) );
  NOR2_X1 U8962 ( .A1(n8585), .A2(n7217), .ZN(n7218) );
  AOI211_X1 U8963 ( .C1(n9821), .C2(n7491), .A(n8317), .B(n7218), .ZN(n7219)
         );
  OAI211_X1 U8964 ( .C1(n7221), .C2(n9807), .A(n7220), .B(n7219), .ZN(P2_U3259) );
  XNOR2_X1 U8965 ( .A(n7201), .B(n7222), .ZN(n9858) );
  OR2_X1 U8966 ( .A1(n7223), .A2(n9853), .ZN(n7224) );
  OAI22_X1 U8967 ( .A1(n8687), .A2(n9854), .B1(n7225), .B2(n8761), .ZN(n7226)
         );
  AOI21_X1 U8968 ( .B1(n8811), .B2(n9858), .A(n7226), .ZN(n7233) );
  OAI21_X1 U8969 ( .B1(n7228), .B2(n7227), .A(n7364), .ZN(n7230) );
  AOI222_X1 U8970 ( .A1(n8871), .A2(n7230), .B1(n8463), .B2(n8817), .C1(n7229), 
        .C2(n8819), .ZN(n9855) );
  MUX2_X1 U8971 ( .A(n7231), .B(n9855), .S(n8772), .Z(n7232) );
  OAI211_X1 U8972 ( .C1(n9853), .C2(n8879), .A(n7233), .B(n7232), .ZN(P2_U3294) );
  OAI211_X1 U8973 ( .C1(n7236), .C2(n7235), .A(n9719), .B(n7234), .ZN(n7237)
         );
  OAI21_X1 U8974 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6065), .A(n7237), .ZN(n7238) );
  AOI21_X1 U8975 ( .B1(n9718), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n7238), .ZN(
        n7243) );
  OAI211_X1 U8976 ( .C1(n7241), .C2(n7240), .A(n9709), .B(n7239), .ZN(n7242)
         );
  OAI211_X1 U8977 ( .C1(n9261), .C2(n7244), .A(n7243), .B(n7242), .ZN(P1_U3242) );
  OAI21_X1 U8978 ( .B1(n7247), .B2(n7246), .A(n7245), .ZN(n7250) );
  AND2_X1 U8979 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7685) );
  INV_X1 U8980 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7248) );
  NOR2_X1 U8981 ( .A1(n9281), .A2(n7248), .ZN(n7249) );
  AOI211_X1 U8982 ( .C1(n9709), .C2(n7250), .A(n7685), .B(n7249), .ZN(n7256)
         );
  AND3_X1 U8983 ( .A1(n9218), .A2(n7252), .A3(n7251), .ZN(n7253) );
  OAI21_X1 U8984 ( .B1(n7254), .B2(n7253), .A(n9719), .ZN(n7255) );
  OAI211_X1 U8985 ( .C1(n9261), .C2(n7257), .A(n7256), .B(n7255), .ZN(P1_U3248) );
  INV_X1 U8986 ( .A(n7267), .ZN(n7262) );
  INV_X1 U8987 ( .A(n7258), .ZN(n7261) );
  INV_X1 U8988 ( .A(n7259), .ZN(n7260) );
  OAI21_X1 U8989 ( .B1(n7262), .B2(n7261), .A(n7260), .ZN(n7272) );
  INV_X1 U8990 ( .A(n7272), .ZN(n9731) );
  INV_X1 U8991 ( .A(n7263), .ZN(n7264) );
  OAI211_X1 U8992 ( .C1(n7265), .C2(n7701), .A(n9627), .B(n7264), .ZN(n9723)
         );
  OAI21_X1 U8993 ( .B1(n9787), .B2(n7265), .A(n9723), .ZN(n7273) );
  AOI22_X1 U8994 ( .A1(n9510), .A2(n9199), .B1(n9506), .B2(n9201), .ZN(n7271)
         );
  OAI21_X1 U8995 ( .B1(n7268), .B2(n7267), .A(n7266), .ZN(n7269) );
  NAND2_X1 U8996 ( .A1(n7269), .A2(n9509), .ZN(n7270) );
  OAI211_X1 U8997 ( .C1(n7272), .C2(n9480), .A(n7271), .B(n7270), .ZN(n9730)
         );
  AOI211_X1 U8998 ( .C1(n9794), .C2(n9731), .A(n7273), .B(n9730), .ZN(n7697)
         );
  NAND2_X1 U8999 ( .A1(n9799), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7274) );
  OAI21_X1 U9000 ( .B1(n7697), .B2(n9799), .A(n7274), .ZN(P1_U3524) );
  INV_X1 U9001 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7465) );
  NAND2_X1 U9002 ( .A1(n9672), .A2(n7465), .ZN(n7275) );
  NAND2_X1 U9003 ( .A1(n9669), .A2(n7275), .ZN(n7279) );
  INV_X1 U9004 ( .A(n7279), .ZN(n7278) );
  OAI21_X1 U9005 ( .B1(n9672), .B2(P1_REG1_REG_0__SCAN_IN), .A(n4650), .ZN(
        n7277) );
  AOI21_X1 U9006 ( .B1(n7278), .B2(n7277), .A(n7276), .ZN(n7280) );
  NAND2_X1 U9007 ( .A1(n7279), .A2(n4650), .ZN(n7409) );
  NAND3_X1 U9008 ( .A1(n7281), .A2(n7280), .A3(n7409), .ZN(n7282) );
  OAI21_X1 U9009 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6070), .A(n7282), .ZN(n7284) );
  NOR3_X1 U9010 ( .A1(n9254), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n4650), .ZN(
        n7283) );
  AOI211_X1 U9011 ( .C1(n9718), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n7284), .B(
        n7283), .ZN(n7285) );
  INV_X1 U9012 ( .A(n7285), .ZN(P1_U3241) );
  INV_X1 U9013 ( .A(n7286), .ZN(n7289) );
  OAI222_X1 U9014 ( .A1(n9040), .A2(n7287), .B1(n9038), .B2(n7289), .C1(n7921), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U9015 ( .A(n7288), .ZN(n9260) );
  OAI222_X1 U9016 ( .A1(n7855), .A2(n7290), .B1(n10109), .B2(n7289), .C1(n9260), .C2(P1_U3084), .ZN(P1_U3337) );
  XOR2_X1 U9017 ( .A(n7292), .B(n7291), .Z(n7302) );
  OAI21_X1 U9018 ( .B1(n7295), .B2(n7294), .A(n7293), .ZN(n7300) );
  INV_X1 U9019 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7298) );
  NAND2_X1 U9020 ( .A1(n9711), .A2(n7296), .ZN(n7297) );
  NAND2_X1 U9021 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8010) );
  OAI211_X1 U9022 ( .C1(n9281), .C2(n7298), .A(n7297), .B(n8010), .ZN(n7299)
         );
  AOI21_X1 U9023 ( .B1(n7300), .B2(n9709), .A(n7299), .ZN(n7301) );
  OAI21_X1 U9024 ( .B1(n9254), .B2(n7302), .A(n7301), .ZN(P1_U3252) );
  INV_X1 U9025 ( .A(n7357), .ZN(n7307) );
  NAND2_X1 U9026 ( .A1(n7407), .A2(n9165), .ZN(n7306) );
  AOI22_X1 U9027 ( .A1(n7462), .A2(n9184), .B1(n9180), .B2(n6587), .ZN(n7305)
         );
  OAI211_X1 U9028 ( .C1(n7307), .C2(n6070), .A(n7306), .B(n7305), .ZN(P1_U3230) );
  XNOR2_X1 U9029 ( .A(n7309), .B(n7308), .ZN(n7310) );
  NAND2_X1 U9030 ( .A1(n7310), .A2(n9165), .ZN(n7313) );
  NOR2_X1 U9031 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6095), .ZN(n7388) );
  OAI22_X1 U9032 ( .A1(n7521), .A2(n9173), .B1(n9178), .B2(n7440), .ZN(n7311)
         );
  AOI211_X1 U9033 ( .C1(n9180), .C2(n9198), .A(n7388), .B(n7311), .ZN(n7312)
         );
  OAI211_X1 U9034 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9182), .A(n7313), .B(
        n7312), .ZN(P1_U3216) );
  NAND2_X1 U9035 ( .A1(n7315), .A2(n7314), .ZN(n7320) );
  XOR2_X1 U9036 ( .A(n7318), .B(n7316), .Z(n8285) );
  NOR2_X1 U9037 ( .A1(n8285), .A2(n8284), .ZN(n8283) );
  AOI21_X1 U9038 ( .B1(n7318), .B2(n5814), .A(n8283), .ZN(n7319) );
  XOR2_X1 U9039 ( .A(n7320), .B(n7319), .Z(n7325) );
  INV_X1 U9040 ( .A(n7330), .ZN(n7321) );
  NAND2_X1 U9041 ( .A1(n7321), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8288) );
  AOI22_X1 U9042 ( .A1(n8288), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n8445), .B2(
        n7322), .ZN(n7324) );
  INV_X1 U9043 ( .A(n8440), .ZN(n7598) );
  INV_X1 U9044 ( .A(n8441), .ZN(n8290) );
  AOI22_X1 U9045 ( .A1(n7598), .A2(n7229), .B1(n8290), .B2(n8463), .ZN(n7323)
         );
  OAI211_X1 U9046 ( .C1(n7325), .C2(n8447), .A(n7324), .B(n7323), .ZN(P2_U3239) );
  OAI21_X1 U9047 ( .B1(n8293), .B2(n7328), .A(n7327), .ZN(n7329) );
  NAND2_X1 U9048 ( .A1(n7326), .A2(n7329), .ZN(n7333) );
  AOI22_X1 U9049 ( .A1(n8290), .A2(n7229), .B1(n9839), .B2(n8445), .ZN(n7332)
         );
  AND2_X1 U9050 ( .A1(P2_U3152), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9809) );
  AOI21_X1 U9051 ( .B1(n7330), .B2(P2_REG3_REG_0__SCAN_IN), .A(n9809), .ZN(
        n7331) );
  OAI211_X1 U9052 ( .C1(n8447), .C2(n7333), .A(n7332), .B(n7331), .ZN(P2_U3234) );
  XNOR2_X1 U9053 ( .A(n7335), .B(n7334), .ZN(n7340) );
  INV_X1 U9054 ( .A(n8426), .ZN(n8376) );
  AOI22_X1 U9055 ( .A1(n8819), .A2(n8462), .B1(n8460), .B2(n8817), .ZN(n7473)
         );
  INV_X1 U9056 ( .A(n7473), .ZN(n7336) );
  AOI22_X1 U9057 ( .A1(n8376), .A2(n7336), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n7339) );
  INV_X1 U9058 ( .A(n7481), .ZN(n7337) );
  AOI22_X1 U9059 ( .A1(n7337), .A2(n8429), .B1(n8445), .B2(n7631), .ZN(n7338)
         );
  OAI211_X1 U9060 ( .C1(n7340), .C2(n8447), .A(n7339), .B(n7338), .ZN(P2_U3229) );
  INV_X1 U9061 ( .A(n7341), .ZN(n7436) );
  AOI22_X1 U9062 ( .A1(n9272), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10113), .ZN(n7342) );
  OAI21_X1 U9063 ( .B1(n7436), .B2(n10109), .A(n7342), .ZN(P1_U3336) );
  AND2_X1 U9064 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7760) );
  XOR2_X1 U9065 ( .A(n7344), .B(n7343), .Z(n7345) );
  NOR2_X1 U9066 ( .A1(n9251), .A2(n7345), .ZN(n7346) );
  AOI211_X1 U9067 ( .C1(n9718), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n7760), .B(
        n7346), .ZN(n7351) );
  OAI211_X1 U9068 ( .C1(n7349), .C2(n7348), .A(n9719), .B(n7347), .ZN(n7350)
         );
  OAI211_X1 U9069 ( .C1(n9261), .C2(n7352), .A(n7351), .B(n7350), .ZN(P1_U3246) );
  XNOR2_X1 U9070 ( .A(n7354), .B(n7353), .ZN(n7355) );
  XNOR2_X1 U9071 ( .A(n7356), .B(n7355), .ZN(n7360) );
  AOI22_X1 U9072 ( .A1(n9180), .A2(n9199), .B1(n9155), .B2(n9201), .ZN(n7359)
         );
  AOI22_X1 U9073 ( .A1(n7357), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n9184), .B2(
        n9724), .ZN(n7358) );
  OAI211_X1 U9074 ( .C1(n7360), .C2(n9186), .A(n7359), .B(n7358), .ZN(P1_U3220) );
  XNOR2_X1 U9075 ( .A(n7361), .B(n4260), .ZN(n7375) );
  INV_X1 U9076 ( .A(n7375), .ZN(n9864) );
  INV_X1 U9077 ( .A(n8867), .ZN(n8087) );
  NAND2_X1 U9078 ( .A1(n9864), .A2(n8087), .ZN(n7371) );
  NAND3_X1 U9079 ( .A1(n7364), .A2(n7363), .A3(n7362), .ZN(n7365) );
  NAND2_X1 U9080 ( .A1(n7366), .A2(n7365), .ZN(n7369) );
  NAND2_X1 U9081 ( .A1(n8462), .A2(n8817), .ZN(n7367) );
  OAI21_X1 U9082 ( .B1(n8282), .B2(n8861), .A(n7367), .ZN(n7368) );
  AOI21_X1 U9083 ( .B1(n7369), .B2(n8871), .A(n7368), .ZN(n7370) );
  AND2_X1 U9084 ( .A1(n7371), .A2(n7370), .ZN(n9865) );
  NAND2_X1 U9085 ( .A1(n7478), .A2(n7372), .ZN(n9862) );
  OAI22_X1 U9086 ( .A1(n8687), .A2(n9862), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8761), .ZN(n7377) );
  INV_X1 U9087 ( .A(n7373), .ZN(n7374) );
  NAND2_X1 U9088 ( .A1(n8772), .A2(n7374), .ZN(n8881) );
  OAI22_X1 U9089 ( .A1(n8879), .A2(n9861), .B1(n7375), .B2(n8881), .ZN(n7376)
         );
  AOI211_X1 U9090 ( .C1(n8886), .C2(P2_REG2_REG_3__SCAN_IN), .A(n7377), .B(
        n7376), .ZN(n7378) );
  OAI21_X1 U9091 ( .B1(n8886), .B2(n9865), .A(n7378), .ZN(P2_U3293) );
  INV_X1 U9092 ( .A(n9840), .ZN(n7383) );
  AOI22_X1 U9093 ( .A1(n9840), .A2(n8871), .B1(n8817), .B2(n7229), .ZN(n9842)
         );
  OAI22_X1 U9094 ( .A1(n8886), .A2(n9842), .B1(n7379), .B2(n8761), .ZN(n7380)
         );
  AOI21_X1 U9095 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n8886), .A(n7380), .ZN(
        n7382) );
  OAI21_X1 U9096 ( .B1(n8765), .B2(n8884), .A(n9839), .ZN(n7381) );
  OAI211_X1 U9097 ( .C1(n7383), .C2(n8854), .A(n7382), .B(n7381), .ZN(P2_U3296) );
  AOI211_X1 U9098 ( .C1(n7386), .C2(n7385), .A(n7384), .B(n9251), .ZN(n7387)
         );
  AOI211_X1 U9099 ( .C1(n9718), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n7388), .B(
        n7387), .ZN(n7393) );
  OAI211_X1 U9100 ( .C1(n7391), .C2(n7390), .A(n9719), .B(n7389), .ZN(n7392)
         );
  OAI211_X1 U9101 ( .C1(n9261), .C2(n7394), .A(n7393), .B(n7392), .ZN(P1_U3244) );
  INV_X1 U9102 ( .A(n7395), .ZN(n7398) );
  MUX2_X1 U9103 ( .A(n6911), .B(P1_REG1_REG_4__SCAN_IN), .S(n7403), .Z(n7397)
         );
  OAI21_X1 U9104 ( .B1(n7398), .B2(n7397), .A(n7396), .ZN(n7406) );
  INV_X1 U9105 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n7399) );
  NAND2_X1 U9106 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n7668) );
  OAI21_X1 U9107 ( .B1(n9281), .B2(n7399), .A(n7668), .ZN(n7405) );
  XNOR2_X1 U9108 ( .A(n7401), .B(n7400), .ZN(n7402) );
  OAI22_X1 U9109 ( .A1(n7403), .A2(n9261), .B1(n9251), .B2(n7402), .ZN(n7404)
         );
  AOI211_X1 U9110 ( .C1(n9719), .C2(n7406), .A(n7405), .B(n7404), .ZN(n7412)
         );
  MUX2_X1 U9111 ( .A(n7408), .B(n7407), .S(n8231), .Z(n7411) );
  OAI211_X1 U9112 ( .C1(n7411), .C2(n7410), .A(n9200), .B(n7409), .ZN(n9212)
         );
  NAND2_X1 U9113 ( .A1(n7412), .A2(n9212), .ZN(P1_U3245) );
  XOR2_X1 U9114 ( .A(n7413), .B(n7414), .Z(n7425) );
  INV_X1 U9115 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n7417) );
  NOR2_X1 U9116 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7415), .ZN(n7877) );
  INV_X1 U9117 ( .A(n7877), .ZN(n7416) );
  OAI21_X1 U9118 ( .B1(n9281), .B2(n7417), .A(n7416), .ZN(n7422) );
  AOI211_X1 U9119 ( .C1(n7420), .C2(n7419), .A(n9251), .B(n7418), .ZN(n7421)
         );
  AOI211_X1 U9120 ( .C1(n9711), .C2(n7423), .A(n7422), .B(n7421), .ZN(n7424)
         );
  OAI21_X1 U9121 ( .B1(n9254), .B2(n7425), .A(n7424), .ZN(P1_U3251) );
  XOR2_X1 U9122 ( .A(n7426), .B(n7427), .Z(n7435) );
  INV_X1 U9123 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10126) );
  NAND2_X1 U9124 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7952) );
  OAI21_X1 U9125 ( .B1(n9281), .B2(n10126), .A(n7952), .ZN(n7432) );
  AOI211_X1 U9126 ( .C1(n7430), .C2(n7429), .A(n9251), .B(n7428), .ZN(n7431)
         );
  AOI211_X1 U9127 ( .C1(n9711), .C2(n7433), .A(n7432), .B(n7431), .ZN(n7434)
         );
  OAI21_X1 U9128 ( .B1(n9254), .B2(n7435), .A(n7434), .ZN(P1_U3250) );
  INV_X1 U9129 ( .A(n8572), .ZN(n7932) );
  OAI222_X1 U9130 ( .A1(n9040), .A2(n7437), .B1(n9038), .B2(n7436), .C1(n7932), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NAND2_X1 U9131 ( .A1(n7440), .A2(n6093), .ZN(n7438) );
  NAND2_X1 U9132 ( .A1(n7439), .A2(n7438), .ZN(n7534) );
  NAND2_X1 U9133 ( .A1(n7534), .A2(n7533), .ZN(n7532) );
  OAI21_X1 U9134 ( .B1(n7534), .B2(n7533), .A(n7532), .ZN(n7523) );
  INV_X1 U9135 ( .A(n7523), .ZN(n7447) );
  INV_X1 U9136 ( .A(n9506), .ZN(n9477) );
  OAI22_X1 U9137 ( .A1(n9477), .A2(n7440), .B1(n7543), .B2(n9474), .ZN(n7444)
         );
  XNOR2_X1 U9138 ( .A(n7533), .B(n7441), .ZN(n7442) );
  NOR2_X1 U9139 ( .A1(n7442), .A2(n7743), .ZN(n7443) );
  AOI211_X1 U9140 ( .C1(n7894), .C2(n7523), .A(n7444), .B(n7443), .ZN(n7525)
         );
  AOI21_X1 U9141 ( .B1(n7529), .B2(n7445), .A(n4929), .ZN(n7518) );
  AOI22_X1 U9142 ( .A1(n7518), .A2(n9627), .B1(n9626), .B2(n7529), .ZN(n7446)
         );
  OAI211_X1 U9143 ( .C1(n7447), .C2(n9632), .A(n7525), .B(n7446), .ZN(n7694)
         );
  NAND2_X1 U9144 ( .A1(n7694), .A2(n9801), .ZN(n7448) );
  OAI21_X1 U9145 ( .B1(n9801), .B2(n6909), .A(n7448), .ZN(P1_U3526) );
  NAND2_X1 U9146 ( .A1(n7450), .A2(n7449), .ZN(n7692) );
  INV_X1 U9147 ( .A(n7692), .ZN(n7452) );
  INV_X1 U9148 ( .A(n7451), .ZN(n9767) );
  NAND2_X1 U9149 ( .A1(n7452), .A2(n9767), .ZN(n7453) );
  INV_X1 U9150 ( .A(n7527), .ZN(n7457) );
  NOR3_X1 U9151 ( .A1(n7457), .A2(n7456), .A3(n7455), .ZN(n7458) );
  AOI21_X1 U9152 ( .B1(n9510), .B2(n6587), .A(n7458), .ZN(n7700) );
  OAI21_X1 U9153 ( .B1(n6070), .B2(n9728), .A(n7700), .ZN(n7459) );
  NAND2_X1 U9154 ( .A1(n7459), .A2(n9733), .ZN(n7464) );
  NOR2_X1 U9155 ( .A1(n7702), .A2(n7460), .ZN(n7461) );
  OAI21_X1 U9156 ( .B1(n9462), .B2(n9494), .A(n7462), .ZN(n7463) );
  OAI211_X1 U9157 ( .C1(n7465), .C2(n9733), .A(n7464), .B(n7463), .ZN(P1_U3291) );
  INV_X1 U9158 ( .A(n8462), .ZN(n8275) );
  NAND2_X1 U9159 ( .A1(n8275), .A2(n9868), .ZN(n7468) );
  XOR2_X1 U9160 ( .A(n7502), .B(n7472), .Z(n7633) );
  NAND2_X1 U9161 ( .A1(n7470), .A2(n7469), .ZN(n7471) );
  XOR2_X1 U9162 ( .A(n7472), .B(n7471), .Z(n7474) );
  OAI21_X1 U9163 ( .B1(n7474), .B2(n8831), .A(n7473), .ZN(n7629) );
  INV_X1 U9164 ( .A(n7629), .ZN(n7476) );
  MUX2_X1 U9165 ( .A(n7476), .B(n7475), .S(n8886), .Z(n7486) );
  NOR2_X1 U9166 ( .A1(n8886), .A2(n7627), .ZN(n8796) );
  INV_X1 U9167 ( .A(n8796), .ZN(n7483) );
  INV_X1 U9168 ( .A(n7479), .ZN(n7480) );
  AOI211_X1 U9169 ( .C1(n7631), .C2(n7480), .A(n9907), .B(n7508), .ZN(n7630)
         );
  INV_X1 U9170 ( .A(n7630), .ZN(n7482) );
  OAI22_X1 U9171 ( .A1(n7483), .A2(n7482), .B1(n7481), .B2(n8761), .ZN(n7484)
         );
  AOI21_X1 U9172 ( .B1(n8765), .B2(n7631), .A(n7484), .ZN(n7485) );
  OAI211_X1 U9173 ( .C1(n7633), .C2(n8854), .A(n7486), .B(n7485), .ZN(P2_U3291) );
  NOR2_X1 U9174 ( .A1(n7488), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7841) );
  AOI21_X1 U9175 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n7488), .A(n7841), .ZN(
        n7499) );
  INV_X1 U9176 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7489) );
  NAND2_X1 U9177 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8438) );
  OAI21_X1 U9178 ( .B1(n8585), .B2(n7489), .A(n8438), .ZN(n7490) );
  AOI21_X1 U9179 ( .B1(n9821), .B2(n7837), .A(n7490), .ZN(n7498) );
  NOR2_X1 U9180 ( .A1(n7491), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7492) );
  XOR2_X1 U9181 ( .A(n7837), .B(n7838), .Z(n7496) );
  INV_X1 U9182 ( .A(n7836), .ZN(n7495) );
  OAI211_X1 U9183 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n7496), .A(n7495), .B(
        n9823), .ZN(n7497) );
  OAI211_X1 U9184 ( .C1(n7499), .C2(n9827), .A(n7498), .B(n7497), .ZN(P2_U3260) );
  NAND2_X1 U9185 ( .A1(n7631), .A2(n8461), .ZN(n7501) );
  XNOR2_X1 U9186 ( .A(n7719), .B(n7504), .ZN(n9879) );
  INV_X1 U9187 ( .A(n9879), .ZN(n7513) );
  OAI21_X1 U9188 ( .B1(n7505), .B2(n7504), .A(n7503), .ZN(n7506) );
  INV_X1 U9189 ( .A(n7771), .ZN(n8459) );
  AOI222_X1 U9190 ( .A1(n8871), .A2(n7506), .B1(n8461), .B2(n8819), .C1(n8459), 
        .C2(n8817), .ZN(n9876) );
  MUX2_X1 U9191 ( .A(n7507), .B(n9876), .S(n8772), .Z(n7512) );
  INV_X1 U9192 ( .A(n7716), .ZN(n9874) );
  NAND2_X1 U9193 ( .A1(n7508), .A2(n9874), .ZN(n7781) );
  OR2_X1 U9194 ( .A1(n7508), .A2(n9874), .ZN(n7509) );
  NAND2_X1 U9195 ( .A1(n7781), .A2(n7509), .ZN(n9875) );
  OAI22_X1 U9196 ( .A1(n8687), .A2(n9875), .B1(n7568), .B2(n8761), .ZN(n7510)
         );
  AOI21_X1 U9197 ( .B1(n8765), .B2(n7716), .A(n7510), .ZN(n7511) );
  OAI211_X1 U9198 ( .C1(n7513), .C2(n8854), .A(n7512), .B(n7511), .ZN(P2_U3290) );
  INV_X1 U9199 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10036) );
  INV_X1 U9200 ( .A(n7514), .ZN(n7515) );
  INV_X1 U9201 ( .A(n9710), .ZN(n9269) );
  OAI222_X1 U9202 ( .A1(n7855), .A2(n10036), .B1(n10109), .B2(n7515), .C1(
        P1_U3084), .C2(n9269), .ZN(P1_U3335) );
  INV_X1 U9203 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7516) );
  INV_X1 U9204 ( .A(n9822), .ZN(n8573) );
  OAI222_X1 U9205 ( .A1(n9040), .A2(n7516), .B1(n9038), .B2(n7515), .C1(
        P2_U3152), .C2(n8573), .ZN(P2_U3340) );
  AND2_X1 U9206 ( .A1(n7517), .A2(n9278), .ZN(n9732) );
  NAND2_X1 U9207 ( .A1(n9733), .A2(n9732), .ZN(n9491) );
  INV_X1 U9208 ( .A(n9491), .ZN(n7942) );
  AOI22_X1 U9209 ( .A1(n9735), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9499), .B2(
        n6095), .ZN(n7520) );
  NAND2_X1 U9210 ( .A1(n9494), .A2(n7518), .ZN(n7519) );
  OAI211_X1 U9211 ( .C1(n7521), .C2(n9502), .A(n7520), .B(n7519), .ZN(n7522)
         );
  AOI21_X1 U9212 ( .B1(n7942), .B2(n7523), .A(n7522), .ZN(n7524) );
  OAI21_X1 U9213 ( .B1(n7525), .B2(n9735), .A(n7524), .ZN(P1_U3288) );
  AND2_X1 U9214 ( .A1(n7527), .A2(n7526), .ZN(n7528) );
  NOR2_X1 U9215 ( .A1(n7530), .A2(n7529), .ZN(n7536) );
  INV_X1 U9216 ( .A(n7536), .ZN(n7531) );
  NAND2_X1 U9217 ( .A1(n7532), .A2(n7531), .ZN(n7644) );
  AND2_X1 U9218 ( .A1(n7644), .A2(n7651), .ZN(n7646) );
  NOR2_X1 U9219 ( .A1(n9198), .A2(n7667), .ZN(n7535) );
  NOR2_X1 U9220 ( .A1(n7646), .A2(n7535), .ZN(n7539) );
  NAND3_X1 U9221 ( .A1(n7534), .A2(n7533), .A3(n7651), .ZN(n7538) );
  AOI21_X1 U9222 ( .B1(n7651), .B2(n7536), .A(n7535), .ZN(n7537) );
  OAI21_X1 U9223 ( .B1(n7539), .B2(n7540), .A(n7604), .ZN(n9779) );
  NOR2_X1 U9224 ( .A1(n7541), .A2(n7540), .ZN(n7735) );
  AOI21_X1 U9225 ( .B1(n7541), .B2(n7540), .A(n7735), .ZN(n7542) );
  OAI222_X1 U9226 ( .A1(n9477), .A2(n7543), .B1(n9474), .B2(n7758), .C1(n7542), 
        .C2(n7743), .ZN(n9782) );
  INV_X1 U9227 ( .A(n7745), .ZN(n7544) );
  OAI211_X1 U9228 ( .C1(n9781), .C2(n7647), .A(n7544), .B(n9627), .ZN(n9780)
         );
  INV_X1 U9229 ( .A(n7545), .ZN(n7763) );
  OAI22_X1 U9230 ( .A1(n9780), .A2(n9278), .B1(n9728), .B2(n7763), .ZN(n7546)
         );
  OAI21_X1 U9231 ( .B1(n9782), .B2(n7546), .A(n9733), .ZN(n7548) );
  AOI22_X1 U9232 ( .A1(n9462), .A2(n7602), .B1(n9735), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n7547) );
  OAI211_X1 U9233 ( .C1(n9516), .C2(n9779), .A(n7548), .B(n7547), .ZN(P1_U3286) );
  XOR2_X1 U9234 ( .A(n7550), .B(n7549), .Z(n7558) );
  INV_X1 U9235 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9990) );
  NAND2_X1 U9236 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8126) );
  OAI21_X1 U9237 ( .B1(n9281), .B2(n9990), .A(n8126), .ZN(n7555) );
  AOI211_X1 U9238 ( .C1(n7553), .C2(n7552), .A(n9251), .B(n7551), .ZN(n7554)
         );
  AOI211_X1 U9239 ( .C1(n9711), .C2(n7556), .A(n7555), .B(n7554), .ZN(n7557)
         );
  OAI21_X1 U9240 ( .B1(n9254), .B2(n7558), .A(n7557), .ZN(P1_U3253) );
  XNOR2_X1 U9241 ( .A(n7559), .B(n7560), .ZN(n7564) );
  INV_X1 U9242 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8529) );
  OAI22_X1 U9243 ( .A1(n8432), .A2(n4846), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8529), .ZN(n7562) );
  OAI22_X1 U9244 ( .A1(n8439), .A2(n7720), .B1(n8441), .B2(n7725), .ZN(n7561)
         );
  AOI211_X1 U9245 ( .C1(n7598), .C2(n8460), .A(n7562), .B(n7561), .ZN(n7563)
         );
  OAI21_X1 U9246 ( .B1(n7564), .B2(n8447), .A(n7563), .ZN(P2_U3215) );
  AOI21_X1 U9247 ( .B1(n7567), .B2(n4388), .A(n7565), .ZN(n7572) );
  OAI22_X1 U9248 ( .A1(n8432), .A2(n9874), .B1(n8441), .B2(n7771), .ZN(n7570)
         );
  NAND2_X1 U9249 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8512) );
  OAI21_X1 U9250 ( .B1(n8439), .B2(n7568), .A(n8512), .ZN(n7569) );
  AOI211_X1 U9251 ( .C1(n7598), .C2(n8461), .A(n7570), .B(n7569), .ZN(n7571)
         );
  OAI21_X1 U9252 ( .B1(n7572), .B2(n8447), .A(n7571), .ZN(P2_U3241) );
  INV_X1 U9253 ( .A(n7573), .ZN(n7574) );
  NOR2_X1 U9254 ( .A1(n7575), .A2(n7574), .ZN(n7576) );
  XNOR2_X1 U9255 ( .A(n7577), .B(n7576), .ZN(n7583) );
  OAI22_X1 U9256 ( .A1(n8432), .A2(n9868), .B1(n8441), .B2(n7578), .ZN(n7581)
         );
  NAND2_X1 U9257 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n8484) );
  OAI21_X1 U9258 ( .B1(n8439), .B2(n7579), .A(n8484), .ZN(n7580) );
  AOI211_X1 U9259 ( .C1(n7598), .C2(n8463), .A(n7581), .B(n7580), .ZN(n7582)
         );
  OAI21_X1 U9260 ( .B1(n7583), .B2(n8447), .A(n7582), .ZN(P2_U3232) );
  INV_X1 U9261 ( .A(n7584), .ZN(n7593) );
  INV_X1 U9262 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7585) );
  NOR2_X1 U9263 ( .A1(n9728), .A2(n7585), .ZN(n7588) );
  INV_X1 U9264 ( .A(n9494), .ZN(n9286) );
  NOR2_X1 U9265 ( .A1(n9286), .A2(n7586), .ZN(n7587) );
  AOI211_X1 U9266 ( .C1(n9735), .C2(P1_REG2_REG_2__SCAN_IN), .A(n7588), .B(
        n7587), .ZN(n7592) );
  AOI22_X1 U9267 ( .A1(n7942), .A2(n7590), .B1(n9462), .B2(n7589), .ZN(n7591)
         );
  OAI211_X1 U9268 ( .C1(n9735), .C2(n7593), .A(n7592), .B(n7591), .ZN(P1_U3289) );
  XNOR2_X1 U9269 ( .A(n7595), .B(n7594), .ZN(n7600) );
  OAI22_X1 U9270 ( .A1(n8432), .A2(n9886), .B1(n8441), .B2(n7984), .ZN(n7597)
         );
  NAND2_X1 U9271 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8537) );
  OAI21_X1 U9272 ( .B1(n8439), .B2(n7784), .A(n8537), .ZN(n7596) );
  AOI211_X1 U9273 ( .C1(n7598), .C2(n8459), .A(n7597), .B(n7596), .ZN(n7599)
         );
  OAI21_X1 U9274 ( .B1(n7600), .B2(n8447), .A(n7599), .ZN(P2_U3223) );
  NAND2_X1 U9275 ( .A1(n8464), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7601) );
  OAI21_X1 U9276 ( .B1(n8268), .B2(n8464), .A(n7601), .ZN(P2_U3581) );
  NAND2_X1 U9277 ( .A1(n7602), .A2(n9197), .ZN(n7603) );
  OR2_X1 U9278 ( .A1(n7605), .A2(n9196), .ZN(n7606) );
  NAND2_X1 U9279 ( .A1(n7739), .A2(n7606), .ZN(n7607) );
  OAI21_X1 U9280 ( .B1(n7607), .B2(n7801), .A(n7793), .ZN(n7608) );
  INV_X1 U9281 ( .A(n7608), .ZN(n7664) );
  NAND2_X1 U9282 ( .A1(n7610), .A2(n7609), .ZN(n7614) );
  AND2_X1 U9283 ( .A1(n7612), .A2(n7611), .ZN(n7613) );
  XNOR2_X1 U9284 ( .A(n7802), .B(n7801), .ZN(n7615) );
  AOI222_X1 U9285 ( .A1(n7615), .A2(n9509), .B1(n9196), .B2(n9506), .C1(n9194), 
        .C2(n9510), .ZN(n7663) );
  MUX2_X1 U9286 ( .A(n6887), .B(n7663), .S(n9733), .Z(n7622) );
  INV_X1 U9287 ( .A(n7797), .ZN(n7617) );
  AOI211_X1 U9288 ( .C1(n7791), .C2(n7616), .A(n9789), .B(n7617), .ZN(n7661)
         );
  NOR2_X1 U9289 ( .A1(n7618), .A2(n9278), .ZN(n9471) );
  INV_X1 U9290 ( .A(n7684), .ZN(n7619) );
  OAI22_X1 U9291 ( .A1(n9502), .A2(n4403), .B1(n9728), .B2(n7619), .ZN(n7620)
         );
  AOI21_X1 U9292 ( .B1(n7661), .B2(n9471), .A(n7620), .ZN(n7621) );
  OAI211_X1 U9293 ( .C1(n7664), .C2(n9516), .A(n7622), .B(n7621), .ZN(P1_U3284) );
  INV_X1 U9294 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7635) );
  AND2_X1 U9295 ( .A1(n7765), .A2(n7627), .ZN(n7628) );
  NAND2_X1 U9296 ( .A1(n5637), .A2(n7628), .ZN(n9860) );
  AOI211_X1 U9297 ( .C1(n8988), .C2(n7631), .A(n7630), .B(n7629), .ZN(n7632)
         );
  OAI21_X1 U9298 ( .B1(n8993), .B2(n7633), .A(n7632), .ZN(n7638) );
  NAND2_X1 U9299 ( .A1(n7638), .A2(n9913), .ZN(n7634) );
  OAI21_X1 U9300 ( .B1(n9913), .B2(n7635), .A(n7634), .ZN(P2_U3466) );
  NAND2_X1 U9301 ( .A1(n7638), .A2(n9926), .ZN(n7639) );
  OAI21_X1 U9302 ( .B1(n9926), .B2(n5092), .A(n7639), .ZN(P2_U3525) );
  INV_X1 U9303 ( .A(n7640), .ZN(n7642) );
  OAI222_X1 U9304 ( .A1(n7855), .A2(n7641), .B1(n10109), .B2(n7642), .C1(
        P1_U3084), .C2(n6576), .ZN(P1_U3334) );
  OAI222_X1 U9305 ( .A1(n9040), .A2(n7643), .B1(n9038), .B2(n7642), .C1(n8758), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  NOR2_X1 U9306 ( .A1(n7644), .A2(n7651), .ZN(n7645) );
  OR2_X1 U9307 ( .A1(n7646), .A2(n7645), .ZN(n9777) );
  AOI21_X1 U9308 ( .B1(n7667), .B2(n7648), .A(n7647), .ZN(n9773) );
  AOI22_X1 U9309 ( .A1(n9494), .A2(n9773), .B1(n7677), .B2(n9499), .ZN(n7649)
         );
  OAI21_X1 U9310 ( .B1(n4931), .B2(n9502), .A(n7649), .ZN(n7659) );
  INV_X1 U9311 ( .A(n7650), .ZN(n7653) );
  AOI21_X1 U9312 ( .B1(n6125), .B2(n7651), .A(n7743), .ZN(n7652) );
  OAI21_X1 U9313 ( .B1(n7654), .B2(n7653), .A(n7652), .ZN(n7657) );
  AOI22_X1 U9314 ( .A1(n9510), .A2(n9197), .B1(n9506), .B2(n7530), .ZN(n7656)
         );
  NAND2_X1 U9315 ( .A1(n9777), .A2(n7894), .ZN(n7655) );
  NAND3_X1 U9316 ( .A1(n7657), .A2(n7656), .A3(n7655), .ZN(n9775) );
  MUX2_X1 U9317 ( .A(n9775), .B(P1_REG2_REG_4__SCAN_IN), .S(n9735), .Z(n7658)
         );
  AOI211_X1 U9318 ( .C1(n7942), .C2(n9777), .A(n7659), .B(n7658), .ZN(n7660)
         );
  INV_X1 U9319 ( .A(n7660), .ZN(P1_U3287) );
  AOI21_X1 U9320 ( .B1(n9626), .B2(n7791), .A(n7661), .ZN(n7662) );
  OAI211_X1 U9321 ( .C1(n9624), .C2(n7664), .A(n7663), .B(n7662), .ZN(n7732)
         );
  NAND2_X1 U9322 ( .A1(n7732), .A2(n9801), .ZN(n7665) );
  OAI21_X1 U9323 ( .B1(n9801), .B2(n7666), .A(n7665), .ZN(P1_U3530) );
  AOI22_X1 U9324 ( .A1(n7667), .A2(n9184), .B1(n9180), .B2(n9197), .ZN(n7669)
         );
  OAI211_X1 U9325 ( .C1(n7670), .C2(n9178), .A(n7669), .B(n7668), .ZN(n7676)
         );
  INV_X1 U9326 ( .A(n7671), .ZN(n7672) );
  AOI211_X1 U9327 ( .C1(n7674), .C2(n7673), .A(n9186), .B(n7672), .ZN(n7675)
         );
  AOI211_X1 U9328 ( .C1(n7677), .C2(n9167), .A(n7676), .B(n7675), .ZN(n7678)
         );
  INV_X1 U9329 ( .A(n7678), .ZN(P1_U3228) );
  INV_X1 U9330 ( .A(n7679), .ZN(n7681) );
  NOR2_X1 U9331 ( .A1(n7681), .A2(n7680), .ZN(n7682) );
  XNOR2_X1 U9332 ( .A(n7683), .B(n7682), .ZN(n7691) );
  NAND2_X1 U9333 ( .A1(n9167), .A2(n7684), .ZN(n7687) );
  AOI21_X1 U9334 ( .B1(n9155), .B2(n9196), .A(n7685), .ZN(n7686) );
  OAI211_X1 U9335 ( .C1(n7688), .C2(n9152), .A(n7687), .B(n7686), .ZN(n7689)
         );
  AOI21_X1 U9336 ( .B1(n7791), .B2(n9184), .A(n7689), .ZN(n7690) );
  OAI21_X1 U9337 ( .B1(n7691), .B2(n9186), .A(n7690), .ZN(P1_U3211) );
  INV_X1 U9338 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7696) );
  NAND2_X1 U9339 ( .A1(n7694), .A2(n9655), .ZN(n7695) );
  OAI21_X1 U9340 ( .B1(n9796), .B2(n7696), .A(n7695), .ZN(P1_U3463) );
  INV_X1 U9341 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7699) );
  OR2_X1 U9342 ( .A1(n7697), .A2(n9795), .ZN(n7698) );
  OAI21_X1 U9343 ( .B1(n9796), .B2(n7699), .A(n7698), .ZN(P1_U3457) );
  INV_X1 U9344 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7704) );
  OAI21_X1 U9345 ( .B1(n7702), .B2(n7701), .A(n7700), .ZN(n9633) );
  NAND2_X1 U9346 ( .A1(n9633), .A2(n9655), .ZN(n7703) );
  OAI21_X1 U9347 ( .B1(n9796), .B2(n7704), .A(n7703), .ZN(P1_U3454) );
  XNOR2_X1 U9348 ( .A(n7706), .B(n7705), .ZN(n7715) );
  INV_X1 U9349 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U9350 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8166) );
  OAI21_X1 U9351 ( .B1(n9281), .B2(n7707), .A(n8166), .ZN(n7712) );
  AOI211_X1 U9352 ( .C1(n7710), .C2(n7709), .A(n9251), .B(n7708), .ZN(n7711)
         );
  AOI211_X1 U9353 ( .C1(n9711), .C2(n7713), .A(n7712), .B(n7711), .ZN(n7714)
         );
  OAI21_X1 U9354 ( .B1(n9254), .B2(n7715), .A(n7714), .ZN(P1_U3254) );
  AND2_X1 U9355 ( .A1(n7716), .A2(n8460), .ZN(n7718) );
  OR2_X1 U9356 ( .A1(n7716), .A2(n8460), .ZN(n7717) );
  XNOR2_X1 U9357 ( .A(n7768), .B(n7767), .ZN(n9884) );
  XNOR2_X1 U9358 ( .A(n7781), .B(n7780), .ZN(n9881) );
  INV_X1 U9359 ( .A(n7720), .ZN(n7721) );
  AOI22_X1 U9360 ( .A1(n8765), .A2(n7780), .B1(n8876), .B2(n7721), .ZN(n7722)
         );
  OAI21_X1 U9361 ( .B1(n8687), .B2(n9881), .A(n7722), .ZN(n7728) );
  XNOR2_X1 U9362 ( .A(n7723), .B(n7767), .ZN(n7724) );
  OAI222_X1 U9363 ( .A1(n8861), .A2(n7726), .B1(n8859), .B2(n7725), .C1(n7724), 
        .C2(n8831), .ZN(n9882) );
  MUX2_X1 U9364 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9882), .S(n8772), .Z(n7727)
         );
  AOI211_X1 U9365 ( .C1(n8811), .C2(n9884), .A(n7728), .B(n7727), .ZN(n7729)
         );
  INV_X1 U9366 ( .A(n7729), .ZN(P2_U3289) );
  INV_X1 U9367 ( .A(n7730), .ZN(n7764) );
  OAI222_X1 U9368 ( .A1(n7855), .A2(n7731), .B1(n10109), .B2(n7764), .C1(n6506), .C2(P1_U3084), .ZN(P1_U3333) );
  INV_X1 U9369 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10082) );
  NAND2_X1 U9370 ( .A1(n7732), .A2(n9796), .ZN(n7733) );
  OAI21_X1 U9371 ( .B1(n9796), .B2(n10082), .A(n7733), .ZN(P1_U3475) );
  NOR2_X1 U9372 ( .A1(n7735), .A2(n4508), .ZN(n7736) );
  XNOR2_X1 U9373 ( .A(n7736), .B(n4279), .ZN(n7744) );
  NAND2_X1 U9374 ( .A1(n7737), .A2(n4279), .ZN(n7738) );
  NAND2_X1 U9375 ( .A1(n7739), .A2(n7738), .ZN(n9793) );
  OAI22_X1 U9376 ( .A1(n9477), .A2(n7740), .B1(n7910), .B2(n9474), .ZN(n7741)
         );
  AOI21_X1 U9377 ( .B1(n9793), .B2(n7894), .A(n7741), .ZN(n7742) );
  OAI21_X1 U9378 ( .B1(n7744), .B2(n7743), .A(n7742), .ZN(n9791) );
  OR2_X1 U9379 ( .A1(n7745), .A2(n9788), .ZN(n7746) );
  NAND2_X1 U9380 ( .A1(n7616), .A2(n7746), .ZN(n9790) );
  NAND2_X1 U9381 ( .A1(n9793), .A2(n7942), .ZN(n7751) );
  NAND2_X1 U9382 ( .A1(n9735), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U9383 ( .A1(n9499), .A2(n7866), .ZN(n7747) );
  OAI211_X1 U9384 ( .C1(n9502), .C2(n9788), .A(n7748), .B(n7747), .ZN(n7749)
         );
  INV_X1 U9385 ( .A(n7749), .ZN(n7750) );
  OAI211_X1 U9386 ( .C1(n9286), .C2(n9790), .A(n7751), .B(n7750), .ZN(n7752)
         );
  AOI21_X1 U9387 ( .B1(n9791), .B2(n9733), .A(n7752), .ZN(n7753) );
  INV_X1 U9388 ( .A(n7753), .ZN(P1_U3285) );
  XNOR2_X1 U9389 ( .A(n7857), .B(n7754), .ZN(n7755) );
  NAND2_X1 U9390 ( .A1(n7755), .A2(n7756), .ZN(n7856) );
  OAI21_X1 U9391 ( .B1(n7756), .B2(n7755), .A(n7856), .ZN(n7757) );
  NAND2_X1 U9392 ( .A1(n7757), .A2(n9165), .ZN(n7762) );
  OAI22_X1 U9393 ( .A1(n9781), .A2(n9173), .B1(n9152), .B2(n7758), .ZN(n7759)
         );
  AOI211_X1 U9394 ( .C1(n9155), .C2(n9198), .A(n7760), .B(n7759), .ZN(n7761)
         );
  OAI211_X1 U9395 ( .C1(n9182), .C2(n7763), .A(n7762), .B(n7761), .ZN(P1_U3225) );
  OAI222_X1 U9396 ( .A1(n9040), .A2(n7766), .B1(P2_U3152), .B2(n7765), .C1(
        n9038), .C2(n7764), .ZN(P2_U3338) );
  OR2_X1 U9397 ( .A1(n7780), .A2(n8459), .ZN(n7985) );
  NAND2_X1 U9398 ( .A1(n7989), .A2(n7985), .ZN(n7769) );
  OR2_X1 U9399 ( .A1(n7769), .A2(n4912), .ZN(n8076) );
  NAND2_X1 U9400 ( .A1(n7769), .A2(n4912), .ZN(n7770) );
  NAND2_X1 U9401 ( .A1(n8076), .A2(n7770), .ZN(n7779) );
  OAI22_X1 U9402 ( .A1(n7771), .A2(n8861), .B1(n7984), .B2(n8859), .ZN(n7772)
         );
  INV_X1 U9403 ( .A(n7772), .ZN(n7777) );
  XNOR2_X1 U9404 ( .A(n7773), .B(n7774), .ZN(n7775) );
  NAND2_X1 U9405 ( .A1(n7775), .A2(n8871), .ZN(n7776) );
  OAI211_X1 U9406 ( .C1(n7779), .C2(n8867), .A(n7777), .B(n7776), .ZN(n9888)
         );
  MUX2_X1 U9407 ( .A(n9888), .B(P2_REG2_REG_8__SCAN_IN), .S(n8886), .Z(n7778)
         );
  INV_X1 U9408 ( .A(n7778), .ZN(n7790) );
  INV_X1 U9409 ( .A(n7779), .ZN(n9890) );
  INV_X1 U9410 ( .A(n8881), .ZN(n8096) );
  NAND2_X1 U9411 ( .A1(n4969), .A2(n7783), .ZN(n7782) );
  NAND2_X1 U9412 ( .A1(n8080), .A2(n7782), .ZN(n9887) );
  NAND2_X1 U9413 ( .A1(n8765), .A2(n7783), .ZN(n7787) );
  INV_X1 U9414 ( .A(n7784), .ZN(n7785) );
  NAND2_X1 U9415 ( .A1(n8876), .A2(n7785), .ZN(n7786) );
  OAI211_X1 U9416 ( .C1(n9887), .C2(n8687), .A(n7787), .B(n7786), .ZN(n7788)
         );
  AOI21_X1 U9417 ( .B1(n9890), .B2(n8096), .A(n7788), .ZN(n7789) );
  NAND2_X1 U9418 ( .A1(n7790), .A2(n7789), .ZN(P2_U3288) );
  OR2_X1 U9419 ( .A1(n7791), .A2(n9195), .ZN(n7792) );
  NAND2_X1 U9420 ( .A1(n7793), .A2(n7792), .ZN(n7795) );
  NAND2_X1 U9421 ( .A1(n7795), .A2(n7804), .ZN(n7796) );
  NAND2_X1 U9422 ( .A1(n7797), .A2(n7936), .ZN(n7798) );
  NAND2_X1 U9423 ( .A1(n7823), .A2(n7798), .ZN(n7938) );
  INV_X1 U9424 ( .A(n7936), .ZN(n7799) );
  OAI22_X1 U9425 ( .A1(n7938), .A2(n9789), .B1(n7799), .B2(n9787), .ZN(n7811)
         );
  INV_X1 U9426 ( .A(n7815), .ZN(n7806) );
  NAND2_X1 U9427 ( .A1(n4292), .A2(n7794), .ZN(n7805) );
  OAI211_X1 U9428 ( .C1(n7885), .C2(n7806), .A(n9509), .B(n7805), .ZN(n7810)
         );
  NAND2_X1 U9429 ( .A1(n9506), .A2(n9195), .ZN(n7807) );
  OAI21_X1 U9430 ( .B1(n7880), .B2(n9474), .A(n7807), .ZN(n7808) );
  AOI21_X1 U9431 ( .B1(n7943), .B2(n7894), .A(n7808), .ZN(n7809) );
  NAND2_X1 U9432 ( .A1(n7810), .A2(n7809), .ZN(n7939) );
  AOI211_X1 U9433 ( .C1(n9794), .C2(n7943), .A(n7811), .B(n7939), .ZN(n7814)
         );
  NAND2_X1 U9434 ( .A1(n9799), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7812) );
  OAI21_X1 U9435 ( .B1(n7814), .B2(n9799), .A(n7812), .ZN(P1_U3531) );
  NAND2_X1 U9436 ( .A1(n9795), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7813) );
  OAI21_X1 U9437 ( .B1(n7814), .B2(n9795), .A(n7813), .ZN(P1_U3478) );
  NAND2_X1 U9438 ( .A1(n7885), .A2(n7815), .ZN(n7816) );
  XNOR2_X1 U9439 ( .A(n7816), .B(n7819), .ZN(n7822) );
  NAND2_X1 U9440 ( .A1(n7936), .A2(n9194), .ZN(n7817) );
  XNOR2_X1 U9441 ( .A(n7896), .B(n7819), .ZN(n9631) );
  AOI22_X1 U9442 ( .A1(n9510), .A2(n9192), .B1(n9506), .B2(n9194), .ZN(n7820)
         );
  OAI21_X1 U9443 ( .B1(n9631), .B2(n9480), .A(n7820), .ZN(n7821) );
  AOI21_X1 U9444 ( .B1(n9509), .B2(n7822), .A(n7821), .ZN(n9630) );
  AOI21_X1 U9445 ( .B1(n9625), .B2(n7823), .A(n7889), .ZN(n9628) );
  INV_X1 U9446 ( .A(n9625), .ZN(n7825) );
  AOI22_X1 U9447 ( .A1(n9735), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7955), .B2(
        n9499), .ZN(n7824) );
  OAI21_X1 U9448 ( .B1(n7825), .B2(n9502), .A(n7824), .ZN(n7827) );
  NOR2_X1 U9449 ( .A1(n9631), .A2(n9491), .ZN(n7826) );
  AOI211_X1 U9450 ( .C1(n9628), .C2(n9494), .A(n7827), .B(n7826), .ZN(n7828)
         );
  OAI21_X1 U9451 ( .B1(n9735), .B2(n9630), .A(n7828), .ZN(P1_U3282) );
  XNOR2_X1 U9452 ( .A(n7830), .B(n7829), .ZN(n7835) );
  OAI22_X1 U9453 ( .A1(n8101), .A2(n8441), .B1(n8440), .B2(n7984), .ZN(n7833)
         );
  OAI21_X1 U9454 ( .B1(n8439), .B2(n7995), .A(n7831), .ZN(n7832) );
  AOI211_X1 U9455 ( .C1(n8028), .C2(n8445), .A(n7833), .B(n7832), .ZN(n7834)
         );
  OAI21_X1 U9456 ( .B1(n7835), .B2(n8447), .A(n7834), .ZN(P2_U3219) );
  XNOR2_X1 U9457 ( .A(n7921), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U9458 ( .A1(n7839), .A2(n7840), .ZN(n7922) );
  OAI21_X1 U9459 ( .B1(n7840), .B2(n7839), .A(n7922), .ZN(n7851) );
  INV_X1 U9460 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7843) );
  MUX2_X1 U9461 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n7843), .S(n7921), .Z(n7844)
         );
  INV_X1 U9462 ( .A(n7844), .ZN(n7845) );
  OAI211_X1 U9463 ( .C1(n7846), .C2(n7845), .A(n8579), .B(n7926), .ZN(n7849)
         );
  NOR2_X1 U9464 ( .A1(n7847), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8368) );
  AOI21_X1 U9465 ( .B1(n9817), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8368), .ZN(
        n7848) );
  OAI211_X1 U9466 ( .C1(n9805), .C2(n7921), .A(n7849), .B(n7848), .ZN(n7850)
         );
  AOI21_X1 U9467 ( .B1(n9823), .B2(n7851), .A(n7850), .ZN(n7852) );
  INV_X1 U9468 ( .A(n7852), .ZN(P2_U3261) );
  INV_X1 U9469 ( .A(n7853), .ZN(n7869) );
  OAI222_X1 U9470 ( .A1(n7855), .A2(n10033), .B1(n10109), .B2(n7869), .C1(
        n7854), .C2(P1_U3084), .ZN(P1_U3332) );
  OAI21_X1 U9471 ( .B1(n7858), .B2(n7857), .A(n7856), .ZN(n7862) );
  XNOR2_X1 U9472 ( .A(n7860), .B(n7859), .ZN(n7861) );
  XNOR2_X1 U9473 ( .A(n7862), .B(n7861), .ZN(n7868) );
  NAND2_X1 U9474 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9224) );
  OAI21_X1 U9475 ( .B1(n9152), .B2(n7910), .A(n9224), .ZN(n7863) );
  AOI21_X1 U9476 ( .B1(n9155), .B2(n9197), .A(n7863), .ZN(n7864) );
  OAI21_X1 U9477 ( .B1(n9788), .B2(n9173), .A(n7864), .ZN(n7865) );
  AOI21_X1 U9478 ( .B1(n7866), .B2(n9167), .A(n7865), .ZN(n7867) );
  OAI21_X1 U9479 ( .B1(n7868), .B2(n9186), .A(n7867), .ZN(P1_U3237) );
  OAI222_X1 U9480 ( .A1(n9040), .A2(n7871), .B1(P2_U3152), .B2(n7870), .C1(
        n9038), .C2(n7869), .ZN(P2_U3337) );
  XNOR2_X1 U9481 ( .A(n7875), .B(n7874), .ZN(n7876) );
  XNOR2_X1 U9482 ( .A(n7873), .B(n7876), .ZN(n7883) );
  NAND2_X1 U9483 ( .A1(n9167), .A2(n7891), .ZN(n7879) );
  AOI21_X1 U9484 ( .B1(n9180), .B2(n9191), .A(n7877), .ZN(n7878) );
  OAI211_X1 U9485 ( .C1(n7880), .C2(n9178), .A(n7879), .B(n7878), .ZN(n7881)
         );
  AOI21_X1 U9486 ( .B1(n9620), .B2(n9184), .A(n7881), .ZN(n7882) );
  OAI21_X1 U9487 ( .B1(n7883), .B2(n9186), .A(n7882), .ZN(P1_U3215) );
  NAND2_X1 U9488 ( .A1(n7885), .A2(n7884), .ZN(n7965) );
  NAND2_X1 U9489 ( .A1(n7965), .A2(n7886), .ZN(n7887) );
  XOR2_X1 U9490 ( .A(n7959), .B(n7887), .Z(n7888) );
  AOI222_X1 U9491 ( .A1(n9191), .A2(n9510), .B1(n9509), .B2(n7888), .C1(n9193), 
        .C2(n9506), .ZN(n9622) );
  INV_X1 U9492 ( .A(n7889), .ZN(n7890) );
  AOI211_X1 U9493 ( .C1(n9620), .C2(n7890), .A(n9789), .B(n7973), .ZN(n9619)
         );
  AOI22_X1 U9494 ( .A1(n9735), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7891), .B2(
        n9499), .ZN(n7892) );
  OAI21_X1 U9495 ( .B1(n7893), .B2(n9502), .A(n7892), .ZN(n7899) );
  NAND2_X1 U9496 ( .A1(n9733), .A2(n7894), .ZN(n7897) );
  AND2_X1 U9497 ( .A1(n9625), .A2(n9193), .ZN(n7895) );
  XOR2_X1 U9498 ( .A(n7960), .B(n7959), .Z(n9623) );
  AOI21_X1 U9499 ( .B1(n9491), .B2(n7897), .A(n9623), .ZN(n7898) );
  AOI211_X1 U9500 ( .C1(n9619), .C2(n9471), .A(n7899), .B(n7898), .ZN(n7900)
         );
  OAI21_X1 U9501 ( .B1(n9622), .B2(n9735), .A(n7900), .ZN(P1_U3281) );
  NOR2_X1 U9502 ( .A1(n7903), .A2(n7902), .ZN(n7947) );
  INV_X1 U9503 ( .A(n7947), .ZN(n7904) );
  NAND2_X1 U9504 ( .A1(n7903), .A2(n7902), .ZN(n7945) );
  NAND2_X1 U9505 ( .A1(n7904), .A2(n7945), .ZN(n7906) );
  XNOR2_X1 U9506 ( .A(n7906), .B(n7905), .ZN(n7913) );
  NAND2_X1 U9507 ( .A1(n9167), .A2(n7935), .ZN(n7909) );
  AOI21_X1 U9508 ( .B1(n9180), .B2(n9193), .A(n7907), .ZN(n7908) );
  OAI211_X1 U9509 ( .C1(n7910), .C2(n9178), .A(n7909), .B(n7908), .ZN(n7911)
         );
  AOI21_X1 U9510 ( .B1(n7936), .B2(n9184), .A(n7911), .ZN(n7912) );
  OAI21_X1 U9511 ( .B1(n7913), .B2(n9186), .A(n7912), .ZN(P1_U3219) );
  XNOR2_X1 U9512 ( .A(n7914), .B(n7915), .ZN(n7920) );
  OAI22_X1 U9513 ( .A1(n8862), .A2(n8441), .B1(n8440), .B2(n8021), .ZN(n7918)
         );
  OAI22_X1 U9514 ( .A1(n8439), .A2(n8025), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7916), .ZN(n7917) );
  AOI211_X1 U9515 ( .C1(n8987), .C2(n8445), .A(n7918), .B(n7917), .ZN(n7919)
         );
  OAI21_X1 U9516 ( .B1(n7920), .B2(n8447), .A(n7919), .ZN(P2_U3238) );
  XNOR2_X1 U9517 ( .A(n8572), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7924) );
  INV_X1 U9518 ( .A(n7921), .ZN(n7925) );
  OAI21_X1 U9519 ( .B1(n7925), .B2(P2_REG1_REG_16__SCAN_IN), .A(n7922), .ZN(
        n7923) );
  NOR2_X1 U9520 ( .A1(n7923), .A2(n7924), .ZN(n8571) );
  AOI211_X1 U9521 ( .C1(n7924), .C2(n7923), .A(n9807), .B(n8571), .ZN(n7934)
         );
  AOI22_X1 U9522 ( .A1(n8572), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n5349), .B2(
        n7932), .ZN(n7929) );
  NAND2_X1 U9523 ( .A1(n7925), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7927) );
  NAND2_X1 U9524 ( .A1(n7927), .A2(n7926), .ZN(n7928) );
  OAI211_X1 U9525 ( .C1(n7929), .C2(n7928), .A(n8579), .B(n8567), .ZN(n7931)
         );
  NOR2_X1 U9526 ( .A1(n9956), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8375) );
  AOI21_X1 U9527 ( .B1(n9817), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8375), .ZN(
        n7930) );
  OAI211_X1 U9528 ( .C1(n9805), .C2(n7932), .A(n7931), .B(n7930), .ZN(n7933)
         );
  OR2_X1 U9529 ( .A1(n7934), .A2(n7933), .ZN(P2_U3262) );
  AOI22_X1 U9530 ( .A1(n9462), .A2(n7936), .B1(n9499), .B2(n7935), .ZN(n7937)
         );
  OAI21_X1 U9531 ( .B1(n7938), .B2(n9286), .A(n7937), .ZN(n7941) );
  MUX2_X1 U9532 ( .A(n7939), .B(P1_REG2_REG_8__SCAN_IN), .S(n9735), .Z(n7940)
         );
  AOI211_X1 U9533 ( .C1(n7943), .C2(n7942), .A(n7941), .B(n7940), .ZN(n7944)
         );
  INV_X1 U9534 ( .A(n7944), .ZN(P1_U3283) );
  OAI21_X1 U9535 ( .B1(n7947), .B2(n7946), .A(n7945), .ZN(n7951) );
  XNOR2_X1 U9536 ( .A(n7949), .B(n7948), .ZN(n7950) );
  XNOR2_X1 U9537 ( .A(n7951), .B(n7950), .ZN(n7958) );
  NAND2_X1 U9538 ( .A1(n9155), .A2(n9194), .ZN(n7953) );
  OAI211_X1 U9539 ( .C1(n7969), .C2(n9152), .A(n7953), .B(n7952), .ZN(n7954)
         );
  AOI21_X1 U9540 ( .B1(n7955), .B2(n9167), .A(n7954), .ZN(n7957) );
  NAND2_X1 U9541 ( .A1(n9184), .A2(n9625), .ZN(n7956) );
  OAI211_X1 U9542 ( .C1(n7958), .C2(n9186), .A(n7957), .B(n7956), .ZN(P1_U3229) );
  OR2_X1 U9543 ( .A1(n9620), .A2(n9192), .ZN(n7961) );
  NAND2_X1 U9544 ( .A1(n7962), .A2(n7961), .ZN(n8045) );
  XNOR2_X1 U9545 ( .A(n8045), .B(n7963), .ZN(n8056) );
  NAND2_X1 U9546 ( .A1(n7965), .A2(n7964), .ZN(n7967) );
  XNOR2_X1 U9547 ( .A(n8038), .B(n7968), .ZN(n7971) );
  OAI22_X1 U9548 ( .A1(n9477), .A2(n7969), .B1(n8136), .B2(n9474), .ZN(n7970)
         );
  AOI21_X1 U9549 ( .B1(n7971), .B2(n9509), .A(n7970), .ZN(n7972) );
  OAI21_X1 U9550 ( .B1(n8056), .B2(n9480), .A(n7972), .ZN(n8059) );
  NAND2_X1 U9551 ( .A1(n8059), .A2(n9733), .ZN(n7979) );
  NOR2_X1 U9552 ( .A1(n7973), .A2(n8057), .ZN(n7974) );
  OR2_X1 U9553 ( .A1(n8049), .A2(n7974), .ZN(n8058) );
  INV_X1 U9554 ( .A(n8058), .ZN(n7977) );
  AOI22_X1 U9555 ( .A1(n9735), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8014), .B2(
        n9499), .ZN(n7975) );
  OAI21_X1 U9556 ( .B1(n8057), .B2(n9502), .A(n7975), .ZN(n7976) );
  AOI21_X1 U9557 ( .B1(n7977), .B2(n9494), .A(n7976), .ZN(n7978) );
  OAI211_X1 U9558 ( .C1(n8056), .C2(n9491), .A(n7979), .B(n7978), .ZN(P1_U3280) );
  INV_X1 U9559 ( .A(n7980), .ZN(n8172) );
  AOI22_X1 U9560 ( .A1(n6530), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n10113), .ZN(n7981) );
  OAI21_X1 U9561 ( .B1(n8172), .B2(n10109), .A(n7981), .ZN(P1_U3331) );
  XNOR2_X1 U9562 ( .A(n7982), .B(n7993), .ZN(n7983) );
  OAI222_X1 U9563 ( .A1(n8861), .A2(n7984), .B1(n8859), .B2(n8101), .C1(n7983), 
        .C2(n8831), .ZN(n9911) );
  MUX2_X1 U9564 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n9911), .S(n8772), .Z(n8000)
         );
  INV_X1 U9565 ( .A(n8028), .ZN(n9906) );
  OAI21_X1 U9566 ( .B1(n8079), .B2(n9906), .A(n8024), .ZN(n9908) );
  INV_X1 U9567 ( .A(n7984), .ZN(n8457) );
  OR2_X1 U9568 ( .A1(n8085), .A2(n8457), .ZN(n7991) );
  INV_X1 U9569 ( .A(n8072), .ZN(n7990) );
  NAND2_X1 U9570 ( .A1(n8074), .A2(n7991), .ZN(n7992) );
  OR2_X1 U9571 ( .A1(n7994), .A2(n7993), .ZN(n9903) );
  NAND3_X1 U9572 ( .A1(n9903), .A2(n8811), .A3(n9904), .ZN(n7998) );
  NOR2_X1 U9573 ( .A1(n8761), .A2(n7995), .ZN(n7996) );
  AOI21_X1 U9574 ( .B1(n8765), .B2(n8028), .A(n7996), .ZN(n7997) );
  OAI211_X1 U9575 ( .C1(n8687), .C2(n9908), .A(n7998), .B(n7997), .ZN(n7999)
         );
  OR2_X1 U9576 ( .A1(n8000), .A2(n7999), .ZN(P2_U3286) );
  XNOR2_X1 U9577 ( .A(n8001), .B(n8002), .ZN(n8007) );
  OAI22_X1 U9578 ( .A1(n8834), .A2(n8441), .B1(n8440), .B2(n8101), .ZN(n8005)
         );
  OAI21_X1 U9579 ( .B1(n8439), .B2(n8114), .A(n8003), .ZN(n8004) );
  AOI211_X1 U9580 ( .C1(n8982), .C2(n8445), .A(n8005), .B(n8004), .ZN(n8006)
         );
  OAI21_X1 U9581 ( .B1(n8007), .B2(n8447), .A(n8006), .ZN(P2_U3226) );
  XNOR2_X1 U9582 ( .A(n8009), .B(n8008), .ZN(n8016) );
  NAND2_X1 U9583 ( .A1(n9155), .A2(n9192), .ZN(n8011) );
  OAI211_X1 U9584 ( .C1(n8136), .C2(n9152), .A(n8011), .B(n8010), .ZN(n8013)
         );
  NOR2_X1 U9585 ( .A1(n8057), .A2(n9173), .ZN(n8012) );
  AOI211_X1 U9586 ( .C1(n8014), .C2(n9167), .A(n8013), .B(n8012), .ZN(n8015)
         );
  OAI21_X1 U9587 ( .B1(n8016), .B2(n9186), .A(n8015), .ZN(P1_U3234) );
  INV_X1 U9588 ( .A(n8017), .ZN(n10110) );
  AOI21_X1 U9589 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9026), .A(n8018), .ZN(
        n8019) );
  OAI21_X1 U9590 ( .B1(n10110), .B2(n9038), .A(n8019), .ZN(P2_U3335) );
  XNOR2_X1 U9591 ( .A(n8020), .B(n8030), .ZN(n8022) );
  INV_X1 U9592 ( .A(n8021), .ZN(n8456) );
  AOI222_X1 U9593 ( .A1(n8871), .A2(n8022), .B1(n8456), .B2(n8819), .C1(n8454), 
        .C2(n8817), .ZN(n8991) );
  INV_X1 U9594 ( .A(n8113), .ZN(n8023) );
  AOI21_X1 U9595 ( .B1(n8987), .B2(n8024), .A(n8023), .ZN(n8989) );
  INV_X1 U9596 ( .A(n8025), .ZN(n8026) );
  AOI22_X1 U9597 ( .A1(n8886), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8026), .B2(
        n8876), .ZN(n8027) );
  OAI21_X1 U9598 ( .B1(n8879), .B2(n4421), .A(n8027), .ZN(n8035) );
  NAND2_X1 U9599 ( .A1(n8028), .A2(n8456), .ZN(n8029) );
  INV_X1 U9600 ( .A(n8030), .ZN(n8031) );
  OR2_X1 U9601 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  NAND2_X1 U9602 ( .A1(n8103), .A2(n8033), .ZN(n8992) );
  NOR2_X1 U9603 ( .A1(n8992), .A2(n8854), .ZN(n8034) );
  AOI211_X1 U9604 ( .C1(n8989), .C2(n8884), .A(n8035), .B(n8034), .ZN(n8036)
         );
  OAI21_X1 U9605 ( .B1(n8991), .B2(n8886), .A(n8036), .ZN(P2_U3285) );
  NAND2_X1 U9606 ( .A1(n8142), .A2(n8039), .ZN(n8040) );
  XNOR2_X1 U9607 ( .A(n8040), .B(n8134), .ZN(n8048) );
  OAI22_X1 U9608 ( .A1(n9477), .A2(n8041), .B1(n9049), .B2(n9474), .ZN(n8047)
         );
  NOR2_X1 U9609 ( .A1(n8042), .A2(n9191), .ZN(n8044) );
  NAND2_X1 U9610 ( .A1(n8042), .A2(n9191), .ZN(n8043) );
  XNOR2_X1 U9611 ( .A(n8135), .B(n8134), .ZN(n9618) );
  NOR2_X1 U9612 ( .A1(n9618), .A2(n9480), .ZN(n8046) );
  AOI211_X1 U9613 ( .C1(n9509), .C2(n8048), .A(n8047), .B(n8046), .ZN(n9617)
         );
  INV_X1 U9614 ( .A(n8049), .ZN(n8051) );
  INV_X1 U9615 ( .A(n8150), .ZN(n8050) );
  AOI211_X1 U9616 ( .C1(n9615), .C2(n8051), .A(n9789), .B(n8050), .ZN(n9614)
         );
  AOI22_X1 U9617 ( .A1(n9735), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n8131), .B2(
        n9499), .ZN(n8052) );
  OAI21_X1 U9618 ( .B1(n8128), .B2(n9502), .A(n8052), .ZN(n8054) );
  NOR2_X1 U9619 ( .A1(n9618), .A2(n9491), .ZN(n8053) );
  AOI211_X1 U9620 ( .C1(n9614), .C2(n9471), .A(n8054), .B(n8053), .ZN(n8055)
         );
  OAI21_X1 U9621 ( .B1(n9617), .B2(n9735), .A(n8055), .ZN(P1_U3279) );
  INV_X1 U9622 ( .A(n8056), .ZN(n8061) );
  OAI22_X1 U9623 ( .A1(n8058), .A2(n9789), .B1(n8057), .B2(n9787), .ZN(n8060)
         );
  AOI211_X1 U9624 ( .C1(n9794), .C2(n8061), .A(n8060), .B(n8059), .ZN(n8064)
         );
  NAND2_X1 U9625 ( .A1(n9799), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8062) );
  OAI21_X1 U9626 ( .B1(n8064), .B2(n9799), .A(n8062), .ZN(P1_U3534) );
  NAND2_X1 U9627 ( .A1(n9795), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8063) );
  OAI21_X1 U9628 ( .B1(n8064), .B2(n9795), .A(n8063), .ZN(P1_U3487) );
  XNOR2_X1 U9629 ( .A(n8065), .B(n8066), .ZN(n8071) );
  OAI22_X1 U9630 ( .A1(n8862), .A2(n8440), .B1(n8441), .B2(n8860), .ZN(n8069)
         );
  OAI21_X1 U9631 ( .B1(n8439), .B2(n8875), .A(n8067), .ZN(n8068) );
  AOI211_X1 U9632 ( .C1(n8977), .C2(n8445), .A(n8069), .B(n8068), .ZN(n8070)
         );
  OAI21_X1 U9633 ( .B1(n8071), .B2(n8447), .A(n8070), .ZN(P2_U3236) );
  NAND2_X1 U9634 ( .A1(n8076), .A2(n8072), .ZN(n8073) );
  NAND2_X1 U9635 ( .A1(n8073), .A2(n8088), .ZN(n8078) );
  INV_X1 U9636 ( .A(n8074), .ZN(n8075) );
  NAND2_X1 U9637 ( .A1(n8076), .A2(n8075), .ZN(n8077) );
  NAND2_X1 U9638 ( .A1(n8078), .A2(n8077), .ZN(n9893) );
  INV_X1 U9639 ( .A(n8079), .ZN(n8082) );
  NAND2_X1 U9640 ( .A1(n8080), .A2(n8085), .ZN(n8081) );
  NAND2_X1 U9641 ( .A1(n8082), .A2(n8081), .ZN(n9895) );
  INV_X1 U9642 ( .A(n8083), .ZN(n8084) );
  AOI22_X1 U9643 ( .A1(n8765), .A2(n8085), .B1(n8876), .B2(n8084), .ZN(n8086)
         );
  OAI21_X1 U9644 ( .B1(n9895), .B2(n8687), .A(n8086), .ZN(n8095) );
  NAND2_X1 U9645 ( .A1(n9893), .A2(n8087), .ZN(n8093) );
  XNOR2_X1 U9646 ( .A(n8089), .B(n8088), .ZN(n8090) );
  NAND2_X1 U9647 ( .A1(n8090), .A2(n8871), .ZN(n8092) );
  AOI22_X1 U9648 ( .A1(n8456), .A2(n8817), .B1(n8819), .B2(n8458), .ZN(n8091)
         );
  NAND3_X1 U9649 ( .A1(n8093), .A2(n8092), .A3(n8091), .ZN(n9900) );
  MUX2_X1 U9650 ( .A(n9900), .B(P2_REG2_REG_9__SCAN_IN), .S(n8886), .Z(n8094)
         );
  AOI211_X1 U9651 ( .C1(n8096), .C2(n9893), .A(n8095), .B(n8094), .ZN(n8097)
         );
  INV_X1 U9652 ( .A(n8097), .ZN(P2_U3287) );
  INV_X1 U9653 ( .A(n8098), .ZN(n8120) );
  AOI22_X1 U9654 ( .A1(n8099), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10113), .ZN(n8100) );
  OAI21_X1 U9655 ( .B1(n8120), .B2(n10109), .A(n8100), .ZN(P1_U3329) );
  INV_X1 U9656 ( .A(n8109), .ZN(n8106) );
  INV_X1 U9657 ( .A(n8101), .ZN(n8455) );
  NAND2_X1 U9658 ( .A1(n8987), .A2(n8455), .ZN(n8102) );
  INV_X1 U9659 ( .A(n8849), .ZN(n8104) );
  AOI21_X1 U9660 ( .B1(n8106), .B2(n8105), .A(n8104), .ZN(n8986) );
  NAND2_X1 U9661 ( .A1(n8108), .A2(n8107), .ZN(n8110) );
  XNOR2_X1 U9662 ( .A(n8110), .B(n8109), .ZN(n8111) );
  AOI222_X1 U9663 ( .A1(n8871), .A2(n8111), .B1(n8455), .B2(n8819), .C1(n8453), 
        .C2(n8817), .ZN(n8985) );
  MUX2_X1 U9664 ( .A(n8112), .B(n8985), .S(n8772), .Z(n8118) );
  AOI21_X1 U9665 ( .B1(n8982), .B2(n8113), .A(n8872), .ZN(n8983) );
  INV_X1 U9666 ( .A(n8982), .ZN(n8115) );
  OAI22_X1 U9667 ( .A1(n8115), .A2(n8879), .B1(n8761), .B2(n8114), .ZN(n8116)
         );
  AOI21_X1 U9668 ( .B1(n8983), .B2(n8884), .A(n8116), .ZN(n8117) );
  OAI211_X1 U9669 ( .C1(n8986), .C2(n8854), .A(n8118), .B(n8117), .ZN(P2_U3284) );
  OAI222_X1 U9670 ( .A1(n8121), .A2(P2_U3152), .B1(n9038), .B2(n8120), .C1(
        n8119), .C2(n9040), .ZN(P2_U3334) );
  INV_X1 U9671 ( .A(n8122), .ZN(n8123) );
  AOI21_X1 U9672 ( .B1(n8125), .B2(n8124), .A(n8123), .ZN(n8133) );
  NAND2_X1 U9673 ( .A1(n9155), .A2(n9191), .ZN(n8127) );
  OAI211_X1 U9674 ( .C1(n9049), .C2(n9152), .A(n8127), .B(n8126), .ZN(n8130)
         );
  NOR2_X1 U9675 ( .A1(n8128), .A2(n9173), .ZN(n8129) );
  AOI211_X1 U9676 ( .C1(n8131), .C2(n9167), .A(n8130), .B(n8129), .ZN(n8132)
         );
  OAI21_X1 U9677 ( .B1(n8133), .B2(n9186), .A(n8132), .ZN(P1_U3222) );
  INV_X1 U9678 ( .A(n8136), .ZN(n9507) );
  NAND2_X1 U9679 ( .A1(n9615), .A2(n9507), .ZN(n8137) );
  AND2_X1 U9680 ( .A1(n9610), .A2(n9190), .ZN(n8140) );
  OR2_X1 U9681 ( .A1(n9610), .A2(n9190), .ZN(n8139) );
  XNOR2_X1 U9682 ( .A(n8175), .B(n8146), .ZN(n9608) );
  INV_X1 U9683 ( .A(n9052), .ZN(n8149) );
  OAI211_X1 U9684 ( .C1(n4949), .C2(n8146), .A(n9509), .B(n8204), .ZN(n8148)
         );
  AOI22_X1 U9685 ( .A1(n9510), .A2(n9458), .B1(n9506), .B2(n9190), .ZN(n8147)
         );
  NAND2_X1 U9686 ( .A1(n8148), .A2(n8147), .ZN(n9604) );
  AOI21_X1 U9687 ( .B1(n8149), .B2(n9499), .A(n9604), .ZN(n8155) );
  AOI22_X1 U9688 ( .A1(n9606), .A2(n9462), .B1(n9735), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n8154) );
  NAND2_X1 U9689 ( .A1(n9497), .A2(n9606), .ZN(n8151) );
  NAND2_X1 U9690 ( .A1(n8151), .A2(n9627), .ZN(n8152) );
  NOR2_X1 U9691 ( .A1(n9484), .A2(n8152), .ZN(n9605) );
  NAND2_X1 U9692 ( .A1(n9605), .A2(n9471), .ZN(n8153) );
  OAI211_X1 U9693 ( .C1(n8155), .C2(n9735), .A(n8154), .B(n8153), .ZN(n8156)
         );
  INV_X1 U9694 ( .A(n8156), .ZN(n8157) );
  OAI21_X1 U9695 ( .B1(n9608), .B2(n9516), .A(n8157), .ZN(P1_U3277) );
  INV_X1 U9696 ( .A(n8158), .ZN(n9037) );
  AOI22_X1 U9697 ( .A1(n8159), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n10113), .ZN(n8160) );
  OAI21_X1 U9698 ( .B1(n9037), .B2(n10109), .A(n8160), .ZN(P1_U3328) );
  INV_X1 U9699 ( .A(n8161), .ZN(n8163) );
  NAND2_X1 U9700 ( .A1(n8163), .A2(n8162), .ZN(n8164) );
  XNOR2_X1 U9701 ( .A(n8165), .B(n8164), .ZN(n8171) );
  NAND2_X1 U9702 ( .A1(n9155), .A2(n9507), .ZN(n8167) );
  OAI211_X1 U9703 ( .C1(n9476), .C2(n9152), .A(n8167), .B(n8166), .ZN(n8168)
         );
  AOI21_X1 U9704 ( .B1(n9500), .B2(n9167), .A(n8168), .ZN(n8170) );
  NAND2_X1 U9705 ( .A1(n9610), .A2(n9184), .ZN(n8169) );
  OAI211_X1 U9706 ( .C1(n8171), .C2(n9186), .A(n8170), .B(n8169), .ZN(P1_U3232) );
  OAI222_X1 U9707 ( .A1(n9040), .A2(n8173), .B1(n9038), .B2(n8172), .C1(n5637), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9708 ( .A(n9606), .ZN(n8174) );
  AND2_X1 U9709 ( .A1(n9599), .A2(n9458), .ZN(n8176) );
  NAND2_X1 U9710 ( .A1(n9595), .A2(n9448), .ZN(n8178) );
  OR2_X1 U9711 ( .A1(n9589), .A2(n9457), .ZN(n8179) );
  NAND2_X1 U9712 ( .A1(n9589), .A2(n9457), .ZN(n8180) );
  NAND2_X1 U9713 ( .A1(n9424), .A2(n9434), .ZN(n8182) );
  NAND2_X1 U9714 ( .A1(n9584), .A2(n9450), .ZN(n8181) );
  OR2_X1 U9715 ( .A1(n9580), .A2(n9436), .ZN(n8183) );
  NAND2_X1 U9716 ( .A1(n9580), .A2(n9436), .ZN(n8184) );
  AND2_X1 U9717 ( .A1(n9574), .A2(n9420), .ZN(n8187) );
  OR2_X1 U9718 ( .A1(n9574), .A2(n9420), .ZN(n8186) );
  OR2_X1 U9719 ( .A1(n9564), .A2(n9392), .ZN(n8188) );
  NAND2_X1 U9720 ( .A1(n9564), .A2(n9392), .ZN(n8189) );
  OR2_X1 U9721 ( .A1(n9559), .A2(n9377), .ZN(n8191) );
  NAND2_X1 U9722 ( .A1(n9559), .A2(n9377), .ZN(n8192) );
  AND2_X1 U9723 ( .A1(n4942), .A2(n9362), .ZN(n8193) );
  NOR2_X1 U9724 ( .A1(n9550), .A2(n9348), .ZN(n8194) );
  NAND2_X1 U9725 ( .A1(n9536), .A2(n9297), .ZN(n9530) );
  NAND2_X1 U9726 ( .A1(n9534), .A2(n9530), .ZN(n8198) );
  XNOR2_X1 U9727 ( .A(n8198), .B(n9531), .ZN(n8238) );
  NAND2_X1 U9728 ( .A1(n9413), .A2(n9404), .ZN(n9398) );
  NOR2_X2 U9729 ( .A1(n9398), .A2(n9570), .ZN(n9383) );
  NAND2_X2 U9730 ( .A1(n9383), .A2(n9373), .ZN(n9367) );
  NOR2_X4 U9731 ( .A1(n9367), .A2(n9559), .ZN(n9353) );
  AOI211_X1 U9732 ( .C1(n9527), .C2(n8296), .A(n9789), .B(n9287), .ZN(n9525)
         );
  NOR2_X1 U9733 ( .A1(n9735), .A2(n9278), .ZN(n9514) );
  INV_X1 U9734 ( .A(n9527), .ZN(n8202) );
  INV_X1 U9735 ( .A(n8199), .ZN(n8200) );
  AOI22_X1 U9736 ( .A1(n8200), .A2(n9499), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9735), .ZN(n8201) );
  OAI21_X1 U9737 ( .B1(n8202), .B2(n9502), .A(n8201), .ZN(n8236) );
  NOR2_X1 U9738 ( .A1(n4907), .A2(n8215), .ZN(n8216) );
  INV_X1 U9739 ( .A(n9358), .ZN(n8218) );
  NAND2_X1 U9740 ( .A1(n9294), .A2(n9296), .ZN(n9295) );
  NAND2_X1 U9741 ( .A1(n9295), .A2(n8225), .ZN(n8304) );
  INV_X1 U9742 ( .A(n8226), .ZN(n8228) );
  XNOR2_X1 U9743 ( .A(n8229), .B(n9532), .ZN(n8235) );
  NOR2_X1 U9744 ( .A1(n8231), .A2(n8230), .ZN(n8232) );
  NOR2_X1 U9745 ( .A1(n9474), .A2(n8232), .ZN(n9283) );
  AOI22_X1 U9746 ( .A1(n9297), .A2(n9506), .B1(n9283), .B2(n9188), .ZN(n8233)
         );
  AOI21_X2 U9747 ( .B1(n8235), .B2(n9509), .A(n8234), .ZN(n9529) );
  OAI21_X1 U9748 ( .B1(n8238), .B2(n9516), .A(n8237), .ZN(P1_U3355) );
  INV_X1 U9749 ( .A(n8977), .ZN(n8880) );
  NOR2_X1 U9750 ( .A1(n8982), .A2(n8454), .ZN(n8844) );
  AOI21_X1 U9751 ( .B1(n8880), .B2(n8834), .A(n8844), .ZN(n8848) );
  INV_X1 U9752 ( .A(n8860), .ZN(n8820) );
  OR2_X1 U9753 ( .A1(n5859), .A2(n8820), .ZN(n8240) );
  AND2_X1 U9754 ( .A1(n8848), .A2(n8240), .ZN(n8243) );
  AND2_X1 U9755 ( .A1(n8977), .A2(n8453), .ZN(n8846) );
  NOR2_X1 U9756 ( .A1(n8239), .A2(n8846), .ZN(n8850) );
  INV_X1 U9757 ( .A(n8240), .ZN(n8241) );
  NOR2_X1 U9758 ( .A1(n8850), .A2(n8241), .ZN(n8242) );
  INV_X1 U9759 ( .A(n8835), .ZN(n8799) );
  OR2_X1 U9760 ( .A1(n8968), .A2(n8799), .ZN(n8807) );
  OR2_X1 U9761 ( .A1(n8804), .A2(n8442), .ZN(n8245) );
  INV_X1 U9762 ( .A(n8415), .ZN(n8800) );
  OR2_X1 U9763 ( .A1(n8958), .A2(n8800), .ZN(n8247) );
  NAND2_X1 U9764 ( .A1(n8791), .A2(n8247), .ZN(n8768) );
  INV_X1 U9765 ( .A(n8372), .ZN(n8452) );
  NOR2_X1 U9766 ( .A1(n8952), .A2(n8452), .ZN(n8248) );
  INV_X1 U9767 ( .A(n8952), .ZN(n8773) );
  AND2_X1 U9768 ( .A1(n8948), .A2(n8776), .ZN(n8249) );
  OR2_X1 U9769 ( .A1(n8948), .A2(n8776), .ZN(n8250) );
  INV_X1 U9770 ( .A(n8250), .ZN(n8251) );
  INV_X1 U9771 ( .A(n8339), .ZN(n8728) );
  NAND2_X1 U9772 ( .A1(n8942), .A2(n8728), .ZN(n8252) );
  INV_X1 U9773 ( .A(n8736), .ZN(n8714) );
  OR2_X1 U9774 ( .A1(n8936), .A2(n8714), .ZN(n8253) );
  NAND2_X1 U9775 ( .A1(n8936), .A2(n8714), .ZN(n8254) );
  INV_X1 U9776 ( .A(n8926), .ZN(n8695) );
  INV_X1 U9777 ( .A(n8655), .ZN(n8668) );
  INV_X1 U9778 ( .A(n8631), .ZN(n8450) );
  INV_X1 U9779 ( .A(n8931), .ZN(n8709) );
  INV_X1 U9780 ( .A(n8948), .ZN(n8259) );
  INV_X1 U9781 ( .A(n8916), .ZN(n8666) );
  AOI21_X1 U9782 ( .B1(n8900), .B2(n8620), .A(n8605), .ZN(n8901) );
  AOI22_X1 U9783 ( .A1(n8261), .A2(n8876), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8886), .ZN(n8262) );
  OAI21_X1 U9784 ( .B1(n8263), .B2(n8879), .A(n8262), .ZN(n8272) );
  INV_X1 U9785 ( .A(n8264), .ZN(n8266) );
  AOI21_X1 U9786 ( .B1(n8266), .B2(n4743), .A(n8831), .ZN(n8270) );
  OAI22_X1 U9787 ( .A1(n8268), .A2(n8859), .B1(n8424), .B2(n8861), .ZN(n8269)
         );
  AOI21_X1 U9788 ( .B1(n8270), .B2(n8267), .A(n8269), .ZN(n8903) );
  NOR2_X1 U9789 ( .A1(n8903), .A2(n8886), .ZN(n8271) );
  AOI211_X1 U9790 ( .C1(n8884), .C2(n8901), .A(n8272), .B(n8271), .ZN(n8273)
         );
  OAI21_X1 U9791 ( .B1(n8904), .B2(n8854), .A(n8273), .ZN(P2_U3268) );
  INV_X1 U9792 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8274) );
  NOR2_X1 U9793 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8274), .ZN(n8470) );
  OAI22_X1 U9794 ( .A1(n8439), .A2(P2_REG3_REG_3__SCAN_IN), .B1(n8441), .B2(
        n8275), .ZN(n8276) );
  AOI211_X1 U9795 ( .C1(n5823), .C2(n8445), .A(n8470), .B(n8276), .ZN(n8281)
         );
  OAI211_X1 U9796 ( .C1(n8279), .C2(n8277), .A(n8314), .B(n8278), .ZN(n8280)
         );
  OAI211_X1 U9797 ( .C1(n8282), .C2(n8440), .A(n8281), .B(n8280), .ZN(P2_U3220) );
  AOI21_X1 U9798 ( .B1(n8285), .B2(n8284), .A(n8283), .ZN(n8286) );
  NOR2_X1 U9799 ( .A1(n8286), .A2(n8447), .ZN(n8287) );
  AOI21_X1 U9800 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8288), .A(n8287), .ZN(
        n8292) );
  AOI22_X1 U9801 ( .A1(n8290), .A2(n7120), .B1(n8289), .B2(n8445), .ZN(n8291)
         );
  OAI211_X1 U9802 ( .C1(n8293), .C2(n8440), .A(n8292), .B(n8291), .ZN(P2_U3224) );
  NAND2_X1 U9803 ( .A1(n8295), .A2(n9534), .ZN(n9540) );
  INV_X1 U9804 ( .A(n9300), .ZN(n8298) );
  INV_X1 U9805 ( .A(n8296), .ZN(n8297) );
  AOI21_X1 U9806 ( .B1(n9536), .B2(n8298), .A(n8297), .ZN(n9537) );
  AOI22_X1 U9807 ( .A1(n8299), .A2(n9499), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9735), .ZN(n8300) );
  OAI21_X1 U9808 ( .B1(n8301), .B2(n9502), .A(n8300), .ZN(n8309) );
  OAI222_X1 U9809 ( .A1(n8307), .A2(n7743), .B1(n8306), .B2(n9477), .C1(n8305), 
        .C2(n9474), .ZN(n8308) );
  OAI21_X1 U9810 ( .B1(n9540), .B2(n9516), .A(n8310), .ZN(P1_U3263) );
  INV_X1 U9811 ( .A(n5859), .ZN(n8843) );
  OAI21_X1 U9812 ( .B1(n8313), .B2(n8312), .A(n8354), .ZN(n8315) );
  NAND2_X1 U9813 ( .A1(n8315), .A2(n8314), .ZN(n8319) );
  OAI22_X1 U9814 ( .A1(n8835), .A2(n8441), .B1(n8440), .B2(n8834), .ZN(n8316)
         );
  AOI211_X1 U9815 ( .C1(n8429), .C2(n8841), .A(n8317), .B(n8316), .ZN(n8318)
         );
  OAI211_X1 U9816 ( .C1(n8843), .C2(n8432), .A(n8319), .B(n8318), .ZN(P2_U3217) );
  XNOR2_X1 U9817 ( .A(n8320), .B(n8382), .ZN(n8326) );
  INV_X1 U9818 ( .A(n8693), .ZN(n8322) );
  OAI22_X1 U9819 ( .A1(n8439), .A2(n8322), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8321), .ZN(n8324) );
  OAI22_X1 U9820 ( .A1(n8349), .A2(n8441), .B1(n8440), .B2(n8340), .ZN(n8323)
         );
  AOI211_X1 U9821 ( .C1(n8926), .C2(n8445), .A(n8324), .B(n8323), .ZN(n8325)
         );
  OAI21_X1 U9822 ( .B1(n8326), .B2(n8447), .A(n8325), .ZN(P2_U3218) );
  INV_X1 U9823 ( .A(n8327), .ZN(n8328) );
  AOI21_X1 U9824 ( .B1(n8330), .B2(n8329), .A(n8328), .ZN(n8334) );
  OAI22_X1 U9825 ( .A1(n8339), .A2(n8859), .B1(n8372), .B2(n8861), .ZN(n8753)
         );
  AOI22_X1 U9826 ( .A1(n8376), .A2(n8753), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8331) );
  OAI21_X1 U9827 ( .B1(n8439), .B2(n8762), .A(n8331), .ZN(n8332) );
  AOI21_X1 U9828 ( .B1(n8948), .B2(n8445), .A(n8332), .ZN(n8333) );
  OAI21_X1 U9829 ( .B1(n8334), .B2(n8447), .A(n8333), .ZN(P2_U3221) );
  XNOR2_X1 U9830 ( .A(n8335), .B(n8336), .ZN(n8344) );
  INV_X1 U9831 ( .A(n8723), .ZN(n8338) );
  OAI22_X1 U9832 ( .A1(n8439), .A2(n8338), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8337), .ZN(n8342) );
  OAI22_X1 U9833 ( .A1(n8340), .A2(n8441), .B1(n8440), .B2(n8339), .ZN(n8341)
         );
  AOI211_X1 U9834 ( .C1(n8936), .C2(n8445), .A(n8342), .B(n8341), .ZN(n8343)
         );
  OAI21_X1 U9835 ( .B1(n8344), .B2(n8447), .A(n8343), .ZN(P2_U3225) );
  XOR2_X1 U9836 ( .A(n8347), .B(n8346), .Z(n8348) );
  XNOR2_X1 U9837 ( .A(n8345), .B(n8348), .ZN(n8353) );
  OAI22_X1 U9838 ( .A1(n8631), .A2(n8859), .B1(n8349), .B2(n8861), .ZN(n8657)
         );
  AOI22_X1 U9839 ( .A1(n8657), .A2(n8376), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8350) );
  OAI21_X1 U9840 ( .B1(n8663), .B2(n8439), .A(n8350), .ZN(n8351) );
  AOI21_X1 U9841 ( .B1(n8916), .B2(n8445), .A(n8351), .ZN(n8352) );
  OAI21_X1 U9842 ( .B1(n8353), .B2(n8447), .A(n8352), .ZN(P2_U3227) );
  INV_X1 U9843 ( .A(n8354), .ZN(n8356) );
  NOR2_X1 U9844 ( .A1(n8356), .A2(n8355), .ZN(n8357) );
  NAND2_X1 U9845 ( .A1(n8357), .A2(n8358), .ZN(n8435) );
  INV_X1 U9846 ( .A(n8435), .ZN(n8362) );
  INV_X1 U9847 ( .A(n8357), .ZN(n8360) );
  INV_X1 U9848 ( .A(n8358), .ZN(n8359) );
  NAND2_X1 U9849 ( .A1(n8360), .A2(n8359), .ZN(n8434) );
  OAI211_X1 U9850 ( .C1(n8362), .C2(n8437), .A(n8434), .B(n8361), .ZN(n8364)
         );
  AOI21_X1 U9851 ( .B1(n8364), .B2(n8363), .A(n8447), .ZN(n8365) );
  INV_X1 U9852 ( .A(n8365), .ZN(n8370) );
  INV_X1 U9853 ( .A(n8366), .ZN(n8802) );
  OAI22_X1 U9854 ( .A1(n8835), .A2(n8440), .B1(n8441), .B2(n8415), .ZN(n8367)
         );
  AOI211_X1 U9855 ( .C1(n8429), .C2(n8802), .A(n8368), .B(n8367), .ZN(n8369)
         );
  OAI211_X1 U9856 ( .C1(n8804), .C2(n8432), .A(n8370), .B(n8369), .ZN(P2_U3228) );
  XNOR2_X1 U9857 ( .A(n8371), .B(n8410), .ZN(n8380) );
  OR2_X1 U9858 ( .A1(n8372), .A2(n8859), .ZN(n8374) );
  NAND2_X1 U9859 ( .A1(n8818), .A2(n8819), .ZN(n8373) );
  NAND2_X1 U9860 ( .A1(n8374), .A2(n8373), .ZN(n8784) );
  AOI21_X1 U9861 ( .B1(n8376), .B2(n8784), .A(n8375), .ZN(n8377) );
  OAI21_X1 U9862 ( .B1(n8439), .B2(n8788), .A(n8377), .ZN(n8378) );
  AOI21_X1 U9863 ( .B1(n8958), .B2(n8445), .A(n8378), .ZN(n8379) );
  OAI21_X1 U9864 ( .B1(n8380), .B2(n8447), .A(n8379), .ZN(P2_U3230) );
  OAI21_X1 U9865 ( .B1(n8320), .B2(n8382), .A(n8381), .ZN(n8386) );
  XOR2_X1 U9866 ( .A(n8384), .B(n8383), .Z(n8385) );
  XNOR2_X1 U9867 ( .A(n8386), .B(n8385), .ZN(n8391) );
  OAI22_X1 U9868 ( .A1(n8439), .A2(n8683), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8387), .ZN(n8389) );
  OAI22_X1 U9869 ( .A1(n8680), .A2(n8441), .B1(n8440), .B2(n8405), .ZN(n8388)
         );
  AOI211_X1 U9870 ( .C1(n8923), .C2(n8445), .A(n8389), .B(n8388), .ZN(n8390)
         );
  OAI21_X1 U9871 ( .B1(n8391), .B2(n8447), .A(n8390), .ZN(P2_U3231) );
  XNOR2_X1 U9872 ( .A(n8392), .B(n8393), .ZN(n8397) );
  OAI22_X1 U9873 ( .A1(n8439), .A2(n8740), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10018), .ZN(n8395) );
  OAI22_X1 U9874 ( .A1(n8736), .A2(n8441), .B1(n8440), .B2(n8735), .ZN(n8394)
         );
  AOI211_X1 U9875 ( .C1(n8942), .C2(n8445), .A(n8395), .B(n8394), .ZN(n8396)
         );
  OAI21_X1 U9876 ( .B1(n8397), .B2(n8447), .A(n8396), .ZN(P2_U3235) );
  NAND2_X1 U9877 ( .A1(n8399), .A2(n8398), .ZN(n8403) );
  XNOR2_X1 U9878 ( .A(n8401), .B(n8400), .ZN(n8402) );
  XNOR2_X1 U9879 ( .A(n8403), .B(n8402), .ZN(n8409) );
  OAI22_X1 U9880 ( .A1(n8439), .A2(n8706), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8404), .ZN(n8407) );
  OAI22_X1 U9881 ( .A1(n8405), .A2(n8441), .B1(n8440), .B2(n8736), .ZN(n8406)
         );
  AOI211_X1 U9882 ( .C1(n8931), .C2(n8445), .A(n8407), .B(n8406), .ZN(n8408)
         );
  OAI21_X1 U9883 ( .B1(n8409), .B2(n8447), .A(n8408), .ZN(P2_U3237) );
  OR2_X1 U9884 ( .A1(n8371), .A2(n8410), .ZN(n8412) );
  NAND2_X1 U9885 ( .A1(n8412), .A2(n8411), .ZN(n8414) );
  XNOR2_X1 U9886 ( .A(n8414), .B(n8413), .ZN(n8419) );
  NOR2_X1 U9887 ( .A1(n10037), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9816) );
  OAI22_X1 U9888 ( .A1(n8415), .A2(n8440), .B1(n8441), .B2(n8735), .ZN(n8416)
         );
  AOI211_X1 U9889 ( .C1(n8429), .C2(n8778), .A(n9816), .B(n8416), .ZN(n8418)
         );
  NAND2_X1 U9890 ( .A1(n8952), .A2(n8445), .ZN(n8417) );
  OAI211_X1 U9891 ( .C1(n8419), .C2(n8447), .A(n8418), .B(n8417), .ZN(P2_U3240) );
  INV_X1 U9892 ( .A(n8911), .ZN(n8433) );
  AOI21_X1 U9893 ( .B1(n8421), .B2(n8420), .A(n8447), .ZN(n8423) );
  NAND2_X1 U9894 ( .A1(n8423), .A2(n8422), .ZN(n8431) );
  OAI22_X1 U9895 ( .A1(n8424), .A2(n8859), .B1(n8680), .B2(n8861), .ZN(n8645)
         );
  INV_X1 U9896 ( .A(n8645), .ZN(n8427) );
  OAI22_X1 U9897 ( .A1(n8427), .A2(n8426), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8425), .ZN(n8428) );
  AOI21_X1 U9898 ( .B1(n8648), .B2(n8429), .A(n8428), .ZN(n8430) );
  OAI211_X1 U9899 ( .C1(n8433), .C2(n8432), .A(n8431), .B(n8430), .ZN(P2_U3242) );
  NAND2_X1 U9900 ( .A1(n8435), .A2(n8434), .ZN(n8436) );
  XOR2_X1 U9901 ( .A(n8437), .B(n8436), .Z(n8448) );
  OAI21_X1 U9902 ( .B1(n8439), .B2(n8822), .A(n8438), .ZN(n8444) );
  OAI22_X1 U9903 ( .A1(n8442), .A2(n8441), .B1(n8440), .B2(n8860), .ZN(n8443)
         );
  AOI211_X1 U9904 ( .C1(n8968), .C2(n8445), .A(n8444), .B(n8443), .ZN(n8446)
         );
  OAI21_X1 U9905 ( .B1(n8448), .B2(n8447), .A(n8446), .ZN(P2_U3243) );
  MUX2_X1 U9906 ( .A(n8599), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8464), .Z(
        P2_U3582) );
  MUX2_X1 U9907 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8601), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9908 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8449), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9909 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8450), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9910 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8451), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9911 ( .A(n8690), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8464), .Z(
        P2_U3576) );
  MUX2_X1 U9912 ( .A(n8713), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8464), .Z(
        P2_U3575) );
  MUX2_X1 U9913 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8727), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9914 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8714), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9915 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8728), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9916 ( .A(n8776), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8464), .Z(
        P2_U3571) );
  MUX2_X1 U9917 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8452), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9918 ( .A(n8800), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8464), .Z(
        P2_U3569) );
  MUX2_X1 U9919 ( .A(n8818), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8464), .Z(
        P2_U3568) );
  MUX2_X1 U9920 ( .A(n8799), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8464), .Z(
        P2_U3567) );
  MUX2_X1 U9921 ( .A(n8820), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8464), .Z(
        P2_U3566) );
  MUX2_X1 U9922 ( .A(n8453), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8464), .Z(
        P2_U3565) );
  MUX2_X1 U9923 ( .A(n8454), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8464), .Z(
        P2_U3564) );
  MUX2_X1 U9924 ( .A(n8455), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8464), .Z(
        P2_U3563) );
  MUX2_X1 U9925 ( .A(n8456), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8464), .Z(
        P2_U3562) );
  MUX2_X1 U9926 ( .A(n8457), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8464), .Z(
        P2_U3561) );
  MUX2_X1 U9927 ( .A(n8458), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8464), .Z(
        P2_U3560) );
  MUX2_X1 U9928 ( .A(n8459), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8464), .Z(
        P2_U3559) );
  MUX2_X1 U9929 ( .A(n8460), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8464), .Z(
        P2_U3558) );
  MUX2_X1 U9930 ( .A(n8461), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8464), .Z(
        P2_U3557) );
  MUX2_X1 U9931 ( .A(n8462), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8464), .Z(
        P2_U3556) );
  MUX2_X1 U9932 ( .A(n8463), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8464), .Z(
        P2_U3555) );
  MUX2_X1 U9933 ( .A(n7120), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8464), .Z(
        P2_U3554) );
  MUX2_X1 U9934 ( .A(n7229), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8464), .Z(
        P2_U3553) );
  MUX2_X1 U9935 ( .A(n8465), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8464), .Z(
        P2_U3552) );
  OR3_X1 U9936 ( .A1(n8468), .A2(n8467), .A3(n8466), .ZN(n8469) );
  NAND3_X1 U9937 ( .A1(n8579), .A2(n8481), .A3(n8469), .ZN(n8478) );
  AOI21_X1 U9938 ( .B1(n9817), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8470), .ZN(
        n8477) );
  NAND2_X1 U9939 ( .A1(n9821), .A2(n8471), .ZN(n8476) );
  OAI211_X1 U9940 ( .C1(n8474), .C2(n8473), .A(n9823), .B(n8472), .ZN(n8475)
         );
  NAND4_X1 U9941 ( .A1(n8478), .A2(n8477), .A3(n8476), .A4(n8475), .ZN(
        P2_U3248) );
  INV_X1 U9942 ( .A(n8496), .ZN(n8483) );
  NAND3_X1 U9943 ( .A1(n8481), .A2(n8480), .A3(n8479), .ZN(n8482) );
  NAND3_X1 U9944 ( .A1(n8579), .A2(n8483), .A3(n8482), .ZN(n8493) );
  INV_X1 U9945 ( .A(n8484), .ZN(n8485) );
  AOI21_X1 U9946 ( .B1(n9817), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8485), .ZN(
        n8492) );
  NAND2_X1 U9947 ( .A1(n9821), .A2(n8486), .ZN(n8491) );
  OAI211_X1 U9948 ( .C1(n8489), .C2(n8488), .A(n9823), .B(n8487), .ZN(n8490)
         );
  NAND4_X1 U9949 ( .A1(n8493), .A2(n8492), .A3(n8491), .A4(n8490), .ZN(
        P2_U3249) );
  OR3_X1 U9950 ( .A1(n8496), .A2(n8495), .A3(n8494), .ZN(n8497) );
  NAND3_X1 U9951 ( .A1(n8579), .A2(n8509), .A3(n8497), .ZN(n8506) );
  NOR2_X1 U9952 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5090), .ZN(n8498) );
  AOI21_X1 U9953 ( .B1(n9817), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8498), .ZN(
        n8505) );
  NAND2_X1 U9954 ( .A1(n9821), .A2(n8499), .ZN(n8504) );
  OAI211_X1 U9955 ( .C1(n8502), .C2(n8501), .A(n9823), .B(n8500), .ZN(n8503)
         );
  NAND4_X1 U9956 ( .A1(n8506), .A2(n8505), .A3(n8504), .A4(n8503), .ZN(
        P2_U3250) );
  INV_X1 U9957 ( .A(n8524), .ZN(n8511) );
  NAND3_X1 U9958 ( .A1(n8509), .A2(n8508), .A3(n8507), .ZN(n8510) );
  NAND3_X1 U9959 ( .A1(n8579), .A2(n8511), .A3(n8510), .ZN(n8521) );
  INV_X1 U9960 ( .A(n8512), .ZN(n8513) );
  AOI21_X1 U9961 ( .B1(n9817), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8513), .ZN(
        n8520) );
  NAND2_X1 U9962 ( .A1(n9821), .A2(n8514), .ZN(n8519) );
  OAI211_X1 U9963 ( .C1(n8517), .C2(n8516), .A(n9823), .B(n8515), .ZN(n8518)
         );
  NAND4_X1 U9964 ( .A1(n8521), .A2(n8520), .A3(n8519), .A4(n8518), .ZN(
        P2_U3251) );
  INV_X1 U9965 ( .A(n8546), .ZN(n8526) );
  NOR3_X1 U9966 ( .A1(n8524), .A2(n8523), .A3(n8522), .ZN(n8525) );
  NOR3_X1 U9967 ( .A1(n9827), .A2(n8526), .A3(n8525), .ZN(n8527) );
  AOI21_X1 U9968 ( .B1(n9821), .B2(n8528), .A(n8527), .ZN(n8536) );
  NOR2_X1 U9969 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8529), .ZN(n8530) );
  AOI21_X1 U9970 ( .B1(n9817), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8530), .ZN(
        n8535) );
  OAI211_X1 U9971 ( .C1(n8533), .C2(n8532), .A(n9823), .B(n8531), .ZN(n8534)
         );
  NAND3_X1 U9972 ( .A1(n8536), .A2(n8535), .A3(n8534), .ZN(P2_U3252) );
  INV_X1 U9973 ( .A(n8537), .ZN(n8540) );
  NOR2_X1 U9974 ( .A1(n9805), .A2(n8538), .ZN(n8539) );
  AOI211_X1 U9975 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n9817), .A(n8540), .B(
        n8539), .ZN(n8551) );
  OAI211_X1 U9976 ( .C1(n8543), .C2(n8542), .A(n9823), .B(n8541), .ZN(n8550)
         );
  INV_X1 U9977 ( .A(n8554), .ZN(n8548) );
  NAND3_X1 U9978 ( .A1(n8546), .A2(n8545), .A3(n8544), .ZN(n8547) );
  NAND3_X1 U9979 ( .A1(n8548), .A2(n8579), .A3(n8547), .ZN(n8549) );
  NAND3_X1 U9980 ( .A1(n8551), .A2(n8550), .A3(n8549), .ZN(P2_U3253) );
  OR3_X1 U9981 ( .A1(n8554), .A2(n8553), .A3(n8552), .ZN(n8555) );
  NAND3_X1 U9982 ( .A1(n8556), .A2(n8579), .A3(n8555), .ZN(n8566) );
  NOR2_X1 U9983 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8557), .ZN(n8558) );
  AOI21_X1 U9984 ( .B1(n9817), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8558), .ZN(
        n8565) );
  OAI211_X1 U9985 ( .C1(n8561), .C2(n8560), .A(n9823), .B(n8559), .ZN(n8564)
         );
  NAND2_X1 U9986 ( .A1(n9821), .A2(n8562), .ZN(n8563) );
  NAND4_X1 U9987 ( .A1(n8566), .A2(n8565), .A3(n8564), .A4(n8563), .ZN(
        P2_U3254) );
  NAND2_X1 U9988 ( .A1(n8572), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8568) );
  NOR2_X1 U9989 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n9815), .ZN(n9814) );
  NOR2_X1 U9990 ( .A1(n9822), .A2(n8569), .ZN(n8570) );
  INV_X1 U9991 ( .A(n8580), .ZN(n8577) );
  AOI22_X1 U9992 ( .A1(n9822), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8574), .B2(
        n8573), .ZN(n9819) );
  NAND2_X1 U9993 ( .A1(n9820), .A2(n9819), .ZN(n9818) );
  OAI21_X1 U9994 ( .B1(n9822), .B2(P2_REG1_REG_18__SCAN_IN), .A(n9818), .ZN(
        n8575) );
  XNOR2_X1 U9995 ( .A(n8575), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8578) );
  OAI21_X1 U9996 ( .B1(n8578), .B2(n9807), .A(n9805), .ZN(n8576) );
  AOI21_X1 U9997 ( .B1(n8577), .B2(n8579), .A(n8576), .ZN(n8582) );
  AOI22_X1 U9998 ( .A1(n8580), .A2(n8579), .B1(n9823), .B2(n8578), .ZN(n8581)
         );
  NAND2_X1 U9999 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8583) );
  OAI211_X1 U10000 ( .C1(n8585), .C2(n4457), .A(n8584), .B(n8583), .ZN(
        P2_U3264) );
  NAND2_X1 U10001 ( .A1(n4406), .A2(n8605), .ZN(n8607) );
  NAND2_X1 U10002 ( .A1(n8592), .A2(n8593), .ZN(n8591) );
  INV_X1 U10003 ( .A(P2_B_REG_SCAN_IN), .ZN(n8586) );
  NOR2_X1 U10004 ( .A1(n9030), .A2(n8586), .ZN(n8587) );
  NOR2_X1 U10005 ( .A1(n8859), .A2(n8587), .ZN(n8600) );
  NAND2_X1 U10006 ( .A1(n8600), .A2(n8588), .ZN(n8891) );
  NOR2_X1 U10007 ( .A1(n8886), .A2(n8891), .ZN(n8595) );
  AOI21_X1 U10008 ( .B1(n8886), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8595), .ZN(
        n8590) );
  NAND2_X1 U10009 ( .A1(n5774), .A2(n8765), .ZN(n8589) );
  OAI211_X1 U10010 ( .C1(n8888), .C2(n8687), .A(n8590), .B(n8589), .ZN(
        P2_U3265) );
  OAI21_X1 U10011 ( .B1(n8592), .B2(n8593), .A(n8591), .ZN(n8892) );
  NOR2_X1 U10012 ( .A1(n8593), .A2(n8879), .ZN(n8594) );
  AOI211_X1 U10013 ( .C1(n8886), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8595), .B(
        n8594), .ZN(n8596) );
  OAI21_X1 U10014 ( .B1(n8687), .B2(n8892), .A(n8596), .ZN(P2_U3266) );
  NOR2_X1 U10015 ( .A1(n8900), .A2(n8601), .ZN(n8896) );
  NOR2_X1 U10016 ( .A1(n8893), .A2(n8896), .ZN(n8597) );
  XNOR2_X1 U10017 ( .A(n8597), .B(n4626), .ZN(n8616) );
  INV_X1 U10018 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8608) );
  OAI22_X1 U10019 ( .A1(n8609), .A2(n8761), .B1(n8608), .B2(n8772), .ZN(n8610)
         );
  AOI21_X1 U10020 ( .B1(n8611), .B2(n8765), .A(n8610), .ZN(n8612) );
  OAI21_X1 U10021 ( .B1(n8895), .B2(n8687), .A(n8612), .ZN(n8613) );
  AOI21_X1 U10022 ( .B1(n8614), .B2(n8772), .A(n8613), .ZN(n8615) );
  OAI21_X1 U10023 ( .B1(n8616), .B2(n8854), .A(n8615), .ZN(P2_U3267) );
  INV_X1 U10024 ( .A(n8617), .ZN(n8619) );
  AOI21_X1 U10025 ( .B1(n8619), .B2(n4552), .A(n8618), .ZN(n8909) );
  INV_X1 U10026 ( .A(n8620), .ZN(n8621) );
  AOI21_X1 U10027 ( .B1(n8905), .B2(n4298), .A(n8621), .ZN(n8906) );
  INV_X1 U10028 ( .A(n8622), .ZN(n8623) );
  AOI22_X1 U10029 ( .A1(n8623), .A2(n8876), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8886), .ZN(n8624) );
  OAI21_X1 U10030 ( .B1(n8625), .B2(n8879), .A(n8624), .ZN(n8636) );
  NAND2_X1 U10031 ( .A1(n8626), .A2(n8655), .ZN(n8659) );
  NAND3_X1 U10032 ( .A1(n8659), .A2(n4551), .A3(n8642), .ZN(n8643) );
  AOI21_X1 U10033 ( .B1(n8643), .B2(n8627), .A(n4552), .ZN(n8630) );
  INV_X1 U10034 ( .A(n8628), .ZN(n8629) );
  NOR3_X1 U10035 ( .A1(n8630), .A2(n8629), .A3(n8831), .ZN(n8634) );
  OAI22_X1 U10036 ( .A1(n8632), .A2(n8859), .B1(n8631), .B2(n8861), .ZN(n8633)
         );
  NOR2_X1 U10037 ( .A1(n8634), .A2(n8633), .ZN(n8908) );
  NOR2_X1 U10038 ( .A1(n8908), .A2(n8886), .ZN(n8635) );
  AOI211_X1 U10039 ( .C1(n8906), .C2(n8884), .A(n8636), .B(n8635), .ZN(n8637)
         );
  OAI21_X1 U10040 ( .B1(n8909), .B2(n8854), .A(n8637), .ZN(P2_U3269) );
  OAI21_X1 U10041 ( .B1(n8640), .B2(n8639), .A(n8638), .ZN(n8641) );
  INV_X1 U10042 ( .A(n8641), .ZN(n8914) );
  AND2_X1 U10043 ( .A1(n8659), .A2(n8642), .ZN(n8644) );
  OAI21_X1 U10044 ( .B1(n8644), .B2(n4551), .A(n8643), .ZN(n8646) );
  AOI21_X1 U10045 ( .B1(n8646), .B2(n8871), .A(n8645), .ZN(n8913) );
  AOI21_X1 U10046 ( .B1(n8660), .B2(n8911), .A(n9907), .ZN(n8647) );
  AOI22_X1 U10047 ( .A1(n8910), .A2(n8758), .B1(n8876), .B2(n8648), .ZN(n8649)
         );
  AOI21_X1 U10048 ( .B1(n8913), .B2(n8649), .A(n8886), .ZN(n8650) );
  INV_X1 U10049 ( .A(n8650), .ZN(n8652) );
  AOI22_X1 U10050 ( .A1(n8911), .A2(n8765), .B1(P2_REG2_REG_26__SCAN_IN), .B2(
        n8886), .ZN(n8651) );
  OAI211_X1 U10051 ( .C1(n8914), .C2(n8854), .A(n8652), .B(n8651), .ZN(
        P2_U3270) );
  NOR2_X1 U10052 ( .A1(n8655), .A2(n4925), .ZN(n8656) );
  AOI21_X1 U10053 ( .B1(n8653), .B2(n8656), .A(n8831), .ZN(n8658) );
  AOI21_X1 U10054 ( .B1(n8659), .B2(n8658), .A(n8657), .ZN(n8918) );
  INV_X1 U10055 ( .A(n8682), .ZN(n8662) );
  INV_X1 U10056 ( .A(n8660), .ZN(n8661) );
  AOI211_X1 U10057 ( .C1(n8916), .C2(n8662), .A(n9907), .B(n8661), .ZN(n8915)
         );
  INV_X1 U10058 ( .A(n8663), .ZN(n8664) );
  AOI22_X1 U10059 ( .A1(n8664), .A2(n8876), .B1(n8886), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8665) );
  OAI21_X1 U10060 ( .B1(n8666), .B2(n8879), .A(n8665), .ZN(n8672) );
  OAI21_X1 U10061 ( .B1(n8669), .B2(n8668), .A(n8667), .ZN(n8670) );
  INV_X1 U10062 ( .A(n8670), .ZN(n8919) );
  NOR2_X1 U10063 ( .A1(n8919), .A2(n8854), .ZN(n8671) );
  AOI211_X1 U10064 ( .C1(n8915), .C2(n8796), .A(n8672), .B(n8671), .ZN(n8673)
         );
  OAI21_X1 U10065 ( .B1(n8886), .B2(n8918), .A(n8673), .ZN(P2_U3271) );
  XNOR2_X1 U10066 ( .A(n8674), .B(n4543), .ZN(n8925) );
  AND2_X1 U10067 ( .A1(n8675), .A2(n8676), .ZN(n8677) );
  NAND2_X1 U10068 ( .A1(n8713), .A2(n8819), .ZN(n8679) );
  AND2_X1 U10069 ( .A1(n8923), .A2(n8692), .ZN(n8681) );
  OR2_X1 U10070 ( .A1(n8682), .A2(n8681), .ZN(n8920) );
  INV_X1 U10071 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8684) );
  OAI22_X1 U10072 ( .A1(n8772), .A2(n8684), .B1(n8683), .B2(n8761), .ZN(n8685)
         );
  AOI21_X1 U10073 ( .B1(n8923), .B2(n8765), .A(n8685), .ZN(n8686) );
  OAI21_X1 U10074 ( .B1(n8920), .B2(n8687), .A(n8686), .ZN(n8688) );
  AOI21_X1 U10075 ( .B1(n8921), .B2(n8772), .A(n8688), .ZN(n8689) );
  OAI21_X1 U10076 ( .B1(n8854), .B2(n8925), .A(n8689), .ZN(P2_U3272) );
  OAI21_X1 U10077 ( .B1(n4287), .B2(n8696), .A(n8675), .ZN(n8691) );
  AOI222_X1 U10078 ( .A1(n8871), .A2(n8691), .B1(n8727), .B2(n8819), .C1(n8690), .C2(n8817), .ZN(n8929) );
  AOI21_X1 U10079 ( .B1(n8926), .B2(n8704), .A(n8260), .ZN(n8927) );
  AOI22_X1 U10080 ( .A1(n8886), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8693), .B2(
        n8876), .ZN(n8694) );
  OAI21_X1 U10081 ( .B1(n8695), .B2(n8879), .A(n8694), .ZN(n8701) );
  NAND2_X1 U10082 ( .A1(n8697), .A2(n8696), .ZN(n8698) );
  NAND2_X1 U10083 ( .A1(n8699), .A2(n8698), .ZN(n8930) );
  NOR2_X1 U10084 ( .A1(n8930), .A2(n8854), .ZN(n8700) );
  AOI211_X1 U10085 ( .C1(n8927), .C2(n8884), .A(n8701), .B(n8700), .ZN(n8702)
         );
  OAI21_X1 U10086 ( .B1(n8929), .B2(n8886), .A(n8702), .ZN(P2_U3273) );
  XOR2_X1 U10087 ( .A(n8703), .B(n8712), .Z(n8935) );
  INV_X1 U10088 ( .A(n8704), .ZN(n8705) );
  AOI21_X1 U10089 ( .B1(n8931), .B2(n4859), .A(n8705), .ZN(n8932) );
  INV_X1 U10090 ( .A(n8706), .ZN(n8707) );
  AOI22_X1 U10091 ( .A1(n8886), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8707), .B2(
        n8876), .ZN(n8708) );
  OAI21_X1 U10092 ( .B1(n8709), .B2(n8879), .A(n8708), .ZN(n8718) );
  OAI211_X1 U10093 ( .C1(n8712), .C2(n8711), .A(n8710), .B(n8871), .ZN(n8716)
         );
  AOI22_X1 U10094 ( .A1(n8819), .A2(n8714), .B1(n8713), .B2(n8817), .ZN(n8715)
         );
  NOR2_X1 U10095 ( .A1(n8934), .A2(n8886), .ZN(n8717) );
  AOI211_X1 U10096 ( .C1(n8932), .C2(n8884), .A(n8718), .B(n8717), .ZN(n8719)
         );
  OAI21_X1 U10097 ( .B1(n8854), .B2(n8935), .A(n8719), .ZN(P2_U3274) );
  XNOR2_X1 U10098 ( .A(n8721), .B(n8720), .ZN(n8940) );
  AOI21_X1 U10099 ( .B1(n8936), .B2(n4970), .A(n8722), .ZN(n8937) );
  AOI22_X1 U10100 ( .A1(n8886), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8723), .B2(
        n8876), .ZN(n8724) );
  OAI21_X1 U10101 ( .B1(n4857), .B2(n8879), .A(n8724), .ZN(n8731) );
  OAI21_X1 U10102 ( .B1(n8726), .B2(n5422), .A(n8725), .ZN(n8729) );
  AOI222_X1 U10103 ( .A1(n8871), .A2(n8729), .B1(n8728), .B2(n8819), .C1(n8727), .C2(n8817), .ZN(n8939) );
  NOR2_X1 U10104 ( .A1(n8939), .A2(n8886), .ZN(n8730) );
  AOI211_X1 U10105 ( .C1(n8937), .C2(n8884), .A(n8731), .B(n8730), .ZN(n8732)
         );
  OAI21_X1 U10106 ( .B1(n8940), .B2(n8854), .A(n8732), .ZN(P2_U3275) );
  AOI21_X1 U10107 ( .B1(n8733), .B2(n8745), .A(n8831), .ZN(n8738) );
  OAI22_X1 U10108 ( .A1(n8736), .A2(n8859), .B1(n8735), .B2(n8861), .ZN(n8737)
         );
  AOI21_X1 U10109 ( .B1(n8738), .B2(n8734), .A(n8737), .ZN(n8945) );
  INV_X1 U10110 ( .A(n4970), .ZN(n8739) );
  AOI21_X1 U10111 ( .B1(n8942), .B2(n8755), .A(n8739), .ZN(n8943) );
  INV_X1 U10112 ( .A(n8942), .ZN(n8743) );
  INV_X1 U10113 ( .A(n8740), .ZN(n8741) );
  AOI22_X1 U10114 ( .A1(n8886), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8741), .B2(
        n8876), .ZN(n8742) );
  OAI21_X1 U10115 ( .B1(n8743), .B2(n8879), .A(n8742), .ZN(n8744) );
  AOI21_X1 U10116 ( .B1(n8943), .B2(n8884), .A(n8744), .ZN(n8749) );
  OR2_X1 U10117 ( .A1(n8746), .A2(n8745), .ZN(n8941) );
  NAND3_X1 U10118 ( .A1(n8941), .A2(n8811), .A3(n8747), .ZN(n8748) );
  OAI211_X1 U10119 ( .C1(n8945), .C2(n8886), .A(n8749), .B(n8748), .ZN(
        P2_U3276) );
  XNOR2_X1 U10120 ( .A(n8750), .B(n4469), .ZN(n8951) );
  XNOR2_X1 U10121 ( .A(n8751), .B(n8752), .ZN(n8754) );
  AOI21_X1 U10122 ( .B1(n8754), .B2(n8871), .A(n8753), .ZN(n8950) );
  INV_X1 U10123 ( .A(n8770), .ZN(n8757) );
  INV_X1 U10124 ( .A(n8755), .ZN(n8756) );
  AOI211_X1 U10125 ( .C1(n8948), .C2(n8757), .A(n9907), .B(n8756), .ZN(n8947)
         );
  NAND2_X1 U10126 ( .A1(n8947), .A2(n8758), .ZN(n8759) );
  OAI211_X1 U10127 ( .C1(n8951), .C2(n8867), .A(n8950), .B(n8759), .ZN(n8760)
         );
  NAND2_X1 U10128 ( .A1(n8760), .A2(n8772), .ZN(n8767) );
  INV_X1 U10129 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8763) );
  OAI22_X1 U10130 ( .A1(n8772), .A2(n8763), .B1(n8762), .B2(n8761), .ZN(n8764)
         );
  AOI21_X1 U10131 ( .B1(n8948), .B2(n8765), .A(n8764), .ZN(n8766) );
  OAI211_X1 U10132 ( .C1(n8951), .C2(n8881), .A(n8767), .B(n8766), .ZN(
        P2_U3277) );
  XOR2_X1 U10133 ( .A(n8768), .B(n8774), .Z(n8956) );
  AND2_X1 U10134 ( .A1(n8952), .A2(n4967), .ZN(n8769) );
  NOR2_X1 U10135 ( .A1(n8770), .A2(n8769), .ZN(n8953) );
  INV_X1 U10136 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8771) );
  OAI22_X1 U10137 ( .A1(n8773), .A2(n8879), .B1(n8772), .B2(n8771), .ZN(n8781)
         );
  XNOR2_X1 U10138 ( .A(n8775), .B(n8774), .ZN(n8777) );
  AOI222_X1 U10139 ( .A1(n8871), .A2(n8777), .B1(n8776), .B2(n8817), .C1(n8800), .C2(n8819), .ZN(n8955) );
  NAND2_X1 U10140 ( .A1(n8876), .A2(n8778), .ZN(n8779) );
  AOI21_X1 U10141 ( .B1(n8955), .B2(n8779), .A(n8886), .ZN(n8780) );
  AOI211_X1 U10142 ( .C1(n8953), .C2(n8884), .A(n8781), .B(n8780), .ZN(n8782)
         );
  OAI21_X1 U10143 ( .B1(n8956), .B2(n8854), .A(n8782), .ZN(P2_U3278) );
  XNOR2_X1 U10144 ( .A(n8783), .B(n4478), .ZN(n8785) );
  AOI21_X1 U10145 ( .B1(n8785), .B2(n8871), .A(n8784), .ZN(n8960) );
  INV_X1 U10146 ( .A(n4967), .ZN(n8786) );
  AOI211_X1 U10147 ( .C1(n8958), .C2(n8787), .A(n9907), .B(n8786), .ZN(n8957)
         );
  INV_X1 U10148 ( .A(n8788), .ZN(n8789) );
  AOI22_X1 U10149 ( .A1(n8886), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8789), .B2(
        n8876), .ZN(n8790) );
  OAI21_X1 U10150 ( .B1(n4419), .B2(n8879), .A(n8790), .ZN(n8795) );
  INV_X1 U10151 ( .A(n8791), .ZN(n8792) );
  AOI21_X1 U10152 ( .B1(n4478), .B2(n8793), .A(n8792), .ZN(n8961) );
  NOR2_X1 U10153 ( .A1(n8961), .A2(n8854), .ZN(n8794) );
  AOI211_X1 U10154 ( .C1(n8957), .C2(n8796), .A(n8795), .B(n8794), .ZN(n8797)
         );
  OAI21_X1 U10155 ( .B1(n8886), .B2(n8960), .A(n8797), .ZN(P2_U3279) );
  XOR2_X1 U10156 ( .A(n8798), .B(n8809), .Z(n8801) );
  AOI222_X1 U10157 ( .A1(n8871), .A2(n8801), .B1(n8800), .B2(n8817), .C1(n8799), .C2(n8819), .ZN(n8967) );
  XNOR2_X1 U10158 ( .A(n8962), .B(n4353), .ZN(n8963) );
  AOI22_X1 U10159 ( .A1(n8886), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8802), .B2(
        n8876), .ZN(n8803) );
  OAI21_X1 U10160 ( .B1(n8804), .B2(n8879), .A(n8803), .ZN(n8805) );
  AOI21_X1 U10161 ( .B1(n8963), .B2(n8884), .A(n8805), .ZN(n8813) );
  NAND2_X1 U10162 ( .A1(n8808), .A2(n8807), .ZN(n8810) );
  NAND2_X1 U10163 ( .A1(n8810), .A2(n8809), .ZN(n8964) );
  NAND3_X1 U10164 ( .A1(n8806), .A2(n8964), .A3(n8811), .ZN(n8812) );
  OAI211_X1 U10165 ( .C1(n8967), .C2(n8886), .A(n8813), .B(n8812), .ZN(
        P2_U3280) );
  NAND2_X1 U10166 ( .A1(n8814), .A2(n8863), .ZN(n8858) );
  NAND3_X1 U10167 ( .A1(n8858), .A2(n8239), .A3(n8830), .ZN(n8829) );
  NAND2_X1 U10168 ( .A1(n8829), .A2(n8815), .ZN(n8816) );
  XNOR2_X1 U10169 ( .A(n8816), .B(n4530), .ZN(n8821) );
  AOI222_X1 U10170 ( .A1(n8871), .A2(n8821), .B1(n8820), .B2(n8819), .C1(n8818), .C2(n8817), .ZN(n8971) );
  AOI21_X1 U10171 ( .B1(n8968), .B2(n8839), .A(n4353), .ZN(n8969) );
  INV_X1 U10172 ( .A(n8822), .ZN(n8823) );
  AOI22_X1 U10173 ( .A1(n8886), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8823), .B2(
        n8876), .ZN(n8824) );
  OAI21_X1 U10174 ( .B1(n4860), .B2(n8879), .A(n8824), .ZN(n8827) );
  XNOR2_X1 U10175 ( .A(n4304), .B(n8825), .ZN(n8972) );
  NOR2_X1 U10176 ( .A1(n8972), .A2(n8854), .ZN(n8826) );
  AOI211_X1 U10177 ( .C1(n8969), .C2(n8884), .A(n8827), .B(n8826), .ZN(n8828)
         );
  OAI21_X1 U10178 ( .B1(n8971), .B2(n8886), .A(n8828), .ZN(P2_U3281) );
  INV_X1 U10179 ( .A(n8829), .ZN(n8833) );
  AOI21_X1 U10180 ( .B1(n8858), .B2(n8830), .A(n8239), .ZN(n8832) );
  NOR3_X1 U10181 ( .A1(n8833), .A2(n8832), .A3(n8831), .ZN(n8837) );
  OAI22_X1 U10182 ( .A1(n8835), .A2(n8859), .B1(n8834), .B2(n8861), .ZN(n8836)
         );
  NOR2_X1 U10183 ( .A1(n8837), .A2(n8836), .ZN(n8975) );
  INV_X1 U10184 ( .A(n8839), .ZN(n8840) );
  AOI21_X1 U10185 ( .B1(n5859), .B2(n8838), .A(n8840), .ZN(n8973) );
  AOI22_X1 U10186 ( .A1(n8886), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8841), .B2(
        n8876), .ZN(n8842) );
  OAI21_X1 U10187 ( .B1(n8843), .B2(n8879), .A(n8842), .ZN(n8856) );
  INV_X1 U10188 ( .A(n8844), .ZN(n8845) );
  NAND2_X1 U10189 ( .A1(n8849), .A2(n8845), .ZN(n8864) );
  OR2_X1 U10190 ( .A1(n8864), .A2(n8863), .ZN(n8866) );
  INV_X1 U10191 ( .A(n8866), .ZN(n8847) );
  OAI21_X1 U10192 ( .B1(n8847), .B2(n8846), .A(n8239), .ZN(n8853) );
  NAND2_X1 U10193 ( .A1(n8849), .A2(n8848), .ZN(n8851) );
  NAND2_X1 U10194 ( .A1(n8851), .A2(n8850), .ZN(n8852) );
  NOR2_X1 U10195 ( .A1(n8976), .A2(n8854), .ZN(n8855) );
  AOI211_X1 U10196 ( .C1(n8973), .C2(n8884), .A(n8856), .B(n8855), .ZN(n8857)
         );
  OAI21_X1 U10197 ( .B1(n8886), .B2(n8975), .A(n8857), .ZN(P2_U3282) );
  OAI21_X1 U10198 ( .B1(n8814), .B2(n8863), .A(n8858), .ZN(n8870) );
  OAI22_X1 U10199 ( .A1(n8862), .A2(n8861), .B1(n8860), .B2(n8859), .ZN(n8869)
         );
  NAND2_X1 U10200 ( .A1(n8864), .A2(n8863), .ZN(n8865) );
  NAND2_X1 U10201 ( .A1(n8866), .A2(n8865), .ZN(n8981) );
  NOR2_X1 U10202 ( .A1(n8981), .A2(n8867), .ZN(n8868) );
  AOI211_X1 U10203 ( .C1(n8871), .C2(n8870), .A(n8869), .B(n8868), .ZN(n8980)
         );
  INV_X1 U10204 ( .A(n8872), .ZN(n8874) );
  INV_X1 U10205 ( .A(n8838), .ZN(n8873) );
  AOI21_X1 U10206 ( .B1(n8977), .B2(n8874), .A(n8873), .ZN(n8978) );
  INV_X1 U10207 ( .A(n8875), .ZN(n8877) );
  AOI22_X1 U10208 ( .A1(n8886), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8877), .B2(
        n8876), .ZN(n8878) );
  OAI21_X1 U10209 ( .B1(n8880), .B2(n8879), .A(n8878), .ZN(n8883) );
  NOR2_X1 U10210 ( .A1(n8981), .A2(n8881), .ZN(n8882) );
  AOI211_X1 U10211 ( .C1(n8978), .C2(n8884), .A(n8883), .B(n8882), .ZN(n8885)
         );
  OAI21_X1 U10212 ( .B1(n8980), .B2(n8886), .A(n8885), .ZN(P2_U3283) );
  NAND2_X1 U10213 ( .A1(n5774), .A2(n8988), .ZN(n8887) );
  OAI211_X1 U10214 ( .C1(n8888), .C2(n9907), .A(n8887), .B(n8891), .ZN(n8994)
         );
  MUX2_X1 U10215 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8994), .S(n9926), .Z(
        P2_U3551) );
  NAND2_X1 U10216 ( .A1(n8889), .A2(n8988), .ZN(n8890) );
  OAI211_X1 U10217 ( .C1(n8892), .C2(n9907), .A(n8891), .B(n8890), .ZN(n8995)
         );
  MUX2_X1 U10218 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8995), .S(n9926), .Z(
        P2_U3550) );
  NAND3_X1 U10219 ( .A1(n8893), .A2(n4626), .A3(n9902), .ZN(n8894) );
  INV_X1 U10220 ( .A(n8896), .ZN(n8897) );
  NOR3_X1 U10221 ( .A1(n8898), .A2(n8993), .A3(n8897), .ZN(n8899) );
  INV_X1 U10222 ( .A(n9907), .ZN(n9846) );
  AOI22_X1 U10223 ( .A1(n8901), .A2(n9846), .B1(n8988), .B2(n8900), .ZN(n8902)
         );
  OAI211_X1 U10224 ( .C1(n8904), .C2(n8993), .A(n8903), .B(n8902), .ZN(n8997)
         );
  MUX2_X1 U10225 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8997), .S(n9926), .Z(
        P2_U3548) );
  AOI22_X1 U10226 ( .A1(n8906), .A2(n9846), .B1(n8988), .B2(n8905), .ZN(n8907)
         );
  OAI211_X1 U10227 ( .C1(n8909), .C2(n8993), .A(n8908), .B(n8907), .ZN(n8998)
         );
  MUX2_X1 U10228 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8998), .S(n9926), .Z(
        P2_U3547) );
  AOI21_X1 U10229 ( .B1(n8988), .B2(n8911), .A(n8910), .ZN(n8912) );
  OAI211_X1 U10230 ( .C1(n8914), .C2(n8993), .A(n8913), .B(n8912), .ZN(n8999)
         );
  MUX2_X1 U10231 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8999), .S(n9926), .Z(
        P2_U3546) );
  AOI21_X1 U10232 ( .B1(n8988), .B2(n8916), .A(n8915), .ZN(n8917) );
  OAI211_X1 U10233 ( .C1(n8919), .C2(n8993), .A(n8918), .B(n8917), .ZN(n9000)
         );
  MUX2_X1 U10234 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9000), .S(n9926), .Z(
        P2_U3545) );
  NOR2_X1 U10235 ( .A1(n8920), .A2(n9907), .ZN(n8922) );
  AOI211_X1 U10236 ( .C1(n8988), .C2(n8923), .A(n8922), .B(n8921), .ZN(n8924)
         );
  MUX2_X1 U10237 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9001), .S(n9926), .Z(
        P2_U3544) );
  AOI22_X1 U10238 ( .A1(n8927), .A2(n9846), .B1(n8988), .B2(n8926), .ZN(n8928)
         );
  OAI211_X1 U10239 ( .C1(n8993), .C2(n8930), .A(n8929), .B(n8928), .ZN(n9002)
         );
  MUX2_X1 U10240 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9002), .S(n9926), .Z(
        P2_U3543) );
  AOI22_X1 U10241 ( .A1(n8932), .A2(n9846), .B1(n8988), .B2(n8931), .ZN(n8933)
         );
  OAI211_X1 U10242 ( .C1(n8935), .C2(n8993), .A(n8934), .B(n8933), .ZN(n9003)
         );
  MUX2_X1 U10243 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9003), .S(n9926), .Z(
        P2_U3542) );
  AOI22_X1 U10244 ( .A1(n8937), .A2(n9846), .B1(n8988), .B2(n8936), .ZN(n8938)
         );
  OAI211_X1 U10245 ( .C1(n8993), .C2(n8940), .A(n8939), .B(n8938), .ZN(n9004)
         );
  MUX2_X1 U10246 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9004), .S(n9926), .Z(
        P2_U3541) );
  NAND3_X1 U10247 ( .A1(n8941), .A2(n8747), .A3(n9902), .ZN(n8946) );
  AOI22_X1 U10248 ( .A1(n8943), .A2(n9846), .B1(n8988), .B2(n8942), .ZN(n8944)
         );
  NAND3_X1 U10249 ( .A1(n8946), .A2(n8945), .A3(n8944), .ZN(n9005) );
  MUX2_X1 U10250 ( .A(n9005), .B(P2_REG1_REG_20__SCAN_IN), .S(n9923), .Z(
        P2_U3540) );
  AOI21_X1 U10251 ( .B1(n8988), .B2(n8948), .A(n8947), .ZN(n8949) );
  OAI211_X1 U10252 ( .C1(n8951), .C2(n8993), .A(n8950), .B(n8949), .ZN(n9006)
         );
  MUX2_X1 U10253 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9006), .S(n9926), .Z(
        P2_U3539) );
  AOI22_X1 U10254 ( .A1(n8953), .A2(n9846), .B1(n8988), .B2(n8952), .ZN(n8954)
         );
  OAI211_X1 U10255 ( .C1(n8993), .C2(n8956), .A(n8955), .B(n8954), .ZN(n9007)
         );
  MUX2_X1 U10256 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9007), .S(n9926), .Z(
        P2_U3538) );
  AOI21_X1 U10257 ( .B1(n8988), .B2(n8958), .A(n8957), .ZN(n8959) );
  OAI211_X1 U10258 ( .C1(n8961), .C2(n8993), .A(n8960), .B(n8959), .ZN(n9008)
         );
  MUX2_X1 U10259 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9008), .S(n9926), .Z(
        P2_U3537) );
  AOI22_X1 U10260 ( .A1(n8963), .A2(n9846), .B1(n8988), .B2(n8962), .ZN(n8966)
         );
  NAND3_X1 U10261 ( .A1(n8806), .A2(n8964), .A3(n9902), .ZN(n8965) );
  NAND3_X1 U10262 ( .A1(n8967), .A2(n8966), .A3(n8965), .ZN(n9009) );
  MUX2_X1 U10263 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9009), .S(n9926), .Z(
        P2_U3536) );
  AOI22_X1 U10264 ( .A1(n8969), .A2(n9846), .B1(n8988), .B2(n8968), .ZN(n8970)
         );
  OAI211_X1 U10265 ( .C1(n8993), .C2(n8972), .A(n8971), .B(n8970), .ZN(n9010)
         );
  MUX2_X1 U10266 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9010), .S(n9926), .Z(
        P2_U3535) );
  AOI22_X1 U10267 ( .A1(n8973), .A2(n9846), .B1(n8988), .B2(n5859), .ZN(n8974)
         );
  OAI211_X1 U10268 ( .C1(n8993), .C2(n8976), .A(n8975), .B(n8974), .ZN(n9011)
         );
  MUX2_X1 U10269 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9011), .S(n9926), .Z(
        P2_U3534) );
  AOI22_X1 U10270 ( .A1(n8978), .A2(n9846), .B1(n8988), .B2(n8977), .ZN(n8979)
         );
  OAI211_X1 U10271 ( .C1(n9860), .C2(n8981), .A(n8980), .B(n8979), .ZN(n9012)
         );
  MUX2_X1 U10272 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9012), .S(n9926), .Z(
        P2_U3533) );
  AOI22_X1 U10273 ( .A1(n8983), .A2(n9846), .B1(n8988), .B2(n8982), .ZN(n8984)
         );
  OAI211_X1 U10274 ( .C1(n8993), .C2(n8986), .A(n8985), .B(n8984), .ZN(n9013)
         );
  MUX2_X1 U10275 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9013), .S(n9926), .Z(
        P2_U3532) );
  AOI22_X1 U10276 ( .A1(n8989), .A2(n9846), .B1(n8988), .B2(n8987), .ZN(n8990)
         );
  OAI211_X1 U10277 ( .C1(n8993), .C2(n8992), .A(n8991), .B(n8990), .ZN(n9014)
         );
  MUX2_X1 U10278 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9014), .S(n9926), .Z(
        P2_U3531) );
  MUX2_X1 U10279 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8994), .S(n9913), .Z(
        P2_U3519) );
  MUX2_X1 U10280 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8995), .S(n9913), .Z(
        P2_U3518) );
  MUX2_X1 U10281 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8997), .S(n9913), .Z(
        P2_U3516) );
  MUX2_X1 U10282 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8998), .S(n9913), .Z(
        P2_U3515) );
  MUX2_X1 U10283 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8999), .S(n9913), .Z(
        P2_U3514) );
  MUX2_X1 U10284 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9000), .S(n9913), .Z(
        P2_U3513) );
  MUX2_X1 U10285 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9002), .S(n9913), .Z(
        P2_U3511) );
  MUX2_X1 U10286 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9003), .S(n9913), .Z(
        P2_U3510) );
  MUX2_X1 U10287 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9004), .S(n9913), .Z(
        P2_U3509) );
  MUX2_X1 U10288 ( .A(n9005), .B(P2_REG0_REG_20__SCAN_IN), .S(n9912), .Z(
        P2_U3508) );
  MUX2_X1 U10289 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9006), .S(n9913), .Z(
        P2_U3507) );
  MUX2_X1 U10290 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9007), .S(n9913), .Z(
        P2_U3505) );
  MUX2_X1 U10291 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9008), .S(n9913), .Z(
        P2_U3502) );
  MUX2_X1 U10292 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9009), .S(n9913), .Z(
        P2_U3499) );
  MUX2_X1 U10293 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9010), .S(n9913), .Z(
        P2_U3496) );
  MUX2_X1 U10294 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9011), .S(n9913), .Z(
        P2_U3493) );
  MUX2_X1 U10295 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9012), .S(n9913), .Z(
        P2_U3490) );
  MUX2_X1 U10296 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n9013), .S(n9913), .Z(
        P2_U3487) );
  MUX2_X1 U10297 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9014), .S(n9913), .Z(
        P2_U3484) );
  INV_X1 U10298 ( .A(n5991), .ZN(n9662) );
  NOR4_X1 U10299 ( .A1(n9016), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9015), .A4(
        P2_U3152), .ZN(n9017) );
  AOI21_X1 U10300 ( .B1(n9026), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9017), .ZN(
        n9018) );
  OAI21_X1 U10301 ( .B1(n9662), .B2(n9038), .A(n9018), .ZN(P2_U3327) );
  INV_X1 U10302 ( .A(n9019), .ZN(n9665) );
  AOI22_X1 U10303 ( .A1(n9020), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9026), .ZN(n9021) );
  OAI21_X1 U10304 ( .B1(n9665), .B2(n9038), .A(n9021), .ZN(P2_U3328) );
  INV_X1 U10305 ( .A(n9022), .ZN(n9668) );
  AOI22_X1 U10306 ( .A1(n9023), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9026), .ZN(n9024) );
  OAI21_X1 U10307 ( .B1(n9668), .B2(n9038), .A(n9024), .ZN(P2_U3329) );
  INV_X1 U10308 ( .A(n9025), .ZN(n9671) );
  AOI22_X1 U10309 ( .A1(n9027), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n9026), .ZN(n9028) );
  OAI21_X1 U10310 ( .B1(n9671), .B2(n9038), .A(n9028), .ZN(P2_U3330) );
  INV_X1 U10311 ( .A(n9029), .ZN(n9674) );
  OAI222_X1 U10312 ( .A1(n9040), .A2(n9031), .B1(P2_U3152), .B2(n9030), .C1(
        n9038), .C2(n9674), .ZN(P2_U3331) );
  INV_X1 U10313 ( .A(n9032), .ZN(n9677) );
  OAI222_X1 U10314 ( .A1(n9034), .A2(P2_U3152), .B1(n9038), .B2(n9677), .C1(
        n9033), .C2(n9040), .ZN(P2_U3332) );
  OAI222_X1 U10315 ( .A1(n9040), .A2(n9039), .B1(n9038), .B2(n9037), .C1(n9036), .C2(P2_U3152), .ZN(P2_U3333) );
  MUX2_X1 U10316 ( .A(n9041), .B(n9813), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10317 ( .A(n9043), .ZN(n9045) );
  NAND2_X1 U10318 ( .A1(n9045), .A2(n9044), .ZN(n9090) );
  NAND2_X1 U10319 ( .A1(n9043), .A2(n9046), .ZN(n9092) );
  NAND2_X1 U10320 ( .A1(n9090), .A2(n9092), .ZN(n9048) );
  XNOR2_X1 U10321 ( .A(n9048), .B(n9047), .ZN(n9055) );
  NAND2_X1 U10322 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9236) );
  OAI21_X1 U10323 ( .B1(n9178), .B2(n9049), .A(n9236), .ZN(n9050) );
  AOI21_X1 U10324 ( .B1(n9180), .B2(n9458), .A(n9050), .ZN(n9051) );
  OAI21_X1 U10325 ( .B1(n9182), .B2(n9052), .A(n9051), .ZN(n9053) );
  AOI21_X1 U10326 ( .B1(n9606), .B2(n9184), .A(n9053), .ZN(n9054) );
  OAI21_X1 U10327 ( .B1(n9055), .B2(n9186), .A(n9054), .ZN(P1_U3213) );
  INV_X1 U10328 ( .A(n9118), .ZN(n9059) );
  AOI21_X1 U10329 ( .B1(n9056), .B2(n9117), .A(n9057), .ZN(n9058) );
  AOI21_X1 U10330 ( .B1(n9059), .B2(n9117), .A(n9058), .ZN(n9064) );
  NAND2_X1 U10331 ( .A1(n9362), .A2(n9180), .ZN(n9061) );
  AOI22_X1 U10332 ( .A1(n9392), .A2(n9155), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9060) );
  OAI211_X1 U10333 ( .C1(n9182), .C2(n9354), .A(n9061), .B(n9060), .ZN(n9062)
         );
  AOI21_X1 U10334 ( .B1(n9559), .B2(n9184), .A(n9062), .ZN(n9063) );
  OAI21_X1 U10335 ( .B1(n9064), .B2(n9186), .A(n9063), .ZN(P1_U3214) );
  XOR2_X1 U10336 ( .A(n9066), .B(n9065), .Z(n9071) );
  AOI22_X1 U10337 ( .A1(n9420), .A2(n9180), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3084), .ZN(n9068) );
  NAND2_X1 U10338 ( .A1(n9155), .A2(n9450), .ZN(n9067) );
  OAI211_X1 U10339 ( .C1(n9182), .C2(n9414), .A(n9068), .B(n9067), .ZN(n9069)
         );
  AOI21_X1 U10340 ( .B1(n9580), .B2(n9184), .A(n9069), .ZN(n9070) );
  OAI21_X1 U10341 ( .B1(n9071), .B2(n9186), .A(n9070), .ZN(P1_U3217) );
  XOR2_X1 U10342 ( .A(n9072), .B(n9073), .Z(n9079) );
  AOI22_X1 U10343 ( .A1(n9420), .A2(n9155), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9075) );
  NAND2_X1 U10344 ( .A1(n9167), .A2(n9384), .ZN(n9074) );
  OAI211_X1 U10345 ( .C1(n9076), .C2(n9152), .A(n9075), .B(n9074), .ZN(n9077)
         );
  AOI21_X1 U10346 ( .B1(n9570), .B2(n9184), .A(n9077), .ZN(n9078) );
  OAI21_X1 U10347 ( .B1(n9079), .B2(n9186), .A(n9078), .ZN(P1_U3221) );
  AOI21_X1 U10348 ( .B1(n9081), .B2(n9080), .A(n9163), .ZN(n9088) );
  NOR2_X1 U10349 ( .A1(n9326), .A2(n9182), .ZN(n9085) );
  OAI22_X1 U10350 ( .A1(n9083), .A2(n9178), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9082), .ZN(n9084) );
  AOI211_X1 U10351 ( .C1(n9180), .C2(n9334), .A(n9085), .B(n9084), .ZN(n9087)
         );
  NAND2_X1 U10352 ( .A1(n9550), .A2(n9184), .ZN(n9086) );
  OAI211_X1 U10353 ( .C1(n9088), .C2(n9186), .A(n9087), .B(n9086), .ZN(
        P1_U3223) );
  NAND2_X1 U10354 ( .A1(n9090), .A2(n9089), .ZN(n9093) );
  NAND3_X1 U10355 ( .A1(n9093), .A2(n9091), .A3(n9092), .ZN(n9174) );
  INV_X1 U10356 ( .A(n9174), .ZN(n9095) );
  NAND2_X1 U10357 ( .A1(n9093), .A2(n9092), .ZN(n9108) );
  NAND2_X1 U10358 ( .A1(n9108), .A2(n9094), .ZN(n9175) );
  OAI21_X1 U10359 ( .B1(n9095), .B2(n9176), .A(n9175), .ZN(n9099) );
  XNOR2_X1 U10360 ( .A(n9097), .B(n9096), .ZN(n9098) );
  XNOR2_X1 U10361 ( .A(n9099), .B(n9098), .ZN(n9104) );
  AOI22_X1 U10362 ( .A1(n9180), .A2(n9457), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n9101) );
  NAND2_X1 U10363 ( .A1(n9155), .A2(n9458), .ZN(n9100) );
  OAI211_X1 U10364 ( .C1(n9182), .C2(n9465), .A(n9101), .B(n9100), .ZN(n9102)
         );
  AOI21_X1 U10365 ( .B1(n9595), .B2(n9184), .A(n9102), .ZN(n9103) );
  OAI21_X1 U10366 ( .B1(n9104), .B2(n9186), .A(n9103), .ZN(P1_U3224) );
  INV_X1 U10367 ( .A(n9105), .ZN(n9107) );
  OAI21_X1 U10368 ( .B1(n9108), .B2(n9107), .A(n9106), .ZN(n9109) );
  XOR2_X1 U10369 ( .A(n9110), .B(n9109), .Z(n9115) );
  NAND2_X1 U10370 ( .A1(n9167), .A2(n9443), .ZN(n9112) );
  AOI22_X1 U10371 ( .A1(n9180), .A2(n9450), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n9111) );
  OAI211_X1 U10372 ( .C1(n9475), .C2(n9178), .A(n9112), .B(n9111), .ZN(n9113)
         );
  AOI21_X1 U10373 ( .B1(n9589), .B2(n9184), .A(n9113), .ZN(n9114) );
  OAI21_X1 U10374 ( .B1(n9115), .B2(n9186), .A(n9114), .ZN(P1_U3226) );
  AND3_X1 U10375 ( .A1(n9118), .A2(n9117), .A3(n9116), .ZN(n9119) );
  OAI21_X1 U10376 ( .B1(n9120), .B2(n9119), .A(n9165), .ZN(n9126) );
  OAI22_X1 U10377 ( .A1(n9122), .A2(n9178), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9121), .ZN(n9124) );
  NOR2_X1 U10378 ( .A1(n9169), .A2(n9152), .ZN(n9123) );
  AOI211_X1 U10379 ( .C1(n9342), .C2(n9167), .A(n9124), .B(n9123), .ZN(n9125)
         );
  OAI211_X1 U10380 ( .C1(n9344), .C2(n9173), .A(n9126), .B(n9125), .ZN(
        P1_U3227) );
  NAND2_X1 U10381 ( .A1(n9128), .A2(n9127), .ZN(n9129) );
  XNOR2_X1 U10382 ( .A(n9130), .B(n9129), .ZN(n9136) );
  OAI22_X1 U10383 ( .A1(n9142), .A2(n9152), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9131), .ZN(n9132) );
  AOI21_X1 U10384 ( .B1(n9155), .B2(n9436), .A(n9132), .ZN(n9133) );
  OAI21_X1 U10385 ( .B1(n9182), .B2(n9401), .A(n9133), .ZN(n9134) );
  AOI21_X1 U10386 ( .B1(n9574), .B2(n9184), .A(n9134), .ZN(n9135) );
  OAI21_X1 U10387 ( .B1(n9136), .B2(n9186), .A(n9135), .ZN(P1_U3231) );
  NAND2_X1 U10388 ( .A1(n9138), .A2(n9137), .ZN(n9139) );
  XOR2_X1 U10389 ( .A(n9140), .B(n9139), .Z(n9147) );
  OAI22_X1 U10390 ( .A1(n9142), .A2(n9178), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9141), .ZN(n9143) );
  AOI21_X1 U10391 ( .B1(n9377), .B2(n9180), .A(n9143), .ZN(n9144) );
  OAI21_X1 U10392 ( .B1(n9182), .B2(n9370), .A(n9144), .ZN(n9145) );
  AOI21_X1 U10393 ( .B1(n9564), .B2(n9184), .A(n9145), .ZN(n9146) );
  OAI21_X1 U10394 ( .B1(n9147), .B2(n9186), .A(n9146), .ZN(P1_U3233) );
  XNOR2_X1 U10395 ( .A(n9149), .B(n9148), .ZN(n9150) );
  XNOR2_X1 U10396 ( .A(n9151), .B(n9150), .ZN(n9159) );
  NAND2_X1 U10397 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9712) );
  OAI21_X1 U10398 ( .B1(n9153), .B2(n9152), .A(n9712), .ZN(n9154) );
  AOI21_X1 U10399 ( .B1(n9155), .B2(n9457), .A(n9154), .ZN(n9156) );
  OAI21_X1 U10400 ( .B1(n9182), .B2(n9428), .A(n9156), .ZN(n9157) );
  AOI21_X1 U10401 ( .B1(n9584), .B2(n9184), .A(n9157), .ZN(n9158) );
  OAI21_X1 U10402 ( .B1(n9159), .B2(n9186), .A(n9158), .ZN(P1_U3236) );
  OAI21_X1 U10403 ( .B1(n9163), .B2(n9162), .A(n9161), .ZN(n9164) );
  NAND3_X1 U10404 ( .A1(n9166), .A2(n9165), .A3(n9164), .ZN(n9172) );
  AOI22_X1 U10405 ( .A1(n9309), .A2(n9167), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9168) );
  OAI21_X1 U10406 ( .B1(n9169), .B2(n9178), .A(n9168), .ZN(n9170) );
  AOI21_X1 U10407 ( .B1(n9316), .B2(n9180), .A(n9170), .ZN(n9171) );
  OAI211_X1 U10408 ( .C1(n9311), .C2(n9173), .A(n9172), .B(n9171), .ZN(
        P1_U3238) );
  NAND2_X1 U10409 ( .A1(n9175), .A2(n9174), .ZN(n9177) );
  XNOR2_X1 U10410 ( .A(n9177), .B(n9176), .ZN(n9187) );
  NAND2_X1 U10411 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9246) );
  OAI21_X1 U10412 ( .B1(n9178), .B2(n9476), .A(n9246), .ZN(n9179) );
  AOI21_X1 U10413 ( .B1(n9180), .B2(n9448), .A(n9179), .ZN(n9181) );
  OAI21_X1 U10414 ( .B1(n9182), .B2(n9487), .A(n9181), .ZN(n9183) );
  AOI21_X1 U10415 ( .B1(n9599), .B2(n9184), .A(n9183), .ZN(n9185) );
  OAI21_X1 U10416 ( .B1(n9187), .B2(n9186), .A(n9185), .ZN(P1_U3239) );
  MUX2_X1 U10417 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9188), .S(n9200), .Z(
        P1_U3585) );
  MUX2_X1 U10418 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9189), .S(n9200), .Z(
        P1_U3584) );
  MUX2_X1 U10419 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9297), .S(n9200), .Z(
        P1_U3583) );
  MUX2_X1 U10420 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9316), .S(n9200), .Z(
        P1_U3582) );
  MUX2_X1 U10421 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9334), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10422 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9348), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10423 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9362), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10424 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9377), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10425 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9392), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10426 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9408), .S(n9200), .Z(
        P1_U3576) );
  MUX2_X1 U10427 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9420), .S(n9200), .Z(
        P1_U3575) );
  MUX2_X1 U10428 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9436), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10429 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9450), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10430 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9457), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10431 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9448), .S(n9200), .Z(
        P1_U3571) );
  MUX2_X1 U10432 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9458), .S(n9200), .Z(
        P1_U3570) );
  MUX2_X1 U10433 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9511), .S(n9200), .Z(
        P1_U3569) );
  MUX2_X1 U10434 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9190), .S(n9200), .Z(
        P1_U3568) );
  MUX2_X1 U10435 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9507), .S(n9200), .Z(
        P1_U3567) );
  MUX2_X1 U10436 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9191), .S(n9200), .Z(
        P1_U3566) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9192), .S(n9200), .Z(
        P1_U3565) );
  MUX2_X1 U10438 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9193), .S(n9200), .Z(
        P1_U3564) );
  MUX2_X1 U10439 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9194), .S(n9200), .Z(
        P1_U3563) );
  MUX2_X1 U10440 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9195), .S(n9200), .Z(
        P1_U3562) );
  MUX2_X1 U10441 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9196), .S(n9200), .Z(
        P1_U3561) );
  MUX2_X1 U10442 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9197), .S(n9200), .Z(
        P1_U3560) );
  MUX2_X1 U10443 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9198), .S(n9200), .Z(
        P1_U3559) );
  MUX2_X1 U10444 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n7530), .S(n9200), .Z(
        P1_U3558) );
  MUX2_X1 U10445 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9199), .S(n9200), .Z(
        P1_U3557) );
  MUX2_X1 U10446 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6587), .S(n9200), .Z(
        P1_U3556) );
  MUX2_X1 U10447 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9201), .S(n9200), .Z(
        P1_U3555) );
  XOR2_X1 U10448 ( .A(n9203), .B(n9202), .Z(n9204) );
  AOI22_X1 U10449 ( .A1(n9205), .A2(n9711), .B1(n9709), .B2(n9204), .ZN(n9211)
         );
  AOI22_X1 U10450 ( .A1(n9718), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(P1_U3084), 
        .B2(P1_REG3_REG_2__SCAN_IN), .ZN(n9210) );
  XOR2_X1 U10451 ( .A(n9207), .B(n9206), .Z(n9208) );
  NAND2_X1 U10452 ( .A1(n9719), .A2(n9208), .ZN(n9209) );
  NAND4_X1 U10453 ( .A1(n9212), .A2(n9211), .A3(n9210), .A4(n9209), .ZN(
        P1_U3243) );
  AOI211_X1 U10454 ( .C1(n9215), .C2(n9214), .A(n9213), .B(n9251), .ZN(n9216)
         );
  AOI21_X1 U10455 ( .B1(n9711), .B2(n9217), .A(n9216), .ZN(n9225) );
  OAI21_X1 U10456 ( .B1(n9220), .B2(n9219), .A(n9218), .ZN(n9221) );
  NAND2_X1 U10457 ( .A1(n9719), .A2(n9221), .ZN(n9223) );
  NAND2_X1 U10458 ( .A1(n9718), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9222) );
  NAND4_X1 U10459 ( .A1(n9225), .A2(n9224), .A3(n9223), .A4(n9222), .ZN(
        P1_U3247) );
  OAI21_X1 U10460 ( .B1(n9228), .B2(n9227), .A(n9226), .ZN(n9229) );
  NAND2_X1 U10461 ( .A1(n9229), .A2(n9719), .ZN(n9238) );
  AOI211_X1 U10462 ( .C1(n9232), .C2(n9231), .A(n9230), .B(n9251), .ZN(n9233)
         );
  AOI21_X1 U10463 ( .B1(n9711), .B2(n9234), .A(n9233), .ZN(n9237) );
  NAND2_X1 U10464 ( .A1(n9718), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n9235) );
  NAND4_X1 U10465 ( .A1(n9238), .A2(n9237), .A3(n9236), .A4(n9235), .ZN(
        P1_U3255) );
  AOI211_X1 U10466 ( .C1(n9240), .C2(n10016), .A(n9239), .B(n9251), .ZN(n9250)
         );
  INV_X1 U10467 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9248) );
  AOI211_X1 U10468 ( .C1(n9243), .C2(n9242), .A(n9241), .B(n9254), .ZN(n9244)
         );
  AOI21_X1 U10469 ( .B1(n9711), .B2(n9245), .A(n9244), .ZN(n9247) );
  OAI211_X1 U10470 ( .C1(n9281), .C2(n9248), .A(n9247), .B(n9246), .ZN(n9249)
         );
  OR2_X1 U10471 ( .A1(n9250), .A2(n9249), .ZN(P1_U3256) );
  AOI211_X1 U10472 ( .C1(n4311), .C2(n9253), .A(n9252), .B(n9251), .ZN(n9264)
         );
  AOI211_X1 U10473 ( .C1(n9257), .C2(n9256), .A(n9255), .B(n9254), .ZN(n9263)
         );
  NAND2_X1 U10474 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n9259) );
  NAND2_X1 U10475 ( .A1(n9718), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9258) );
  OAI211_X1 U10476 ( .C1(n9261), .C2(n9260), .A(n9259), .B(n9258), .ZN(n9262)
         );
  OR3_X1 U10477 ( .A1(n9264), .A2(n9263), .A3(n9262), .ZN(P1_U3257) );
  OR2_X1 U10478 ( .A1(n9710), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U10479 ( .A1(n9710), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9266) );
  NAND2_X1 U10480 ( .A1(n9267), .A2(n9266), .ZN(n9707) );
  NOR2_X1 U10481 ( .A1(n9706), .A2(n9707), .ZN(n9705) );
  AOI21_X1 U10482 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9710), .A(n9705), .ZN(
        n9268) );
  AOI22_X1 U10483 ( .A1(n9710), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9270), .B2(
        n9269), .ZN(n9717) );
  NAND2_X1 U10484 ( .A1(n9717), .A2(n9716), .ZN(n9715) );
  OAI21_X1 U10485 ( .B1(n9710), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9715), .ZN(
        n9273) );
  XNOR2_X1 U10486 ( .A(n9273), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9274) );
  AOI22_X1 U10487 ( .A1(n9276), .A2(n9709), .B1(n9719), .B2(n9274), .ZN(n9279)
         );
  INV_X1 U10488 ( .A(n9274), .ZN(n9277) );
  NAND2_X1 U10489 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3084), .ZN(n9280) );
  NAND2_X1 U10490 ( .A1(n9524), .A2(n9287), .ZN(n9520) );
  XNOR2_X1 U10491 ( .A(n9520), .B(n9517), .ZN(n9519) );
  NAND2_X1 U10492 ( .A1(n9283), .A2(n9282), .ZN(n9522) );
  NOR2_X1 U10493 ( .A1(n9735), .A2(n9522), .ZN(n9290) );
  AOI21_X1 U10494 ( .B1(n9735), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9290), .ZN(
        n9285) );
  NAND2_X1 U10495 ( .A1(n9517), .A2(n9462), .ZN(n9284) );
  OAI211_X1 U10496 ( .C1(n9519), .C2(n9286), .A(n9285), .B(n9284), .ZN(
        P1_U3261) );
  INV_X1 U10497 ( .A(n9287), .ZN(n9289) );
  NAND2_X1 U10498 ( .A1(n9289), .A2(n9288), .ZN(n9521) );
  NAND3_X1 U10499 ( .A1(n9521), .A2(n9494), .A3(n9520), .ZN(n9292) );
  AOI21_X1 U10500 ( .B1(n9735), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9290), .ZN(
        n9291) );
  OAI211_X1 U10501 ( .C1(n9524), .C2(n9502), .A(n9292), .B(n9291), .ZN(
        P1_U3262) );
  XOR2_X1 U10502 ( .A(n9296), .B(n9293), .Z(n9545) );
  OAI211_X1 U10503 ( .C1(n9294), .C2(n9296), .A(n9295), .B(n9509), .ZN(n9299)
         );
  AOI22_X1 U10504 ( .A1(n9297), .A2(n9510), .B1(n9506), .B2(n9334), .ZN(n9298)
         );
  AOI211_X1 U10505 ( .C1(n9543), .C2(n9307), .A(n9789), .B(n9300), .ZN(n9541)
         );
  NAND2_X1 U10506 ( .A1(n9541), .A2(n9514), .ZN(n9303) );
  AOI22_X1 U10507 ( .A1(n9301), .A2(n9499), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9735), .ZN(n9302) );
  OAI211_X1 U10508 ( .C1(n4938), .C2(n9502), .A(n9303), .B(n9302), .ZN(n9304)
         );
  AOI21_X1 U10509 ( .B1(n9542), .B2(n9733), .A(n9304), .ZN(n9305) );
  OAI21_X1 U10510 ( .B1(n9545), .B2(n9516), .A(n9305), .ZN(P1_U3264) );
  XOR2_X1 U10511 ( .A(n9306), .B(n9315), .Z(n9549) );
  INV_X1 U10512 ( .A(n9307), .ZN(n9308) );
  AOI21_X1 U10513 ( .B1(n4943), .B2(n4944), .A(n9308), .ZN(n9546) );
  AOI22_X1 U10514 ( .A1(n9309), .A2(n9499), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9735), .ZN(n9310) );
  OAI21_X1 U10515 ( .B1(n9311), .B2(n9502), .A(n9310), .ZN(n9322) );
  NAND2_X1 U10516 ( .A1(n9313), .A2(n9312), .ZN(n9314) );
  XOR2_X1 U10517 ( .A(n9315), .B(n9314), .Z(n9320) );
  AOI211_X1 U10518 ( .C1(n9494), .C2(n9546), .A(n9322), .B(n9321), .ZN(n9323)
         );
  OAI21_X1 U10519 ( .B1(n9516), .B2(n9549), .A(n9323), .ZN(P1_U3265) );
  XOR2_X1 U10520 ( .A(n9324), .B(n9333), .Z(n9554) );
  AOI21_X1 U10521 ( .B1(n9550), .B2(n9339), .A(n9325), .ZN(n9551) );
  INV_X1 U10522 ( .A(n9550), .ZN(n9329) );
  INV_X1 U10523 ( .A(n9326), .ZN(n9327) );
  AOI22_X1 U10524 ( .A1(n9327), .A2(n9499), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9735), .ZN(n9328) );
  OAI21_X1 U10525 ( .B1(n9329), .B2(n9502), .A(n9328), .ZN(n9336) );
  NAND2_X1 U10526 ( .A1(n9331), .A2(n9330), .ZN(n9332) );
  NOR2_X1 U10527 ( .A1(n9553), .A2(n9735), .ZN(n9335) );
  AOI211_X1 U10528 ( .C1(n9551), .C2(n9494), .A(n9336), .B(n9335), .ZN(n9337)
         );
  OAI21_X1 U10529 ( .B1(n9554), .B2(n9516), .A(n9337), .ZN(P1_U3266) );
  XNOR2_X1 U10530 ( .A(n9338), .B(n9346), .ZN(n9558) );
  INV_X1 U10531 ( .A(n9353), .ZN(n9341) );
  INV_X1 U10532 ( .A(n9339), .ZN(n9340) );
  AOI21_X1 U10533 ( .B1(n4942), .B2(n9341), .A(n9340), .ZN(n9555) );
  AOI22_X1 U10534 ( .A1(n9342), .A2(n9499), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9735), .ZN(n9343) );
  OAI21_X1 U10535 ( .B1(n9344), .B2(n9502), .A(n9343), .ZN(n9350) );
  XNOR2_X1 U10536 ( .A(n9345), .B(n9346), .ZN(n9347) );
  NOR2_X1 U10537 ( .A1(n9557), .A2(n9735), .ZN(n9349) );
  OAI21_X1 U10538 ( .B1(n9558), .B2(n9516), .A(n9351), .ZN(P1_U3267) );
  XNOR2_X1 U10539 ( .A(n9352), .B(n9360), .ZN(n9563) );
  AOI21_X1 U10540 ( .B1(n9559), .B2(n9367), .A(n9353), .ZN(n9560) );
  INV_X1 U10541 ( .A(n9559), .ZN(n9357) );
  INV_X1 U10542 ( .A(n9354), .ZN(n9355) );
  AOI22_X1 U10543 ( .A1(n9355), .A2(n9499), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9735), .ZN(n9356) );
  OAI21_X1 U10544 ( .B1(n9357), .B2(n9502), .A(n9356), .ZN(n9364) );
  NAND2_X1 U10545 ( .A1(n9374), .A2(n9358), .ZN(n9359) );
  XOR2_X1 U10546 ( .A(n9360), .B(n9359), .Z(n9361) );
  AOI222_X1 U10547 ( .A1(n9362), .A2(n9510), .B1(n9509), .B2(n9361), .C1(n9392), .C2(n9506), .ZN(n9562) );
  NOR2_X1 U10548 ( .A1(n9562), .A2(n9735), .ZN(n9363) );
  AOI211_X1 U10549 ( .C1(n9560), .C2(n9494), .A(n9364), .B(n9363), .ZN(n9365)
         );
  OAI21_X1 U10550 ( .B1(n9516), .B2(n9563), .A(n9365), .ZN(P1_U3268) );
  XOR2_X1 U10551 ( .A(n9366), .B(n9376), .Z(n9568) );
  INV_X1 U10552 ( .A(n9383), .ZN(n9369) );
  INV_X1 U10553 ( .A(n9367), .ZN(n9368) );
  AOI21_X1 U10554 ( .B1(n9564), .B2(n9369), .A(n9368), .ZN(n9565) );
  INV_X1 U10555 ( .A(n9370), .ZN(n9371) );
  AOI22_X1 U10556 ( .A1(n9371), .A2(n9499), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9735), .ZN(n9372) );
  OAI21_X1 U10557 ( .B1(n9373), .B2(n9502), .A(n9372), .ZN(n9380) );
  OAI21_X1 U10558 ( .B1(n9376), .B2(n9375), .A(n9374), .ZN(n9378) );
  AOI222_X1 U10559 ( .A1(n9378), .A2(n9509), .B1(n9408), .B2(n9506), .C1(n9377), .C2(n9510), .ZN(n9567) );
  NOR2_X1 U10560 ( .A1(n9567), .A2(n9735), .ZN(n9379) );
  AOI211_X1 U10561 ( .C1(n9565), .C2(n9494), .A(n9380), .B(n9379), .ZN(n9381)
         );
  OAI21_X1 U10562 ( .B1(n9516), .B2(n9568), .A(n9381), .ZN(P1_U3269) );
  OAI21_X1 U10563 ( .B1(n4318), .B2(n4907), .A(n9382), .ZN(n9573) );
  AOI211_X1 U10564 ( .C1(n9570), .C2(n9398), .A(n9789), .B(n9383), .ZN(n9569)
         );
  INV_X1 U10565 ( .A(n9570), .ZN(n9386) );
  AOI22_X1 U10566 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n9735), .B1(n9384), .B2(
        n9499), .ZN(n9385) );
  OAI21_X1 U10567 ( .B1(n9386), .B2(n9502), .A(n9385), .ZN(n9395) );
  AND2_X1 U10568 ( .A1(n9388), .A2(n9387), .ZN(n9391) );
  OAI21_X1 U10569 ( .B1(n9391), .B2(n9390), .A(n9389), .ZN(n9393) );
  AOI222_X1 U10570 ( .A1(n9393), .A2(n9509), .B1(n9420), .B2(n9506), .C1(n9392), .C2(n9510), .ZN(n9572) );
  NOR2_X1 U10571 ( .A1(n9572), .A2(n9735), .ZN(n9394) );
  AOI211_X1 U10572 ( .C1(n9569), .C2(n9514), .A(n9395), .B(n9394), .ZN(n9396)
         );
  OAI21_X1 U10573 ( .B1(n9516), .B2(n9573), .A(n9396), .ZN(P1_U3270) );
  XNOR2_X1 U10574 ( .A(n9397), .B(n9405), .ZN(n9578) );
  INV_X1 U10575 ( .A(n9413), .ZN(n9400) );
  INV_X1 U10576 ( .A(n9398), .ZN(n9399) );
  AOI21_X1 U10577 ( .B1(n9574), .B2(n9400), .A(n9399), .ZN(n9575) );
  INV_X1 U10578 ( .A(n9401), .ZN(n9402) );
  AOI22_X1 U10579 ( .A1(n9735), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9402), .B2(
        n9499), .ZN(n9403) );
  OAI21_X1 U10580 ( .B1(n9404), .B2(n9502), .A(n9403), .ZN(n9410) );
  XOR2_X1 U10581 ( .A(n9406), .B(n9405), .Z(n9407) );
  AOI222_X1 U10582 ( .A1(n9408), .A2(n9510), .B1(n9509), .B2(n9407), .C1(n9436), .C2(n9506), .ZN(n9577) );
  NOR2_X1 U10583 ( .A1(n9577), .A2(n9735), .ZN(n9409) );
  AOI211_X1 U10584 ( .C1(n9575), .C2(n9494), .A(n9410), .B(n9409), .ZN(n9411)
         );
  OAI21_X1 U10585 ( .B1(n9516), .B2(n9578), .A(n9411), .ZN(P1_U3271) );
  XOR2_X1 U10586 ( .A(n9412), .B(n9418), .Z(n9583) );
  AOI211_X1 U10587 ( .C1(n9580), .C2(n4356), .A(n9789), .B(n9413), .ZN(n9579)
         );
  INV_X1 U10588 ( .A(n9414), .ZN(n9415) );
  AOI22_X1 U10589 ( .A1(n9735), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9415), .B2(
        n9499), .ZN(n9416) );
  OAI21_X1 U10590 ( .B1(n4934), .B2(n9502), .A(n9416), .ZN(n9422) );
  XNOR2_X1 U10591 ( .A(n9417), .B(n9418), .ZN(n9419) );
  AOI222_X1 U10592 ( .A1(n9420), .A2(n9510), .B1(n9509), .B2(n9419), .C1(n9450), .C2(n9506), .ZN(n9582) );
  NOR2_X1 U10593 ( .A1(n9582), .A2(n9735), .ZN(n9421) );
  AOI211_X1 U10594 ( .C1(n9579), .C2(n9514), .A(n9422), .B(n9421), .ZN(n9423)
         );
  OAI21_X1 U10595 ( .B1(n9516), .B2(n9583), .A(n9423), .ZN(P1_U3272) );
  XNOR2_X1 U10596 ( .A(n9425), .B(n9434), .ZN(n9588) );
  INV_X1 U10597 ( .A(n9442), .ZN(n9427) );
  INV_X1 U10598 ( .A(n4356), .ZN(n9426) );
  AOI21_X1 U10599 ( .B1(n9584), .B2(n9427), .A(n9426), .ZN(n9585) );
  INV_X1 U10600 ( .A(n9428), .ZN(n9429) );
  AOI22_X1 U10601 ( .A1(n9735), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9429), .B2(
        n9499), .ZN(n9430) );
  OAI21_X1 U10602 ( .B1(n9431), .B2(n9502), .A(n9430), .ZN(n9439) );
  NAND2_X1 U10603 ( .A1(n9433), .A2(n9432), .ZN(n9435) );
  XNOR2_X1 U10604 ( .A(n9435), .B(n9434), .ZN(n9437) );
  AOI222_X1 U10605 ( .A1(n9437), .A2(n9509), .B1(n9457), .B2(n9506), .C1(n9436), .C2(n9510), .ZN(n9587) );
  NOR2_X1 U10606 ( .A1(n9587), .A2(n9735), .ZN(n9438) );
  AOI211_X1 U10607 ( .C1(n9585), .C2(n9494), .A(n9439), .B(n9438), .ZN(n9440)
         );
  OAI21_X1 U10608 ( .B1(n9516), .B2(n9588), .A(n9440), .ZN(P1_U3273) );
  XOR2_X1 U10609 ( .A(n9441), .B(n9447), .Z(n9593) );
  AOI21_X1 U10610 ( .B1(n9589), .B2(n4354), .A(n9442), .ZN(n9590) );
  INV_X1 U10611 ( .A(n9589), .ZN(n9445) );
  AOI22_X1 U10612 ( .A1(n9735), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9443), .B2(
        n9499), .ZN(n9444) );
  OAI21_X1 U10613 ( .B1(n9445), .B2(n9502), .A(n9444), .ZN(n9452) );
  XNOR2_X1 U10614 ( .A(n9446), .B(n9447), .ZN(n9449) );
  AOI222_X1 U10615 ( .A1(n9450), .A2(n9510), .B1(n9509), .B2(n9449), .C1(n9448), .C2(n9506), .ZN(n9592) );
  NOR2_X1 U10616 ( .A1(n9592), .A2(n9735), .ZN(n9451) );
  AOI211_X1 U10617 ( .C1(n9590), .C2(n9494), .A(n9452), .B(n9451), .ZN(n9453)
         );
  OAI21_X1 U10618 ( .B1(n9516), .B2(n9593), .A(n9453), .ZN(P1_U3274) );
  NAND2_X1 U10619 ( .A1(n9454), .A2(n9455), .ZN(n9456) );
  XNOR2_X1 U10620 ( .A(n9456), .B(n9467), .ZN(n9459) );
  AOI222_X1 U10621 ( .A1(n9459), .A2(n9509), .B1(n9458), .B2(n9506), .C1(n9457), .C2(n9510), .ZN(n9597) );
  AOI21_X1 U10622 ( .B1(n9460), .B2(n9595), .A(n9789), .ZN(n9461) );
  AND2_X1 U10623 ( .A1(n9461), .A2(n4354), .ZN(n9594) );
  NAND2_X1 U10624 ( .A1(n9595), .A2(n9462), .ZN(n9464) );
  NAND2_X1 U10625 ( .A1(n9735), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9463) );
  OAI211_X1 U10626 ( .C1(n9728), .C2(n9465), .A(n9464), .B(n9463), .ZN(n9470)
         );
  OAI21_X1 U10627 ( .B1(n9468), .B2(n9467), .A(n9466), .ZN(n9598) );
  NOR2_X1 U10628 ( .A1(n9598), .A2(n9516), .ZN(n9469) );
  AOI211_X1 U10629 ( .C1(n9594), .C2(n9471), .A(n9470), .B(n9469), .ZN(n9472)
         );
  OAI21_X1 U10630 ( .B1(n9735), .B2(n9597), .A(n9472), .ZN(P1_U3275) );
  XNOR2_X1 U10631 ( .A(n9473), .B(n9479), .ZN(n9483) );
  OAI22_X1 U10632 ( .A1(n9477), .A2(n9476), .B1(n9475), .B2(n9474), .ZN(n9482)
         );
  XNOR2_X1 U10633 ( .A(n9478), .B(n9479), .ZN(n9603) );
  NOR2_X1 U10634 ( .A1(n9603), .A2(n9480), .ZN(n9481) );
  AOI211_X1 U10635 ( .C1(n9509), .C2(n9483), .A(n9482), .B(n9481), .ZN(n9602)
         );
  INV_X1 U10636 ( .A(n9484), .ZN(n9486) );
  INV_X1 U10637 ( .A(n9460), .ZN(n9485) );
  AOI21_X1 U10638 ( .B1(n9599), .B2(n9486), .A(n9485), .ZN(n9600) );
  INV_X1 U10639 ( .A(n9487), .ZN(n9488) );
  AOI22_X1 U10640 ( .A1(n9735), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9488), .B2(
        n9499), .ZN(n9489) );
  OAI21_X1 U10641 ( .B1(n9490), .B2(n9502), .A(n9489), .ZN(n9493) );
  NOR2_X1 U10642 ( .A1(n9603), .A2(n9491), .ZN(n9492) );
  AOI211_X1 U10643 ( .C1(n9600), .C2(n9494), .A(n9493), .B(n9492), .ZN(n9495)
         );
  OAI21_X1 U10644 ( .B1(n9602), .B2(n9735), .A(n9495), .ZN(P1_U3276) );
  XOR2_X1 U10645 ( .A(n9504), .B(n9496), .Z(n9613) );
  INV_X1 U10646 ( .A(n9497), .ZN(n9498) );
  AOI211_X1 U10647 ( .C1(n9610), .C2(n8150), .A(n9789), .B(n9498), .ZN(n9609)
         );
  AOI22_X1 U10648 ( .A1(n9735), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9500), .B2(
        n9499), .ZN(n9501) );
  OAI21_X1 U10649 ( .B1(n4948), .B2(n9502), .A(n9501), .ZN(n9513) );
  XNOR2_X1 U10650 ( .A(n9505), .B(n9504), .ZN(n9508) );
  AOI222_X1 U10651 ( .A1(n9511), .A2(n9510), .B1(n9509), .B2(n9508), .C1(n9507), .C2(n9506), .ZN(n9612) );
  NOR2_X1 U10652 ( .A1(n9612), .A2(n9735), .ZN(n9512) );
  AOI211_X1 U10653 ( .C1(n9609), .C2(n9514), .A(n9513), .B(n9512), .ZN(n9515)
         );
  OAI21_X1 U10654 ( .B1(n9516), .B2(n9613), .A(n9515), .ZN(P1_U3278) );
  NAND2_X1 U10655 ( .A1(n9517), .A2(n9626), .ZN(n9518) );
  OAI211_X1 U10656 ( .C1(n9519), .C2(n9789), .A(n9518), .B(n9522), .ZN(n9634)
         );
  MUX2_X1 U10657 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9634), .S(n9801), .Z(
        P1_U3554) );
  NAND3_X1 U10658 ( .A1(n9521), .A2(n9627), .A3(n9520), .ZN(n9523) );
  OAI211_X1 U10659 ( .C1(n9524), .C2(n9787), .A(n9523), .B(n9522), .ZN(n9635)
         );
  MUX2_X1 U10660 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9635), .S(n9801), .Z(
        P1_U3553) );
  NOR3_X1 U10661 ( .A1(n9531), .A2(n9624), .A3(n9530), .ZN(n9526) );
  INV_X1 U10662 ( .A(n9624), .ZN(n9784) );
  NAND4_X1 U10663 ( .A1(n9534), .A2(n9531), .A3(n9784), .A4(n9530), .ZN(n9535)
         );
  NAND2_X1 U10664 ( .A1(n9532), .A2(n9784), .ZN(n9533) );
  MUX2_X1 U10665 ( .A(n9636), .B(P1_REG1_REG_29__SCAN_IN), .S(n9799), .Z(
        P1_U3552) );
  AOI22_X1 U10666 ( .A1(n9537), .A2(n9627), .B1(n9626), .B2(n9536), .ZN(n9538)
         );
  MUX2_X1 U10667 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9637), .S(n9801), .Z(
        P1_U3551) );
  OAI21_X1 U10668 ( .B1(n9545), .B2(n9624), .A(n9544), .ZN(n9638) );
  MUX2_X1 U10669 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9638), .S(n9801), .Z(
        P1_U3550) );
  AOI22_X1 U10670 ( .A1(n9546), .A2(n9627), .B1(n9626), .B2(n4943), .ZN(n9547)
         );
  OAI211_X1 U10671 ( .C1(n9549), .C2(n9624), .A(n9548), .B(n9547), .ZN(n9639)
         );
  MUX2_X1 U10672 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9639), .S(n9801), .Z(
        P1_U3549) );
  AOI22_X1 U10673 ( .A1(n9551), .A2(n9627), .B1(n9626), .B2(n9550), .ZN(n9552)
         );
  OAI211_X1 U10674 ( .C1(n9554), .C2(n9624), .A(n9553), .B(n9552), .ZN(n9640)
         );
  MUX2_X1 U10675 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9640), .S(n9801), .Z(
        P1_U3548) );
  AOI22_X1 U10676 ( .A1(n9555), .A2(n9627), .B1(n9626), .B2(n4942), .ZN(n9556)
         );
  OAI211_X1 U10677 ( .C1(n9558), .C2(n9624), .A(n9557), .B(n9556), .ZN(n9641)
         );
  MUX2_X1 U10678 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9641), .S(n9801), .Z(
        P1_U3547) );
  AOI22_X1 U10679 ( .A1(n9560), .A2(n9627), .B1(n9626), .B2(n9559), .ZN(n9561)
         );
  OAI211_X1 U10680 ( .C1(n9624), .C2(n9563), .A(n9562), .B(n9561), .ZN(n9642)
         );
  MUX2_X1 U10681 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9642), .S(n9801), .Z(
        P1_U3546) );
  AOI22_X1 U10682 ( .A1(n9565), .A2(n9627), .B1(n9626), .B2(n9564), .ZN(n9566)
         );
  OAI211_X1 U10683 ( .C1(n9568), .C2(n9624), .A(n9567), .B(n9566), .ZN(n9643)
         );
  MUX2_X1 U10684 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9643), .S(n9801), .Z(
        P1_U3545) );
  AOI21_X1 U10685 ( .B1(n9626), .B2(n9570), .A(n9569), .ZN(n9571) );
  OAI211_X1 U10686 ( .C1(n9573), .C2(n9624), .A(n9572), .B(n9571), .ZN(n9644)
         );
  MUX2_X1 U10687 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9644), .S(n9801), .Z(
        P1_U3544) );
  AOI22_X1 U10688 ( .A1(n9575), .A2(n9627), .B1(n9626), .B2(n9574), .ZN(n9576)
         );
  OAI211_X1 U10689 ( .C1(n9624), .C2(n9578), .A(n9577), .B(n9576), .ZN(n9645)
         );
  MUX2_X1 U10690 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9645), .S(n9801), .Z(
        P1_U3543) );
  AOI21_X1 U10691 ( .B1(n9626), .B2(n9580), .A(n9579), .ZN(n9581) );
  OAI211_X1 U10692 ( .C1(n9583), .C2(n9624), .A(n9582), .B(n9581), .ZN(n9646)
         );
  MUX2_X1 U10693 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9646), .S(n9801), .Z(
        P1_U3542) );
  AOI22_X1 U10694 ( .A1(n9585), .A2(n9627), .B1(n9626), .B2(n9584), .ZN(n9586)
         );
  OAI211_X1 U10695 ( .C1(n9588), .C2(n9624), .A(n9587), .B(n9586), .ZN(n9647)
         );
  MUX2_X1 U10696 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9647), .S(n9801), .Z(
        P1_U3541) );
  AOI22_X1 U10697 ( .A1(n9590), .A2(n9627), .B1(n9626), .B2(n9589), .ZN(n9591)
         );
  OAI211_X1 U10698 ( .C1(n9593), .C2(n9624), .A(n9592), .B(n9591), .ZN(n9648)
         );
  MUX2_X1 U10699 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9648), .S(n9801), .Z(
        P1_U3540) );
  AOI21_X1 U10700 ( .B1(n9626), .B2(n9595), .A(n9594), .ZN(n9596) );
  OAI211_X1 U10701 ( .C1(n9624), .C2(n9598), .A(n9597), .B(n9596), .ZN(n9649)
         );
  MUX2_X1 U10702 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9649), .S(n9801), .Z(
        P1_U3539) );
  AOI22_X1 U10703 ( .A1(n9600), .A2(n9627), .B1(n9626), .B2(n9599), .ZN(n9601)
         );
  OAI211_X1 U10704 ( .C1(n9632), .C2(n9603), .A(n9602), .B(n9601), .ZN(n9650)
         );
  MUX2_X1 U10705 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9650), .S(n9801), .Z(
        P1_U3538) );
  AOI211_X1 U10706 ( .C1(n9626), .C2(n9606), .A(n9605), .B(n9604), .ZN(n9607)
         );
  OAI21_X1 U10707 ( .B1(n9624), .B2(n9608), .A(n9607), .ZN(n9651) );
  MUX2_X1 U10708 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9651), .S(n9801), .Z(
        P1_U3537) );
  AOI21_X1 U10709 ( .B1(n9626), .B2(n9610), .A(n9609), .ZN(n9611) );
  OAI211_X1 U10710 ( .C1(n9624), .C2(n9613), .A(n9612), .B(n9611), .ZN(n9652)
         );
  MUX2_X1 U10711 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9652), .S(n9801), .Z(
        P1_U3536) );
  AOI21_X1 U10712 ( .B1(n9626), .B2(n9615), .A(n9614), .ZN(n9616) );
  OAI211_X1 U10713 ( .C1(n9632), .C2(n9618), .A(n9617), .B(n9616), .ZN(n9653)
         );
  MUX2_X1 U10714 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9653), .S(n9801), .Z(
        P1_U3535) );
  AOI21_X1 U10715 ( .B1(n9626), .B2(n9620), .A(n9619), .ZN(n9621) );
  OAI211_X1 U10716 ( .C1(n9624), .C2(n9623), .A(n9622), .B(n9621), .ZN(n9654)
         );
  MUX2_X1 U10717 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n9654), .S(n9801), .Z(
        P1_U3533) );
  AOI22_X1 U10718 ( .A1(n9628), .A2(n9627), .B1(n9626), .B2(n9625), .ZN(n9629)
         );
  OAI211_X1 U10719 ( .C1(n9632), .C2(n9631), .A(n9630), .B(n9629), .ZN(n9656)
         );
  MUX2_X1 U10720 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9656), .S(n9801), .Z(
        P1_U3532) );
  MUX2_X1 U10721 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9633), .S(n9801), .Z(
        P1_U3523) );
  MUX2_X1 U10722 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9634), .S(n9796), .Z(
        P1_U3522) );
  MUX2_X1 U10723 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9635), .S(n9796), .Z(
        P1_U3521) );
  MUX2_X1 U10724 ( .A(n9636), .B(P1_REG0_REG_29__SCAN_IN), .S(n9795), .Z(
        P1_U3520) );
  MUX2_X1 U10725 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9638), .S(n9796), .Z(
        P1_U3518) );
  MUX2_X1 U10726 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9639), .S(n9796), .Z(
        P1_U3517) );
  MUX2_X1 U10727 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9640), .S(n9796), .Z(
        P1_U3516) );
  MUX2_X1 U10728 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9641), .S(n9796), .Z(
        P1_U3515) );
  MUX2_X1 U10729 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9642), .S(n9796), .Z(
        P1_U3514) );
  MUX2_X1 U10730 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9643), .S(n9796), .Z(
        P1_U3513) );
  MUX2_X1 U10731 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9644), .S(n9796), .Z(
        P1_U3512) );
  MUX2_X1 U10732 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9645), .S(n9796), .Z(
        P1_U3511) );
  MUX2_X1 U10733 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9646), .S(n9796), .Z(
        P1_U3510) );
  MUX2_X1 U10734 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9647), .S(n9796), .Z(
        P1_U3508) );
  MUX2_X1 U10735 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9648), .S(n9796), .Z(
        P1_U3505) );
  MUX2_X1 U10736 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9649), .S(n9796), .Z(
        P1_U3502) );
  MUX2_X1 U10737 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9650), .S(n9796), .Z(
        P1_U3499) );
  MUX2_X1 U10738 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9651), .S(n9655), .Z(
        P1_U3496) );
  MUX2_X1 U10739 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9652), .S(n9655), .Z(
        P1_U3493) );
  MUX2_X1 U10740 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9653), .S(n9655), .Z(
        P1_U3490) );
  MUX2_X1 U10741 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n9654), .S(n9655), .Z(
        P1_U3484) );
  MUX2_X1 U10742 ( .A(P1_REG0_REG_9__SCAN_IN), .B(n9656), .S(n9655), .Z(
        P1_U3481) );
  MUX2_X1 U10743 ( .A(n9657), .B(P1_D_REG_0__SCAN_IN), .S(n9738), .Z(P1_U3440)
         );
  NOR4_X1 U10744 ( .A1(n5980), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9659), .A4(
        P1_U3084), .ZN(n9660) );
  AOI21_X1 U10745 ( .B1(n10113), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9660), 
        .ZN(n9661) );
  OAI21_X1 U10746 ( .B1(n9662), .B2(n10109), .A(n9661), .ZN(P1_U3322) );
  AOI22_X1 U10747 ( .A1(n9663), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10113), .ZN(n9664) );
  OAI21_X1 U10748 ( .B1(n9665), .B2(n10109), .A(n9664), .ZN(P1_U3323) );
  AOI22_X1 U10749 ( .A1(n9666), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10113), .ZN(n9667) );
  OAI21_X1 U10750 ( .B1(n9668), .B2(n10109), .A(n9667), .ZN(P1_U3324) );
  AOI22_X1 U10751 ( .A1(n9669), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10113), .ZN(n9670) );
  OAI21_X1 U10752 ( .B1(n9671), .B2(n10109), .A(n9670), .ZN(P1_U3325) );
  AOI22_X1 U10753 ( .A1(n9672), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n10113), .ZN(n9673) );
  OAI21_X1 U10754 ( .B1(n9674), .B2(n10109), .A(n9673), .ZN(P1_U3326) );
  AOI22_X1 U10755 ( .A1(n9675), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10113), .ZN(n9676) );
  OAI21_X1 U10756 ( .B1(n9677), .B2(n10109), .A(n9676), .ZN(P1_U3327) );
  MUX2_X1 U10757 ( .A(n9678), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10758 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10122) );
  NOR2_X1 U10759 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9679) );
  AOI21_X1 U10760 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9679), .ZN(n9933) );
  NOR2_X1 U10761 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(P2_ADDR_REG_16__SCAN_IN), 
        .ZN(n9680) );
  AOI21_X1 U10762 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9680), .ZN(n9936) );
  NOR2_X1 U10763 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9681) );
  AOI21_X1 U10764 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9681), .ZN(n9939) );
  NAND2_X1 U10765 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9682) );
  OAI21_X1 U10766 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9682), .ZN(n9945) );
  NAND2_X1 U10767 ( .A1(n9990), .A2(n9987), .ZN(n9967) );
  AOI22_X1 U10768 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n7399), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n10089), .ZN(n10136) );
  NAND2_X1 U10769 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9687) );
  XOR2_X1 U10770 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10134) );
  NAND2_X1 U10771 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9685) );
  XOR2_X1 U10772 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10132) );
  AOI21_X1 U10773 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9927) );
  INV_X1 U10774 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9683) );
  NAND3_X1 U10775 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9929) );
  NAND2_X1 U10776 ( .A1(n10132), .A2(n10131), .ZN(n9684) );
  NAND2_X1 U10777 ( .A1(n9685), .A2(n9684), .ZN(n10133) );
  NAND2_X1 U10778 ( .A1(n10134), .A2(n10133), .ZN(n9686) );
  NAND2_X1 U10779 ( .A1(n9687), .A2(n9686), .ZN(n10135) );
  NOR2_X1 U10780 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9688), .ZN(n10118) );
  NAND2_X1 U10781 ( .A1(n9690), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9691) );
  NAND2_X1 U10782 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9692), .ZN(n9693) );
  XOR2_X1 U10783 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9692), .Z(n10130) );
  INV_X1 U10784 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10129) );
  XNOR2_X1 U10785 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9694), .ZN(n10128) );
  INV_X1 U10786 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10019) );
  NOR2_X1 U10787 ( .A1(n9696), .A2(n10019), .ZN(n9697) );
  XNOR2_X1 U10788 ( .A(n10019), .B(n9696), .ZN(n10125) );
  NAND2_X1 U10789 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9698) );
  OAI21_X1 U10790 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9698), .ZN(n9954) );
  NAND2_X1 U10791 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9699) );
  OAI21_X1 U10792 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9699), .ZN(n9951) );
  NAND2_X1 U10793 ( .A1(n9967), .A2(n9947), .ZN(n9944) );
  NOR2_X1 U10794 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9700) );
  AOI21_X1 U10795 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9700), .ZN(n9941) );
  NAND2_X1 U10796 ( .A1(n9942), .A2(n9941), .ZN(n9940) );
  NAND2_X1 U10797 ( .A1(n9939), .A2(n9938), .ZN(n9937) );
  NAND2_X1 U10798 ( .A1(n9933), .A2(n9932), .ZN(n9931) );
  NOR2_X1 U10799 ( .A1(n10122), .A2(n10121), .ZN(n9701) );
  NAND2_X1 U10800 ( .A1(n10122), .A2(n10121), .ZN(n10120) );
  XNOR2_X1 U10801 ( .A(n9702), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n9703) );
  XNOR2_X1 U10802 ( .A(n9704), .B(n9703), .ZN(ADD_1071_U4) );
  INV_X1 U10803 ( .A(P1_WR_REG_SCAN_IN), .ZN(n10070) );
  INV_X1 U10804 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10020) );
  AOI22_X1 U10805 ( .A1(P2_WR_REG_SCAN_IN), .A2(n10070), .B1(P1_WR_REG_SCAN_IN), .B2(n10020), .ZN(U123) );
  XNOR2_X1 U10806 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U10807 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9708) );
  NAND2_X1 U10808 ( .A1(n9709), .A2(n9708), .ZN(n9714) );
  NAND2_X1 U10809 ( .A1(n9711), .A2(n9710), .ZN(n9713) );
  AND3_X1 U10810 ( .A1(n9714), .A2(n9713), .A3(n9712), .ZN(n9722) );
  OAI21_X1 U10811 ( .B1(n9717), .B2(n9716), .A(n9715), .ZN(n9720) );
  AOI22_X1 U10812 ( .A1(n9720), .A2(n9719), .B1(n9718), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U10813 ( .A1(n9722), .A2(n9721), .ZN(P1_U3259) );
  INV_X1 U10814 ( .A(n9723), .ZN(n9726) );
  AOI22_X1 U10815 ( .A1(n9726), .A2(n6576), .B1(n9725), .B2(n9724), .ZN(n9727)
         );
  OAI21_X1 U10816 ( .B1(n6065), .B2(n9728), .A(n9727), .ZN(n9729) );
  AOI211_X1 U10817 ( .C1(n9732), .C2(n9731), .A(n9730), .B(n9729), .ZN(n9734)
         );
  AOI22_X1 U10818 ( .A1(n9735), .A2(n6883), .B1(n9734), .B2(n9733), .ZN(
        P1_U3290) );
  INV_X1 U10819 ( .A(n9736), .ZN(n9737) );
  INV_X1 U10820 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10094) );
  NOR2_X1 U10821 ( .A1(n9754), .A2(n10094), .ZN(P1_U3292) );
  INV_X1 U10822 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9739) );
  NOR2_X1 U10823 ( .A1(n9754), .A2(n9739), .ZN(P1_U3293) );
  INV_X1 U10824 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9740) );
  NOR2_X1 U10825 ( .A1(n9754), .A2(n9740), .ZN(P1_U3294) );
  INV_X1 U10826 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9741) );
  NOR2_X1 U10827 ( .A1(n9754), .A2(n9741), .ZN(P1_U3295) );
  INV_X1 U10828 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9742) );
  NOR2_X1 U10829 ( .A1(n9754), .A2(n9742), .ZN(P1_U3296) );
  INV_X1 U10830 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9743) );
  NOR2_X1 U10831 ( .A1(n9754), .A2(n9743), .ZN(P1_U3297) );
  INV_X1 U10832 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U10833 ( .A1(n9754), .A2(n10047), .ZN(P1_U3298) );
  INV_X1 U10834 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9744) );
  NOR2_X1 U10835 ( .A1(n9754), .A2(n9744), .ZN(P1_U3299) );
  INV_X1 U10836 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9745) );
  NOR2_X1 U10837 ( .A1(n9754), .A2(n9745), .ZN(P1_U3300) );
  INV_X1 U10838 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9746) );
  NOR2_X1 U10839 ( .A1(n9754), .A2(n9746), .ZN(P1_U3301) );
  INV_X1 U10840 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9747) );
  NOR2_X1 U10841 ( .A1(n9754), .A2(n9747), .ZN(P1_U3302) );
  INV_X1 U10842 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10052) );
  NOR2_X1 U10843 ( .A1(n9754), .A2(n10052), .ZN(P1_U3303) );
  INV_X1 U10844 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9748) );
  NOR2_X1 U10845 ( .A1(n9754), .A2(n9748), .ZN(P1_U3304) );
  INV_X1 U10846 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U10847 ( .A1(n9754), .A2(n10063), .ZN(P1_U3305) );
  INV_X1 U10848 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9749) );
  NOR2_X1 U10849 ( .A1(n9754), .A2(n9749), .ZN(P1_U3306) );
  INV_X1 U10850 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9750) );
  NOR2_X1 U10851 ( .A1(n9754), .A2(n9750), .ZN(P1_U3307) );
  INV_X1 U10852 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9751) );
  NOR2_X1 U10853 ( .A1(n9754), .A2(n9751), .ZN(P1_U3308) );
  INV_X1 U10854 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9752) );
  NOR2_X1 U10855 ( .A1(n9754), .A2(n9752), .ZN(P1_U3309) );
  INV_X1 U10856 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9753) );
  NOR2_X1 U10857 ( .A1(n9754), .A2(n9753), .ZN(P1_U3310) );
  INV_X1 U10858 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9755) );
  NOR2_X1 U10859 ( .A1(n9766), .A2(n9755), .ZN(P1_U3311) );
  INV_X1 U10860 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9756) );
  NOR2_X1 U10861 ( .A1(n9766), .A2(n9756), .ZN(P1_U3312) );
  INV_X1 U10862 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9757) );
  NOR2_X1 U10863 ( .A1(n9766), .A2(n9757), .ZN(P1_U3313) );
  INV_X1 U10864 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9758) );
  NOR2_X1 U10865 ( .A1(n9766), .A2(n9758), .ZN(P1_U3314) );
  INV_X1 U10866 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9759) );
  NOR2_X1 U10867 ( .A1(n9766), .A2(n9759), .ZN(P1_U3315) );
  INV_X1 U10868 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n9760) );
  NOR2_X1 U10869 ( .A1(n9766), .A2(n9760), .ZN(P1_U3316) );
  INV_X1 U10870 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9761) );
  NOR2_X1 U10871 ( .A1(n9766), .A2(n9761), .ZN(P1_U3317) );
  INV_X1 U10872 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9762) );
  NOR2_X1 U10873 ( .A1(n9766), .A2(n9762), .ZN(P1_U3318) );
  INV_X1 U10874 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9763) );
  NOR2_X1 U10875 ( .A1(n9766), .A2(n9763), .ZN(P1_U3319) );
  INV_X1 U10876 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9764) );
  NOR2_X1 U10877 ( .A1(n9766), .A2(n9764), .ZN(P1_U3320) );
  INV_X1 U10878 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9765) );
  NOR2_X1 U10879 ( .A1(n9766), .A2(n9765), .ZN(P1_U3321) );
  INV_X1 U10880 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9770) );
  NAND2_X1 U10881 ( .A1(n9767), .A2(n9769), .ZN(n9768) );
  OAI21_X1 U10882 ( .B1(n9770), .B2(n9769), .A(n9768), .ZN(P1_U3441) );
  INV_X1 U10883 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9771) );
  AOI22_X1 U10884 ( .A1(n9796), .A2(n9772), .B1(n9771), .B2(n9795), .ZN(
        P1_U3460) );
  INV_X1 U10885 ( .A(n9773), .ZN(n9774) );
  OAI22_X1 U10886 ( .A1(n9774), .A2(n9789), .B1(n4931), .B2(n9787), .ZN(n9776)
         );
  AOI211_X1 U10887 ( .C1(n9794), .C2(n9777), .A(n9776), .B(n9775), .ZN(n9797)
         );
  INV_X1 U10888 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U10889 ( .A1(n9796), .A2(n9797), .B1(n9778), .B2(n9795), .ZN(
        P1_U3466) );
  INV_X1 U10890 ( .A(n9779), .ZN(n9785) );
  OAI21_X1 U10891 ( .B1(n9781), .B2(n9787), .A(n9780), .ZN(n9783) );
  AOI211_X1 U10892 ( .C1(n9785), .C2(n9784), .A(n9783), .B(n9782), .ZN(n9798)
         );
  INV_X1 U10893 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9786) );
  AOI22_X1 U10894 ( .A1(n9796), .A2(n9798), .B1(n9786), .B2(n9795), .ZN(
        P1_U3469) );
  OAI22_X1 U10895 ( .A1(n9790), .A2(n9789), .B1(n9788), .B2(n9787), .ZN(n9792)
         );
  AOI211_X1 U10896 ( .C1(n9794), .C2(n9793), .A(n9792), .B(n9791), .ZN(n9800)
         );
  INV_X1 U10897 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10083) );
  AOI22_X1 U10898 ( .A1(n9796), .A2(n9800), .B1(n10083), .B2(n9795), .ZN(
        P1_U3472) );
  AOI22_X1 U10899 ( .A1(n9801), .A2(n9797), .B1(n6911), .B2(n9799), .ZN(
        P1_U3527) );
  AOI22_X1 U10900 ( .A1(n9801), .A2(n9798), .B1(n6914), .B2(n9799), .ZN(
        P1_U3528) );
  AOI22_X1 U10901 ( .A1(n9801), .A2(n9800), .B1(n9984), .B2(n9799), .ZN(
        P1_U3529) );
  OAI22_X1 U10902 ( .A1(n9827), .A2(n9803), .B1(n9807), .B2(n9802), .ZN(n9804)
         );
  INV_X1 U10903 ( .A(n9804), .ZN(n9812) );
  INV_X1 U10904 ( .A(n9813), .ZN(n10002) );
  OR2_X1 U10905 ( .A1(n9827), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9806) );
  OAI211_X1 U10906 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n9807), .A(n9806), .B(
        n9805), .ZN(n9808) );
  INV_X1 U10907 ( .A(n9808), .ZN(n9811) );
  AOI21_X1 U10908 ( .B1(n9817), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n9809), .ZN(
        n9810) );
  OAI221_X1 U10909 ( .B1(n9813), .B2(n9812), .C1(n10002), .C2(n9811), .A(n9810), .ZN(P2_U3245) );
  AOI21_X1 U10910 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n9815), .A(n9814), .ZN(
        n9828) );
  AOI21_X1 U10911 ( .B1(n9817), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n9816), .ZN(
        n9826) );
  OAI21_X1 U10912 ( .B1(n9820), .B2(n9819), .A(n9818), .ZN(n9824) );
  AOI22_X1 U10913 ( .A1(n9824), .A2(n9823), .B1(n9822), .B2(n9821), .ZN(n9825)
         );
  OAI211_X1 U10914 ( .C1(n9828), .C2(n9827), .A(n9826), .B(n9825), .ZN(
        P2_U3263) );
  AND2_X1 U10915 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9834), .ZN(P2_U3297) );
  AND2_X1 U10916 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9834), .ZN(P2_U3298) );
  AND2_X1 U10917 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9834), .ZN(P2_U3299) );
  AND2_X1 U10918 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9834), .ZN(P2_U3300) );
  AND2_X1 U10919 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9834), .ZN(P2_U3301) );
  AND2_X1 U10920 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9834), .ZN(P2_U3302) );
  INV_X1 U10921 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10029) );
  NOR2_X1 U10922 ( .A1(n9831), .A2(n10029), .ZN(P2_U3303) );
  INV_X1 U10923 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10068) );
  NOR2_X1 U10924 ( .A1(n9831), .A2(n10068), .ZN(P2_U3304) );
  INV_X1 U10925 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10061) );
  NOR2_X1 U10926 ( .A1(n9831), .A2(n10061), .ZN(P2_U3305) );
  AND2_X1 U10927 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9834), .ZN(P2_U3306) );
  AND2_X1 U10928 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9834), .ZN(P2_U3307) );
  AND2_X1 U10929 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9834), .ZN(P2_U3308) );
  AND2_X1 U10930 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9834), .ZN(P2_U3309) );
  AND2_X1 U10931 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9834), .ZN(P2_U3310) );
  INV_X1 U10932 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10013) );
  NOR2_X1 U10933 ( .A1(n9831), .A2(n10013), .ZN(P2_U3311) );
  AND2_X1 U10934 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9834), .ZN(P2_U3312) );
  AND2_X1 U10935 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9834), .ZN(P2_U3313) );
  AND2_X1 U10936 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9834), .ZN(P2_U3314) );
  AND2_X1 U10937 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n9834), .ZN(P2_U3315) );
  AND2_X1 U10938 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9834), .ZN(P2_U3316) );
  AND2_X1 U10939 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9834), .ZN(P2_U3317) );
  AND2_X1 U10940 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9834), .ZN(P2_U3318) );
  AND2_X1 U10941 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9834), .ZN(P2_U3319) );
  AND2_X1 U10942 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9834), .ZN(P2_U3320) );
  AND2_X1 U10943 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9834), .ZN(P2_U3321) );
  AND2_X1 U10944 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9834), .ZN(P2_U3322) );
  AND2_X1 U10945 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9834), .ZN(P2_U3323) );
  AND2_X1 U10946 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9834), .ZN(P2_U3324) );
  AND2_X1 U10947 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9834), .ZN(P2_U3325) );
  AND2_X1 U10948 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n9834), .ZN(P2_U3326) );
  AOI22_X1 U10949 ( .A1(n9837), .A2(n9833), .B1(n9832), .B2(n9834), .ZN(
        P2_U3437) );
  AOI22_X1 U10950 ( .A1(n9837), .A2(n9836), .B1(n9835), .B2(n9834), .ZN(
        P2_U3438) );
  AOI22_X1 U10951 ( .A1(n9840), .A2(n9902), .B1(n9839), .B2(n9838), .ZN(n9841)
         );
  AND2_X1 U10952 ( .A1(n9842), .A2(n9841), .ZN(n9914) );
  INV_X1 U10953 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9843) );
  AOI22_X1 U10954 ( .A1(n9913), .A2(n9914), .B1(n9843), .B2(n9912), .ZN(
        P2_U3451) );
  INV_X1 U10955 ( .A(n9844), .ZN(n9852) );
  NAND3_X1 U10956 ( .A1(n9847), .A2(n9846), .A3(n9845), .ZN(n9848) );
  OAI21_X1 U10957 ( .B1(n7199), .B2(n9905), .A(n9848), .ZN(n9851) );
  INV_X1 U10958 ( .A(n9849), .ZN(n9850) );
  AOI211_X1 U10959 ( .C1(n9902), .C2(n9852), .A(n9851), .B(n9850), .ZN(n9915)
         );
  AOI22_X1 U10960 ( .A1(n9913), .A2(n9915), .B1(n4988), .B2(n9912), .ZN(
        P2_U3454) );
  OAI22_X1 U10961 ( .A1(n9854), .A2(n9907), .B1(n9853), .B2(n9905), .ZN(n9857)
         );
  INV_X1 U10962 ( .A(n9855), .ZN(n9856) );
  AOI211_X1 U10963 ( .C1(n9902), .C2(n9858), .A(n9857), .B(n9856), .ZN(n9916)
         );
  INV_X1 U10964 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9859) );
  AOI22_X1 U10965 ( .A1(n9913), .A2(n9916), .B1(n9859), .B2(n9912), .ZN(
        P2_U3457) );
  INV_X1 U10966 ( .A(n9860), .ZN(n9892) );
  OAI22_X1 U10967 ( .A1(n9862), .A2(n9907), .B1(n9861), .B2(n9905), .ZN(n9863)
         );
  AOI21_X1 U10968 ( .B1(n9864), .B2(n9892), .A(n9863), .ZN(n9866) );
  AND2_X1 U10969 ( .A1(n9866), .A2(n9865), .ZN(n9917) );
  INV_X1 U10970 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9867) );
  AOI22_X1 U10971 ( .A1(n9913), .A2(n9917), .B1(n9867), .B2(n9912), .ZN(
        P2_U3460) );
  OAI22_X1 U10972 ( .A1(n9869), .A2(n9907), .B1(n9868), .B2(n9905), .ZN(n9871)
         );
  AOI211_X1 U10973 ( .C1(n9902), .C2(n9872), .A(n9871), .B(n9870), .ZN(n9918)
         );
  INV_X1 U10974 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9873) );
  AOI22_X1 U10975 ( .A1(n9913), .A2(n9918), .B1(n9873), .B2(n9912), .ZN(
        P2_U3463) );
  OAI22_X1 U10976 ( .A1(n9875), .A2(n9907), .B1(n9874), .B2(n9905), .ZN(n9878)
         );
  INV_X1 U10977 ( .A(n9876), .ZN(n9877) );
  AOI211_X1 U10978 ( .C1(n9902), .C2(n9879), .A(n9878), .B(n9877), .ZN(n9919)
         );
  INV_X1 U10979 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9880) );
  AOI22_X1 U10980 ( .A1(n9913), .A2(n9919), .B1(n9880), .B2(n9912), .ZN(
        P2_U3469) );
  OAI22_X1 U10981 ( .A1(n9881), .A2(n9907), .B1(n4846), .B2(n9905), .ZN(n9883)
         );
  AOI211_X1 U10982 ( .C1(n9902), .C2(n9884), .A(n9883), .B(n9882), .ZN(n9920)
         );
  INV_X1 U10983 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9885) );
  AOI22_X1 U10984 ( .A1(n9913), .A2(n9920), .B1(n9885), .B2(n9912), .ZN(
        P2_U3472) );
  OAI22_X1 U10985 ( .A1(n9887), .A2(n9907), .B1(n9886), .B2(n9905), .ZN(n9889)
         );
  AOI211_X1 U10986 ( .C1(n9892), .C2(n9890), .A(n9889), .B(n9888), .ZN(n9921)
         );
  INV_X1 U10987 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9891) );
  AOI22_X1 U10988 ( .A1(n9913), .A2(n9921), .B1(n9891), .B2(n9912), .ZN(
        P2_U3475) );
  NAND2_X1 U10989 ( .A1(n9893), .A2(n9892), .ZN(n9898) );
  OAI22_X1 U10990 ( .A1(n9895), .A2(n9907), .B1(n9894), .B2(n9905), .ZN(n9896)
         );
  INV_X1 U10991 ( .A(n9896), .ZN(n9897) );
  NAND2_X1 U10992 ( .A1(n9898), .A2(n9897), .ZN(n9899) );
  NOR2_X1 U10993 ( .A1(n9900), .A2(n9899), .ZN(n9922) );
  INV_X1 U10994 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9901) );
  AOI22_X1 U10995 ( .A1(n9913), .A2(n9922), .B1(n9901), .B2(n9912), .ZN(
        P2_U3478) );
  AND3_X1 U10996 ( .A1(n9904), .A2(n9903), .A3(n9902), .ZN(n9910) );
  OAI22_X1 U10997 ( .A1(n9908), .A2(n9907), .B1(n9906), .B2(n9905), .ZN(n9909)
         );
  NOR3_X1 U10998 ( .A1(n9911), .A2(n9910), .A3(n9909), .ZN(n9925) );
  AOI22_X1 U10999 ( .A1(n9913), .A2(n9925), .B1(n5197), .B2(n9912), .ZN(
        P2_U3481) );
  AOI22_X1 U11000 ( .A1(n9926), .A2(n9914), .B1(n9802), .B2(n9923), .ZN(
        P2_U3520) );
  AOI22_X1 U11001 ( .A1(n9926), .A2(n9915), .B1(n4986), .B2(n9923), .ZN(
        P2_U3521) );
  AOI22_X1 U11002 ( .A1(n9926), .A2(n9916), .B1(n5020), .B2(n9923), .ZN(
        P2_U3522) );
  AOI22_X1 U11003 ( .A1(n9926), .A2(n9917), .B1(n5042), .B2(n9923), .ZN(
        P2_U3523) );
  AOI22_X1 U11004 ( .A1(n9926), .A2(n9918), .B1(n5063), .B2(n9923), .ZN(
        P2_U3524) );
  AOI22_X1 U11005 ( .A1(n9926), .A2(n9919), .B1(n7045), .B2(n9923), .ZN(
        P2_U3526) );
  AOI22_X1 U11006 ( .A1(n9926), .A2(n9920), .B1(n5129), .B2(n9923), .ZN(
        P2_U3527) );
  AOI22_X1 U11007 ( .A1(n9926), .A2(n9921), .B1(n5156), .B2(n9923), .ZN(
        P2_U3528) );
  AOI22_X1 U11008 ( .A1(n9926), .A2(n9922), .B1(n5173), .B2(n9923), .ZN(
        P2_U3529) );
  AOI22_X1 U11009 ( .A1(n9926), .A2(n9925), .B1(n9924), .B2(n9923), .ZN(
        P2_U3530) );
  INV_X1 U11010 ( .A(n9927), .ZN(n9928) );
  NAND2_X1 U11011 ( .A1(n9929), .A2(n9928), .ZN(n9930) );
  XNOR2_X1 U11012 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9930), .ZN(ADD_1071_U5) );
  XOR2_X1 U11013 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11014 ( .B1(n9933), .B2(n9932), .A(n9931), .ZN(ADD_1071_U56) );
  OAI21_X1 U11015 ( .B1(n9936), .B2(n9935), .A(n9934), .ZN(ADD_1071_U57) );
  OAI21_X1 U11016 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(ADD_1071_U58) );
  OAI21_X1 U11017 ( .B1(n9942), .B2(n9941), .A(n9940), .ZN(ADD_1071_U59) );
  AOI21_X1 U11018 ( .B1(n9945), .B2(n9944), .A(n9943), .ZN(ADD_1071_U60) );
  OAI21_X1 U11019 ( .B1(n9987), .B2(n9990), .A(n9967), .ZN(n9946) );
  INV_X1 U11020 ( .A(n9946), .ZN(n9949) );
  OAI21_X1 U11021 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(ADD_1071_U61) );
  AOI21_X1 U11022 ( .B1(n9952), .B2(n9951), .A(n9950), .ZN(ADD_1071_U62) );
  AOI21_X1 U11023 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(ADD_1071_U63) );
  INV_X1 U11024 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10077) );
  NAND4_X1 U11025 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(P2_DATAO_REG_8__SCAN_IN), 
        .A3(n10077), .A4(n9956), .ZN(n9957) );
  NOR2_X1 U11026 ( .A1(n9958), .A2(n9957), .ZN(n9959) );
  NAND4_X1 U11027 ( .A1(n9959), .A2(P1_REG0_REG_7__SCAN_IN), .A3(
        P1_REG0_REG_6__SCAN_IN), .A4(n10090), .ZN(n9964) );
  NAND4_X1 U11028 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_REG1_REG_26__SCAN_IN), .A4(n6024), .ZN(n9963) );
  INV_X1 U11029 ( .A(SI_7_), .ZN(n9961) );
  INV_X1 U11030 ( .A(SI_0_), .ZN(n9960) );
  NAND4_X1 U11031 ( .A1(n9961), .A2(n9960), .A3(P2_DATAO_REG_0__SCAN_IN), .A4(
        P2_REG3_REG_6__SCAN_IN), .ZN(n9962) );
  NOR3_X1 U11032 ( .A1(n9964), .A2(n9963), .A3(n9962), .ZN(n10108) );
  NAND2_X1 U11033 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n7399), .ZN(n9968) );
  INV_X1 U11034 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10053) );
  NAND4_X1 U11035 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(SI_15_), .A3(
        P2_ADDR_REG_13__SCAN_IN), .A4(n10053), .ZN(n9966) );
  NAND4_X1 U11036 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .A3(P2_REG1_REG_13__SCAN_IN), .A4(P2_REG1_REG_5__SCAN_IN), .ZN(n9965)
         );
  NOR4_X1 U11037 ( .A1(n9968), .A2(n9967), .A3(n9966), .A4(n9965), .ZN(n9969)
         );
  NAND4_X1 U11038 ( .A1(n9970), .A2(P2_ADDR_REG_9__SCAN_IN), .A3(
        P2_ADDR_REG_18__SCAN_IN), .A4(n9969), .ZN(n9982) );
  NOR4_X1 U11039 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .A3(P2_REG1_REG_2__SCAN_IN), .A4(n10029), .ZN(n9975) );
  NOR4_X1 U11040 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(P1_REG0_REG_12__SCAN_IN), 
        .A3(n9999), .A4(n5616), .ZN(n9974) );
  NOR4_X1 U11041 ( .A1(SI_29_), .A2(n10002), .A3(n10005), .A4(n10004), .ZN(
        n9971) );
  NAND3_X1 U11042 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(n9971), .A3(
        P1_REG2_REG_15__SCAN_IN), .ZN(n9972) );
  NOR3_X1 U11043 ( .A1(n9972), .A2(n10015), .A3(P2_WR_REG_SCAN_IN), .ZN(n9973)
         );
  NAND3_X1 U11044 ( .A1(n9975), .A2(n9974), .A3(n9973), .ZN(n9981) );
  NAND4_X1 U11045 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .A3(P2_REG2_REG_12__SCAN_IN), .A4(P1_WR_REG_SCAN_IN), .ZN(n9980) );
  INV_X1 U11046 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10034) );
  INV_X1 U11047 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10031) );
  NOR3_X1 U11048 ( .A1(P2_REG0_REG_10__SCAN_IN), .A2(n10034), .A3(n10031), 
        .ZN(n9978) );
  NOR4_X1 U11049 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(P1_DATAO_REG_13__SCAN_IN), .A3(n10036), .A4(n10037), .ZN(n9977) );
  NOR4_X1 U11050 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P2_REG3_REG_5__SCAN_IN), .A4(n10050), .ZN(n9976) );
  NAND4_X1 U11051 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(n9978), .A3(n9977), .A4(
        n9976), .ZN(n9979) );
  NOR4_X1 U11052 ( .A1(n9982), .A2(n9981), .A3(n9980), .A4(n9979), .ZN(n10107)
         );
  AOI22_X1 U11053 ( .A1(n9985), .A2(keyinput34), .B1(keyinput14), .B2(n9984), 
        .ZN(n9983) );
  OAI221_X1 U11054 ( .B1(n9985), .B2(keyinput34), .C1(n9984), .C2(keyinput14), 
        .A(n9983), .ZN(n9997) );
  INV_X1 U11055 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U11056 ( .A1(n9988), .A2(keyinput4), .B1(keyinput15), .B2(n9987), 
        .ZN(n9986) );
  OAI221_X1 U11057 ( .B1(n9988), .B2(keyinput4), .C1(n9987), .C2(keyinput15), 
        .A(n9986), .ZN(n9996) );
  AOI22_X1 U11058 ( .A1(n9991), .A2(keyinput31), .B1(keyinput8), .B2(n9990), 
        .ZN(n9989) );
  OAI221_X1 U11059 ( .B1(n9991), .B2(keyinput31), .C1(n9990), .C2(keyinput8), 
        .A(n9989), .ZN(n9995) );
  AOI22_X1 U11060 ( .A1(n9993), .A2(keyinput22), .B1(keyinput44), .B2(n5092), 
        .ZN(n9992) );
  OAI221_X1 U11061 ( .B1(n9993), .B2(keyinput22), .C1(n5092), .C2(keyinput44), 
        .A(n9992), .ZN(n9994) );
  NOR4_X1 U11062 ( .A1(n9997), .A2(n9996), .A3(n9995), .A4(n9994), .ZN(n10045)
         );
  AOI22_X1 U11063 ( .A1(n5616), .A2(keyinput41), .B1(n9999), .B2(keyinput23), 
        .ZN(n9998) );
  OAI221_X1 U11064 ( .B1(n5616), .B2(keyinput41), .C1(n9999), .C2(keyinput23), 
        .A(n9998), .ZN(n10011) );
  INV_X1 U11065 ( .A(SI_29_), .ZN(n10001) );
  AOI22_X1 U11066 ( .A1(n10002), .A2(keyinput25), .B1(keyinput63), .B2(n10001), 
        .ZN(n10000) );
  OAI221_X1 U11067 ( .B1(n10002), .B2(keyinput25), .C1(n10001), .C2(keyinput63), .A(n10000), .ZN(n10010) );
  AOI22_X1 U11068 ( .A1(n10005), .A2(keyinput7), .B1(keyinput17), .B2(n10004), 
        .ZN(n10003) );
  OAI221_X1 U11069 ( .B1(n10005), .B2(keyinput7), .C1(n10004), .C2(keyinput17), 
        .A(n10003), .ZN(n10009) );
  XNOR2_X1 U11070 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput21), .ZN(n10007)
         );
  XNOR2_X1 U11071 ( .A(P1_REG0_REG_12__SCAN_IN), .B(keyinput37), .ZN(n10006)
         );
  NAND2_X1 U11072 ( .A1(n10007), .A2(n10006), .ZN(n10008) );
  NOR4_X1 U11073 ( .A1(n10011), .A2(n10010), .A3(n10009), .A4(n10008), .ZN(
        n10044) );
  AOI22_X1 U11074 ( .A1(n10013), .A2(keyinput24), .B1(keyinput61), .B2(n5020), 
        .ZN(n10012) );
  OAI221_X1 U11075 ( .B1(n10013), .B2(keyinput24), .C1(n5020), .C2(keyinput61), 
        .A(n10012), .ZN(n10026) );
  AOI22_X1 U11076 ( .A1(n10016), .A2(keyinput49), .B1(n10015), .B2(keyinput19), 
        .ZN(n10014) );
  OAI221_X1 U11077 ( .B1(n10016), .B2(keyinput49), .C1(n10015), .C2(keyinput19), .A(n10014), .ZN(n10025) );
  AOI22_X1 U11078 ( .A1(n10019), .A2(keyinput36), .B1(n10018), .B2(keyinput13), 
        .ZN(n10017) );
  OAI221_X1 U11079 ( .B1(n10019), .B2(keyinput36), .C1(n10018), .C2(keyinput13), .A(n10017), .ZN(n10024) );
  XOR2_X1 U11080 ( .A(n10020), .B(keyinput0), .Z(n10022) );
  XNOR2_X1 U11081 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput26), .ZN(n10021) );
  NAND2_X1 U11082 ( .A1(n10022), .A2(n10021), .ZN(n10023) );
  NOR4_X1 U11083 ( .A1(n10026), .A2(n10025), .A3(n10024), .A4(n10023), .ZN(
        n10043) );
  INV_X1 U11084 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10028) );
  AOI22_X1 U11085 ( .A1(n10029), .A2(keyinput57), .B1(n10028), .B2(keyinput28), 
        .ZN(n10027) );
  OAI221_X1 U11086 ( .B1(n10029), .B2(keyinput57), .C1(n10028), .C2(keyinput28), .A(n10027), .ZN(n10041) );
  AOI22_X1 U11087 ( .A1(n10031), .A2(keyinput10), .B1(n5197), .B2(keyinput58), 
        .ZN(n10030) );
  OAI221_X1 U11088 ( .B1(n10031), .B2(keyinput10), .C1(n5197), .C2(keyinput58), 
        .A(n10030), .ZN(n10040) );
  AOI22_X1 U11089 ( .A1(n10034), .A2(keyinput48), .B1(n10033), .B2(keyinput27), 
        .ZN(n10032) );
  OAI221_X1 U11090 ( .B1(n10034), .B2(keyinput48), .C1(n10033), .C2(keyinput27), .A(n10032), .ZN(n10039) );
  AOI22_X1 U11091 ( .A1(n10037), .A2(keyinput54), .B1(n10036), .B2(keyinput3), 
        .ZN(n10035) );
  OAI221_X1 U11092 ( .B1(n10037), .B2(keyinput54), .C1(n10036), .C2(keyinput3), 
        .A(n10035), .ZN(n10038) );
  NOR4_X1 U11093 ( .A1(n10041), .A2(n10040), .A3(n10039), .A4(n10038), .ZN(
        n10042) );
  NAND4_X1 U11094 ( .A1(n10045), .A2(n10044), .A3(n10043), .A4(n10042), .ZN(
        n10106) );
  AOI22_X1 U11095 ( .A1(n10047), .A2(keyinput35), .B1(keyinput42), .B2(n7399), 
        .ZN(n10046) );
  OAI221_X1 U11096 ( .B1(n10047), .B2(keyinput35), .C1(n7399), .C2(keyinput42), 
        .A(n10046), .ZN(n10059) );
  INV_X1 U11097 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10049) );
  AOI22_X1 U11098 ( .A1(n10050), .A2(keyinput16), .B1(keyinput46), .B2(n10049), 
        .ZN(n10048) );
  OAI221_X1 U11099 ( .B1(n10050), .B2(keyinput16), .C1(n10049), .C2(keyinput46), .A(n10048), .ZN(n10058) );
  AOI22_X1 U11100 ( .A1(n10053), .A2(keyinput62), .B1(n10052), .B2(keyinput20), 
        .ZN(n10051) );
  OAI221_X1 U11101 ( .B1(n10053), .B2(keyinput62), .C1(n10052), .C2(keyinput20), .A(n10051), .ZN(n10057) );
  XOR2_X1 U11102 ( .A(n10122), .B(keyinput29), .Z(n10055) );
  XNOR2_X1 U11103 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput2), .ZN(n10054) );
  NAND2_X1 U11104 ( .A1(n10055), .A2(n10054), .ZN(n10056) );
  NOR4_X1 U11105 ( .A1(n10059), .A2(n10058), .A3(n10057), .A4(n10056), .ZN(
        n10104) );
  AOI22_X1 U11106 ( .A1(n5090), .A2(keyinput53), .B1(n10061), .B2(keyinput45), 
        .ZN(n10060) );
  OAI221_X1 U11107 ( .B1(n5090), .B2(keyinput53), .C1(n10061), .C2(keyinput45), 
        .A(n10060), .ZN(n10066) );
  XNOR2_X1 U11108 ( .A(n10062), .B(keyinput38), .ZN(n10065) );
  XNOR2_X1 U11109 ( .A(n10063), .B(keyinput56), .ZN(n10064) );
  OR3_X1 U11110 ( .A1(n10066), .A2(n10065), .A3(n10064), .ZN(n10074) );
  AOI22_X1 U11111 ( .A1(n10068), .A2(keyinput18), .B1(keyinput39), .B2(n8112), 
        .ZN(n10067) );
  OAI221_X1 U11112 ( .B1(n10068), .B2(keyinput18), .C1(n8112), .C2(keyinput39), 
        .A(n10067), .ZN(n10073) );
  AOI22_X1 U11113 ( .A1(n10071), .A2(keyinput60), .B1(keyinput50), .B2(n10070), 
        .ZN(n10069) );
  OAI221_X1 U11114 ( .B1(n10071), .B2(keyinput60), .C1(n10070), .C2(keyinput50), .A(n10069), .ZN(n10072) );
  NOR3_X1 U11115 ( .A1(n10074), .A2(n10073), .A3(n10072), .ZN(n10103) );
  AOI22_X1 U11116 ( .A1(n10077), .A2(keyinput33), .B1(n10076), .B2(keyinput32), 
        .ZN(n10075) );
  OAI221_X1 U11117 ( .B1(n10077), .B2(keyinput33), .C1(n10076), .C2(keyinput32), .A(n10075), .ZN(n10087) );
  XNOR2_X1 U11118 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput1), .ZN(n10081) );
  XNOR2_X1 U11119 ( .A(SI_7_), .B(keyinput59), .ZN(n10080) );
  XNOR2_X1 U11120 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput11), .ZN(n10079)
         );
  XNOR2_X1 U11121 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput12), .ZN(n10078)
         );
  NAND4_X1 U11122 ( .A1(n10081), .A2(n10080), .A3(n10079), .A4(n10078), .ZN(
        n10086) );
  XNOR2_X1 U11123 ( .A(keyinput43), .B(n10082), .ZN(n10085) );
  XNOR2_X1 U11124 ( .A(keyinput52), .B(n10083), .ZN(n10084) );
  NOR4_X1 U11125 ( .A1(n10087), .A2(n10086), .A3(n10085), .A4(n10084), .ZN(
        n10102) );
  AOI22_X1 U11126 ( .A1(n10090), .A2(keyinput30), .B1(keyinput55), .B2(n10089), 
        .ZN(n10088) );
  OAI221_X1 U11127 ( .B1(n10090), .B2(keyinput30), .C1(n10089), .C2(keyinput55), .A(n10088), .ZN(n10100) );
  AOI22_X1 U11128 ( .A1(n10092), .A2(keyinput51), .B1(keyinput5), .B2(n6024), 
        .ZN(n10091) );
  OAI221_X1 U11129 ( .B1(n10092), .B2(keyinput51), .C1(n6024), .C2(keyinput5), 
        .A(n10091), .ZN(n10099) );
  AOI22_X1 U11130 ( .A1(n10094), .A2(keyinput6), .B1(keyinput40), .B2(n9958), 
        .ZN(n10093) );
  OAI221_X1 U11131 ( .B1(n10094), .B2(keyinput6), .C1(n9958), .C2(keyinput40), 
        .A(n10093), .ZN(n10098) );
  XNOR2_X1 U11132 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput47), .ZN(n10096) );
  XNOR2_X1 U11133 ( .A(SI_0_), .B(keyinput9), .ZN(n10095) );
  NAND2_X1 U11134 ( .A1(n10096), .A2(n10095), .ZN(n10097) );
  NOR4_X1 U11135 ( .A1(n10100), .A2(n10099), .A3(n10098), .A4(n10097), .ZN(
        n10101) );
  NAND4_X1 U11136 ( .A1(n10104), .A2(n10103), .A3(n10102), .A4(n10101), .ZN(
        n10105) );
  AOI211_X1 U11137 ( .C1(n10108), .C2(n10107), .A(n10106), .B(n10105), .ZN(
        n10115) );
  NOR2_X1 U11138 ( .A1(n10110), .A2(n10109), .ZN(n10111) );
  AOI211_X1 U11139 ( .C1(P2_DATAO_REG_23__SCAN_IN), .C2(n10113), .A(n10112), 
        .B(n10111), .ZN(n10114) );
  XNOR2_X1 U11140 ( .A(n10115), .B(n10114), .ZN(P1_U3330) );
  XOR2_X1 U11141 ( .A(n10116), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11142 ( .A1(n10118), .A2(n10117), .ZN(n10119) );
  XOR2_X1 U11143 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10119), .Z(ADD_1071_U51) );
  OAI21_X1 U11144 ( .B1(n10122), .B2(n10121), .A(n10120), .ZN(n10123) );
  XNOR2_X1 U11145 ( .A(n10123), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11146 ( .B1(n10126), .B2(n10125), .A(n10124), .ZN(ADD_1071_U47) );
  AOI21_X1 U11147 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(ADD_1071_U48) );
  XOR2_X1 U11148 ( .A(n10130), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11149 ( .A(n10131), .B(n10132), .Z(ADD_1071_U54) );
  XOR2_X1 U11150 ( .A(n10133), .B(n10134), .Z(ADD_1071_U53) );
  XNOR2_X1 U11151 ( .A(n10136), .B(n10135), .ZN(ADD_1071_U52) );
  INV_X1 U4773 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9659) );
  CLKBUF_X1 U4800 ( .A(n8145), .Z(n4371) );
  CLKBUF_X1 U4837 ( .A(n5302), .Z(n5579) );
  CLKBUF_X1 U4838 ( .A(n5065), .Z(n5350) );
  CLKBUF_X1 U4961 ( .A(n6944), .Z(n4256) );
  CLKBUF_X1 U5051 ( .A(n6064), .Z(n6021) );
  CLKBUF_X1 U5156 ( .A(n6841), .Z(n5928) );
  NAND2_X1 U5939 ( .A1(n7210), .A2(n7209), .ZN(n7494) );
endmodule

