

module b22_C_AntiSAT_k_128_6 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310;

  AOI211_X1 U7225 ( .C1(n13695), .C2(n14951), .A(n13694), .B(n13693), .ZN(
        n13771) );
  AND2_X1 U7226 ( .A1(n8195), .A2(n8197), .ZN(n11145) );
  NAND2_X1 U7227 ( .A1(n10305), .A2(n10818), .ZN(n8280) );
  NAND2_X2 U7228 ( .A1(n12205), .A2(n14294), .ZN(n12228) );
  AND4_X1 U7229 ( .A1(n7569), .A2(n7568), .A3(n7567), .A4(n7566), .ZN(n10753)
         );
  INV_X1 U7230 ( .A(n7646), .ZN(n8118) );
  INV_X1 U7231 ( .A(n10032), .ZN(n10029) );
  INV_X1 U7233 ( .A(n6483), .ZN(n12467) );
  CLKBUF_X2 U7234 ( .A(n12223), .Z(n12440) );
  INV_X1 U7235 ( .A(n12449), .ZN(n12451) );
  INV_X2 U7236 ( .A(n8731), .ZN(n9065) );
  INV_X2 U7237 ( .A(n8648), .ZN(n8731) );
  CLKBUF_X2 U7238 ( .A(n8839), .Z(n9023) );
  AND2_X1 U7239 ( .A1(n12001), .A2(n9175), .ZN(n9936) );
  INV_X1 U7240 ( .A(n6636), .ZN(n9249) );
  OR2_X1 U7241 ( .A1(n9191), .A2(n9168), .ZN(n6668) );
  BUF_X1 U7242 ( .A(n14824), .Z(n6482) );
  INV_X1 U7243 ( .A(n8482), .ZN(n13809) );
  NAND2_X1 U7244 ( .A1(n9922), .A2(n15025), .ZN(n6477) );
  NAND2_X1 U7245 ( .A1(n9922), .A2(n15025), .ZN(n6478) );
  CLKBUF_X1 U7246 ( .A(n13904), .Z(n6479) );
  NOR2_X1 U7247 ( .A1(n12462), .A2(n9616), .ZN(n13904) );
  OR2_X1 U7248 ( .A1(n12814), .A2(n12813), .ZN(n12815) );
  NOR2_X1 U7249 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n8433) );
  INV_X2 U7250 ( .A(n12205), .ZN(n12231) );
  INV_X1 U7251 ( .A(n13222), .ZN(n13178) );
  NAND2_X1 U7252 ( .A1(n13496), .A2(n13495), .ZN(n13494) );
  INV_X1 U7253 ( .A(n9936), .ZN(n12049) );
  INV_X2 U7254 ( .A(n10523), .ZN(n10532) );
  AND2_X1 U7255 ( .A1(n7482), .A2(n7483), .ZN(n7564) );
  INV_X1 U7256 ( .A(n7550), .ZN(n7797) );
  INV_X2 U7257 ( .A(n7828), .ZN(n7559) );
  OAI21_X1 U7258 ( .B1(n7778), .B2(n6993), .A(n6991), .ZN(n7819) );
  OR2_X1 U7259 ( .A1(n7776), .A2(n7775), .ZN(n7778) );
  NAND2_X1 U7260 ( .A1(n8608), .A2(n8607), .ZN(n10433) );
  OAI21_X1 U7261 ( .B1(n10940), .B2(n10939), .A(n10938), .ZN(n11037) );
  OAI21_X1 U7263 ( .B1(n13288), .B2(n13249), .A(n13494), .ZN(n13471) );
  OR2_X1 U7264 ( .A1(n10112), .A2(n9712), .ZN(n9828) );
  INV_X2 U7265 ( .A(n13521), .ZN(n13221) );
  NAND2_X1 U7266 ( .A1(n8440), .A2(n8469), .ZN(n9724) );
  AND2_X1 U7267 ( .A1(n10590), .A2(n10589), .ZN(n12292) );
  NAND2_X1 U7268 ( .A1(n8342), .A2(n8341), .ZN(n8669) );
  INV_X1 U7269 ( .A(n8328), .ZN(n9257) );
  NAND2_X1 U7270 ( .A1(n13233), .A2(n13235), .ZN(n13234) );
  INV_X1 U7271 ( .A(n13773), .ZN(n13475) );
  OR2_X1 U7272 ( .A1(n13411), .A2(n13408), .ZN(n13410) );
  NAND2_X1 U7273 ( .A1(n12164), .A2(n12163), .ZN(n14320) );
  AOI21_X1 U7274 ( .B1(n7207), .B2(n7204), .A(n6619), .ZN(n11084) );
  NAND2_X1 U7275 ( .A1(n7919), .A2(n7918), .ZN(n12906) );
  BUF_X1 U7277 ( .A(n9109), .Z(n13359) );
  INV_X1 U7278 ( .A(n10873), .ZN(n9869) );
  INV_X1 U7279 ( .A(n9579), .ZN(n12254) );
  NAND3_X1 U7280 ( .A1(n13759), .A2(n8731), .A3(n13404), .ZN(n6480) );
  OAI21_X2 U7281 ( .B1(n11704), .B2(n11703), .A(n11702), .ZN(n11871) );
  NAND2_X2 U7282 ( .A1(n11585), .A2(n11584), .ZN(n11704) );
  NAND2_X1 U7283 ( .A1(n14248), .A2(n14053), .ZN(n14233) );
  CLKBUF_X1 U7284 ( .A(n10447), .Z(n6481) );
  NAND2_X1 U7285 ( .A1(n6682), .A2(n8547), .ZN(n10447) );
  NOR2_X4 U7286 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9214) );
  OAI21_X2 U7287 ( .B1(n8919), .B2(n7029), .A(n7026), .ZN(n8393) );
  NAND2_X2 U7288 ( .A1(n8387), .A2(n8386), .ZN(n8919) );
  AOI21_X2 U7289 ( .B1(n11357), .B2(n11356), .A(n7435), .ZN(n11358) );
  XNOR2_X2 U7290 ( .A(n14483), .B(n6852), .ZN(n15302) );
  NAND2_X2 U7291 ( .A1(n14479), .A2(n14480), .ZN(n14483) );
  XNOR2_X2 U7292 ( .A(n14736), .B(n13972), .ZN(n12473) );
  NAND2_X2 U7293 ( .A1(n7480), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7474) );
  OAI21_X2 U7294 ( .B1(n11948), .B2(n11947), .A(n11946), .ZN(n13627) );
  OR2_X2 U7295 ( .A1(n14263), .A2(n14070), .ZN(n14072) );
  NAND2_X2 U7296 ( .A1(n9709), .A2(n13400), .ZN(n9792) );
  AND2_X2 U7297 ( .A1(n6913), .A2(n6912), .ZN(n10696) );
  OAI22_X2 U7298 ( .A1(n6651), .A2(n6650), .B1(n12878), .B2(n13092), .ZN(
        n12876) );
  NAND2_X2 U7299 ( .A1(n11823), .A2(n11822), .ZN(n14069) );
  AOI22_X2 U7300 ( .A1(n12456), .A2(n12455), .B1(n12454), .B2(n7306), .ZN(
        n12511) );
  XNOR2_X2 U7301 ( .A(n11923), .B(n11922), .ZN(n14989) );
  AND2_X2 U7302 ( .A1(n7087), .A2(n7086), .ZN(n11923) );
  AOI21_X2 U7303 ( .B1(n12880), .B2(n8297), .A(n8079), .ZN(n8106) );
  NOR2_X1 U7304 ( .A1(n10072), .A2(n10071), .ZN(n10529) );
  AOI21_X2 U7306 ( .B1(n14406), .B2(n14405), .A(n14404), .ZN(n14408) );
  OAI21_X2 U7307 ( .B1(n14459), .B2(n14401), .A(n6866), .ZN(n14406) );
  AOI21_X2 U7308 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n15143), .A(n8082), .ZN(
        n8116) );
  NAND2_X1 U7309 ( .A1(n10856), .A2(n12479), .ZN(n10894) );
  AOI21_X2 U7310 ( .B1(n14693), .B2(n10855), .A(n10854), .ZN(n10856) );
  NOR2_X2 U7311 ( .A1(n14233), .A2(n14076), .ZN(n14232) );
  XNOR2_X2 U7312 ( .A(n11539), .B(n11552), .ZN(n11258) );
  AND2_X2 U7313 ( .A1(n6924), .A2(n6923), .ZN(n11539) );
  AOI21_X1 U7314 ( .B1(n8544), .B2(n8543), .A(n8322), .ZN(n8569) );
  XNOR2_X2 U7315 ( .A(n7105), .B(P3_IR_REG_2__SCAN_IN), .ZN(n7529) );
  NOR2_X2 U7316 ( .A1(n10148), .A2(n7083), .ZN(n7105) );
  XNOR2_X2 U7317 ( .A(n7536), .B(P3_IR_REG_1__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U7318 ( .A1(n6697), .A2(n8349), .ZN(n8725) );
  NAND2_X1 U7319 ( .A1(n7984), .A2(n15067), .ZN(n8202) );
  NAND2_X1 U7320 ( .A1(n10421), .A2(n10420), .ZN(n10505) );
  NAND2_X2 U7321 ( .A1(n8179), .A2(n8174), .ZN(n10099) );
  INV_X2 U7322 ( .A(n12292), .ZN(n14736) );
  OAI21_X1 U7323 ( .B1(n12739), .B2(n6917), .A(n12738), .ZN(n12737) );
  AND4_X1 U7324 ( .A1(n7490), .A2(n7489), .A3(n7488), .A4(n7487), .ZN(n11270)
         );
  INV_X1 U7325 ( .A(n12287), .ZN(n12285) );
  AND3_X1 U7326 ( .A1(n7577), .A2(n7576), .A3(n7575), .ZN(n15051) );
  INV_X2 U7327 ( .A(n7596), .ZN(n8109) );
  INV_X1 U7328 ( .A(n15044), .ZN(n10559) );
  INV_X1 U7329 ( .A(n7595), .ZN(n7579) );
  BUF_X4 U7330 ( .A(n9794), .Z(n13222) );
  INV_X4 U7331 ( .A(n12228), .ZN(n12216) );
  INV_X1 U7332 ( .A(n13973), .ZN(n12286) );
  INV_X2 U7333 ( .A(n12230), .ZN(n9767) );
  BUF_X4 U7334 ( .A(n12449), .Z(n6483) );
  INV_X4 U7335 ( .A(n8280), .ZN(n10001) );
  INV_X1 U7336 ( .A(n14279), .ZN(n10475) );
  MUX2_X1 U7338 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8470), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n8471) );
  BUF_X1 U7339 ( .A(n7475), .Z(n7493) );
  AOI21_X1 U7340 ( .B1(n7361), .B2(n7496), .A(n7497), .ZN(n6877) );
  OR2_X1 U7341 ( .A1(n7495), .A2(n6879), .ZN(n6878) );
  CLKBUF_X2 U7342 ( .A(n7529), .Z(n10216) );
  XNOR2_X1 U7343 ( .A(n6848), .B(n6847), .ZN(n14824) );
  INV_X2 U7344 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7083) );
  AND2_X1 U7345 ( .A1(n12872), .A2(n14581), .ZN(n6638) );
  NAND2_X1 U7346 ( .A1(n12678), .A2(n12679), .ZN(n12677) );
  AOI21_X1 U7347 ( .B1(n11975), .B2(n13625), .A(n11974), .ZN(n13676) );
  NOR2_X1 U7348 ( .A1(n12875), .A2(n6649), .ZN(n6648) );
  INV_X1 U7349 ( .A(n6907), .ZN(n12875) );
  AND2_X1 U7350 ( .A1(n13677), .A2(n13675), .ZN(n6683) );
  AOI21_X1 U7351 ( .B1(n12417), .B2(n12416), .A(n6516), .ZN(n12420) );
  OR2_X1 U7352 ( .A1(n12876), .A2(n12881), .ZN(n6907) );
  XNOR2_X1 U7353 ( .A(n13174), .B(n13173), .ZN(n13199) );
  NAND3_X1 U7354 ( .A1(n12546), .A2(n12961), .A3(n12547), .ZN(n12657) );
  INV_X1 U7355 ( .A(n13418), .ZN(n13680) );
  NAND2_X1 U7356 ( .A1(n6739), .A2(n12543), .ZN(n12546) );
  NAND2_X1 U7357 ( .A1(n7792), .A2(n13000), .ZN(n13073) );
  NAND2_X1 U7358 ( .A1(n12545), .A2(n12544), .ZN(n12547) );
  AOI21_X2 U7359 ( .B1(n12972), .B2(n8007), .A(n7450), .ZN(n12958) );
  INV_X1 U7360 ( .A(n12598), .ZN(n12599) );
  NAND2_X1 U7361 ( .A1(n12665), .A2(n7060), .ZN(n6754) );
  NAND2_X1 U7362 ( .A1(n14072), .A2(n14071), .ZN(n14247) );
  NAND2_X1 U7363 ( .A1(n6637), .A2(n7177), .ZN(n14599) );
  NAND2_X1 U7364 ( .A1(n11801), .A2(n7146), .ZN(n14610) );
  INV_X1 U7365 ( .A(n12906), .ZN(n12878) );
  NAND2_X1 U7366 ( .A1(n6681), .A2(n6680), .ZN(n11801) );
  AND2_X1 U7367 ( .A1(n12037), .A2(n12036), .ZN(n14366) );
  AND2_X1 U7368 ( .A1(n7893), .A2(n7875), .ZN(n7892) );
  NAND2_X1 U7369 ( .A1(n11481), .A2(n11480), .ZN(n12008) );
  AND2_X1 U7370 ( .A1(n8852), .A2(n8851), .ZN(n11788) );
  NAND2_X1 U7371 ( .A1(n11059), .A2(n11058), .ZN(n11060) );
  NAND2_X1 U7372 ( .A1(n10824), .A2(n7979), .ZN(n10823) );
  OR2_X1 U7373 ( .A1(n11549), .A2(n11548), .ZN(n7087) );
  NAND2_X1 U7374 ( .A1(n11213), .A2(n11212), .ZN(n12329) );
  NOR2_X1 U7375 ( .A1(n11247), .A2(n11248), .ZN(n11545) );
  NAND2_X1 U7376 ( .A1(n8768), .A2(n8767), .ZN(n14813) );
  INV_X1 U7377 ( .A(n12320), .ZN(n14643) );
  NAND2_X1 U7378 ( .A1(n8790), .A2(n8789), .ZN(n13644) );
  AOI21_X1 U7379 ( .B1(n11873), .B2(n6491), .A(n6750), .ZN(n6749) );
  AND2_X1 U7380 ( .A1(n11057), .A2(n7443), .ZN(n11058) );
  XNOR2_X1 U7381 ( .A(n8749), .B(n8748), .ZN(n10976) );
  NAND2_X1 U7382 ( .A1(n7044), .A2(n7042), .ZN(n8786) );
  NAND2_X1 U7383 ( .A1(n8353), .A2(n7046), .ZN(n7044) );
  NAND2_X1 U7384 ( .A1(n6915), .A2(n6914), .ZN(n6913) );
  XNOR2_X1 U7385 ( .A(n8725), .B(n8724), .ZN(n10884) );
  NAND2_X1 U7386 ( .A1(n8725), .A2(n8350), .ZN(n8353) );
  NAND2_X1 U7387 ( .A1(n8713), .A2(n8712), .ZN(n11100) );
  NAND2_X1 U7388 ( .A1(n6673), .A2(n6867), .ZN(n14717) );
  AND2_X1 U7389 ( .A1(n8194), .A2(n8189), .ZN(n10822) );
  AND2_X1 U7390 ( .A1(n8180), .A2(n8184), .ZN(n10317) );
  NAND2_X1 U7391 ( .A1(n10029), .A2(n10031), .ZN(n8168) );
  NAND2_X1 U7392 ( .A1(n9947), .A2(n12285), .ZN(n10771) );
  NAND2_X1 U7393 ( .A1(n7968), .A2(n10032), .ZN(n8169) );
  OR2_X1 U7394 ( .A1(n7697), .A2(n11215), .ZN(n6934) );
  NAND2_X1 U7395 ( .A1(n14102), .A2(n14252), .ZN(n14282) );
  AND4_X1 U7396 ( .A1(n7524), .A2(n7523), .A3(n7522), .A4(n7521), .ZN(n7971)
         );
  AND3_X1 U7397 ( .A1(n7520), .A2(n7519), .A3(n7518), .ZN(n11073) );
  NAND2_X1 U7398 ( .A1(n6746), .A2(n6496), .ZN(n10028) );
  CLKBUF_X1 U7399 ( .A(n7595), .Z(n7596) );
  NAND2_X1 U7400 ( .A1(n7552), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n7539) );
  OAI211_X1 U7401 ( .C1(n7646), .C2(SI_3_), .A(n7425), .B(n6497), .ZN(n15044)
         );
  NAND4_X1 U7402 ( .A1(n8567), .A2(n7448), .A3(n8566), .A4(n8565), .ZN(n13358)
         );
  AOI21_X1 U7403 ( .B1(n7046), .B2(n7048), .A(n7043), .ZN(n7042) );
  INV_X1 U7404 ( .A(n10065), .ZN(n10466) );
  OR2_X1 U7405 ( .A1(n10217), .A2(n6522), .ZN(n7094) );
  AND2_X1 U7406 ( .A1(n7550), .A2(n12101), .ZN(n7535) );
  NAND2_X1 U7407 ( .A1(n7640), .A2(n7639), .ZN(n7654) );
  NAND2_X1 U7408 ( .A1(n7481), .A2(n7480), .ZN(n13137) );
  NAND2_X1 U7409 ( .A1(n7479), .A2(n7478), .ZN(n7481) );
  NAND2_X2 U7410 ( .A1(n10491), .A2(n9770), .ZN(n12230) );
  OR2_X1 U7411 ( .A1(n7638), .A2(n7637), .ZN(n7640) );
  AOI21_X1 U7412 ( .B1(n10181), .B2(n10153), .A(n10154), .ZN(n10217) );
  NAND4_X1 U7414 ( .A1(n9657), .A2(n9656), .A3(n9655), .A4(n9654), .ZN(n13974)
         );
  OAI21_X1 U7415 ( .B1(n12445), .B2(n9578), .A(n12258), .ZN(n12449) );
  NAND2_X1 U7416 ( .A1(n11732), .A2(n9166), .ZN(n9770) );
  AOI22_X1 U7417 ( .A1(n9062), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n6482), .B2(
        n8909), .ZN(n6682) );
  AND2_X1 U7418 ( .A1(n8477), .A2(n9124), .ZN(n9708) );
  INV_X2 U7419 ( .A(n9003), .ZN(n9061) );
  NAND2_X1 U7420 ( .A1(n12447), .A2(n12257), .ZN(n12262) );
  NAND2_X1 U7421 ( .A1(n8467), .A2(n9090), .ZN(n11348) );
  AOI21_X1 U7422 ( .B1(n8668), .B2(n8345), .A(n8685), .ZN(n7039) );
  OAI21_X1 U7423 ( .B1(n12833), .B2(n10305), .A(n10521), .ZN(n6660) );
  OR2_X2 U7424 ( .A1(n12461), .A2(n12447), .ZN(n14294) );
  AND2_X1 U7425 ( .A1(n8461), .A2(n8463), .ZN(n9124) );
  INV_X1 U7426 ( .A(n8361), .ZN(n7043) );
  XNOR2_X1 U7427 ( .A(n7950), .B(P3_IR_REG_22__SCAN_IN), .ZN(n10818) );
  INV_X1 U7428 ( .A(n14394), .ZN(n9175) );
  NAND2_X1 U7429 ( .A1(n8444), .A2(n8443), .ZN(n13816) );
  NAND2_X1 U7430 ( .A1(n7418), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7417) );
  NAND2_X1 U7431 ( .A1(n9173), .A2(n14387), .ZN(n14394) );
  OAI21_X1 U7432 ( .B1(n12101), .B2(n9261), .A(n8333), .ZN(n8335) );
  NAND2_X2 U7433 ( .A1(n6636), .A2(P1_U3086), .ZN(n14391) );
  XNOR2_X1 U7434 ( .A(n8321), .B(SI_1_), .ZN(n8544) );
  NAND2_X2 U7435 ( .A1(n12101), .A2(P1_U3086), .ZN(n14396) );
  OAI21_X1 U7436 ( .B1(n7558), .B2(n7506), .A(n7507), .ZN(n7571) );
  MUX2_X1 U7437 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8439), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n8440) );
  INV_X2 U7438 ( .A(n10968), .ZN(n6484) );
  OR2_X1 U7439 ( .A1(n9172), .A2(n14386), .ZN(n9169) );
  BUF_X2 U7440 ( .A(n9257), .Z(n6636) );
  NOR2_X2 U7441 ( .A1(n8818), .A2(n8450), .ZN(n8796) );
  INV_X4 U7442 ( .A(n9257), .ZN(n12101) );
  XNOR2_X1 U7443 ( .A(n14408), .B(n14407), .ZN(n14467) );
  OAI21_X1 U7444 ( .B1(n8328), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n8318), .ZN(
        n8321) );
  AND2_X1 U7445 ( .A1(n8460), .A2(n8459), .ZN(n8466) );
  NAND2_X1 U7446 ( .A1(n8454), .A2(n8448), .ZN(n8818) );
  OR2_X1 U7447 ( .A1(n7597), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7599) );
  AND2_X1 U7448 ( .A1(n8454), .A2(n8456), .ZN(n8460) );
  AND3_X2 U7449 ( .A1(n6868), .A2(n6523), .A3(n6869), .ZN(n9157) );
  AND2_X1 U7450 ( .A1(n7421), .A2(n8436), .ZN(n7419) );
  AND2_X1 U7451 ( .A1(n7438), .A2(n7422), .ZN(n7421) );
  INV_X1 U7452 ( .A(n7560), .ZN(n7457) );
  NOR2_X1 U7453 ( .A1(n6489), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n7358) );
  AND2_X1 U7454 ( .A1(n7290), .A2(n8433), .ZN(n7289) );
  NAND2_X1 U7455 ( .A1(n7477), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7478) );
  AND2_X1 U7456 ( .A1(n9299), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7637) );
  XNOR2_X1 U7457 ( .A(n14402), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n14459) );
  INV_X1 U7458 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6998) );
  INV_X1 U7459 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8831) );
  INV_X1 U7460 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9215) );
  INV_X1 U7461 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8449) );
  NOR2_X1 U7462 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8430) );
  INV_X1 U7463 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14402) );
  INV_X1 U7464 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8459) );
  INV_X1 U7465 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9445) );
  NOR2_X1 U7466 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n8420) );
  NOR2_X1 U7467 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n8421) );
  INV_X1 U7468 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8465) );
  INV_X4 U7469 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7470 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6689) );
  INV_X2 U7471 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7472 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7655) );
  INV_X1 U7473 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7624) );
  INV_X1 U7474 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n7359) );
  INV_X4 U7475 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  OR2_X2 U7476 ( .A1(n7750), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n6509) );
  NOR2_X2 U7477 ( .A1(n12781), .A2(n6921), .ZN(n12805) );
  NOR2_X2 U7478 ( .A1(n12751), .A2(n12750), .ZN(n12781) );
  NAND2_X1 U7479 ( .A1(n7424), .A2(n14083), .ZN(n14200) );
  AOI21_X1 U7480 ( .B1(n7020), .B2(n6538), .A(n7022), .ZN(n7019) );
  NOR2_X2 U7481 ( .A1(n10241), .A2(n15100), .ZN(n10273) );
  NOR2_X1 U7482 ( .A1(n14996), .A2(n15259), .ZN(n14995) );
  NOR2_X4 U7483 ( .A1(n6507), .A2(n14320), .ZN(n14168) );
  OR2_X4 U7484 ( .A1(n6502), .A2(n14327), .ZN(n6507) );
  OAI222_X1 U7485 ( .A1(P1_U3086), .A2(n11945), .B1(n14391), .B2(n11944), .C1(
        n15143), .C2(n14396), .ZN(P1_U3327) );
  NOR2_X2 U7486 ( .A1(n14995), .A2(n11918), .ZN(n11919) );
  AOI21_X2 U7487 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n12752), .A(n12746), .ZN(
        n12747) );
  NOR2_X2 U7488 ( .A1(n11919), .A2(n11929), .ZN(n12746) );
  OAI21_X2 U7489 ( .B1(n10853), .B2(n10852), .A(n10851), .ZN(n14693) );
  AND2_X1 U7490 ( .A1(n13490), .A2(n6758), .ZN(n13417) );
  NOR2_X2 U7491 ( .A1(n13700), .A2(n13505), .ZN(n13490) );
  NOR2_X2 U7492 ( .A1(n10005), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10087) );
  NOR2_X2 U7493 ( .A1(n14223), .A2(n14346), .ZN(n14208) );
  NOR3_X4 U7494 ( .A1(n10897), .A2(n6870), .A3(n6871), .ZN(n11483) );
  INV_X1 U7495 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n6910) );
  AOI21_X1 U7496 ( .B1(n7372), .B2(n7373), .A(n11979), .ZN(n7371) );
  AND3_X1 U7497 ( .A1(n8428), .A2(n8427), .A3(n8426), .ZN(n7438) );
  INV_X1 U7498 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8426) );
  INV_X1 U7499 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8424) );
  INV_X1 U7500 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8423) );
  INV_X1 U7501 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8448) );
  NAND2_X1 U7502 ( .A1(n8817), .A2(n6736), .ZN(n6738) );
  NOR2_X1 U7503 ( .A1(n7035), .A2(n6737), .ZN(n6736) );
  INV_X1 U7504 ( .A(n8816), .ZN(n6737) );
  INV_X1 U7505 ( .A(n8107), .ZN(n7965) );
  CLKBUF_X3 U7506 ( .A(n7563), .Z(n8108) );
  AND2_X2 U7507 ( .A1(n11943), .A2(n7483), .ZN(n7563) );
  INV_X1 U7508 ( .A(n7535), .ZN(n7646) );
  AOI21_X1 U7509 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14430), .A(n14429), .ZN(
        n14447) );
  NOR2_X1 U7510 ( .A1(n14449), .A2(n14448), .ZN(n14429) );
  INV_X1 U7511 ( .A(n8594), .ZN(n7267) );
  NOR2_X1 U7512 ( .A1(n8597), .A2(n8594), .ZN(n7268) );
  NAND2_X1 U7513 ( .A1(n6822), .A2(n12316), .ZN(n6821) );
  NAND2_X1 U7514 ( .A1(n7307), .A2(n6823), .ZN(n6822) );
  NOR2_X1 U7515 ( .A1(n6820), .A2(n12316), .ZN(n6819) );
  INV_X1 U7516 ( .A(n6823), .ZN(n6820) );
  INV_X1 U7517 ( .A(n12398), .ZN(n6827) );
  INV_X1 U7518 ( .A(n10737), .ZN(n7232) );
  NAND2_X1 U7519 ( .A1(n13526), .A2(n13340), .ZN(n7401) );
  INV_X1 U7520 ( .A(n8336), .ZN(n6722) );
  AOI21_X1 U7521 ( .B1(n7064), .B2(n7062), .A(n7061), .ZN(n7060) );
  INV_X1 U7522 ( .A(n12647), .ZN(n7061) );
  INV_X1 U7523 ( .A(n7065), .ZN(n7062) );
  NAND2_X1 U7524 ( .A1(n10407), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6912) );
  NOR2_X1 U7525 ( .A1(n12896), .A2(n12906), .ZN(n6650) );
  NAND2_X1 U7526 ( .A1(n11943), .A2(n13137), .ZN(n7595) );
  NAND2_X1 U7527 ( .A1(n12720), .A2(n15044), .ZN(n8184) );
  BUF_X1 U7528 ( .A(n6757), .Z(n6755) );
  AND2_X1 U7529 ( .A1(n7780), .A2(n7777), .ZN(n6994) );
  NAND2_X1 U7530 ( .A1(n6934), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6933) );
  AND2_X1 U7531 ( .A1(n9348), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7677) );
  INV_X1 U7532 ( .A(n6984), .ZN(n6980) );
  INV_X1 U7533 ( .A(n6510), .ZN(n6978) );
  NOR2_X1 U7534 ( .A1(n7642), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7656) );
  NAND2_X1 U7535 ( .A1(n9070), .A2(n9069), .ZN(n7278) );
  OR2_X1 U7536 ( .A1(n13680), .A2(n13436), .ZN(n11968) );
  AND2_X1 U7537 ( .A1(n7246), .A2(n6567), .ZN(n7244) );
  NOR2_X1 U7538 ( .A1(n11951), .A2(n7250), .ZN(n7249) );
  INV_X1 U7539 ( .A(n11950), .ZN(n7250) );
  NAND2_X1 U7540 ( .A1(n13571), .A2(n13576), .ZN(n11981) );
  XNOR2_X1 U7541 ( .A(n9109), .B(n10447), .ZN(n9712) );
  INV_X1 U7542 ( .A(n8584), .ZN(n8435) );
  AND2_X1 U7543 ( .A1(n8431), .A2(n8430), .ZN(n8432) );
  INV_X1 U7544 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6997) );
  NAND2_X1 U7545 ( .A1(n14310), .A2(n14090), .ZN(n7127) );
  NOR2_X1 U7546 ( .A1(n6506), .A2(n7132), .ZN(n7131) );
  INV_X1 U7547 ( .A(n9933), .ZN(n7132) );
  AND2_X1 U7548 ( .A1(n7165), .A2(n10765), .ZN(n7162) );
  OR2_X1 U7549 ( .A1(n7168), .A2(n7170), .ZN(n7165) );
  NAND2_X1 U7550 ( .A1(n8418), .A2(n8417), .ZN(n8500) );
  OAI21_X1 U7551 ( .B1(n9000), .B2(n7052), .A(n7051), .ZN(n9031) );
  INV_X1 U7552 ( .A(n7053), .ZN(n7052) );
  AOI21_X1 U7553 ( .B1(n8401), .B2(n7053), .A(n6613), .ZN(n7051) );
  NOR2_X1 U7554 ( .A1(n7054), .A2(n8526), .ZN(n7053) );
  INV_X1 U7555 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6828) );
  NOR2_X2 U7556 ( .A1(n9143), .A2(n9140), .ZN(n6869) );
  NAND4_X1 U7557 ( .A1(n9255), .A2(n9266), .A3(n9139), .A4(n9138), .ZN(n9140)
         );
  INV_X1 U7558 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9139) );
  INV_X1 U7559 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9138) );
  AND2_X1 U7560 ( .A1(n8377), .A2(n8376), .ZN(n8816) );
  NAND2_X1 U7561 ( .A1(n8372), .A2(n8371), .ZN(n8817) );
  NAND2_X1 U7562 ( .A1(n8830), .A2(n8829), .ZN(n8372) );
  INV_X4 U7563 ( .A(n10532), .ZN(n12567) );
  NAND2_X1 U7564 ( .A1(n6754), .A2(n6752), .ZN(n12598) );
  NOR2_X1 U7565 ( .A1(n6753), .A2(n12601), .ZN(n6752) );
  INV_X1 U7566 ( .A(n7058), .ZN(n6753) );
  OR2_X1 U7567 ( .A1(n8101), .A2(n12572), .ZN(n8301) );
  AOI21_X1 U7568 ( .B1(n12852), .B2(n8130), .A(n8137), .ZN(n8308) );
  OR2_X1 U7569 ( .A1(n8130), .A2(n12852), .ZN(n6990) );
  AND2_X1 U7570 ( .A1(n7088), .A2(n7089), .ZN(n10394) );
  NAND2_X1 U7571 ( .A1(n7090), .A2(n11138), .ZN(n7089) );
  NAND2_X1 U7572 ( .A1(n12766), .A2(n12765), .ZN(n7091) );
  NAND2_X1 U7573 ( .A1(n7093), .A2(n12765), .ZN(n7092) );
  INV_X1 U7574 ( .A(n11924), .ZN(n7093) );
  AND2_X1 U7575 ( .A1(n7891), .A2(n8279), .ZN(n7352) );
  NAND2_X1 U7576 ( .A1(n7890), .A2(n8281), .ZN(n12924) );
  INV_X1 U7577 ( .A(n7994), .ZN(n6904) );
  NOR2_X1 U7578 ( .A1(n11678), .A2(n7449), .ZN(n7337) );
  NAND2_X1 U7579 ( .A1(n11313), .A2(n7989), .ZN(n11383) );
  INV_X1 U7580 ( .A(n12960), .ZN(n13019) );
  NAND2_X1 U7581 ( .A1(n10040), .A2(n10001), .ZN(n12964) );
  AND2_X1 U7582 ( .A1(n8135), .A2(n8064), .ZN(n12960) );
  AND2_X1 U7583 ( .A1(n9908), .A2(n13131), .ZN(n9998) );
  AND2_X1 U7584 ( .A1(n7894), .A2(n7893), .ZN(n7909) );
  INV_X1 U7585 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7461) );
  AOI21_X1 U7586 ( .B1(n6929), .B2(n6931), .A(n6599), .ZN(n6927) );
  NAND2_X1 U7587 ( .A1(n6732), .A2(n13177), .ZN(n6731) );
  NAND2_X1 U7588 ( .A1(n13234), .A2(n6711), .ZN(n6719) );
  NOR2_X1 U7589 ( .A1(n6526), .A2(n13172), .ZN(n6711) );
  NAND2_X2 U7590 ( .A1(n8472), .A2(n13809), .ZN(n8589) );
  BUF_X1 U7591 ( .A(n8481), .Z(n8472) );
  NAND2_X1 U7592 ( .A1(n13804), .A2(n13809), .ZN(n8839) );
  NAND2_X1 U7593 ( .A1(n8796), .A2(n6521), .ZN(n8890) );
  NOR2_X1 U7594 ( .A1(n13680), .A2(n6759), .ZN(n6758) );
  INV_X1 U7595 ( .A(n6760), .ZN(n6759) );
  NAND2_X1 U7596 ( .A1(n13482), .A2(n11964), .ZN(n7234) );
  INV_X1 U7597 ( .A(n7398), .ZN(n7397) );
  OAI21_X1 U7598 ( .B1(n13535), .B2(n7399), .A(n7402), .ZN(n7398) );
  NAND2_X1 U7599 ( .A1(n7403), .A2(n11984), .ZN(n7399) );
  AOI21_X1 U7600 ( .B1(n7371), .B2(n7368), .A(n6564), .ZN(n7367) );
  INV_X1 U7601 ( .A(n7373), .ZN(n7368) );
  OR2_X1 U7602 ( .A1(n11977), .A2(n7369), .ZN(n7366) );
  INV_X1 U7603 ( .A(n7371), .ZN(n7369) );
  OR2_X1 U7604 ( .A1(n11172), .A2(n11171), .ZN(n7253) );
  NAND2_X1 U7605 ( .A1(n9098), .A2(n12101), .ZN(n9003) );
  NAND2_X2 U7606 ( .A1(n9724), .A2(n13816), .ZN(n9098) );
  OR2_X1 U7607 ( .A1(n13554), .A2(n6694), .ZN(n6693) );
  INV_X1 U7608 ( .A(n6695), .ZN(n6694) );
  INV_X1 U7609 ( .A(n13590), .ZN(n13733) );
  INV_X2 U7610 ( .A(n9098), .ZN(n8909) );
  INV_X1 U7611 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U7612 ( .A1(n7222), .A2(n6539), .ZN(n7221) );
  NAND2_X1 U7613 ( .A1(n11720), .A2(n7223), .ZN(n7222) );
  NAND2_X1 U7614 ( .A1(n11425), .A2(n7224), .ZN(n7220) );
  AND2_X1 U7615 ( .A1(n6505), .A2(n11720), .ZN(n7224) );
  OR2_X1 U7616 ( .A1(n14003), .A2(n6781), .ZN(n6780) );
  AND2_X1 U7617 ( .A1(n14004), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6781) );
  NAND2_X1 U7618 ( .A1(n12424), .A2(n12423), .ZN(n14297) );
  INV_X1 U7619 ( .A(n14062), .ZN(n14303) );
  NAND2_X1 U7620 ( .A1(n14151), .A2(n7173), .ZN(n7172) );
  NOR2_X1 U7621 ( .A1(n14133), .A2(n7176), .ZN(n7173) );
  XNOR2_X1 U7622 ( .A(n14310), .B(n13959), .ZN(n14133) );
  NAND2_X1 U7623 ( .A1(n14200), .A2(n7181), .ZN(n7183) );
  NOR2_X1 U7624 ( .A1(n14183), .A2(n7182), .ZN(n7181) );
  INV_X1 U7625 ( .A(n14085), .ZN(n7182) );
  AOI21_X1 U7626 ( .B1(n6642), .B2(n6493), .A(n6641), .ZN(n7424) );
  INV_X1 U7627 ( .A(n7160), .ZN(n6641) );
  AOI21_X1 U7628 ( .B1(n14081), .B2(n7161), .A(n6515), .ZN(n7160) );
  NAND2_X1 U7629 ( .A1(n14366), .A2(n14051), .ZN(n14052) );
  NAND2_X1 U7630 ( .A1(n14265), .A2(n14366), .ZN(n14264) );
  INV_X1 U7631 ( .A(n14366), .ZN(n14267) );
  AND2_X1 U7632 ( .A1(n12487), .A2(n12344), .ZN(n7146) );
  OR2_X1 U7633 ( .A1(n13953), .A2(n11631), .ZN(n12344) );
  INV_X2 U7634 ( .A(n12141), .ZN(n12457) );
  NAND2_X1 U7635 ( .A1(n12287), .A2(n13973), .ZN(n7170) );
  INV_X1 U7636 ( .A(n9157), .ZN(n9164) );
  OR2_X1 U7637 ( .A1(n8886), .A2(n8885), .ZN(n8906) );
  OAI22_X1 U7638 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14992), .B1(n14447), 
        .B2(n14431), .ZN(n14510) );
  NAND2_X1 U7639 ( .A1(n7861), .A2(n7860), .ZN(n12940) );
  AOI21_X1 U7640 ( .B1(n12868), .B2(n7787), .A(n7946), .ZN(n12877) );
  INV_X1 U7641 ( .A(n7001), .ZN(n7000) );
  INV_X1 U7642 ( .A(n7004), .ZN(n7002) );
  NAND2_X1 U7643 ( .A1(n14660), .A2(n14659), .ZN(n14507) );
  NAND2_X1 U7644 ( .A1(n6849), .A2(n6625), .ZN(n14509) );
  INV_X1 U7645 ( .A(n14659), .ZN(n6625) );
  NAND2_X1 U7646 ( .A1(n8611), .A2(n8612), .ZN(n8610) );
  NOR2_X1 U7647 ( .A1(n12276), .A2(n12275), .ZN(n12283) );
  NAND2_X1 U7648 ( .A1(n12300), .A2(n7324), .ZN(n7323) );
  INV_X1 U7649 ( .A(n12299), .ZN(n7324) );
  AND2_X1 U7650 ( .A1(n12313), .A2(n7308), .ZN(n7307) );
  AND2_X1 U7651 ( .A1(n8757), .A2(n7274), .ZN(n7273) );
  INV_X1 U7652 ( .A(n8755), .ZN(n7274) );
  NAND2_X1 U7653 ( .A1(n8758), .A2(n8755), .ZN(n7272) );
  NAND2_X1 U7654 ( .A1(n12312), .A2(n6816), .ZN(n6815) );
  NAND2_X1 U7655 ( .A1(n6818), .A2(n6817), .ZN(n6816) );
  NAND2_X1 U7656 ( .A1(n6814), .A2(n6821), .ZN(n6813) );
  INV_X1 U7657 ( .A(n6818), .ZN(n6814) );
  NAND2_X1 U7658 ( .A1(n6789), .A2(n6788), .ZN(n12338) );
  NAND2_X1 U7659 ( .A1(n12330), .A2(n12332), .ZN(n6788) );
  NAND2_X1 U7660 ( .A1(n12338), .A2(n12337), .ZN(n6787) );
  AOI21_X1 U7661 ( .B1(n12376), .B2(n6792), .A(n6797), .ZN(n6796) );
  OAI21_X1 U7662 ( .B1(n12376), .B2(n6795), .A(n6790), .ZN(n6794) );
  INV_X1 U7663 ( .A(n12387), .ZN(n7319) );
  OR2_X1 U7664 ( .A1(n12402), .A2(n12400), .ZN(n7316) );
  OR2_X1 U7665 ( .A1(n6827), .A2(n12399), .ZN(n6825) );
  NAND2_X1 U7666 ( .A1(n12399), .A2(n6827), .ZN(n6826) );
  NAND2_X1 U7667 ( .A1(n12408), .A2(n12407), .ZN(n7328) );
  AOI21_X1 U7668 ( .B1(n12404), .B2(n6801), .A(n6799), .ZN(n6798) );
  NOR2_X1 U7669 ( .A1(n7870), .A2(n6956), .ZN(n6955) );
  INV_X1 U7670 ( .A(n7858), .ZN(n6956) );
  INV_X1 U7671 ( .A(n7621), .ZN(n6942) );
  MUX2_X1 U7672 ( .A(n13426), .B(n13672), .S(n9065), .Z(n8508) );
  NAND2_X1 U7673 ( .A1(n12256), .A2(n12255), .ZN(n12445) );
  INV_X1 U7674 ( .A(n7169), .ZN(n7168) );
  INV_X1 U7675 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6811) );
  INV_X1 U7676 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U7677 ( .A1(n6703), .A2(n6702), .ZN(n6701) );
  INV_X1 U7678 ( .A(n6705), .ZN(n6703) );
  INV_X1 U7679 ( .A(n6707), .ZN(n6702) );
  AOI21_X1 U7680 ( .B1(n6709), .B2(n6708), .A(n8847), .ZN(n6705) );
  NAND2_X1 U7681 ( .A1(n8358), .A2(n9287), .ZN(n8361) );
  OR2_X1 U7682 ( .A1(n9298), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9346) );
  OAI21_X1 U7683 ( .B1(n12101), .B2(n6663), .A(n6662), .ZN(n8344) );
  NAND2_X1 U7684 ( .A1(n12101), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6662) );
  INV_X1 U7685 ( .A(n9257), .ZN(n7149) );
  NAND2_X1 U7686 ( .A1(n12101), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8333) );
  INV_X1 U7687 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14403) );
  NAND2_X1 U7688 ( .A1(n12657), .A2(n12547), .ZN(n12551) );
  INV_X1 U7689 ( .A(n11061), .ZN(n7076) );
  INV_X1 U7690 ( .A(n11374), .ZN(n7077) );
  INV_X1 U7691 ( .A(n11943), .ZN(n7482) );
  INV_X1 U7692 ( .A(n13137), .ZN(n7483) );
  NAND2_X1 U7693 ( .A1(n12772), .A2(n6614), .ZN(n7113) );
  NOR2_X1 U7694 ( .A1(n12897), .A2(n7357), .ZN(n7356) );
  AND2_X1 U7695 ( .A1(n6518), .A2(n8139), .ZN(n6894) );
  NOR2_X1 U7696 ( .A1(n6885), .A2(n6884), .ZN(n6883) );
  INV_X1 U7697 ( .A(n6503), .ZN(n6885) );
  NOR2_X1 U7698 ( .A1(n13000), .A2(n6887), .ZN(n6886) );
  NAND2_X1 U7699 ( .A1(n7767), .A2(n12632), .ZN(n7785) );
  INV_X1 U7700 ( .A(n7768), .ZN(n7767) );
  NAND2_X1 U7701 ( .A1(n7705), .A2(n11707), .ZN(n7723) );
  INV_X1 U7702 ( .A(n7335), .ZN(n7334) );
  OAI21_X1 U7703 ( .B1(n11145), .B2(n7336), .A(n7613), .ZN(n7335) );
  INV_X1 U7704 ( .A(n8195), .ZN(n7336) );
  INV_X1 U7705 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10225) );
  NAND2_X1 U7706 ( .A1(n7970), .A2(n7969), .ZN(n10100) );
  OR2_X1 U7707 ( .A1(n7550), .A2(n10012), .ZN(n7537) );
  NAND2_X1 U7708 ( .A1(n8030), .A2(n11579), .ZN(n6747) );
  XNOR2_X1 U7709 ( .A(n8032), .B(P3_B_REG_SCAN_IN), .ZN(n8030) );
  NAND2_X1 U7710 ( .A1(n7082), .A2(n7084), .ZN(n7081) );
  NAND2_X1 U7711 ( .A1(n7949), .A2(n7083), .ZN(n7080) );
  NOR2_X1 U7712 ( .A1(n7949), .A2(n7083), .ZN(n7082) );
  OR2_X1 U7713 ( .A1(n7694), .A2(n7693), .ZN(n7696) );
  NOR2_X1 U7714 ( .A1(n7604), .A2(n6948), .ZN(n6947) );
  INV_X1 U7715 ( .A(n7510), .ZN(n6948) );
  NAND2_X1 U7716 ( .A1(n9276), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7512) );
  INV_X1 U7717 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7515) );
  AND2_X1 U7718 ( .A1(n13434), .A2(n7384), .ZN(n7383) );
  NAND2_X1 U7719 ( .A1(n7386), .A2(n7385), .ZN(n7384) );
  INV_X1 U7720 ( .A(n7389), .ZN(n7385) );
  NAND2_X1 U7721 ( .A1(n6513), .A2(n11987), .ZN(n7388) );
  XNOR2_X1 U7722 ( .A(n6764), .B(n13325), .ZN(n13434) );
  NOR2_X1 U7723 ( .A1(n13475), .A2(n13688), .ZN(n6762) );
  NOR2_X1 U7724 ( .A1(n6768), .A2(n13526), .ZN(n6767) );
  INV_X1 U7725 ( .A(n6769), .ZN(n6768) );
  INV_X1 U7726 ( .A(n11566), .ZN(n7410) );
  NOR2_X1 U7727 ( .A1(n6517), .A2(n7408), .ZN(n7407) );
  INV_X1 U7728 ( .A(n7439), .ZN(n7408) );
  AOI21_X1 U7729 ( .B1(n6490), .B2(n7230), .A(n6560), .ZN(n7229) );
  INV_X1 U7730 ( .A(n10736), .ZN(n7230) );
  INV_X1 U7731 ( .A(n6490), .ZN(n7231) );
  INV_X1 U7732 ( .A(n10356), .ZN(n7377) );
  OR2_X1 U7733 ( .A1(n7394), .A2(n7392), .ZN(n7391) );
  INV_X1 U7734 ( .A(n7401), .ZN(n7392) );
  INV_X1 U7735 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7282) );
  OR2_X1 U7736 ( .A1(n8584), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n8619) );
  OR2_X1 U7737 ( .A1(n13883), .A2(n12017), .ZN(n7210) );
  INV_X1 U7738 ( .A(n13902), .ZN(n7199) );
  AND2_X1 U7739 ( .A1(n13855), .A2(n6530), .ZN(n7201) );
  NAND2_X1 U7740 ( .A1(n12426), .A2(n12425), .ZN(n7305) );
  NAND2_X1 U7741 ( .A1(n12430), .A2(n12429), .ZN(n7304) );
  NOR2_X1 U7742 ( .A1(n12482), .A2(n7158), .ZN(n7157) );
  NOR2_X1 U7743 ( .A1(n11207), .A2(n7159), .ZN(n7158) );
  INV_X1 U7744 ( .A(n11209), .ZN(n7159) );
  NOR2_X1 U7745 ( .A1(n12478), .A2(n10892), .ZN(n10893) );
  OAI21_X1 U7746 ( .B1(n10615), .B2(n6506), .A(n10617), .ZN(n7135) );
  NAND2_X1 U7747 ( .A1(n7168), .A2(n10765), .ZN(n7166) );
  OR2_X1 U7748 ( .A1(n14088), .A2(n14087), .ZN(n7431) );
  NAND2_X1 U7749 ( .A1(n9881), .A2(n12279), .ZN(n9934) );
  NOR2_X1 U7750 ( .A1(n7314), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n7313) );
  NAND2_X1 U7751 ( .A1(n9167), .A2(n9193), .ZN(n7314) );
  AND3_X1 U7752 ( .A1(n9150), .A2(n9149), .A3(n9148), .ZN(n9155) );
  NAND2_X1 U7753 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n6809) );
  AND2_X1 U7754 ( .A1(n6488), .A2(n6811), .ZN(n6807) );
  OAI22_X1 U7755 ( .A1(n6488), .A2(n6809), .B1(P1_IR_REG_31__SCAN_IN), .B2(
        P1_IR_REG_22__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U7756 ( .A1(n6738), .A2(n6500), .ZN(n8905) );
  OR2_X1 U7757 ( .A1(n8786), .A2(n8366), .ZN(n6698) );
  AOI21_X1 U7758 ( .B1(n6708), .B2(n8365), .A(SI_14_), .ZN(n6707) );
  NAND2_X1 U7759 ( .A1(n8786), .A2(n8785), .ZN(n6704) );
  AND2_X1 U7760 ( .A1(n8365), .A2(SI_14_), .ZN(n6709) );
  NOR2_X1 U7761 ( .A1(n8748), .A2(n7050), .ZN(n7049) );
  INV_X1 U7762 ( .A(n8352), .ZN(n7050) );
  OR2_X1 U7763 ( .A1(n10342), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n9298) );
  OR2_X1 U7764 ( .A1(n9259), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9264) );
  NAND2_X1 U7765 ( .A1(n14402), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6866) );
  NOR2_X1 U7766 ( .A1(n14413), .A2(n14412), .ZN(n14415) );
  XNOR2_X1 U7767 ( .A(n14415), .B(n14414), .ZN(n14471) );
  OAI22_X1 U7768 ( .A1(n14477), .A2(n14418), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14476), .ZN(n14419) );
  AOI21_X1 U7769 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n10279), .A(n14422), .ZN(
        n14489) );
  NOR2_X1 U7770 ( .A1(n14454), .A2(n14453), .ZN(n14422) );
  AOI21_X1 U7771 ( .B1(n14424), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n14423), .ZN(
        n14425) );
  AND2_X1 U7772 ( .A1(n14490), .A2(n14489), .ZN(n14423) );
  AOI21_X1 U7773 ( .B1(n7060), .B2(n7063), .A(n6558), .ZN(n7058) );
  INV_X1 U7774 ( .A(n7064), .ZN(n7063) );
  AND2_X1 U7775 ( .A1(n12561), .A2(n12559), .ZN(n12610) );
  INV_X1 U7776 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10156) );
  INV_X1 U7777 ( .A(n11267), .ZN(n11052) );
  NOR2_X1 U7778 ( .A1(n12590), .A2(n7066), .ZN(n7065) );
  NOR2_X1 U7779 ( .A1(n12667), .A2(n12537), .ZN(n7066) );
  AND4_X1 U7780 ( .A1(n7603), .A2(n7602), .A3(n7601), .A4(n7600), .ZN(n11074)
         );
  NAND2_X1 U7781 ( .A1(n10015), .A2(n10016), .ZN(n10161) );
  NAND2_X1 U7782 ( .A1(n10282), .A2(n10281), .ZN(n7090) );
  NOR2_X1 U7783 ( .A1(n10245), .A2(n11138), .ZN(n10284) );
  INV_X1 U7784 ( .A(n10276), .ZN(n6914) );
  AND2_X1 U7785 ( .A1(n10407), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10393) );
  INV_X1 U7786 ( .A(n11256), .ZN(n10702) );
  OR2_X1 U7787 ( .A1(n10395), .A2(n10396), .ZN(n7109) );
  NAND2_X1 U7788 ( .A1(n11256), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n6923) );
  NOR2_X1 U7789 ( .A1(n11258), .A2(n14582), .ZN(n11540) );
  NAND2_X1 U7790 ( .A1(n11921), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7086) );
  NOR2_X1 U7791 ( .A1(n11916), .A2(n6922), .ZN(n11917) );
  AND2_X1 U7792 ( .A1(n11921), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6922) );
  OAI21_X1 U7793 ( .B1(n12792), .B2(n12791), .A(n12790), .ZN(n12793) );
  AND2_X1 U7794 ( .A1(n12783), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U7795 ( .A1(n12816), .A2(n12815), .ZN(n12817) );
  INV_X1 U7796 ( .A(n12838), .ZN(n7101) );
  NAND2_X1 U7797 ( .A1(n6963), .A2(n6966), .ZN(n6962) );
  NAND2_X1 U7798 ( .A1(n7925), .A2(n12579), .ZN(n7941) );
  AND2_X1 U7799 ( .A1(n12876), .A2(n12881), .ZN(n6649) );
  NOR2_X1 U7800 ( .A1(n12877), .A2(n12962), .ZN(n6647) );
  NOR2_X1 U7801 ( .A1(n12878), .A2(n12964), .ZN(n6646) );
  INV_X1 U7802 ( .A(n12920), .ZN(n12890) );
  OAI21_X1 U7803 ( .B1(n12586), .B2(n13100), .A(n12917), .ZN(n12905) );
  INV_X1 U7804 ( .A(n12904), .ZN(n12910) );
  NAND2_X1 U7805 ( .A1(n6893), .A2(n6518), .ZN(n6892) );
  INV_X1 U7806 ( .A(n6895), .ZN(n6893) );
  AOI21_X1 U7807 ( .B1(n8139), .B2(n8138), .A(n6514), .ZN(n6895) );
  NAND2_X1 U7808 ( .A1(n12958), .A2(n6894), .ZN(n6888) );
  OAI21_X1 U7809 ( .B1(n12958), .B2(n6891), .A(n6889), .ZN(n12932) );
  INV_X1 U7810 ( .A(n6890), .ZN(n6889) );
  OAI21_X1 U7811 ( .B1(n6894), .B2(n6891), .A(n12939), .ZN(n6890) );
  INV_X1 U7812 ( .A(n6892), .ZN(n6891) );
  INV_X1 U7813 ( .A(n12976), .ZN(n12950) );
  AOI21_X1 U7814 ( .B1(n7343), .B2(n7345), .A(n7342), .ZN(n7341) );
  INV_X1 U7815 ( .A(n8271), .ZN(n7342) );
  INV_X1 U7816 ( .A(n7344), .ZN(n7343) );
  OR2_X1 U7817 ( .A1(n12983), .A2(n12963), .ZN(n8266) );
  AND2_X1 U7818 ( .A1(n8263), .A2(n8262), .ZN(n12993) );
  AND2_X1 U7819 ( .A1(n7998), .A2(n7996), .ZN(n6902) );
  AND2_X1 U7820 ( .A1(n8235), .A2(n8245), .ZN(n11886) );
  AND2_X1 U7821 ( .A1(n7712), .A2(n8225), .ZN(n7339) );
  OR2_X1 U7822 ( .A1(n14573), .A2(n12713), .ZN(n8225) );
  AND2_X1 U7823 ( .A1(n7669), .A2(n7668), .ZN(n11510) );
  NOR2_X1 U7824 ( .A1(n6542), .A2(n6901), .ZN(n6900) );
  INV_X1 U7825 ( .A(n7985), .ZN(n6901) );
  INV_X1 U7826 ( .A(n7427), .ZN(n6896) );
  NAND2_X1 U7827 ( .A1(n6899), .A2(n6897), .ZN(n11313) );
  NOR2_X1 U7828 ( .A1(n7427), .A2(n6898), .ZN(n6897) );
  NAND2_X1 U7829 ( .A1(n11133), .A2(n11132), .ZN(n11131) );
  AND2_X1 U7830 ( .A1(n7982), .A2(n7981), .ZN(n6908) );
  AND2_X1 U7831 ( .A1(n10455), .A2(n7978), .ZN(n10824) );
  INV_X1 U7832 ( .A(n13022), .ZN(n12962) );
  NAND2_X1 U7833 ( .A1(n9699), .A2(n9698), .ZN(n9705) );
  NAND2_X1 U7834 ( .A1(n7924), .A2(n7923), .ZN(n13036) );
  INV_X1 U7835 ( .A(n9246), .ZN(n6911) );
  AND2_X1 U7836 ( .A1(n9919), .A2(n10001), .ZN(n13022) );
  NOR2_X2 U7837 ( .A1(n8013), .A2(n7360), .ZN(n7497) );
  NAND2_X1 U7838 ( .A1(n7471), .A2(n7361), .ZN(n7360) );
  NOR2_X1 U7839 ( .A1(n8022), .A2(n7083), .ZN(n8023) );
  INV_X1 U7840 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8022) );
  INV_X1 U7841 ( .A(n8025), .ZN(n8027) );
  AND2_X1 U7842 ( .A1(n15118), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6938) );
  NOR2_X1 U7843 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), .ZN(
        n6756) );
  INV_X1 U7844 ( .A(n6953), .ZN(n6952) );
  INV_X1 U7845 ( .A(n7825), .ZN(n7823) );
  INV_X1 U7846 ( .A(n6992), .ZN(n6991) );
  OAI22_X1 U7847 ( .A1(n6994), .A2(n6993), .B1(n11187), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6992) );
  NAND2_X1 U7848 ( .A1(n6608), .A2(n7793), .ZN(n6993) );
  AND2_X1 U7849 ( .A1(n7793), .A2(n7779), .ZN(n7780) );
  NAND2_X1 U7850 ( .A1(n7778), .A2(n6994), .ZN(n7794) );
  NAND2_X1 U7851 ( .A1(n7731), .A2(n7730), .ZN(n7733) );
  NAND2_X1 U7852 ( .A1(n6933), .A2(n7713), .ZN(n7731) );
  INV_X1 U7853 ( .A(n6933), .ZN(n6932) );
  INV_X1 U7854 ( .A(n7653), .ZN(n6986) );
  INV_X1 U7855 ( .A(n7654), .ZN(n6982) );
  AOI21_X1 U7856 ( .B1(n6985), .B2(n7662), .A(n6562), .ZN(n6984) );
  INV_X1 U7857 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7664) );
  OR2_X1 U7858 ( .A1(n7658), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n7680) );
  NOR2_X1 U7859 ( .A1(n9304), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n6985) );
  XNOR2_X1 U7860 ( .A(n7643), .B(P3_IR_REG_9__SCAN_IN), .ZN(n10697) );
  OR2_X1 U7861 ( .A1(n7701), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7642) );
  INV_X1 U7862 ( .A(n6947), .ZN(n6946) );
  XNOR2_X1 U7863 ( .A(n6663), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n7621) );
  AOI21_X1 U7864 ( .B1(n6947), .B2(n6945), .A(n6944), .ZN(n6943) );
  INV_X1 U7865 ( .A(n7512), .ZN(n6944) );
  INV_X1 U7866 ( .A(n7586), .ZN(n6945) );
  OR2_X1 U7867 ( .A1(n7607), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7701) );
  XNOR2_X1 U7868 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7586) );
  AND2_X1 U7869 ( .A1(n9250), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7506) );
  INV_X1 U7870 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7456) );
  AND2_X1 U7871 ( .A1(n13192), .A2(n13189), .ZN(n7009) );
  NAND2_X1 U7872 ( .A1(n6729), .A2(n13243), .ZN(n6728) );
  INV_X1 U7873 ( .A(n10581), .ZN(n7022) );
  INV_X1 U7874 ( .A(n11897), .ZN(n7013) );
  AND2_X1 U7875 ( .A1(n13146), .A2(n11897), .ZN(n7011) );
  NAND2_X1 U7876 ( .A1(n13162), .A2(n7006), .ZN(n6735) );
  NAND2_X1 U7877 ( .A1(n11614), .A2(n7017), .ZN(n14804) );
  INV_X1 U7878 ( .A(n13172), .ZN(n6718) );
  NOR2_X1 U7879 ( .A1(n6526), .A2(n13172), .ZN(n6717) );
  AND2_X1 U7880 ( .A1(n7008), .A2(n13156), .ZN(n7007) );
  INV_X1 U7881 ( .A(n13314), .ZN(n7008) );
  AOI21_X1 U7882 ( .B1(n9067), .B2(n9066), .A(n7451), .ZN(n7275) );
  OR2_X1 U7883 ( .A1(n9071), .A2(n7446), .ZN(n7451) );
  NAND2_X1 U7884 ( .A1(n9039), .A2(n9038), .ZN(n9066) );
  AND3_X1 U7885 ( .A1(n8882), .A2(n8881), .A3(n8880), .ZN(n13263) );
  OR3_X1 U7886 ( .A1(n9745), .A2(n9746), .A3(n11908), .ZN(n9137) );
  OAI21_X1 U7887 ( .B1(n6482), .B2(P2_REG2_REG_1__SCAN_IN), .A(n6644), .ZN(
        n14826) );
  NAND2_X1 U7888 ( .A1(n6482), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6644) );
  AOI21_X1 U7889 ( .B1(n11860), .B2(P2_REG2_REG_13__SCAN_IN), .A(n11852), .ZN(
        n11854) );
  AND2_X1 U7890 ( .A1(n8427), .A2(n8428), .ZN(n7290) );
  INV_X1 U7891 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8451) );
  XNOR2_X1 U7892 ( .A(n6829), .B(n13395), .ZN(n13396) );
  NOR2_X1 U7893 ( .A1(n13394), .A2(n13393), .ZN(n6829) );
  INV_X1 U7894 ( .A(n11990), .ZN(n11969) );
  NAND2_X1 U7895 ( .A1(n13432), .A2(n13438), .ZN(n13433) );
  AND2_X1 U7896 ( .A1(n8519), .A2(n8518), .ZN(n13418) );
  AND4_X1 U7897 ( .A1(n8515), .A2(n8514), .A3(n8513), .A4(n8512), .ZN(n13436)
         );
  INV_X1 U7898 ( .A(n13434), .ZN(n13438) );
  NOR2_X1 U7899 ( .A1(n7241), .A2(n7240), .ZN(n7239) );
  AND2_X1 U7900 ( .A1(n13495), .A2(n11964), .ZN(n7240) );
  INV_X1 U7901 ( .A(n13470), .ZN(n7241) );
  NAND2_X1 U7902 ( .A1(n11963), .A2(n11962), .ZN(n13482) );
  OR2_X1 U7903 ( .A1(n13482), .A2(n13495), .ZN(n13484) );
  NOR2_X1 U7904 ( .A1(n13535), .A2(n7404), .ZN(n7400) );
  AND2_X1 U7905 ( .A1(n7397), .A2(n11958), .ZN(n7394) );
  AND2_X1 U7906 ( .A1(n7366), .A2(n7364), .ZN(n13577) );
  INV_X1 U7907 ( .A(n7367), .ZN(n7365) );
  OR2_X1 U7908 ( .A1(n13626), .A2(n7374), .ZN(n7372) );
  NAND2_X1 U7909 ( .A1(n13744), .A2(n13345), .ZN(n7373) );
  INV_X1 U7910 ( .A(n13575), .ZN(n13628) );
  NOR2_X1 U7911 ( .A1(n11976), .A2(n13629), .ZN(n7374) );
  OR2_X1 U7912 ( .A1(n14594), .A2(n11621), .ZN(n7439) );
  OR2_X1 U7913 ( .A1(n14813), .A2(n13348), .ZN(n11566) );
  NOR2_X1 U7914 ( .A1(n7254), .A2(n7252), .ZN(n7251) );
  INV_X1 U7915 ( .A(n11173), .ZN(n7252) );
  AOI21_X1 U7916 ( .B1(n11180), .B2(n11179), .A(n11178), .ZN(n11565) );
  AND2_X1 U7917 ( .A1(n11310), .A2(n13349), .ZN(n11178) );
  NAND2_X1 U7918 ( .A1(n11161), .A2(n11160), .ZN(n11172) );
  NAND2_X1 U7919 ( .A1(n11156), .A2(n11155), .ZN(n11180) );
  NAND2_X1 U7920 ( .A1(n9953), .A2(n10358), .ZN(n10357) );
  XNOR2_X1 U7921 ( .A(n10355), .B(n13356), .ZN(n10358) );
  INV_X1 U7922 ( .A(n13631), .ZN(n13466) );
  INV_X1 U7923 ( .A(n9641), .ZN(n6635) );
  NAND2_X1 U7924 ( .A1(n8505), .A2(n8504), .ZN(n8507) );
  NAND2_X1 U7925 ( .A1(n13796), .A2(n9061), .ZN(n8505) );
  NAND2_X1 U7926 ( .A1(n8446), .A2(n8445), .ZN(n13411) );
  NAND2_X1 U7927 ( .A1(n9005), .A2(n9004), .ZN(n13700) );
  OR2_X1 U7928 ( .A1(n12142), .A2(n9003), .ZN(n9005) );
  INV_X1 U7929 ( .A(n14967), .ZN(n14939) );
  INV_X1 U7930 ( .A(n14951), .ZN(n13751) );
  INV_X1 U7931 ( .A(n8765), .ZN(n8447) );
  NAND2_X1 U7932 ( .A1(n7194), .A2(n7192), .ZN(n13837) );
  AOI21_X1 U7933 ( .B1(n6492), .B2(n6519), .A(n7193), .ZN(n7192) );
  INV_X1 U7934 ( .A(n13838), .ZN(n7193) );
  AOI21_X1 U7935 ( .B1(n13824), .B2(n12201), .A(n12221), .ZN(n7190) );
  INV_X1 U7936 ( .A(n7190), .ZN(n7188) );
  NAND2_X1 U7937 ( .A1(n13901), .A2(n13902), .ZN(n7202) );
  INV_X1 U7938 ( .A(n13875), .ZN(n7213) );
  NAND2_X1 U7939 ( .A1(n7202), .A2(n7201), .ZN(n13913) );
  NOR2_X1 U7940 ( .A1(n7219), .A2(n7221), .ZN(n7218) );
  INV_X1 U7941 ( .A(n11722), .ZN(n7219) );
  OR2_X1 U7942 ( .A1(n10673), .A2(n7204), .ZN(n6561) );
  OR2_X1 U7943 ( .A1(n10674), .A2(n10673), .ZN(n7207) );
  NAND2_X1 U7944 ( .A1(n13867), .A2(n12182), .ZN(n13935) );
  NAND2_X1 U7945 ( .A1(n13828), .A2(n12014), .ZN(n12016) );
  OR2_X1 U7946 ( .A1(n12016), .A2(n12017), .ZN(n7216) );
  OR2_X1 U7947 ( .A1(n9404), .A2(n9403), .ZN(n6777) );
  OR2_X1 U7948 ( .A1(n9628), .A2(n9627), .ZN(n6775) );
  NOR2_X1 U7949 ( .A1(n13982), .A2(n13981), .ZN(n14003) );
  XNOR2_X1 U7950 ( .A(n6780), .B(n14019), .ZN(n14005) );
  NAND2_X1 U7951 ( .A1(n12460), .A2(n12459), .ZN(n14035) );
  NAND2_X1 U7952 ( .A1(n12434), .A2(n12433), .ZN(n14034) );
  NAND2_X1 U7953 ( .A1(n14145), .A2(n7118), .ZN(n7116) );
  NOR2_X1 U7954 ( .A1(n7119), .A2(n7120), .ZN(n7118) );
  INV_X1 U7955 ( .A(n7123), .ZN(n7120) );
  AND2_X1 U7956 ( .A1(n7115), .A2(n7126), .ZN(n6670) );
  NAND2_X1 U7957 ( .A1(n14303), .A2(n14065), .ZN(n7126) );
  NAND2_X1 U7958 ( .A1(n7117), .A2(n14063), .ZN(n7115) );
  INV_X1 U7959 ( .A(n7122), .ZN(n7117) );
  NAND2_X1 U7960 ( .A1(n7172), .A2(n6540), .ZN(n14117) );
  AND2_X1 U7961 ( .A1(n12236), .A2(n12208), .ZN(n14136) );
  NAND2_X1 U7962 ( .A1(n14168), .A2(n14156), .ZN(n14142) );
  NOR2_X1 U7963 ( .A1(n14351), .A2(n14077), .ZN(n14055) );
  NAND2_X1 U7964 ( .A1(n6642), .A2(n14220), .ZN(n14217) );
  NAND2_X1 U7965 ( .A1(n14247), .A2(n14073), .ZN(n7179) );
  AND2_X1 U7966 ( .A1(n12380), .A2(n14053), .ZN(n14249) );
  OAI21_X1 U7967 ( .B1(n14050), .B2(n14049), .A(n14048), .ZN(n14273) );
  XNOR2_X1 U7968 ( .A(n14267), .B(n14051), .ZN(n14272) );
  INV_X1 U7969 ( .A(n12486), .ZN(n6680) );
  OR2_X1 U7970 ( .A1(n14778), .A2(n10888), .ZN(n10980) );
  NAND2_X1 U7971 ( .A1(n10894), .A2(n10893), .ZN(n10981) );
  NAND2_X1 U7972 ( .A1(n9934), .A2(n9933), .ZN(n10616) );
  NAND2_X1 U7973 ( .A1(n12285), .A2(n12286), .ZN(n7169) );
  AOI21_X1 U7974 ( .B1(n14297), .B2(n14735), .A(n14296), .ZN(n6875) );
  NAND2_X1 U7975 ( .A1(n12204), .A2(n12203), .ZN(n14310) );
  NAND2_X1 U7976 ( .A1(n12084), .A2(n12083), .ZN(n14346) );
  NAND2_X1 U7977 ( .A1(n11488), .A2(n12485), .ZN(n14638) );
  INV_X1 U7978 ( .A(n11489), .ZN(n11488) );
  INV_X1 U7979 ( .A(n14294), .ZN(n14749) );
  NAND2_X1 U7980 ( .A1(n10488), .A2(n10495), .ZN(n14735) );
  INV_X1 U7981 ( .A(n14770), .ZN(n14710) );
  NAND2_X1 U7982 ( .A1(n7171), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9191) );
  NAND2_X1 U7983 ( .A1(n9157), .A2(n7312), .ZN(n7171) );
  INV_X1 U7984 ( .A(n7314), .ZN(n7312) );
  INV_X1 U7985 ( .A(n9170), .ZN(n6667) );
  XNOR2_X1 U7986 ( .A(n9031), .B(n9030), .ZN(n12183) );
  NAND2_X1 U7987 ( .A1(n7030), .A2(n7031), .ZN(n8387) );
  INV_X1 U7988 ( .A(n8391), .ZN(n7029) );
  INV_X1 U7989 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9185) );
  INV_X1 U7990 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9145) );
  NAND2_X1 U7991 ( .A1(n6868), .A2(n6869), .ZN(n9156) );
  NAND2_X1 U7992 ( .A1(n8378), .A2(n8377), .ZN(n8795) );
  NOR2_X1 U7993 ( .A1(n9264), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9267) );
  NAND2_X1 U7994 ( .A1(n9267), .A2(n9266), .ZN(n10342) );
  XNOR2_X1 U7995 ( .A(n14471), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14472) );
  NAND2_X1 U7996 ( .A1(n14469), .A2(n14470), .ZN(n14473) );
  OAI21_X1 U7997 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n14433), .A(n14432), .ZN(
        n14444) );
  NAND2_X1 U7998 ( .A1(n12677), .A2(n12564), .ZN(n6743) );
  INV_X1 U7999 ( .A(n11874), .ZN(n11879) );
  NAND2_X1 U8000 ( .A1(n7940), .A2(n7939), .ZN(n12575) );
  NAND2_X1 U8001 ( .A1(n12692), .A2(n12688), .ZN(n12621) );
  NAND2_X1 U8002 ( .A1(n7754), .A2(n7753), .ZN(n12627) );
  NAND2_X1 U8003 ( .A1(n9922), .A2(n15025), .ZN(n12674) );
  AND4_X1 U8004 ( .A1(n7585), .A2(n7584), .A3(n7583), .A4(n7582), .ZN(n11147)
         );
  AND4_X1 U8005 ( .A1(n7760), .A2(n7759), .A3(n7758), .A4(n7757), .ZN(n12698)
         );
  AOI21_X1 U8006 ( .B1(n8133), .B2(n8132), .A(n7437), .ZN(n8134) );
  NOR2_X1 U8007 ( .A1(n8158), .A2(n6987), .ZN(n8159) );
  INV_X1 U8008 ( .A(n7349), .ZN(n7348) );
  OAI21_X1 U8009 ( .B1(n8312), .B2(n10970), .A(n8316), .ZN(n7349) );
  INV_X1 U8010 ( .A(n8311), .ZN(n8312) );
  NAND2_X1 U8011 ( .A1(n7888), .A2(n7887), .ZN(n12935) );
  INV_X1 U8012 ( .A(n8001), .ZN(n13004) );
  NAND4_X1 U8013 ( .A1(n7652), .A2(n7651), .A3(n7650), .A4(n7649), .ZN(n11505)
         );
  NOR2_X1 U8014 ( .A1(n11543), .A2(n11542), .ZN(n11916) );
  AOI21_X1 U8015 ( .B1(n12810), .B2(n12809), .A(n12808), .ZN(n12829) );
  XNOR2_X1 U8016 ( .A(n6684), .B(n12843), .ZN(n12844) );
  NAND2_X1 U8017 ( .A1(n6686), .A2(n6685), .ZN(n6684) );
  NOR2_X1 U8018 ( .A1(n8098), .A2(n8097), .ZN(n8099) );
  NAND2_X1 U8019 ( .A1(n8012), .A2(n6639), .ZN(n12867) );
  NOR2_X1 U8020 ( .A1(n6589), .A2(n6640), .ZN(n6639) );
  INV_X1 U8021 ( .A(n13036), .ZN(n12885) );
  NAND2_X1 U8022 ( .A1(n7912), .A2(n7911), .ZN(n12896) );
  NAND2_X1 U8023 ( .A1(n7353), .A2(n8279), .ZN(n12923) );
  NAND2_X1 U8024 ( .A1(n15106), .A2(n15065), .ZN(n13087) );
  NAND2_X1 U8025 ( .A1(n8085), .A2(n8084), .ZN(n8101) );
  INV_X1 U8026 ( .A(n12575), .ZN(n12870) );
  NAND2_X1 U8027 ( .A1(n7799), .A2(n7798), .ZN(n13120) );
  NAND2_X1 U8028 ( .A1(n15089), .A2(n15065), .ZN(n13129) );
  XNOR2_X1 U8029 ( .A(n7796), .B(n7085), .ZN(n12833) );
  OAI21_X1 U8030 ( .B1(n7781), .B2(n6623), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7796) );
  NAND2_X1 U8031 ( .A1(n7795), .A2(n7465), .ZN(n6623) );
  OR2_X1 U8032 ( .A1(n7719), .A2(n7718), .ZN(n12752) );
  NAND2_X1 U8033 ( .A1(n8911), .A2(n8910), .ZN(n6696) );
  OR2_X1 U8034 ( .A1(n13214), .A2(n13215), .ZN(n6690) );
  INV_X1 U8035 ( .A(n7015), .ZN(n7014) );
  OAI21_X1 U8036 ( .B1(n7017), .B2(n7016), .A(n11620), .ZN(n7015) );
  INV_X1 U8037 ( .A(n14805), .ZN(n7016) );
  NAND2_X1 U8038 ( .A1(n9807), .A2(n13639), .ZN(n14812) );
  INV_X1 U8039 ( .A(n13436), .ZN(n13338) );
  INV_X1 U8040 ( .A(n7363), .ZN(n8540) );
  OR2_X1 U8041 ( .A1(P2_U3088), .A2(n9137), .ZN(n13360) );
  INV_X1 U8042 ( .A(n13396), .ZN(n13398) );
  NOR2_X1 U8043 ( .A1(n9458), .A2(n9455), .ZN(n14876) );
  NAND2_X1 U8044 ( .A1(n7263), .A2(n7261), .ZN(n13682) );
  INV_X1 U8045 ( .A(n7262), .ZN(n7261) );
  NAND2_X1 U8046 ( .A1(n7264), .A2(n13625), .ZN(n7263) );
  OAI22_X1 U8047 ( .A1(n13436), .A2(n13631), .B1(n13575), .B2(n13437), .ZN(
        n7262) );
  NAND2_X1 U8048 ( .A1(n8948), .A2(n8947), .ZN(n13539) );
  OR2_X1 U8049 ( .A1(n12081), .A2(n9003), .ZN(n8948) );
  NAND2_X1 U8050 ( .A1(n7245), .A2(n7246), .ZN(n13563) );
  OR2_X1 U8051 ( .A1(n13624), .A2(n7248), .ZN(n7245) );
  AND2_X1 U8052 ( .A1(n8893), .A2(n8892), .ZN(n13590) );
  NAND2_X2 U8053 ( .A1(n14925), .A2(n9806), .ZN(n13639) );
  NAND2_X1 U8054 ( .A1(n8546), .A2(n8545), .ZN(n8547) );
  CLKBUF_X1 U8055 ( .A(n8441), .Z(n8444) );
  INV_X1 U8056 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10949) );
  OAI22_X1 U8057 ( .A1(n11084), .A2(n11083), .B1(n11082), .B2(n11081), .ZN(
        n11357) );
  NAND2_X1 U8058 ( .A1(n12125), .A2(n12124), .ZN(n14332) );
  NAND2_X1 U8059 ( .A1(n13935), .A2(n13936), .ZN(n13934) );
  NOR2_X1 U8060 ( .A1(n10654), .A2(n10655), .ZN(n10674) );
  XNOR2_X1 U8061 ( .A(n10672), .B(n10671), .ZN(n10654) );
  AOI21_X1 U8062 ( .B1(n12040), .B2(n9930), .A(n6556), .ZN(n9931) );
  INV_X1 U8063 ( .A(n13955), .ZN(n13937) );
  NAND2_X1 U8064 ( .A1(n11630), .A2(n11629), .ZN(n13953) );
  AND2_X1 U8065 ( .A1(n6777), .A2(n6776), .ZN(n9628) );
  NAND2_X1 U8066 ( .A1(n7152), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6776) );
  NOR2_X1 U8067 ( .A1(n9389), .A2(n9388), .ZN(n9475) );
  INV_X1 U8068 ( .A(n14034), .ZN(n14293) );
  NAND2_X1 U8069 ( .A1(n14096), .A2(n6876), .ZN(n14295) );
  OR2_X1 U8070 ( .A1(n14097), .A2(n14107), .ZN(n6876) );
  INV_X1 U8071 ( .A(n14150), .ZN(n14609) );
  OR2_X1 U8072 ( .A1(n11732), .A2(n9293), .ZN(n9584) );
  INV_X1 U8073 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10948) );
  NAND2_X1 U8074 ( .A1(n6861), .A2(n6860), .ZN(n14667) );
  NAND2_X1 U8075 ( .A1(n14663), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U8076 ( .A1(n6863), .A2(n14887), .ZN(n6862) );
  INV_X1 U8077 ( .A(n14529), .ZN(n6856) );
  NAND2_X1 U8078 ( .A1(n6859), .A2(n6858), .ZN(n6857) );
  INV_X1 U8079 ( .A(n8632), .ZN(n7298) );
  OR2_X1 U8080 ( .A1(n7295), .A2(n8675), .ZN(n7294) );
  INV_X1 U8081 ( .A(n8674), .ZN(n7295) );
  NAND2_X1 U8082 ( .A1(n7301), .A2(n8714), .ZN(n7300) );
  NAND2_X1 U8083 ( .A1(n12299), .A2(n12301), .ZN(n7325) );
  INV_X1 U8084 ( .A(n12311), .ZN(n7308) );
  INV_X1 U8085 ( .A(n6819), .ZN(n6817) );
  AOI21_X1 U8086 ( .B1(n7273), .B2(n7272), .A(n7271), .ZN(n7270) );
  INV_X1 U8087 ( .A(n8791), .ZN(n7287) );
  AND2_X1 U8088 ( .A1(n12319), .A2(n7310), .ZN(n7309) );
  INV_X1 U8089 ( .A(n12317), .ZN(n7310) );
  AND2_X1 U8090 ( .A1(n8854), .A2(n7285), .ZN(n7284) );
  NAND2_X1 U8091 ( .A1(n7286), .A2(n8791), .ZN(n7285) );
  AOI21_X1 U8092 ( .B1(n6787), .B2(n12346), .A(n12345), .ZN(n12347) );
  NAND2_X1 U8093 ( .A1(n8912), .A2(n8914), .ZN(n7292) );
  INV_X1 U8094 ( .A(n6791), .ZN(n6790) );
  INV_X1 U8095 ( .A(n14070), .ZN(n6795) );
  NOR2_X1 U8096 ( .A1(n14071), .A2(n6793), .ZN(n6792) );
  INV_X1 U8097 ( .A(n7434), .ZN(n6793) );
  INV_X1 U8098 ( .A(n12377), .ZN(n6797) );
  NAND2_X1 U8099 ( .A1(n8951), .A2(n8949), .ZN(n7303) );
  NAND2_X1 U8100 ( .A1(n12387), .A2(n12389), .ZN(n7321) );
  NAND2_X1 U8101 ( .A1(n8991), .A2(n8990), .ZN(n9008) );
  AND2_X1 U8102 ( .A1(n12405), .A2(n6803), .ZN(n6802) );
  NAND2_X1 U8103 ( .A1(n12400), .A2(n12402), .ZN(n7317) );
  NAND2_X1 U8104 ( .A1(n6800), .A2(n12410), .ZN(n6799) );
  INV_X1 U8105 ( .A(n6802), .ZN(n6800) );
  NAND2_X1 U8106 ( .A1(n12403), .A2(n12406), .ZN(n6801) );
  INV_X1 U8107 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7024) );
  INV_X1 U8108 ( .A(n8402), .ZN(n7054) );
  INV_X1 U8109 ( .A(n7047), .ZN(n7046) );
  OAI21_X1 U8110 ( .B1(n7049), .B2(n7048), .A(n7447), .ZN(n7047) );
  INV_X1 U8111 ( .A(n8357), .ZN(n7048) );
  NOR2_X1 U8112 ( .A1(n14410), .A2(n14409), .ZN(n14411) );
  NAND2_X1 U8113 ( .A1(n12598), .A2(n12542), .ZN(n12545) );
  INV_X1 U8114 ( .A(n12523), .ZN(n6750) );
  NAND2_X1 U8115 ( .A1(n12858), .A2(n12707), .ZN(n8136) );
  OAI21_X1 U8116 ( .B1(n13141), .B2(P3_REG2_REG_1__SCAN_IN), .A(n6688), .ZN(
        n10016) );
  NAND2_X1 U8117 ( .A1(n13141), .A2(n15090), .ZN(n6688) );
  AOI21_X1 U8118 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n10251), .A(n12723), .ZN(
        n10280) );
  NAND2_X1 U8119 ( .A1(n12755), .A2(n12754), .ZN(n12756) );
  OAI21_X1 U8120 ( .B1(n12815), .B2(n7104), .A(n12831), .ZN(n7103) );
  OR2_X1 U8121 ( .A1(n7941), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n7961) );
  OR2_X1 U8122 ( .A1(n12575), .A2(n12877), .ZN(n8298) );
  INV_X1 U8123 ( .A(n8266), .ZN(n7345) );
  OAI21_X1 U8124 ( .B1(n7816), .B2(n7345), .A(n8270), .ZN(n7344) );
  NAND2_X1 U8125 ( .A1(n7686), .A2(n7685), .ZN(n7706) );
  INV_X1 U8126 ( .A(n7687), .ZN(n7686) );
  AND2_X1 U8127 ( .A1(n11442), .A2(n7986), .ZN(n7987) );
  NAND2_X1 U8128 ( .A1(n7972), .A2(n12721), .ZN(n8174) );
  INV_X1 U8129 ( .A(n10818), .ZN(n7960) );
  INV_X1 U8130 ( .A(n7873), .ZN(n6954) );
  OAI21_X1 U8131 ( .B1(n6955), .B2(n6954), .A(P2_DATAO_REG_24__SCAN_IN), .ZN(
        n6953) );
  OR2_X1 U8132 ( .A1(n7874), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n7893) );
  NAND2_X1 U8133 ( .A1(n7859), .A2(n6955), .ZN(n6950) );
  INV_X1 U8134 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n8373) );
  INV_X1 U8135 ( .A(n6930), .ZN(n6929) );
  OAI21_X1 U8136 ( .B1(n7746), .B2(n6931), .A(n7761), .ZN(n6930) );
  INV_X1 U8137 ( .A(n7748), .ZN(n6931) );
  INV_X1 U8138 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8317) );
  XNOR2_X1 U8139 ( .A(n6696), .B(n13222), .ZN(n13163) );
  NOR2_X1 U8140 ( .A1(n6713), .A2(n13305), .ZN(n6712) );
  INV_X1 U8141 ( .A(n6716), .ZN(n6713) );
  INV_X1 U8142 ( .A(n13275), .ZN(n6734) );
  INV_X1 U8143 ( .A(n7007), .ZN(n7006) );
  OAI21_X1 U8144 ( .B1(n11861), .B2(n6831), .A(n6830), .ZN(n13376) );
  OR2_X1 U8145 ( .A1(n6832), .A2(n6607), .ZN(n6831) );
  NAND2_X1 U8146 ( .A1(n6833), .A2(n11862), .ZN(n6830) );
  AND2_X1 U8147 ( .A1(n14909), .A2(n13368), .ZN(n13371) );
  NOR2_X1 U8148 ( .A1(n6764), .A2(n6761), .ZN(n6760) );
  INV_X1 U8149 ( .A(n6762), .ZN(n6761) );
  INV_X1 U8150 ( .A(n11965), .ZN(n7236) );
  NOR2_X1 U8151 ( .A1(n13724), .A2(n13539), .ZN(n6769) );
  NOR2_X1 U8152 ( .A1(n11793), .A2(n11976), .ZN(n11993) );
  NOR2_X1 U8153 ( .A1(n11310), .A2(n14813), .ZN(n6772) );
  AND2_X1 U8154 ( .A1(n6772), .A2(n6771), .ZN(n6770) );
  AND2_X1 U8155 ( .A1(n11106), .A2(n14968), .ZN(n11163) );
  AND2_X1 U8156 ( .A1(n8660), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U8157 ( .A1(n13624), .A2(n11949), .ZN(n13604) );
  NOR2_X1 U8158 ( .A1(n10961), .A2(n11100), .ZN(n11106) );
  OR2_X1 U8159 ( .A1(n10778), .A2(n10954), .ZN(n10961) );
  INV_X1 U8160 ( .A(n9956), .ZN(n9891) );
  NOR2_X1 U8161 ( .A1(n8709), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8727) );
  OR2_X1 U8162 ( .A1(n8687), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8709) );
  AND2_X1 U8163 ( .A1(n8643), .A2(n8642), .ZN(n8670) );
  NOR2_X1 U8164 ( .A1(n8619), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8643) );
  INV_X1 U8165 ( .A(n11524), .ZN(n7223) );
  NAND2_X1 U8166 ( .A1(n11736), .A2(n6784), .ZN(n11737) );
  OR2_X1 U8167 ( .A1(n11745), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6784) );
  INV_X1 U8168 ( .A(n14080), .ZN(n7161) );
  AND2_X1 U8169 ( .A1(n11232), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n11491) );
  NOR2_X1 U8170 ( .A1(n11221), .A2(n11220), .ZN(n11232) );
  INV_X1 U8171 ( .A(n7144), .ZN(n7143) );
  INV_X1 U8172 ( .A(n10980), .ZN(n7145) );
  NAND2_X1 U8173 ( .A1(n14643), .A2(n6872), .ZN(n6871) );
  INV_X1 U8174 ( .A(n13969), .ZN(n11350) );
  INV_X1 U8175 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10608) );
  INV_X1 U8176 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U8177 ( .A1(n6674), .A2(n12292), .ZN(n10770) );
  INV_X1 U8178 ( .A(n10771), .ZN(n6674) );
  NAND2_X1 U8179 ( .A1(n12101), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7148) );
  AND2_X1 U8180 ( .A1(n13977), .A2(n10475), .ZN(n12261) );
  OR2_X1 U8181 ( .A1(n9031), .A2(n12252), .ZN(n8407) );
  AOI21_X1 U8182 ( .B1(n8391), .B2(n7028), .A(n7027), .ZN(n7026) );
  INV_X1 U8183 ( .A(n8388), .ZN(n7028) );
  INV_X1 U8184 ( .A(n8392), .ZN(n7027) );
  AOI21_X1 U8185 ( .B1(n6499), .B2(n7035), .A(n6592), .ZN(n7031) );
  AND2_X1 U8186 ( .A1(n7033), .A2(n8381), .ZN(n7032) );
  NAND2_X1 U8187 ( .A1(n7034), .A2(n8380), .ZN(n7033) );
  INV_X1 U8188 ( .A(n8377), .ZN(n7034) );
  NAND2_X1 U8189 ( .A1(n8374), .A2(n9678), .ZN(n8377) );
  NAND2_X1 U8190 ( .A1(n6700), .A2(n6699), .ZN(n8830) );
  AOI22_X1 U8191 ( .A1(n6705), .A2(n6706), .B1(n6707), .B2(n8366), .ZN(n6699)
         );
  INV_X1 U8192 ( .A(n6709), .ZN(n6706) );
  NOR2_X1 U8193 ( .A1(n9346), .A2(n9345), .ZN(n9446) );
  AOI21_X1 U8194 ( .B1(n7039), .B2(n7040), .A(n6557), .ZN(n7037) );
  INV_X1 U8195 ( .A(n8345), .ZN(n7040) );
  NAND2_X1 U8196 ( .A1(n6720), .A2(n6721), .ZN(n8641) );
  AOI21_X1 U8197 ( .B1(n8337), .B2(n6722), .A(n6559), .ZN(n6721) );
  INV_X1 U8198 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14407) );
  XNOR2_X1 U8199 ( .A(n14411), .B(n6865), .ZN(n14455) );
  NOR2_X1 U8200 ( .A1(n14421), .A2(n14420), .ZN(n14454) );
  NOR2_X1 U8201 ( .A1(n14481), .A2(n14482), .ZN(n14420) );
  INV_X2 U8202 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n15238) );
  NAND2_X1 U8203 ( .A1(n14496), .A2(n14426), .ZN(n14451) );
  NAND2_X1 U8204 ( .A1(n7801), .A2(n7800), .ZN(n7811) );
  AOI21_X1 U8205 ( .B1(n12578), .B2(n12563), .A(n12566), .ZN(n7073) );
  INV_X1 U8206 ( .A(n7073), .ZN(n7070) );
  XNOR2_X1 U8207 ( .A(n11463), .B(n10532), .ZN(n11055) );
  AND2_X1 U8208 ( .A1(n12609), .A2(n12555), .ZN(n12639) );
  NAND2_X1 U8209 ( .A1(n7880), .A2(n7879), .ZN(n7900) );
  INV_X1 U8210 ( .A(n7881), .ZN(n7880) );
  INV_X1 U8211 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n10409) );
  AOI21_X1 U8212 ( .B1(n7065), .B2(n12537), .A(n6524), .ZN(n7064) );
  INV_X1 U8213 ( .A(n7075), .ZN(n7074) );
  NAND2_X1 U8214 ( .A1(n11060), .A2(n7077), .ZN(n6744) );
  OAI21_X1 U8215 ( .B1(n11374), .B2(n7076), .A(n11507), .ZN(n7075) );
  OR2_X1 U8216 ( .A1(n7670), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7687) );
  INV_X1 U8217 ( .A(n6990), .ZN(n8306) );
  NOR2_X1 U8218 ( .A1(n8157), .A2(n6989), .ZN(n6988) );
  AND2_X1 U8219 ( .A1(n8114), .A2(n8113), .ZN(n12852) );
  AND2_X1 U8220 ( .A1(n8114), .A2(n8094), .ZN(n8129) );
  CLKBUF_X1 U8221 ( .A(P3_IR_REG_1__SCAN_IN), .Z(n10138) );
  AND2_X1 U8222 ( .A1(n10148), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10149) );
  AND2_X1 U8223 ( .A1(n10151), .A2(n6653), .ZN(n6672) );
  NAND2_X1 U8224 ( .A1(n10182), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10181) );
  AND2_X1 U8225 ( .A1(n6652), .A2(n10145), .ZN(n10185) );
  NAND2_X1 U8226 ( .A1(n6654), .A2(n6653), .ZN(n6652) );
  NAND2_X1 U8227 ( .A1(n10185), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10184) );
  AND3_X1 U8228 ( .A1(n6919), .A2(P3_REG1_REG_5__SCAN_IN), .A3(n6918), .ZN(
        n12739) );
  AOI21_X1 U8229 ( .B1(n12725), .B2(n6504), .A(n12724), .ZN(n12723) );
  OR2_X1 U8230 ( .A1(n10273), .A2(n6531), .ZN(n6915) );
  INV_X1 U8231 ( .A(n6924), .ZN(n11255) );
  NOR2_X1 U8232 ( .A1(n11545), .A2(n11546), .ZN(n11549) );
  OR3_X1 U8233 ( .A1(n14997), .A2(n11931), .A3(n11930), .ZN(n12755) );
  NOR2_X1 U8234 ( .A1(n14998), .A2(n14999), .ZN(n14997) );
  INV_X1 U8235 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n12694) );
  XNOR2_X1 U8236 ( .A(n12756), .B(n6687), .ZN(n14554) );
  INV_X1 U8237 ( .A(n7103), .ZN(n7102) );
  NOR2_X1 U8238 ( .A1(n7104), .A2(n7101), .ZN(n7096) );
  OAI21_X1 U8239 ( .B1(n7103), .B2(n7099), .A(n7098), .ZN(n7097) );
  NOR2_X1 U8240 ( .A1(n12818), .A2(n12838), .ZN(n7099) );
  NAND2_X1 U8241 ( .A1(n7103), .A2(n7101), .ZN(n7098) );
  INV_X1 U8242 ( .A(n6965), .ZN(n6960) );
  OR2_X1 U8243 ( .A1(n12852), .A2(n12851), .ZN(n14563) );
  AOI21_X1 U8244 ( .B1(n6486), .B2(n12881), .A(n6553), .ZN(n6906) );
  NAND2_X1 U8245 ( .A1(n6907), .A2(n6486), .ZN(n8088) );
  NAND2_X1 U8246 ( .A1(n8298), .A2(n8078), .ZN(n12568) );
  NOR2_X1 U8247 ( .A1(n12572), .A2(n12962), .ZN(n6640) );
  AND2_X1 U8248 ( .A1(n8164), .A2(n8163), .ZN(n12946) );
  AND3_X1 U8249 ( .A1(n7815), .A2(n7814), .A3(n7813), .ZN(n12963) );
  NAND2_X1 U8250 ( .A1(n7817), .A2(n7816), .ZN(n12979) );
  NAND2_X1 U8251 ( .A1(n6503), .A2(n6881), .ZN(n6880) );
  INV_X1 U8252 ( .A(n6886), .ZN(n6881) );
  INV_X1 U8253 ( .A(n12993), .ZN(n8004) );
  NAND2_X1 U8254 ( .A1(n8000), .A2(n7999), .ZN(n13020) );
  AND4_X1 U8255 ( .A1(n7711), .A2(n7710), .A3(n7709), .A4(n7708), .ZN(n11677)
         );
  OR2_X1 U8256 ( .A1(n7647), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7670) );
  NAND2_X1 U8257 ( .A1(n7630), .A2(n10409), .ZN(n7647) );
  INV_X1 U8258 ( .A(n7631), .ZN(n7630) );
  AOI21_X1 U8259 ( .B1(n7334), .B2(n7336), .A(n7331), .ZN(n7330) );
  INV_X1 U8260 ( .A(n8201), .ZN(n7331) );
  OR2_X1 U8261 ( .A1(n7614), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n7631) );
  AND2_X1 U8262 ( .A1(n11131), .A2(n7985), .ZN(n11459) );
  NAND2_X1 U8263 ( .A1(n7485), .A2(n10242), .ZN(n7614) );
  INV_X1 U8264 ( .A(n7599), .ZN(n7485) );
  NAND2_X1 U8265 ( .A1(n7484), .A2(n10225), .ZN(n7597) );
  NAND2_X1 U8266 ( .A1(n10569), .A2(n10156), .ZN(n7580) );
  AND4_X1 U8267 ( .A1(n7556), .A2(n7555), .A3(n7554), .A4(n7553), .ZN(n10538)
         );
  NAND2_X1 U8268 ( .A1(n7976), .A2(n7975), .ZN(n10320) );
  CLKBUF_X1 U8269 ( .A(n10031), .Z(n10310) );
  CLKBUF_X1 U8270 ( .A(n7971), .Z(n10560) );
  CLKBUF_X1 U8271 ( .A(n8143), .Z(n10303) );
  CLKBUF_X1 U8272 ( .A(n8145), .Z(n10304) );
  NAND2_X1 U8273 ( .A1(n8120), .A2(n8119), .ZN(n14566) );
  INV_X1 U8274 ( .A(n14563), .ZN(n14565) );
  NAND2_X1 U8275 ( .A1(n11144), .A2(n11145), .ZN(n7333) );
  AND2_X1 U8276 ( .A1(n6748), .A2(n6747), .ZN(n8034) );
  NAND2_X1 U8277 ( .A1(n6967), .A2(n6974), .ZN(n6966) );
  INV_X1 U8278 ( .A(n6972), .ZN(n6967) );
  NOR2_X1 U8279 ( .A1(n6969), .A2(n6974), .ZN(n6965) );
  OR2_X1 U8280 ( .A1(n6973), .A2(n6616), .ZN(n6972) );
  INV_X1 U8281 ( .A(n8121), .ZN(n6973) );
  NAND2_X1 U8282 ( .A1(n12432), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6975) );
  NAND2_X1 U8283 ( .A1(n6971), .A2(n8121), .ZN(n6970) );
  INV_X1 U8284 ( .A(n8115), .ZN(n6971) );
  AOI21_X1 U8285 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n15230), .A(n7937), .ZN(
        n8081) );
  NOR2_X1 U8286 ( .A1(n7936), .A2(n7935), .ZN(n7937) );
  AOI21_X1 U8287 ( .B1(n6937), .B2(n6936), .A(n6935), .ZN(n7936) );
  AND2_X1 U8288 ( .A1(n12184), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6935) );
  INV_X1 U8289 ( .A(n8015), .ZN(n8017) );
  XNOR2_X1 U8290 ( .A(n8039), .B(n8038), .ZN(n10000) );
  NOR2_X1 U8291 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_20__SCAN_IN), .ZN(
        n7466) );
  CLKBUF_X1 U8292 ( .A(n8013), .Z(n7953) );
  AOI21_X1 U8293 ( .B1(n7781), .B2(n7082), .A(n7079), .ZN(n7078) );
  NAND2_X1 U8294 ( .A1(n7081), .A2(n7080), .ZN(n7079) );
  AND2_X1 U8295 ( .A1(n6529), .A2(n7464), .ZN(n6661) );
  AOI21_X1 U8296 ( .B1(n6978), .B2(n6979), .A(n6596), .ZN(n6977) );
  NAND2_X1 U8297 ( .A1(n6941), .A2(n6939), .ZN(n7638) );
  AOI21_X1 U8298 ( .B1(n6563), .B2(n6943), .A(n6940), .ZN(n6939) );
  NOR2_X1 U8299 ( .A1(n9279), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n6940) );
  XNOR2_X1 U8300 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7570) );
  NAND2_X1 U8301 ( .A1(n6925), .A2(n7505), .ZN(n7558) );
  NAND2_X1 U8302 ( .A1(n7526), .A2(n7504), .ZN(n6925) );
  NAND2_X1 U8303 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7536) );
  XNOR2_X1 U8304 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7533) );
  AND2_X1 U8305 ( .A1(n8536), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7548) );
  INV_X1 U8306 ( .A(n11197), .ZN(n7005) );
  NOR2_X1 U8307 ( .A1(n8931), .A2(n13237), .ZN(n8952) );
  OR2_X1 U8308 ( .A1(n8840), .A2(n14875), .ZN(n8842) );
  OR2_X1 U8309 ( .A1(n10505), .A2(n10504), .ZN(n10430) );
  NAND2_X1 U8310 ( .A1(n6656), .A2(n6552), .ZN(n13289) );
  INV_X1 U8311 ( .A(n13290), .ZN(n6656) );
  NOR2_X1 U8312 ( .A1(n7018), .A2(n14809), .ZN(n7017) );
  INV_X1 U8313 ( .A(n11613), .ZN(n7018) );
  NAND2_X1 U8314 ( .A1(n6526), .A2(n13172), .ZN(n6716) );
  NAND2_X1 U8315 ( .A1(n7363), .A2(n10060), .ZN(n9827) );
  XNOR2_X1 U8316 ( .A(n9796), .B(n9812), .ZN(n10113) );
  NOR2_X1 U8317 ( .A1(n14920), .A2(n9788), .ZN(n9809) );
  NAND2_X1 U8318 ( .A1(n6485), .A2(n13400), .ZN(n9751) );
  OR2_X1 U8319 ( .A1(n7277), .A2(n9068), .ZN(n7276) );
  NAND4_X1 U8320 ( .A1(n8553), .A2(n8552), .A3(n8551), .A4(n8550), .ZN(n9109)
         );
  NOR2_X1 U8321 ( .A1(n9547), .A2(n6841), .ZN(n9549) );
  AND2_X1 U8322 ( .A1(n9550), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6841) );
  NOR2_X1 U8323 ( .A1(n9549), .A2(n9548), .ZN(n9564) );
  NOR2_X1 U8324 ( .A1(n11861), .A2(n6607), .ZN(n6834) );
  INV_X1 U8325 ( .A(n14878), .ZN(n6833) );
  AND2_X1 U8326 ( .A1(n13384), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n13394) );
  AND2_X1 U8327 ( .A1(n13371), .A2(n13370), .ZN(n13391) );
  NOR2_X1 U8328 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13372), .ZN(n13390) );
  AOI21_X1 U8329 ( .B1(n13807), .B2(n9061), .A(n7444), .ZN(n11994) );
  AOI21_X1 U8330 ( .B1(n7383), .B2(n7387), .A(n6555), .ZN(n7381) );
  NAND2_X1 U8331 ( .A1(n11968), .A2(n9102), .ZN(n13415) );
  OR2_X1 U8332 ( .A1(n9050), .A2(n13227), .ZN(n11995) );
  NAND2_X1 U8333 ( .A1(n7265), .A2(n13433), .ZN(n7264) );
  NAND2_X1 U8334 ( .A1(n13435), .A2(n13434), .ZN(n7265) );
  NOR2_X1 U8335 ( .A1(n11988), .A2(n7390), .ZN(n7389) );
  INV_X1 U8336 ( .A(n11987), .ZN(n7390) );
  OAI21_X1 U8337 ( .B1(n13482), .B2(n7238), .A(n7235), .ZN(n13456) );
  AOI21_X1 U8338 ( .B1(n7239), .B2(n7237), .A(n7236), .ZN(n7235) );
  INV_X1 U8339 ( .A(n7239), .ZN(n7238) );
  INV_X1 U8340 ( .A(n11964), .ZN(n7237) );
  NAND2_X1 U8341 ( .A1(n13456), .A2(n13457), .ZN(n13455) );
  AND2_X1 U8342 ( .A1(n13490), .A2(n6762), .ZN(n13450) );
  NAND2_X1 U8343 ( .A1(n13490), .A2(n13773), .ZN(n13472) );
  NAND2_X1 U8344 ( .A1(n13554), .A2(n6765), .ZN(n13505) );
  AND2_X1 U8345 ( .A1(n6767), .A2(n6766), .ZN(n6765) );
  NAND2_X1 U8346 ( .A1(n13554), .A2(n6767), .ZN(n13522) );
  OR2_X1 U8347 ( .A1(n11347), .A2(n9003), .ZN(n8961) );
  NAND2_X1 U8348 ( .A1(n13554), .A2(n11983), .ZN(n13555) );
  NAND2_X1 U8349 ( .A1(n7244), .A2(n7248), .ZN(n7242) );
  INV_X1 U8350 ( .A(n11953), .ZN(n13549) );
  INV_X1 U8351 ( .A(n7249), .ZN(n7248) );
  AOI21_X1 U8352 ( .B1(n7249), .B2(n7247), .A(n6544), .ZN(n7246) );
  INV_X1 U8353 ( .A(n11949), .ZN(n7247) );
  NAND2_X1 U8354 ( .A1(n13604), .A2(n11950), .ZN(n13574) );
  OR2_X1 U8355 ( .A1(n6517), .A2(n7409), .ZN(n7406) );
  NOR2_X1 U8356 ( .A1(n11656), .A2(n7410), .ZN(n7409) );
  NAND3_X1 U8357 ( .A1(n11788), .A2(n6770), .A3(n11163), .ZN(n11793) );
  NAND2_X1 U8358 ( .A1(n11163), .A2(n6772), .ZN(n11567) );
  AOI21_X1 U8359 ( .B1(n7229), .B2(n7231), .A(n11098), .ZN(n7228) );
  AND2_X1 U8360 ( .A1(n11155), .A2(n9107), .ZN(n11157) );
  OAI21_X1 U8361 ( .B1(n10783), .B2(n7231), .A(n7229), .ZN(n11099) );
  NOR2_X1 U8362 ( .A1(n10738), .A2(n7413), .ZN(n7412) );
  INV_X1 U8363 ( .A(n10731), .ZN(n7413) );
  NAND2_X1 U8364 ( .A1(n10783), .A2(n10736), .ZN(n7233) );
  INV_X1 U8365 ( .A(n10730), .ZN(n10782) );
  NOR2_X1 U8366 ( .A1(n10377), .A2(n14938), .ZN(n10779) );
  NOR2_X1 U8367 ( .A1(n10382), .A2(n10375), .ZN(n7379) );
  AND2_X1 U8368 ( .A1(n7378), .A2(n7376), .ZN(n7375) );
  OR2_X1 U8369 ( .A1(n14932), .A2(n13355), .ZN(n7378) );
  NAND2_X1 U8370 ( .A1(n10734), .A2(n9110), .ZN(n10726) );
  NAND2_X1 U8371 ( .A1(n10363), .A2(n10362), .ZN(n10381) );
  XNOR2_X1 U8372 ( .A(n10502), .B(n7226), .ZN(n9956) );
  INV_X1 U8373 ( .A(n9827), .ZN(n10112) );
  CLKBUF_X1 U8374 ( .A(n9712), .Z(n6618) );
  AND2_X1 U8375 ( .A1(n13680), .A2(n14939), .ZN(n6632) );
  NAND2_X1 U8376 ( .A1(n7396), .A2(n7403), .ZN(n13531) );
  OR2_X1 U8377 ( .A1(n13550), .A2(n11984), .ZN(n7396) );
  AND2_X1 U8378 ( .A1(n9727), .A2(n9742), .ZN(n14917) );
  OR2_X1 U8379 ( .A1(n12102), .A2(n8957), .ZN(n8959) );
  INV_X1 U8380 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n7281) );
  AND2_X1 U8381 ( .A1(n8433), .A2(n8427), .ZN(n7288) );
  INV_X1 U8382 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8429) );
  INV_X1 U8383 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8536) );
  OR2_X1 U8384 ( .A1(n9258), .A2(n12141), .ZN(n9757) );
  OR2_X1 U8385 ( .A1(n10609), .A2(n10608), .ZN(n10624) );
  OR2_X1 U8386 ( .A1(n10983), .A2(n10982), .ZN(n11221) );
  AND2_X1 U8387 ( .A1(n12182), .A2(n12180), .ZN(n13865) );
  NAND2_X1 U8388 ( .A1(n11491), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11634) );
  OR2_X1 U8389 ( .A1(n11634), .A2(n11633), .ZN(n11810) );
  NAND2_X1 U8390 ( .A1(n6494), .A2(n7210), .ZN(n7208) );
  CLKBUF_X1 U8391 ( .A(n11425), .Z(n11421) );
  INV_X1 U8392 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10843) );
  OR2_X1 U8393 ( .A1(n10624), .A2(n10623), .ZN(n10844) );
  OR2_X1 U8394 ( .A1(n12069), .A2(n13907), .ZN(n12085) );
  OR2_X1 U8395 ( .A1(n12045), .A2(n12044), .ZN(n12069) );
  NAND2_X1 U8396 ( .A1(n7196), .A2(n7203), .ZN(n7195) );
  INV_X1 U8397 ( .A(n7198), .ZN(n7196) );
  AOI21_X1 U8398 ( .B1(n7201), .B2(n7199), .A(n12100), .ZN(n7198) );
  INV_X1 U8399 ( .A(n7201), .ZN(n7200) );
  NOR2_X1 U8400 ( .A1(n10844), .A2(n10843), .ZN(n10901) );
  INV_X1 U8401 ( .A(n12165), .ZN(n12187) );
  INV_X1 U8402 ( .A(n9937), .ZN(n12092) );
  AND4_X1 U8403 ( .A1(n11237), .A2(n11236), .A3(n11235), .A4(n11234), .ZN(
        n12010) );
  AND2_X1 U8404 ( .A1(n9414), .A2(n6579), .ZN(n9415) );
  NOR2_X1 U8405 ( .A1(n10331), .A2(n6779), .ZN(n10334) );
  AND2_X1 U8406 ( .A1(n10885), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6779) );
  NAND2_X1 U8407 ( .A1(n10334), .A2(n10333), .ZN(n10545) );
  NAND2_X1 U8408 ( .A1(n10545), .A2(n6778), .ZN(n10546) );
  OR2_X1 U8409 ( .A1(n10977), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8410 ( .A1(n10546), .A2(n10547), .ZN(n11000) );
  XNOR2_X1 U8411 ( .A(n11737), .B(n14682), .ZN(n14679) );
  NOR2_X1 U8412 ( .A1(n13978), .A2(n6782), .ZN(n13982) );
  AND2_X1 U8413 ( .A1(n13989), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6782) );
  NOR2_X1 U8414 ( .A1(n7124), .A2(n7129), .ZN(n7123) );
  INV_X1 U8415 ( .A(n7127), .ZN(n7124) );
  NAND2_X1 U8416 ( .A1(n6565), .A2(n7127), .ZN(n7122) );
  NAND2_X1 U8417 ( .A1(n14152), .A2(n7128), .ZN(n7125) );
  NAND2_X1 U8418 ( .A1(n14091), .A2(n14090), .ZN(n7174) );
  AND2_X1 U8419 ( .A1(n14320), .A2(n14087), .ZN(n6626) );
  NAND2_X1 U8420 ( .A1(n7138), .A2(n7137), .ZN(n7136) );
  INV_X1 U8421 ( .A(n14055), .ZN(n7137) );
  NAND2_X1 U8422 ( .A1(n14207), .A2(n14206), .ZN(n14205) );
  AOI21_X1 U8423 ( .B1(n7178), .B2(n11490), .A(n6550), .ZN(n7177) );
  NAND2_X1 U8424 ( .A1(n11489), .A2(n7178), .ZN(n6637) );
  OR2_X1 U8425 ( .A1(n12329), .A2(n12339), .ZN(n6870) );
  NAND2_X1 U8426 ( .A1(n11483), .A2(n14636), .ZN(n11824) );
  AOI21_X1 U8427 ( .B1(n7157), .B2(n7159), .A(n6548), .ZN(n7155) );
  INV_X1 U8428 ( .A(n13917), .ZN(n14064) );
  NOR2_X1 U8429 ( .A1(n10897), .A2(n6871), .ZN(n11277) );
  NOR2_X1 U8430 ( .A1(n10897), .A2(n14778), .ZN(n10993) );
  NAND2_X1 U8431 ( .A1(n10619), .A2(n10618), .ZN(n14708) );
  INV_X1 U8432 ( .A(n7135), .ZN(n7134) );
  NOR2_X1 U8433 ( .A1(n9939), .A2(n9938), .ZN(n10596) );
  AND2_X1 U8434 ( .A1(n7166), .A2(n10591), .ZN(n7163) );
  NAND2_X1 U8435 ( .A1(n7150), .A2(n9645), .ZN(n10873) );
  NAND2_X1 U8436 ( .A1(n9644), .A2(n7147), .ZN(n7150) );
  OR2_X1 U8437 ( .A1(n9644), .A2(n9643), .ZN(n9645) );
  OAI21_X1 U8438 ( .B1(n9641), .B2(n9249), .A(n7148), .ZN(n7147) );
  NAND2_X1 U8439 ( .A1(n12265), .A2(n12259), .ZN(n9880) );
  CLKBUF_X1 U8440 ( .A(n10477), .Z(n12471) );
  OR2_X1 U8441 ( .A1(n10487), .A2(n12514), .ZN(n14102) );
  NAND2_X1 U8442 ( .A1(n12186), .A2(n12185), .ZN(n14315) );
  INV_X1 U8443 ( .A(n14735), .ZN(n14780) );
  INV_X1 U8444 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7311) );
  XNOR2_X1 U8445 ( .A(n8503), .B(n8502), .ZN(n13796) );
  OAI21_X1 U8446 ( .B1(n8500), .B2(n8499), .A(n8498), .ZN(n8503) );
  XNOR2_X1 U8447 ( .A(n8500), .B(n8419), .ZN(n12431) );
  XNOR2_X1 U8448 ( .A(n8496), .B(n8495), .ZN(n13807) );
  XNOR2_X1 U8449 ( .A(n9194), .B(n9193), .ZN(n9201) );
  NAND2_X1 U8450 ( .A1(n9192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9194) );
  NAND2_X1 U8451 ( .A1(n9002), .A2(n8402), .ZN(n8527) );
  NAND2_X1 U8452 ( .A1(n8981), .A2(n8399), .ZN(n9000) );
  NAND2_X1 U8453 ( .A1(n8959), .A2(n8396), .ZN(n8979) );
  NAND2_X1 U8454 ( .A1(n8979), .A2(n8978), .ZN(n8981) );
  NAND2_X1 U8455 ( .A1(n8394), .A2(n8396), .ZN(n12102) );
  OR2_X1 U8456 ( .A1(n8393), .A2(SI_22_), .ZN(n8394) );
  INV_X1 U8457 ( .A(n6805), .ZN(n6804) );
  OR2_X1 U8458 ( .A1(n9183), .A2(n6809), .ZN(n6808) );
  XNOR2_X1 U8459 ( .A(n8944), .B(n8939), .ZN(n12065) );
  XNOR2_X1 U8460 ( .A(n8908), .B(n8907), .ZN(n12039) );
  NAND2_X1 U8461 ( .A1(n7041), .A2(n8367), .ZN(n8848) );
  NAND2_X1 U8462 ( .A1(n6704), .A2(n6709), .ZN(n8367) );
  NAND2_X1 U8463 ( .A1(n6698), .A2(n6707), .ZN(n7041) );
  NAND2_X1 U8464 ( .A1(n7045), .A2(n8357), .ZN(n8764) );
  NAND2_X1 U8465 ( .A1(n8353), .A2(n7049), .ZN(n7045) );
  NAND2_X1 U8466 ( .A1(n8353), .A2(n8352), .ZN(n8749) );
  NAND2_X1 U8467 ( .A1(n7038), .A2(n8345), .ZN(n8686) );
  NAND2_X1 U8468 ( .A1(n8669), .A2(n8343), .ZN(n7038) );
  NAND2_X1 U8469 ( .A1(n6723), .A2(n8336), .ZN(n8618) );
  NAND2_X1 U8470 ( .A1(n8605), .A2(n8334), .ZN(n6723) );
  NAND2_X1 U8471 ( .A1(n8327), .A2(n8326), .ZN(n8587) );
  INV_X1 U8472 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14461) );
  NAND2_X1 U8473 ( .A1(n15309), .A2(n15310), .ZN(n14463) );
  INV_X1 U8474 ( .A(n14406), .ZN(n14458) );
  XNOR2_X1 U8475 ( .A(n14455), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14456) );
  INV_X1 U8476 ( .A(n6850), .ZN(n14475) );
  OAI21_X1 U8477 ( .B1(n15299), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6545), .ZN(
        n6850) );
  NOR2_X1 U8478 ( .A1(n14417), .A2(n14416), .ZN(n14477) );
  NOR2_X1 U8479 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14471), .ZN(n14416) );
  INV_X1 U8480 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14476) );
  NAND2_X1 U8481 ( .A1(n6851), .A2(n14484), .ZN(n14485) );
  NAND2_X1 U8482 ( .A1(n15302), .A2(n15303), .ZN(n6851) );
  OR2_X1 U8483 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14425), .ZN(n14496) );
  INV_X1 U8484 ( .A(n14663), .ZN(n6863) );
  NAND2_X1 U8485 ( .A1(n6854), .A2(n6853), .ZN(n14534) );
  NAND2_X1 U8486 ( .A1(n14529), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6853) );
  NAND2_X1 U8487 ( .A1(n6856), .A2(n14915), .ZN(n6855) );
  AND4_X1 U8488 ( .A1(n7620), .A2(n7619), .A3(n7618), .A4(n7617), .ZN(n11077)
         );
  INV_X1 U8489 ( .A(n12935), .ZN(n12586) );
  INV_X1 U8490 ( .A(n7057), .ZN(n7056) );
  AND4_X1 U8491 ( .A1(n7675), .A2(n7674), .A3(n7673), .A4(n7672), .ZN(n11588)
         );
  AOI21_X1 U8492 ( .B1(n12666), .B2(n12667), .A(n12537), .ZN(n12591) );
  XNOR2_X1 U8493 ( .A(n11055), .B(n11077), .ZN(n11267) );
  NAND2_X1 U8494 ( .A1(n10068), .A2(n10033), .ZN(n10038) );
  NAND2_X1 U8495 ( .A1(n6754), .A2(n7058), .ZN(n12600) );
  NAND2_X1 U8496 ( .A1(n7830), .A2(n7829), .ZN(n12605) );
  OR2_X1 U8497 ( .A1(n10573), .A2(n7828), .ZN(n7830) );
  INV_X1 U8498 ( .A(n12710), .ZN(n12625) );
  NAND2_X1 U8499 ( .A1(n12621), .A2(n12619), .ZN(n6740) );
  OAI21_X1 U8500 ( .B1(n12621), .B2(n12619), .A(n13024), .ZN(n6741) );
  NAND2_X1 U8501 ( .A1(n7766), .A2(n7765), .ZN(n13028) );
  NAND2_X1 U8502 ( .A1(n7059), .A2(n7064), .ZN(n12648) );
  NAND2_X1 U8503 ( .A1(n12666), .A2(n7065), .ZN(n7059) );
  NAND2_X1 U8504 ( .A1(n7810), .A2(n7809), .ZN(n12983) );
  CLKBUF_X1 U8505 ( .A(n11871), .Z(n6622) );
  NAND2_X1 U8506 ( .A1(n7848), .A2(n7847), .ZN(n12662) );
  CLKBUF_X1 U8507 ( .A(n12665), .Z(n12666) );
  AND2_X1 U8508 ( .A1(n7933), .A2(n7932), .ZN(n12891) );
  NAND2_X1 U8509 ( .A1(n10041), .A2(n9919), .ZN(n12697) );
  NAND2_X1 U8510 ( .A1(n12686), .A2(n12687), .ZN(n12692) );
  INV_X1 U8511 ( .A(n12672), .ZN(n12700) );
  INV_X1 U8512 ( .A(n12891), .ZN(n12708) );
  NAND2_X1 U8513 ( .A1(n7906), .A2(n7905), .ZN(n12920) );
  NAND2_X1 U8514 ( .A1(n7840), .A2(n7839), .ZN(n12976) );
  INV_X1 U8515 ( .A(n12963), .ZN(n12990) );
  INV_X1 U8516 ( .A(n11588), .ZN(n12714) );
  OR2_X1 U8517 ( .A1(n9908), .A2(n9353), .ZN(n12718) );
  INV_X1 U8518 ( .A(n10538), .ZN(n12720) );
  NAND2_X1 U8519 ( .A1(n7563), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7541) );
  NOR2_X1 U8520 ( .A1(n10017), .A2(n10085), .ZN(n10211) );
  AOI21_X1 U8521 ( .B1(n10208), .B2(n10191), .A(n10190), .ZN(n10193) );
  XNOR2_X1 U8522 ( .A(n7094), .B(n6920), .ZN(n10218) );
  NAND2_X1 U8523 ( .A1(n10218), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n12725) );
  AND2_X1 U8524 ( .A1(n7609), .A2(n7701), .ZN(n12736) );
  AOI21_X1 U8525 ( .B1(n12730), .B2(n10259), .A(n10258), .ZN(n10297) );
  INV_X1 U8526 ( .A(n7090), .ZN(n10283) );
  INV_X1 U8527 ( .A(n6913), .ZN(n10406) );
  INV_X1 U8528 ( .A(n6915), .ZN(n10277) );
  INV_X1 U8529 ( .A(n7109), .ZN(n10683) );
  NAND2_X1 U8530 ( .A1(n7110), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7107) );
  INV_X1 U8531 ( .A(n10685), .ZN(n7110) );
  INV_X1 U8532 ( .A(n10684), .ZN(n7108) );
  NOR2_X1 U8533 ( .A1(n11540), .A2(n11541), .ZN(n11543) );
  NOR2_X1 U8534 ( .A1(n14988), .A2(n11924), .ZN(n12767) );
  NOR2_X1 U8535 ( .A1(n14546), .A2(n12770), .ZN(n12773) );
  NAND2_X1 U8536 ( .A1(n12817), .A2(n12818), .ZN(n12832) );
  AND2_X1 U8537 ( .A1(n7354), .A2(n8291), .ZN(n12882) );
  OAI21_X1 U8538 ( .B1(n6648), .B2(n12960), .A(n6645), .ZN(n12879) );
  NOR2_X1 U8539 ( .A1(n6647), .A2(n6646), .ZN(n6645) );
  AND2_X1 U8540 ( .A1(n7354), .A2(n12899), .ZN(n13041) );
  NAND2_X1 U8541 ( .A1(n6888), .A2(n6892), .ZN(n12933) );
  NAND2_X1 U8542 ( .A1(n13073), .A2(n8254), .ZN(n12994) );
  NAND2_X1 U8543 ( .A1(n7784), .A2(n7783), .ZN(n13074) );
  AND2_X1 U8544 ( .A1(n6903), .A2(n7996), .ZN(n11882) );
  NAND2_X1 U8545 ( .A1(n7995), .A2(n7994), .ZN(n11756) );
  AND2_X1 U8546 ( .A1(n7338), .A2(n7340), .ZN(n11680) );
  NAND2_X1 U8547 ( .A1(n11386), .A2(n8225), .ZN(n11601) );
  AND2_X1 U8548 ( .A1(n6899), .A2(n6896), .ZN(n11314) );
  OR2_X1 U8549 ( .A1(n9705), .A2(n9704), .ZN(n13031) );
  NAND2_X1 U8550 ( .A1(n10823), .A2(n7981), .ZN(n11146) );
  NAND2_X1 U8551 ( .A1(n7592), .A2(n7591), .ZN(n7593) );
  NAND2_X1 U8552 ( .A1(n9998), .A2(n9700), .ZN(n15025) );
  NAND2_X1 U8553 ( .A1(n9705), .A2(n15025), .ZN(n15030) );
  AND2_X1 U8554 ( .A1(n7897), .A2(n7896), .ZN(n13096) );
  AND2_X1 U8555 ( .A1(n7878), .A2(n7877), .ZN(n13100) );
  OR2_X1 U8556 ( .A1(n13050), .A2(n13049), .ZN(n13097) );
  INV_X1 U8557 ( .A(n12662), .ZN(n13108) );
  INV_X1 U8558 ( .A(n12605), .ZN(n13112) );
  AND2_X1 U8559 ( .A1(n7722), .A2(n7721), .ZN(n11874) );
  AND2_X1 U8560 ( .A1(n10000), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13131) );
  OAI22_X1 U8561 ( .A1(n6969), .A2(n6964), .B1(n6974), .B2(n6968), .ZN(n6963)
         );
  AND2_X1 U8562 ( .A1(n6972), .A2(n8123), .ZN(n6964) );
  INV_X1 U8563 ( .A(n7496), .ZN(n6879) );
  NOR2_X1 U8564 ( .A1(n8027), .A2(n8026), .ZN(n8028) );
  NAND2_X1 U8565 ( .A1(n8024), .A2(n8023), .ZN(n8029) );
  NOR2_X1 U8566 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n8026) );
  INV_X1 U8567 ( .A(n6937), .ZN(n7921) );
  NAND2_X1 U8568 ( .A1(n8015), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U8569 ( .A1(n7859), .A2(n7858), .ZN(n7871) );
  NAND2_X1 U8570 ( .A1(n7794), .A2(n7793), .ZN(n7808) );
  NAND2_X1 U8571 ( .A1(n6928), .A2(n7748), .ZN(n7762) );
  NAND2_X1 U8572 ( .A1(n7747), .A2(n7746), .ZN(n6928) );
  INV_X1 U8573 ( .A(SI_15_), .ZN(n9597) );
  INV_X1 U8574 ( .A(SI_13_), .ZN(n9327) );
  NAND2_X1 U8575 ( .A1(n6932), .A2(n7713), .ZN(n7714) );
  NAND2_X1 U8576 ( .A1(n6934), .A2(n7713), .ZN(n7698) );
  INV_X1 U8577 ( .A(SI_12_), .ZN(n9287) );
  XNOR2_X1 U8578 ( .A(n7682), .B(n7681), .ZN(n11921) );
  NAND2_X1 U8579 ( .A1(n6981), .A2(n6984), .ZN(n7678) );
  NAND2_X1 U8580 ( .A1(n6982), .A2(n6510), .ZN(n6981) );
  INV_X1 U8581 ( .A(SI_11_), .ZN(n9278) );
  NAND2_X1 U8582 ( .A1(n7659), .A2(n7680), .ZN(n11256) );
  OAI21_X1 U8583 ( .B1(n7654), .B2(n7653), .A(n6983), .ZN(n7663) );
  INV_X1 U8584 ( .A(n6985), .ZN(n6983) );
  XNOR2_X1 U8585 ( .A(n7625), .B(n7624), .ZN(n10407) );
  OAI21_X1 U8586 ( .B1(n7587), .B2(n6946), .A(n6943), .ZN(n7622) );
  NAND2_X1 U8587 ( .A1(n6949), .A2(n7510), .ZN(n7606) );
  NAND2_X1 U8588 ( .A1(n7587), .A2(n7586), .ZN(n6949) );
  NAND2_X1 U8589 ( .A1(n7457), .A2(n7456), .ZN(n7572) );
  INV_X1 U8590 ( .A(n13467), .ZN(n13437) );
  AND2_X1 U8591 ( .A1(n13322), .A2(n13189), .ZN(n13193) );
  NAND2_X1 U8592 ( .A1(n6724), .A2(n6726), .ZN(n13220) );
  NAND2_X1 U8593 ( .A1(n6999), .A2(n7004), .ZN(n11199) );
  NAND2_X1 U8594 ( .A1(n11037), .A2(n6511), .ZN(n6999) );
  OAI21_X1 U8595 ( .B1(n13242), .B2(n6727), .A(n6725), .ZN(n13226) );
  AOI21_X1 U8596 ( .B1(n6726), .B2(n6730), .A(n13219), .ZN(n6725) );
  INV_X1 U8597 ( .A(n10447), .ZN(n10110) );
  NAND2_X1 U8598 ( .A1(n13149), .A2(n6587), .ZN(n13256) );
  INV_X1 U8599 ( .A(n10429), .ZN(n7023) );
  AOI21_X1 U8600 ( .B1(n13148), .B2(n7011), .A(n13257), .ZN(n7010) );
  OR2_X1 U8601 ( .A1(n13146), .A2(n7013), .ZN(n7012) );
  NAND2_X1 U8602 ( .A1(n7003), .A2(n11032), .ZN(n11198) );
  NAND2_X1 U8603 ( .A1(n11037), .A2(n11031), .ZN(n7003) );
  OR2_X1 U8604 ( .A1(n14808), .A2(n13521), .ZN(n13329) );
  NAND2_X1 U8605 ( .A1(n14804), .A2(n14805), .ZN(n11619) );
  NAND2_X1 U8606 ( .A1(n11300), .A2(n11299), .ZN(n11614) );
  OR2_X1 U8607 ( .A1(n13282), .A2(n13631), .ZN(n14800) );
  OR2_X1 U8608 ( .A1(n13282), .A2(n13575), .ZN(n14801) );
  NAND2_X1 U8609 ( .A1(n10431), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14816) );
  NAND2_X1 U8610 ( .A1(n13275), .A2(n13156), .ZN(n13315) );
  NAND2_X1 U8611 ( .A1(n9033), .A2(n9032), .ZN(n13688) );
  NAND2_X1 U8612 ( .A1(n11898), .A2(n11897), .ZN(n13149) );
  XNOR2_X1 U8613 ( .A(n13148), .B(n13146), .ZN(n11898) );
  INV_X1 U8614 ( .A(n14808), .ZN(n13276) );
  NOR2_X1 U8615 ( .A1(n9457), .A2(n9456), .ZN(n9547) );
  NOR2_X1 U8616 ( .A1(n9521), .A2(n6842), .ZN(n9457) );
  AND2_X1 U8617 ( .A1(n9463), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6842) );
  NOR2_X1 U8618 ( .A1(n9849), .A2(n9848), .ZN(n10120) );
  NOR2_X1 U8619 ( .A1(n9846), .A2(n6844), .ZN(n9849) );
  AND2_X1 U8620 ( .A1(n9850), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6844) );
  NOR2_X1 U8621 ( .A1(n10120), .A2(n6843), .ZN(n10123) );
  AND2_X1 U8622 ( .A1(n10126), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U8623 ( .A1(n10123), .A2(n10122), .ZN(n10660) );
  NOR2_X1 U8624 ( .A1(n14856), .A2(n14855), .ZN(n14854) );
  NOR2_X1 U8625 ( .A1(n11394), .A2(n6846), .ZN(n14856) );
  AND2_X1 U8626 ( .A1(n11395), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6846) );
  NOR2_X1 U8627 ( .A1(n14854), .A2(n6845), .ZN(n14867) );
  AND2_X1 U8628 ( .A1(n14859), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U8629 ( .A1(n14867), .A2(n14868), .ZN(n14866) );
  NAND2_X1 U8630 ( .A1(n8796), .A2(n8451), .ZN(n8888) );
  XNOR2_X1 U8631 ( .A(n13410), .B(n13759), .ZN(n13403) );
  XNOR2_X1 U8632 ( .A(n11970), .B(n11969), .ZN(n11975) );
  OAI21_X1 U8633 ( .B1(n13471), .B2(n6513), .A(n11987), .ZN(n13449) );
  NAND2_X1 U8634 ( .A1(n7234), .A2(n7239), .ZN(n13464) );
  NAND2_X1 U8635 ( .A1(n7395), .A2(n7397), .ZN(n13519) );
  NAND2_X1 U8636 ( .A1(n13550), .A2(n7400), .ZN(n7395) );
  INV_X1 U8637 ( .A(n6693), .ZN(n13729) );
  NAND2_X1 U8638 ( .A1(n7366), .A2(n7367), .ZN(n13578) );
  AND2_X1 U8639 ( .A1(n7370), .A2(n7373), .ZN(n13596) );
  OR2_X1 U8640 ( .A1(n11977), .A2(n7372), .ZN(n7370) );
  NAND2_X1 U8641 ( .A1(n8800), .A2(n8799), .ZN(n13608) );
  NAND2_X1 U8642 ( .A1(n8821), .A2(n8820), .ZN(n13744) );
  NAND2_X1 U8643 ( .A1(n11565), .A2(n7439), .ZN(n7411) );
  NAND2_X1 U8644 ( .A1(n7253), .A2(n11173), .ZN(n11175) );
  NAND2_X1 U8645 ( .A1(n10357), .A2(n10356), .ZN(n10376) );
  INV_X1 U8646 ( .A(n7256), .ZN(n7255) );
  NAND2_X1 U8647 ( .A1(n9062), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7257) );
  OAI22_X1 U8648 ( .A1(n9003), .A2(n9258), .B1(n9546), .B2(n9098), .ZN(n7256)
         );
  NAND2_X1 U8649 ( .A1(n13591), .A2(n10345), .ZN(n13656) );
  INV_X1 U8650 ( .A(n13656), .ZN(n13636) );
  NAND2_X1 U8651 ( .A1(n13642), .A2(n13400), .ZN(n13659) );
  AND2_X1 U8652 ( .A1(n13642), .A2(n10059), .ZN(n13655) );
  NAND2_X1 U8653 ( .A1(n8546), .A2(n6635), .ZN(n6634) );
  INV_X2 U8654 ( .A(n14984), .ZN(n14986) );
  INV_X1 U8655 ( .A(n8507), .ZN(n13759) );
  AND2_X1 U8656 ( .A1(n13664), .A2(n13667), .ZN(n13756) );
  NAND2_X1 U8657 ( .A1(n6633), .A2(n6630), .ZN(n13765) );
  INV_X1 U8658 ( .A(n13678), .ZN(n6633) );
  INV_X1 U8659 ( .A(n6631), .ZN(n6630) );
  OAI21_X1 U8660 ( .B1(n13681), .B2(n13751), .A(n6549), .ZN(n6631) );
  NAND2_X1 U8661 ( .A1(n7260), .A2(n7259), .ZN(n7258) );
  INV_X1 U8662 ( .A(n13683), .ZN(n7259) );
  NOR2_X1 U8663 ( .A1(n13728), .A2(n6691), .ZN(n13730) );
  NAND2_X1 U8664 ( .A1(n6693), .A2(n6692), .ZN(n6691) );
  INV_X1 U8665 ( .A(n9108), .ZN(n10502) );
  AND2_X1 U8666 ( .A1(n9801), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14925) );
  AND2_X1 U8667 ( .A1(n8437), .A2(n7416), .ZN(n7415) );
  INV_X1 U8668 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7416) );
  XNOR2_X1 U8669 ( .A(n9097), .B(n7422), .ZN(n11908) );
  XNOR2_X1 U8670 ( .A(n9091), .B(P2_IR_REG_24__SCAN_IN), .ZN(n11537) );
  OAI21_X1 U8671 ( .B1(n9090), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9091) );
  INV_X1 U8672 ( .A(n9124), .ZN(n11111) );
  INV_X1 U8673 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10453) );
  INV_X1 U8674 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10272) );
  INV_X1 U8675 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9841) );
  INV_X1 U8676 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9444) );
  INV_X1 U8677 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9304) );
  INV_X1 U8678 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9301) );
  INV_X1 U8679 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9279) );
  INV_X1 U8680 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9276) );
  INV_X1 U8681 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9250) );
  INV_X1 U8682 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9263) );
  INV_X1 U8683 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6847) );
  NOR2_X1 U8684 ( .A1(n9459), .A2(n8468), .ZN(n6848) );
  NAND2_X1 U8685 ( .A1(n11525), .A2(n11524), .ZN(n11721) );
  AOI21_X1 U8686 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9769) );
  NOR2_X1 U8687 ( .A1(n9759), .A2(n9760), .ZN(n9761) );
  NOR2_X1 U8688 ( .A1(n12234), .A2(n7188), .ZN(n7185) );
  INV_X1 U8689 ( .A(n12234), .ZN(n7189) );
  OAI22_X1 U8690 ( .A1(n7188), .A2(n7187), .B1(n12234), .B2(n7190), .ZN(n7186)
         );
  NOR2_X1 U8691 ( .A1(n13824), .A2(n12234), .ZN(n7187) );
  NAND2_X1 U8692 ( .A1(n7055), .A2(n12222), .ZN(n14062) );
  NAND2_X1 U8693 ( .A1(n13811), .A2(n12457), .ZN(n7055) );
  AOI21_X1 U8694 ( .B1(n9611), .B2(n12020), .A(n9610), .ZN(n9649) );
  AND2_X1 U8695 ( .A1(n7202), .A2(n6530), .ZN(n13856) );
  AND2_X1 U8696 ( .A1(n7216), .A2(n7213), .ZN(n7212) );
  NAND2_X1 U8697 ( .A1(n7214), .A2(n7216), .ZN(n13874) );
  AND2_X1 U8698 ( .A1(n11808), .A2(n11807), .ZN(n14619) );
  NAND2_X1 U8699 ( .A1(n11421), .A2(n6505), .ZN(n11525) );
  AOI21_X1 U8700 ( .B1(n9774), .B2(P1_STATE_REG_SCAN_IN), .A(n11433), .ZN(
        n13920) );
  NAND2_X1 U8701 ( .A1(n7197), .A2(n7195), .ZN(n13915) );
  OR2_X1 U8702 ( .A1(n13901), .A2(n6519), .ZN(n7197) );
  INV_X1 U8703 ( .A(n7221), .ZN(n7217) );
  NOR2_X1 U8704 ( .A1(n12514), .A2(n9588), .ZN(n13923) );
  INV_X1 U8705 ( .A(n7205), .ZN(n6619) );
  OAI21_X1 U8706 ( .B1(n10674), .B2(n6561), .A(n7206), .ZN(n7205) );
  INV_X1 U8707 ( .A(n11015), .ZN(n7206) );
  INV_X1 U8708 ( .A(n13920), .ZN(n13947) );
  NAND2_X1 U8709 ( .A1(n12016), .A2(n12017), .ZN(n7211) );
  OR2_X1 U8710 ( .A1(n14735), .A2(n9587), .ZN(n13955) );
  NAND2_X1 U8711 ( .A1(n10489), .A2(n9771), .ZN(n12514) );
  INV_X1 U8712 ( .A(n14038), .ZN(n13957) );
  CLKBUF_X1 U8713 ( .A(n9682), .Z(n13975) );
  NOR2_X1 U8714 ( .A1(n6786), .A2(n9415), .ZN(n9226) );
  NOR2_X1 U8715 ( .A1(n9606), .A2(n14787), .ZN(n6786) );
  INV_X1 U8716 ( .A(n6777), .ZN(n9402) );
  INV_X1 U8717 ( .A(n6775), .ZN(n9626) );
  NAND2_X1 U8718 ( .A1(n9930), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6774) );
  NOR2_X1 U8719 ( .A1(n9426), .A2(n6591), .ZN(n9389) );
  NOR2_X1 U8720 ( .A1(n9475), .A2(n6783), .ZN(n9478) );
  AND2_X1 U8721 ( .A1(n10605), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6783) );
  NAND2_X1 U8722 ( .A1(n9478), .A2(n9477), .ZN(n9667) );
  NOR2_X1 U8723 ( .A1(n11113), .A2(n6785), .ZN(n11116) );
  AND2_X1 U8724 ( .A1(n11217), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U8725 ( .A1(n11116), .A2(n11115), .ZN(n11736) );
  INV_X1 U8726 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14033) );
  INV_X1 U8727 ( .A(n6780), .ZN(n14013) );
  INV_X1 U8728 ( .A(n14035), .ZN(n14290) );
  NAND2_X1 U8729 ( .A1(n14042), .A2(n6677), .ZN(n14292) );
  AND2_X1 U8730 ( .A1(n6678), .A2(n14749), .ZN(n6677) );
  OR2_X1 U8731 ( .A1(n14043), .A2(n14293), .ZN(n6678) );
  NAND2_X1 U8732 ( .A1(n14151), .A2(n7175), .ZN(n14132) );
  INV_X1 U8733 ( .A(n7172), .ZN(n14131) );
  INV_X1 U8734 ( .A(n14315), .ZN(n14156) );
  AND2_X1 U8735 ( .A1(n7180), .A2(n6520), .ZN(n14174) );
  NAND2_X1 U8736 ( .A1(n14200), .A2(n14085), .ZN(n14182) );
  NAND2_X1 U8737 ( .A1(n14217), .A2(n14080), .ZN(n14204) );
  OR2_X1 U8738 ( .A1(n14232), .A2(n14055), .ZN(n7140) );
  NAND2_X1 U8739 ( .A1(n7179), .A2(n14075), .ZN(n14244) );
  AND2_X1 U8740 ( .A1(n14271), .A2(n14052), .ZN(n14250) );
  OR3_X1 U8741 ( .A1(n14275), .A2(n14710), .A3(n14274), .ZN(n14367) );
  NAND2_X1 U8742 ( .A1(n11804), .A2(n11803), .ZN(n14607) );
  NAND2_X1 U8743 ( .A1(n11801), .A2(n12344), .ZN(n14612) );
  NAND2_X1 U8744 ( .A1(n14638), .A2(n7178), .ZN(n11821) );
  NAND2_X1 U8745 ( .A1(n14282), .A2(n14606), .ZN(n14258) );
  NAND2_X1 U8746 ( .A1(n7156), .A2(n11209), .ZN(n11276) );
  NAND2_X1 U8747 ( .A1(n11208), .A2(n11207), .ZN(n7156) );
  NAND2_X1 U8748 ( .A1(n10981), .A2(n10980), .ZN(n11227) );
  INV_X1 U8749 ( .A(n7133), .ZN(n10766) );
  AOI21_X1 U8750 ( .B1(n10616), .B2(n10615), .A(n6506), .ZN(n7133) );
  NAND2_X1 U8751 ( .A1(n7167), .A2(n7169), .ZN(n10764) );
  NAND2_X1 U8752 ( .A1(n10586), .A2(n7170), .ZN(n7167) );
  INV_X1 U8753 ( .A(n14258), .ZN(n14715) );
  INV_X1 U8754 ( .A(n14252), .ZN(n14713) );
  NAND2_X1 U8755 ( .A1(n14292), .A2(n6675), .ZN(n14373) );
  INV_X1 U8756 ( .A(n6676), .ZN(n6675) );
  OAI21_X1 U8757 ( .B1(n14293), .B2(n14780), .A(n14291), .ZN(n6676) );
  OR2_X1 U8758 ( .A1(n14295), .A2(n14294), .ZN(n6669) );
  INV_X1 U8759 ( .A(n6874), .ZN(n6873) );
  NAND2_X1 U8760 ( .A1(n7445), .A2(n14784), .ZN(n14307) );
  INV_X1 U8761 ( .A(n9174), .ZN(n12001) );
  INV_X1 U8762 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15143) );
  NOR2_X1 U8763 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6666) );
  INV_X1 U8764 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n15230) );
  CLKBUF_X1 U8765 ( .A(n9201), .Z(n14398) );
  AND2_X1 U8766 ( .A1(n9158), .A2(n9164), .ZN(n11732) );
  NAND2_X1 U8767 ( .A1(n9163), .A2(n9162), .ZN(n11596) );
  MUX2_X1 U8768 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9161), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9163) );
  INV_X1 U8769 ( .A(n7025), .ZN(n8945) );
  AOI21_X1 U8770 ( .B1(n8919), .B2(n8388), .A(n7029), .ZN(n7025) );
  XNOR2_X1 U8771 ( .A(n9186), .B(n9185), .ZN(n12257) );
  INV_X1 U8772 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11187) );
  XNOR2_X1 U8773 ( .A(n9496), .B(n9495), .ZN(n14150) );
  NAND2_X1 U8774 ( .A1(n8906), .A2(n8887), .ZN(n12035) );
  INV_X1 U8775 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10642) );
  INV_X1 U8776 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n11215) );
  INV_X1 U8777 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9447) );
  INV_X1 U8778 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9348) );
  INV_X1 U8779 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9299) );
  INV_X1 U8780 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9284) );
  INV_X1 U8781 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9270) );
  OR2_X1 U8782 ( .A1(n9269), .A2(n9268), .ZN(n9390) );
  INV_X1 U8783 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9755) );
  XNOR2_X1 U8784 ( .A(n14462), .B(n6624), .ZN(n15309) );
  INV_X1 U8785 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6624) );
  AOI21_X1 U8786 ( .B1(n14848), .B2(n14518), .A(n14519), .ZN(n15305) );
  XNOR2_X1 U8787 ( .A(n14456), .B(n6864), .ZN(n15298) );
  INV_X1 U8788 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6864) );
  XNOR2_X1 U8789 ( .A(n14473), .B(n14472), .ZN(n15299) );
  INV_X1 U8790 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6852) );
  INV_X1 U8791 ( .A(n14491), .ZN(n14492) );
  NOR2_X1 U8792 ( .A1(n14667), .A2(n14668), .ZN(n14512) );
  NOR2_X1 U8793 ( .A1(n14673), .A2(n14672), .ZN(n14671) );
  XNOR2_X1 U8794 ( .A(n14533), .B(n14534), .ZN(n14532) );
  AND2_X1 U8795 ( .A1(n12582), .A2(n6600), .ZN(n6620) );
  OR2_X1 U8796 ( .A1(n8135), .A2(n10970), .ZN(n7351) );
  INV_X1 U8797 ( .A(n12810), .ZN(n12804) );
  XNOR2_X1 U8798 ( .A(n6655), .B(n12839), .ZN(n12850) );
  OR2_X1 U8799 ( .A1(n12829), .A2(n12828), .ZN(n6655) );
  OAI22_X1 U8800 ( .A1(n12862), .A2(n13087), .B1(n15106), .B2(n9133), .ZN(
        n9134) );
  OAI22_X1 U8801 ( .A1(n12870), .A2(n13087), .B1(n15106), .B2(n8059), .ZN(
        n8060) );
  AOI21_X1 U8802 ( .B1(n8101), .B2(n8104), .A(n8103), .ZN(n8105) );
  OAI22_X1 U8803 ( .A1(n12870), .A2(n13129), .B1(n15089), .B2(n8073), .ZN(
        n8074) );
  OAI222_X1 U8804 ( .A1(P3_U3151), .A2(n12752), .B1(n13143), .B2(n9443), .C1(
        n6484), .C2(n9442), .ZN(P3_U3281) );
  NAND2_X1 U8805 ( .A1(n13208), .A2(n13162), .ZN(n13218) );
  NAND2_X1 U8806 ( .A1(n13360), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7362) );
  OR2_X1 U8807 ( .A1(n13401), .A2(n9710), .ZN(n6835) );
  INV_X1 U8808 ( .A(n6628), .ZN(n6627) );
  OAI22_X1 U8809 ( .A1(n13773), .A2(n13794), .B1(n14974), .B2(n13772), .ZN(
        n6628) );
  INV_X1 U8810 ( .A(n6658), .ZN(n6657) );
  OAI21_X1 U8811 ( .B1(n14091), .B2(n13943), .A(n13827), .ZN(n6658) );
  INV_X1 U8812 ( .A(n14509), .ZN(n14658) );
  NOR2_X1 U8813 ( .A1(n14664), .A2(n14663), .ZN(n14662) );
  AND2_X1 U8814 ( .A1(n14509), .A2(n14508), .ZN(n14664) );
  INV_X1 U8815 ( .A(n6857), .ZN(n14530) );
  AND2_X1 U8816 ( .A1(n12568), .A2(n8009), .ZN(n6486) );
  INV_X2 U8817 ( .A(n7629), .ZN(n7787) );
  INV_X1 U8818 ( .A(n10196), .ZN(n6653) );
  AND2_X1 U8819 ( .A1(n7056), .A2(n12638), .ZN(n6487) );
  NAND4_X1 U8820 ( .A1(n8593), .A2(n8592), .A3(n8591), .A4(n8590), .ZN(n13357)
         );
  INV_X1 U8821 ( .A(n13357), .ZN(n7226) );
  AND2_X1 U8822 ( .A1(n9185), .A2(n6810), .ZN(n6488) );
  NAND4_X1 U8823 ( .A1(n7467), .A2(n7466), .A3(n7465), .A4(n7751), .ZN(n6489)
         );
  NAND2_X1 U8824 ( .A1(n8836), .A2(n8835), .ZN(n11976) );
  NOR2_X1 U8825 ( .A1(n10955), .A2(n7232), .ZN(n6490) );
  INV_X1 U8826 ( .A(n13243), .ZN(n6732) );
  NOR2_X1 U8827 ( .A1(n11872), .A2(n12712), .ZN(n6491) );
  NAND2_X2 U8828 ( .A1(n10058), .A2(n11348), .ZN(n8648) );
  AND2_X1 U8829 ( .A1(n7195), .A2(n12121), .ZN(n6492) );
  AND2_X1 U8830 ( .A1(n14081), .A2(n14220), .ZN(n6493) );
  OR2_X1 U8831 ( .A1(n6532), .A2(n13883), .ZN(n6494) );
  OR3_X1 U8832 ( .A1(n13759), .A2(n8731), .A3(n13404), .ZN(n6495) );
  INV_X1 U8833 ( .A(n7387), .ZN(n7386) );
  OAI22_X1 U8834 ( .A1(n11988), .A2(n7388), .B1(n13454), .B2(n13437), .ZN(
        n7387) );
  AND2_X1 U8835 ( .A1(n8077), .A2(n7934), .ZN(n12881) );
  INV_X1 U8836 ( .A(n6730), .ZN(n6729) );
  NAND2_X1 U8837 ( .A1(n6554), .A2(n6731), .ZN(n6730) );
  AND2_X1 U8838 ( .A1(n8033), .A2(n6745), .ZN(n6496) );
  NAND2_X1 U8839 ( .A1(n6671), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n12816) );
  OR2_X1 U8840 ( .A1(n7828), .A2(n6911), .ZN(n6497) );
  AND2_X1 U8841 ( .A1(n8365), .A2(n8364), .ZN(n8785) );
  INV_X1 U8842 ( .A(n8785), .ZN(n6708) );
  INV_X1 U8843 ( .A(n8792), .ZN(n7286) );
  INV_X1 U8844 ( .A(n11788), .ZN(n11697) );
  INV_X1 U8845 ( .A(n12330), .ZN(n7326) );
  INV_X1 U8846 ( .A(n12403), .ZN(n6803) );
  AND2_X1 U8847 ( .A1(n13147), .A2(n7012), .ZN(n6498) );
  AND2_X1 U8848 ( .A1(n7032), .A2(n6594), .ZN(n6499) );
  AND2_X1 U8849 ( .A1(n7032), .A2(SI_18_), .ZN(n6500) );
  OR3_X1 U8850 ( .A1(n10897), .A2(n6871), .A3(n12329), .ZN(n6501) );
  INV_X1 U8851 ( .A(n7153), .ZN(n14339) );
  OR2_X2 U8852 ( .A1(n14209), .A2(n14332), .ZN(n6502) );
  NAND2_X1 U8853 ( .A1(n8003), .A2(n12593), .ZN(n6503) );
  INV_X1 U8854 ( .A(n11270), .ZN(n7984) );
  INV_X1 U8855 ( .A(n9758), .ZN(n7152) );
  NAND2_X1 U8856 ( .A1(n7094), .A2(n10240), .ZN(n6504) );
  AND2_X1 U8857 ( .A1(n11426), .A2(n11424), .ZN(n6505) );
  AND2_X1 U8858 ( .A1(n12286), .A2(n12287), .ZN(n6506) );
  AND2_X1 U8859 ( .A1(n13554), .A2(n6769), .ZN(n6508) );
  INV_X1 U8860 ( .A(n11016), .ZN(n7204) );
  INV_X1 U8861 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9459) );
  AND2_X1 U8862 ( .A1(n6986), .A2(n7662), .ZN(n6510) );
  AND2_X1 U8863 ( .A1(n11031), .A2(n11197), .ZN(n6511) );
  NAND2_X1 U8864 ( .A1(n7257), .A2(n7255), .ZN(n9108) );
  OR2_X1 U8865 ( .A1(n14505), .A2(n14504), .ZN(n6512) );
  NOR2_X1 U8866 ( .A1(n13773), .A2(n13279), .ZN(n6513) );
  AND2_X1 U8867 ( .A1(n12662), .A2(n12934), .ZN(n6514) );
  NOR2_X1 U8868 ( .A1(n14339), .A2(n14082), .ZN(n6515) );
  AND3_X1 U8869 ( .A1(n7328), .A2(n12415), .A3(n7327), .ZN(n6516) );
  INV_X1 U8870 ( .A(n11318), .ZN(n6898) );
  AND2_X1 U8871 ( .A1(n13644), .A2(n13347), .ZN(n6517) );
  OR2_X1 U8872 ( .A1(n12662), .A2(n12934), .ZN(n6518) );
  OR2_X1 U8873 ( .A1(n7200), .A2(n13911), .ZN(n6519) );
  OR2_X1 U8874 ( .A1(n12896), .A2(n12878), .ZN(n8291) );
  OR2_X1 U8875 ( .A1(n14327), .A2(n14086), .ZN(n6520) );
  AND2_X1 U8876 ( .A1(n8451), .A2(n7282), .ZN(n6521) );
  INV_X1 U8877 ( .A(n7971), .ZN(n12721) );
  NAND2_X1 U8878 ( .A1(n7216), .A2(n7211), .ZN(n13944) );
  OAI21_X1 U8879 ( .B1(n12981), .B2(n7344), .A(n7341), .ZN(n12951) );
  AND2_X1 U8880 ( .A1(n10219), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6522) );
  NAND2_X1 U8881 ( .A1(n12979), .A2(n8266), .ZN(n12965) );
  AND2_X1 U8882 ( .A1(n9155), .A2(n9154), .ZN(n6523) );
  AND2_X1 U8883 ( .A1(n12538), .A2(n13005), .ZN(n6524) );
  INV_X1 U8884 ( .A(n9003), .ZN(n8546) );
  AND2_X1 U8885 ( .A1(n14173), .A2(n6520), .ZN(n6525) );
  INV_X1 U8886 ( .A(n13824), .ZN(n7191) );
  XNOR2_X1 U8887 ( .A(n8014), .B(n8016), .ZN(n8032) );
  NAND2_X1 U8888 ( .A1(n8922), .A2(n8921), .ZN(n13724) );
  AND2_X1 U8889 ( .A1(n13171), .A2(n13170), .ZN(n6526) );
  AND2_X1 U8890 ( .A1(n7214), .A2(n7212), .ZN(n6527) );
  NAND2_X1 U8891 ( .A1(n8753), .A2(n8752), .ZN(n11310) );
  INV_X1 U8892 ( .A(n12482), .ZN(n11283) );
  INV_X1 U8893 ( .A(n7999), .ZN(n6884) );
  NAND2_X1 U8894 ( .A1(n12552), .A2(n12638), .ZN(n12583) );
  XNOR2_X1 U8895 ( .A(n9210), .B(n9211), .ZN(n9606) );
  AND2_X1 U8896 ( .A1(n7213), .A2(n12017), .ZN(n6528) );
  AND2_X1 U8897 ( .A1(n7456), .A2(n7573), .ZN(n6529) );
  NAND2_X1 U8898 ( .A1(n12079), .A2(n12080), .ZN(n6530) );
  AND2_X1 U8899 ( .A1(n10274), .A2(n10281), .ZN(n6531) );
  AND2_X1 U8900 ( .A1(n7213), .A2(n13945), .ZN(n6532) );
  AND2_X1 U8901 ( .A1(n12101), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6533) );
  AND2_X1 U8902 ( .A1(n12068), .A2(n12067), .ZN(n14241) );
  INV_X1 U8903 ( .A(n14241), .ZN(n14351) );
  AND2_X1 U8904 ( .A1(n14076), .A2(n14075), .ZN(n6534) );
  AND2_X1 U8905 ( .A1(n12881), .A2(n8291), .ZN(n6535) );
  NAND2_X1 U8906 ( .A1(n8961), .A2(n8960), .ZN(n13526) );
  OR2_X1 U8907 ( .A1(n7550), .A2(n7530), .ZN(n6536) );
  INV_X1 U8908 ( .A(n8772), .ZN(n7271) );
  NAND2_X1 U8909 ( .A1(n13490), .A2(n6760), .ZN(n6763) );
  INV_X1 U8910 ( .A(n14219), .ZN(n6642) );
  AND2_X1 U8911 ( .A1(n8254), .A2(n8253), .ZN(n13000) );
  NOR2_X1 U8912 ( .A1(n12773), .A2(n12772), .ZN(n6537) );
  INV_X1 U8913 ( .A(n8715), .ZN(n7301) );
  NAND2_X1 U8914 ( .A1(n10575), .A2(n10574), .ZN(n6538) );
  NAND2_X1 U8915 ( .A1(n11719), .A2(n11718), .ZN(n6539) );
  AND2_X1 U8916 ( .A1(n14114), .A2(n7174), .ZN(n6540) );
  AND2_X1 U8917 ( .A1(n14332), .A2(n14057), .ZN(n6541) );
  NAND2_X1 U8918 ( .A1(n11458), .A2(n7987), .ZN(n6542) );
  AND2_X1 U8919 ( .A1(n6775), .A2(n6774), .ZN(n6543) );
  AND2_X1 U8920 ( .A1(n13590), .A2(n13344), .ZN(n6544) );
  INV_X1 U8921 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9193) );
  OR2_X1 U8922 ( .A1(n14473), .A2(n14472), .ZN(n6545) );
  INV_X1 U8923 ( .A(n14063), .ZN(n7119) );
  AND2_X1 U8924 ( .A1(n12486), .A2(n11644), .ZN(n7178) );
  OR3_X1 U8925 ( .A1(n7781), .A2(P3_IR_REG_20__SCAN_IN), .A3(n7084), .ZN(n6546) );
  AND2_X1 U8926 ( .A1(n7395), .A2(n7394), .ZN(n6547) );
  NOR2_X1 U8927 ( .A1(n12329), .A2(n13965), .ZN(n6548) );
  NOR2_X1 U8928 ( .A1(n13679), .A2(n6632), .ZN(n6549) );
  NOR2_X1 U8929 ( .A1(n13953), .A2(n13962), .ZN(n6550) );
  INV_X1 U8930 ( .A(n7129), .ZN(n7128) );
  NOR2_X1 U8931 ( .A1(n14156), .A2(n14060), .ZN(n7129) );
  AND2_X1 U8932 ( .A1(n7140), .A2(n7139), .ZN(n6551) );
  INV_X1 U8933 ( .A(n13911), .ZN(n7203) );
  NAND2_X1 U8934 ( .A1(n13166), .A2(n13167), .ZN(n6552) );
  INV_X1 U8935 ( .A(n7176), .ZN(n7175) );
  NOR2_X1 U8936 ( .A1(n14156), .A2(n14089), .ZN(n7176) );
  INV_X1 U8937 ( .A(n7404), .ZN(n7403) );
  NOR2_X1 U8938 ( .A1(n11983), .A2(n13300), .ZN(n7404) );
  INV_X1 U8939 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8038) );
  AND2_X1 U8940 ( .A1(n12575), .A2(n8087), .ZN(n6553) );
  NOR2_X1 U8941 ( .A1(n13328), .A2(n13185), .ZN(n6554) );
  INV_X1 U8942 ( .A(n12453), .ZN(n7306) );
  AND2_X1 U8943 ( .A1(n6764), .A2(n13459), .ZN(n6555) );
  AND2_X1 U8944 ( .A1(n9644), .A2(n6533), .ZN(n6556) );
  AND2_X1 U8945 ( .A1(n8346), .A2(SI_8_), .ZN(n6557) );
  AND2_X1 U8946 ( .A1(n12540), .A2(n12990), .ZN(n6558) );
  AND2_X1 U8947 ( .A1(n8338), .A2(SI_5_), .ZN(n6559) );
  NOR2_X1 U8948 ( .A1(n10954), .A2(n11040), .ZN(n6560) );
  INV_X1 U8949 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9261) );
  INV_X1 U8950 ( .A(n6727), .ZN(n6726) );
  NAND2_X1 U8951 ( .A1(n7009), .A2(n6728), .ZN(n6727) );
  AND2_X1 U8952 ( .A1(n7664), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6562) );
  AND2_X1 U8953 ( .A1(n6946), .A2(n6942), .ZN(n6563) );
  INV_X1 U8954 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7361) );
  INV_X1 U8955 ( .A(n6849), .ZN(n14660) );
  OAI21_X1 U8956 ( .B1(n14657), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6512), .ZN(
        n6849) );
  NOR2_X1 U8957 ( .A1(n13789), .A2(n13632), .ZN(n6564) );
  NAND2_X1 U8958 ( .A1(n7125), .A2(n14133), .ZN(n6565) );
  INV_X1 U8959 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6663) );
  OR2_X1 U8960 ( .A1(n7590), .A2(n7589), .ZN(n10240) );
  INV_X1 U8961 ( .A(n10240), .ZN(n6920) );
  AND2_X1 U8962 ( .A1(n6943), .A2(n6942), .ZN(n6566) );
  OR2_X1 U8963 ( .A1(n6696), .A2(n13576), .ZN(n6567) );
  AOI21_X1 U8964 ( .B1(n14066), .B2(n14770), .A(n7441), .ZN(n14298) );
  AND2_X1 U8965 ( .A1(n7400), .A2(n7401), .ZN(n6568) );
  AND2_X1 U8966 ( .A1(n7313), .A2(n7311), .ZN(n6569) );
  AND2_X1 U8967 ( .A1(n7778), .A2(n7777), .ZN(n6570) );
  AND2_X1 U8968 ( .A1(n14249), .A2(n14052), .ZN(n6571) );
  NOR2_X1 U8969 ( .A1(n6980), .A2(n7677), .ZN(n6979) );
  AND2_X1 U8970 ( .A1(n6898), .A2(n8218), .ZN(n6572) );
  AND2_X1 U8971 ( .A1(n9064), .A2(n9063), .ZN(n13769) );
  INV_X1 U8972 ( .A(n13769), .ZN(n6764) );
  INV_X1 U8973 ( .A(n14056), .ZN(n7138) );
  NOR2_X1 U8974 ( .A1(n14346), .A2(n13918), .ZN(n14056) );
  OR2_X1 U8975 ( .A1(n8914), .A2(n8912), .ZN(n6573) );
  OR2_X1 U8976 ( .A1(n7301), .A2(n8714), .ZN(n6574) );
  OR2_X1 U8977 ( .A1(n8951), .A2(n8949), .ZN(n6575) );
  OR2_X1 U8978 ( .A1(n8634), .A2(n8632), .ZN(n6576) );
  AND2_X1 U8979 ( .A1(n6857), .A2(n6856), .ZN(n6577) );
  OR2_X1 U8980 ( .A1(n8674), .A2(n8676), .ZN(n6578) );
  AND2_X1 U8981 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6579) );
  NAND2_X1 U8982 ( .A1(n6819), .A2(n7307), .ZN(n6580) );
  NAND2_X1 U8983 ( .A1(n8792), .A2(n7287), .ZN(n6581) );
  NAND2_X1 U8984 ( .A1(n12331), .A2(n7326), .ZN(n6582) );
  AND2_X1 U8985 ( .A1(n7316), .A2(n6825), .ZN(n6583) );
  NAND2_X1 U8986 ( .A1(n13165), .A2(n13164), .ZN(n6584) );
  INV_X1 U8987 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9168) );
  OR2_X1 U8988 ( .A1(n6494), .A2(n6528), .ZN(n6585) );
  OR2_X1 U8989 ( .A1(n7191), .A2(n7189), .ZN(n6586) );
  NAND2_X1 U8991 ( .A1(n8983), .A2(n8982), .ZN(n13507) );
  INV_X1 U8992 ( .A(n13507), .ZN(n6766) );
  INV_X1 U8993 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7085) );
  NAND2_X1 U8994 ( .A1(n13275), .A2(n7007), .ZN(n13208) );
  OR2_X1 U8995 ( .A1(n13148), .A2(n13147), .ZN(n6587) );
  NAND2_X1 U8996 ( .A1(n11614), .A2(n11613), .ZN(n14803) );
  NAND2_X1 U8997 ( .A1(n7411), .A2(n11566), .ZN(n11657) );
  NOR2_X1 U8998 ( .A1(n11977), .A2(n7374), .ZN(n6588) );
  AND2_X1 U8999 ( .A1(n12708), .A2(n13023), .ZN(n6589) );
  AND2_X1 U9000 ( .A1(n7513), .A2(n7463), .ZN(n7716) );
  AND3_X1 U9001 ( .A1(n6958), .A2(n6957), .A3(n6963), .ZN(n6590) );
  AND2_X1 U9002 ( .A1(n10593), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6591) );
  OR2_X1 U9003 ( .A1(n8907), .A2(n8383), .ZN(n6592) );
  OR2_X1 U9004 ( .A1(n6834), .A2(n6833), .ZN(n6593) );
  INV_X1 U9005 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n6865) );
  OR2_X1 U9006 ( .A1(n8382), .A2(SI_18_), .ZN(n6594) );
  INV_X1 U9007 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9642) );
  INV_X1 U9008 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9598) );
  OR2_X1 U9009 ( .A1(n7781), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6595) );
  INV_X1 U9010 ( .A(n8380), .ZN(n7035) );
  AND2_X1 U9011 ( .A1(n9350), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n6596) );
  OR2_X1 U9012 ( .A1(n9143), .A2(n9144), .ZN(n6597) );
  NAND2_X1 U9013 ( .A1(n13020), .A2(n6886), .ZN(n6598) );
  AND2_X1 U9014 ( .A1(n8373), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n6599) );
  NAND2_X1 U9015 ( .A1(n11487), .A2(n11486), .ZN(n11489) );
  OR2_X1 U9016 ( .A1(n12885), .A2(n12704), .ZN(n6600) );
  AND2_X1 U9017 ( .A1(n8262), .A2(n8254), .ZN(n6601) );
  NOR2_X1 U9018 ( .A1(n7997), .A2(n6904), .ZN(n6602) );
  AND2_X1 U9019 ( .A1(n14638), .A2(n11644), .ZN(n6603) );
  AND2_X1 U9020 ( .A1(n7220), .A2(n7217), .ZN(n6604) );
  AND2_X1 U9021 ( .A1(n10051), .A2(n13639), .ZN(n13595) );
  NAND2_X1 U9023 ( .A1(n6746), .A2(n8033), .ZN(n10027) );
  OR3_X1 U9024 ( .A1(n9966), .A2(n9750), .A3(n10046), .ZN(n14973) );
  INV_X1 U9025 ( .A(n11174), .ZN(n7254) );
  OAI21_X1 U9026 ( .B1(n11037), .B2(n7002), .A(n7000), .ZN(n11300) );
  OAI21_X1 U9027 ( .B1(n11614), .B2(n7016), .A(n7014), .ZN(n11687) );
  AND2_X1 U9028 ( .A1(n10430), .A2(n10429), .ZN(n6605) );
  AND2_X1 U9029 ( .A1(n11163), .A2(n11293), .ZN(n6606) );
  AND2_X1 U9030 ( .A1(n11860), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6607) );
  NOR2_X1 U9031 ( .A1(n11060), .A2(n11061), .ZN(n11375) );
  XOR2_X1 U9032 ( .A(n11187), .B(P1_DATAO_REG_19__SCAN_IN), .Z(n6608) );
  NAND2_X1 U9033 ( .A1(n7333), .A2(n8195), .ZN(n11130) );
  NAND2_X1 U9034 ( .A1(n7346), .A2(n8218), .ZN(n11317) );
  NAND2_X1 U9035 ( .A1(n7225), .A2(n9958), .ZN(n10360) );
  NAND2_X1 U9036 ( .A1(n7164), .A2(n7163), .ZN(n14706) );
  NAND2_X1 U9037 ( .A1(n7233), .A2(n10737), .ZN(n10956) );
  NAND2_X1 U9038 ( .A1(n7414), .A2(n10731), .ZN(n10732) );
  NOR2_X1 U9039 ( .A1(n11375), .A2(n11374), .ZN(n6609) );
  NOR2_X1 U9040 ( .A1(n10284), .A2(n10283), .ZN(n6610) );
  NAND2_X1 U9041 ( .A1(n11163), .A2(n6770), .ZN(n6773) );
  NAND2_X1 U9042 ( .A1(n8029), .A2(n8028), .ZN(n12251) );
  INV_X1 U9043 ( .A(n12251), .ZN(n6748) );
  AND2_X1 U9044 ( .A1(n7109), .A2(n7108), .ZN(n6611) );
  INV_X1 U9045 ( .A(n11862), .ZN(n6832) );
  INV_X1 U9046 ( .A(SI_18_), .ZN(n9971) );
  NAND3_X1 U9047 ( .A1(n6755), .A2(n6909), .A3(n7469), .ZN(n6612) );
  AND2_X1 U9048 ( .A1(n8404), .A2(n11580), .ZN(n6613) );
  INV_X1 U9049 ( .A(n7449), .ZN(n7340) );
  INV_X1 U9050 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7422) );
  INV_X1 U9051 ( .A(n14716), .ZN(n6867) );
  AND2_X1 U9052 ( .A1(n15030), .A2(n15010), .ZN(n13033) );
  OR3_X1 U9053 ( .A1(n10113), .A2(n9795), .A3(n10111), .ZN(n9814) );
  INV_X1 U9054 ( .A(n7920), .ZN(n6936) );
  INV_X1 U9055 ( .A(n13644), .ZN(n6771) );
  INV_X1 U9056 ( .A(n13625), .ZN(n13603) );
  NAND2_X1 U9057 ( .A1(n9722), .A2(n9721), .ZN(n13625) );
  NAND2_X1 U9058 ( .A1(n12783), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n6614) );
  INV_X1 U9059 ( .A(n12818), .ZN(n7104) );
  NAND2_X2 U9060 ( .A1(n10887), .A2(n10886), .ZN(n14778) );
  INV_X1 U9061 ( .A(n14778), .ZN(n6872) );
  AND2_X1 U9062 ( .A1(n6960), .A2(n6963), .ZN(n6615) );
  INV_X1 U9063 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7469) );
  INV_X1 U9064 ( .A(n12769), .ZN(n6687) );
  AND2_X1 U9065 ( .A1(n13808), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6616) );
  INV_X1 U9066 ( .A(n6969), .ZN(n6968) );
  OAI21_X1 U9067 ( .B1(n6616), .B2(n6970), .A(n6975), .ZN(n6969) );
  OR2_X1 U9068 ( .A1(n8063), .A2(n10305), .ZN(n10026) );
  INV_X1 U9069 ( .A(n10026), .ZN(n6745) );
  INV_X1 U9070 ( .A(n9710), .ZN(n13400) );
  XNOR2_X1 U9071 ( .A(n8462), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9710) );
  INV_X1 U9072 ( .A(n8481), .ZN(n13804) );
  NAND2_X1 U9073 ( .A1(n10222), .A2(n10240), .ZN(n6918) );
  INV_X1 U9074 ( .A(n6918), .ZN(n6917) );
  AND2_X1 U9075 ( .A1(n6745), .A2(n8313), .ZN(n6617) );
  NOR2_X1 U9076 ( .A1(n12748), .A2(n14550), .ZN(n12751) );
  XNOR2_X1 U9077 ( .A(n11917), .B(n11922), .ZN(n14996) );
  INV_X1 U9078 ( .A(n10142), .ZN(n6654) );
  NOR2_X1 U9079 ( .A1(n14552), .A2(n14551), .ZN(n14550) );
  NAND2_X1 U9080 ( .A1(n13684), .A2(n14951), .ZN(n7260) );
  NAND2_X1 U9081 ( .A1(n7382), .A2(n7386), .ZN(n13439) );
  NAND2_X1 U9082 ( .A1(n9952), .A2(n9951), .ZN(n9953) );
  NOR2_X1 U9083 ( .A1(n13682), .A2(n7258), .ZN(n13766) );
  NOR2_X1 U9084 ( .A1(n11791), .A2(n11792), .ZN(n11977) );
  OAI21_X1 U9085 ( .B1(n13561), .B2(n11982), .A(n11981), .ZN(n13550) );
  NAND2_X1 U9086 ( .A1(n10777), .A2(n10782), .ZN(n7414) );
  NAND2_X1 U9087 ( .A1(n9714), .A2(n9719), .ZN(n9889) );
  OAI22_X1 U9088 ( .A1(n11790), .A2(n11789), .B1(n11788), .B2(n11787), .ZN(
        n11791) );
  NOR2_X1 U9089 ( .A1(n10666), .A2(n10665), .ZN(n11404) );
  INV_X1 U9090 ( .A(n6840), .ZN(n6839) );
  AOI21_X1 U9091 ( .B1(n9853), .B2(n9852), .A(n9851), .ZN(n10125) );
  AOI21_X1 U9092 ( .B1(n6838), .B2(n9710), .A(n6837), .ZN(n6836) );
  AOI21_X1 U9093 ( .B1(n9536), .B2(n9525), .A(n9524), .ZN(n9527) );
  NOR2_X1 U9094 ( .A1(n11409), .A2(n14849), .ZN(n14864) );
  NOR2_X1 U9095 ( .A1(n11411), .A2(n14862), .ZN(n11414) );
  NOR2_X1 U9096 ( .A1(n14844), .A2(n14843), .ZN(n14842) );
  NAND2_X1 U9097 ( .A1(n10148), .A2(n7528), .ZN(n7560) );
  NAND4_X1 U9098 ( .A1(n7358), .A2(n6909), .A3(n7514), .A4(n7471), .ZN(n8025)
         );
  NAND2_X2 U9099 ( .A1(n7355), .A2(n6535), .ZN(n12880) );
  INV_X1 U9100 ( .A(n10099), .ZN(n8171) );
  NAND2_X1 U9101 ( .A1(n12938), .A2(n8276), .ZN(n7353) );
  NAND2_X1 U9102 ( .A1(n7676), .A2(n8215), .ZN(n11388) );
  NAND2_X1 U9103 ( .A1(n7562), .A2(n8180), .ZN(n10454) );
  NAND2_X1 U9104 ( .A1(n7332), .A2(n7330), .ZN(n11456) );
  NAND2_X1 U9105 ( .A1(n7594), .A2(n8194), .ZN(n11144) );
  NOR2_X1 U9106 ( .A1(n12867), .A2(n6638), .ZN(n8072) );
  NAND2_X1 U9107 ( .A1(n11437), .A2(n11438), .ZN(n7346) );
  OR2_X2 U9108 ( .A1(n9132), .A2(n15104), .ZN(n9136) );
  NAND2_X1 U9109 ( .A1(n7338), .A2(n7337), .ZN(n11679) );
  NAND2_X1 U9110 ( .A1(n13848), .A2(n7433), .ZN(n13901) );
  AOI21_X2 U9111 ( .B1(n12007), .B2(n12006), .A(n7430), .ZN(n13829) );
  NAND2_X1 U9112 ( .A1(n7112), .A2(n6614), .ZN(n7111) );
  AOI21_X1 U9113 ( .B1(P3_REG2_REG_2__SCAN_IN), .B2(n10216), .A(n10200), .ZN(
        n10151) );
  NOR2_X2 U9114 ( .A1(n10394), .A2(n10393), .ZN(n10682) );
  OAI21_X1 U9115 ( .B1(n10012), .B2(n10086), .A(n10011), .ZN(n10013) );
  NOR2_X1 U9116 ( .A1(n10150), .A2(n10149), .ZN(n10201) );
  XNOR2_X1 U9117 ( .A(n11544), .B(n11552), .ZN(n11247) );
  NOR2_X1 U9118 ( .A1(n6672), .A2(n10152), .ZN(n10182) );
  NAND3_X1 U9119 ( .A1(n6868), .A2(n6869), .A3(n6828), .ZN(n10946) );
  NAND2_X1 U9120 ( .A1(n8143), .A2(n8169), .ZN(n10034) );
  NOR2_X1 U9121 ( .A1(n12722), .A2(n10084), .ZN(n8143) );
  NAND2_X1 U9122 ( .A1(n6621), .A2(n6620), .ZN(P3_U3154) );
  NAND2_X1 U9123 ( .A1(n6742), .A2(n12680), .ZN(n6621) );
  NAND2_X1 U9124 ( .A1(n12552), .A2(n12949), .ZN(n7057) );
  NAND2_X1 U9125 ( .A1(n10751), .A2(n10752), .ZN(n11049) );
  NOR2_X1 U9126 ( .A1(n10070), .A2(n10069), .ZN(n10072) );
  NAND2_X1 U9127 ( .A1(n10536), .A2(n10535), .ZN(n10750) );
  NAND2_X1 U9128 ( .A1(n12722), .A2(n9923), .ZN(n10306) );
  NAND2_X1 U9129 ( .A1(n6903), .A2(n6902), .ZN(n13017) );
  XNOR2_X1 U9130 ( .A(n6743), .B(n12578), .ZN(n6742) );
  NAND2_X1 U9131 ( .A1(n6905), .A2(n6906), .ZN(n8090) );
  NAND2_X1 U9132 ( .A1(n14273), .A2(n14272), .ZN(n14271) );
  XNOR2_X1 U9133 ( .A(n14113), .B(n14112), .ZN(n14300) );
  NAND2_X1 U9134 ( .A1(n14178), .A2(n14183), .ZN(n14177) );
  NAND2_X1 U9135 ( .A1(n14145), .A2(n7123), .ZN(n7121) );
  OAI21_X1 U9136 ( .B1(n11627), .B2(n11626), .A(n12333), .ZN(n11632) );
  OAI22_X1 U9137 ( .A1(n14232), .A2(n7136), .B1(n14056), .B2(n7139), .ZN(
        n14207) );
  XNOR2_X1 U9138 ( .A(n14493), .B(n14492), .ZN(n14524) );
  XNOR2_X1 U9139 ( .A(n14505), .B(n14504), .ZN(n14657) );
  NAND3_X1 U9140 ( .A1(n14508), .A2(n6862), .A3(n14509), .ZN(n6861) );
  AND4_X2 U9141 ( .A1(n9178), .A2(n9177), .A3(n9176), .A4(n9179), .ZN(n7455)
         );
  NOR2_X2 U9142 ( .A1(n14161), .A2(n6626), .ZN(n14145) );
  NAND3_X1 U9143 ( .A1(n7419), .A2(n9093), .A3(n7420), .ZN(n8441) );
  NAND2_X1 U9144 ( .A1(n13484), .A2(n11964), .ZN(n13465) );
  OAI21_X1 U9145 ( .B1(n10381), .B2(n10380), .A(n10383), .ZN(n10384) );
  OAI21_X1 U9146 ( .B1(n13536), .B2(n11957), .A(n11956), .ZN(n13515) );
  NAND2_X1 U9147 ( .A1(n11102), .A2(n11101), .ZN(n11159) );
  AOI222_X2 U9148 ( .A1(n13625), .A2(n13469), .B1(n13468), .B2(n13628), .C1(
        n13467), .C2(n13466), .ZN(n13692) );
  OAI22_X2 U9149 ( .A1(n11784), .A2(n11783), .B1(n11788), .B2(n13346), .ZN(
        n11948) );
  NAND2_X2 U9150 ( .A1(n13627), .A2(n13626), .ZN(n13624) );
  NAND2_X1 U9151 ( .A1(n6629), .A2(n6627), .ZN(P2_U3492) );
  OR2_X1 U9152 ( .A1(n13771), .A2(n14973), .ZN(n6629) );
  NAND3_X2 U9153 ( .A1(n8573), .A2(n8574), .A3(n6634), .ZN(n10065) );
  NAND2_X1 U9154 ( .A1(n7253), .A2(n7251), .ZN(n11571) );
  NAND2_X1 U9155 ( .A1(n13927), .A2(n13928), .ZN(n13926) );
  INV_X1 U9156 ( .A(n9719), .ZN(n9892) );
  NAND2_X1 U9157 ( .A1(n9183), .A2(n6488), .ZN(n6812) );
  NAND2_X1 U9158 ( .A1(n6643), .A2(n12270), .ZN(n9881) );
  INV_X1 U9159 ( .A(n14729), .ZN(n9679) );
  NAND2_X1 U9160 ( .A1(n8708), .A2(n8347), .ZN(n6697) );
  NOR2_X2 U9161 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9142) );
  NAND2_X1 U9162 ( .A1(n9879), .A2(n9880), .ZN(n6643) );
  AND2_X2 U9163 ( .A1(n9157), .A2(n6569), .ZN(n9172) );
  NOR2_X1 U9164 ( .A1(n6667), .A2(n6666), .ZN(n6665) );
  AOI21_X2 U9165 ( .B1(n14130), .B2(n14770), .A(n14129), .ZN(n14312) );
  AND2_X4 U9166 ( .A1(n9098), .A2(n6636), .ZN(n9062) );
  NOR2_X1 U9167 ( .A1(n13390), .A2(n13391), .ZN(n13392) );
  NAND2_X1 U9168 ( .A1(n13397), .A2(n6839), .ZN(n6838) );
  NAND2_X1 U9169 ( .A1(n7266), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8442) );
  NAND2_X1 U9170 ( .A1(n6836), .A2(n6835), .ZN(P2_U3233) );
  OAI21_X1 U9171 ( .B1(n13399), .B2(n14852), .A(n14839), .ZN(n6840) );
  INV_X1 U9172 ( .A(n12888), .ZN(n6651) );
  OAI211_X1 U9173 ( .C1(n8011), .C2(n12568), .A(n8088), .B(n13019), .ZN(n8012)
         );
  NAND2_X2 U9174 ( .A1(n13289), .A2(n13291), .ZN(n13233) );
  NAND2_X1 U9175 ( .A1(n13162), .A2(n6734), .ZN(n6733) );
  OR2_X2 U9176 ( .A1(n13234), .A2(n6718), .ZN(n6715) );
  OAI21_X2 U9177 ( .B1(n13242), .B2(n13243), .A(n6729), .ZN(n13322) );
  NAND2_X1 U9178 ( .A1(n10429), .A2(n10504), .ZN(n7020) );
  OAI21_X1 U9179 ( .B1(n13148), .B2(n6498), .A(n7010), .ZN(n13254) );
  NAND2_X2 U9180 ( .A1(n13152), .A2(n13268), .ZN(n13275) );
  NAND2_X1 U9181 ( .A1(n11687), .A2(n11686), .ZN(n11896) );
  AOI21_X1 U9182 ( .B1(n10505), .B2(n7021), .A(n7019), .ZN(n10714) );
  NAND2_X1 U9183 ( .A1(n6659), .A2(n6657), .ZN(P1_U3214) );
  NAND2_X1 U9184 ( .A1(n13825), .A2(n13937), .ZN(n6659) );
  NAND4_X1 U9185 ( .A1(n6868), .A2(n6869), .A3(n9145), .A4(n6828), .ZN(n9494)
         );
  NAND2_X1 U9186 ( .A1(n13823), .A2(n13824), .ZN(n13822) );
  NAND2_X1 U9187 ( .A1(n10651), .A2(n7442), .ZN(n10672) );
  NAND2_X1 U9188 ( .A1(n9183), .A2(n9185), .ZN(n9180) );
  NAND2_X1 U9189 ( .A1(n7209), .A2(n7208), .ZN(n7215) );
  INV_X1 U9190 ( .A(n12981), .ZN(n7817) );
  NAND2_X2 U9191 ( .A1(n11388), .A2(n11387), .ZN(n11386) );
  NAND2_X1 U9192 ( .A1(n11885), .A2(n8245), .ZN(n13027) );
  NAND2_X1 U9193 ( .A1(n12612), .A2(n12561), .ZN(n12678) );
  NAND2_X2 U9194 ( .A1(n6660), .A2(n10028), .ZN(n10523) );
  NAND3_X1 U9195 ( .A1(n7463), .A2(n7457), .A3(n6661), .ZN(n7750) );
  NOR2_X1 U9196 ( .A1(n10564), .A2(n7436), .ZN(n10536) );
  NAND2_X2 U9197 ( .A1(n10979), .A2(n10978), .ZN(n12320) );
  AOI21_X2 U9198 ( .B1(n14192), .B2(n14199), .A(n6541), .ZN(n14178) );
  NAND4_X2 U9199 ( .A1(n9142), .A2(n6664), .A3(n9141), .A4(n9445), .ZN(n9144)
         );
  NOR2_X2 U9200 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n6664) );
  NAND2_X2 U9201 ( .A1(n6668), .A2(n6665), .ZN(n11945) );
  OR2_X2 U9202 ( .A1(n12458), .A2(n9605), .ZN(n9608) );
  NAND2_X1 U9203 ( .A1(n7116), .A2(n6670), .ZN(n7114) );
  NAND2_X1 U9204 ( .A1(n14271), .A2(n6571), .ZN(n14248) );
  NAND3_X1 U9205 ( .A1(n6873), .A2(n14298), .A3(n6669), .ZN(n14374) );
  NAND2_X1 U9206 ( .A1(n13676), .A2(n6683), .ZN(n13764) );
  NAND2_X1 U9207 ( .A1(n7393), .A2(n7391), .ZN(n13510) );
  NAND2_X1 U9208 ( .A1(n7995), .A2(n6602), .ZN(n6903) );
  NAND2_X1 U9209 ( .A1(n11149), .A2(n7983), .ZN(n11133) );
  NAND2_X1 U9210 ( .A1(n12932), .A2(n8008), .ZN(n12918) );
  NAND2_X1 U9211 ( .A1(n6882), .A2(n6880), .ZN(n12989) );
  NAND2_X1 U9212 ( .A1(n8438), .A2(n8437), .ZN(n8469) );
  NAND2_X2 U9213 ( .A1(n12270), .A2(n12277), .ZN(n9878) );
  NAND2_X1 U9214 ( .A1(n14205), .A2(n7432), .ZN(n14192) );
  INV_X1 U9215 ( .A(n11632), .ZN(n6681) );
  NAND2_X1 U9216 ( .A1(n6741), .A2(n6740), .ZN(n12631) );
  NAND2_X1 U9217 ( .A1(n10684), .A2(n7110), .ZN(n7106) );
  OAI21_X1 U9218 ( .B1(n10395), .B2(n7107), .A(n7106), .ZN(n11246) );
  NOR2_X1 U9219 ( .A1(n10202), .A2(n10201), .ZN(n10200) );
  INV_X1 U9220 ( .A(n12786), .ZN(n6671) );
  INV_X1 U9221 ( .A(n12770), .ZN(n7112) );
  NOR2_X2 U9222 ( .A1(n14990), .A2(n14989), .ZN(n14988) );
  OAI21_X2 U9223 ( .B1(n14988), .B2(n7092), .A(n7091), .ZN(n12768) );
  NAND2_X4 U9224 ( .A1(n9644), .A2(n12101), .ZN(n12458) );
  NOR2_X2 U9225 ( .A1(n14264), .A2(n12379), .ZN(n14251) );
  AND3_X4 U9226 ( .A1(n9609), .A2(n9608), .A3(n9607), .ZN(n14729) );
  NOR2_X2 U9227 ( .A1(n14607), .A2(n14600), .ZN(n14601) );
  NOR2_X2 U9228 ( .A1(n14034), .A2(n14096), .ZN(n14041) );
  INV_X1 U9229 ( .A(n10770), .ZN(n6673) );
  OR2_X2 U9230 ( .A1(n14700), .A2(n12314), .ZN(n10897) );
  NAND2_X1 U9231 ( .A1(n6679), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7501) );
  NAND3_X1 U9232 ( .A1(n14033), .A2(n6689), .A3(n7024), .ZN(n6679) );
  OR2_X1 U9233 ( .A1(n14300), .A2(n14710), .ZN(n14306) );
  NAND2_X1 U9234 ( .A1(n7121), .A2(n7122), .ZN(n14113) );
  NAND2_X1 U9235 ( .A1(n7143), .A2(n7145), .ZN(n7141) );
  OAI21_X1 U9236 ( .B1(n10893), .B2(n7145), .A(n12480), .ZN(n7144) );
  NAND2_X2 U9237 ( .A1(n10980), .A2(n10889), .ZN(n12478) );
  NOR2_X1 U9238 ( .A1(n10698), .A2(n10699), .ZN(n10701) );
  XNOR2_X1 U9239 ( .A(n12805), .B(n12813), .ZN(n12782) );
  NAND2_X2 U9240 ( .A1(n10735), .A2(n10734), .ZN(n10783) );
  NAND2_X1 U9241 ( .A1(n11654), .A2(n11653), .ZN(n11784) );
  NAND2_X1 U9242 ( .A1(n9957), .A2(n9956), .ZN(n7225) );
  NAND2_X1 U9243 ( .A1(n12842), .A2(n12841), .ZN(n6685) );
  INV_X1 U9244 ( .A(n12840), .ZN(n6686) );
  NAND2_X1 U9245 ( .A1(n9873), .A2(n12470), .ZN(n9928) );
  NAND2_X1 U9246 ( .A1(n9680), .A2(n9679), .ZN(n12259) );
  NOR2_X4 U9247 ( .A1(n9144), .A2(n9259), .ZN(n6868) );
  NAND2_X4 U9248 ( .A1(n9201), .A2(n11945), .ZN(n9644) );
  OAI21_X1 U9249 ( .B1(n14299), .B2(n14363), .A(n6875), .ZN(n6874) );
  OAI21_X1 U9250 ( .B1(n14916), .B2(n6689), .A(n13402), .ZN(n6837) );
  NAND2_X1 U9251 ( .A1(n6696), .A2(n13576), .ZN(n11952) );
  INV_X1 U9252 ( .A(n6696), .ZN(n13571) );
  NAND2_X1 U9253 ( .A1(n6696), .A2(n13343), .ZN(n11980) );
  AOI21_X1 U9254 ( .B1(n6696), .B2(n14812), .A(n6690), .ZN(n13216) );
  NOR2_X1 U9255 ( .A1(n13583), .A2(n6696), .ZN(n13554) );
  MUX2_X1 U9256 ( .A(n13343), .B(n6696), .S(n8754), .Z(n8913) );
  MUX2_X1 U9257 ( .A(n13343), .B(n6696), .S(n9065), .Z(n8912) );
  NAND2_X1 U9258 ( .A1(n6696), .A2(n14939), .ZN(n6692) );
  AOI21_X1 U9259 ( .B1(n13583), .B2(n6696), .A(n13221), .ZN(n6695) );
  NAND2_X1 U9260 ( .A1(n8786), .A2(n6701), .ZN(n6700) );
  NAND3_X1 U9261 ( .A1(n6715), .A2(n6714), .A3(n6712), .ZN(n6710) );
  NAND2_X1 U9262 ( .A1(n13234), .A2(n6717), .ZN(n6714) );
  NAND2_X1 U9263 ( .A1(n6710), .A2(n6719), .ZN(n13174) );
  NAND3_X1 U9264 ( .A1(n6715), .A2(n6714), .A3(n6716), .ZN(n13307) );
  NAND3_X1 U9265 ( .A1(n8605), .A2(n8334), .A3(n8337), .ZN(n6720) );
  NAND2_X1 U9266 ( .A1(n13242), .A2(n6729), .ZN(n6724) );
  AOI21_X1 U9267 ( .B1(n13242), .B2(n13183), .A(n13243), .ZN(n13247) );
  NAND3_X1 U9268 ( .A1(n6735), .A2(n6733), .A3(n6584), .ZN(n13290) );
  NAND2_X1 U9269 ( .A1(n6738), .A2(n7032), .ZN(n8883) );
  NAND2_X1 U9270 ( .A1(n8817), .A2(n8816), .ZN(n8378) );
  NAND2_X1 U9271 ( .A1(n8884), .A2(n8905), .ZN(n8886) );
  INV_X1 U9272 ( .A(n12545), .ZN(n6739) );
  XNOR2_X2 U9273 ( .A(n11582), .B(n11508), .ZN(n11581) );
  NAND2_X2 U9274 ( .A1(n6744), .A2(n7074), .ZN(n11582) );
  NAND3_X1 U9275 ( .A1(n6747), .A2(n6748), .A3(n8031), .ZN(n6746) );
  OAI21_X1 U9276 ( .B1(n6622), .B2(n6491), .A(n11873), .ZN(n12524) );
  NAND2_X1 U9277 ( .A1(n6751), .A2(n6749), .ZN(n12528) );
  NAND2_X1 U9278 ( .A1(n11871), .A2(n11873), .ZN(n6751) );
  NAND2_X1 U9279 ( .A1(n6909), .A2(n6757), .ZN(n8013) );
  AND2_X2 U9280 ( .A1(n7513), .A2(n7358), .ZN(n6757) );
  NAND3_X1 U9281 ( .A1(n6755), .A2(n6909), .A3(n6756), .ZN(n8015) );
  INV_X1 U9282 ( .A(n6763), .ZN(n13440) );
  INV_X1 U9283 ( .A(n6773), .ZN(n11658) );
  MUX2_X1 U9284 ( .A(n14787), .B(P1_REG1_REG_1__SCAN_IN), .S(n9606), .Z(n9414)
         );
  NAND3_X1 U9285 ( .A1(n12328), .A2(n12327), .A3(n6582), .ZN(n6789) );
  OAI21_X1 U9286 ( .B1(n6795), .B2(n7434), .A(n14249), .ZN(n6791) );
  OAI21_X1 U9287 ( .B1(n6796), .B2(n6794), .A(n12381), .ZN(n12384) );
  OAI21_X1 U9288 ( .B1(n12404), .B2(n6802), .A(n6801), .ZN(n12409) );
  INV_X1 U9289 ( .A(n6798), .ZN(n12408) );
  NAND2_X1 U9290 ( .A1(n9183), .A2(n6807), .ZN(n6806) );
  NAND3_X1 U9291 ( .A1(n6808), .A2(n6806), .A3(n6804), .ZN(n9579) );
  OR2_X1 U9292 ( .A1(n7308), .A2(n12313), .ZN(n6823) );
  NAND3_X1 U9293 ( .A1(n6815), .A2(n6813), .A3(n6580), .ZN(n12318) );
  OAI21_X1 U9294 ( .B1(n6821), .B2(n6823), .A(n12315), .ZN(n6818) );
  NAND2_X1 U9295 ( .A1(n6824), .A2(n6583), .ZN(n7315) );
  NAND3_X1 U9296 ( .A1(n12397), .A2(n6826), .A3(n12396), .ZN(n6824) );
  INV_X1 U9297 ( .A(n6834), .ZN(n14877) );
  MUX2_X1 U9298 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9449), .S(n6482), .Z(n14823)
         );
  NAND3_X1 U9299 ( .A1(n6859), .A2(n6858), .A3(n6855), .ZN(n6854) );
  NAND2_X1 U9300 ( .A1(n14513), .A2(n14900), .ZN(n6858) );
  INV_X1 U9301 ( .A(n14671), .ZN(n6859) );
  NOR2_X2 U9302 ( .A1(n14142), .A2(n14310), .ZN(n14135) );
  AND2_X1 U9303 ( .A1(n9875), .A2(n12280), .ZN(n9947) );
  INV_X2 U9304 ( .A(n12458), .ZN(n12041) );
  NAND4_X1 U9305 ( .A1(n6523), .A2(n9167), .A3(n6868), .A4(n6869), .ZN(n9192)
         );
  NAND2_X4 U9306 ( .A1(n6878), .A2(n6877), .ZN(n13141) );
  NAND2_X1 U9307 ( .A1(n8000), .A2(n6883), .ZN(n6882) );
  NAND2_X1 U9308 ( .A1(n13020), .A2(n8002), .ZN(n13001) );
  INV_X1 U9309 ( .A(n8002), .ZN(n6887) );
  OAI21_X1 U9310 ( .B1(n12958), .B2(n8138), .A(n8139), .ZN(n12947) );
  NAND2_X1 U9311 ( .A1(n11131), .A2(n6900), .ZN(n6899) );
  NAND2_X1 U9312 ( .A1(n12876), .A2(n6486), .ZN(n6905) );
  NOR2_X1 U9313 ( .A1(n12875), .A2(n8010), .ZN(n8011) );
  NAND2_X1 U9314 ( .A1(n10823), .A2(n6908), .ZN(n11149) );
  AND2_X2 U9315 ( .A1(n7463), .A2(n6910), .ZN(n6909) );
  NAND3_X1 U9316 ( .A1(n7513), .A2(n7358), .A3(n7463), .ZN(n7951) );
  INV_X2 U9317 ( .A(n7646), .ZN(n8124) );
  NAND2_X1 U9318 ( .A1(n10184), .A2(n10145), .ZN(n10143) );
  NAND2_X1 U9319 ( .A1(n10142), .A2(n10196), .ZN(n10145) );
  NAND2_X1 U9320 ( .A1(n6916), .A2(n6920), .ZN(n6919) );
  INV_X1 U9321 ( .A(n10222), .ZN(n6916) );
  NAND2_X1 U9322 ( .A1(n6918), .A2(n6919), .ZN(n10223) );
  OR2_X2 U9323 ( .A1(n12782), .A2(n13081), .ZN(n12810) );
  OR2_X2 U9324 ( .A1(n10701), .A2(n10700), .ZN(n6924) );
  NAND2_X1 U9325 ( .A1(n7747), .A2(n6929), .ZN(n6926) );
  NAND2_X1 U9326 ( .A1(n6926), .A2(n6927), .ZN(n7776) );
  OR2_X2 U9327 ( .A1(n7910), .A2(n6938), .ZN(n6937) );
  NAND2_X1 U9328 ( .A1(n7587), .A2(n6566), .ZN(n6941) );
  OR2_X1 U9329 ( .A1(n7859), .A2(n6954), .ZN(n6951) );
  NAND2_X1 U9330 ( .A1(n6950), .A2(n7873), .ZN(n7874) );
  NAND2_X1 U9331 ( .A1(n6951), .A2(n6952), .ZN(n7875) );
  AOI21_X1 U9332 ( .B1(n8116), .B2(n8115), .A(n6616), .ZN(n8122) );
  NAND2_X1 U9333 ( .A1(n8116), .A2(n6965), .ZN(n6957) );
  OR2_X1 U9334 ( .A1(n8116), .A2(n6966), .ZN(n6958) );
  NAND3_X1 U9335 ( .A1(n6961), .A2(n6959), .A3(n7559), .ZN(n8126) );
  NAND2_X1 U9336 ( .A1(n8116), .A2(n6615), .ZN(n6959) );
  OR2_X1 U9337 ( .A1(n8116), .A2(n6962), .ZN(n6961) );
  INV_X1 U9338 ( .A(n8123), .ZN(n6974) );
  NAND2_X1 U9339 ( .A1(n7654), .A2(n6979), .ZN(n6976) );
  NAND2_X1 U9340 ( .A1(n6976), .A2(n6977), .ZN(n7694) );
  NAND3_X1 U9341 ( .A1(n6990), .A2(n8305), .A3(n6988), .ZN(n6987) );
  NAND3_X1 U9342 ( .A1(n7947), .A2(n8156), .A3(n12881), .ZN(n6989) );
  NOR2_X2 U9343 ( .A1(n6995), .A2(n8584), .ZN(n7420) );
  NAND4_X1 U9344 ( .A1(n8434), .A2(n8431), .A3(n8430), .A4(n8433), .ZN(n6995)
         );
  AND3_X2 U9345 ( .A1(n6998), .A2(n6996), .A3(n6997), .ZN(n8434) );
  INV_X1 U9346 ( .A(n7420), .ZN(n8765) );
  INV_X2 U9347 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6996) );
  OAI21_X1 U9348 ( .B1(n6511), .B2(n7002), .A(n11200), .ZN(n7001) );
  OR2_X1 U9349 ( .A1(n11032), .A2(n7005), .ZN(n7004) );
  XNOR2_X1 U9350 ( .A(n10110), .B(n9794), .ZN(n9812) );
  NOR2_X1 U9351 ( .A1(n7023), .A2(n7022), .ZN(n7021) );
  NAND2_X1 U9352 ( .A1(n8378), .A2(n6499), .ZN(n7030) );
  NAND2_X1 U9353 ( .A1(n8669), .A2(n7039), .ZN(n7036) );
  NAND2_X1 U9354 ( .A1(n7036), .A2(n7037), .ZN(n8708) );
  NAND2_X1 U9355 ( .A1(n9000), .A2(n8999), .ZN(n9002) );
  XNOR2_X1 U9356 ( .A(n8517), .B(n8516), .ZN(n13811) );
  NAND2_X1 U9357 ( .A1(n8408), .A2(n8407), .ZN(n9060) );
  NAND2_X1 U9358 ( .A1(n8496), .A2(n8495), .ZN(n8418) );
  NAND2_X1 U9359 ( .A1(n9077), .A2(n7278), .ZN(n7277) );
  NAND2_X1 U9360 ( .A1(n7696), .A2(n7695), .ZN(n7697) );
  NAND2_X1 U9361 ( .A1(n7824), .A2(n7823), .ZN(n7842) );
  NOR2_X1 U9362 ( .A1(n8081), .A2(n8080), .ZN(n8082) );
  NAND2_X1 U9363 ( .A1(n7509), .A2(n7508), .ZN(n7587) );
  NAND2_X1 U9364 ( .A1(n8415), .A2(n8414), .ZN(n8496) );
  OAI21_X1 U9365 ( .B1(n7276), .B2(n7275), .A(n9080), .ZN(n9081) );
  NAND2_X1 U9366 ( .A1(n7845), .A2(n7844), .ZN(n7859) );
  NAND2_X1 U9367 ( .A1(n7842), .A2(n7841), .ZN(n7845) );
  NAND2_X1 U9368 ( .A1(n7697), .A2(n11215), .ZN(n7713) );
  NAND2_X1 U9369 ( .A1(n7503), .A2(n7502), .ZN(n7526) );
  NAND2_X1 U9370 ( .A1(n7821), .A2(n7820), .ZN(n7826) );
  NAND2_X1 U9371 ( .A1(n7733), .A2(n7732), .ZN(n7747) );
  INV_X1 U9372 ( .A(n7826), .ZN(n7824) );
  NOR2_X4 U9373 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n10148) );
  AND3_X1 U9374 ( .A1(n10068), .A2(n10033), .A3(n10036), .ZN(n10070) );
  NAND2_X1 U9375 ( .A1(n7057), .A2(n12638), .ZN(n12556) );
  NAND2_X1 U9376 ( .A1(n12546), .A2(n12547), .ZN(n12656) );
  OAI211_X1 U9377 ( .C1(n12677), .C2(n7072), .A(n7069), .B(n7067), .ZN(n12577)
         );
  NAND2_X1 U9378 ( .A1(n12677), .A2(n7068), .ZN(n7067) );
  NOR2_X1 U9379 ( .A1(n7070), .A2(n12569), .ZN(n7068) );
  OAI22_X1 U9380 ( .A1(n7071), .A2(n7070), .B1(n12569), .B2(n7073), .ZN(n7069)
         );
  NOR2_X1 U9381 ( .A1(n12569), .A2(n12578), .ZN(n7071) );
  NAND2_X1 U9382 ( .A1(n12578), .A2(n12569), .ZN(n7072) );
  NAND2_X1 U9383 ( .A1(n6546), .A2(n7078), .ZN(n8063) );
  NAND3_X1 U9384 ( .A1(n7795), .A2(n7465), .A3(n7085), .ZN(n7084) );
  AND2_X2 U9385 ( .A1(n7457), .A2(n6529), .ZN(n7513) );
  INV_X1 U9386 ( .A(n7087), .ZN(n11920) );
  AOI21_X1 U9387 ( .B1(n7090), .B2(n10245), .A(n10286), .ZN(n7088) );
  XNOR2_X2 U9388 ( .A(n12768), .B(n12769), .ZN(n14547) );
  NAND2_X1 U9389 ( .A1(n12784), .A2(n7096), .ZN(n7095) );
  NAND3_X1 U9390 ( .A1(n7100), .A2(n7097), .A3(n7095), .ZN(n12836) );
  NAND3_X1 U9391 ( .A1(n7102), .A2(n12816), .A3(n7101), .ZN(n7100) );
  XNOR2_X1 U9392 ( .A(n10682), .B(n10697), .ZN(n10395) );
  OAI21_X1 U9393 ( .B1(n14546), .B2(n7111), .A(n7113), .ZN(n12814) );
  XNOR2_X1 U9394 ( .A(n12814), .B(n12813), .ZN(n12786) );
  XNOR2_X1 U9395 ( .A(n7114), .B(n14094), .ZN(n14066) );
  OAI21_X1 U9396 ( .B1(n14145), .B2(n14152), .A(n7128), .ZN(n14127) );
  NAND2_X1 U9397 ( .A1(n7130), .A2(n7134), .ZN(n10619) );
  NAND2_X1 U9398 ( .A1(n9934), .A2(n7131), .ZN(n7130) );
  INV_X1 U9399 ( .A(n7140), .ZN(n14221) );
  INV_X1 U9400 ( .A(n14220), .ZN(n7139) );
  NAND2_X1 U9401 ( .A1(n10894), .A2(n7143), .ZN(n7142) );
  NAND3_X1 U9402 ( .A1(n7142), .A2(n11228), .A3(n7141), .ZN(n11282) );
  NAND2_X1 U9403 ( .A1(n9157), .A2(n7313), .ZN(n9170) );
  NAND2_X2 U9404 ( .A1(n9644), .A2(n6636), .ZN(n12141) );
  OR2_X1 U9405 ( .A1(n9644), .A2(n9606), .ZN(n9607) );
  MUX2_X1 U9406 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14400), .S(n9644), .Z(n14279)
         );
  NAND3_X1 U9407 ( .A1(n9757), .A2(n9756), .A3(n7151), .ZN(n12268) );
  NAND2_X1 U9408 ( .A1(n12040), .A2(n7152), .ZN(n7151) );
  INV_X2 U9409 ( .A(n9644), .ZN(n12040) );
  NAND2_X1 U9410 ( .A1(n9207), .A2(n9644), .ZN(n9227) );
  NAND2_X1 U9411 ( .A1(n14399), .A2(n9644), .ZN(n7153) );
  NAND2_X1 U9412 ( .A1(n11208), .A2(n7157), .ZN(n7154) );
  NAND2_X1 U9413 ( .A1(n7154), .A2(n7155), .ZN(n11485) );
  NAND2_X1 U9414 ( .A1(n10586), .A2(n7162), .ZN(n7164) );
  AND2_X1 U9415 ( .A1(n7172), .A2(n7174), .ZN(n14115) );
  NAND2_X2 U9416 ( .A1(n7179), .A2(n6534), .ZN(n14353) );
  CLKBUF_X1 U9417 ( .A(n7183), .Z(n7180) );
  NAND2_X2 U9418 ( .A1(n7183), .A2(n6525), .ZN(n14321) );
  INV_X1 U9419 ( .A(n7180), .ZN(n14181) );
  NAND2_X1 U9420 ( .A1(n13934), .A2(n12202), .ZN(n13823) );
  OAI211_X1 U9421 ( .C1(n13934), .C2(n6586), .A(n7186), .B(n7184), .ZN(n12246)
         );
  NAND2_X1 U9422 ( .A1(n13934), .A2(n7185), .ZN(n7184) );
  NAND2_X1 U9423 ( .A1(n13901), .A2(n6492), .ZN(n7194) );
  INV_X1 U9424 ( .A(n7207), .ZN(n11014) );
  NAND2_X1 U9425 ( .A1(n12016), .A2(n6585), .ZN(n7209) );
  OR2_X1 U9426 ( .A1(n13944), .A2(n13945), .ZN(n7214) );
  NAND2_X1 U9427 ( .A1(n7215), .A2(n13882), .ZN(n13881) );
  NAND2_X1 U9428 ( .A1(n7220), .A2(n7218), .ZN(n11773) );
  NAND2_X1 U9429 ( .A1(n9156), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10641) );
  NAND2_X1 U9430 ( .A1(n10783), .A2(n7229), .ZN(n7227) );
  NAND2_X1 U9431 ( .A1(n7227), .A2(n7228), .ZN(n11102) );
  NAND2_X1 U9432 ( .A1(n13624), .A2(n7244), .ZN(n7243) );
  NAND3_X1 U9433 ( .A1(n7243), .A2(n11952), .A3(n7242), .ZN(n13546) );
  OR2_X1 U9434 ( .A1(n10384), .A2(n10726), .ZN(n10735) );
  NAND3_X1 U9435 ( .A1(n7420), .A2(n7421), .A3(n9093), .ZN(n7266) );
  OAI22_X1 U9436 ( .A1(n7268), .A2(n8595), .B1(n8596), .B2(n7267), .ZN(n8611)
         );
  OAI21_X1 U9437 ( .B1(n8756), .B2(n7273), .A(n7272), .ZN(n8771) );
  NAND2_X1 U9438 ( .A1(n7269), .A2(n7270), .ZN(n8770) );
  NAND2_X1 U9439 ( .A1(n8756), .A2(n7272), .ZN(n7269) );
  NAND2_X1 U9440 ( .A1(n8796), .A2(n7280), .ZN(n7279) );
  NAND2_X1 U9441 ( .A1(n7279), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8453) );
  AND2_X1 U9442 ( .A1(n6521), .A2(n7281), .ZN(n7280) );
  NAND2_X1 U9443 ( .A1(n7283), .A2(n7284), .ZN(n8873) );
  NAND3_X1 U9444 ( .A1(n8775), .A2(n8774), .A3(n6581), .ZN(n7283) );
  NAND4_X1 U9445 ( .A1(n8434), .A2(n8432), .A3(n8435), .A4(n7288), .ZN(n8787)
         );
  AND4_X2 U9446 ( .A1(n8435), .A2(n8432), .A3(n8434), .A4(n7289), .ZN(n8454)
         );
  NAND3_X1 U9447 ( .A1(n8898), .A2(n8897), .A3(n6573), .ZN(n7291) );
  NAND2_X1 U9448 ( .A1(n7291), .A2(n7292), .ZN(n8925) );
  NAND2_X1 U9449 ( .A1(n7293), .A2(n7294), .ZN(n8693) );
  NAND3_X1 U9450 ( .A1(n8656), .A2(n6578), .A3(n8655), .ZN(n7293) );
  NAND3_X1 U9451 ( .A1(n8616), .A2(n6576), .A3(n8615), .ZN(n7296) );
  NAND2_X1 U9452 ( .A1(n7296), .A2(n7297), .ZN(n8651) );
  OR2_X1 U9453 ( .A1(n7298), .A2(n8633), .ZN(n7297) );
  NAND2_X1 U9454 ( .A1(n7299), .A2(n7300), .ZN(n8734) );
  NAND3_X1 U9455 ( .A1(n8698), .A2(n6574), .A3(n8697), .ZN(n7299) );
  NAND2_X1 U9456 ( .A1(n7302), .A2(n7303), .ZN(n8964) );
  NAND3_X1 U9457 ( .A1(n8930), .A2(n6575), .A3(n8929), .ZN(n7302) );
  NAND2_X1 U9458 ( .A1(n7305), .A2(n7304), .ZN(n12454) );
  NAND3_X1 U9459 ( .A1(n7305), .A2(n7304), .A3(n12453), .ZN(n12456) );
  OAI22_X1 U9460 ( .A1(n12318), .A2(n7309), .B1(n12319), .B2(n7310), .ZN(
        n12323) );
  NAND2_X1 U9461 ( .A1(n12323), .A2(n12324), .ZN(n12322) );
  NAND2_X1 U9462 ( .A1(n7315), .A2(n7317), .ZN(n12404) );
  NAND3_X1 U9463 ( .A1(n12386), .A2(n12385), .A3(n7318), .ZN(n7320) );
  NAND2_X1 U9464 ( .A1(n12388), .A2(n7319), .ZN(n7318) );
  NAND2_X1 U9465 ( .A1(n7320), .A2(n7321), .ZN(n12392) );
  NAND2_X1 U9466 ( .A1(n7322), .A2(n7325), .ZN(n12305) );
  NAND3_X1 U9467 ( .A1(n12298), .A2(n7323), .A3(n12297), .ZN(n7322) );
  OAI22_X1 U9468 ( .A1(n12338), .A2(n12335), .B1(n12334), .B2(n12449), .ZN(
        n12336) );
  NAND2_X1 U9469 ( .A1(n12412), .A2(n12411), .ZN(n7327) );
  NAND2_X1 U9470 ( .A1(n7328), .A2(n7327), .ZN(n12413) );
  NAND2_X1 U9471 ( .A1(n7329), .A2(n8179), .ZN(n10316) );
  NAND2_X1 U9472 ( .A1(n8171), .A2(n10098), .ZN(n7329) );
  NAND2_X1 U9473 ( .A1(n11144), .A2(n7334), .ZN(n7332) );
  NAND2_X1 U9474 ( .A1(n11386), .A2(n7339), .ZN(n7338) );
  NAND2_X1 U9475 ( .A1(n7346), .A2(n6572), .ZN(n7676) );
  OAI211_X1 U9476 ( .C1(n7350), .C2(n7351), .A(n7348), .B(n7347), .ZN(P3_U3296) );
  NAND2_X1 U9477 ( .A1(n8160), .A2(n6617), .ZN(n7347) );
  XNOR2_X1 U9478 ( .A(n8134), .B(n12848), .ZN(n7350) );
  NAND2_X1 U9479 ( .A1(n7353), .A2(n7352), .ZN(n12926) );
  NAND2_X1 U9480 ( .A1(n12909), .A2(n7356), .ZN(n7355) );
  CLKBUF_X1 U9481 ( .A(n7355), .Z(n7354) );
  NAND2_X1 U9482 ( .A1(n12909), .A2(n8287), .ZN(n12898) );
  INV_X1 U9483 ( .A(n8287), .ZN(n7357) );
  NAND2_X1 U9484 ( .A1(n13073), .A2(n6601), .ZN(n7807) );
  XNOR2_X2 U9485 ( .A(n7474), .B(n7359), .ZN(n11943) );
  NAND2_X1 U9486 ( .A1(n7497), .A2(n7472), .ZN(n7475) );
  NAND4_X2 U9487 ( .A1(n8533), .A2(n8535), .A3(n8534), .A4(n8532), .ZN(n7363)
         );
  NAND2_X1 U9488 ( .A1(n7363), .A2(n9831), .ZN(n9821) );
  OAI21_X1 U9489 ( .B1(n8540), .B2(n13360), .A(n7362), .ZN(P2_U3531) );
  AOI22_X1 U9490 ( .A1(n13466), .A2(n13358), .B1(n13628), .B2(n7363), .ZN(
        n10109) );
  NOR2_X1 U9491 ( .A1(n7365), .A2(n13579), .ZN(n7364) );
  OAI21_X2 U9492 ( .B1(n10357), .B2(n7379), .A(n7375), .ZN(n10727) );
  OAI21_X1 U9493 ( .B1(n10382), .B2(n10375), .A(n7377), .ZN(n7376) );
  NAND2_X1 U9494 ( .A1(n10727), .A2(n10726), .ZN(n10729) );
  NAND2_X1 U9495 ( .A1(n13471), .A2(n7383), .ZN(n7380) );
  NAND2_X1 U9496 ( .A1(n7380), .A2(n7381), .ZN(n13416) );
  NAND2_X1 U9497 ( .A1(n13471), .A2(n7389), .ZN(n7382) );
  NAND2_X1 U9498 ( .A1(n13550), .A2(n6568), .ZN(n7393) );
  OR2_X1 U9499 ( .A1(n13539), .A2(n13341), .ZN(n7402) );
  NAND2_X1 U9500 ( .A1(n11565), .A2(n7407), .ZN(n7405) );
  NAND2_X1 U9501 ( .A1(n7405), .A2(n7406), .ZN(n11790) );
  NAND2_X1 U9502 ( .A1(n7414), .A2(n7412), .ZN(n10951) );
  NAND2_X1 U9503 ( .A1(n8438), .A2(n7415), .ZN(n7418) );
  XNOR2_X2 U9504 ( .A(n7417), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8481) );
  NAND3_X1 U9505 ( .A1(n8447), .A2(n9093), .A3(n7438), .ZN(n9092) );
  INV_X1 U9506 ( .A(n13322), .ZN(n13323) );
  NAND2_X1 U9507 ( .A1(n8517), .A2(n8516), .ZN(n8415) );
  NAND2_X1 U9508 ( .A1(n9035), .A2(n9034), .ZN(n9067) );
  NAND2_X1 U9509 ( .A1(n8412), .A2(n8411), .ZN(n8517) );
  OR2_X1 U9510 ( .A1(n13359), .A2(n6481), .ZN(n9713) );
  NAND2_X1 U9511 ( .A1(n11896), .A2(n11895), .ZN(n13148) );
  NAND2_X1 U9512 ( .A1(n8319), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8539) );
  AOI21_X1 U9513 ( .B1(n12864), .B2(n14581), .A(n12859), .ZN(n9132) );
  NAND2_X2 U9514 ( .A1(n12256), .A2(n12262), .ZN(n12020) );
  XNOR2_X1 U9515 ( .A(n9060), .B(n9059), .ZN(n13815) );
  INV_X1 U9516 ( .A(n9060), .ZN(n8410) );
  INV_X4 U9517 ( .A(n9793), .ZN(n13521) );
  NAND2_X2 U9518 ( .A1(n6485), .A2(n10052), .ZN(n9793) );
  OR2_X1 U9519 ( .A1(n7595), .A2(n7551), .ZN(n7556) );
  NAND3_X1 U9520 ( .A1(n7498), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7499) );
  OR2_X1 U9521 ( .A1(n12035), .A2(n12141), .ZN(n12037) );
  OR2_X1 U9522 ( .A1(n12035), .A2(n9003), .ZN(n8893) );
  NAND2_X1 U9523 ( .A1(n7579), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7540) );
  NAND2_X1 U9524 ( .A1(n15238), .A2(n7499), .ZN(n7500) );
  AND2_X1 U9525 ( .A1(n12513), .A2(n12512), .ZN(n12518) );
  OR2_X1 U9526 ( .A1(n12254), .A2(n14150), .ZN(n12255) );
  NAND2_X1 U9527 ( .A1(n12254), .A2(n14150), .ZN(n12256) );
  NAND2_X1 U9528 ( .A1(n8328), .A2(n8317), .ZN(n8318) );
  INV_X1 U9529 ( .A(n9708), .ZN(n9791) );
  AND2_X1 U9530 ( .A1(n9708), .A2(n9710), .ZN(n10058) );
  XNOR2_X1 U9531 ( .A(n9708), .B(n11348), .ZN(n9709) );
  XNOR2_X1 U9532 ( .A(n14095), .B(n14094), .ZN(n14299) );
  NAND2_X1 U9533 ( .A1(n12880), .A2(n8077), .ZN(n7948) );
  INV_X2 U9534 ( .A(n13976), .ZN(n9680) );
  XNOR2_X1 U9535 ( .A(n8106), .B(n8086), .ZN(n12864) );
  INV_X1 U9536 ( .A(n8441), .ZN(n8438) );
  NAND2_X1 U9537 ( .A1(n8562), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8550) );
  NAND2_X2 U9538 ( .A1(n9932), .A2(n9931), .ZN(n12287) );
  OR2_X1 U9539 ( .A1(n13096), .A2(n12890), .ZN(n7423) );
  INV_X2 U9540 ( .A(n15087), .ZN(n15089) );
  INV_X2 U9541 ( .A(n15030), .ZN(n15032) );
  OR2_X1 U9542 ( .A1(n7550), .A2(n6653), .ZN(n7425) );
  AND2_X1 U9543 ( .A1(n6495), .A2(n6480), .ZN(n7426) );
  OR2_X1 U9544 ( .A1(n9862), .A2(n10485), .ZN(n14796) );
  CLKBUF_X3 U9545 ( .A(n9767), .Z(n12175) );
  NOR2_X1 U9546 ( .A1(n7988), .A2(n11441), .ZN(n7427) );
  NAND2_X1 U9547 ( .A1(n13680), .A2(n13338), .ZN(n7428) );
  AND2_X1 U9548 ( .A1(n14306), .A2(n14305), .ZN(n7429) );
  AND2_X1 U9549 ( .A1(n12005), .A2(n12004), .ZN(n7430) );
  OR2_X1 U9550 ( .A1(n7153), .A2(n14082), .ZN(n7432) );
  OR2_X1 U9551 ( .A1(n12064), .A2(n12063), .ZN(n7433) );
  AND2_X1 U9552 ( .A1(n12375), .A2(n12374), .ZN(n7434) );
  AND2_X1 U9553 ( .A1(n11355), .A2(n11354), .ZN(n7435) );
  AND2_X1 U9554 ( .A1(n10531), .A2(n12720), .ZN(n7436) );
  AND2_X1 U9555 ( .A1(n8131), .A2(n8130), .ZN(n7437) );
  NAND2_X1 U9556 ( .A1(n7856), .A2(n7855), .ZN(n12934) );
  INV_X1 U9557 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8427) );
  AND4_X1 U9558 ( .A1(n9056), .A2(n9055), .A3(n9054), .A4(n9053), .ZN(n13325)
         );
  OR2_X1 U9559 ( .A1(n11840), .A2(n11839), .ZN(n7440) );
  AND2_X1 U9560 ( .A1(n14065), .A2(n14064), .ZN(n7441) );
  OR2_X1 U9561 ( .A1(n10650), .A2(n10649), .ZN(n7442) );
  OR2_X1 U9562 ( .A1(n11056), .A2(n11077), .ZN(n7443) );
  AND2_X1 U9563 ( .A1(n9062), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7444) );
  AND2_X1 U9564 ( .A1(n14117), .A2(n14116), .ZN(n7445) );
  AND2_X1 U9565 ( .A1(n9072), .A2(n9073), .ZN(n7446) );
  AND2_X1 U9566 ( .A1(n8361), .A2(n8360), .ZN(n7447) );
  OAI21_X1 U9567 ( .B1(n14224), .B2(n12092), .A(n12091), .ZN(n14079) );
  NAND2_X1 U9568 ( .A1(n8563), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7448) );
  AND2_X1 U9569 ( .A1(n14569), .A2(n12712), .ZN(n7449) );
  NOR2_X1 U9570 ( .A1(n8006), .A2(n12982), .ZN(n7450) );
  INV_X1 U9571 ( .A(n12982), .ZN(n7816) );
  INV_X1 U9572 ( .A(n8101), .ZN(n12862) );
  INV_X1 U9573 ( .A(n12711), .ZN(n12526) );
  NAND2_X1 U9574 ( .A1(n10034), .A2(n8168), .ZN(n10098) );
  INV_X1 U9575 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7477) );
  INV_X1 U9576 ( .A(n12924), .ZN(n7891) );
  INV_X1 U9577 ( .A(n12487), .ZN(n14613) );
  INV_X1 U9578 ( .A(n11886), .ZN(n7998) );
  AND2_X1 U9579 ( .A1(n12282), .A2(n12281), .ZN(n7452) );
  AND4_X1 U9580 ( .A1(n12277), .A2(n6483), .A3(n12279), .A4(n12260), .ZN(n7453) );
  AND4_X1 U9581 ( .A1(n12279), .A2(n12451), .A3(n12270), .A4(n12259), .ZN(
        n7454) );
  MUX2_X1 U9582 ( .A(n6481), .B(n13359), .S(n8648), .Z(n8556) );
  NAND2_X1 U9583 ( .A1(n8561), .A2(n8560), .ZN(n8578) );
  AND2_X1 U9584 ( .A1(n8855), .A2(n8853), .ZN(n8854) );
  INV_X1 U9585 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7460) );
  INV_X1 U9586 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7465) );
  INV_X1 U9587 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8428) );
  INV_X1 U9588 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9141) );
  INV_X1 U9589 ( .A(n7833), .ZN(n7832) );
  INV_X1 U9590 ( .A(n7706), .ZN(n7705) );
  INV_X1 U9591 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7468) );
  INV_X1 U9592 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9167) );
  INV_X1 U9593 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7498) );
  OR2_X1 U9594 ( .A1(n11377), .A2(n11373), .ZN(n11374) );
  INV_X1 U9595 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U9596 ( .A1(n7832), .A2(n7831), .ZN(n7849) );
  INV_X1 U9597 ( .A(n10822), .ZN(n7979) );
  OR2_X1 U9598 ( .A1(n7828), .A2(n7527), .ZN(n7532) );
  AND4_X1 U9599 ( .A1(n7470), .A2(n8038), .A3(n7469), .A4(n7468), .ZN(n7471)
         );
  AND2_X1 U9600 ( .A1(n8801), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8876) );
  AND2_X1 U9601 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(n8952), .ZN(n8970) );
  NOR2_X1 U9602 ( .A1(n8808), .A2(n15265), .ZN(n8801) );
  AND2_X1 U9603 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8598) );
  NOR2_X1 U9604 ( .A1(n13644), .A2(n13347), .ZN(n11656) );
  INV_X1 U9605 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8437) );
  INV_X1 U9606 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11220) );
  INV_X1 U9607 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10623) );
  AND2_X1 U9608 ( .A1(n14403), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n14404) );
  INV_X1 U9609 ( .A(n7802), .ZN(n7801) );
  INV_X1 U9610 ( .A(n7900), .ZN(n7899) );
  INV_X1 U9611 ( .A(n7739), .ZN(n7738) );
  INV_X1 U9612 ( .A(n12816), .ZN(n12784) );
  INV_X1 U9613 ( .A(n11678), .ZN(n7729) );
  INV_X1 U9614 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10242) );
  INV_X1 U9615 ( .A(n11445), .ZN(n11438) );
  INV_X1 U9616 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7472) );
  AND2_X1 U9617 ( .A1(n8677), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8699) );
  AND2_X1 U9618 ( .A1(n10937), .A2(n10944), .ZN(n10938) );
  AND2_X1 U9619 ( .A1(n8876), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8915) );
  INV_X1 U9620 ( .A(n11994), .ZN(n13672) );
  OR2_X1 U9621 ( .A1(n8842), .A2(n8486), .ZN(n8808) );
  INV_X1 U9622 ( .A(n13744), .ZN(n11992) );
  INV_X1 U9623 ( .A(n11521), .ZN(n11522) );
  INV_X1 U9624 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10982) );
  INV_X1 U9625 ( .A(n12147), .ZN(n12146) );
  OR2_X1 U9626 ( .A1(n14115), .A2(n14114), .ZN(n14116) );
  NAND2_X1 U9627 ( .A1(n14208), .A2(n7153), .ZN(n14209) );
  INV_X1 U9628 ( .A(n14271), .ZN(n14275) );
  INV_X1 U9629 ( .A(n12262), .ZN(n10491) );
  INV_X1 U9630 ( .A(n14304), .ZN(n14305) );
  INV_X1 U9631 ( .A(n14199), .ZN(n14083) );
  NAND2_X1 U9632 ( .A1(n8393), .A2(SI_22_), .ZN(n8396) );
  NAND2_X1 U9633 ( .A1(n8368), .A2(n9597), .ZN(n8371) );
  NAND2_X1 U9634 ( .A1(n8354), .A2(n9278), .ZN(n8357) );
  NAND2_X1 U9635 ( .A1(n7899), .A2(n7898), .ZN(n7913) );
  OR2_X1 U9636 ( .A1(n9695), .A2(n8068), .ZN(n9918) );
  OR2_X1 U9637 ( .A1(n7913), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U9638 ( .A1(n7738), .A2(n12694), .ZN(n7755) );
  INV_X1 U9639 ( .A(n7961), .ZN(n12853) );
  AOI21_X1 U9640 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11256), .A(n11246), .ZN(
        n11544) );
  INV_X1 U9641 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11707) );
  INV_X1 U9642 ( .A(n14987), .ZN(n14991) );
  INV_X1 U9643 ( .A(n12568), .ZN(n7947) );
  AND2_X1 U9644 ( .A1(n8234), .A2(n8244), .ZN(n11758) );
  INV_X1 U9645 ( .A(n12964), .ZN(n13023) );
  INV_X1 U9646 ( .A(n10571), .ZN(n10305) );
  NAND2_X1 U9647 ( .A1(n8126), .A2(n8125), .ZN(n8130) );
  INV_X1 U9648 ( .A(n11510), .ZN(n14577) );
  NAND2_X1 U9649 ( .A1(n7361), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7496) );
  INV_X1 U9650 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8016) );
  AND2_X1 U9651 ( .A1(n9304), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n7653) );
  INV_X1 U9652 ( .A(n13351), .ZN(n11202) );
  INV_X1 U9653 ( .A(n13629), .ZN(n13258) );
  NAND2_X1 U9654 ( .A1(n8915), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8931) );
  INV_X1 U9655 ( .A(n8562), .ZN(n9052) );
  INV_X1 U9656 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n14875) );
  INV_X1 U9657 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n15265) );
  AOI22_X1 U9658 ( .A1(n13338), .A2(n13628), .B1(n13405), .B2(n13337), .ZN(
        n11973) );
  AND2_X1 U9659 ( .A1(n11965), .A2(n9104), .ZN(n13470) );
  INV_X1 U9660 ( .A(n11958), .ZN(n13520) );
  INV_X1 U9661 ( .A(n11947), .ZN(n11792) );
  INV_X1 U9662 ( .A(n13349), .ZN(n14802) );
  INV_X1 U9663 ( .A(n13655), .ZN(n13589) );
  AND2_X1 U9664 ( .A1(n13674), .A2(n13673), .ZN(n13675) );
  NAND2_X1 U9665 ( .A1(n11993), .A2(n11992), .ZN(n13620) );
  NAND2_X1 U9666 ( .A1(n9751), .A2(n10052), .ZN(n14967) );
  INV_X1 U9667 ( .A(n10433), .ZN(n10355) );
  OR2_X1 U9668 ( .A1(n9726), .A2(n9739), .ZN(n9727) );
  NAND2_X1 U9669 ( .A1(n11523), .A2(n11522), .ZN(n11524) );
  AND2_X1 U9670 ( .A1(n13849), .A2(n13847), .ZN(n12061) );
  NAND2_X1 U9671 ( .A1(n12146), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n12165) );
  AND2_X1 U9672 ( .A1(n13864), .A2(n12160), .ZN(n13892) );
  INV_X1 U9673 ( .A(n13923), .ZN(n13949) );
  NAND2_X1 U9674 ( .A1(n14749), .A2(n14609), .ZN(n10488) );
  NOR2_X1 U9675 ( .A1(n12085), .A2(n13859), .ZN(n12104) );
  NOR2_X1 U9676 ( .A1(n11810), .A2(n11809), .ZN(n11814) );
  OR2_X1 U9677 ( .A1(n11007), .A2(n11006), .ZN(n11118) );
  INV_X1 U9678 ( .A(n14208), .ZN(n14222) );
  INV_X1 U9679 ( .A(n14243), .ZN(n14076) );
  NAND2_X1 U9680 ( .A1(n10490), .A2(n10489), .ZN(n14252) );
  INV_X1 U9681 ( .A(n14058), .ZN(n14183) );
  INV_X1 U9682 ( .A(n12488), .ZN(n14049) );
  AND2_X1 U9683 ( .A1(n8371), .A2(n8370), .ZN(n8829) );
  OAI22_X1 U9684 ( .A1(n14428), .A2(n14451), .B1(P3_ADDR_REG_11__SCAN_IN), 
        .B2(n14427), .ZN(n14449) );
  INV_X1 U9685 ( .A(n12697), .ZN(n12649) );
  INV_X1 U9686 ( .A(n12689), .ZN(n12680) );
  AND2_X1 U9687 ( .A1(n7869), .A2(n7868), .ZN(n12949) );
  AND4_X1 U9688 ( .A1(n7773), .A2(n7772), .A3(n7771), .A4(n7770), .ZN(n8001)
         );
  INV_X1 U9689 ( .A(n12833), .ZN(n12848) );
  INV_X1 U9690 ( .A(n15025), .ZN(n15014) );
  AND2_X1 U9691 ( .A1(n8051), .A2(n8050), .ZN(n9699) );
  OR2_X1 U9692 ( .A1(n15085), .A2(n15041), .ZN(n14581) );
  INV_X1 U9693 ( .A(n15079), .ZN(n15065) );
  AND2_X1 U9694 ( .A1(n8036), .A2(n8035), .ZN(n9695) );
  INV_X1 U9695 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7751) );
  AND2_X1 U9696 ( .A1(n11690), .A2(n11685), .ZN(n11686) );
  OR2_X1 U9697 ( .A1(n8741), .A2(n8740), .ZN(n8778) );
  INV_X1 U9698 ( .A(n11348), .ZN(n9101) );
  AND4_X1 U9699 ( .A1(n8525), .A2(n8524), .A3(n8523), .A4(n8522), .ZN(n13279)
         );
  AND4_X1 U9700 ( .A1(n8846), .A2(n8845), .A3(n8844), .A4(n8843), .ZN(n11787)
         );
  NAND2_X1 U9701 ( .A1(n8530), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8535) );
  AND2_X1 U9702 ( .A1(n9137), .A2(n9099), .ZN(n9469) );
  INV_X1 U9703 ( .A(n14876), .ZN(n14901) );
  NOR2_X1 U9704 ( .A1(n9458), .A2(n13816), .ZN(n14910) );
  INV_X1 U9705 ( .A(n11973), .ZN(n11974) );
  INV_X1 U9706 ( .A(n11966), .ZN(n13457) );
  OR2_X1 U9707 ( .A1(n13607), .A2(n13606), .ZN(n13737) );
  INV_X1 U9709 ( .A(n13659), .ZN(n13646) );
  INV_X1 U9710 ( .A(n9804), .ZN(n10052) );
  AND2_X1 U9711 ( .A1(n9711), .A2(n6485), .ZN(n14972) );
  NAND2_X1 U9712 ( .A1(n9792), .A2(n14942), .ZN(n14951) );
  AND2_X1 U9713 ( .A1(n9748), .A2(n9747), .ZN(n9801) );
  NAND2_X1 U9714 ( .A1(n8466), .A2(n8465), .ZN(n9090) );
  AND3_X1 U9715 ( .A1(n9773), .A2(n10489), .A3(n14735), .ZN(n13952) );
  AND4_X1 U9716 ( .A1(n12227), .A2(n12226), .A3(n12225), .A4(n12224), .ZN(
        n14061) );
  AND2_X1 U9717 ( .A1(n12077), .A2(n12076), .ZN(n14077) );
  AND2_X1 U9718 ( .A1(n9228), .A2(n9208), .ZN(n9320) );
  INV_X1 U9719 ( .A(n14680), .ZN(n13980) );
  AND2_X1 U9720 ( .A1(n9320), .A2(n14398), .ZN(n14680) );
  INV_X1 U9721 ( .A(n12484), .ZN(n11475) );
  AND2_X1 U9722 ( .A1(n14282), .A2(n10763), .ZN(n14703) );
  NAND2_X1 U9723 ( .A1(n9519), .A2(n9518), .ZN(n10485) );
  AND2_X1 U9724 ( .A1(n9877), .A2(n14773), .ZN(n14363) );
  NAND2_X1 U9725 ( .A1(n9497), .A2(n12450), .ZN(n14770) );
  INV_X1 U9726 ( .A(n14363), .ZN(n14784) );
  INV_X1 U9727 ( .A(n10485), .ZN(n9861) );
  OAI21_X1 U9728 ( .B1(n11732), .B2(n9290), .A(n9289), .ZN(n9583) );
  AND2_X1 U9729 ( .A1(n9842), .A2(n9602), .ZN(n11217) );
  INV_X1 U9730 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9255) );
  AND2_X1 U9731 ( .A1(n10019), .A2(n10018), .ZN(n14987) );
  AND2_X1 U9732 ( .A1(n9916), .A2(n9915), .ZN(n12672) );
  NAND2_X1 U9733 ( .A1(n9905), .A2(n9998), .ZN(n12689) );
  AND2_X1 U9734 ( .A1(n8114), .A2(n7967), .ZN(n12572) );
  INV_X1 U9735 ( .A(n12949), .ZN(n12709) );
  INV_X1 U9736 ( .A(n11677), .ZN(n12712) );
  OR2_X1 U9737 ( .A1(n10009), .A2(n10008), .ZN(n15008) );
  OR2_X1 U9738 ( .A1(n10009), .A2(n12837), .ZN(n15002) );
  INV_X1 U9739 ( .A(n13033), .ZN(n11466) );
  INV_X1 U9740 ( .A(n8060), .ZN(n8061) );
  INV_X1 U9741 ( .A(n15106), .ZN(n15104) );
  AND2_X2 U9742 ( .A1(n9699), .A2(n8058), .ZN(n15106) );
  INV_X1 U9743 ( .A(n12896), .ZN(n13092) );
  OR2_X1 U9744 ( .A1(n13078), .A2(n13077), .ZN(n13121) );
  AND2_X1 U9745 ( .A1(n8071), .A2(n8070), .ZN(n15087) );
  INV_X1 U9746 ( .A(SI_16_), .ZN(n9678) );
  INV_X1 U9747 ( .A(n13526), .ZN(n13713) );
  INV_X1 U9748 ( .A(n14812), .ZN(n13321) );
  INV_X1 U9749 ( .A(n13228), .ZN(n13426) );
  INV_X1 U9750 ( .A(n13263), .ZN(n13344) );
  AND4_X1 U9751 ( .A1(n8806), .A2(n8805), .A3(n8804), .A4(n8803), .ZN(n13632)
         );
  OR2_X1 U9752 ( .A1(n9469), .A2(n9468), .ZN(n14839) );
  NAND2_X1 U9753 ( .A1(n13403), .A2(n13521), .ZN(n13664) );
  NAND2_X1 U9754 ( .A1(n14986), .A2(n14939), .ZN(n13755) );
  OR3_X1 U9755 ( .A1(n14920), .A2(n9966), .A3(n9965), .ZN(n14984) );
  NAND2_X1 U9756 ( .A1(n14974), .A2(n14939), .ZN(n13794) );
  INV_X2 U9757 ( .A(n14973), .ZN(n14974) );
  INV_X1 U9758 ( .A(n14918), .ZN(n14919) );
  OR2_X1 U9759 ( .A1(n14922), .A2(n10048), .ZN(n14920) );
  INV_X1 U9760 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10644) );
  INV_X1 U9761 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9350) );
  INV_X1 U9762 ( .A(n14697), .ZN(n14760) );
  INV_X1 U9763 ( .A(n13952), .ZN(n13943) );
  INV_X1 U9764 ( .A(n14061), .ZN(n14065) );
  INV_X1 U9765 ( .A(n14077), .ZN(n14054) );
  INV_X1 U9766 ( .A(n14720), .ZN(n14270) );
  AND2_X1 U9767 ( .A1(n14180), .A2(n14179), .ZN(n14329) );
  INV_X1 U9768 ( .A(n14703), .ZN(n14262) );
  INV_X2 U9769 ( .A(n14282), .ZN(n14724) );
  INV_X2 U9770 ( .A(n14796), .ZN(n14798) );
  OR2_X1 U9771 ( .A1(n9862), .A2(n9861), .ZN(n14785) );
  AND2_X1 U9772 ( .A1(n9206), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9295) );
  INV_X1 U9773 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10270) );
  XNOR2_X1 U9774 ( .A(n14475), .B(n14474), .ZN(n14522) );
  INV_X2 U9775 ( .A(n12718), .ZN(P3_U3897) );
  OAI21_X1 U9776 ( .B1(n9132), .B2(n15087), .A(n8105), .ZN(P3_U3456) );
  INV_X1 U9777 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7528) );
  NOR2_X1 U9778 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7459) );
  NOR2_X2 U9779 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7458) );
  NAND4_X1 U9780 ( .A1(n7459), .A2(n7458), .A3(n7655), .A4(n7624), .ZN(n7700)
         );
  NAND3_X1 U9781 ( .A1(n7515), .A2(n7461), .A3(n7460), .ZN(n7462) );
  NOR2_X2 U9782 ( .A1(n7700), .A2(n7462), .ZN(n7463) );
  INV_X1 U9783 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7464) );
  NOR2_X1 U9784 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), .ZN(
        n7467) );
  NOR2_X1 U9785 ( .A1(P3_IR_REG_26__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n7470) );
  INV_X1 U9786 ( .A(n7475), .ZN(n7473) );
  NAND2_X1 U9787 ( .A1(n7473), .A2(n7477), .ZN(n7480) );
  NAND2_X1 U9788 ( .A1(n7493), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7476) );
  NAND2_X1 U9789 ( .A1(n7476), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n7479) );
  NAND2_X1 U9790 ( .A1(n7579), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7490) );
  NAND2_X1 U9791 ( .A1(n7563), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7489) );
  INV_X1 U9792 ( .A(n7564), .ZN(n7629) );
  INV_X2 U9793 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10569) );
  INV_X1 U9794 ( .A(n7580), .ZN(n7484) );
  NAND2_X1 U9795 ( .A1(n7599), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7486) );
  NAND2_X1 U9796 ( .A1(n7614), .A2(n7486), .ZN(n11137) );
  NAND2_X1 U9797 ( .A1(n7616), .A2(n11137), .ZN(n7488) );
  AND2_X2 U9798 ( .A1(n7482), .A2(n13137), .ZN(n7552) );
  NAND2_X1 U9799 ( .A1(n8107), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7487) );
  INV_X1 U9800 ( .A(n7497), .ZN(n7491) );
  NAND2_X1 U9801 ( .A1(n7491), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7492) );
  MUX2_X1 U9802 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7492), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7494) );
  NAND2_X2 U9803 ( .A1(n7494), .A2(n7493), .ZN(n12521) );
  NAND2_X1 U9804 ( .A1(n8025), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7495) );
  NAND2_X2 U9805 ( .A1(n7501), .A2(n7500), .ZN(n8328) );
  NAND2_X2 U9806 ( .A1(n7550), .A2(n6636), .ZN(n7828) );
  NAND2_X1 U9807 ( .A1(n7533), .A2(n7548), .ZN(n7503) );
  NAND2_X1 U9808 ( .A1(n8317), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7502) );
  NAND2_X1 U9809 ( .A1(n9642), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7504) );
  NAND2_X1 U9810 ( .A1(n9263), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7505) );
  NAND2_X1 U9811 ( .A1(n9755), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7507) );
  NAND2_X1 U9812 ( .A1(n7571), .A2(n7570), .ZN(n7509) );
  NAND2_X1 U9813 ( .A1(n9261), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n7508) );
  NAND2_X1 U9814 ( .A1(n9270), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n7510) );
  NAND2_X1 U9815 ( .A1(n9284), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7511) );
  NAND2_X1 U9816 ( .A1(n7512), .A2(n7511), .ZN(n7604) );
  XNOR2_X1 U9817 ( .A(n7622), .B(n7621), .ZN(n9244) );
  NAND2_X1 U9818 ( .A1(n7559), .A2(n9244), .ZN(n7520) );
  INV_X1 U9819 ( .A(SI_7_), .ZN(n9243) );
  NAND2_X1 U9820 ( .A1(n8124), .A2(n9243), .ZN(n7519) );
  BUF_X1 U9821 ( .A(n7513), .Z(n7514) );
  NAND2_X1 U9822 ( .A1(n7514), .A2(n7515), .ZN(n7607) );
  NAND2_X1 U9823 ( .A1(n7701), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7517) );
  INV_X1 U9824 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7516) );
  XNOR2_X1 U9825 ( .A(n7517), .B(n7516), .ZN(n10281) );
  NAND2_X1 U9826 ( .A1(n7797), .A2(n10281), .ZN(n7518) );
  NAND2_X1 U9827 ( .A1(n11270), .A2(n11073), .ZN(n8201) );
  NAND2_X1 U9828 ( .A1(n7579), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7524) );
  NAND2_X1 U9829 ( .A1(n7552), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7523) );
  NAND2_X1 U9830 ( .A1(n7563), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7522) );
  NAND2_X1 U9831 ( .A1(n7564), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7521) );
  XNOR2_X1 U9832 ( .A(n9263), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n7525) );
  XNOR2_X1 U9833 ( .A(n7526), .B(n7525), .ZN(n9240) );
  INV_X1 U9834 ( .A(n9240), .ZN(n7527) );
  INV_X1 U9835 ( .A(SI_2_), .ZN(n9239) );
  NAND2_X1 U9836 ( .A1(n7535), .A2(n9239), .ZN(n7531) );
  INV_X1 U9837 ( .A(n10216), .ZN(n7530) );
  AND3_X2 U9838 ( .A1(n7532), .A2(n7531), .A3(n6536), .ZN(n10106) );
  INV_X1 U9839 ( .A(n10106), .ZN(n7972) );
  NAND2_X1 U9840 ( .A1(n7971), .A2(n10106), .ZN(n8179) );
  INV_X1 U9841 ( .A(n7548), .ZN(n7534) );
  XNOR2_X1 U9842 ( .A(n7534), .B(n7533), .ZN(n9238) );
  NAND2_X1 U9843 ( .A1(n7535), .A2(SI_1_), .ZN(n7538) );
  OAI211_X2 U9844 ( .C1(n7828), .C2(n9238), .A(n7538), .B(n7537), .ZN(n10031)
         );
  INV_X1 U9845 ( .A(n10031), .ZN(n7968) );
  NAND2_X1 U9846 ( .A1(n7564), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7542) );
  NAND4_X4 U9847 ( .A1(n7542), .A2(n7541), .A3(n7540), .A4(n7539), .ZN(n10032)
         );
  NAND2_X1 U9848 ( .A1(n7579), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U9849 ( .A1(n7563), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7545) );
  NAND2_X1 U9850 ( .A1(n7564), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7544) );
  NAND2_X1 U9851 ( .A1(n7552), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7543) );
  NAND4_X1 U9852 ( .A1(n7543), .A2(n7545), .A3(n7544), .A4(n7546), .ZN(n12722)
         );
  INV_X1 U9853 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9187) );
  AND2_X1 U9854 ( .A1(n9187), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7547) );
  NOR2_X1 U9855 ( .A1(n7548), .A2(n7547), .ZN(n7549) );
  NAND2_X1 U9856 ( .A1(n8328), .A2(SI_0_), .ZN(n8537) );
  OAI21_X1 U9857 ( .B1(n12101), .B2(n7549), .A(n8537), .ZN(n13145) );
  MUX2_X1 U9858 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13145), .S(n7550), .Z(n9923)
         );
  INV_X1 U9859 ( .A(n9923), .ZN(n10084) );
  INV_X1 U9860 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n7551) );
  NAND2_X1 U9861 ( .A1(n7563), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U9862 ( .A1(n7552), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7554) );
  NAND2_X1 U9863 ( .A1(n7564), .A2(n10569), .ZN(n7553) );
  INV_X1 U9864 ( .A(SI_3_), .ZN(n9245) );
  XNOR2_X1 U9865 ( .A(n9250), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n7557) );
  XNOR2_X1 U9866 ( .A(n7558), .B(n7557), .ZN(n9246) );
  NAND2_X1 U9867 ( .A1(n7560), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7561) );
  XNOR2_X1 U9868 ( .A(n7561), .B(n7456), .ZN(n10196) );
  NAND2_X1 U9869 ( .A1(n10538), .A2(n10559), .ZN(n8180) );
  NAND2_X1 U9870 ( .A1(n10316), .A2(n10317), .ZN(n7562) );
  NAND2_X1 U9871 ( .A1(n8108), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7569) );
  NAND2_X1 U9872 ( .A1(n7579), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7568) );
  NAND2_X1 U9873 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7565) );
  NAND2_X1 U9874 ( .A1(n7580), .A2(n7565), .ZN(n10522) );
  NAND2_X1 U9875 ( .A1(n7616), .A2(n10522), .ZN(n7567) );
  NAND2_X1 U9876 ( .A1(n8107), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7566) );
  INV_X1 U9877 ( .A(SI_4_), .ZN(n9236) );
  NAND2_X1 U9878 ( .A1(n8124), .A2(n9236), .ZN(n7577) );
  XNOR2_X1 U9879 ( .A(n7571), .B(n7570), .ZN(n9235) );
  NAND2_X1 U9880 ( .A1(n7559), .A2(n9235), .ZN(n7576) );
  NAND2_X1 U9881 ( .A1(n7572), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7574) );
  INV_X1 U9882 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7573) );
  XNOR2_X1 U9883 ( .A(n7574), .B(n7573), .ZN(n10219) );
  NAND2_X1 U9884 ( .A1(n7797), .A2(n10219), .ZN(n7575) );
  NAND2_X1 U9885 ( .A1(n10753), .A2(n15051), .ZN(n8188) );
  INV_X2 U9886 ( .A(n10753), .ZN(n12719) );
  INV_X1 U9887 ( .A(n15051), .ZN(n10533) );
  NAND2_X1 U9888 ( .A1(n12719), .A2(n10533), .ZN(n8192) );
  NAND2_X2 U9889 ( .A1(n8188), .A2(n8192), .ZN(n10456) );
  INV_X1 U9890 ( .A(n10456), .ZN(n8141) );
  NAND2_X1 U9891 ( .A1(n10454), .A2(n8141), .ZN(n7578) );
  NAND2_X1 U9892 ( .A1(n7578), .A2(n8188), .ZN(n10821) );
  NAND2_X1 U9893 ( .A1(n7579), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7585) );
  NAND2_X1 U9894 ( .A1(n8107), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7584) );
  NAND2_X1 U9895 ( .A1(n7580), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n7581) );
  NAND2_X1 U9896 ( .A1(n7597), .A2(n7581), .ZN(n10827) );
  NAND2_X1 U9897 ( .A1(n7616), .A2(n10827), .ZN(n7583) );
  NAND2_X1 U9898 ( .A1(n8108), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7582) );
  XNOR2_X1 U9899 ( .A(n7587), .B(n7586), .ZN(n9233) );
  INV_X1 U9900 ( .A(SI_5_), .ZN(n9234) );
  NAND2_X1 U9901 ( .A1(n8118), .A2(n9234), .ZN(n7592) );
  NOR2_X1 U9902 ( .A1(n7514), .A2(n7083), .ZN(n7588) );
  MUX2_X1 U9903 ( .A(n7083), .B(n7588), .S(P3_IR_REG_5__SCAN_IN), .Z(n7590) );
  INV_X1 U9904 ( .A(n7607), .ZN(n7589) );
  NAND2_X1 U9905 ( .A1(n7797), .A2(n10240), .ZN(n7591) );
  AOI21_X2 U9906 ( .B1(n7559), .B2(n9233), .A(n7593), .ZN(n15057) );
  NAND2_X1 U9907 ( .A1(n11147), .A2(n15057), .ZN(n8194) );
  INV_X1 U9908 ( .A(n11147), .ZN(n12717) );
  INV_X1 U9909 ( .A(n15057), .ZN(n7980) );
  NAND2_X1 U9910 ( .A1(n12717), .A2(n7980), .ZN(n8189) );
  NAND2_X1 U9911 ( .A1(n10821), .A2(n10822), .ZN(n7594) );
  NAND2_X1 U9912 ( .A1(n8109), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9913 ( .A1(n8108), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7602) );
  NAND2_X1 U9914 ( .A1(n7597), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7598) );
  NAND2_X1 U9915 ( .A1(n7599), .A2(n7598), .ZN(n11152) );
  NAND2_X1 U9916 ( .A1(n7616), .A2(n11152), .ZN(n7601) );
  NAND2_X1 U9917 ( .A1(n8107), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7600) );
  INV_X1 U9918 ( .A(n7604), .ZN(n7605) );
  XNOR2_X1 U9919 ( .A(n7606), .B(n7605), .ZN(n9242) );
  NAND2_X1 U9920 ( .A1(n8124), .A2(SI_6_), .ZN(n7611) );
  NAND2_X1 U9921 ( .A1(n7607), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7608) );
  MUX2_X1 U9922 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7608), .S(
        P3_IR_REG_6__SCAN_IN), .Z(n7609) );
  NAND2_X1 U9923 ( .A1(n7797), .A2(n12736), .ZN(n7610) );
  OAI211_X1 U9924 ( .C1(n7828), .C2(n9242), .A(n7611), .B(n7610), .ZN(n15064)
         );
  NAND2_X1 U9925 ( .A1(n11074), .A2(n15064), .ZN(n8195) );
  INV_X2 U9926 ( .A(n11074), .ZN(n11134) );
  INV_X1 U9927 ( .A(n15064), .ZN(n7612) );
  NAND2_X1 U9928 ( .A1(n11134), .A2(n7612), .ZN(n8197) );
  INV_X1 U9929 ( .A(n11073), .ZN(n15067) );
  NAND2_X2 U9930 ( .A1(n8201), .A2(n8202), .ZN(n11132) );
  INV_X1 U9931 ( .A(n11132), .ZN(n7613) );
  NAND2_X1 U9932 ( .A1(n8108), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7620) );
  NAND2_X1 U9933 ( .A1(n8109), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7619) );
  INV_X1 U9934 ( .A(n7629), .ZN(n7616) );
  NAND2_X1 U9935 ( .A1(n7614), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n7615) );
  NAND2_X1 U9936 ( .A1(n7631), .A2(n7615), .ZN(n11462) );
  NAND2_X1 U9937 ( .A1(n7616), .A2(n11462), .ZN(n7618) );
  NAND2_X1 U9938 ( .A1(n8107), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7617) );
  XNOR2_X1 U9939 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7623) );
  XNOR2_X1 U9940 ( .A(n7638), .B(n7623), .ZN(n9247) );
  NAND2_X1 U9941 ( .A1(n8124), .A2(SI_8_), .ZN(n7627) );
  NAND2_X1 U9942 ( .A1(n7642), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7625) );
  INV_X1 U9943 ( .A(n10407), .ZN(n10291) );
  NAND2_X1 U9944 ( .A1(n7797), .A2(n10291), .ZN(n7626) );
  OAI211_X1 U9945 ( .C1(n7828), .C2(n9247), .A(n7627), .B(n7626), .ZN(n11463)
         );
  NAND2_X1 U9946 ( .A1(n11077), .A2(n11463), .ZN(n8206) );
  INV_X1 U9947 ( .A(n11077), .ZN(n12716) );
  INV_X1 U9948 ( .A(n11463), .ZN(n15072) );
  NAND2_X1 U9949 ( .A1(n12716), .A2(n15072), .ZN(n8207) );
  NAND2_X1 U9950 ( .A1(n8206), .A2(n8207), .ZN(n11458) );
  INV_X1 U9951 ( .A(n11458), .ZN(n8204) );
  NAND2_X1 U9952 ( .A1(n11456), .A2(n8204), .ZN(n7628) );
  NAND2_X1 U9953 ( .A1(n7628), .A2(n8206), .ZN(n11335) );
  NAND2_X1 U9954 ( .A1(n8109), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7636) );
  NAND2_X1 U9955 ( .A1(n7631), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n7632) );
  NAND2_X1 U9956 ( .A1(n7647), .A2(n7632), .ZN(n11342) );
  NAND2_X1 U9957 ( .A1(n7616), .A2(n11342), .ZN(n7635) );
  NAND2_X1 U9958 ( .A1(n8108), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7634) );
  NAND2_X1 U9959 ( .A1(n8107), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7633) );
  NAND4_X1 U9960 ( .A1(n7636), .A2(n7635), .A3(n7634), .A4(n7633), .ZN(n12715)
         );
  NAND2_X1 U9961 ( .A1(n9301), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n7639) );
  XNOR2_X1 U9962 ( .A(n9304), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n7641) );
  XNOR2_X1 U9963 ( .A(n7654), .B(n7641), .ZN(n9254) );
  NAND2_X1 U9964 ( .A1(n7559), .A2(n9254), .ZN(n7645) );
  OR2_X1 U9965 ( .A1(n7656), .A2(n7083), .ZN(n7643) );
  INV_X1 U9966 ( .A(n10697), .ZN(n10399) );
  NAND2_X1 U9967 ( .A1(n7797), .A2(n10399), .ZN(n7644) );
  OAI211_X1 U9968 ( .C1(n7646), .C2(SI_9_), .A(n7645), .B(n7644), .ZN(n15080)
         );
  NOR2_X1 U9969 ( .A1(n12715), .A2(n15080), .ZN(n8212) );
  NAND2_X1 U9970 ( .A1(n12715), .A2(n15080), .ZN(n8211) );
  OAI21_X1 U9971 ( .B1(n11335), .B2(n8212), .A(n8211), .ZN(n11437) );
  NAND2_X1 U9972 ( .A1(n8108), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7652) );
  NAND2_X1 U9973 ( .A1(n8109), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7651) );
  NAND2_X1 U9974 ( .A1(n7647), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7648) );
  NAND2_X1 U9975 ( .A1(n7670), .A2(n7648), .ZN(n15015) );
  NAND2_X1 U9976 ( .A1(n7616), .A2(n15015), .ZN(n7650) );
  NAND2_X1 U9977 ( .A1(n8107), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7649) );
  XNOR2_X1 U9978 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n7662) );
  XNOR2_X1 U9979 ( .A(n7663), .B(n7662), .ZN(n9273) );
  NAND2_X1 U9980 ( .A1(n9273), .A2(n7559), .ZN(n7661) );
  INV_X1 U9981 ( .A(SI_10_), .ZN(n9274) );
  NAND2_X1 U9982 ( .A1(n7656), .A2(n7655), .ZN(n7658) );
  NAND2_X1 U9983 ( .A1(n7658), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7657) );
  MUX2_X1 U9984 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7657), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n7659) );
  AOI22_X1 U9985 ( .A1(n8118), .A2(n9274), .B1(n7797), .B2(n11256), .ZN(n7660)
         );
  NAND2_X1 U9986 ( .A1(n7661), .A2(n7660), .ZN(n11452) );
  XNOR2_X1 U9987 ( .A(n11505), .B(n11452), .ZN(n11445) );
  NAND2_X1 U9988 ( .A1(n11505), .A2(n11452), .ZN(n8218) );
  XNOR2_X1 U9989 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n7665) );
  XNOR2_X1 U9990 ( .A(n7678), .B(n7665), .ZN(n9277) );
  NAND2_X1 U9991 ( .A1(n9277), .A2(n7559), .ZN(n7669) );
  NAND2_X1 U9992 ( .A1(n7680), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7667) );
  INV_X1 U9993 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7666) );
  XNOR2_X1 U9994 ( .A(n7667), .B(n7666), .ZN(n11257) );
  AOI22_X1 U9995 ( .A1(n8118), .A2(n9278), .B1(n7797), .B2(n11257), .ZN(n7668)
         );
  NAND2_X1 U9996 ( .A1(n8108), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U9997 ( .A1(n8109), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U9998 ( .A1(n7670), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U9999 ( .A1(n7687), .A2(n7671), .ZN(n11517) );
  NAND2_X1 U10000 ( .A1(n7787), .A2(n11517), .ZN(n7673) );
  NAND2_X1 U10001 ( .A1(n8107), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7672) );
  NAND2_X1 U10002 ( .A1(n11510), .A2(n11588), .ZN(n8215) );
  NAND2_X1 U10003 ( .A1(n14577), .A2(n12714), .ZN(n8217) );
  NAND2_X1 U10004 ( .A1(n8215), .A2(n8217), .ZN(n11318) );
  NAND2_X1 U10005 ( .A1(n9447), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7695) );
  NAND2_X1 U10006 ( .A1(n9444), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7679) );
  NAND2_X1 U10007 ( .A1(n7695), .A2(n7679), .ZN(n7693) );
  XNOR2_X1 U10008 ( .A(n7694), .B(n7693), .ZN(n9286) );
  NAND2_X1 U10009 ( .A1(n9286), .A2(n7559), .ZN(n7684) );
  OAI21_X1 U10010 ( .B1(n7680), .B2(P3_IR_REG_11__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7682) );
  INV_X1 U10011 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7681) );
  AOI22_X1 U10012 ( .A1(n8118), .A2(n9287), .B1(n7797), .B2(n11921), .ZN(n7683) );
  NAND2_X1 U10013 ( .A1(n7684), .A2(n7683), .ZN(n14573) );
  NAND2_X1 U10014 ( .A1(n8108), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U10015 ( .A1(n8109), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U10016 ( .A1(n7687), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7688) );
  NAND2_X1 U10017 ( .A1(n7706), .A2(n7688), .ZN(n11389) );
  NAND2_X1 U10018 ( .A1(n7787), .A2(n11389), .ZN(n7690) );
  NAND2_X1 U10019 ( .A1(n8107), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7689) );
  NAND4_X1 U10020 ( .A1(n7692), .A2(n7691), .A3(n7690), .A4(n7689), .ZN(n12713) );
  NAND2_X1 U10021 ( .A1(n14573), .A2(n12713), .ZN(n8224) );
  NAND2_X1 U10022 ( .A1(n8225), .A2(n8224), .ZN(n11382) );
  INV_X1 U10023 ( .A(n11382), .ZN(n11387) );
  NAND2_X1 U10024 ( .A1(n7698), .A2(n9598), .ZN(n7699) );
  NAND2_X1 U10025 ( .A1(n7714), .A2(n7699), .ZN(n9326) );
  NAND2_X1 U10026 ( .A1(n9326), .A2(n7559), .ZN(n7704) );
  OAI21_X1 U10027 ( .B1(n7701), .B2(n7700), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7702) );
  XNOR2_X1 U10028 ( .A(n7702), .B(P3_IR_REG_13__SCAN_IN), .ZN(n11922) );
  INV_X1 U10029 ( .A(n11922), .ZN(n14993) );
  AOI22_X1 U10030 ( .A1(n8118), .A2(n9327), .B1(n7797), .B2(n14993), .ZN(n7703) );
  NAND2_X1 U10031 ( .A1(n7704), .A2(n7703), .ZN(n14569) );
  NAND2_X1 U10032 ( .A1(n8109), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7711) );
  NAND2_X1 U10033 ( .A1(n8108), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7710) );
  NAND2_X1 U10034 ( .A1(n7706), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U10035 ( .A1(n7723), .A2(n7707), .ZN(n11706) );
  NAND2_X1 U10036 ( .A1(n7787), .A2(n11706), .ZN(n7709) );
  NAND2_X1 U10037 ( .A1(n8107), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7708) );
  NOR2_X1 U10038 ( .A1(n14569), .A2(n12712), .ZN(n8229) );
  INV_X1 U10039 ( .A(n8229), .ZN(n7712) );
  XNOR2_X1 U10040 ( .A(n9841), .B(P2_DATAO_REG_14__SCAN_IN), .ZN(n7715) );
  XNOR2_X1 U10041 ( .A(n7731), .B(n7715), .ZN(n9441) );
  NAND2_X1 U10042 ( .A1(n9441), .A2(n7559), .ZN(n7722) );
  NOR2_X1 U10043 ( .A1(n7716), .A2(n7083), .ZN(n7717) );
  MUX2_X1 U10044 ( .A(n7083), .B(n7717), .S(P3_IR_REG_14__SCAN_IN), .Z(n7719)
         );
  INV_X1 U10045 ( .A(n7750), .ZN(n7718) );
  INV_X1 U10046 ( .A(n12752), .ZN(n7720) );
  AOI22_X1 U10047 ( .A1(n8118), .A2(SI_14_), .B1(n7797), .B2(n7720), .ZN(n7721) );
  NAND2_X1 U10048 ( .A1(n8109), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7728) );
  OR2_X2 U10049 ( .A1(n7723), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U10050 ( .A1(n7723), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7724) );
  NAND2_X1 U10051 ( .A1(n7739), .A2(n7724), .ZN(n11875) );
  NAND2_X1 U10052 ( .A1(n7787), .A2(n11875), .ZN(n7727) );
  NAND2_X1 U10053 ( .A1(n8108), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7726) );
  NAND2_X1 U10054 ( .A1(n8107), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7725) );
  NAND4_X1 U10055 ( .A1(n7728), .A2(n7727), .A3(n7726), .A4(n7725), .ZN(n12711) );
  NAND2_X1 U10056 ( .A1(n11874), .A2(n12711), .ZN(n8233) );
  NAND2_X1 U10057 ( .A1(n11879), .A2(n12526), .ZN(n8238) );
  NAND2_X1 U10058 ( .A1(n8233), .A2(n8238), .ZN(n11678) );
  NAND2_X1 U10059 ( .A1(n11679), .A2(n8238), .ZN(n11759) );
  NAND2_X1 U10060 ( .A1(n9841), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n7730) );
  INV_X1 U10061 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9844) );
  NAND2_X1 U10062 ( .A1(n9844), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7732) );
  XNOR2_X1 U10063 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n7746) );
  INV_X1 U10064 ( .A(n7746), .ZN(n7734) );
  XNOR2_X1 U10065 ( .A(n7747), .B(n7734), .ZN(n9595) );
  NAND2_X1 U10066 ( .A1(n9595), .A2(n7559), .ZN(n7737) );
  NAND2_X1 U10067 ( .A1(n7750), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7735) );
  XNOR2_X1 U10068 ( .A(n7735), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U10069 ( .A1(n8118), .A2(SI_15_), .B1(n7797), .B2(n12769), .ZN(
        n7736) );
  NAND2_X1 U10070 ( .A1(n7737), .A2(n7736), .ZN(n12529) );
  NAND2_X1 U10071 ( .A1(n8109), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7744) );
  NAND2_X1 U10072 ( .A1(n7739), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7740) );
  NAND2_X1 U10073 ( .A1(n7755), .A2(n7740), .ZN(n12701) );
  NAND2_X1 U10074 ( .A1(n7787), .A2(n12701), .ZN(n7743) );
  NAND2_X1 U10075 ( .A1(n8108), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U10076 ( .A1(n8107), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7741) );
  NAND4_X1 U10077 ( .A1(n7744), .A2(n7743), .A3(n7742), .A4(n7741), .ZN(n12710) );
  OR2_X1 U10078 ( .A1(n12529), .A2(n12625), .ZN(n8234) );
  NAND2_X1 U10079 ( .A1(n12529), .A2(n12625), .ZN(n8244) );
  NAND2_X1 U10080 ( .A1(n11759), .A2(n11758), .ZN(n7745) );
  NAND2_X1 U10081 ( .A1(n7745), .A2(n8244), .ZN(n11887) );
  NAND2_X1 U10082 ( .A1(n10270), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7748) );
  XNOR2_X1 U10083 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n7761) );
  INV_X1 U10084 ( .A(n7761), .ZN(n7749) );
  XNOR2_X1 U10085 ( .A(n7762), .B(n7749), .ZN(n9676) );
  NAND2_X1 U10086 ( .A1(n9676), .A2(n7559), .ZN(n7754) );
  NAND2_X1 U10087 ( .A1(n6509), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7752) );
  XNOR2_X1 U10088 ( .A(n7752), .B(n7751), .ZN(n12783) );
  INV_X1 U10089 ( .A(n12783), .ZN(n12759) );
  AOI22_X1 U10090 ( .A1(n8118), .A2(SI_16_), .B1(n7797), .B2(n12759), .ZN(
        n7753) );
  NAND2_X1 U10091 ( .A1(n8108), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7760) );
  NAND2_X1 U10092 ( .A1(n8109), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7759) );
  OR2_X2 U10093 ( .A1(n7755), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7768) );
  NAND2_X1 U10094 ( .A1(n7755), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U10095 ( .A1(n7768), .A2(n7756), .ZN(n12622) );
  NAND2_X1 U10096 ( .A1(n7787), .A2(n12622), .ZN(n7758) );
  NAND2_X1 U10097 ( .A1(n8107), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7757) );
  OR2_X1 U10098 ( .A1(n12627), .A2(n12698), .ZN(n8235) );
  NAND2_X1 U10099 ( .A1(n12627), .A2(n12698), .ZN(n8245) );
  NAND2_X1 U10100 ( .A1(n11887), .A2(n11886), .ZN(n11885) );
  XNOR2_X1 U10101 ( .A(n10644), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n7763) );
  XNOR2_X1 U10102 ( .A(n7776), .B(n7763), .ZN(n9838) );
  NAND2_X1 U10103 ( .A1(n9838), .A2(n7559), .ZN(n7766) );
  OR2_X2 U10104 ( .A1(n6509), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n7781) );
  NAND2_X1 U10105 ( .A1(n7781), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7764) );
  XNOR2_X1 U10106 ( .A(n7764), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U10107 ( .A1(n8118), .A2(SI_17_), .B1(n7797), .B2(n12813), .ZN(
        n7765) );
  NAND2_X1 U10108 ( .A1(n8108), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7773) );
  NAND2_X1 U10109 ( .A1(n8109), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7772) );
  INV_X1 U10110 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12632) );
  NAND2_X1 U10111 ( .A1(n7768), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U10112 ( .A1(n7785), .A2(n7769), .ZN(n13029) );
  NAND2_X1 U10113 ( .A1(n7787), .A2(n13029), .ZN(n7771) );
  NAND2_X1 U10114 ( .A1(n8107), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7770) );
  OR2_X1 U10115 ( .A1(n13028), .A2(n8001), .ZN(n8255) );
  NAND2_X1 U10116 ( .A1(n13028), .A2(n8001), .ZN(n8250) );
  NAND2_X1 U10117 ( .A1(n8255), .A2(n8250), .ZN(n7999) );
  NAND2_X1 U10118 ( .A1(n13027), .A2(n6884), .ZN(n7774) );
  NAND2_X1 U10119 ( .A1(n7774), .A2(n8250), .ZN(n13012) );
  INV_X1 U10120 ( .A(n13012), .ZN(n7792) );
  AND2_X1 U10121 ( .A1(n10642), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U10122 ( .A1(n10644), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n7777) );
  NAND2_X1 U10123 ( .A1(n10948), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n7793) );
  NAND2_X1 U10124 ( .A1(n10949), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n7779) );
  OAI21_X1 U10125 ( .B1(n6570), .B2(n7780), .A(n7794), .ZN(n9970) );
  OR2_X1 U10126 ( .A1(n9970), .A2(n7828), .ZN(n7784) );
  NAND2_X1 U10127 ( .A1(n6595), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7782) );
  XNOR2_X1 U10128 ( .A(n7782), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U10129 ( .A1(n8118), .A2(SI_18_), .B1(n7797), .B2(n12841), .ZN(
        n7783) );
  INV_X1 U10130 ( .A(n13074), .ZN(n8003) );
  OR2_X2 U10131 ( .A1(n7785), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U10132 ( .A1(n7785), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U10133 ( .A1(n7802), .A2(n7786), .ZN(n12668) );
  NAND2_X1 U10134 ( .A1(n12668), .A2(n7787), .ZN(n7791) );
  NAND2_X1 U10135 ( .A1(n8109), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U10136 ( .A1(n8107), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7789) );
  NAND2_X1 U10137 ( .A1(n8108), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7788) );
  NAND4_X1 U10138 ( .A1(n7791), .A2(n7790), .A3(n7789), .A4(n7788), .ZN(n13021) );
  NAND2_X1 U10139 ( .A1(n8003), .A2(n13021), .ZN(n8254) );
  INV_X1 U10140 ( .A(n13021), .ZN(n12593) );
  NAND2_X1 U10141 ( .A1(n13074), .A2(n12593), .ZN(n8253) );
  INV_X1 U10142 ( .A(n13000), .ZN(n13011) );
  XNOR2_X1 U10143 ( .A(n7808), .B(n6608), .ZN(n10136) );
  NAND2_X1 U10144 ( .A1(n10136), .A2(n7559), .ZN(n7799) );
  INV_X1 U10145 ( .A(SI_19_), .ZN(n10135) );
  INV_X1 U10146 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7795) );
  AOI22_X1 U10147 ( .A1(n8118), .A2(n10135), .B1(n7797), .B2(n12833), .ZN(
        n7798) );
  INV_X1 U10148 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n7806) );
  INV_X1 U10149 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U10150 ( .A1(n7802), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7803) );
  NAND2_X1 U10151 ( .A1(n7811), .A2(n7803), .ZN(n12995) );
  NAND2_X1 U10152 ( .A1(n12995), .A2(n7787), .ZN(n7805) );
  AOI22_X1 U10153 ( .A1(n8109), .A2(P3_REG0_REG_19__SCAN_IN), .B1(n8108), .B2(
        P3_REG1_REG_19__SCAN_IN), .ZN(n7804) );
  OAI211_X1 U10154 ( .C1(n7965), .C2(n7806), .A(n7805), .B(n7804), .ZN(n13005)
         );
  NAND2_X1 U10155 ( .A1(n13120), .A2(n13005), .ZN(n8262) );
  OR2_X1 U10156 ( .A1(n13120), .A2(n13005), .ZN(n8263) );
  NAND2_X1 U10157 ( .A1(n7807), .A2(n8263), .ZN(n12981) );
  XNOR2_X1 U10158 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .ZN(n7818) );
  XNOR2_X1 U10159 ( .A(n7819), .B(n7818), .ZN(n10518) );
  NAND2_X1 U10160 ( .A1(n10518), .A2(n7559), .ZN(n7810) );
  NAND2_X1 U10161 ( .A1(n8124), .A2(SI_20_), .ZN(n7809) );
  OR2_X2 U10162 ( .A1(n7811), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7833) );
  NAND2_X1 U10163 ( .A1(n7811), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7812) );
  NAND2_X1 U10164 ( .A1(n7833), .A2(n7812), .ZN(n12984) );
  NAND2_X1 U10165 ( .A1(n12984), .A2(n7787), .ZN(n7815) );
  AOI22_X1 U10166 ( .A1(n8109), .A2(P3_REG0_REG_20__SCAN_IN), .B1(n8108), .B2(
        P3_REG1_REG_20__SCAN_IN), .ZN(n7814) );
  NAND2_X1 U10167 ( .A1(n8107), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U10168 ( .A1(n12983), .A2(n12963), .ZN(n8267) );
  NAND2_X1 U10169 ( .A1(n8266), .A2(n8267), .ZN(n12982) );
  NAND2_X1 U10170 ( .A1(n7819), .A2(n7818), .ZN(n7821) );
  INV_X1 U10171 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U10172 ( .A1(n11324), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7820) );
  INV_X1 U10173 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12082) );
  NAND2_X1 U10174 ( .A1(n12082), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7841) );
  INV_X1 U10175 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11112) );
  NAND2_X1 U10176 ( .A1(n11112), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n7822) );
  NAND2_X1 U10177 ( .A1(n7841), .A2(n7822), .ZN(n7825) );
  NAND2_X1 U10178 ( .A1(n7826), .A2(n7825), .ZN(n7827) );
  NAND2_X1 U10179 ( .A1(n7842), .A2(n7827), .ZN(n10573) );
  NAND2_X1 U10180 ( .A1(n8124), .A2(SI_21_), .ZN(n7829) );
  INV_X1 U10181 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n7831) );
  NAND2_X1 U10182 ( .A1(n7833), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U10183 ( .A1(n7849), .A2(n7834), .ZN(n12967) );
  NAND2_X1 U10184 ( .A1(n12967), .A2(n7787), .ZN(n7840) );
  INV_X1 U10185 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U10186 ( .A1(n8109), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n7836) );
  NAND2_X1 U10187 ( .A1(n8108), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n7835) );
  OAI211_X1 U10188 ( .C1(n7837), .C2(n7965), .A(n7836), .B(n7835), .ZN(n7838)
         );
  INV_X1 U10189 ( .A(n7838), .ZN(n7839) );
  NAND2_X1 U10190 ( .A1(n12605), .A2(n12950), .ZN(n8270) );
  NAND2_X1 U10191 ( .A1(n13112), .A2(n12976), .ZN(n8271) );
  INV_X1 U10192 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10193 ( .A1(n8395), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7858) );
  INV_X1 U10194 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11349) );
  NAND2_X1 U10195 ( .A1(n11349), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7843) );
  AND2_X1 U10196 ( .A1(n7858), .A2(n7843), .ZN(n7844) );
  OR2_X1 U10197 ( .A1(n7845), .A2(n7844), .ZN(n7846) );
  AND2_X1 U10198 ( .A1(n7859), .A2(n7846), .ZN(n10817) );
  NAND2_X1 U10199 ( .A1(n10817), .A2(n7559), .ZN(n7848) );
  NAND2_X1 U10200 ( .A1(n8124), .A2(SI_22_), .ZN(n7847) );
  OR2_X2 U10201 ( .A1(n7849), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7862) );
  NAND2_X1 U10202 ( .A1(n7849), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U10203 ( .A1(n7862), .A2(n7850), .ZN(n12953) );
  NAND2_X1 U10204 ( .A1(n12953), .A2(n7787), .ZN(n7856) );
  INV_X1 U10205 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n7853) );
  NAND2_X1 U10206 ( .A1(n8108), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n7852) );
  NAND2_X1 U10207 ( .A1(n8109), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n7851) );
  OAI211_X1 U10208 ( .C1(n7853), .C2(n7965), .A(n7852), .B(n7851), .ZN(n7854)
         );
  INV_X1 U10209 ( .A(n7854), .ZN(n7855) );
  INV_X1 U10210 ( .A(n12934), .ZN(n12961) );
  NAND2_X1 U10211 ( .A1(n12662), .A2(n12961), .ZN(n8163) );
  NAND2_X1 U10212 ( .A1(n12951), .A2(n8163), .ZN(n7857) );
  NAND2_X1 U10213 ( .A1(n13108), .A2(n12934), .ZN(n8164) );
  NAND2_X1 U10214 ( .A1(n7857), .A2(n8164), .ZN(n12938) );
  INV_X1 U10215 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7872) );
  XNOR2_X1 U10216 ( .A(n7872), .B(P2_DATAO_REG_23__SCAN_IN), .ZN(n7870) );
  XNOR2_X1 U10217 ( .A(n7871), .B(n7870), .ZN(n10969) );
  NAND2_X1 U10218 ( .A1(n10969), .A2(n7559), .ZN(n7861) );
  NAND2_X1 U10219 ( .A1(n8124), .A2(SI_23_), .ZN(n7860) );
  OR2_X2 U10220 ( .A1(n7862), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7881) );
  NAND2_X1 U10221 ( .A1(n7862), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U10222 ( .A1(n7881), .A2(n7863), .ZN(n12941) );
  NAND2_X1 U10223 ( .A1(n12941), .A2(n7787), .ZN(n7869) );
  INV_X1 U10224 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n7866) );
  NAND2_X1 U10225 ( .A1(n8108), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n7865) );
  NAND2_X1 U10226 ( .A1(n8109), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n7864) );
  OAI211_X1 U10227 ( .C1(n7866), .C2(n7965), .A(n7865), .B(n7864), .ZN(n7867)
         );
  INV_X1 U10228 ( .A(n7867), .ZN(n7868) );
  XNOR2_X1 U10229 ( .A(n12940), .B(n12949), .ZN(n12939) );
  INV_X1 U10230 ( .A(n12939), .ZN(n8276) );
  OR2_X1 U10231 ( .A1(n12940), .A2(n12949), .ZN(n8279) );
  NAND2_X1 U10232 ( .A1(n7872), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7873) );
  INV_X1 U10233 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7876) );
  XNOR2_X1 U10234 ( .A(n7892), .B(n7876), .ZN(n12247) );
  NAND2_X1 U10235 ( .A1(n12247), .A2(n7559), .ZN(n7878) );
  NAND2_X1 U10236 ( .A1(n8118), .A2(SI_24_), .ZN(n7877) );
  INV_X1 U10237 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n7879) );
  NAND2_X1 U10238 ( .A1(n7881), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7882) );
  NAND2_X1 U10239 ( .A1(n7900), .A2(n7882), .ZN(n12927) );
  NAND2_X1 U10240 ( .A1(n12927), .A2(n7787), .ZN(n7888) );
  INV_X1 U10241 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U10242 ( .A1(n8109), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n7884) );
  NAND2_X1 U10243 ( .A1(n8108), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n7883) );
  OAI211_X1 U10244 ( .C1(n7885), .C2(n7965), .A(n7884), .B(n7883), .ZN(n7886)
         );
  INV_X1 U10245 ( .A(n7886), .ZN(n7887) );
  NAND2_X1 U10246 ( .A1(n13100), .A2(n12935), .ZN(n7890) );
  INV_X1 U10247 ( .A(n13100), .ZN(n7889) );
  NAND2_X1 U10248 ( .A1(n7889), .A2(n12586), .ZN(n8281) );
  NAND2_X1 U10249 ( .A1(n12926), .A2(n8281), .ZN(n12911) );
  NAND2_X1 U10250 ( .A1(n7892), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n7894) );
  INV_X1 U10251 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11731) );
  INV_X1 U10252 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15118) );
  AOI22_X1 U10253 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n11731), .B2(n15118), .ZN(n7908) );
  INV_X1 U10254 ( .A(n7908), .ZN(n7895) );
  XNOR2_X1 U10255 ( .A(n7909), .B(n7895), .ZN(n11577) );
  NAND2_X1 U10256 ( .A1(n11577), .A2(n7559), .ZN(n7897) );
  NAND2_X1 U10257 ( .A1(n8124), .A2(SI_25_), .ZN(n7896) );
  INV_X1 U10258 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n7898) );
  NAND2_X1 U10259 ( .A1(n7900), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7901) );
  NAND2_X1 U10260 ( .A1(n7913), .A2(n7901), .ZN(n12912) );
  NAND2_X1 U10261 ( .A1(n12912), .A2(n7787), .ZN(n7906) );
  INV_X1 U10262 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n15109) );
  NAND2_X1 U10263 ( .A1(n8108), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U10264 ( .A1(n8109), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n7902) );
  OAI211_X1 U10265 ( .C1(n15109), .C2(n7965), .A(n7903), .B(n7902), .ZN(n7904)
         );
  INV_X1 U10266 ( .A(n7904), .ZN(n7905) );
  NAND2_X1 U10267 ( .A1(n13096), .A2(n12920), .ZN(n8286) );
  INV_X1 U10268 ( .A(n13096), .ZN(n7907) );
  NAND2_X1 U10269 ( .A1(n7907), .A2(n12890), .ZN(n8287) );
  NAND2_X1 U10270 ( .A1(n8286), .A2(n8287), .ZN(n12904) );
  NAND2_X1 U10271 ( .A1(n12911), .A2(n12910), .ZN(n12909) );
  NOR2_X1 U10272 ( .A1(n7909), .A2(n7908), .ZN(n7910) );
  INV_X1 U10273 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n11909) );
  INV_X1 U10274 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U10275 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n11909), .B2(n12184), .ZN(n7920) );
  XNOR2_X1 U10276 ( .A(n7921), .B(n6936), .ZN(n12250) );
  NAND2_X1 U10277 ( .A1(n12250), .A2(n7559), .ZN(n7912) );
  NAND2_X1 U10278 ( .A1(n8124), .A2(SI_26_), .ZN(n7911) );
  NAND2_X1 U10279 ( .A1(n7913), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7914) );
  NAND2_X1 U10280 ( .A1(n7926), .A2(n7914), .ZN(n12892) );
  NAND2_X1 U10281 ( .A1(n12892), .A2(n7787), .ZN(n7919) );
  INV_X1 U10282 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12894) );
  NAND2_X1 U10283 ( .A1(n8108), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n7916) );
  NAND2_X1 U10284 ( .A1(n8109), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n7915) );
  OAI211_X1 U10285 ( .C1(n12894), .C2(n7965), .A(n7916), .B(n7915), .ZN(n7917)
         );
  INV_X1 U10286 ( .A(n7917), .ZN(n7918) );
  NAND2_X1 U10287 ( .A1(n12896), .A2(n12878), .ZN(n8290) );
  NAND2_X1 U10288 ( .A1(n8291), .A2(n8290), .ZN(n12897) );
  INV_X1 U10289 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13818) );
  AOI22_X1 U10290 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13818), .B2(n15230), .ZN(n7935) );
  INV_X1 U10291 ( .A(n7935), .ZN(n7922) );
  XNOR2_X1 U10292 ( .A(n7936), .B(n7922), .ZN(n13140) );
  NAND2_X1 U10293 ( .A1(n13140), .A2(n7559), .ZN(n7924) );
  NAND2_X1 U10294 ( .A1(n8124), .A2(SI_27_), .ZN(n7923) );
  INV_X1 U10295 ( .A(n7926), .ZN(n7925) );
  INV_X1 U10296 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n12579) );
  NAND2_X1 U10297 ( .A1(n7926), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n7927) );
  NAND2_X1 U10298 ( .A1(n7941), .A2(n7927), .ZN(n12883) );
  NAND2_X1 U10299 ( .A1(n12883), .A2(n7787), .ZN(n7933) );
  INV_X1 U10300 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10301 ( .A1(n8109), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U10302 ( .A1(n8108), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n7928) );
  OAI211_X1 U10303 ( .C1(n7930), .C2(n7965), .A(n7929), .B(n7928), .ZN(n7931)
         );
  INV_X1 U10304 ( .A(n7931), .ZN(n7932) );
  NAND2_X1 U10305 ( .A1(n13036), .A2(n12891), .ZN(n8077) );
  OR2_X1 U10306 ( .A1(n13036), .A2(n12891), .ZN(n7934) );
  INV_X1 U10307 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13814) );
  AOI22_X1 U10308 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n13814), .B2(n15143), .ZN(n8080) );
  INV_X1 U10309 ( .A(n8080), .ZN(n7938) );
  XNOR2_X1 U10310 ( .A(n8081), .B(n7938), .ZN(n12519) );
  NAND2_X1 U10311 ( .A1(n12519), .A2(n7559), .ZN(n7940) );
  NAND2_X1 U10312 ( .A1(n8118), .A2(SI_28_), .ZN(n7939) );
  NAND2_X1 U10313 ( .A1(n7941), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U10314 ( .A1(n7961), .A2(n7942), .ZN(n12868) );
  INV_X1 U10315 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n7945) );
  NAND2_X1 U10316 ( .A1(n8109), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U10317 ( .A1(n8108), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7943) );
  OAI211_X1 U10318 ( .C1(n7965), .C2(n7945), .A(n7944), .B(n7943), .ZN(n7946)
         );
  NAND2_X1 U10319 ( .A1(n12575), .A2(n12877), .ZN(n8078) );
  XNOR2_X2 U10320 ( .A(n7948), .B(n7947), .ZN(n12872) );
  INV_X1 U10321 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U10322 ( .A1(n7953), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7950) );
  NAND2_X1 U10323 ( .A1(n10521), .A2(n10818), .ZN(n7955) );
  NAND2_X1 U10324 ( .A1(n7951), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7952) );
  MUX2_X1 U10325 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7952), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n7954) );
  NAND2_X1 U10326 ( .A1(n7954), .A2(n7953), .ZN(n10571) );
  AOI21_X1 U10327 ( .B1(n7955), .B2(n12848), .A(n10305), .ZN(n7957) );
  AOI21_X1 U10328 ( .B1(n10521), .B2(n10571), .A(n10818), .ZN(n7956) );
  OR2_X1 U10329 ( .A1(n7957), .A2(n7956), .ZN(n9906) );
  NAND2_X1 U10330 ( .A1(n10521), .A2(n12833), .ZN(n8161) );
  NAND2_X1 U10331 ( .A1(n7960), .A2(n10571), .ZN(n15079) );
  NOR2_X1 U10332 ( .A1(n8161), .A2(n15065), .ZN(n7958) );
  NAND2_X1 U10333 ( .A1(n9906), .A2(n7958), .ZN(n7959) );
  NAND2_X1 U10334 ( .A1(n12833), .A2(n10818), .ZN(n8053) );
  OR2_X1 U10335 ( .A1(n8053), .A2(n10521), .ZN(n8052) );
  NAND2_X1 U10336 ( .A1(n7959), .A2(n8052), .ZN(n15085) );
  AND2_X1 U10337 ( .A1(n10521), .A2(n12848), .ZN(n15023) );
  AND2_X1 U10338 ( .A1(n15023), .A2(n7960), .ZN(n15041) );
  NAND2_X1 U10339 ( .A1(n12853), .A2(n7787), .ZN(n8114) );
  INV_X1 U10340 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n7964) );
  NAND2_X1 U10341 ( .A1(n8109), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U10342 ( .A1(n8108), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7962) );
  OAI211_X1 U10343 ( .C1(n7965), .C2(n7964), .A(n7963), .B(n7962), .ZN(n7966)
         );
  INV_X1 U10344 ( .A(n7966), .ZN(n7967) );
  INV_X1 U10345 ( .A(n12521), .ZN(n8095) );
  INV_X1 U10346 ( .A(n13141), .ZN(n12837) );
  NAND2_X1 U10347 ( .A1(n8095), .A2(n12837), .ZN(n10008) );
  NAND2_X1 U10348 ( .A1(n10008), .A2(n7550), .ZN(n9919) );
  NAND2_X1 U10349 ( .A1(n8168), .A2(n8169), .ZN(n8145) );
  NAND2_X1 U10350 ( .A1(n8145), .A2(n10306), .ZN(n7970) );
  NAND2_X1 U10351 ( .A1(n10029), .A2(n7968), .ZN(n7969) );
  NAND2_X1 U10352 ( .A1(n10100), .A2(n10099), .ZN(n7974) );
  NAND2_X1 U10353 ( .A1(n10560), .A2(n7972), .ZN(n7973) );
  NAND2_X1 U10354 ( .A1(n7974), .A2(n7973), .ZN(n10318) );
  INV_X1 U10355 ( .A(n10318), .ZN(n7976) );
  INV_X1 U10356 ( .A(n10317), .ZN(n7975) );
  NAND2_X1 U10357 ( .A1(n12720), .A2(n10559), .ZN(n7977) );
  NAND2_X1 U10358 ( .A1(n10320), .A2(n7977), .ZN(n10457) );
  NAND2_X1 U10359 ( .A1(n10457), .A2(n10456), .ZN(n10455) );
  NAND2_X1 U10360 ( .A1(n12719), .A2(n15051), .ZN(n7978) );
  NAND2_X1 U10361 ( .A1(n11147), .A2(n7980), .ZN(n7981) );
  INV_X1 U10362 ( .A(n11145), .ZN(n7982) );
  NAND2_X1 U10363 ( .A1(n11134), .A2(n15064), .ZN(n7983) );
  NAND2_X1 U10364 ( .A1(n7984), .A2(n11073), .ZN(n7985) );
  INV_X1 U10365 ( .A(n15080), .ZN(n11064) );
  NAND2_X1 U10366 ( .A1(n12715), .A2(n11064), .ZN(n11439) );
  OR2_X1 U10367 ( .A1(n11438), .A2(n11439), .ZN(n11442) );
  INV_X1 U10368 ( .A(n11452), .ZN(n15017) );
  NAND2_X1 U10369 ( .A1(n11505), .A2(n15017), .ZN(n7986) );
  INV_X1 U10370 ( .A(n7987), .ZN(n7988) );
  XNOR2_X1 U10371 ( .A(n12715), .B(n15080), .ZN(n11338) );
  NAND2_X1 U10372 ( .A1(n11077), .A2(n15072), .ZN(n11336) );
  AND2_X1 U10373 ( .A1(n11338), .A2(n11336), .ZN(n11337) );
  AND2_X1 U10374 ( .A1(n11337), .A2(n11445), .ZN(n11441) );
  NAND2_X1 U10375 ( .A1(n11510), .A2(n12714), .ZN(n7989) );
  NAND2_X1 U10376 ( .A1(n11383), .A2(n11382), .ZN(n11381) );
  INV_X1 U10377 ( .A(n12713), .ZN(n11700) );
  OR2_X1 U10378 ( .A1(n14573), .A2(n11700), .ZN(n7990) );
  NAND2_X1 U10379 ( .A1(n11381), .A2(n7990), .ZN(n11597) );
  NAND2_X1 U10380 ( .A1(n14569), .A2(n11677), .ZN(n7991) );
  NAND2_X1 U10381 ( .A1(n11597), .A2(n7991), .ZN(n7993) );
  INV_X1 U10382 ( .A(n14569), .ZN(n11711) );
  NAND2_X1 U10383 ( .A1(n11711), .A2(n12712), .ZN(n7992) );
  NAND2_X1 U10384 ( .A1(n7993), .A2(n7992), .ZN(n11675) );
  NAND2_X1 U10385 ( .A1(n11675), .A2(n11678), .ZN(n7995) );
  NAND2_X1 U10386 ( .A1(n11879), .A2(n12711), .ZN(n7994) );
  AND2_X1 U10387 ( .A1(n12529), .A2(n12710), .ZN(n7997) );
  OR2_X1 U10388 ( .A1(n12529), .A2(n12710), .ZN(n7996) );
  INV_X1 U10389 ( .A(n12698), .ZN(n13024) );
  NAND2_X1 U10390 ( .A1(n12627), .A2(n13024), .ZN(n13016) );
  NAND2_X1 U10391 ( .A1(n13017), .A2(n13016), .ZN(n8000) );
  NAND2_X1 U10392 ( .A1(n13028), .A2(n13004), .ZN(n8002) );
  NAND2_X1 U10393 ( .A1(n12989), .A2(n8004), .ZN(n12972) );
  INV_X1 U10394 ( .A(n13005), .ZN(n12669) );
  OR2_X1 U10395 ( .A1(n13120), .A2(n12669), .ZN(n12973) );
  NAND2_X1 U10396 ( .A1(n12983), .A2(n12990), .ZN(n8005) );
  AND2_X1 U10397 ( .A1(n12973), .A2(n8005), .ZN(n8007) );
  INV_X1 U10398 ( .A(n8005), .ZN(n8006) );
  AND2_X1 U10399 ( .A1(n12605), .A2(n12976), .ZN(n8138) );
  NAND2_X1 U10400 ( .A1(n13112), .A2(n12950), .ZN(n8139) );
  NAND2_X1 U10401 ( .A1(n12940), .A2(n12709), .ZN(n8008) );
  NAND2_X1 U10402 ( .A1(n12918), .A2(n12924), .ZN(n12917) );
  NAND2_X1 U10403 ( .A1(n12905), .A2(n12904), .ZN(n12903) );
  NAND2_X1 U10404 ( .A1(n12903), .A2(n7423), .ZN(n12888) );
  NAND2_X1 U10405 ( .A1(n12885), .A2(n12891), .ZN(n8009) );
  INV_X1 U10406 ( .A(n8009), .ZN(n8010) );
  INV_X1 U10407 ( .A(n10521), .ZN(n8054) );
  NAND2_X1 U10408 ( .A1(n8054), .A2(n10305), .ZN(n8135) );
  NAND2_X1 U10409 ( .A1(n12848), .A2(n10818), .ZN(n8064) );
  INV_X1 U10410 ( .A(n9919), .ZN(n10040) );
  NAND2_X1 U10411 ( .A1(n8017), .A2(n8016), .ZN(n8019) );
  NAND2_X1 U10412 ( .A1(n8019), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8018) );
  MUX2_X1 U10413 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8018), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8021) );
  INV_X1 U10414 ( .A(n8019), .ZN(n8020) );
  NAND2_X1 U10415 ( .A1(n8020), .A2(n7468), .ZN(n8024) );
  NAND2_X1 U10416 ( .A1(n8021), .A2(n8024), .ZN(n11579) );
  INV_X1 U10417 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U10418 ( .A1(n12251), .A2(n8032), .ZN(n8033) );
  INV_X1 U10419 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9303) );
  NAND2_X1 U10420 ( .A1(n8034), .A2(n9303), .ZN(n8036) );
  NAND2_X1 U10421 ( .A1(n12251), .A2(n11579), .ZN(n8035) );
  XNOR2_X1 U10422 ( .A(n10027), .B(n9695), .ZN(n8051) );
  NOR2_X1 U10423 ( .A1(n11579), .A2(n8032), .ZN(n8037) );
  NAND2_X1 U10424 ( .A1(n6748), .A2(n8037), .ZN(n9908) );
  NAND2_X1 U10425 ( .A1(n6612), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8039) );
  NOR2_X1 U10426 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .ZN(
        n8043) );
  NOR4_X1 U10427 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n8042) );
  NOR4_X1 U10428 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8041) );
  NOR4_X1 U10429 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n8040) );
  NAND4_X1 U10430 ( .A1(n8043), .A2(n8042), .A3(n8041), .A4(n8040), .ZN(n8049)
         );
  NOR4_X1 U10431 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8047) );
  NOR4_X1 U10432 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_12__SCAN_IN), .ZN(n8046) );
  NOR4_X1 U10433 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8045) );
  NOR4_X1 U10434 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8044) );
  NAND4_X1 U10435 ( .A1(n8047), .A2(n8046), .A3(n8045), .A4(n8044), .ZN(n8048)
         );
  OAI21_X1 U10436 ( .B1(n8049), .B2(n8048), .A(n8034), .ZN(n8067) );
  AND2_X1 U10437 ( .A1(n9998), .A2(n8067), .ZN(n8050) );
  NAND2_X1 U10438 ( .A1(n8052), .A2(n8280), .ZN(n9693) );
  NAND2_X1 U10439 ( .A1(n8161), .A2(n10001), .ZN(n9907) );
  AND2_X1 U10440 ( .A1(n9693), .A2(n9907), .ZN(n8057) );
  OAI21_X1 U10441 ( .B1(n8054), .B2(n15079), .A(n8053), .ZN(n8055) );
  AOI21_X1 U10442 ( .B1(n8055), .B2(n8161), .A(n10001), .ZN(n8056) );
  INV_X1 U10443 ( .A(n9695), .ZN(n9692) );
  MUX2_X1 U10444 ( .A(n8057), .B(n8056), .S(n9692), .Z(n8058) );
  OR2_X1 U10445 ( .A1(n8072), .A2(n15104), .ZN(n8062) );
  INV_X1 U10446 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U10447 ( .A1(n8062), .A2(n8061), .ZN(P3_U3487) );
  INV_X1 U10448 ( .A(n10027), .ZN(n13132) );
  AND3_X1 U10449 ( .A1(n13132), .A2(n9695), .A3(n8067), .ZN(n9921) );
  NOR2_X1 U10450 ( .A1(n8161), .A2(n8280), .ZN(n9701) );
  NAND2_X1 U10451 ( .A1(n9998), .A2(n9701), .ZN(n9917) );
  NOR2_X1 U10452 ( .A1(n10026), .A2(n8064), .ZN(n9909) );
  NAND2_X1 U10453 ( .A1(n9998), .A2(n9909), .ZN(n8065) );
  NAND2_X1 U10454 ( .A1(n9917), .A2(n8065), .ZN(n8066) );
  NAND2_X1 U10455 ( .A1(n9921), .A2(n8066), .ZN(n8071) );
  NAND2_X1 U10456 ( .A1(n10027), .A2(n8067), .ZN(n8068) );
  INV_X1 U10457 ( .A(n9918), .ZN(n9902) );
  AND2_X1 U10458 ( .A1(n9998), .A2(n9906), .ZN(n8069) );
  NAND2_X1 U10459 ( .A1(n9902), .A2(n8069), .ZN(n8070) );
  OR2_X1 U10460 ( .A1(n8072), .A2(n15087), .ZN(n8076) );
  INV_X1 U10461 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8073) );
  INV_X1 U10462 ( .A(n8074), .ZN(n8075) );
  NAND2_X1 U10463 ( .A1(n8076), .A2(n8075), .ZN(P3_U3455) );
  AND2_X1 U10464 ( .A1(n8078), .A2(n8077), .ZN(n8297) );
  INV_X1 U10465 ( .A(n8298), .ZN(n8079) );
  INV_X1 U10466 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13808) );
  INV_X1 U10467 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14393) );
  AOI22_X1 U10468 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n13808), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n14393), .ZN(n8083) );
  XNOR2_X1 U10469 ( .A(n8116), .B(n8083), .ZN(n13136) );
  NAND2_X1 U10470 ( .A1(n13136), .A2(n7559), .ZN(n8085) );
  NAND2_X1 U10471 ( .A1(n8124), .A2(SI_29_), .ZN(n8084) );
  NAND2_X1 U10472 ( .A1(n8101), .A2(n12572), .ZN(n8127) );
  NAND2_X1 U10473 ( .A1(n8301), .A2(n8127), .ZN(n8089) );
  INV_X1 U10474 ( .A(n8089), .ZN(n8086) );
  INV_X1 U10475 ( .A(n12877), .ZN(n8087) );
  XNOR2_X1 U10476 ( .A(n8090), .B(n8089), .ZN(n8100) );
  NOR2_X1 U10477 ( .A1(n12877), .A2(n12964), .ZN(n8098) );
  INV_X1 U10478 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14585) );
  NAND2_X1 U10479 ( .A1(n8108), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U10480 ( .A1(n8107), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8091) );
  OAI211_X1 U10481 ( .C1(n7596), .C2(n14585), .A(n8092), .B(n8091), .ZN(n8093)
         );
  INV_X1 U10482 ( .A(n8093), .ZN(n8094) );
  NAND2_X1 U10483 ( .A1(n8095), .A2(P3_B_REG_SCAN_IN), .ZN(n8096) );
  NAND2_X1 U10484 ( .A1(n13022), .A2(n8096), .ZN(n12851) );
  NOR2_X1 U10485 ( .A1(n8129), .A2(n12851), .ZN(n8097) );
  OAI21_X1 U10486 ( .B1(n8100), .B2(n12960), .A(n8099), .ZN(n12859) );
  INV_X1 U10487 ( .A(n13129), .ZN(n8104) );
  INV_X1 U10488 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8102) );
  NOR2_X1 U10489 ( .A1(n15089), .A2(n8102), .ZN(n8103) );
  NAND2_X1 U10490 ( .A1(n8106), .A2(n8301), .ZN(n8133) );
  NAND2_X1 U10491 ( .A1(n8107), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n8112) );
  NAND2_X1 U10492 ( .A1(n8108), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8111) );
  NAND2_X1 U10493 ( .A1(n8109), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n8110) );
  AND3_X1 U10494 ( .A1(n8112), .A2(n8111), .A3(n8110), .ZN(n8113) );
  NAND2_X1 U10495 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n14393), .ZN(n8115) );
  INV_X1 U10496 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13805) );
  INV_X1 U10497 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U10498 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(
        P1_DATAO_REG_30__SCAN_IN), .B1(n13805), .B2(n12432), .ZN(n8117) );
  XNOR2_X1 U10499 ( .A(n8122), .B(n8117), .ZN(n11940) );
  NAND2_X1 U10500 ( .A1(n11940), .A2(n7559), .ZN(n8120) );
  NAND2_X1 U10501 ( .A1(n8118), .A2(SI_30_), .ZN(n8119) );
  NAND2_X1 U10502 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n13805), .ZN(n8121) );
  INV_X1 U10503 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13799) );
  INV_X1 U10504 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9352) );
  AOI22_X1 U10505 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n13799), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n9352), .ZN(n8123) );
  NAND2_X1 U10506 ( .A1(n8124), .A2(SI_31_), .ZN(n8125) );
  NAND2_X1 U10507 ( .A1(n14566), .A2(n8129), .ZN(n8128) );
  NAND2_X1 U10508 ( .A1(n8128), .A2(n8127), .ZN(n8162) );
  AOI211_X1 U10509 ( .C1(n12852), .C2(n14566), .A(n8306), .B(n8162), .ZN(n8132) );
  INV_X1 U10510 ( .A(n14566), .ZN(n12858) );
  INV_X1 U10511 ( .A(n8129), .ZN(n12707) );
  INV_X1 U10512 ( .A(n12852), .ZN(n12706) );
  NAND2_X1 U10513 ( .A1(n8136), .A2(n12706), .ZN(n8131) );
  INV_X1 U10514 ( .A(n8136), .ZN(n8137) );
  INV_X1 U10515 ( .A(n8308), .ZN(n8158) );
  INV_X1 U10516 ( .A(n12946), .ZN(n12952) );
  INV_X1 U10517 ( .A(n8138), .ZN(n8140) );
  NAND2_X1 U10518 ( .A1(n8140), .A2(n8139), .ZN(n12966) );
  OR2_X1 U10519 ( .A1(n7449), .A2(n8229), .ZN(n11598) );
  NOR2_X1 U10520 ( .A1(n11132), .A2(n10099), .ZN(n8142) );
  NAND4_X1 U10521 ( .A1(n8142), .A2(n8141), .A3(n10822), .A4(n8204), .ZN(n8147) );
  NAND2_X1 U10522 ( .A1(n12722), .A2(n10084), .ZN(n8165) );
  INV_X1 U10523 ( .A(n8165), .ZN(n8144) );
  NOR2_X1 U10524 ( .A1(n10303), .A2(n8144), .ZN(n9926) );
  INV_X1 U10525 ( .A(n10304), .ZN(n10307) );
  NAND4_X1 U10526 ( .A1(n9926), .A2(n10307), .A3(n10317), .A4(n11145), .ZN(
        n8146) );
  NOR3_X1 U10527 ( .A1(n8147), .A2(n8146), .A3(n11338), .ZN(n8148) );
  NAND4_X1 U10528 ( .A1(n8148), .A2(n11438), .A3(n6898), .A4(n11387), .ZN(
        n8149) );
  NOR3_X1 U10529 ( .A1(n11678), .A2(n11598), .A3(n8149), .ZN(n8150) );
  AND2_X1 U10530 ( .A1(n11758), .A2(n8150), .ZN(n8151) );
  AND4_X1 U10531 ( .A1(n13000), .A2(n11886), .A3(n6884), .A4(n8151), .ZN(n8152) );
  NAND4_X1 U10532 ( .A1(n12966), .A2(n12993), .A3(n7816), .A4(n8152), .ZN(
        n8153) );
  NOR2_X1 U10533 ( .A1(n12952), .A2(n8153), .ZN(n8154) );
  NAND4_X1 U10534 ( .A1(n12910), .A2(n7891), .A3(n8154), .A4(n8276), .ZN(n8155) );
  NOR2_X1 U10535 ( .A1(n12897), .A2(n8155), .ZN(n8156) );
  INV_X1 U10536 ( .A(n8301), .ZN(n8157) );
  XNOR2_X1 U10537 ( .A(n8159), .B(n12833), .ZN(n8160) );
  INV_X1 U10538 ( .A(n8161), .ZN(n8310) );
  INV_X1 U10539 ( .A(n8162), .ZN(n8305) );
  MUX2_X1 U10540 ( .A(n8164), .B(n8163), .S(n8280), .Z(n8275) );
  AOI21_X1 U10541 ( .B1(n8169), .B2(n10818), .A(n10571), .ZN(n8166) );
  MUX2_X1 U10542 ( .A(n10001), .B(n8166), .S(n8165), .Z(n8173) );
  NAND2_X1 U10543 ( .A1(n10303), .A2(n10571), .ZN(n8167) );
  NAND2_X1 U10544 ( .A1(n8167), .A2(n8168), .ZN(n8172) );
  MUX2_X1 U10545 ( .A(n8169), .B(n8168), .S(n10001), .Z(n8170) );
  OAI211_X1 U10546 ( .C1(n8173), .C2(n8172), .A(n8171), .B(n8170), .ZN(n8177)
         );
  NAND2_X1 U10547 ( .A1(n8184), .A2(n8174), .ZN(n8175) );
  NAND2_X1 U10548 ( .A1(n8175), .A2(n10001), .ZN(n8176) );
  NAND2_X1 U10549 ( .A1(n8177), .A2(n8176), .ZN(n8178) );
  NAND2_X1 U10550 ( .A1(n8178), .A2(n8180), .ZN(n8183) );
  NAND2_X1 U10551 ( .A1(n8180), .A2(n8179), .ZN(n8181) );
  NAND2_X1 U10552 ( .A1(n8181), .A2(n8280), .ZN(n8182) );
  NAND2_X1 U10553 ( .A1(n8183), .A2(n8182), .ZN(n8187) );
  NOR2_X1 U10554 ( .A1(n8184), .A2(n10001), .ZN(n8185) );
  NOR2_X1 U10555 ( .A1(n10456), .A2(n8185), .ZN(n8186) );
  NAND2_X1 U10556 ( .A1(n8187), .A2(n8186), .ZN(n8193) );
  NAND3_X1 U10557 ( .A1(n8193), .A2(n10822), .A3(n8188), .ZN(n8190) );
  NAND3_X1 U10558 ( .A1(n8190), .A2(n8189), .A3(n8197), .ZN(n8191) );
  NAND2_X1 U10559 ( .A1(n8191), .A2(n8195), .ZN(n8200) );
  NAND3_X1 U10560 ( .A1(n8193), .A2(n10822), .A3(n8192), .ZN(n8196) );
  NAND3_X1 U10561 ( .A1(n8196), .A2(n8195), .A3(n8194), .ZN(n8198) );
  NAND2_X1 U10562 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  MUX2_X1 U10563 ( .A(n8200), .B(n8199), .S(n10001), .Z(n8205) );
  MUX2_X1 U10564 ( .A(n8202), .B(n8201), .S(n10001), .Z(n8203) );
  OAI211_X1 U10565 ( .C1(n8205), .C2(n11132), .A(n8204), .B(n8203), .ZN(n8210)
         );
  INV_X1 U10566 ( .A(n11338), .ZN(n8209) );
  MUX2_X1 U10567 ( .A(n8207), .B(n8206), .S(n8280), .Z(n8208) );
  NAND3_X1 U10568 ( .A1(n8210), .A2(n8209), .A3(n8208), .ZN(n8223) );
  INV_X1 U10569 ( .A(n8211), .ZN(n8213) );
  MUX2_X1 U10570 ( .A(n8213), .B(n8212), .S(n10001), .Z(n8214) );
  NOR3_X1 U10571 ( .A1(n8214), .A2(n11318), .A3(n11445), .ZN(n8222) );
  INV_X1 U10572 ( .A(n11505), .ZN(n11509) );
  NAND2_X1 U10573 ( .A1(n11509), .A2(n15017), .ZN(n8216) );
  OAI211_X1 U10574 ( .C1(n11318), .C2(n8216), .A(n8225), .B(n8215), .ZN(n8220)
         );
  OAI211_X1 U10575 ( .C1(n11318), .C2(n8218), .A(n8217), .B(n8224), .ZN(n8219)
         );
  MUX2_X1 U10576 ( .A(n8220), .B(n8219), .S(n10001), .Z(n8221) );
  AOI21_X1 U10577 ( .B1(n8223), .B2(n8222), .A(n8221), .ZN(n8228) );
  INV_X1 U10578 ( .A(n11598), .ZN(n11600) );
  MUX2_X1 U10579 ( .A(n8225), .B(n8224), .S(n8280), .Z(n8226) );
  NAND2_X1 U10580 ( .A1(n11600), .A2(n8226), .ZN(n8227) );
  OR2_X1 U10581 ( .A1(n8228), .A2(n8227), .ZN(n8232) );
  AND2_X1 U10582 ( .A1(n8229), .A2(n8280), .ZN(n8230) );
  NOR2_X1 U10583 ( .A1(n11678), .A2(n8230), .ZN(n8231) );
  NAND2_X1 U10584 ( .A1(n8232), .A2(n8231), .ZN(n8239) );
  INV_X1 U10585 ( .A(n11758), .ZN(n11755) );
  AOI21_X1 U10586 ( .B1(n8239), .B2(n8233), .A(n11755), .ZN(n8237) );
  NAND2_X1 U10587 ( .A1(n8235), .A2(n8234), .ZN(n8236) );
  OAI21_X1 U10588 ( .B1(n8237), .B2(n8236), .A(n8280), .ZN(n8243) );
  OAI22_X1 U10589 ( .A1(n8239), .A2(n7449), .B1(n8280), .B2(n8238), .ZN(n8240)
         );
  NAND2_X1 U10590 ( .A1(n8240), .A2(n11758), .ZN(n8242) );
  INV_X1 U10591 ( .A(n8245), .ZN(n8241) );
  AOI21_X1 U10592 ( .B1(n8243), .B2(n8242), .A(n8241), .ZN(n8248) );
  AOI21_X1 U10593 ( .B1(n8245), .B2(n8244), .A(n8280), .ZN(n8247) );
  OR2_X1 U10594 ( .A1(n12698), .A2(n8280), .ZN(n8246) );
  OAI22_X1 U10595 ( .A1(n8248), .A2(n8247), .B1(n12627), .B2(n8246), .ZN(n8249) );
  NAND3_X1 U10596 ( .A1(n8249), .A2(n6884), .A3(n13000), .ZN(n8261) );
  INV_X1 U10597 ( .A(n8250), .ZN(n8251) );
  NAND2_X1 U10598 ( .A1(n13000), .A2(n8251), .ZN(n8252) );
  NAND3_X1 U10599 ( .A1(n8252), .A2(n8263), .A3(n8253), .ZN(n8258) );
  INV_X1 U10600 ( .A(n8253), .ZN(n8256) );
  OAI211_X1 U10601 ( .C1(n8256), .C2(n8255), .A(n8262), .B(n8254), .ZN(n8257)
         );
  MUX2_X1 U10602 ( .A(n8258), .B(n8257), .S(n10001), .Z(n8259) );
  INV_X1 U10603 ( .A(n8259), .ZN(n8260) );
  NAND2_X1 U10604 ( .A1(n8261), .A2(n8260), .ZN(n8265) );
  MUX2_X1 U10605 ( .A(n8263), .B(n8262), .S(n8280), .Z(n8264) );
  NAND3_X1 U10606 ( .A1(n8265), .A2(n7816), .A3(n8264), .ZN(n8269) );
  MUX2_X1 U10607 ( .A(n8267), .B(n8266), .S(n10001), .Z(n8268) );
  NAND3_X1 U10608 ( .A1(n8269), .A2(n12966), .A3(n8268), .ZN(n8273) );
  MUX2_X1 U10609 ( .A(n8271), .B(n8270), .S(n10001), .Z(n8272) );
  NAND3_X1 U10610 ( .A1(n8273), .A2(n12946), .A3(n8272), .ZN(n8274) );
  NAND3_X1 U10611 ( .A1(n8276), .A2(n8275), .A3(n8274), .ZN(n8278) );
  NAND3_X1 U10612 ( .A1(n12940), .A2(n12949), .A3(n10001), .ZN(n8277) );
  AND2_X1 U10613 ( .A1(n8278), .A2(n8277), .ZN(n8285) );
  INV_X1 U10614 ( .A(n8279), .ZN(n8283) );
  XNOR2_X1 U10615 ( .A(n8281), .B(n8280), .ZN(n8282) );
  OAI21_X1 U10616 ( .B1(n12924), .B2(n8283), .A(n8282), .ZN(n8284) );
  OAI211_X1 U10617 ( .C1(n8285), .C2(n12924), .A(n12910), .B(n8284), .ZN(n8289) );
  MUX2_X1 U10618 ( .A(n8287), .B(n8286), .S(n10001), .Z(n8288) );
  NAND2_X1 U10619 ( .A1(n8289), .A2(n8288), .ZN(n8293) );
  MUX2_X1 U10620 ( .A(n8291), .B(n8290), .S(n10001), .Z(n8292) );
  OAI21_X1 U10621 ( .B1(n8293), .B2(n12897), .A(n8292), .ZN(n8295) );
  NOR2_X1 U10622 ( .A1(n12891), .A2(n10001), .ZN(n8294) );
  AOI22_X1 U10623 ( .A1(n12881), .A2(n8295), .B1(n12885), .B2(n8294), .ZN(
        n8296) );
  OR2_X1 U10624 ( .A1(n12568), .A2(n8296), .ZN(n8303) );
  NAND2_X1 U10625 ( .A1(n8297), .A2(n10001), .ZN(n8299) );
  NAND2_X1 U10626 ( .A1(n8299), .A2(n8298), .ZN(n8300) );
  NAND2_X1 U10627 ( .A1(n8300), .A2(n8303), .ZN(n8302) );
  OAI211_X1 U10628 ( .C1(n10001), .C2(n8303), .A(n8302), .B(n8301), .ZN(n8304)
         );
  NAND2_X1 U10629 ( .A1(n8305), .A2(n8304), .ZN(n8307) );
  AOI21_X1 U10630 ( .B1(n8308), .B2(n8307), .A(n8306), .ZN(n8309) );
  MUX2_X1 U10631 ( .A(n8310), .B(n15023), .S(n8309), .Z(n8311) );
  OR2_X1 U10632 ( .A1(n10000), .A2(P3_U3151), .ZN(n10970) );
  INV_X1 U10633 ( .A(n10970), .ZN(n8313) );
  NOR3_X1 U10634 ( .A1(n9917), .A2(n12837), .A3(n12521), .ZN(n8315) );
  OAI21_X1 U10635 ( .B1(n10970), .B2(n10818), .A(P3_B_REG_SCAN_IN), .ZN(n8314)
         );
  OR2_X1 U10636 ( .A1(n8315), .A2(n8314), .ZN(n8316) );
  INV_X1 U10637 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9605) );
  INV_X1 U10638 ( .A(n8537), .ZN(n8319) );
  AND2_X1 U10639 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8320) );
  NAND2_X1 U10640 ( .A1(n9257), .A2(n8320), .ZN(n9190) );
  NAND2_X1 U10641 ( .A1(n8539), .A2(n9190), .ZN(n8543) );
  INV_X1 U10642 ( .A(SI_1_), .ZN(n9237) );
  NOR2_X1 U10643 ( .A1(n8321), .A2(n9237), .ZN(n8322) );
  INV_X1 U10644 ( .A(n8569), .ZN(n8324) );
  MUX2_X1 U10645 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8328), .Z(n8325) );
  XNOR2_X1 U10646 ( .A(n8325), .B(SI_2_), .ZN(n8568) );
  INV_X1 U10647 ( .A(n8568), .ZN(n8323) );
  NAND2_X1 U10648 ( .A1(n8324), .A2(n8323), .ZN(n8327) );
  NAND2_X1 U10649 ( .A1(n8325), .A2(SI_2_), .ZN(n8326) );
  MUX2_X1 U10650 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n8328), .Z(n8330) );
  XNOR2_X1 U10651 ( .A(n8330), .B(SI_3_), .ZN(n8586) );
  INV_X1 U10652 ( .A(n8586), .ZN(n8329) );
  NAND2_X1 U10653 ( .A1(n8587), .A2(n8329), .ZN(n8332) );
  NAND2_X1 U10654 ( .A1(n8330), .A2(SI_3_), .ZN(n8331) );
  NAND2_X2 U10655 ( .A1(n8332), .A2(n8331), .ZN(n8605) );
  XNOR2_X1 U10656 ( .A(n8335), .B(SI_4_), .ZN(n8604) );
  INV_X1 U10657 ( .A(n8604), .ZN(n8334) );
  NAND2_X1 U10658 ( .A1(n8335), .A2(SI_4_), .ZN(n8336) );
  MUX2_X1 U10659 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7149), .Z(n8338) );
  XNOR2_X1 U10660 ( .A(n8338), .B(SI_5_), .ZN(n8617) );
  INV_X1 U10661 ( .A(n8617), .ZN(n8337) );
  MUX2_X1 U10662 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9249), .Z(n8340) );
  XNOR2_X1 U10663 ( .A(n8340), .B(SI_6_), .ZN(n8640) );
  INV_X1 U10664 ( .A(n8640), .ZN(n8339) );
  NAND2_X1 U10665 ( .A1(n8641), .A2(n8339), .ZN(n8342) );
  NAND2_X1 U10666 ( .A1(n8340), .A2(SI_6_), .ZN(n8341) );
  XNOR2_X1 U10667 ( .A(n8344), .B(SI_7_), .ZN(n8668) );
  INV_X1 U10668 ( .A(n8668), .ZN(n8343) );
  NAND2_X1 U10669 ( .A1(n8344), .A2(SI_7_), .ZN(n8345) );
  MUX2_X1 U10670 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n12101), .Z(n8346) );
  XNOR2_X1 U10671 ( .A(n8346), .B(SI_8_), .ZN(n8685) );
  MUX2_X1 U10672 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n12101), .Z(n8348) );
  XNOR2_X1 U10673 ( .A(n8348), .B(SI_9_), .ZN(n8707) );
  INV_X1 U10674 ( .A(n8707), .ZN(n8347) );
  NAND2_X1 U10675 ( .A1(n8348), .A2(SI_9_), .ZN(n8349) );
  MUX2_X1 U10676 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n12101), .Z(n8351) );
  XNOR2_X1 U10677 ( .A(n8351), .B(SI_10_), .ZN(n8724) );
  INV_X1 U10678 ( .A(n8724), .ZN(n8350) );
  NAND2_X1 U10679 ( .A1(n8351), .A2(SI_10_), .ZN(n8352) );
  MUX2_X1 U10680 ( .A(n9348), .B(n9350), .S(n12101), .Z(n8354) );
  INV_X1 U10681 ( .A(n8354), .ZN(n8355) );
  NAND2_X1 U10682 ( .A1(n8355), .A2(SI_11_), .ZN(n8356) );
  NAND2_X1 U10683 ( .A1(n8357), .A2(n8356), .ZN(n8748) );
  MUX2_X1 U10684 ( .A(n9447), .B(n9444), .S(n12101), .Z(n8358) );
  INV_X1 U10685 ( .A(n8358), .ZN(n8359) );
  NAND2_X1 U10686 ( .A1(n8359), .A2(SI_12_), .ZN(n8360) );
  MUX2_X1 U10687 ( .A(n11215), .B(n9598), .S(n12101), .Z(n8362) );
  NAND2_X1 U10688 ( .A1(n8362), .A2(n9327), .ZN(n8365) );
  INV_X1 U10689 ( .A(n8362), .ZN(n8363) );
  NAND2_X1 U10690 ( .A1(n8363), .A2(SI_13_), .ZN(n8364) );
  INV_X1 U10691 ( .A(n8365), .ZN(n8366) );
  INV_X1 U10692 ( .A(SI_14_), .ZN(n9443) );
  MUX2_X1 U10693 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n12101), .Z(n8847) );
  MUX2_X1 U10694 ( .A(n10270), .B(n10272), .S(n12101), .Z(n8368) );
  INV_X1 U10695 ( .A(n8368), .ZN(n8369) );
  NAND2_X1 U10696 ( .A1(n8369), .A2(SI_15_), .ZN(n8370) );
  MUX2_X1 U10697 ( .A(n8373), .B(n10453), .S(n12101), .Z(n8374) );
  INV_X1 U10698 ( .A(n8374), .ZN(n8375) );
  NAND2_X1 U10699 ( .A1(n8375), .A2(SI_16_), .ZN(n8376) );
  MUX2_X1 U10700 ( .A(n10642), .B(n10644), .S(n12101), .Z(n8793) );
  INV_X1 U10701 ( .A(n8793), .ZN(n8379) );
  NAND2_X1 U10702 ( .A1(n8379), .A2(SI_17_), .ZN(n8380) );
  INV_X1 U10703 ( .A(SI_17_), .ZN(n9840) );
  NAND2_X1 U10704 ( .A1(n8793), .A2(n9840), .ZN(n8381) );
  MUX2_X1 U10705 ( .A(n10948), .B(n10949), .S(n12101), .Z(n8885) );
  INV_X1 U10706 ( .A(n8885), .ZN(n8382) );
  MUX2_X1 U10707 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n12101), .Z(n8384) );
  XNOR2_X1 U10708 ( .A(n8384), .B(SI_19_), .ZN(n8907) );
  NOR2_X1 U10709 ( .A1(n8885), .A2(n9971), .ZN(n8383) );
  INV_X1 U10710 ( .A(n8384), .ZN(n8385) );
  NAND2_X1 U10711 ( .A1(n8385), .A2(n10135), .ZN(n8386) );
  MUX2_X1 U10712 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n12101), .Z(n8939) );
  NAND2_X1 U10713 ( .A1(n8939), .A2(SI_20_), .ZN(n8388) );
  MUX2_X1 U10714 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9249), .Z(n8389) );
  NAND2_X1 U10715 ( .A1(n8389), .A2(SI_21_), .ZN(n8392) );
  OAI21_X1 U10716 ( .B1(SI_21_), .B2(n8389), .A(n8392), .ZN(n8940) );
  NOR2_X1 U10717 ( .A1(n8939), .A2(SI_20_), .ZN(n8390) );
  NOR2_X1 U10718 ( .A1(n8940), .A2(n8390), .ZN(n8391) );
  MUX2_X1 U10719 ( .A(n8395), .B(n11349), .S(n9249), .Z(n8957) );
  MUX2_X1 U10720 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n12101), .Z(n8397) );
  NAND2_X1 U10721 ( .A1(n8397), .A2(SI_23_), .ZN(n8399) );
  OAI21_X1 U10722 ( .B1(SI_23_), .B2(n8397), .A(n8399), .ZN(n8398) );
  INV_X1 U10723 ( .A(n8398), .ZN(n8978) );
  MUX2_X1 U10724 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n12101), .Z(n8400) );
  NAND2_X1 U10725 ( .A1(n8400), .A2(SI_24_), .ZN(n8402) );
  OAI21_X1 U10726 ( .B1(SI_24_), .B2(n8400), .A(n8402), .ZN(n8401) );
  INV_X1 U10727 ( .A(n8401), .ZN(n8999) );
  MUX2_X1 U10728 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9249), .Z(n8403) );
  XNOR2_X1 U10729 ( .A(n8403), .B(SI_25_), .ZN(n8526) );
  INV_X1 U10730 ( .A(n8403), .ZN(n8404) );
  INV_X1 U10731 ( .A(SI_25_), .ZN(n11580) );
  INV_X1 U10732 ( .A(SI_26_), .ZN(n12252) );
  NAND2_X1 U10733 ( .A1(n9031), .A2(n12252), .ZN(n8406) );
  MUX2_X1 U10734 ( .A(n12184), .B(n11909), .S(n9249), .Z(n9029) );
  INV_X1 U10735 ( .A(n9029), .ZN(n8405) );
  NAND2_X1 U10736 ( .A1(n8406), .A2(n8405), .ZN(n8408) );
  NAND2_X1 U10737 ( .A1(n9060), .A2(SI_27_), .ZN(n8409) );
  MUX2_X1 U10738 ( .A(n15230), .B(n13818), .S(n9249), .Z(n9057) );
  NAND2_X1 U10739 ( .A1(n8409), .A2(n9057), .ZN(n8412) );
  NAND2_X1 U10740 ( .A1(n8410), .A2(n13142), .ZN(n8411) );
  MUX2_X1 U10741 ( .A(n15143), .B(n13814), .S(n12101), .Z(n8413) );
  XNOR2_X1 U10742 ( .A(n8413), .B(SI_28_), .ZN(n8516) );
  INV_X1 U10743 ( .A(SI_28_), .ZN(n12522) );
  NAND2_X1 U10744 ( .A1(n8413), .A2(n12522), .ZN(n8414) );
  MUX2_X1 U10745 ( .A(n14393), .B(n13808), .S(n12101), .Z(n8416) );
  XNOR2_X1 U10746 ( .A(n8416), .B(SI_29_), .ZN(n8495) );
  INV_X1 U10747 ( .A(SI_29_), .ZN(n13139) );
  NAND2_X1 U10748 ( .A1(n8416), .A2(n13139), .ZN(n8417) );
  MUX2_X1 U10749 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9249), .Z(n8497) );
  XNOR2_X1 U10750 ( .A(n8497), .B(SI_30_), .ZN(n8499) );
  INV_X1 U10751 ( .A(n8499), .ZN(n8419) );
  NOR2_X1 U10752 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8422) );
  NAND4_X1 U10753 ( .A1(n8422), .A2(n8421), .A3(n8420), .A4(n8449), .ZN(n8455)
         );
  NAND4_X1 U10754 ( .A1(n8465), .A2(n8459), .A3(n8424), .A4(n8423), .ZN(n8425)
         );
  NOR2_X2 U10755 ( .A1(n8455), .A2(n8425), .ZN(n9093) );
  NOR2_X2 U10756 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8570) );
  NAND2_X1 U10757 ( .A1(n8570), .A2(n8429), .ZN(n8584) );
  NOR2_X1 U10758 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8431) );
  NAND2_X1 U10759 ( .A1(n8441), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8439) );
  MUX2_X1 U10760 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8442), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n8443) );
  NAND2_X1 U10761 ( .A1(n12431), .A2(n9061), .ZN(n8446) );
  NAND2_X1 U10762 ( .A1(n9062), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10763 ( .A1(n8831), .A2(n8449), .ZN(n8450) );
  INV_X1 U10764 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8452) );
  XNOR2_X1 U10765 ( .A(n8453), .B(n8452), .ZN(n8477) );
  INV_X1 U10766 ( .A(n8455), .ZN(n8456) );
  INV_X1 U10767 ( .A(n8460), .ZN(n8457) );
  NAND2_X1 U10768 ( .A1(n8457), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8458) );
  MUX2_X1 U10769 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8458), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8461) );
  INV_X1 U10770 ( .A(n8466), .ZN(n8463) );
  NAND2_X1 U10771 ( .A1(n8890), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U10772 ( .A1(n8463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8464) );
  MUX2_X1 U10773 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8464), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n8467) );
  INV_X1 U10774 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U10775 ( .A1(n8469), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8470) );
  AND2_X2 U10776 ( .A1(n8471), .A2(n7418), .ZN(n8482) );
  INV_X1 U10777 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n13761) );
  NAND2_X1 U10778 ( .A1(n8530), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8474) );
  AND2_X4 U10779 ( .A1(n8482), .A2(n13804), .ZN(n8562) );
  NAND2_X1 U10780 ( .A1(n8562), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8473) );
  OAI211_X1 U10781 ( .C1(n9023), .C2(n13761), .A(n8474), .B(n8473), .ZN(n13337) );
  INV_X1 U10782 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13757) );
  NAND2_X1 U10783 ( .A1(n8530), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U10784 ( .A1(n8562), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8475) );
  OAI211_X1 U10785 ( .C1(n9023), .C2(n13757), .A(n8476), .B(n8475), .ZN(n13404) );
  NAND2_X1 U10786 ( .A1(n8648), .A2(n13404), .ZN(n8506) );
  AND2_X1 U10787 ( .A1(n9710), .A2(n9101), .ZN(n9720) );
  AOI21_X1 U10788 ( .B1(n9720), .B2(n6485), .A(n11111), .ZN(n8478) );
  NAND3_X1 U10789 ( .A1(n8506), .A2(n8478), .A3(n9751), .ZN(n8479) );
  AOI22_X1 U10790 ( .A1(n13411), .A2(n8731), .B1(n13337), .B2(n8479), .ZN(
        n9078) );
  MUX2_X1 U10791 ( .A(n13337), .B(n13411), .S(n9065), .Z(n9079) );
  NAND2_X1 U10792 ( .A1(n8562), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8494) );
  INV_X1 U10793 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8480) );
  OR2_X1 U10794 ( .A1(n9023), .A2(n8480), .ZN(n8493) );
  AND2_X2 U10795 ( .A1(n8482), .A2(n8481), .ZN(n8563) );
  INV_X4 U10796 ( .A(n8563), .ZN(n9051) );
  NAND2_X1 U10797 ( .A1(n8598), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U10798 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n8483) );
  NOR2_X1 U10799 ( .A1(n8659), .A2(n8483), .ZN(n8660) );
  NAND2_X1 U10800 ( .A1(n8699), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8741) );
  INV_X1 U10801 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8740) );
  INV_X1 U10802 ( .A(n8778), .ZN(n8485) );
  AND2_X1 U10803 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n8484) );
  NAND2_X1 U10804 ( .A1(n8485), .A2(n8484), .ZN(n8840) );
  NAND2_X1 U10805 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n8486) );
  INV_X1 U10806 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13237) );
  NAND2_X1 U10807 ( .A1(n8970), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8992) );
  INV_X1 U10808 ( .A(n8992), .ZN(n8487) );
  NAND2_X1 U10809 ( .A1(n8487), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n9020) );
  INV_X1 U10810 ( .A(n9020), .ZN(n8489) );
  AND2_X1 U10811 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8488) );
  NAND2_X1 U10812 ( .A1(n8489), .A2(n8488), .ZN(n9048) );
  INV_X1 U10813 ( .A(n9048), .ZN(n8490) );
  NAND2_X1 U10814 ( .A1(n8490), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9050) );
  INV_X1 U10815 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13227) );
  OR2_X1 U10816 ( .A1(n9051), .A2(n11995), .ZN(n8492) );
  INV_X1 U10817 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n11996) );
  OR2_X1 U10818 ( .A1(n9046), .A2(n11996), .ZN(n8491) );
  AND4_X1 U10819 ( .A1(n8494), .A2(n8493), .A3(n8492), .A4(n8491), .ZN(n13228)
         );
  MUX2_X1 U10820 ( .A(n13228), .B(n11994), .S(n8754), .Z(n8509) );
  OAI22_X1 U10821 ( .A1(n9078), .A2(n9079), .B1(n8509), .B2(n8508), .ZN(n9070)
         );
  NAND2_X1 U10822 ( .A1(n8497), .A2(SI_30_), .ZN(n8498) );
  MUX2_X1 U10823 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n12101), .Z(n8501) );
  XNOR2_X1 U10824 ( .A(n8501), .B(SI_31_), .ZN(n8502) );
  NAND2_X1 U10825 ( .A1(n9062), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8504) );
  MUX2_X1 U10826 ( .A(n8506), .B(n13404), .S(n8507), .Z(n9069) );
  XNOR2_X1 U10827 ( .A(n8507), .B(n13404), .ZN(n9122) );
  INV_X1 U10828 ( .A(n9122), .ZN(n8521) );
  NAND2_X1 U10829 ( .A1(n8509), .A2(n8508), .ZN(n9043) );
  INV_X1 U10830 ( .A(n9043), .ZN(n8520) );
  NAND2_X1 U10831 ( .A1(n8562), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8515) );
  INV_X1 U10832 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8510) );
  OR2_X1 U10833 ( .A1(n9023), .A2(n8510), .ZN(n8514) );
  NAND2_X1 U10834 ( .A1(n9050), .A2(n13227), .ZN(n8511) );
  NAND2_X1 U10835 ( .A1(n11995), .A2(n8511), .ZN(n13419) );
  OR2_X1 U10836 ( .A1(n9051), .A2(n13419), .ZN(n8513) );
  INV_X1 U10837 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13420) );
  OR2_X1 U10838 ( .A1(n9046), .A2(n13420), .ZN(n8512) );
  NAND2_X1 U10839 ( .A1(n13811), .A2(n8546), .ZN(n8519) );
  NAND2_X1 U10840 ( .A1(n9062), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8518) );
  MUX2_X1 U10841 ( .A(n13436), .B(n13418), .S(n8731), .Z(n9041) );
  MUX2_X1 U10842 ( .A(n13338), .B(n13680), .S(n8648), .Z(n9040) );
  NOR4_X1 U10843 ( .A1(n8521), .A2(n8520), .A3(n9041), .A4(n9040), .ZN(n9068)
         );
  NAND2_X1 U10844 ( .A1(n8562), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8525) );
  INV_X1 U10845 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n13772) );
  OR2_X1 U10846 ( .A1(n9023), .A2(n13772), .ZN(n8524) );
  INV_X1 U10847 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n13248) );
  XNOR2_X1 U10848 ( .A(n9020), .B(n13248), .ZN(n13476) );
  OR2_X1 U10849 ( .A1(n9051), .A2(n13476), .ZN(n8523) );
  INV_X1 U10850 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13477) );
  OR2_X1 U10851 ( .A1(n9046), .A2(n13477), .ZN(n8522) );
  XNOR2_X1 U10852 ( .A(n8527), .B(n8526), .ZN(n12162) );
  NAND2_X1 U10853 ( .A1(n12162), .A2(n9061), .ZN(n8529) );
  NAND2_X1 U10854 ( .A1(n9062), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8528) );
  AND2_X2 U10855 ( .A1(n8529), .A2(n8528), .ZN(n13773) );
  MUX2_X1 U10856 ( .A(n13279), .B(n13773), .S(n8754), .Z(n9015) );
  INV_X1 U10857 ( .A(n9015), .ZN(n9019) );
  INV_X1 U10858 ( .A(n8589), .ZN(n8530) );
  NAND2_X1 U10859 ( .A1(n8563), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U10860 ( .A1(n8562), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8533) );
  INV_X1 U10861 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8531) );
  OR2_X1 U10862 ( .A1(n8839), .A2(n8531), .ZN(n8532) );
  NAND2_X1 U10863 ( .A1(n8537), .A2(n8536), .ZN(n8538) );
  NAND2_X1 U10864 ( .A1(n8539), .A2(n8538), .ZN(n13820) );
  MUX2_X1 U10865 ( .A(n9459), .B(n13820), .S(n9098), .Z(n9831) );
  XNOR2_X1 U10866 ( .A(n9821), .B(n8648), .ZN(n8542) );
  INV_X1 U10867 ( .A(n9831), .ZN(n10060) );
  NAND2_X1 U10868 ( .A1(n8540), .A2(n10060), .ZN(n9832) );
  NAND2_X1 U10869 ( .A1(n9832), .A2(n9791), .ZN(n8541) );
  NAND2_X1 U10870 ( .A1(n8542), .A2(n8541), .ZN(n8557) );
  XNOR2_X1 U10871 ( .A(n8544), .B(n8543), .ZN(n9604) );
  INV_X1 U10872 ( .A(n9604), .ZN(n8545) );
  INV_X1 U10873 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n8548) );
  OR2_X1 U10874 ( .A1(n8589), .A2(n8548), .ZN(n8553) );
  INV_X1 U10875 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n8549) );
  OR2_X1 U10876 ( .A1(n8839), .A2(n8549), .ZN(n8552) );
  NAND2_X1 U10877 ( .A1(n8563), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U10878 ( .A1(n8557), .A2(n8556), .ZN(n8555) );
  MUX2_X1 U10879 ( .A(n13359), .B(n6481), .S(n8648), .Z(n8554) );
  NAND2_X1 U10880 ( .A1(n8555), .A2(n8554), .ZN(n8561) );
  INV_X1 U10881 ( .A(n8556), .ZN(n8559) );
  INV_X1 U10882 ( .A(n8557), .ZN(n8558) );
  NAND2_X1 U10883 ( .A1(n8559), .A2(n8558), .ZN(n8560) );
  NAND2_X1 U10884 ( .A1(n8562), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8567) );
  INV_X1 U10885 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8564) );
  OR2_X1 U10886 ( .A1(n8839), .A2(n8564), .ZN(n8566) );
  OR2_X1 U10887 ( .A1(n8589), .A2(n10465), .ZN(n8565) );
  XNOR2_X1 U10888 ( .A(n8569), .B(n8568), .ZN(n9641) );
  NAND2_X1 U10889 ( .A1(n9062), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8574) );
  INV_X1 U10890 ( .A(n8570), .ZN(n8571) );
  NAND2_X1 U10891 ( .A1(n8571), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8572) );
  XNOR2_X1 U10892 ( .A(n8572), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U10893 ( .A1(n8909), .A2(n9461), .ZN(n8573) );
  MUX2_X1 U10895 ( .A(n13358), .B(n10065), .S(n8648), .Z(n8579) );
  NAND2_X1 U10896 ( .A1(n8578), .A2(n8579), .ZN(n8577) );
  MUX2_X1 U10897 ( .A(n10065), .B(n13358), .S(n8648), .Z(n8576) );
  NAND2_X1 U10898 ( .A1(n8577), .A2(n8576), .ZN(n8583) );
  INV_X1 U10899 ( .A(n8578), .ZN(n8581) );
  INV_X1 U10900 ( .A(n8579), .ZN(n8580) );
  NAND2_X1 U10901 ( .A1(n8581), .A2(n8580), .ZN(n8582) );
  NAND2_X1 U10902 ( .A1(n8583), .A2(n8582), .ZN(n8595) );
  NAND2_X1 U10903 ( .A1(n8584), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8585) );
  XNOR2_X1 U10904 ( .A(n8585), .B(n6996), .ZN(n9546) );
  XNOR2_X1 U10905 ( .A(n8587), .B(n8586), .ZN(n9754) );
  NAND2_X1 U10906 ( .A1(n8562), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8593) );
  OR2_X1 U10907 ( .A1(n9051), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8592) );
  INV_X1 U10908 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8588) );
  OR2_X1 U10909 ( .A1(n8839), .A2(n8588), .ZN(n8591) );
  INV_X1 U10910 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n13653) );
  OR2_X1 U10911 ( .A1(n8589), .A2(n13653), .ZN(n8590) );
  MUX2_X1 U10912 ( .A(n9108), .B(n13357), .S(n8648), .Z(n8596) );
  MUX2_X1 U10913 ( .A(n13357), .B(n9108), .S(n8648), .Z(n8594) );
  INV_X1 U10914 ( .A(n8596), .ZN(n8597) );
  NAND2_X1 U10915 ( .A1(n8562), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n8603) );
  INV_X1 U10916 ( .A(n8598), .ZN(n8625) );
  OAI21_X1 U10917 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n8625), .ZN(n10432) );
  OR2_X1 U10918 ( .A1(n9051), .A2(n10432), .ZN(n8602) );
  INV_X1 U10919 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8599) );
  OR2_X1 U10920 ( .A1(n8839), .A2(n8599), .ZN(n8601) );
  INV_X1 U10921 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10349) );
  OR2_X1 U10922 ( .A1(n8589), .A2(n10349), .ZN(n8600) );
  NAND4_X1 U10923 ( .A1(n8603), .A2(n8602), .A3(n8601), .A4(n8600), .ZN(n13356) );
  XNOR2_X1 U10924 ( .A(n8604), .B(n8605), .ZN(n9929) );
  NAND2_X1 U10925 ( .A1(n9929), .A2(n9061), .ZN(n8608) );
  NAND2_X1 U10926 ( .A1(n8619), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8606) );
  XNOR2_X1 U10927 ( .A(n8606), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9463) );
  AOI22_X1 U10928 ( .A1(n9062), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8909), .B2(
        n9463), .ZN(n8607) );
  MUX2_X1 U10929 ( .A(n13356), .B(n10433), .S(n9065), .Z(n8612) );
  MUX2_X1 U10930 ( .A(n10433), .B(n13356), .S(n9065), .Z(n8609) );
  NAND2_X1 U10931 ( .A1(n8610), .A2(n8609), .ZN(n8616) );
  INV_X1 U10932 ( .A(n8611), .ZN(n8614) );
  INV_X1 U10933 ( .A(n8612), .ZN(n8613) );
  NAND2_X1 U10934 ( .A1(n8614), .A2(n8613), .ZN(n8615) );
  XNOR2_X1 U10935 ( .A(n8618), .B(n8617), .ZN(n10587) );
  NAND2_X1 U10936 ( .A1(n10587), .A2(n9061), .ZN(n8623) );
  INV_X1 U10937 ( .A(n8643), .ZN(n8620) );
  NAND2_X1 U10938 ( .A1(n8620), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8621) );
  XNOR2_X1 U10939 ( .A(n8621), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9550) );
  AOI22_X1 U10940 ( .A1(n9062), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8909), .B2(
        n9550), .ZN(n8622) );
  NAND2_X1 U10941 ( .A1(n8623), .A2(n8622), .ZN(n14932) );
  NAND2_X1 U10942 ( .A1(n8562), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8631) );
  INV_X1 U10943 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8624) );
  NAND2_X1 U10944 ( .A1(n8625), .A2(n8624), .ZN(n8626) );
  NAND2_X1 U10945 ( .A1(n8659), .A2(n8626), .ZN(n10579) );
  OR2_X1 U10946 ( .A1(n9051), .A2(n10579), .ZN(n8630) );
  INV_X1 U10947 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n8627) );
  OR2_X1 U10948 ( .A1(n9023), .A2(n8627), .ZN(n8629) );
  INV_X1 U10949 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10369) );
  OR2_X1 U10950 ( .A1(n9046), .A2(n10369), .ZN(n8628) );
  NAND4_X1 U10951 ( .A1(n8631), .A2(n8630), .A3(n8629), .A4(n8628), .ZN(n13355) );
  MUX2_X1 U10952 ( .A(n14932), .B(n13355), .S(n9065), .Z(n8633) );
  MUX2_X1 U10953 ( .A(n13355), .B(n14932), .S(n9065), .Z(n8632) );
  INV_X1 U10954 ( .A(n8633), .ZN(n8634) );
  NAND2_X1 U10955 ( .A1(n8562), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8639) );
  INV_X1 U10956 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8658) );
  XNOR2_X1 U10957 ( .A(n8659), .B(n8658), .ZN(n10719) );
  OR2_X1 U10958 ( .A1(n9051), .A2(n10719), .ZN(n8638) );
  INV_X1 U10959 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8635) );
  OR2_X1 U10960 ( .A1(n9023), .A2(n8635), .ZN(n8637) );
  INV_X1 U10961 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10390) );
  OR2_X1 U10962 ( .A1(n9046), .A2(n10390), .ZN(n8636) );
  NAND4_X1 U10963 ( .A1(n8639), .A2(n8638), .A3(n8637), .A4(n8636), .ZN(n13354) );
  XNOR2_X1 U10964 ( .A(n8641), .B(n8640), .ZN(n10592) );
  NAND2_X1 U10965 ( .A1(n10592), .A2(n9061), .ZN(n8647) );
  INV_X1 U10966 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8642) );
  INV_X1 U10967 ( .A(n8670), .ZN(n8644) );
  NAND2_X1 U10968 ( .A1(n8644), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8645) );
  XNOR2_X1 U10969 ( .A(n8645), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9569) );
  AOI22_X1 U10970 ( .A1(n9062), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8909), .B2(
        n9569), .ZN(n8646) );
  NAND2_X1 U10971 ( .A1(n8647), .A2(n8646), .ZN(n14938) );
  MUX2_X1 U10972 ( .A(n13354), .B(n14938), .S(n9065), .Z(n8652) );
  NAND2_X1 U10973 ( .A1(n8651), .A2(n8652), .ZN(n8650) );
  MUX2_X1 U10974 ( .A(n13354), .B(n14938), .S(n8731), .Z(n8649) );
  NAND2_X1 U10975 ( .A1(n8650), .A2(n8649), .ZN(n8656) );
  INV_X1 U10976 ( .A(n8651), .ZN(n8654) );
  INV_X1 U10977 ( .A(n8652), .ZN(n8653) );
  NAND2_X1 U10978 ( .A1(n8654), .A2(n8653), .ZN(n8655) );
  NAND2_X1 U10979 ( .A1(n8562), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8667) );
  INV_X1 U10980 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8657) );
  OAI21_X1 U10981 ( .B1(n8659), .B2(n8658), .A(n8657), .ZN(n8661) );
  INV_X1 U10982 ( .A(n8660), .ZN(n8678) );
  NAND2_X1 U10983 ( .A1(n8661), .A2(n8678), .ZN(n10800) );
  OR2_X1 U10984 ( .A1(n9051), .A2(n10800), .ZN(n8666) );
  INV_X1 U10985 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8662) );
  OR2_X1 U10986 ( .A1(n9023), .A2(n8662), .ZN(n8665) );
  INV_X1 U10987 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8663) );
  OR2_X1 U10988 ( .A1(n9046), .A2(n8663), .ZN(n8664) );
  NAND4_X1 U10989 ( .A1(n8667), .A2(n8666), .A3(n8665), .A4(n8664), .ZN(n13353) );
  XNOR2_X1 U10990 ( .A(n8669), .B(n8668), .ZN(n10604) );
  NAND2_X1 U10991 ( .A1(n10604), .A2(n9061), .ZN(n8673) );
  NAND2_X1 U10992 ( .A1(n8670), .A2(n6998), .ZN(n8687) );
  NAND2_X1 U10993 ( .A1(n8687), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8671) );
  XNOR2_X1 U10994 ( .A(n8671), .B(P2_IR_REG_7__SCAN_IN), .ZN(n9850) );
  AOI22_X1 U10995 ( .A1(n9062), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8909), .B2(
        n9850), .ZN(n8672) );
  NAND2_X1 U10996 ( .A1(n8673), .A2(n8672), .ZN(n10804) );
  MUX2_X1 U10997 ( .A(n13353), .B(n10804), .S(n8731), .Z(n8675) );
  MUX2_X1 U10998 ( .A(n13353), .B(n10804), .S(n9065), .Z(n8674) );
  INV_X1 U10999 ( .A(n8675), .ZN(n8676) );
  NAND2_X1 U11000 ( .A1(n8562), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n8684) );
  INV_X1 U11001 ( .A(n8677), .ZN(n8700) );
  INV_X1 U11002 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10927) );
  NAND2_X1 U11003 ( .A1(n8678), .A2(n10927), .ZN(n8679) );
  NAND2_X1 U11004 ( .A1(n8700), .A2(n8679), .ZN(n10928) );
  OR2_X1 U11005 ( .A1(n9051), .A2(n10928), .ZN(n8683) );
  INV_X1 U11006 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8680) );
  OR2_X1 U11007 ( .A1(n9023), .A2(n8680), .ZN(n8682) );
  INV_X1 U11008 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10742) );
  OR2_X1 U11009 ( .A1(n9046), .A2(n10742), .ZN(n8681) );
  NAND4_X1 U11010 ( .A1(n8684), .A2(n8683), .A3(n8682), .A4(n8681), .ZN(n13352) );
  XNOR2_X1 U11011 ( .A(n8686), .B(n8685), .ZN(n10833) );
  NAND2_X1 U11012 ( .A1(n10833), .A2(n9061), .ZN(n8690) );
  NAND2_X1 U11013 ( .A1(n8709), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8688) );
  XNOR2_X1 U11014 ( .A(n8688), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U11015 ( .A1(n9062), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n8909), .B2(
        n10126), .ZN(n8689) );
  NAND2_X1 U11016 ( .A1(n8690), .A2(n8689), .ZN(n10954) );
  MUX2_X1 U11017 ( .A(n13352), .B(n10954), .S(n9065), .Z(n8694) );
  NAND2_X1 U11018 ( .A1(n8693), .A2(n8694), .ZN(n8692) );
  MUX2_X1 U11019 ( .A(n13352), .B(n10954), .S(n8731), .Z(n8691) );
  NAND2_X1 U11020 ( .A1(n8692), .A2(n8691), .ZN(n8698) );
  INV_X1 U11021 ( .A(n8693), .ZN(n8696) );
  INV_X1 U11022 ( .A(n8694), .ZN(n8695) );
  NAND2_X1 U11023 ( .A1(n8696), .A2(n8695), .ZN(n8697) );
  NAND2_X1 U11024 ( .A1(n8562), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8706) );
  INV_X1 U11025 ( .A(n8699), .ZN(n8717) );
  INV_X1 U11026 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11038) );
  NAND2_X1 U11027 ( .A1(n8700), .A2(n11038), .ZN(n8701) );
  NAND2_X1 U11028 ( .A1(n8717), .A2(n8701), .ZN(n11039) );
  OR2_X1 U11029 ( .A1(n9051), .A2(n11039), .ZN(n8705) );
  INV_X1 U11030 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n8702) );
  OR2_X1 U11031 ( .A1(n9023), .A2(n8702), .ZN(n8704) );
  INV_X1 U11032 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10960) );
  OR2_X1 U11033 ( .A1(n9046), .A2(n10960), .ZN(n8703) );
  NAND4_X1 U11034 ( .A1(n8706), .A2(n8705), .A3(n8704), .A4(n8703), .ZN(n13351) );
  XNOR2_X1 U11035 ( .A(n8708), .B(n8707), .ZN(n10839) );
  NAND2_X1 U11036 ( .A1(n10839), .A2(n9061), .ZN(n8713) );
  INV_X1 U11037 ( .A(n8727), .ZN(n8710) );
  NAND2_X1 U11038 ( .A1(n8710), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8711) );
  XNOR2_X1 U11039 ( .A(n8711), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U11040 ( .A1(n9062), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8909), .B2(
        n10664), .ZN(n8712) );
  MUX2_X1 U11041 ( .A(n13351), .B(n11100), .S(n8731), .Z(n8715) );
  MUX2_X1 U11042 ( .A(n13351), .B(n11100), .S(n9065), .Z(n8714) );
  NAND2_X1 U11043 ( .A1(n8562), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8723) );
  INV_X1 U11044 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U11045 ( .A1(n8717), .A2(n8716), .ZN(n8718) );
  NAND2_X1 U11046 ( .A1(n8741), .A2(n8718), .ZN(n11201) );
  OR2_X1 U11047 ( .A1(n9051), .A2(n11201), .ZN(n8722) );
  INV_X1 U11048 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n8719) );
  OR2_X1 U11049 ( .A1(n9023), .A2(n8719), .ZN(n8721) );
  INV_X1 U11050 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n11407) );
  OR2_X1 U11051 ( .A1(n9046), .A2(n11407), .ZN(n8720) );
  NAND4_X1 U11052 ( .A1(n8723), .A2(n8722), .A3(n8721), .A4(n8720), .ZN(n13350) );
  NAND2_X1 U11053 ( .A1(n10884), .A2(n9061), .ZN(n8730) );
  INV_X1 U11054 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8726) );
  NAND2_X1 U11055 ( .A1(n8727), .A2(n8726), .ZN(n8750) );
  NAND2_X1 U11056 ( .A1(n8750), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8728) );
  XNOR2_X1 U11057 ( .A(n8728), .B(P2_IR_REG_10__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U11058 ( .A1(n8909), .A2(n11395), .B1(n9062), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U11059 ( .A1(n8730), .A2(n8729), .ZN(n11189) );
  MUX2_X1 U11060 ( .A(n13350), .B(n11189), .S(n9065), .Z(n8735) );
  NAND2_X1 U11061 ( .A1(n8734), .A2(n8735), .ZN(n8733) );
  MUX2_X1 U11062 ( .A(n13350), .B(n11189), .S(n8731), .Z(n8732) );
  NAND2_X1 U11063 ( .A1(n8733), .A2(n8732), .ZN(n8739) );
  INV_X1 U11064 ( .A(n8734), .ZN(n8737) );
  INV_X1 U11065 ( .A(n8735), .ZN(n8736) );
  NAND2_X1 U11066 ( .A1(n8737), .A2(n8736), .ZN(n8738) );
  NAND2_X1 U11067 ( .A1(n8739), .A2(n8738), .ZN(n8756) );
  NAND2_X1 U11068 ( .A1(n8562), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U11069 ( .A1(n8741), .A2(n8740), .ZN(n8742) );
  NAND2_X1 U11070 ( .A1(n8778), .A2(n8742), .ZN(n11307) );
  OR2_X1 U11071 ( .A1(n9051), .A2(n11307), .ZN(n8746) );
  INV_X1 U11072 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8743) );
  OR2_X1 U11073 ( .A1(n9023), .A2(n8743), .ZN(n8745) );
  INV_X1 U11074 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11165) );
  OR2_X1 U11075 ( .A1(n9046), .A2(n11165), .ZN(n8744) );
  NAND4_X1 U11076 ( .A1(n8747), .A2(n8746), .A3(n8745), .A4(n8744), .ZN(n13349) );
  NAND2_X1 U11077 ( .A1(n10976), .A2(n9061), .ZN(n8753) );
  OAI21_X1 U11078 ( .B1(n8750), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8751) );
  XNOR2_X1 U11079 ( .A(n8751), .B(P2_IR_REG_11__SCAN_IN), .ZN(n14859) );
  AOI22_X1 U11080 ( .A1(n14859), .A2(n8909), .B1(n9062), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8752) );
  MUX2_X1 U11081 ( .A(n13349), .B(n11310), .S(n8754), .Z(n8757) );
  MUX2_X1 U11082 ( .A(n13349), .B(n11310), .S(n9065), .Z(n8755) );
  INV_X1 U11083 ( .A(n8757), .ZN(n8758) );
  NAND2_X1 U11084 ( .A1(n8562), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8763) );
  INV_X1 U11085 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8777) );
  XNOR2_X1 U11086 ( .A(n8778), .B(n8777), .ZN(n14815) );
  OR2_X1 U11087 ( .A1(n9051), .A2(n14815), .ZN(n8762) );
  INV_X1 U11088 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8759) );
  OR2_X1 U11089 ( .A1(n9023), .A2(n8759), .ZN(n8761) );
  INV_X1 U11090 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11181) );
  OR2_X1 U11091 ( .A1(n9046), .A2(n11181), .ZN(n8760) );
  NAND4_X1 U11092 ( .A1(n8763), .A2(n8762), .A3(n8761), .A4(n8760), .ZN(n13348) );
  XNOR2_X1 U11093 ( .A(n8764), .B(n7447), .ZN(n11210) );
  NAND2_X1 U11094 ( .A1(n11210), .A2(n9061), .ZN(n8768) );
  NAND2_X1 U11095 ( .A1(n8765), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8766) );
  XNOR2_X1 U11096 ( .A(n8766), .B(P2_IR_REG_12__SCAN_IN), .ZN(n14869) );
  AOI22_X1 U11097 ( .A1(n9062), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8909), 
        .B2(n14869), .ZN(n8767) );
  MUX2_X1 U11098 ( .A(n13348), .B(n14813), .S(n9065), .Z(n8772) );
  MUX2_X1 U11099 ( .A(n13348), .B(n14813), .S(n8731), .Z(n8769) );
  NAND2_X1 U11100 ( .A1(n8770), .A2(n8769), .ZN(n8775) );
  INV_X1 U11101 ( .A(n8771), .ZN(n8773) );
  NAND2_X1 U11102 ( .A1(n8773), .A2(n7271), .ZN(n8774) );
  NAND2_X1 U11103 ( .A1(n8562), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8784) );
  INV_X1 U11104 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8776) );
  OAI21_X1 U11105 ( .B1(n8778), .B2(n8777), .A(n8776), .ZN(n8779) );
  NAND2_X1 U11106 ( .A1(n8779), .A2(n8840), .ZN(n13640) );
  OR2_X1 U11107 ( .A1(n9051), .A2(n13640), .ZN(n8783) );
  INV_X1 U11108 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8780) );
  OR2_X1 U11109 ( .A1(n9023), .A2(n8780), .ZN(n8782) );
  INV_X1 U11110 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n13641) );
  OR2_X1 U11111 ( .A1(n9046), .A2(n13641), .ZN(n8781) );
  NAND4_X1 U11112 ( .A1(n8784), .A2(n8783), .A3(n8782), .A4(n8781), .ZN(n13347) );
  XNOR2_X1 U11113 ( .A(n8786), .B(n8785), .ZN(n11214) );
  NAND2_X1 U11114 ( .A1(n11214), .A2(n9061), .ZN(n8790) );
  NAND2_X1 U11115 ( .A1(n8787), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8788) );
  XNOR2_X1 U11116 ( .A(n8788), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U11117 ( .A1(n9062), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8909), 
        .B2(n11860), .ZN(n8789) );
  MUX2_X1 U11118 ( .A(n13347), .B(n13644), .S(n8731), .Z(n8792) );
  MUX2_X1 U11119 ( .A(n13347), .B(n13644), .S(n9065), .Z(n8791) );
  XNOR2_X1 U11120 ( .A(n8793), .B(SI_17_), .ZN(n8794) );
  XNOR2_X1 U11121 ( .A(n8795), .B(n8794), .ZN(n11806) );
  NAND2_X1 U11122 ( .A1(n11806), .A2(n9061), .ZN(n8800) );
  INV_X1 U11123 ( .A(n8796), .ZN(n8797) );
  NAND2_X1 U11124 ( .A1(n8797), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8798) );
  XNOR2_X1 U11125 ( .A(n8798), .B(P2_IR_REG_17__SCAN_IN), .ZN(n14907) );
  AOI22_X1 U11126 ( .A1(n9062), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8909), 
        .B2(n14907), .ZN(n8799) );
  NAND2_X1 U11127 ( .A1(n8562), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8806) );
  INV_X1 U11128 ( .A(n8801), .ZN(n8878) );
  NAND2_X1 U11129 ( .A1(n8808), .A2(n15265), .ZN(n8802) );
  NAND2_X1 U11130 ( .A1(n8878), .A2(n8802), .ZN(n13597) );
  OR2_X1 U11131 ( .A1(n13597), .A2(n9051), .ZN(n8805) );
  INV_X1 U11132 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n13787) );
  OR2_X1 U11133 ( .A1(n9023), .A2(n13787), .ZN(n8804) );
  INV_X1 U11134 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13598) );
  OR2_X1 U11135 ( .A1(n9046), .A2(n13598), .ZN(n8803) );
  OR2_X1 U11136 ( .A1(n13608), .A2(n13632), .ZN(n9106) );
  NAND2_X1 U11137 ( .A1(n13608), .A2(n13632), .ZN(n11950) );
  INV_X1 U11138 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11864) );
  INV_X1 U11139 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8807) );
  OAI21_X1 U11140 ( .B1(n8842), .B2(n11864), .A(n8807), .ZN(n8809) );
  NAND2_X1 U11141 ( .A1(n8809), .A2(n8808), .ZN(n13616) );
  OR2_X1 U11142 ( .A1(n9051), .A2(n13616), .ZN(n8815) );
  INV_X1 U11143 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8810) );
  OR2_X1 U11144 ( .A1(n9052), .A2(n8810), .ZN(n8814) );
  INV_X1 U11145 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8811) );
  OR2_X1 U11146 ( .A1(n9023), .A2(n8811), .ZN(n8813) );
  INV_X1 U11147 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n13617) );
  OR2_X1 U11148 ( .A1(n9046), .A2(n13617), .ZN(n8812) );
  NAND4_X1 U11149 ( .A1(n8815), .A2(n8814), .A3(n8813), .A4(n8812), .ZN(n13345) );
  INV_X1 U11150 ( .A(n13345), .ZN(n13269) );
  NOR2_X1 U11151 ( .A1(n9065), .A2(n13269), .ZN(n8823) );
  XNOR2_X1 U11152 ( .A(n8817), .B(n8816), .ZN(n11802) );
  NAND2_X1 U11153 ( .A1(n11802), .A2(n9061), .ZN(n8821) );
  NAND2_X1 U11154 ( .A1(n8818), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8832) );
  NAND2_X1 U11155 ( .A1(n8832), .A2(n8831), .ZN(n8834) );
  NAND2_X1 U11156 ( .A1(n8834), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8819) );
  XNOR2_X1 U11157 ( .A(n8819), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14894) );
  AOI22_X1 U11158 ( .A1(n9062), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8909), 
        .B2(n14894), .ZN(n8820) );
  OAI21_X1 U11159 ( .B1(n8731), .B2(n13345), .A(n13744), .ZN(n8822) );
  OAI21_X1 U11160 ( .B1(n8823), .B2(n13744), .A(n8822), .ZN(n8824) );
  NAND3_X1 U11161 ( .A1(n9106), .A2(n11950), .A3(n8824), .ZN(n8860) );
  INV_X1 U11162 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15131) );
  OR2_X1 U11163 ( .A1(n9052), .A2(n15131), .ZN(n8828) );
  XNOR2_X1 U11164 ( .A(n8842), .B(n11864), .ZN(n11901) );
  OR2_X1 U11165 ( .A1(n9051), .A2(n11901), .ZN(n8827) );
  INV_X1 U11166 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n13792) );
  OR2_X1 U11167 ( .A1(n9023), .A2(n13792), .ZN(n8826) );
  INV_X1 U11168 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n11795) );
  OR2_X1 U11169 ( .A1(n9046), .A2(n11795), .ZN(n8825) );
  NAND4_X1 U11170 ( .A1(n8828), .A2(n8827), .A3(n8826), .A4(n8825), .ZN(n13629) );
  XNOR2_X1 U11171 ( .A(n8830), .B(n8829), .ZN(n11628) );
  NAND2_X1 U11172 ( .A1(n11628), .A2(n9061), .ZN(n8836) );
  OR2_X1 U11173 ( .A1(n8832), .A2(n8831), .ZN(n8833) );
  AND2_X1 U11174 ( .A1(n8834), .A2(n8833), .ZN(n13364) );
  AOI22_X1 U11175 ( .A1(n9062), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8909), 
        .B2(n13364), .ZN(n8835) );
  MUX2_X1 U11176 ( .A(n13629), .B(n11976), .S(n8731), .Z(n8861) );
  OR2_X1 U11177 ( .A1(n9065), .A2(n13629), .ZN(n8837) );
  OAI21_X1 U11178 ( .B1(n11976), .B2(n8754), .A(n8837), .ZN(n8862) );
  NOR2_X1 U11179 ( .A1(n8861), .A2(n8862), .ZN(n8838) );
  NOR2_X1 U11180 ( .A1(n8860), .A2(n8838), .ZN(n8855) );
  INV_X1 U11181 ( .A(n9023), .ZN(n9045) );
  NAND2_X1 U11182 ( .A1(n9045), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8846) );
  INV_X1 U11183 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n11857) );
  OR2_X1 U11184 ( .A1(n9052), .A2(n11857), .ZN(n8845) );
  NAND2_X1 U11185 ( .A1(n8840), .A2(n14875), .ZN(n8841) );
  NAND2_X1 U11186 ( .A1(n8842), .A2(n8841), .ZN(n11693) );
  OR2_X1 U11187 ( .A1(n9051), .A2(n11693), .ZN(n8844) );
  INV_X1 U11188 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11660) );
  OR2_X1 U11189 ( .A1(n9046), .A2(n11660), .ZN(n8843) );
  XNOR2_X1 U11190 ( .A(n8848), .B(n8847), .ZN(n11479) );
  NAND2_X1 U11191 ( .A1(n11479), .A2(n9061), .ZN(n8852) );
  INV_X1 U11192 ( .A(n8454), .ZN(n8849) );
  NAND2_X1 U11193 ( .A1(n8849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8850) );
  XNOR2_X1 U11194 ( .A(n8850), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14882) );
  AOI22_X1 U11195 ( .A1(n9062), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8909), 
        .B2(n14882), .ZN(n8851) );
  MUX2_X1 U11196 ( .A(n11787), .B(n11788), .S(n8754), .Z(n8857) );
  INV_X1 U11197 ( .A(n11787), .ZN(n13346) );
  MUX2_X1 U11198 ( .A(n13346), .B(n11697), .S(n9065), .Z(n8856) );
  NAND2_X1 U11199 ( .A1(n8857), .A2(n8856), .ZN(n8853) );
  INV_X1 U11200 ( .A(n8855), .ZN(n8870) );
  INV_X1 U11201 ( .A(n8856), .ZN(n8859) );
  INV_X1 U11202 ( .A(n8857), .ZN(n8858) );
  NAND2_X1 U11203 ( .A1(n8859), .A2(n8858), .ZN(n8869) );
  MUX2_X1 U11204 ( .A(n11950), .B(n9106), .S(n9065), .Z(n8868) );
  INV_X1 U11205 ( .A(n8860), .ZN(n8866) );
  INV_X1 U11206 ( .A(n8861), .ZN(n8864) );
  INV_X1 U11207 ( .A(n8862), .ZN(n8863) );
  XNOR2_X1 U11208 ( .A(n13744), .B(n13345), .ZN(n13626) );
  OAI21_X1 U11209 ( .B1(n8864), .B2(n8863), .A(n13626), .ZN(n8865) );
  NAND2_X1 U11210 ( .A1(n8866), .A2(n8865), .ZN(n8867) );
  OAI211_X1 U11211 ( .C1(n8870), .C2(n8869), .A(n8868), .B(n8867), .ZN(n8871)
         );
  INV_X1 U11212 ( .A(n8871), .ZN(n8872) );
  NAND2_X1 U11213 ( .A1(n8873), .A2(n8872), .ZN(n8896) );
  NAND2_X1 U11214 ( .A1(n8562), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U11215 ( .A1(n9045), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8874) );
  AND2_X1 U11216 ( .A1(n8875), .A2(n8874), .ZN(n8882) );
  INV_X1 U11217 ( .A(n8876), .ZN(n8900) );
  INV_X1 U11218 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8877) );
  NAND2_X1 U11219 ( .A1(n8878), .A2(n8877), .ZN(n8879) );
  NAND2_X1 U11220 ( .A1(n8900), .A2(n8879), .ZN(n13586) );
  OR2_X1 U11221 ( .A1(n13586), .A2(n9051), .ZN(n8881) );
  NAND2_X1 U11222 ( .A1(n8530), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U11223 ( .A1(n8883), .A2(n9971), .ZN(n8884) );
  NAND2_X1 U11224 ( .A1(n8886), .A2(n8885), .ZN(n8887) );
  NAND2_X1 U11225 ( .A1(n8888), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8889) );
  MUX2_X1 U11226 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8889), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n8891) );
  AND2_X1 U11227 ( .A1(n8891), .A2(n8890), .ZN(n13385) );
  AOI22_X1 U11228 ( .A1(n13385), .A2(n8909), .B1(n9062), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n8892) );
  MUX2_X1 U11229 ( .A(n13263), .B(n13590), .S(n9065), .Z(n8895) );
  MUX2_X1 U11230 ( .A(n13344), .B(n13733), .S(n8731), .Z(n8894) );
  OAI21_X1 U11231 ( .B1(n8896), .B2(n8895), .A(n8894), .ZN(n8898) );
  NAND2_X1 U11232 ( .A1(n8896), .A2(n8895), .ZN(n8897) );
  INV_X1 U11233 ( .A(n8915), .ZN(n8902) );
  INV_X1 U11234 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U11235 ( .A1(n8900), .A2(n8899), .ZN(n8901) );
  NAND2_X1 U11236 ( .A1(n8902), .A2(n8901), .ZN(n13567) );
  AOI22_X1 U11237 ( .A1(n9045), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n8562), .B2(
        P2_REG1_REG_19__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U11238 ( .A1(n8530), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8903) );
  OAI211_X1 U11239 ( .C1(n13567), .C2(n9051), .A(n8904), .B(n8903), .ZN(n13343) );
  NAND2_X1 U11240 ( .A1(n8906), .A2(n8905), .ZN(n8908) );
  NAND2_X1 U11241 ( .A1(n12039), .A2(n9061), .ZN(n8911) );
  AOI22_X1 U11242 ( .A1(n9710), .A2(n8909), .B1(n9062), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n8910) );
  INV_X1 U11243 ( .A(n8913), .ZN(n8914) );
  OR2_X1 U11244 ( .A1(n8915), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U11245 ( .A1(n8931), .A2(n8916), .ZN(n13551) );
  AOI22_X1 U11246 ( .A1(n9045), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n8562), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U11247 ( .A1(n8530), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8917) );
  OAI211_X1 U11248 ( .C1(n13551), .C2(n9051), .A(n8918), .B(n8917), .ZN(n13342) );
  INV_X1 U11249 ( .A(SI_20_), .ZN(n10519) );
  OR2_X1 U11250 ( .A1(n8919), .A2(n10519), .ZN(n8941) );
  NAND2_X1 U11251 ( .A1(n8919), .A2(n10519), .ZN(n8920) );
  NAND2_X1 U11252 ( .A1(n8941), .A2(n8920), .ZN(n8944) );
  NAND2_X1 U11253 ( .A1(n12065), .A2(n9061), .ZN(n8922) );
  NAND2_X1 U11254 ( .A1(n9062), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8921) );
  MUX2_X1 U11255 ( .A(n13342), .B(n13724), .S(n9065), .Z(n8926) );
  NAND2_X1 U11256 ( .A1(n8925), .A2(n8926), .ZN(n8924) );
  MUX2_X1 U11257 ( .A(n13342), .B(n13724), .S(n8731), .Z(n8923) );
  NAND2_X1 U11258 ( .A1(n8924), .A2(n8923), .ZN(n8930) );
  INV_X1 U11259 ( .A(n8925), .ZN(n8928) );
  INV_X1 U11260 ( .A(n8926), .ZN(n8927) );
  NAND2_X1 U11261 ( .A1(n8928), .A2(n8927), .ZN(n8929) );
  NAND2_X1 U11262 ( .A1(n8931), .A2(n13237), .ZN(n8933) );
  INV_X1 U11263 ( .A(n8952), .ZN(n8932) );
  NAND2_X1 U11264 ( .A1(n8933), .A2(n8932), .ZN(n13532) );
  OR2_X1 U11265 ( .A1(n13532), .A2(n9051), .ZN(n8938) );
  INV_X1 U11266 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13780) );
  NAND2_X1 U11267 ( .A1(n8530), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8935) );
  NAND2_X1 U11268 ( .A1(n8562), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8934) );
  OAI211_X1 U11269 ( .C1(n9023), .C2(n13780), .A(n8935), .B(n8934), .ZN(n8936)
         );
  INV_X1 U11270 ( .A(n8936), .ZN(n8937) );
  NAND2_X1 U11271 ( .A1(n8938), .A2(n8937), .ZN(n13341) );
  INV_X1 U11272 ( .A(n8939), .ZN(n8943) );
  AND2_X1 U11273 ( .A1(n8941), .A2(n8940), .ZN(n8942) );
  OAI21_X1 U11274 ( .B1(n8944), .B2(n8943), .A(n8942), .ZN(n8946) );
  NAND2_X1 U11275 ( .A1(n8946), .A2(n8945), .ZN(n12081) );
  NAND2_X1 U11276 ( .A1(n9062), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8947) );
  MUX2_X1 U11277 ( .A(n13341), .B(n13539), .S(n8754), .Z(n8950) );
  MUX2_X1 U11278 ( .A(n13341), .B(n13539), .S(n9065), .Z(n8949) );
  INV_X1 U11279 ( .A(n8950), .ZN(n8951) );
  INV_X1 U11280 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n15248) );
  OR2_X1 U11281 ( .A1(n9052), .A2(n15248), .ZN(n8956) );
  XNOR2_X1 U11282 ( .A(P2_REG3_REG_22__SCAN_IN), .B(n8952), .ZN(n13523) );
  OR2_X1 U11283 ( .A1(n9051), .A2(n13523), .ZN(n8955) );
  INV_X1 U11284 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n15260) );
  OR2_X1 U11285 ( .A1(n9023), .A2(n15260), .ZN(n8954) );
  INV_X1 U11286 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n13524) );
  OR2_X1 U11287 ( .A1(n9046), .A2(n13524), .ZN(n8953) );
  NAND4_X1 U11288 ( .A1(n8956), .A2(n8955), .A3(n8954), .A4(n8953), .ZN(n13340) );
  NAND2_X1 U11289 ( .A1(n12102), .A2(n8957), .ZN(n8958) );
  NAND2_X1 U11290 ( .A1(n8959), .A2(n8958), .ZN(n11347) );
  NAND2_X1 U11291 ( .A1(n9062), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8960) );
  MUX2_X1 U11292 ( .A(n13340), .B(n13526), .S(n9065), .Z(n8965) );
  NAND2_X1 U11293 ( .A1(n8964), .A2(n8965), .ZN(n8963) );
  MUX2_X1 U11294 ( .A(n13340), .B(n13526), .S(n8754), .Z(n8962) );
  NAND2_X1 U11295 ( .A1(n8963), .A2(n8962), .ZN(n8969) );
  INV_X1 U11296 ( .A(n8964), .ZN(n8967) );
  INV_X1 U11297 ( .A(n8965), .ZN(n8966) );
  NAND2_X1 U11298 ( .A1(n8967), .A2(n8966), .ZN(n8968) );
  NAND2_X1 U11299 ( .A1(n8969), .A2(n8968), .ZN(n8986) );
  NAND2_X1 U11300 ( .A1(n8562), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8977) );
  INV_X1 U11301 ( .A(n8970), .ZN(n8972) );
  INV_X1 U11302 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U11303 ( .A1(n8972), .A2(n8971), .ZN(n8973) );
  NAND2_X1 U11304 ( .A1(n8992), .A2(n8973), .ZN(n13501) );
  OR2_X1 U11305 ( .A1(n9051), .A2(n13501), .ZN(n8976) );
  INV_X1 U11306 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n13776) );
  OR2_X1 U11307 ( .A1(n9023), .A2(n13776), .ZN(n8975) );
  INV_X1 U11308 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13508) );
  OR2_X1 U11309 ( .A1(n9046), .A2(n13508), .ZN(n8974) );
  NAND4_X1 U11310 ( .A1(n8977), .A2(n8976), .A3(n8975), .A4(n8974), .ZN(n13339) );
  OR2_X1 U11311 ( .A1(n8979), .A2(n8978), .ZN(n8980) );
  NAND2_X1 U11312 ( .A1(n8981), .A2(n8980), .ZN(n12122) );
  OR2_X1 U11313 ( .A1(n12122), .A2(n9003), .ZN(n8983) );
  NAND2_X1 U11314 ( .A1(n9062), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8982) );
  MUX2_X1 U11315 ( .A(n13339), .B(n13507), .S(n8754), .Z(n8987) );
  NAND2_X1 U11316 ( .A1(n8986), .A2(n8987), .ZN(n8985) );
  MUX2_X1 U11317 ( .A(n13339), .B(n13507), .S(n9065), .Z(n8984) );
  NAND2_X1 U11318 ( .A1(n8985), .A2(n8984), .ZN(n8991) );
  INV_X1 U11319 ( .A(n8986), .ZN(n8989) );
  INV_X1 U11320 ( .A(n8987), .ZN(n8988) );
  NAND2_X1 U11321 ( .A1(n8989), .A2(n8988), .ZN(n8990) );
  NAND2_X1 U11322 ( .A1(n8562), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8998) );
  INV_X1 U11323 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n15141) );
  NAND2_X1 U11324 ( .A1(n8992), .A2(n15141), .ZN(n8993) );
  NAND2_X1 U11325 ( .A1(n9020), .A2(n8993), .ZN(n13487) );
  OR2_X1 U11326 ( .A1(n9051), .A2(n13487), .ZN(n8997) );
  INV_X1 U11327 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8994) );
  OR2_X1 U11328 ( .A1(n9023), .A2(n8994), .ZN(n8996) );
  INV_X1 U11329 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13491) );
  OR2_X1 U11330 ( .A1(n9046), .A2(n13491), .ZN(n8995) );
  NAND4_X1 U11331 ( .A1(n8998), .A2(n8997), .A3(n8996), .A4(n8995), .ZN(n13468) );
  OR2_X1 U11332 ( .A1(n9000), .A2(n8999), .ZN(n9001) );
  NAND2_X1 U11333 ( .A1(n9002), .A2(n9001), .ZN(n12142) );
  NAND2_X1 U11334 ( .A1(n9062), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9004) );
  MUX2_X1 U11335 ( .A(n13468), .B(n13700), .S(n8648), .Z(n9009) );
  NAND2_X1 U11336 ( .A1(n9008), .A2(n9009), .ZN(n9007) );
  MUX2_X1 U11337 ( .A(n13468), .B(n13700), .S(n8731), .Z(n9006) );
  NAND2_X1 U11338 ( .A1(n9007), .A2(n9006), .ZN(n9013) );
  INV_X1 U11339 ( .A(n9008), .ZN(n9011) );
  INV_X1 U11340 ( .A(n9009), .ZN(n9010) );
  NAND2_X1 U11341 ( .A1(n9011), .A2(n9010), .ZN(n9012) );
  NAND2_X1 U11342 ( .A1(n9013), .A2(n9012), .ZN(n9018) );
  INV_X1 U11343 ( .A(n9018), .ZN(n9016) );
  INV_X1 U11344 ( .A(n13279), .ZN(n13458) );
  MUX2_X1 U11345 ( .A(n13458), .B(n13475), .S(n9065), .Z(n9014) );
  OAI21_X1 U11346 ( .B1(n9016), .B2(n9015), .A(n9014), .ZN(n9017) );
  OAI21_X1 U11347 ( .B1(n9019), .B2(n9018), .A(n9017), .ZN(n9036) );
  NAND2_X1 U11348 ( .A1(n8562), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n9028) );
  INV_X1 U11349 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n13324) );
  OAI21_X1 U11350 ( .B1(n9020), .B2(n13248), .A(n13324), .ZN(n9021) );
  NAND2_X1 U11351 ( .A1(n9021), .A2(n9048), .ZN(n13451) );
  OR2_X1 U11352 ( .A1(n9051), .A2(n13451), .ZN(n9027) );
  INV_X1 U11353 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9022) );
  OR2_X1 U11354 ( .A1(n9023), .A2(n9022), .ZN(n9026) );
  INV_X1 U11355 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9024) );
  OR2_X1 U11356 ( .A1(n9046), .A2(n9024), .ZN(n9025) );
  NAND4_X1 U11357 ( .A1(n9028), .A2(n9027), .A3(n9026), .A4(n9025), .ZN(n13467) );
  XNOR2_X1 U11358 ( .A(n9029), .B(SI_26_), .ZN(n9030) );
  NAND2_X1 U11359 ( .A1(n12183), .A2(n9061), .ZN(n9033) );
  NAND2_X1 U11360 ( .A1(n9062), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9032) );
  MUX2_X1 U11361 ( .A(n13467), .B(n13688), .S(n8648), .Z(n9037) );
  NAND2_X1 U11362 ( .A1(n9036), .A2(n9037), .ZN(n9035) );
  MUX2_X1 U11363 ( .A(n13688), .B(n13467), .S(n9065), .Z(n9034) );
  INV_X1 U11364 ( .A(n9036), .ZN(n9039) );
  INV_X1 U11365 ( .A(n9037), .ZN(n9038) );
  NAND2_X1 U11366 ( .A1(n9041), .A2(n9040), .ZN(n9042) );
  AND2_X1 U11367 ( .A1(n9043), .A2(n9042), .ZN(n9044) );
  NAND2_X1 U11368 ( .A1(n9122), .A2(n9044), .ZN(n9071) );
  NAND2_X1 U11369 ( .A1(n9045), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9056) );
  INV_X1 U11370 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13443) );
  OR2_X1 U11371 ( .A1(n9046), .A2(n13443), .ZN(n9055) );
  INV_X1 U11372 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U11373 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  NAND2_X1 U11374 ( .A1(n9050), .A2(n9049), .ZN(n13442) );
  OR2_X1 U11375 ( .A1(n9051), .A2(n13442), .ZN(n9054) );
  INV_X1 U11376 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13685) );
  OR2_X1 U11377 ( .A1(n9052), .A2(n13685), .ZN(n9053) );
  INV_X1 U11378 ( .A(n13325), .ZN(n13459) );
  INV_X1 U11379 ( .A(n9057), .ZN(n9058) );
  XNOR2_X1 U11380 ( .A(n9058), .B(SI_27_), .ZN(n9059) );
  NAND2_X1 U11381 ( .A1(n13815), .A2(n9061), .ZN(n9064) );
  NAND2_X1 U11382 ( .A1(n9062), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9063) );
  MUX2_X1 U11383 ( .A(n13459), .B(n6764), .S(n8648), .Z(n9072) );
  MUX2_X1 U11384 ( .A(n13769), .B(n13325), .S(n9065), .Z(n9073) );
  INV_X1 U11385 ( .A(n9071), .ZN(n9076) );
  INV_X1 U11386 ( .A(n9072), .ZN(n9075) );
  INV_X1 U11387 ( .A(n9073), .ZN(n9074) );
  NAND3_X1 U11388 ( .A1(n9076), .A2(n9075), .A3(n9074), .ZN(n9077) );
  NAND2_X1 U11389 ( .A1(n9079), .A2(n9078), .ZN(n9080) );
  NAND2_X1 U11390 ( .A1(n9081), .A2(n7426), .ZN(n9128) );
  OAI21_X1 U11391 ( .B1(n9710), .B2(n11111), .A(n9751), .ZN(n9082) );
  AOI21_X1 U11392 ( .B1(n9708), .B2(n11348), .A(n9082), .ZN(n9083) );
  INV_X1 U11393 ( .A(n9083), .ZN(n9089) );
  INV_X1 U11394 ( .A(n6485), .ZN(n9127) );
  MUX2_X1 U11395 ( .A(n9101), .B(n9124), .S(n9127), .Z(n9084) );
  NAND2_X1 U11396 ( .A1(n9084), .A2(n9710), .ZN(n9085) );
  NAND2_X1 U11397 ( .A1(n9128), .A2(n9085), .ZN(n9088) );
  NAND2_X1 U11398 ( .A1(n9090), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9086) );
  XNOR2_X1 U11399 ( .A(n9086), .B(P2_IR_REG_23__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U11400 ( .A1(n9746), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11436) );
  INV_X1 U11401 ( .A(n11436), .ZN(n9087) );
  OAI211_X1 U11402 ( .C1(n9128), .C2(n9089), .A(n9088), .B(n9087), .ZN(n9131)
         );
  NAND2_X1 U11403 ( .A1(n8454), .A2(n9093), .ZN(n9094) );
  NAND2_X1 U11404 ( .A1(n9094), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9095) );
  MUX2_X1 U11405 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9095), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9096) );
  AND2_X1 U11406 ( .A1(n9092), .A2(n9096), .ZN(n9739) );
  NAND2_X1 U11407 ( .A1(n11537), .A2(n9739), .ZN(n9745) );
  NAND2_X1 U11408 ( .A1(n9092), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U11409 ( .A1(n9101), .A2(n9124), .ZN(n9789) );
  OAI21_X1 U11410 ( .B1(n9789), .B2(n9746), .A(n9098), .ZN(n9099) );
  AND2_X1 U11411 ( .A1(n9469), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14821) );
  INV_X1 U11412 ( .A(n9724), .ZN(n9723) );
  INV_X1 U11413 ( .A(n13816), .ZN(n9455) );
  INV_X1 U11414 ( .A(n9751), .ZN(n9808) );
  NAND4_X1 U11415 ( .A1(n14821), .A2(n9723), .A3(n9455), .A4(n9808), .ZN(n9100) );
  OAI211_X1 U11416 ( .C1(n9101), .C2(n11436), .A(n9100), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9130) );
  NAND2_X1 U11417 ( .A1(n13680), .A2(n13436), .ZN(n9102) );
  NAND2_X1 U11418 ( .A1(n13688), .A2(n13437), .ZN(n11967) );
  OR2_X1 U11419 ( .A1(n13688), .A2(n13437), .ZN(n9103) );
  NAND2_X1 U11420 ( .A1(n11967), .A2(n9103), .ZN(n11966) );
  NAND2_X1 U11421 ( .A1(n13475), .A2(n13279), .ZN(n11965) );
  OR2_X1 U11422 ( .A1(n13475), .A2(n13279), .ZN(n9104) );
  INV_X1 U11423 ( .A(n13468), .ZN(n13249) );
  NAND2_X1 U11424 ( .A1(n13700), .A2(n13249), .ZN(n11964) );
  OR2_X1 U11425 ( .A1(n13700), .A2(n13249), .ZN(n9105) );
  NAND2_X1 U11426 ( .A1(n11964), .A2(n9105), .ZN(n13495) );
  INV_X1 U11427 ( .A(n13342), .ZN(n13300) );
  XNOR2_X1 U11428 ( .A(n13724), .B(n13300), .ZN(n11953) );
  INV_X1 U11429 ( .A(n13340), .ZN(n11959) );
  XNOR2_X1 U11430 ( .A(n13526), .B(n11959), .ZN(n11958) );
  NAND2_X1 U11431 ( .A1(n11981), .A2(n11980), .ZN(n13562) );
  NAND2_X1 U11432 ( .A1(n9106), .A2(n11950), .ZN(n13600) );
  INV_X1 U11433 ( .A(n13626), .ZN(n11978) );
  XNOR2_X1 U11434 ( .A(n11976), .B(n13258), .ZN(n11947) );
  XNOR2_X1 U11435 ( .A(n11697), .B(n13346), .ZN(n11789) );
  NAND2_X1 U11436 ( .A1(n11189), .A2(n13350), .ZN(n11155) );
  OR2_X1 U11437 ( .A1(n11189), .A2(n13350), .ZN(n9107) );
  XNOR2_X1 U11438 ( .A(n11310), .B(n14802), .ZN(n11171) );
  XNOR2_X1 U11439 ( .A(n11100), .B(n11202), .ZN(n11098) );
  XNOR2_X2 U11440 ( .A(n10466), .B(n13358), .ZN(n9719) );
  AND2_X1 U11441 ( .A1(n9832), .A2(n9821), .ZN(n14928) );
  NAND4_X1 U11442 ( .A1(n9892), .A2(n14928), .A3(n9127), .A4(n6618), .ZN(n9111) );
  INV_X1 U11443 ( .A(n13354), .ZN(n10790) );
  NAND2_X1 U11444 ( .A1(n14938), .A2(n10790), .ZN(n10734) );
  OR2_X1 U11445 ( .A1(n14938), .A2(n10790), .ZN(n9110) );
  NOR4_X1 U11446 ( .A1(n9891), .A2(n10358), .A3(n9111), .A4(n10726), .ZN(n9112) );
  XNOR2_X1 U11447 ( .A(n10954), .B(n13352), .ZN(n10738) );
  XNOR2_X1 U11448 ( .A(n10804), .B(n13353), .ZN(n10730) );
  XNOR2_X1 U11449 ( .A(n13355), .B(n14932), .ZN(n10364) );
  NAND4_X1 U11450 ( .A1(n9112), .A2(n10738), .A3(n10730), .A4(n10364), .ZN(
        n9113) );
  NOR4_X1 U11451 ( .A1(n11157), .A2(n11171), .A3(n11098), .A4(n9113), .ZN(
        n9114) );
  XNOR2_X1 U11452 ( .A(n13644), .B(n13347), .ZN(n11651) );
  XNOR2_X1 U11453 ( .A(n14813), .B(n13348), .ZN(n11174) );
  NAND4_X1 U11454 ( .A1(n11789), .A2(n9114), .A3(n11651), .A4(n11174), .ZN(
        n9115) );
  NOR4_X1 U11455 ( .A1(n13600), .A2(n11978), .A3(n11947), .A4(n9115), .ZN(
        n9116) );
  XNOR2_X1 U11456 ( .A(n13539), .B(n13341), .ZN(n13535) );
  XNOR2_X1 U11457 ( .A(n13733), .B(n13344), .ZN(n13579) );
  NAND4_X1 U11458 ( .A1(n13562), .A2(n9116), .A3(n13535), .A4(n13579), .ZN(
        n9117) );
  NOR4_X1 U11459 ( .A1(n13495), .A2(n11953), .A3(n11958), .A4(n9117), .ZN(
        n9118) );
  XNOR2_X1 U11460 ( .A(n13507), .B(n13339), .ZN(n13509) );
  NAND3_X1 U11461 ( .A1(n13470), .A2(n9118), .A3(n13509), .ZN(n9119) );
  NOR4_X1 U11462 ( .A1(n13415), .A2(n13434), .A3(n11966), .A4(n9119), .ZN(
        n9121) );
  XNOR2_X1 U11463 ( .A(n13411), .B(n13337), .ZN(n9120) );
  XNOR2_X1 U11464 ( .A(n13672), .B(n13426), .ZN(n11990) );
  NAND4_X1 U11465 ( .A1(n9122), .A2(n9121), .A3(n9120), .A4(n11990), .ZN(n9123) );
  XOR2_X1 U11466 ( .A(n9710), .B(n9123), .Z(n9125) );
  NOR3_X1 U11467 ( .A1(n9125), .A2(n9124), .A3(n11436), .ZN(n9126) );
  OAI21_X1 U11468 ( .B1(n9128), .B2(n9127), .A(n9126), .ZN(n9129) );
  NAND3_X1 U11469 ( .A1(n9131), .A2(n9130), .A3(n9129), .ZN(P2_U3328) );
  INV_X1 U11470 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9133) );
  INV_X1 U11471 ( .A(n9134), .ZN(n9135) );
  NAND2_X1 U11472 ( .A1(n9136), .A2(n9135), .ZN(P3_U3488) );
  INV_X1 U11473 ( .A(n13131), .ZN(n9353) );
  INV_X2 U11474 ( .A(n13360), .ZN(P2_U3947) );
  NAND2_X2 U11475 ( .A1(n9214), .A2(n9215), .ZN(n9259) );
  INV_X2 U11476 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9266) );
  INV_X2 U11477 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10266) );
  INV_X2 U11478 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10265) );
  INV_X2 U11479 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9310) );
  INV_X2 U11480 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9305) );
  NAND4_X1 U11481 ( .A1(n10266), .A2(n10265), .A3(n9310), .A4(n9305), .ZN(
        n9143) );
  NOR2_X2 U11482 ( .A1(n9494), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n9183) );
  OAI21_X1 U11483 ( .B1(n6812), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9147) );
  INV_X1 U11484 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9146) );
  XNOR2_X1 U11485 ( .A(n9147), .B(n9146), .ZN(n9206) );
  NOR2_X1 U11486 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n9150) );
  NOR2_X1 U11487 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n9149) );
  NOR2_X1 U11488 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n9148) );
  INV_X1 U11489 ( .A(n9155), .ZN(n9151) );
  NOR2_X1 U11490 ( .A1(n10946), .A2(n9151), .ZN(n9159) );
  INV_X1 U11491 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9152) );
  NAND2_X1 U11492 ( .A1(n9159), .A2(n9152), .ZN(n9162) );
  NAND2_X1 U11493 ( .A1(n9162), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9153) );
  MUX2_X1 U11494 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9153), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n9158) );
  NOR3_X1 U11495 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .A3(P1_IR_REG_25__SCAN_IN), .ZN(n9154) );
  INV_X1 U11496 ( .A(n9159), .ZN(n9160) );
  NAND2_X1 U11497 ( .A1(n9160), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9161) );
  NAND2_X1 U11498 ( .A1(n9164), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9165) );
  XNOR2_X1 U11499 ( .A(n9165), .B(n9167), .ZN(n11906) );
  NOR2_X1 U11500 ( .A1(n11596), .A2(n11906), .ZN(n9166) );
  INV_X1 U11501 ( .A(n9770), .ZN(n9197) );
  AND2_X2 U11502 ( .A1(n9295), .A2(n9197), .ZN(P1_U4016) );
  AND2_X1 U11503 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9418) );
  XNOR2_X2 U11504 ( .A(n9169), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U11505 ( .A1(n9170), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9171) );
  MUX2_X1 U11506 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9171), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n9173) );
  INV_X1 U11507 ( .A(n9172), .ZN(n14387) );
  AND2_X4 U11508 ( .A1(n9174), .A2(n9175), .ZN(n9937) );
  NAND2_X1 U11509 ( .A1(n9937), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9179) );
  AND2_X4 U11510 ( .A1(n12001), .A2(n14394), .ZN(n12441) );
  NAND2_X1 U11511 ( .A1(n12441), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9178) );
  AND2_X2 U11512 ( .A1(n9174), .A2(n14394), .ZN(n12223) );
  NAND2_X1 U11513 ( .A1(n12223), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U11514 ( .A1(n9936), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9176) );
  NAND2_X1 U11515 ( .A1(n9180), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9181) );
  MUX2_X1 U11516 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9181), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n9182) );
  AND2_X2 U11517 ( .A1(n9182), .A2(n6812), .ZN(n12447) );
  INV_X1 U11518 ( .A(n9183), .ZN(n9184) );
  NAND2_X1 U11519 ( .A1(n9184), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9186) );
  OR2_X1 U11520 ( .A1(n7455), .A2(n12230), .ZN(n9196) );
  INV_X1 U11521 ( .A(SI_0_), .ZN(n9188) );
  OAI21_X1 U11522 ( .B1(n12101), .B2(n9188), .A(n9187), .ZN(n9189) );
  AND2_X1 U11523 ( .A1(n9190), .A2(n9189), .ZN(n14400) );
  AND2_X4 U11524 ( .A1(n12262), .A2(n9770), .ZN(n12205) );
  AOI22_X1 U11525 ( .A1(n14279), .A2(n12205), .B1(n9197), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9195) );
  AND2_X1 U11526 ( .A1(n9196), .A2(n9195), .ZN(n9611) );
  NAND2_X1 U11527 ( .A1(n9579), .A2(n12257), .ZN(n12461) );
  OR2_X1 U11528 ( .A1(n7455), .A2(n12228), .ZN(n9199) );
  AOI22_X1 U11529 ( .A1(n9767), .A2(n14279), .B1(n9197), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9198) );
  NAND2_X1 U11530 ( .A1(n9199), .A2(n9198), .ZN(n9200) );
  NOR2_X1 U11531 ( .A1(n9611), .A2(n9200), .ZN(n9610) );
  AOI21_X1 U11532 ( .B1(n9611), .B2(n9200), .A(n9610), .ZN(n9594) );
  MUX2_X1 U11533 ( .A(n9418), .B(n9594), .S(n14398), .Z(n9204) );
  INV_X1 U11534 ( .A(n11945), .ZN(n9616) );
  INV_X1 U11535 ( .A(n14398), .ZN(n9202) );
  INV_X1 U11536 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9213) );
  AOI21_X1 U11537 ( .B1(n9202), .B2(n9213), .A(n11945), .ZN(n9315) );
  OAI21_X1 U11538 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9315), .A(P1_U4016), .ZN(
        n9203) );
  AOI21_X1 U11539 ( .B1(n9204), .B2(n9616), .A(n9203), .ZN(n9640) );
  AND2_X1 U11540 ( .A1(n9295), .A2(n9770), .ZN(n10489) );
  INV_X1 U11541 ( .A(n9206), .ZN(n9205) );
  NAND2_X1 U11542 ( .A1(n9205), .A2(P1_STATE_REG_SCAN_IN), .ZN(n12517) );
  INV_X1 U11543 ( .A(n12517), .ZN(n11433) );
  OR2_X1 U11544 ( .A1(n10489), .A2(n11433), .ZN(n9228) );
  NAND2_X1 U11545 ( .A1(n12254), .A2(n12447), .ZN(n12462) );
  INV_X1 U11546 ( .A(n12462), .ZN(n9617) );
  NAND2_X1 U11547 ( .A1(n9617), .A2(n9206), .ZN(n9207) );
  INV_X1 U11548 ( .A(n9227), .ZN(n9208) );
  NOR2_X1 U11549 ( .A1(n11945), .A2(n14398), .ZN(n9209) );
  NAND2_X1 U11550 ( .A1(n9320), .A2(n9209), .ZN(n14686) );
  INV_X1 U11551 ( .A(n14686), .ZN(n14027) );
  INV_X1 U11552 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10494) );
  INV_X1 U11553 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U11554 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9210) );
  MUX2_X1 U11555 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10494), .S(n9606), .Z(n9420) );
  INV_X1 U11556 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9212) );
  NOR3_X1 U11557 ( .A1(n9420), .A2(n9213), .A3(n9212), .ZN(n9419) );
  NOR2_X1 U11558 ( .A1(n9606), .A2(n10494), .ZN(n9219) );
  INV_X1 U11559 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9217) );
  INV_X1 U11560 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14386) );
  OR2_X1 U11561 ( .A1(n9214), .A2(n14386), .ZN(n9216) );
  XNOR2_X1 U11562 ( .A(n9216), .B(n9215), .ZN(n9643) );
  MUX2_X1 U11563 ( .A(n9217), .B(P1_REG2_REG_2__SCAN_IN), .S(n9643), .Z(n9218)
         );
  OAI21_X1 U11564 ( .B1(n9419), .B2(n9219), .A(n9218), .ZN(n9407) );
  INV_X1 U11565 ( .A(n9419), .ZN(n9222) );
  INV_X1 U11566 ( .A(n9219), .ZN(n9221) );
  MUX2_X1 U11567 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9217), .S(n9643), .Z(n9220)
         );
  NAND3_X1 U11568 ( .A1(n9222), .A2(n9221), .A3(n9220), .ZN(n9223) );
  AND3_X1 U11569 ( .A1(n14027), .A2(n9407), .A3(n9223), .ZN(n9232) );
  INV_X1 U11570 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14787) );
  INV_X1 U11571 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9224) );
  MUX2_X1 U11572 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9224), .S(n9643), .Z(n9225)
         );
  NOR2_X1 U11573 ( .A1(n9226), .A2(n9225), .ZN(n9328) );
  AOI211_X1 U11574 ( .C1(n9226), .C2(n9225), .A(n9328), .B(n13980), .ZN(n9231)
         );
  NAND2_X1 U11575 ( .A1(n9320), .A2(n11945), .ZN(n14023) );
  NAND2_X1 U11576 ( .A1(n9228), .A2(n9227), .ZN(n14691) );
  INV_X1 U11577 ( .A(n14691), .ZN(n13986) );
  AOI22_X1 U11578 ( .A1(n13986), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9229) );
  OAI21_X1 U11579 ( .B1(n9643), .B2(n14023), .A(n9229), .ZN(n9230) );
  OR4_X1 U11580 ( .A1(n9640), .A2(n9232), .A3(n9231), .A4(n9230), .ZN(P1_U3245) );
  NAND2_X2 U11581 ( .A1(n12101), .A2(P3_U3151), .ZN(n13143) );
  AND2_X1 U11582 ( .A1(n6636), .A2(P3_U3151), .ZN(n10968) );
  OAI222_X1 U11583 ( .A1(P3_U3151), .A2(n10240), .B1(n13143), .B2(n9234), .C1(
        n6484), .C2(n9233), .ZN(P3_U3290) );
  OAI222_X1 U11584 ( .A1(P3_U3151), .A2(n10219), .B1(n13143), .B2(n9236), .C1(
        n6484), .C2(n9235), .ZN(P3_U3291) );
  OAI222_X1 U11585 ( .A1(n6484), .A2(n9238), .B1(n13143), .B2(n9237), .C1(
        P3_U3151), .C2(n10012), .ZN(P3_U3294) );
  OAI222_X1 U11586 ( .A1(n10216), .A2(P3_U3151), .B1(n6484), .B2(n9240), .C1(
        n9239), .C2(n13143), .ZN(P3_U3293) );
  INV_X1 U11587 ( .A(n12736), .ZN(n10251) );
  INV_X1 U11588 ( .A(SI_6_), .ZN(n9241) );
  OAI222_X1 U11589 ( .A1(P3_U3151), .A2(n10251), .B1(n6484), .B2(n9242), .C1(
        n9241), .C2(n13143), .ZN(P3_U3289) );
  OAI222_X1 U11590 ( .A1(n10281), .A2(P3_U3151), .B1(n6484), .B2(n9244), .C1(
        n9243), .C2(n13143), .ZN(P3_U3288) );
  OAI222_X1 U11591 ( .A1(n10196), .A2(P3_U3151), .B1(n6484), .B2(n9246), .C1(
        n9245), .C2(n13143), .ZN(P3_U3292) );
  INV_X1 U11592 ( .A(SI_8_), .ZN(n9248) );
  OAI222_X1 U11593 ( .A1(P3_U3151), .A2(n10407), .B1(n13143), .B2(n9248), .C1(
        n6484), .C2(n9247), .ZN(P3_U3287) );
  NAND2_X1 U11594 ( .A1(n6636), .A2(P2_U3088), .ZN(n13798) );
  NAND2_X1 U11595 ( .A1(n9249), .A2(P2_U3088), .ZN(n13803) );
  INV_X1 U11596 ( .A(n9754), .ZN(n9258) );
  OAI222_X1 U11597 ( .A1(n13798), .A2(n9250), .B1(n13803), .B2(n9258), .C1(
        P2_U3088), .C2(n9546), .ZN(P2_U3324) );
  INV_X1 U11598 ( .A(n13798), .ZN(n11536) );
  AOI22_X1 U11599 ( .A1(n11536), .A2(P1_DATAO_REG_1__SCAN_IN), .B1(n6482), 
        .B2(P2_STATE_REG_SCAN_IN), .ZN(n9251) );
  OAI21_X1 U11600 ( .B1(n9604), .B2(n13803), .A(n9251), .ZN(P2_U3326) );
  INV_X1 U11601 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9252) );
  INV_X1 U11602 ( .A(n9929), .ZN(n9262) );
  INV_X1 U11603 ( .A(n9463), .ZN(n9532) );
  OAI222_X1 U11604 ( .A1(n13798), .A2(n9252), .B1(n13803), .B2(n9262), .C1(
        P2_U3088), .C2(n9532), .ZN(P2_U3323) );
  INV_X1 U11605 ( .A(SI_9_), .ZN(n9253) );
  OAI222_X1 U11606 ( .A1(n10399), .A2(P3_U3151), .B1(n6484), .B2(n9254), .C1(
        n9253), .C2(n13143), .ZN(P3_U3286) );
  NAND2_X1 U11607 ( .A1(n9259), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9256) );
  XNOR2_X1 U11608 ( .A(n9256), .B(n9255), .ZN(n9758) );
  OAI222_X1 U11609 ( .A1(n9758), .A2(P1_U3086), .B1(n14391), .B2(n9258), .C1(
        n9755), .C2(n14396), .ZN(P1_U3352) );
  NAND2_X1 U11610 ( .A1(n9264), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9260) );
  XNOR2_X1 U11611 ( .A(n9260), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9930) );
  INV_X1 U11612 ( .A(n9930), .ZN(n9636) );
  OAI222_X1 U11613 ( .A1(n9636), .A2(P1_U3086), .B1(n14391), .B2(n9262), .C1(
        n9261), .C2(n14396), .ZN(P1_U3351) );
  INV_X1 U11614 ( .A(n11536), .ZN(n13819) );
  INV_X1 U11615 ( .A(n9461), .ZN(n14838) );
  OAI222_X1 U11616 ( .A1(n13819), .A2(n9263), .B1(n13803), .B2(n9641), .C1(
        P2_U3088), .C2(n14838), .ZN(P2_U3325) );
  NOR2_X1 U11617 ( .A1(n9267), .A2(n14386), .ZN(n9265) );
  MUX2_X1 U11618 ( .A(n14386), .B(n9265), .S(P1_IR_REG_5__SCAN_IN), .Z(n9269)
         );
  INV_X1 U11619 ( .A(n10342), .ZN(n9268) );
  INV_X1 U11620 ( .A(n10587), .ZN(n9271) );
  OAI222_X1 U11621 ( .A1(n9390), .A2(P1_U3086), .B1(n14391), .B2(n9271), .C1(
        n9270), .C2(n14396), .ZN(P1_U3350) );
  INV_X1 U11622 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9272) );
  INV_X1 U11623 ( .A(n9550), .ZN(n9471) );
  OAI222_X1 U11624 ( .A1(n13798), .A2(n9272), .B1(n13803), .B2(n9271), .C1(
        P2_U3088), .C2(n9471), .ZN(P2_U3322) );
  OAI222_X1 U11625 ( .A1(P3_U3151), .A2(n11256), .B1(n13143), .B2(n9274), .C1(
        n6484), .C2(n9273), .ZN(P3_U3285) );
  INV_X1 U11626 ( .A(n10592), .ZN(n9285) );
  INV_X1 U11627 ( .A(n9569), .ZN(n9560) );
  OAI222_X1 U11628 ( .A1(n13798), .A2(n9276), .B1(n13803), .B2(n9285), .C1(
        P2_U3088), .C2(n9560), .ZN(P2_U3321) );
  OAI222_X1 U11629 ( .A1(P3_U3151), .A2(n11257), .B1(n13143), .B2(n9278), .C1(
        n6484), .C2(n9277), .ZN(P3_U3284) );
  OAI222_X1 U11630 ( .A1(n9606), .A2(P1_U3086), .B1(n14391), .B2(n9604), .C1(
        n9605), .C2(n14396), .ZN(P1_U3354) );
  INV_X1 U11631 ( .A(n13803), .ZN(n13810) );
  INV_X1 U11632 ( .A(n13810), .ZN(n13817) );
  INV_X1 U11633 ( .A(n10604), .ZN(n9281) );
  INV_X1 U11634 ( .A(n9850), .ZN(n9577) );
  OAI222_X1 U11635 ( .A1(n13798), .A2(n9279), .B1(n13817), .B2(n9281), .C1(
        P2_U3088), .C2(n9577), .ZN(P2_U3320) );
  NAND2_X1 U11636 ( .A1(n9298), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9280) );
  XNOR2_X1 U11637 ( .A(n9280), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10605) );
  INV_X1 U11638 ( .A(n10605), .ZN(n9480) );
  OAI222_X1 U11639 ( .A1(n9480), .A2(P1_U3086), .B1(n14391), .B2(n9281), .C1(
        n6663), .C2(n14396), .ZN(P1_U3348) );
  OAI222_X1 U11640 ( .A1(n9643), .A2(P1_U3086), .B1(n14391), .B2(n9641), .C1(
        n9642), .C2(n14396), .ZN(P1_U3353) );
  NAND2_X1 U11641 ( .A1(n10342), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9282) );
  MUX2_X1 U11642 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9282), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n9283) );
  AND2_X1 U11643 ( .A1(n9283), .A2(n9298), .ZN(n10593) );
  INV_X1 U11644 ( .A(n10593), .ZN(n9440) );
  OAI222_X1 U11645 ( .A1(n9440), .A2(P1_U3086), .B1(n14391), .B2(n9285), .C1(
        n9284), .C2(n14396), .ZN(P1_U3349) );
  OAI222_X1 U11646 ( .A1(P3_U3151), .A2(n11921), .B1(n13143), .B2(n9287), .C1(
        n6484), .C2(n9286), .ZN(P3_U3283) );
  NAND2_X1 U11647 ( .A1(n11596), .A2(P1_B_REG_SCAN_IN), .ZN(n9290) );
  INV_X1 U11648 ( .A(n11596), .ZN(n9288) );
  INV_X1 U11649 ( .A(P1_B_REG_SCAN_IN), .ZN(n14037) );
  AOI21_X1 U11650 ( .B1(n9288), .B2(n14037), .A(n11906), .ZN(n9289) );
  NAND2_X1 U11651 ( .A1(n10489), .A2(n9583), .ZN(n14726) );
  INV_X1 U11652 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U11653 ( .A1(n11596), .A2(n11906), .ZN(n9518) );
  INV_X1 U11654 ( .A(n9518), .ZN(n9291) );
  AOI22_X1 U11655 ( .A1(n14726), .A2(n9292), .B1(n9295), .B2(n9291), .ZN(
        P1_U3445) );
  INV_X1 U11656 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9296) );
  INV_X1 U11657 ( .A(n11906), .ZN(n9293) );
  INV_X1 U11658 ( .A(n9584), .ZN(n9294) );
  AOI22_X1 U11659 ( .A1(n14726), .A2(n9296), .B1(n9295), .B2(n9294), .ZN(
        P1_U3446) );
  NAND2_X1 U11660 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n13360), .ZN(n9297) );
  OAI21_X1 U11661 ( .B1(n13632), .B2(n13360), .A(n9297), .ZN(P2_U3548) );
  NAND2_X1 U11662 ( .A1(n9346), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9306) );
  XNOR2_X1 U11663 ( .A(n9306), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10834) );
  INV_X1 U11664 ( .A(n10834), .ZN(n9489) );
  INV_X1 U11665 ( .A(n10833), .ZN(n9300) );
  OAI222_X1 U11666 ( .A1(n9489), .A2(P1_U3086), .B1(n14391), .B2(n9300), .C1(
        n9299), .C2(n14396), .ZN(P1_U3347) );
  INV_X1 U11667 ( .A(n10126), .ZN(n9857) );
  OAI222_X1 U11668 ( .A1(n13798), .A2(n9301), .B1(n13803), .B2(n9300), .C1(
        P2_U3088), .C2(n9857), .ZN(P2_U3319) );
  NOR2_X1 U11669 ( .A1(n13986), .A2(P1_U4016), .ZN(P1_U3085) );
  NAND2_X1 U11670 ( .A1(n9695), .A2(n13131), .ZN(n9302) );
  OAI21_X1 U11671 ( .B1(n13131), .B2(n9303), .A(n9302), .ZN(P3_U3377) );
  INV_X1 U11672 ( .A(n10839), .ZN(n9309) );
  INV_X1 U11673 ( .A(n10664), .ZN(n10134) );
  OAI222_X1 U11674 ( .A1(n13798), .A2(n9304), .B1(n13817), .B2(n9309), .C1(
        P2_U3088), .C2(n10134), .ZN(P2_U3318) );
  NAND2_X1 U11675 ( .A1(n9306), .A2(n9305), .ZN(n9307) );
  NAND2_X1 U11676 ( .A1(n9307), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9311) );
  XNOR2_X1 U11677 ( .A(n9311), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10840) );
  INV_X1 U11678 ( .A(n10840), .ZN(n9984) );
  INV_X1 U11679 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9308) );
  OAI222_X1 U11680 ( .A1(n9984), .A2(P1_U3086), .B1(n14391), .B2(n9309), .C1(
        n9308), .C2(n14396), .ZN(P1_U3346) );
  INV_X1 U11681 ( .A(n10884), .ZN(n9324) );
  NAND2_X1 U11682 ( .A1(n9311), .A2(n9310), .ZN(n9312) );
  NAND2_X1 U11683 ( .A1(n9312), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9313) );
  XNOR2_X1 U11684 ( .A(n9313), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10885) );
  INV_X1 U11685 ( .A(n14396), .ZN(n14389) );
  AOI22_X1 U11686 ( .A1(n10885), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n14389), .ZN(n9314) );
  OAI21_X1 U11687 ( .B1(n9324), .B2(n14391), .A(n9314), .ZN(P1_U3345) );
  INV_X1 U11688 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9323) );
  INV_X1 U11689 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9316) );
  NAND3_X1 U11690 ( .A1(n14680), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9316), .ZN(
        n9322) );
  INV_X1 U11691 ( .A(n9315), .ZN(n9317) );
  AOI21_X1 U11692 ( .B1(n14398), .B2(n9316), .A(n9317), .ZN(n9318) );
  MUX2_X1 U11693 ( .A(n9318), .B(n9317), .S(P1_IR_REG_0__SCAN_IN), .Z(n9319)
         );
  AOI22_X1 U11694 ( .A1(n9320), .A2(n9319), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9321) );
  OAI211_X1 U11695 ( .C1(n14691), .C2(n9323), .A(n9322), .B(n9321), .ZN(
        P1_U3243) );
  INV_X1 U11696 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9325) );
  INV_X1 U11697 ( .A(n11395), .ZN(n11406) );
  OAI222_X1 U11698 ( .A1(n13798), .A2(n9325), .B1(n13817), .B2(n9324), .C1(
        P2_U3088), .C2(n11406), .ZN(P2_U3317) );
  OAI222_X1 U11699 ( .A1(P3_U3151), .A2(n14993), .B1(n13143), .B2(n9327), .C1(
        n6484), .C2(n9326), .ZN(P3_U3282) );
  XNOR2_X1 U11700 ( .A(n9390), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9331) );
  INV_X1 U11701 ( .A(n9643), .ZN(n9332) );
  AOI21_X1 U11702 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n9332), .A(n9328), .ZN(
        n9404) );
  INV_X1 U11703 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9329) );
  MUX2_X1 U11704 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9329), .S(n9758), .Z(n9403)
         );
  INV_X1 U11705 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9330) );
  MUX2_X1 U11706 ( .A(n9330), .B(P1_REG1_REG_4__SCAN_IN), .S(n9930), .Z(n9627)
         );
  NAND2_X1 U11707 ( .A1(n6543), .A2(n9331), .ZN(n9386) );
  OAI21_X1 U11708 ( .B1(n9331), .B2(n6543), .A(n9386), .ZN(n9340) );
  NAND2_X1 U11709 ( .A1(n9332), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9406) );
  INV_X1 U11710 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9333) );
  MUX2_X1 U11711 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9333), .S(n9758), .Z(n9405)
         );
  AOI21_X1 U11712 ( .B1(n9407), .B2(n9406), .A(n9405), .ZN(n9632) );
  NOR2_X1 U11713 ( .A1(n9758), .A2(n9333), .ZN(n9631) );
  INV_X1 U11714 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9334) );
  MUX2_X1 U11715 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9334), .S(n9930), .Z(n9630)
         );
  OAI21_X1 U11716 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(n9629) );
  NAND2_X1 U11717 ( .A1(n9930), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9337) );
  INV_X1 U11718 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9335) );
  MUX2_X1 U11719 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n9335), .S(n9390), .Z(n9336)
         );
  AOI21_X1 U11720 ( .B1(n9629), .B2(n9337), .A(n9336), .ZN(n9432) );
  AND3_X1 U11721 ( .A1(n9629), .A2(n9337), .A3(n9336), .ZN(n9338) );
  NOR3_X1 U11722 ( .A1(n14686), .A2(n9432), .A3(n9338), .ZN(n9339) );
  AOI21_X1 U11723 ( .B1(n9340), .B2(n14680), .A(n9339), .ZN(n9343) );
  NAND2_X1 U11724 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10677) );
  INV_X1 U11725 ( .A(n10677), .ZN(n9341) );
  AOI21_X1 U11726 ( .B1(n13986), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9341), .ZN(
        n9342) );
  OAI211_X1 U11727 ( .C1(n9390), .C2(n14023), .A(n9343), .B(n9342), .ZN(
        P1_U3248) );
  INV_X1 U11728 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n9344) );
  NAND3_X1 U11729 ( .A1(n9310), .A2(n9305), .A3(n9344), .ZN(n9345) );
  OR2_X1 U11730 ( .A1(n9446), .A2(n14386), .ZN(n9347) );
  XNOR2_X1 U11731 ( .A(n9347), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10977) );
  INV_X1 U11732 ( .A(n10977), .ZN(n10336) );
  INV_X1 U11733 ( .A(n10976), .ZN(n9349) );
  OAI222_X1 U11734 ( .A1(n10336), .A2(P1_U3086), .B1(n14391), .B2(n9349), .C1(
        n9348), .C2(n14396), .ZN(P1_U3344) );
  INV_X1 U11735 ( .A(n14859), .ZN(n11408) );
  OAI222_X1 U11736 ( .A1(n13798), .A2(n9350), .B1(n13817), .B2(n9349), .C1(
        P2_U3088), .C2(n11408), .ZN(P2_U3316) );
  NAND2_X1 U11737 ( .A1(n13404), .A2(P2_U3947), .ZN(n9351) );
  OAI21_X1 U11738 ( .B1(P2_U3947), .B2(n9352), .A(n9351), .ZN(P2_U3562) );
  NOR2_X1 U11739 ( .A1(n8034), .A2(n9353), .ZN(n9355) );
  CLKBUF_X1 U11740 ( .A(n9355), .Z(n9385) );
  INV_X1 U11741 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n9354) );
  NOR2_X1 U11742 ( .A1(n9385), .A2(n9354), .ZN(P3_U3261) );
  INV_X1 U11743 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n9356) );
  NOR2_X1 U11744 ( .A1(n9385), .A2(n9356), .ZN(P3_U3260) );
  INV_X1 U11745 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n9357) );
  NOR2_X1 U11746 ( .A1(n9385), .A2(n9357), .ZN(P3_U3263) );
  INV_X1 U11747 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n9358) );
  NOR2_X1 U11748 ( .A1(n9355), .A2(n9358), .ZN(P3_U3262) );
  INV_X1 U11749 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n9359) );
  NOR2_X1 U11750 ( .A1(n9385), .A2(n9359), .ZN(P3_U3257) );
  INV_X1 U11751 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n9360) );
  NOR2_X1 U11752 ( .A1(n9385), .A2(n9360), .ZN(P3_U3251) );
  INV_X1 U11753 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n9361) );
  NOR2_X1 U11754 ( .A1(n9385), .A2(n9361), .ZN(P3_U3259) );
  INV_X1 U11755 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n9362) );
  NOR2_X1 U11756 ( .A1(n9355), .A2(n9362), .ZN(P3_U3258) );
  INV_X1 U11757 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n9363) );
  NOR2_X1 U11758 ( .A1(n9385), .A2(n9363), .ZN(P3_U3255) );
  INV_X1 U11759 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n9364) );
  NOR2_X1 U11760 ( .A1(n9385), .A2(n9364), .ZN(P3_U3254) );
  INV_X1 U11761 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n9365) );
  NOR2_X1 U11762 ( .A1(n9385), .A2(n9365), .ZN(P3_U3253) );
  INV_X1 U11763 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n9366) );
  NOR2_X1 U11764 ( .A1(n9385), .A2(n9366), .ZN(P3_U3252) );
  INV_X1 U11765 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n9367) );
  NOR2_X1 U11766 ( .A1(n9355), .A2(n9367), .ZN(P3_U3234) );
  INV_X1 U11767 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n9368) );
  NOR2_X1 U11768 ( .A1(n9355), .A2(n9368), .ZN(P3_U3235) );
  INV_X1 U11769 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n9369) );
  NOR2_X1 U11770 ( .A1(n9355), .A2(n9369), .ZN(P3_U3236) );
  INV_X1 U11771 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n9370) );
  NOR2_X1 U11772 ( .A1(n9355), .A2(n9370), .ZN(P3_U3237) );
  INV_X1 U11773 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n9371) );
  NOR2_X1 U11774 ( .A1(n9355), .A2(n9371), .ZN(P3_U3238) );
  INV_X1 U11775 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n9372) );
  NOR2_X1 U11776 ( .A1(n9355), .A2(n9372), .ZN(P3_U3239) );
  INV_X1 U11777 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n9373) );
  NOR2_X1 U11778 ( .A1(n9355), .A2(n9373), .ZN(P3_U3240) );
  INV_X1 U11779 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n9374) );
  NOR2_X1 U11780 ( .A1(n9355), .A2(n9374), .ZN(P3_U3241) );
  INV_X1 U11781 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n9375) );
  NOR2_X1 U11782 ( .A1(n9355), .A2(n9375), .ZN(P3_U3242) );
  INV_X1 U11783 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n9376) );
  NOR2_X1 U11784 ( .A1(n9385), .A2(n9376), .ZN(P3_U3243) );
  INV_X1 U11785 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n9377) );
  NOR2_X1 U11786 ( .A1(n9385), .A2(n9377), .ZN(P3_U3244) );
  INV_X1 U11787 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n9378) );
  NOR2_X1 U11788 ( .A1(n9385), .A2(n9378), .ZN(P3_U3245) );
  INV_X1 U11789 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n9379) );
  NOR2_X1 U11790 ( .A1(n9385), .A2(n9379), .ZN(P3_U3246) );
  INV_X1 U11791 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n9380) );
  NOR2_X1 U11792 ( .A1(n9385), .A2(n9380), .ZN(P3_U3247) );
  INV_X1 U11793 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n9381) );
  NOR2_X1 U11794 ( .A1(n9385), .A2(n9381), .ZN(P3_U3248) );
  INV_X1 U11795 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n9382) );
  NOR2_X1 U11796 ( .A1(n9385), .A2(n9382), .ZN(P3_U3249) );
  INV_X1 U11797 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n9383) );
  NOR2_X1 U11798 ( .A1(n9385), .A2(n9383), .ZN(P3_U3250) );
  INV_X1 U11799 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n9384) );
  NOR2_X1 U11800 ( .A1(n9385), .A2(n9384), .ZN(P3_U3256) );
  INV_X1 U11801 ( .A(n9390), .ZN(n10588) );
  OAI21_X1 U11802 ( .B1(n10588), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9386), .ZN(
        n9427) );
  XNOR2_X1 U11803 ( .A(n10593), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n9428) );
  NOR2_X1 U11804 ( .A1(n9427), .A2(n9428), .ZN(n9426) );
  INV_X1 U11805 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9387) );
  MUX2_X1 U11806 ( .A(n9387), .B(P1_REG1_REG_7__SCAN_IN), .S(n10605), .Z(n9388) );
  AOI211_X1 U11807 ( .C1(n9389), .C2(n9388), .A(n13980), .B(n9475), .ZN(n9401)
         );
  NOR2_X1 U11808 ( .A1(n9390), .A2(n9335), .ZN(n9431) );
  INV_X1 U11809 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9391) );
  MUX2_X1 U11810 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9391), .S(n10593), .Z(n9430) );
  OAI21_X1 U11811 ( .B1(n9432), .B2(n9431), .A(n9430), .ZN(n9429) );
  NAND2_X1 U11812 ( .A1(n10593), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9394) );
  INV_X1 U11813 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9392) );
  MUX2_X1 U11814 ( .A(n9392), .B(P1_REG2_REG_7__SCAN_IN), .S(n10605), .Z(n9393) );
  AOI21_X1 U11815 ( .B1(n9429), .B2(n9394), .A(n9393), .ZN(n9486) );
  INV_X1 U11816 ( .A(n9486), .ZN(n9396) );
  NAND3_X1 U11817 ( .A1(n9429), .A2(n9394), .A3(n9393), .ZN(n9395) );
  NAND3_X1 U11818 ( .A1(n9396), .A2(n14027), .A3(n9395), .ZN(n9399) );
  NAND2_X1 U11819 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11088) );
  INV_X1 U11820 ( .A(n11088), .ZN(n9397) );
  AOI21_X1 U11821 ( .B1(n13986), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9397), .ZN(
        n9398) );
  OAI211_X1 U11822 ( .C1(n14023), .C2(n9480), .A(n9399), .B(n9398), .ZN(n9400)
         );
  OR2_X1 U11823 ( .A1(n9401), .A2(n9400), .ZN(P1_U3250) );
  AOI211_X1 U11824 ( .C1(n9404), .C2(n9403), .A(n9402), .B(n13980), .ZN(n9410)
         );
  AND3_X1 U11825 ( .A1(n9407), .A2(n9406), .A3(n9405), .ZN(n9408) );
  NOR3_X1 U11826 ( .A1(n14686), .A2(n9632), .A3(n9408), .ZN(n9409) );
  NOR2_X1 U11827 ( .A1(n9410), .A2(n9409), .ZN(n9413) );
  NOR2_X1 U11828 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9776), .ZN(n9411) );
  AOI21_X1 U11829 ( .B1(n13986), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9411), .ZN(
        n9412) );
  OAI211_X1 U11830 ( .C1(n9758), .C2(n14023), .A(n9413), .B(n9412), .ZN(
        P1_U3246) );
  NAND2_X1 U11831 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9417) );
  INV_X1 U11832 ( .A(n9414), .ZN(n9416) );
  AOI211_X1 U11833 ( .C1(n9417), .C2(n9416), .A(n9415), .B(n13980), .ZN(n9423)
         );
  INV_X1 U11834 ( .A(n9418), .ZN(n9421) );
  AOI211_X1 U11835 ( .C1(n9421), .C2(n9420), .A(n9419), .B(n14686), .ZN(n9422)
         );
  NOR2_X1 U11836 ( .A1(n9423), .A2(n9422), .ZN(n9425) );
  AOI22_X1 U11837 ( .A1(n13986), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9424) );
  OAI211_X1 U11838 ( .C1(n9606), .C2(n14023), .A(n9425), .B(n9424), .ZN(
        P1_U3244) );
  AOI211_X1 U11839 ( .C1(n9428), .C2(n9427), .A(n13980), .B(n9426), .ZN(n9436)
         );
  INV_X1 U11840 ( .A(n9429), .ZN(n9434) );
  NOR3_X1 U11841 ( .A1(n9432), .A2(n9431), .A3(n9430), .ZN(n9433) );
  NOR3_X1 U11842 ( .A1(n14686), .A2(n9434), .A3(n9433), .ZN(n9435) );
  NOR2_X1 U11843 ( .A1(n9436), .A2(n9435), .ZN(n9439) );
  INV_X1 U11844 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n11023) );
  NOR2_X1 U11845 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11023), .ZN(n9437) );
  AOI21_X1 U11846 ( .B1(n13986), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9437), .ZN(
        n9438) );
  OAI211_X1 U11847 ( .C1(n9440), .C2(n14023), .A(n9439), .B(n9438), .ZN(
        P1_U3249) );
  INV_X1 U11848 ( .A(n9441), .ZN(n9442) );
  INV_X1 U11849 ( .A(n11210), .ZN(n9448) );
  INV_X1 U11850 ( .A(n14869), .ZN(n11410) );
  OAI222_X1 U11851 ( .A1(n13798), .A2(n9444), .B1(n13817), .B2(n9448), .C1(
        n11410), .C2(P2_U3088), .ZN(P2_U3315) );
  NAND2_X1 U11852 ( .A1(n9446), .A2(n9445), .ZN(n10268) );
  NAND2_X1 U11853 ( .A1(n10268), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9599) );
  XNOR2_X1 U11854 ( .A(n9599), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11211) );
  INV_X1 U11855 ( .A(n11211), .ZN(n10553) );
  OAI222_X1 U11856 ( .A1(P1_U3086), .A2(n10553), .B1(n14391), .B2(n9448), .C1(
        n9447), .C2(n14396), .ZN(P1_U3343) );
  INV_X1 U11857 ( .A(n9546), .ZN(n9462) );
  INV_X1 U11858 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9449) );
  NAND2_X1 U11859 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14822) );
  INV_X1 U11860 ( .A(n14822), .ZN(n9450) );
  AOI22_X1 U11861 ( .A1(n14823), .A2(n9450), .B1(P2_REG1_REG_1__SCAN_IN), .B2(
        n6482), .ZN(n14836) );
  INV_X1 U11862 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9451) );
  MUX2_X1 U11863 ( .A(n9451), .B(P2_REG1_REG_2__SCAN_IN), .S(n9461), .Z(n14835) );
  NOR2_X1 U11864 ( .A1(n14836), .A2(n14835), .ZN(n14834) );
  AOI21_X1 U11865 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n9461), .A(n14834), .ZN(
        n9535) );
  INV_X1 U11866 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9452) );
  MUX2_X1 U11867 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9452), .S(n9546), .Z(n9534)
         );
  NOR2_X1 U11868 ( .A1(n9535), .A2(n9534), .ZN(n9533) );
  AOI21_X1 U11869 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n9462), .A(n9533), .ZN(
        n9523) );
  INV_X1 U11870 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9453) );
  MUX2_X1 U11871 ( .A(n9453), .B(P2_REG1_REG_4__SCAN_IN), .S(n9463), .Z(n9522)
         );
  NOR2_X1 U11872 ( .A1(n9523), .A2(n9522), .ZN(n9521) );
  INV_X1 U11873 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9454) );
  MUX2_X1 U11874 ( .A(n9454), .B(P2_REG1_REG_5__SCAN_IN), .S(n9550), .Z(n9456)
         );
  NAND2_X1 U11875 ( .A1(n9723), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13812) );
  OR2_X1 U11876 ( .A1(n9469), .A2(n13812), .ZN(n9458) );
  AOI211_X1 U11877 ( .C1(n9457), .C2(n9456), .A(n14901), .B(n9547), .ZN(n9474)
         );
  INV_X1 U11878 ( .A(n14910), .ZN(n14852) );
  INV_X1 U11879 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9460) );
  NOR3_X1 U11880 ( .A1(n14826), .A2(n9460), .A3(n9459), .ZN(n14827) );
  AOI21_X1 U11881 ( .B1(n6482), .B2(P2_REG2_REG_1__SCAN_IN), .A(n14827), .ZN(
        n14844) );
  INV_X1 U11882 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10465) );
  MUX2_X1 U11883 ( .A(n10465), .B(P2_REG2_REG_2__SCAN_IN), .S(n9461), .Z(
        n14843) );
  NOR2_X1 U11884 ( .A1(n14838), .A2(n10465), .ZN(n9538) );
  MUX2_X1 U11885 ( .A(n13653), .B(P2_REG2_REG_3__SCAN_IN), .S(n9546), .Z(n9537) );
  OAI21_X1 U11886 ( .B1(n14842), .B2(n9538), .A(n9537), .ZN(n9536) );
  NAND2_X1 U11887 ( .A1(n9462), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9525) );
  MUX2_X1 U11888 ( .A(n10349), .B(P2_REG2_REG_4__SCAN_IN), .S(n9463), .Z(n9524) );
  NOR2_X1 U11889 ( .A1(n9532), .A2(n10349), .ZN(n9465) );
  MUX2_X1 U11890 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10369), .S(n9550), .Z(n9464) );
  OAI21_X1 U11891 ( .B1(n9527), .B2(n9465), .A(n9464), .ZN(n9553) );
  INV_X1 U11892 ( .A(n9553), .ZN(n9467) );
  NOR3_X1 U11893 ( .A1(n9527), .A2(n9465), .A3(n9464), .ZN(n9466) );
  NOR3_X1 U11894 ( .A1(n14852), .A2(n9467), .A3(n9466), .ZN(n9473) );
  NAND2_X1 U11895 ( .A1(n9724), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9468) );
  NAND2_X1 U11896 ( .A1(n14821), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U11897 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10577) );
  OAI211_X1 U11898 ( .C1(n14839), .C2(n9471), .A(n9470), .B(n10577), .ZN(n9472) );
  OR3_X1 U11899 ( .A1(n9474), .A2(n9473), .A3(n9472), .ZN(P2_U3219) );
  INV_X1 U11900 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9476) );
  MUX2_X1 U11901 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9476), .S(n10834), .Z(n9477) );
  OAI21_X1 U11902 ( .B1(n9478), .B2(n9477), .A(n9667), .ZN(n9491) );
  INV_X1 U11903 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9479) );
  MUX2_X1 U11904 ( .A(n9479), .B(P1_REG2_REG_8__SCAN_IN), .S(n10834), .Z(n9482) );
  NOR2_X1 U11905 ( .A1(n9480), .A2(n9392), .ZN(n9484) );
  INV_X1 U11906 ( .A(n9484), .ZN(n9481) );
  NAND2_X1 U11907 ( .A1(n9482), .A2(n9481), .ZN(n9485) );
  MUX2_X1 U11908 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9479), .S(n10834), .Z(n9483) );
  OAI21_X1 U11909 ( .B1(n9486), .B2(n9484), .A(n9483), .ZN(n9664) );
  OAI211_X1 U11910 ( .C1(n9486), .C2(n9485), .A(n9664), .B(n14027), .ZN(n9488)
         );
  AND2_X1 U11911 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11365) );
  AOI21_X1 U11912 ( .B1(n13986), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n11365), .ZN(
        n9487) );
  OAI211_X1 U11913 ( .C1(n14023), .C2(n9489), .A(n9488), .B(n9487), .ZN(n9490)
         );
  AOI21_X1 U11914 ( .B1(n9491), .B2(n14680), .A(n9490), .ZN(n9492) );
  INV_X1 U11915 ( .A(n9492), .ZN(P1_U3251) );
  NAND2_X1 U11916 ( .A1(n7455), .A2(n14279), .ZN(n12263) );
  INV_X1 U11917 ( .A(n7455), .ZN(n13977) );
  INV_X1 U11918 ( .A(n12261), .ZN(n9493) );
  NAND2_X1 U11919 ( .A1(n12263), .A2(n9493), .ZN(n14283) );
  NAND2_X1 U11920 ( .A1(n9494), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9496) );
  INV_X1 U11921 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9495) );
  OAI21_X1 U11922 ( .B1(n12256), .B2(n12262), .A(n12020), .ZN(n10762) );
  OR2_X1 U11923 ( .A1(n10762), .A2(n14609), .ZN(n9877) );
  OR2_X1 U11924 ( .A1(n12461), .A2(n14150), .ZN(n14773) );
  NAND2_X1 U11925 ( .A1(n12254), .A2(n14609), .ZN(n9497) );
  INV_X1 U11926 ( .A(n12257), .ZN(n9578) );
  NAND2_X1 U11927 ( .A1(n12447), .A2(n9578), .ZN(n12450) );
  NAND2_X1 U11928 ( .A1(n14363), .A2(n14710), .ZN(n9503) );
  NOR3_X1 U11929 ( .A1(n10475), .A2(n12447), .A3(n12254), .ZN(n9502) );
  NAND2_X1 U11930 ( .A1(n12441), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n9501) );
  NAND2_X1 U11931 ( .A1(n9937), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n9500) );
  NAND2_X1 U11932 ( .A1(n12223), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U11933 ( .A1(n9936), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9498) );
  NAND4_X2 U11934 ( .A1(n9501), .A2(n9500), .A3(n9499), .A4(n9498), .ZN(n13976) );
  INV_X1 U11935 ( .A(n6479), .ZN(n13916) );
  NOR2_X1 U11936 ( .A1(n9680), .A2(n13916), .ZN(n14281) );
  AOI211_X1 U11937 ( .C1(n14283), .C2(n9503), .A(n9502), .B(n14281), .ZN(n9863) );
  OAI21_X1 U11938 ( .B1(n9583), .B2(P1_D_REG_1__SCAN_IN), .A(n9584), .ZN(n9515) );
  NOR4_X1 U11939 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n9507) );
  NOR4_X1 U11940 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n9506) );
  NOR4_X1 U11941 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n9505) );
  NOR4_X1 U11942 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n9504) );
  NAND4_X1 U11943 ( .A1(n9507), .A2(n9506), .A3(n9505), .A4(n9504), .ZN(n9513)
         );
  NOR2_X1 U11944 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .ZN(
        n9511) );
  NOR4_X1 U11945 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9510) );
  NOR4_X1 U11946 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9509) );
  NOR4_X1 U11947 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n9508) );
  NAND4_X1 U11948 ( .A1(n9511), .A2(n9510), .A3(n9509), .A4(n9508), .ZN(n9512)
         );
  NOR2_X1 U11949 ( .A1(n9513), .A2(n9512), .ZN(n9581) );
  OR2_X1 U11950 ( .A1(n9583), .A2(n9581), .ZN(n9514) );
  AND2_X1 U11951 ( .A1(n9515), .A2(n9514), .ZN(n9516) );
  NAND2_X1 U11952 ( .A1(n10488), .A2(n9516), .ZN(n9517) );
  NAND2_X1 U11953 ( .A1(n14770), .A2(n9617), .ZN(n9771) );
  OR2_X1 U11954 ( .A1(n9517), .A2(n12514), .ZN(n9862) );
  OR2_X1 U11955 ( .A1(n9583), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9519) );
  NAND2_X1 U11956 ( .A1(n14796), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9520) );
  OAI21_X1 U11957 ( .B1(n9863), .B2(n14796), .A(n9520), .ZN(P1_U3528) );
  AOI211_X1 U11958 ( .C1(n9523), .C2(n9522), .A(n9521), .B(n14901), .ZN(n9529)
         );
  AND3_X1 U11959 ( .A1(n9536), .A2(n9525), .A3(n9524), .ZN(n9526) );
  NOR3_X1 U11960 ( .A1(n14852), .A2(n9527), .A3(n9526), .ZN(n9528) );
  NOR2_X1 U11961 ( .A1(n9529), .A2(n9528), .ZN(n9531) );
  AND2_X1 U11962 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10434) );
  AOI21_X1 U11963 ( .B1(n14821), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n10434), .ZN(
        n9530) );
  OAI211_X1 U11964 ( .C1(n9532), .C2(n14839), .A(n9531), .B(n9530), .ZN(
        P2_U3218) );
  AOI211_X1 U11965 ( .C1(n9535), .C2(n9534), .A(n9533), .B(n14901), .ZN(n9542)
         );
  INV_X1 U11966 ( .A(n9536), .ZN(n9540) );
  NOR3_X1 U11967 ( .A1(n14842), .A2(n9538), .A3(n9537), .ZN(n9539) );
  NOR3_X1 U11968 ( .A1(n14852), .A2(n9540), .A3(n9539), .ZN(n9541) );
  NOR2_X1 U11969 ( .A1(n9542), .A2(n9541), .ZN(n9545) );
  INV_X1 U11970 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n15241) );
  NOR2_X1 U11971 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15241), .ZN(n9543) );
  AOI21_X1 U11972 ( .B1(n14821), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n9543), .ZN(
        n9544) );
  OAI211_X1 U11973 ( .C1(n9546), .C2(n14839), .A(n9545), .B(n9544), .ZN(
        P2_U3217) );
  MUX2_X1 U11974 ( .A(n14978), .B(P2_REG1_REG_6__SCAN_IN), .S(n9569), .Z(n9548) );
  AOI211_X1 U11975 ( .C1(n9549), .C2(n9548), .A(n14901), .B(n9564), .ZN(n9556)
         );
  NAND2_X1 U11976 ( .A1(n9550), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9552) );
  MUX2_X1 U11977 ( .A(n10390), .B(P2_REG2_REG_6__SCAN_IN), .S(n9569), .Z(n9551) );
  AOI21_X1 U11978 ( .B1(n9553), .B2(n9552), .A(n9551), .ZN(n9568) );
  AND3_X1 U11979 ( .A1(n9553), .A2(n9552), .A3(n9551), .ZN(n9554) );
  NOR3_X1 U11980 ( .A1(n14852), .A2(n9568), .A3(n9554), .ZN(n9555) );
  NOR2_X1 U11981 ( .A1(n9556), .A2(n9555), .ZN(n9559) );
  NAND2_X1 U11982 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10720) );
  INV_X1 U11983 ( .A(n10720), .ZN(n9557) );
  AOI21_X1 U11984 ( .B1(n14821), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9557), .ZN(
        n9558) );
  OAI211_X1 U11985 ( .C1(n9560), .C2(n14839), .A(n9559), .B(n9558), .ZN(
        P2_U3220) );
  INV_X1 U11986 ( .A(P3_DATAO_REG_10__SCAN_IN), .ZN(n15140) );
  NAND2_X1 U11987 ( .A1(P3_U3897), .A2(n11505), .ZN(n9561) );
  OAI21_X1 U11988 ( .B1(P3_U3897), .B2(n15140), .A(n9561), .ZN(P3_U3501) );
  INV_X1 U11989 ( .A(P3_DATAO_REG_6__SCAN_IN), .ZN(n15249) );
  NAND2_X1 U11990 ( .A1(n11134), .A2(P3_U3897), .ZN(n9562) );
  OAI21_X1 U11991 ( .B1(P3_U3897), .B2(n15249), .A(n9562), .ZN(P3_U3497) );
  INV_X1 U11992 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n15146) );
  NAND2_X1 U11993 ( .A1(n10032), .A2(P3_U3897), .ZN(n9563) );
  OAI21_X1 U11994 ( .B1(P3_U3897), .B2(n15146), .A(n9563), .ZN(P3_U3492) );
  AOI21_X1 U11995 ( .B1(n9569), .B2(P2_REG1_REG_6__SCAN_IN), .A(n9564), .ZN(
        n9566) );
  MUX2_X1 U11996 ( .A(n14980), .B(P2_REG1_REG_7__SCAN_IN), .S(n9850), .Z(n9565) );
  NOR2_X1 U11997 ( .A1(n9566), .A2(n9565), .ZN(n9846) );
  AOI211_X1 U11998 ( .C1(n9566), .C2(n9565), .A(n14901), .B(n9846), .ZN(n9567)
         );
  INV_X1 U11999 ( .A(n9567), .ZN(n9576) );
  AOI21_X1 U12000 ( .B1(n9569), .B2(P2_REG2_REG_6__SCAN_IN), .A(n9568), .ZN(
        n9571) );
  MUX2_X1 U12001 ( .A(n8663), .B(P2_REG2_REG_7__SCAN_IN), .S(n9850), .Z(n9570)
         );
  AOI21_X1 U12002 ( .B1(n9571), .B2(n9570), .A(n14852), .ZN(n9572) );
  OR2_X1 U12003 ( .A1(n9571), .A2(n9570), .ZN(n9853) );
  NAND2_X1 U12004 ( .A1(n9572), .A2(n9853), .ZN(n9573) );
  OAI21_X1 U12005 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n8657), .A(n9573), .ZN(
        n9574) );
  AOI21_X1 U12006 ( .B1(n14821), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n9574), .ZN(
        n9575) );
  OAI211_X1 U12007 ( .C1(n14839), .C2(n9577), .A(n9576), .B(n9575), .ZN(
        P2_U3221) );
  INV_X1 U12008 ( .A(n12447), .ZN(n11069) );
  NAND2_X1 U12009 ( .A1(n11069), .A2(n9578), .ZN(n12508) );
  INV_X1 U12010 ( .A(n12508), .ZN(n9580) );
  NAND2_X1 U12011 ( .A1(n9580), .A2(n9579), .ZN(n10495) );
  AND2_X1 U12012 ( .A1(n9581), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9582) );
  OR2_X1 U12013 ( .A1(n9583), .A2(n9582), .ZN(n9585) );
  AND2_X1 U12014 ( .A1(n9585), .A2(n9584), .ZN(n10486) );
  NAND2_X1 U12015 ( .A1(n9861), .A2(n10486), .ZN(n9588) );
  INV_X1 U12016 ( .A(n9588), .ZN(n9586) );
  NAND3_X1 U12017 ( .A1(n9586), .A2(n10489), .A3(n12462), .ZN(n9587) );
  NAND2_X1 U12018 ( .A1(n9588), .A2(n10488), .ZN(n9773) );
  INV_X1 U12019 ( .A(n14281), .ZN(n9591) );
  INV_X1 U12020 ( .A(n12514), .ZN(n9589) );
  NAND2_X1 U12021 ( .A1(n9589), .A2(n9773), .ZN(n9658) );
  NAND2_X1 U12022 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n9658), .ZN(n9590) );
  OAI21_X1 U12023 ( .B1(n13949), .B2(n9591), .A(n9590), .ZN(n9592) );
  AOI21_X1 U12024 ( .B1(n14279), .B2(n13952), .A(n9592), .ZN(n9593) );
  OAI21_X1 U12025 ( .B1(n9594), .B2(n13955), .A(n9593), .ZN(P1_U3232) );
  INV_X1 U12026 ( .A(n9595), .ZN(n9596) );
  OAI222_X1 U12027 ( .A1(P3_U3151), .A2(n6687), .B1(n13143), .B2(n9597), .C1(
        n6484), .C2(n9596), .ZN(P3_U3280) );
  INV_X1 U12028 ( .A(n11860), .ZN(n11412) );
  INV_X1 U12029 ( .A(n11214), .ZN(n9603) );
  OAI222_X1 U12030 ( .A1(P2_U3088), .A2(n11412), .B1(n13817), .B2(n9603), .C1(
        n9598), .C2(n13819), .ZN(P2_U3314) );
  NAND2_X1 U12031 ( .A1(n9599), .A2(n10265), .ZN(n9600) );
  NAND2_X1 U12032 ( .A1(n9600), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U12033 ( .A1(n9601), .A2(n10266), .ZN(n9842) );
  OR2_X1 U12034 ( .A1(n9601), .A2(n10266), .ZN(n9602) );
  INV_X1 U12035 ( .A(n11217), .ZN(n11010) );
  OAI222_X1 U12036 ( .A1(P1_U3086), .A2(n11010), .B1(n14391), .B2(n9603), .C1(
        n11215), .C2(n14396), .ZN(P1_U3342) );
  OR2_X1 U12037 ( .A1(n12141), .A2(n9604), .ZN(n9609) );
  OAI22_X1 U12038 ( .A1(n9680), .A2(n12230), .B1(n14729), .B2(n12231), .ZN(
        n9612) );
  XNOR2_X1 U12039 ( .A(n9612), .B(n12020), .ZN(n9647) );
  NAND2_X1 U12040 ( .A1(n13976), .A2(n12216), .ZN(n9614) );
  NAND2_X1 U12041 ( .A1(n9679), .A2(n9767), .ZN(n9613) );
  NAND2_X1 U12042 ( .A1(n9614), .A2(n9613), .ZN(n9646) );
  XNOR2_X1 U12043 ( .A(n9647), .B(n9646), .ZN(n9648) );
  XNOR2_X1 U12044 ( .A(n9649), .B(n9648), .ZN(n9615) );
  NAND2_X1 U12045 ( .A1(n9615), .A2(n13937), .ZN(n9625) );
  NAND2_X1 U12046 ( .A1(n9617), .A2(n9616), .ZN(n13917) );
  OR2_X1 U12047 ( .A1(n7455), .A2(n13917), .ZN(n9623) );
  NAND2_X1 U12048 ( .A1(n9937), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U12049 ( .A1(n12223), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9620) );
  NAND2_X1 U12050 ( .A1(n12441), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n9619) );
  NAND2_X1 U12051 ( .A1(n9936), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9618) );
  NAND4_X1 U12052 ( .A1(n9621), .A2(n9619), .A3(n9620), .A4(n9618), .ZN(n9682)
         );
  NAND2_X1 U12053 ( .A1(n13975), .A2(n6479), .ZN(n9622) );
  NAND2_X1 U12054 ( .A1(n9623), .A2(n9622), .ZN(n10482) );
  AOI22_X1 U12055 ( .A1(n13923), .A2(n10482), .B1(n9658), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n9624) );
  OAI211_X1 U12056 ( .C1(n14729), .C2(n13943), .A(n9625), .B(n9624), .ZN(
        P1_U3222) );
  AOI211_X1 U12057 ( .C1(n9628), .C2(n9627), .A(n9626), .B(n13980), .ZN(n9639)
         );
  INV_X1 U12058 ( .A(n9629), .ZN(n9634) );
  NOR3_X1 U12059 ( .A1(n9632), .A2(n9631), .A3(n9630), .ZN(n9633) );
  NOR3_X1 U12060 ( .A1(n14686), .A2(n9634), .A3(n9633), .ZN(n9638) );
  NAND2_X1 U12061 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10645) );
  NAND2_X1 U12062 ( .A1(n13986), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9635) );
  OAI211_X1 U12063 ( .C1(n14023), .C2(n9636), .A(n10645), .B(n9635), .ZN(n9637) );
  OR4_X1 U12064 ( .A1(n9640), .A2(n9639), .A3(n9638), .A4(n9637), .ZN(P1_U3247) );
  OAI22_X1 U12065 ( .A1(n9649), .A2(n9648), .B1(n9647), .B2(n9646), .ZN(n9763)
         );
  NAND2_X1 U12066 ( .A1(n13975), .A2(n12216), .ZN(n9651) );
  NAND2_X1 U12067 ( .A1(n10873), .A2(n9767), .ZN(n9650) );
  NAND2_X1 U12068 ( .A1(n9651), .A2(n9650), .ZN(n9759) );
  INV_X1 U12069 ( .A(n9682), .ZN(n9870) );
  OAI22_X1 U12070 ( .A1(n9870), .A2(n12230), .B1(n9869), .B2(n12231), .ZN(
        n9652) );
  XNOR2_X1 U12071 ( .A(n9652), .B(n12020), .ZN(n9760) );
  XOR2_X1 U12072 ( .A(n9759), .B(n9760), .Z(n9762) );
  XNOR2_X1 U12073 ( .A(n9763), .B(n9762), .ZN(n9653) );
  NAND2_X1 U12074 ( .A1(n9653), .A2(n13937), .ZN(n9661) );
  INV_X1 U12075 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U12076 ( .A1(n9937), .A2(n9776), .ZN(n9657) );
  NAND2_X1 U12077 ( .A1(n12441), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9656) );
  NAND2_X1 U12078 ( .A1(n12223), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9655) );
  NAND2_X1 U12079 ( .A1(n9936), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9654) );
  AOI22_X1 U12080 ( .A1(n14064), .A2(n13976), .B1(n13974), .B2(n6479), .ZN(
        n9687) );
  INV_X1 U12081 ( .A(n9687), .ZN(n9659) );
  AOI22_X1 U12082 ( .A1(n9659), .A2(n13923), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9658), .ZN(n9660) );
  OAI211_X1 U12083 ( .C1(n9869), .C2(n13943), .A(n9661), .B(n9660), .ZN(
        P1_U3237) );
  NAND2_X1 U12084 ( .A1(n10834), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9663) );
  INV_X1 U12085 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10865) );
  MUX2_X1 U12086 ( .A(n10865), .B(P1_REG2_REG_9__SCAN_IN), .S(n10840), .Z(
        n9662) );
  AOI21_X1 U12087 ( .B1(n9664), .B2(n9663), .A(n9662), .ZN(n9990) );
  NAND3_X1 U12088 ( .A1(n9664), .A2(n9663), .A3(n9662), .ZN(n9665) );
  NAND2_X1 U12089 ( .A1(n9665), .A2(n14027), .ZN(n9675) );
  INV_X1 U12090 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9666) );
  MUX2_X1 U12091 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9666), .S(n10840), .Z(n9669) );
  OAI21_X1 U12092 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10834), .A(n9667), .ZN(
        n9668) );
  NAND2_X1 U12093 ( .A1(n9668), .A2(n9669), .ZN(n9980) );
  OAI21_X1 U12094 ( .B1(n9669), .B2(n9668), .A(n9980), .ZN(n9670) );
  NAND2_X1 U12095 ( .A1(n9670), .A2(n14680), .ZN(n9674) );
  NAND2_X1 U12096 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11428) );
  INV_X1 U12097 ( .A(n11428), .ZN(n9672) );
  NOR2_X1 U12098 ( .A1(n14023), .A2(n9984), .ZN(n9671) );
  AOI211_X1 U12099 ( .C1(n13986), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n9672), .B(
        n9671), .ZN(n9673) );
  OAI211_X1 U12100 ( .C1(n9990), .C2(n9675), .A(n9674), .B(n9673), .ZN(
        P1_U3252) );
  INV_X1 U12101 ( .A(n9676), .ZN(n9677) );
  OAI222_X1 U12102 ( .A1(P3_U3151), .A2(n12783), .B1(n13143), .B2(n9678), .C1(
        n6484), .C2(n9677), .ZN(P3_U3279) );
  NAND2_X1 U12103 ( .A1(n13976), .A2(n14729), .ZN(n12260) );
  NAND2_X1 U12104 ( .A1(n12259), .A2(n12260), .ZN(n10477) );
  OR2_X1 U12105 ( .A1(n7455), .A2(n10475), .ZN(n10481) );
  NAND2_X1 U12106 ( .A1(n10477), .A2(n10481), .ZN(n10480) );
  NAND2_X1 U12107 ( .A1(n9680), .A2(n14729), .ZN(n9681) );
  NAND2_X1 U12108 ( .A1(n10480), .A2(n9681), .ZN(n9683) );
  NAND2_X1 U12109 ( .A1(n9870), .A2(n10873), .ZN(n12270) );
  NAND2_X1 U12110 ( .A1(n9682), .A2(n9869), .ZN(n12277) );
  NAND2_X1 U12111 ( .A1(n9683), .A2(n9878), .ZN(n9872) );
  OAI21_X1 U12112 ( .B1(n9683), .B2(n9878), .A(n9872), .ZN(n10877) );
  NAND2_X1 U12113 ( .A1(n10475), .A2(n14729), .ZN(n10474) );
  NOR2_X2 U12114 ( .A1(n10474), .A2(n10873), .ZN(n9875) );
  NAND2_X1 U12115 ( .A1(n10474), .A2(n10873), .ZN(n9684) );
  NAND2_X1 U12116 ( .A1(n9684), .A2(n14749), .ZN(n9685) );
  OR2_X1 U12117 ( .A1(n9875), .A2(n9685), .ZN(n10875) );
  OAI21_X1 U12118 ( .B1(n9869), .B2(n14780), .A(n10875), .ZN(n9689) );
  INV_X1 U12119 ( .A(n12263), .ZN(n9686) );
  NAND2_X1 U12120 ( .A1(n9686), .A2(n12260), .ZN(n12265) );
  XNOR2_X1 U12121 ( .A(n9878), .B(n9880), .ZN(n9688) );
  OAI21_X1 U12122 ( .B1(n9688), .B2(n14710), .A(n9687), .ZN(n10870) );
  AOI211_X1 U12123 ( .C1(n14784), .C2(n10877), .A(n9689), .B(n10870), .ZN(
        n9866) );
  NAND2_X1 U12124 ( .A1(n14796), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9690) );
  OAI21_X1 U12125 ( .B1(n9866), .B2(n14796), .A(n9690), .ZN(P1_U3530) );
  INV_X1 U12126 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10010) );
  INV_X1 U12127 ( .A(n9693), .ZN(n9691) );
  NAND2_X1 U12128 ( .A1(n9692), .A2(n9691), .ZN(n9697) );
  INV_X1 U12129 ( .A(n9907), .ZN(n9694) );
  OAI21_X1 U12130 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(n9696) );
  AND2_X1 U12131 ( .A1(n9697), .A2(n9696), .ZN(n9698) );
  AND2_X1 U12132 ( .A1(n15023), .A2(n15065), .ZN(n9700) );
  NOR3_X1 U12133 ( .A1(n9926), .A2(n15065), .A3(n9701), .ZN(n9702) );
  AOI21_X1 U12134 ( .B1(n13022), .B2(n10032), .A(n9702), .ZN(n10081) );
  INV_X1 U12135 ( .A(n10081), .ZN(n9703) );
  NAND2_X1 U12136 ( .A1(n9703), .A2(n15030), .ZN(n9707) );
  OR2_X1 U12137 ( .A1(n15023), .A2(n15079), .ZN(n9704) );
  INV_X1 U12138 ( .A(n13031), .ZN(n15016) );
  AOI22_X1 U12139 ( .A1(n15016), .A2(n9923), .B1(n15014), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n9706) );
  OAI211_X1 U12140 ( .C1(n10010), .C2(n15030), .A(n9707), .B(n9706), .ZN(
        P3_U3233) );
  AND2_X1 U12141 ( .A1(n9710), .A2(n11348), .ZN(n9711) );
  INV_X1 U12142 ( .A(n14972), .ZN(n14942) );
  NAND2_X1 U12143 ( .A1(n9828), .A2(n9713), .ZN(n9714) );
  OAI21_X1 U12144 ( .B1(n9714), .B2(n9719), .A(n9889), .ZN(n10470) );
  NAND2_X1 U12145 ( .A1(n10110), .A2(n9831), .ZN(n9830) );
  NOR2_X2 U12146 ( .A1(n9830), .A2(n10065), .ZN(n9898) );
  NAND2_X1 U12147 ( .A1(n9830), .A2(n10065), .ZN(n9715) );
  NAND2_X1 U12148 ( .A1(n11348), .A2(n11111), .ZN(n9804) );
  NAND2_X1 U12149 ( .A1(n9715), .A2(n13521), .ZN(n9716) );
  NOR2_X1 U12150 ( .A1(n9898), .A2(n9716), .ZN(n10469) );
  INV_X1 U12151 ( .A(n9832), .ZN(n9819) );
  NAND2_X1 U12152 ( .A1(n9819), .A2(n9712), .ZN(n9718) );
  INV_X1 U12153 ( .A(n13359), .ZN(n9822) );
  NAND2_X1 U12154 ( .A1(n9822), .A2(n6481), .ZN(n9717) );
  NAND2_X1 U12155 ( .A1(n9718), .A2(n9717), .ZN(n9893) );
  XNOR2_X1 U12156 ( .A(n9893), .B(n9719), .ZN(n9725) );
  INV_X1 U12157 ( .A(n9720), .ZN(n9722) );
  OR2_X1 U12158 ( .A1(n6485), .A2(n11111), .ZN(n9721) );
  INV_X1 U12159 ( .A(n9789), .ZN(n9749) );
  NAND2_X1 U12160 ( .A1(n9749), .A2(n9723), .ZN(n13575) );
  NAND2_X1 U12161 ( .A1(n9749), .A2(n9724), .ZN(n13631) );
  AOI22_X1 U12162 ( .A1(n13628), .A2(n13359), .B1(n13357), .B2(n13466), .ZN(
        n9810) );
  OAI21_X1 U12163 ( .B1(n9725), .B2(n13603), .A(n9810), .ZN(n10464) );
  AOI211_X1 U12164 ( .C1(n14951), .C2(n10470), .A(n10469), .B(n10464), .ZN(
        n10067) );
  XNOR2_X1 U12165 ( .A(n11537), .B(P2_B_REG_SCAN_IN), .ZN(n9726) );
  INV_X1 U12166 ( .A(n11908), .ZN(n9742) );
  NOR2_X1 U12167 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .ZN(
        n9731) );
  NOR4_X1 U12168 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n9730) );
  NOR4_X1 U12169 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9729) );
  NOR4_X1 U12170 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n9728) );
  AND4_X1 U12171 ( .A1(n9731), .A2(n9730), .A3(n9729), .A4(n9728), .ZN(n9737)
         );
  NOR4_X1 U12172 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n9735) );
  NOR4_X1 U12173 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n9734) );
  NOR4_X1 U12174 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9733) );
  NOR4_X1 U12175 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n9732) );
  AND4_X1 U12176 ( .A1(n9735), .A2(n9734), .A3(n9733), .A4(n9732), .ZN(n9736)
         );
  NAND2_X1 U12177 ( .A1(n9737), .A2(n9736), .ZN(n9738) );
  AND2_X1 U12178 ( .A1(n14917), .A2(n9738), .ZN(n9799) );
  INV_X1 U12179 ( .A(n9799), .ZN(n10047) );
  INV_X1 U12180 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14923) );
  NAND2_X1 U12181 ( .A1(n14917), .A2(n14923), .ZN(n9741) );
  INV_X1 U12182 ( .A(n9739), .ZN(n11730) );
  NAND2_X1 U12183 ( .A1(n11730), .A2(n11908), .ZN(n9740) );
  NAND2_X1 U12184 ( .A1(n9741), .A2(n9740), .ZN(n14924) );
  NAND2_X1 U12185 ( .A1(n14972), .A2(n11111), .ZN(n9805) );
  NAND3_X1 U12186 ( .A1(n10047), .A2(n14924), .A3(n9805), .ZN(n9966) );
  INV_X1 U12187 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14921) );
  NAND2_X1 U12188 ( .A1(n14917), .A2(n14921), .ZN(n9744) );
  OR2_X1 U12189 ( .A1(n11537), .A2(n9742), .ZN(n9743) );
  NAND2_X1 U12190 ( .A1(n9744), .A2(n9743), .ZN(n10048) );
  INV_X1 U12191 ( .A(n10048), .ZN(n9750) );
  OR2_X1 U12192 ( .A1(n9745), .A2(n11908), .ZN(n9748) );
  INV_X1 U12193 ( .A(n9746), .ZN(n9747) );
  NAND2_X1 U12194 ( .A1(n9751), .A2(n9749), .ZN(n9964) );
  NAND2_X1 U12195 ( .A1(n14925), .A2(n9964), .ZN(n10046) );
  OAI22_X1 U12196 ( .A1(n13794), .A2(n10466), .B1(n14974), .B2(n8564), .ZN(
        n9752) );
  INV_X1 U12197 ( .A(n9752), .ZN(n9753) );
  OAI21_X1 U12198 ( .B1(n10067), .B2(n14973), .A(n9753), .ZN(P2_U3436) );
  OR2_X1 U12199 ( .A1(n12458), .A2(n9755), .ZN(n9756) );
  INV_X1 U12200 ( .A(n12268), .ZN(n12280) );
  NAND2_X1 U12201 ( .A1(n13974), .A2(n9767), .ZN(n9765) );
  NAND2_X1 U12202 ( .A1(n12268), .A2(n12205), .ZN(n9764) );
  NAND2_X1 U12203 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  XNOR2_X1 U12204 ( .A(n9766), .B(n12020), .ZN(n10648) );
  AOI22_X1 U12205 ( .A1(n13974), .A2(n12216), .B1(n12175), .B2(n12268), .ZN(
        n10650) );
  XNOR2_X1 U12206 ( .A(n10648), .B(n10650), .ZN(n9768) );
  NAND2_X1 U12207 ( .A1(n9769), .A2(n9768), .ZN(n10651) );
  OAI211_X1 U12208 ( .C1(n9769), .C2(n9768), .A(n10651), .B(n13937), .ZN(n9787) );
  AND2_X1 U12209 ( .A1(n9771), .A2(n9770), .ZN(n9772) );
  NAND2_X1 U12210 ( .A1(n9773), .A2(n9772), .ZN(n9774) );
  NAND2_X1 U12211 ( .A1(n13975), .A2(n14064), .ZN(n9783) );
  NAND2_X1 U12212 ( .A1(n9936), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U12213 ( .A1(n12223), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9780) );
  INV_X1 U12214 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U12215 ( .A1(n9776), .A2(n9775), .ZN(n9777) );
  NAND2_X1 U12216 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9939) );
  AND2_X1 U12217 ( .A1(n9777), .A2(n9939), .ZN(n10807) );
  NAND2_X1 U12218 ( .A1(n9937), .A2(n10807), .ZN(n9779) );
  NAND2_X1 U12219 ( .A1(n12441), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9778) );
  NAND4_X1 U12220 ( .A1(n9781), .A2(n9780), .A3(n9779), .A4(n9778), .ZN(n13973) );
  NAND2_X1 U12221 ( .A1(n13973), .A2(n6479), .ZN(n9782) );
  NAND2_X1 U12222 ( .A1(n9783), .A2(n9782), .ZN(n9882) );
  INV_X1 U12223 ( .A(n9882), .ZN(n9784) );
  OAI22_X1 U12224 ( .A1(n13949), .A2(n9784), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9776), .ZN(n9785) );
  AOI21_X1 U12225 ( .B1(n9776), .B2(n13947), .A(n9785), .ZN(n9786) );
  OAI211_X1 U12226 ( .C1(n12280), .C2(n13943), .A(n9787), .B(n9786), .ZN(
        P1_U3218) );
  INV_X1 U12227 ( .A(n14925), .ZN(n14922) );
  OR2_X1 U12228 ( .A1(n14924), .A2(n9799), .ZN(n9788) );
  AND2_X1 U12229 ( .A1(n14967), .A2(n9789), .ZN(n9790) );
  NAND2_X2 U12230 ( .A1(n9809), .A2(n9790), .ZN(n14808) );
  NAND2_X2 U12231 ( .A1(n9792), .A2(n9791), .ZN(n9794) );
  NAND2_X1 U12232 ( .A1(n13359), .A2(n9793), .ZN(n9796) );
  NOR2_X1 U12233 ( .A1(n9827), .A2(n13521), .ZN(n9795) );
  NOR2_X1 U12234 ( .A1(n13222), .A2(n10060), .ZN(n10111) );
  NAND2_X1 U12235 ( .A1(n9812), .A2(n9796), .ZN(n9797) );
  NAND2_X1 U12236 ( .A1(n9814), .A2(n9797), .ZN(n9798) );
  XNOR2_X1 U12237 ( .A(n13222), .B(n10065), .ZN(n10417) );
  NAND2_X1 U12238 ( .A1(n13358), .A2(n13221), .ZN(n10418) );
  XNOR2_X1 U12239 ( .A(n10417), .B(n10418), .ZN(n9813) );
  NAND2_X1 U12240 ( .A1(n9798), .A2(n9813), .ZN(n10421) );
  OR3_X1 U12241 ( .A1(n9799), .A2(n14924), .A3(n10048), .ZN(n9800) );
  NAND2_X1 U12242 ( .A1(n9800), .A2(n9805), .ZN(n9803) );
  AND2_X1 U12243 ( .A1(n9801), .A2(n9964), .ZN(n9802) );
  NAND2_X1 U12244 ( .A1(n9803), .A2(n9802), .ZN(n10431) );
  OR2_X1 U12245 ( .A1(n10431), .A2(P2_U3088), .ZN(n10118) );
  NOR2_X1 U12246 ( .A1(n6485), .A2(n9804), .ZN(n10059) );
  NAND2_X1 U12247 ( .A1(n9809), .A2(n10059), .ZN(n9807) );
  INV_X1 U12248 ( .A(n9805), .ZN(n9806) );
  NAND2_X1 U12249 ( .A1(n9809), .A2(n9808), .ZN(n13282) );
  OAI22_X1 U12250 ( .A1(n13321), .A2(n10466), .B1(n9810), .B2(n13282), .ZN(
        n9811) );
  AOI21_X1 U12251 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n10118), .A(n9811), .ZN(
        n9818) );
  OAI22_X1 U12252 ( .A1(n13329), .A2(n9822), .B1(n9812), .B2(n14808), .ZN(
        n9816) );
  INV_X1 U12253 ( .A(n9813), .ZN(n9815) );
  NAND3_X1 U12254 ( .A1(n9816), .A2(n9815), .A3(n9814), .ZN(n9817) );
  OAI211_X1 U12255 ( .C1(n14808), .C2(n10421), .A(n9818), .B(n9817), .ZN(
        P2_U3209) );
  AOI21_X1 U12256 ( .B1(n10060), .B2(n13521), .A(n9819), .ZN(n9820) );
  OAI22_X1 U12257 ( .A1(n13321), .A2(n9831), .B1(n9820), .B2(n14808), .ZN(
        n9824) );
  OAI22_X1 U12258 ( .A1(n9822), .A2(n14800), .B1(n13329), .B2(n9821), .ZN(
        n9823) );
  AOI211_X1 U12259 ( .C1(P2_REG3_REG_0__SCAN_IN), .C2(n10118), .A(n9824), .B(
        n9823), .ZN(n9825) );
  INV_X1 U12260 ( .A(n9825), .ZN(P2_U3204) );
  INV_X1 U12261 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n15232) );
  NAND2_X1 U12262 ( .A1(n12976), .A2(P3_U3897), .ZN(n9826) );
  OAI21_X1 U12263 ( .B1(P3_U3897), .B2(n15232), .A(n9826), .ZN(P3_U3512) );
  INV_X1 U12264 ( .A(n9828), .ZN(n9829) );
  AOI21_X1 U12265 ( .B1(n10112), .B2(n6618), .A(n9829), .ZN(n10451) );
  OAI211_X1 U12266 ( .C1(n10110), .C2(n9831), .A(n13521), .B(n9830), .ZN(
        n10444) );
  OAI21_X1 U12267 ( .B1(n10451), .B2(n13751), .A(n10444), .ZN(n9834) );
  XNOR2_X1 U12268 ( .A(n6618), .B(n9832), .ZN(n9833) );
  OAI21_X1 U12269 ( .B1(n9833), .B2(n13603), .A(n10109), .ZN(n10448) );
  NOR2_X1 U12270 ( .A1(n9834), .A2(n10448), .ZN(n9997) );
  INV_X1 U12271 ( .A(n13794), .ZN(n9835) );
  AOI22_X1 U12272 ( .A1(n9835), .A2(n6481), .B1(n14973), .B2(
        P2_REG0_REG_1__SCAN_IN), .ZN(n9836) );
  OAI21_X1 U12273 ( .B1(n9997), .B2(n14973), .A(n9836), .ZN(P2_U3433) );
  INV_X1 U12274 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10005) );
  MUX2_X1 U12275 ( .A(n10005), .B(n10081), .S(n15106), .Z(n9837) );
  OAI21_X1 U12276 ( .B1(n10084), .B2(n13087), .A(n9837), .ZN(P3_U3459) );
  INV_X1 U12277 ( .A(n12813), .ZN(n12800) );
  INV_X1 U12278 ( .A(n9838), .ZN(n9839) );
  OAI222_X1 U12279 ( .A1(P3_U3151), .A2(n12800), .B1(n13143), .B2(n9840), .C1(
        n6484), .C2(n9839), .ZN(P3_U3278) );
  INV_X1 U12280 ( .A(n14882), .ZN(n11853) );
  INV_X1 U12281 ( .A(n11479), .ZN(n9845) );
  OAI222_X1 U12282 ( .A1(P2_U3088), .A2(n11853), .B1(n13817), .B2(n9845), .C1(
        n9841), .C2(n13819), .ZN(P2_U3313) );
  NAND2_X1 U12283 ( .A1(n9842), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9843) );
  XNOR2_X1 U12284 ( .A(n9843), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11745) );
  INV_X1 U12285 ( .A(n11745), .ZN(n11126) );
  OAI222_X1 U12286 ( .A1(P1_U3086), .A2(n11126), .B1(n14391), .B2(n9845), .C1(
        n9844), .C2(n14396), .ZN(P1_U3341) );
  INV_X1 U12287 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9847) );
  MUX2_X1 U12288 ( .A(n9847), .B(P2_REG1_REG_8__SCAN_IN), .S(n10126), .Z(n9848) );
  AOI211_X1 U12289 ( .C1(n9849), .C2(n9848), .A(n14901), .B(n10120), .ZN(n9860) );
  NAND2_X1 U12290 ( .A1(n9850), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9852) );
  MUX2_X1 U12291 ( .A(n10742), .B(P2_REG2_REG_8__SCAN_IN), .S(n10126), .Z(
        n9851) );
  AND3_X1 U12292 ( .A1(n9853), .A2(n9852), .A3(n9851), .ZN(n9854) );
  NOR3_X1 U12293 ( .A1(n10125), .A2(n9854), .A3(n14852), .ZN(n9859) );
  NOR2_X1 U12294 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10927), .ZN(n9855) );
  AOI21_X1 U12295 ( .B1(n14821), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n9855), .ZN(
        n9856) );
  OAI21_X1 U12296 ( .B1(n9857), .B2(n14839), .A(n9856), .ZN(n9858) );
  OR3_X1 U12297 ( .A1(n9860), .A2(n9859), .A3(n9858), .ZN(P2_U3222) );
  INV_X2 U12298 ( .A(n14785), .ZN(n14748) );
  INV_X1 U12299 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9865) );
  OR2_X1 U12300 ( .A1(n9863), .A2(n14785), .ZN(n9864) );
  OAI21_X1 U12301 ( .B1(n14748), .B2(n9865), .A(n9864), .ZN(P1_U3459) );
  INV_X1 U12302 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9868) );
  OR2_X1 U12303 ( .A1(n9866), .A2(n14785), .ZN(n9867) );
  OAI21_X1 U12304 ( .B1(n14748), .B2(n9868), .A(n9867), .ZN(P1_U3465) );
  INV_X1 U12305 ( .A(n14773), .ZN(n14754) );
  NAND2_X1 U12306 ( .A1(n9870), .A2(n9869), .ZN(n9871) );
  NAND2_X1 U12307 ( .A1(n9872), .A2(n9871), .ZN(n9873) );
  XNOR2_X2 U12308 ( .A(n13974), .B(n12268), .ZN(n12279) );
  INV_X1 U12309 ( .A(n12279), .ZN(n12470) );
  OR2_X1 U12310 ( .A1(n9873), .A2(n12470), .ZN(n9874) );
  NAND2_X1 U12311 ( .A1(n9928), .A2(n9874), .ZN(n10509) );
  NOR2_X1 U12312 ( .A1(n9875), .A2(n12280), .ZN(n9876) );
  OR2_X1 U12313 ( .A1(n9947), .A2(n9876), .ZN(n10512) );
  OAI22_X1 U12314 ( .A1(n10512), .A2(n14294), .B1(n12280), .B2(n14780), .ZN(
        n9886) );
  INV_X1 U12315 ( .A(n9877), .ZN(n14777) );
  NAND2_X1 U12316 ( .A1(n10509), .A2(n14777), .ZN(n9885) );
  INV_X1 U12317 ( .A(n9878), .ZN(n9879) );
  OAI21_X1 U12318 ( .B1(n9881), .B2(n12279), .A(n9934), .ZN(n9883) );
  AOI21_X1 U12319 ( .B1(n9883), .B2(n14770), .A(n9882), .ZN(n9884) );
  NAND2_X1 U12320 ( .A1(n9885), .A2(n9884), .ZN(n10510) );
  AOI211_X1 U12321 ( .C1(n14754), .C2(n10509), .A(n9886), .B(n10510), .ZN(
        n9976) );
  NAND2_X1 U12322 ( .A1(n14796), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9887) );
  OAI21_X1 U12323 ( .B1(n9976), .B2(n14796), .A(n9887), .ZN(P1_U3531) );
  INV_X1 U12324 ( .A(n13358), .ZN(n9896) );
  NAND2_X1 U12325 ( .A1(n9896), .A2(n10466), .ZN(n9888) );
  NAND2_X1 U12326 ( .A1(n9889), .A2(n9888), .ZN(n9890) );
  NAND2_X1 U12327 ( .A1(n9890), .A2(n9891), .ZN(n9952) );
  OAI21_X1 U12328 ( .B1(n9890), .B2(n9891), .A(n9952), .ZN(n13657) );
  INV_X1 U12329 ( .A(n13657), .ZN(n9899) );
  NAND2_X1 U12330 ( .A1(n9893), .A2(n9892), .ZN(n9895) );
  NAND2_X1 U12331 ( .A1(n9896), .A2(n10065), .ZN(n9894) );
  NAND2_X1 U12332 ( .A1(n9895), .A2(n9894), .ZN(n9957) );
  XNOR2_X1 U12333 ( .A(n9956), .B(n9957), .ZN(n9897) );
  INV_X1 U12334 ( .A(n13356), .ZN(n10361) );
  OAI22_X1 U12335 ( .A1(n10361), .A2(n13631), .B1(n9896), .B2(n13575), .ZN(
        n10500) );
  AOI21_X1 U12336 ( .B1(n9897), .B2(n13625), .A(n10500), .ZN(n13652) );
  NAND2_X1 U12337 ( .A1(n9898), .A2(n10502), .ZN(n9954) );
  OAI211_X1 U12338 ( .C1(n9898), .C2(n10502), .A(n13521), .B(n9954), .ZN(
        n13658) );
  OAI211_X1 U12339 ( .C1(n9899), .C2(n13751), .A(n13652), .B(n13658), .ZN(
        n9974) );
  OAI22_X1 U12340 ( .A1(n13794), .A2(n10502), .B1(n14974), .B2(n8588), .ZN(
        n9900) );
  AOI21_X1 U12341 ( .B1(n9974), .B2(n14974), .A(n9900), .ZN(n9901) );
  INV_X1 U12342 ( .A(n9901), .ZN(P2_U3439) );
  NAND3_X1 U12343 ( .A1(n9921), .A2(n9906), .A3(n15079), .ZN(n9904) );
  NAND2_X1 U12344 ( .A1(n9902), .A2(n9909), .ZN(n9903) );
  NAND2_X1 U12345 ( .A1(n9904), .A2(n9903), .ZN(n9905) );
  INV_X1 U12346 ( .A(n9906), .ZN(n9912) );
  AND3_X1 U12347 ( .A1(n9908), .A2(n10000), .A3(n9907), .ZN(n9911) );
  NAND2_X1 U12348 ( .A1(n9918), .A2(n9909), .ZN(n9910) );
  OAI211_X1 U12349 ( .C1(n9921), .C2(n9912), .A(n9911), .B(n9910), .ZN(n9913)
         );
  NAND2_X1 U12350 ( .A1(n9913), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9916) );
  INV_X1 U12351 ( .A(n9917), .ZN(n9914) );
  NAND2_X1 U12352 ( .A1(n9914), .A2(n9918), .ZN(n9915) );
  NAND2_X1 U12353 ( .A1(n12672), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10075) );
  NAND2_X1 U12354 ( .A1(n10075), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n9925) );
  NOR2_X1 U12355 ( .A1(n9918), .A2(n9917), .ZN(n10041) );
  AND2_X1 U12356 ( .A1(n9998), .A2(n15065), .ZN(n9920) );
  NAND2_X1 U12357 ( .A1(n9921), .A2(n9920), .ZN(n9922) );
  AOI22_X1 U12358 ( .A1(n12649), .A2(n10032), .B1(n9923), .B2(n6477), .ZN(
        n9924) );
  OAI211_X1 U12359 ( .C1(n9926), .C2(n12689), .A(n9925), .B(n9924), .ZN(
        P3_U3172) );
  INV_X1 U12360 ( .A(n13974), .ZN(n12269) );
  NAND2_X1 U12361 ( .A1(n12269), .A2(n12280), .ZN(n9927) );
  NAND2_X1 U12362 ( .A1(n9928), .A2(n9927), .ZN(n10586) );
  NAND2_X1 U12363 ( .A1(n9929), .A2(n12457), .ZN(n9932) );
  XNOR2_X1 U12364 ( .A(n13973), .B(n12287), .ZN(n12472) );
  XOR2_X1 U12365 ( .A(n10586), .B(n12472), .Z(n10815) );
  NAND2_X1 U12366 ( .A1(n12269), .A2(n12268), .ZN(n9933) );
  XNOR2_X1 U12367 ( .A(n10616), .B(n12472), .ZN(n9935) );
  NAND2_X1 U12368 ( .A1(n9935), .A2(n14770), .ZN(n10811) );
  NAND2_X1 U12369 ( .A1(n12440), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9944) );
  NAND2_X1 U12370 ( .A1(n12439), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9943) );
  AND2_X1 U12371 ( .A1(n9939), .A2(n9938), .ZN(n9940) );
  NOR2_X1 U12372 ( .A1(n10596), .A2(n9940), .ZN(n10772) );
  NAND2_X1 U12373 ( .A1(n9937), .A2(n10772), .ZN(n9942) );
  NAND2_X1 U12374 ( .A1(n12441), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9941) );
  AND4_X2 U12375 ( .A1(n9944), .A2(n9943), .A3(n9942), .A4(n9941), .ZN(n12293)
         );
  OR2_X1 U12376 ( .A1(n12293), .A2(n13916), .ZN(n9946) );
  NAND2_X1 U12377 ( .A1(n13974), .A2(n14064), .ZN(n9945) );
  AND2_X1 U12378 ( .A1(n9946), .A2(n9945), .ZN(n10810) );
  OAI211_X1 U12379 ( .C1(n9947), .C2(n12285), .A(n14749), .B(n10771), .ZN(
        n10809) );
  NAND2_X1 U12380 ( .A1(n14735), .A2(n12287), .ZN(n9948) );
  NAND4_X1 U12381 ( .A1(n10811), .A2(n10810), .A3(n10809), .A4(n9948), .ZN(
        n9949) );
  AOI21_X1 U12382 ( .B1(n10815), .B2(n14784), .A(n9949), .ZN(n10080) );
  NAND2_X1 U12383 ( .A1(n14796), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9950) );
  OAI21_X1 U12384 ( .B1(n10080), .B2(n14796), .A(n9950), .ZN(P1_U3532) );
  NAND2_X1 U12385 ( .A1(n7226), .A2(n10502), .ZN(n9951) );
  OAI21_X1 U12386 ( .B1(n9953), .B2(n10358), .A(n10357), .ZN(n10346) );
  AOI21_X1 U12387 ( .B1(n9954), .B2(n10433), .A(n9793), .ZN(n9955) );
  OR2_X1 U12388 ( .A1(n9954), .A2(n10433), .ZN(n10371) );
  AND2_X1 U12389 ( .A1(n9955), .A2(n10371), .ZN(n10351) );
  NAND2_X1 U12390 ( .A1(n7226), .A2(n9108), .ZN(n9958) );
  XNOR2_X1 U12391 ( .A(n10360), .B(n10358), .ZN(n9961) );
  NAND2_X1 U12392 ( .A1(n13357), .A2(n13628), .ZN(n9960) );
  NAND2_X1 U12393 ( .A1(n13355), .A2(n13466), .ZN(n9959) );
  AND2_X1 U12394 ( .A1(n9960), .A2(n9959), .ZN(n10437) );
  OAI21_X1 U12395 ( .B1(n9961), .B2(n13603), .A(n10437), .ZN(n10347) );
  AOI211_X1 U12396 ( .C1(n14951), .C2(n10346), .A(n10351), .B(n10347), .ZN(
        n9969) );
  OAI22_X1 U12397 ( .A1(n13794), .A2(n10355), .B1(n14974), .B2(n8599), .ZN(
        n9962) );
  INV_X1 U12398 ( .A(n9962), .ZN(n9963) );
  OAI21_X1 U12399 ( .B1(n9969), .B2(n14973), .A(n9963), .ZN(P2_U3442) );
  INV_X1 U12400 ( .A(n9964), .ZN(n9965) );
  OAI22_X1 U12401 ( .A1(n13755), .A2(n10355), .B1(n14986), .B2(n9453), .ZN(
        n9967) );
  INV_X1 U12402 ( .A(n9967), .ZN(n9968) );
  OAI21_X1 U12403 ( .B1(n9969), .B2(n14984), .A(n9968), .ZN(P2_U3503) );
  INV_X1 U12404 ( .A(n12841), .ZN(n9972) );
  OAI222_X1 U12405 ( .A1(P3_U3151), .A2(n9972), .B1(n13143), .B2(n9971), .C1(
        n6484), .C2(n9970), .ZN(P3_U3277) );
  OAI22_X1 U12406 ( .A1(n13755), .A2(n10502), .B1(n14986), .B2(n9452), .ZN(
        n9973) );
  AOI21_X1 U12407 ( .B1(n9974), .B2(n14986), .A(n9973), .ZN(n9975) );
  INV_X1 U12408 ( .A(n9975), .ZN(P2_U3502) );
  INV_X1 U12409 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9978) );
  OR2_X1 U12410 ( .A1(n9976), .A2(n14785), .ZN(n9977) );
  OAI21_X1 U12411 ( .B1(n14748), .B2(n9978), .A(n9977), .ZN(P1_U3468) );
  INV_X1 U12412 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9979) );
  MUX2_X1 U12413 ( .A(n9979), .B(P1_REG1_REG_10__SCAN_IN), .S(n10885), .Z(
        n9982) );
  OAI21_X1 U12414 ( .B1(n10840), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9980), .ZN(
        n9981) );
  NOR2_X1 U12415 ( .A1(n9981), .A2(n9982), .ZN(n10331) );
  AOI211_X1 U12416 ( .C1(n9982), .C2(n9981), .A(n13980), .B(n10331), .ZN(n9995) );
  INV_X1 U12417 ( .A(n10885), .ZN(n9993) );
  INV_X1 U12418 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9983) );
  MUX2_X1 U12419 ( .A(n9983), .B(P1_REG2_REG_10__SCAN_IN), .S(n10885), .Z(
        n9986) );
  NOR2_X1 U12420 ( .A1(n9984), .A2(n10865), .ZN(n9988) );
  INV_X1 U12421 ( .A(n9988), .ZN(n9985) );
  NAND2_X1 U12422 ( .A1(n9986), .A2(n9985), .ZN(n9989) );
  MUX2_X1 U12423 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n9983), .S(n10885), .Z(
        n9987) );
  OAI21_X1 U12424 ( .B1(n9990), .B2(n9988), .A(n9987), .ZN(n10329) );
  OAI211_X1 U12425 ( .C1(n9990), .C2(n9989), .A(n10329), .B(n14027), .ZN(n9992) );
  AND2_X1 U12426 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11531) );
  AOI21_X1 U12427 ( .B1(n13986), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n11531), 
        .ZN(n9991) );
  OAI211_X1 U12428 ( .C1(n14023), .C2(n9993), .A(n9992), .B(n9991), .ZN(n9994)
         );
  OR2_X1 U12429 ( .A1(n9995), .A2(n9994), .ZN(P1_U3253) );
  INV_X1 U12430 ( .A(n13755), .ZN(n11672) );
  AOI22_X1 U12431 ( .A1(n11672), .A2(n6481), .B1(n14984), .B2(
        P2_REG1_REG_1__SCAN_IN), .ZN(n9996) );
  OAI21_X1 U12432 ( .B1(n9997), .B2(n14984), .A(n9996), .ZN(P2_U3500) );
  INV_X1 U12433 ( .A(n9998), .ZN(n9999) );
  NAND2_X1 U12434 ( .A1(n9999), .A2(n10970), .ZN(n10019) );
  NAND2_X1 U12435 ( .A1(n10001), .A2(n10000), .ZN(n10002) );
  NAND2_X1 U12436 ( .A1(n7550), .A2(n10002), .ZN(n10018) );
  INV_X1 U12437 ( .A(n10018), .ZN(n10003) );
  NAND2_X1 U12438 ( .A1(n10019), .A2(n10003), .ZN(n10009) );
  INV_X1 U12439 ( .A(n10009), .ZN(n10004) );
  MUX2_X1 U12440 ( .A(P3_U3897), .B(n10004), .S(n12521), .Z(n12847) );
  INV_X1 U12441 ( .A(n12847), .ZN(n14994) );
  INV_X1 U12442 ( .A(n15002), .ZN(n12811) );
  INV_X1 U12443 ( .A(n10087), .ZN(n10137) );
  NAND2_X1 U12444 ( .A1(n10138), .A2(n10087), .ZN(n10006) );
  OAI21_X1 U12445 ( .B1(n10015), .B2(n10087), .A(n10006), .ZN(n10007) );
  INV_X1 U12446 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15090) );
  NAND2_X1 U12447 ( .A1(n10007), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10140) );
  OAI21_X1 U12448 ( .B1(n10007), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10140), .ZN(
        n10024) );
  INV_X1 U12449 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10314) );
  INV_X1 U12450 ( .A(n10015), .ZN(n10012) );
  NOR2_X1 U12451 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10010), .ZN(n10086) );
  NAND2_X1 U12452 ( .A1(n10148), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10011) );
  NOR2_X1 U12453 ( .A1(n10013), .A2(n10314), .ZN(n10150) );
  AOI21_X1 U12454 ( .B1(n10314), .B2(n10013), .A(n10150), .ZN(n10014) );
  NOR2_X1 U12455 ( .A1(n15008), .A2(n10014), .ZN(n10023) );
  MUX2_X1 U12456 ( .A(n10010), .B(n10005), .S(n13141), .Z(n10091) );
  NAND2_X1 U12457 ( .A1(n10091), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10085) );
  OAI21_X1 U12458 ( .B1(n10016), .B2(n10015), .A(n10161), .ZN(n10017) );
  AOI21_X1 U12459 ( .B1(n10085), .B2(n10017), .A(n10211), .ZN(n10021) );
  NAND2_X1 U12460 ( .A1(P3_U3897), .A2(n12521), .ZN(n15000) );
  AOI22_X1 U12461 ( .A1(n14987), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10020) );
  OAI21_X1 U12462 ( .B1(n10021), .B2(n15000), .A(n10020), .ZN(n10022) );
  AOI211_X1 U12463 ( .C1(n12811), .C2(n10024), .A(n10023), .B(n10022), .ZN(
        n10025) );
  OAI21_X1 U12464 ( .B1(n10012), .B2(n14994), .A(n10025), .ZN(P3_U3183) );
  INV_X1 U12465 ( .A(n10306), .ZN(n10039) );
  XNOR2_X1 U12466 ( .A(n10523), .B(n10031), .ZN(n10030) );
  NAND2_X1 U12467 ( .A1(n10030), .A2(n10029), .ZN(n10068) );
  NAND3_X1 U12468 ( .A1(n10310), .A2(n10532), .A3(n10032), .ZN(n10033) );
  NOR3_X1 U12469 ( .A1(n10307), .A2(n10532), .A3(n10303), .ZN(n10037) );
  NAND2_X1 U12470 ( .A1(n10532), .A2(n10306), .ZN(n10035) );
  NAND2_X1 U12471 ( .A1(n10035), .A2(n10034), .ZN(n10036) );
  AOI211_X1 U12472 ( .C1(n10039), .C2(n10038), .A(n10037), .B(n10070), .ZN(
        n10045) );
  INV_X1 U12473 ( .A(n12722), .ZN(n10309) );
  NAND2_X1 U12474 ( .A1(n10041), .A2(n10040), .ZN(n12652) );
  AOI22_X1 U12475 ( .A1(n12649), .A2(n12721), .B1(n10310), .B2(n12674), .ZN(
        n10042) );
  OAI21_X1 U12476 ( .B1(n10309), .B2(n12652), .A(n10042), .ZN(n10043) );
  AOI21_X1 U12477 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n10075), .A(n10043), .ZN(
        n10044) );
  OAI21_X1 U12478 ( .B1(n10045), .B2(n12689), .A(n10044), .ZN(P3_U3162) );
  INV_X1 U12479 ( .A(n14924), .ZN(n10050) );
  INV_X1 U12480 ( .A(n10046), .ZN(n10049) );
  NAND4_X1 U12481 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        n10051) );
  NAND2_X1 U12482 ( .A1(n10060), .A2(n10052), .ZN(n14926) );
  AND2_X1 U12483 ( .A1(n9792), .A2(n13603), .ZN(n10053) );
  OR2_X1 U12484 ( .A1(n14928), .A2(n10053), .ZN(n10055) );
  NAND2_X1 U12485 ( .A1(n13359), .A2(n13466), .ZN(n10054) );
  AND2_X1 U12486 ( .A1(n10055), .A2(n10054), .ZN(n14927) );
  INV_X1 U12487 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10056) );
  OAI22_X1 U12488 ( .A1(n13595), .A2(n14927), .B1(n10056), .B2(n13639), .ZN(
        n10057) );
  AOI21_X1 U12489 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n13595), .A(n10057), .ZN(
        n10064) );
  NAND2_X1 U12490 ( .A1(n13642), .A2(n10058), .ZN(n13591) );
  INV_X1 U12491 ( .A(n13591), .ZN(n10062) );
  INV_X1 U12492 ( .A(n14928), .ZN(n10061) );
  AOI22_X1 U12493 ( .A1(n10062), .A2(n10061), .B1(n13655), .B2(n10060), .ZN(
        n10063) );
  OAI211_X1 U12494 ( .C1(n13659), .C2(n14926), .A(n10064), .B(n10063), .ZN(
        P2_U3265) );
  AOI22_X1 U12495 ( .A1(n11672), .A2(n10065), .B1(n14984), .B2(
        P2_REG1_REG_2__SCAN_IN), .ZN(n10066) );
  OAI21_X1 U12496 ( .B1(n10067), .B2(n14984), .A(n10066), .ZN(P2_U3501) );
  INV_X1 U12497 ( .A(n10068), .ZN(n10069) );
  XNOR2_X1 U12498 ( .A(n10523), .B(n10106), .ZN(n10524) );
  XNOR2_X1 U12499 ( .A(n10524), .B(n10560), .ZN(n10071) );
  AOI21_X1 U12500 ( .B1(n10072), .B2(n10071), .A(n10529), .ZN(n10077) );
  AOI22_X1 U12501 ( .A1(n12649), .A2(n12720), .B1(n10106), .B2(n6477), .ZN(
        n10073) );
  OAI21_X1 U12502 ( .B1(n10029), .B2(n12652), .A(n10073), .ZN(n10074) );
  AOI21_X1 U12503 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10075), .A(n10074), .ZN(
        n10076) );
  OAI21_X1 U12504 ( .B1(n10077), .B2(n12689), .A(n10076), .ZN(P3_U3177) );
  INV_X1 U12505 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10078) );
  OR2_X1 U12506 ( .A1(n14748), .A2(n10078), .ZN(n10079) );
  OAI21_X1 U12507 ( .B1(n10080), .B2(n14785), .A(n10079), .ZN(P1_U3471) );
  INV_X1 U12508 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10082) );
  MUX2_X1 U12509 ( .A(n10082), .B(n10081), .S(n15089), .Z(n10083) );
  OAI21_X1 U12510 ( .B1(n10084), .B2(n13129), .A(n10083), .ZN(P3_U3390) );
  INV_X1 U12511 ( .A(n10085), .ZN(n10096) );
  NAND3_X1 U12512 ( .A1(n15008), .A2(n15002), .A3(n15000), .ZN(n10095) );
  INV_X1 U12513 ( .A(n10086), .ZN(n10090) );
  NAND2_X1 U12514 ( .A1(n12811), .A2(n10087), .ZN(n10089) );
  AOI22_X1 U12515 ( .A1(n14987), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10088) );
  OAI211_X1 U12516 ( .C1(n10090), .C2(n15008), .A(n10089), .B(n10088), .ZN(
        n10094) );
  NOR2_X1 U12517 ( .A1(n15000), .A2(n10091), .ZN(n10092) );
  MUX2_X1 U12518 ( .A(n10092), .B(n12847), .S(P3_IR_REG_0__SCAN_IN), .Z(n10093) );
  AOI211_X1 U12519 ( .C1(n10096), .C2(n10095), .A(n10094), .B(n10093), .ZN(
        n10097) );
  INV_X1 U12520 ( .A(n10097), .ZN(P3_U3182) );
  INV_X1 U12521 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n10162) );
  XNOR2_X1 U12522 ( .A(n10099), .B(n10098), .ZN(n15021) );
  INV_X1 U12523 ( .A(n15085), .ZN(n15061) );
  OR2_X1 U12524 ( .A1(n15021), .A2(n15061), .ZN(n10105) );
  XNOR2_X1 U12525 ( .A(n10100), .B(n10099), .ZN(n10101) );
  NAND2_X1 U12526 ( .A1(n10101), .A2(n13019), .ZN(n10104) );
  OAI22_X1 U12527 ( .A1(n10029), .A2(n12964), .B1(n10538), .B2(n12962), .ZN(
        n10102) );
  INV_X1 U12528 ( .A(n10102), .ZN(n10103) );
  NAND3_X1 U12529 ( .A1(n10105), .A2(n10104), .A3(n10103), .ZN(n15026) );
  INV_X1 U12530 ( .A(n15041), .ZN(n15081) );
  NAND2_X1 U12531 ( .A1(n10106), .A2(n15065), .ZN(n15022) );
  OAI21_X1 U12532 ( .B1(n15021), .B2(n15081), .A(n15022), .ZN(n10107) );
  NOR2_X1 U12533 ( .A1(n15026), .A2(n10107), .ZN(n15040) );
  MUX2_X1 U12534 ( .A(n10162), .B(n15040), .S(n15106), .Z(n10108) );
  INV_X1 U12535 ( .A(n10108), .ZN(P3_U3461) );
  OAI22_X1 U12536 ( .A1(n13321), .A2(n10110), .B1(n10109), .B2(n13282), .ZN(
        n10117) );
  INV_X1 U12537 ( .A(n13329), .ZN(n13306) );
  AOI22_X1 U12538 ( .A1(n13306), .A2(n10112), .B1(n10111), .B2(n13276), .ZN(
        n10115) );
  INV_X1 U12539 ( .A(n10113), .ZN(n10114) );
  NOR2_X1 U12540 ( .A1(n10115), .A2(n10114), .ZN(n10116) );
  AOI211_X1 U12541 ( .C1(P2_REG3_REG_1__SCAN_IN), .C2(n10118), .A(n10117), .B(
        n10116), .ZN(n10119) );
  OAI21_X1 U12542 ( .B1(n9814), .B2(n14808), .A(n10119), .ZN(P2_U3194) );
  INV_X1 U12543 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10121) );
  MUX2_X1 U12544 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10121), .S(n10664), .Z(
        n10122) );
  OAI21_X1 U12545 ( .B1(n10123), .B2(n10122), .A(n10660), .ZN(n10124) );
  NAND2_X1 U12546 ( .A1(n10124), .A2(n14876), .ZN(n10133) );
  MUX2_X1 U12547 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10960), .S(n10664), .Z(
        n10128) );
  AOI21_X1 U12548 ( .B1(n10126), .B2(P2_REG2_REG_8__SCAN_IN), .A(n10125), .ZN(
        n10127) );
  NAND2_X1 U12549 ( .A1(n10127), .A2(n10128), .ZN(n10663) );
  OAI21_X1 U12550 ( .B1(n10128), .B2(n10127), .A(n10663), .ZN(n10129) );
  INV_X1 U12551 ( .A(n10129), .ZN(n10130) );
  OAI22_X1 U12552 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11038), .B1(n10130), .B2(
        n14852), .ZN(n10131) );
  AOI21_X1 U12553 ( .B1(n14821), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n10131), .ZN(
        n10132) );
  OAI211_X1 U12554 ( .C1(n14839), .C2(n10134), .A(n10133), .B(n10132), .ZN(
        P2_U3223) );
  OAI222_X1 U12555 ( .A1(n6484), .A2(n10136), .B1(n13143), .B2(n10135), .C1(
        P3_U3151), .C2(n12833), .ZN(P3_U3276) );
  INV_X1 U12556 ( .A(n10219), .ZN(n10171) );
  XNOR2_X1 U12557 ( .A(n7529), .B(n10162), .ZN(n10199) );
  OR2_X1 U12558 ( .A1(n10138), .A2(n10137), .ZN(n10139) );
  NAND2_X1 U12559 ( .A1(n10140), .A2(n10139), .ZN(n10198) );
  NAND2_X1 U12560 ( .A1(n10199), .A2(n10198), .ZN(n10197) );
  NAND2_X1 U12561 ( .A1(n10216), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10141) );
  NAND2_X1 U12562 ( .A1(n10197), .A2(n10141), .ZN(n10142) );
  INV_X1 U12563 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15092) );
  INV_X1 U12564 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15094) );
  XNOR2_X1 U12565 ( .A(n10219), .B(n15094), .ZN(n10144) );
  NAND2_X1 U12566 ( .A1(n10143), .A2(n10144), .ZN(n10221) );
  INV_X1 U12567 ( .A(n10144), .ZN(n10146) );
  NAND3_X1 U12568 ( .A1(n10184), .A2(n10146), .A3(n10145), .ZN(n10147) );
  AND2_X1 U12569 ( .A1(n10221), .A2(n10147), .ZN(n10159) );
  XNOR2_X1 U12570 ( .A(n10216), .B(P3_REG2_REG_2__SCAN_IN), .ZN(n10202) );
  NOR2_X1 U12571 ( .A1(n10151), .A2(n6653), .ZN(n10152) );
  INV_X1 U12572 ( .A(n10152), .ZN(n10153) );
  XNOR2_X1 U12573 ( .A(n10219), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n10154) );
  AND3_X1 U12574 ( .A1(n10181), .A2(n10154), .A3(n10153), .ZN(n10155) );
  INV_X1 U12575 ( .A(n15008), .ZN(n12820) );
  OAI21_X1 U12576 ( .B1(n10217), .B2(n10155), .A(n12820), .ZN(n10158) );
  NOR2_X1 U12577 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10156), .ZN(n10540) );
  AOI21_X1 U12578 ( .B1(n14987), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10540), .ZN(
        n10157) );
  OAI211_X1 U12579 ( .C1(n10159), .C2(n15002), .A(n10158), .B(n10157), .ZN(
        n10160) );
  AOI21_X1 U12580 ( .B1(n10171), .B2(n12847), .A(n10160), .ZN(n10180) );
  INV_X1 U12581 ( .A(n10161), .ZN(n10210) );
  INV_X1 U12582 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10163) );
  MUX2_X1 U12583 ( .A(n10163), .B(n10162), .S(n13141), .Z(n10164) );
  NAND2_X1 U12584 ( .A1(n10164), .A2(n7530), .ZN(n10191) );
  INV_X1 U12585 ( .A(n10164), .ZN(n10165) );
  NAND2_X1 U12586 ( .A1(n10165), .A2(n10216), .ZN(n10166) );
  AND2_X1 U12587 ( .A1(n10191), .A2(n10166), .ZN(n10209) );
  OAI21_X1 U12588 ( .B1(n10211), .B2(n10210), .A(n10209), .ZN(n10208) );
  INV_X1 U12589 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10322) );
  MUX2_X1 U12590 ( .A(n10322), .B(n15092), .S(n13141), .Z(n10167) );
  NAND2_X1 U12591 ( .A1(n10167), .A2(n6653), .ZN(n10170) );
  INV_X1 U12592 ( .A(n10167), .ZN(n10168) );
  NAND2_X1 U12593 ( .A1(n10168), .A2(n10196), .ZN(n10169) );
  NAND2_X1 U12594 ( .A1(n10170), .A2(n10169), .ZN(n10190) );
  INV_X1 U12595 ( .A(n10170), .ZN(n10176) );
  INV_X1 U12596 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10461) );
  MUX2_X1 U12597 ( .A(n10461), .B(n15094), .S(n13141), .Z(n10172) );
  NAND2_X1 U12598 ( .A1(n10172), .A2(n10171), .ZN(n10235) );
  INV_X1 U12599 ( .A(n10172), .ZN(n10173) );
  NAND2_X1 U12600 ( .A1(n10173), .A2(n10219), .ZN(n10174) );
  AND2_X1 U12601 ( .A1(n10235), .A2(n10174), .ZN(n10175) );
  OAI21_X1 U12602 ( .B1(n10193), .B2(n10176), .A(n10175), .ZN(n10236) );
  INV_X1 U12603 ( .A(n10236), .ZN(n10178) );
  NOR3_X1 U12604 ( .A1(n10193), .A2(n10176), .A3(n10175), .ZN(n10177) );
  INV_X1 U12605 ( .A(n15000), .ZN(n12778) );
  OAI21_X1 U12606 ( .B1(n10178), .B2(n10177), .A(n12778), .ZN(n10179) );
  NAND2_X1 U12607 ( .A1(n10180), .A2(n10179), .ZN(P3_U3186) );
  OAI21_X1 U12608 ( .B1(n10182), .B2(P3_REG2_REG_3__SCAN_IN), .A(n10181), .ZN(
        n10183) );
  NAND2_X1 U12609 ( .A1(n12820), .A2(n10183), .ZN(n10189) );
  NOR2_X1 U12610 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10569), .ZN(n10558) );
  AOI21_X1 U12611 ( .B1(n14987), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10558), .ZN(
        n10188) );
  OAI21_X1 U12612 ( .B1(n10185), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10184), .ZN(
        n10186) );
  NAND2_X1 U12613 ( .A1(n12811), .A2(n10186), .ZN(n10187) );
  AND3_X1 U12614 ( .A1(n10189), .A2(n10188), .A3(n10187), .ZN(n10195) );
  AND3_X1 U12615 ( .A1(n10208), .A2(n10191), .A3(n10190), .ZN(n10192) );
  OAI21_X1 U12616 ( .B1(n10193), .B2(n10192), .A(n12778), .ZN(n10194) );
  OAI211_X1 U12617 ( .C1(n14994), .C2(n10196), .A(n10195), .B(n10194), .ZN(
        P3_U3185) );
  OAI21_X1 U12618 ( .B1(n10199), .B2(n10198), .A(n10197), .ZN(n10207) );
  AOI21_X1 U12619 ( .B1(n10202), .B2(n10201), .A(n10200), .ZN(n10203) );
  NOR2_X1 U12620 ( .A1(n15008), .A2(n10203), .ZN(n10206) );
  INV_X1 U12621 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10204) );
  INV_X1 U12622 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15024) );
  OAI22_X1 U12623 ( .A1(n14991), .A2(n10204), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15024), .ZN(n10205) );
  AOI211_X1 U12624 ( .C1(n12811), .C2(n10207), .A(n10206), .B(n10205), .ZN(
        n10215) );
  INV_X1 U12625 ( .A(n10208), .ZN(n10213) );
  NOR3_X1 U12626 ( .A1(n10211), .A2(n10210), .A3(n10209), .ZN(n10212) );
  OAI21_X1 U12627 ( .B1(n10213), .B2(n10212), .A(n12778), .ZN(n10214) );
  OAI211_X1 U12628 ( .C1(n14994), .C2(n10216), .A(n10215), .B(n10214), .ZN(
        P3_U3184) );
  OAI21_X1 U12629 ( .B1(n10218), .B2(P3_REG2_REG_5__SCAN_IN), .A(n12725), .ZN(
        n10230) );
  NAND2_X1 U12630 ( .A1(n10219), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10220) );
  NAND2_X1 U12631 ( .A1(n10221), .A2(n10220), .ZN(n10222) );
  INV_X1 U12632 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15096) );
  AND2_X1 U12633 ( .A1(n10223), .A2(n15096), .ZN(n10224) );
  NOR2_X1 U12634 ( .A1(n12739), .A2(n10224), .ZN(n10228) );
  NOR2_X1 U12635 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10225), .ZN(n10755) );
  INV_X1 U12636 ( .A(n10755), .ZN(n10227) );
  NAND2_X1 U12637 ( .A1(n14987), .A2(P3_ADDR_REG_5__SCAN_IN), .ZN(n10226) );
  OAI211_X1 U12638 ( .C1(n15002), .C2(n10228), .A(n10227), .B(n10226), .ZN(
        n10229) );
  AOI21_X1 U12639 ( .B1(n10230), .B2(n12820), .A(n10229), .ZN(n10239) );
  INV_X1 U12640 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10826) );
  MUX2_X1 U12641 ( .A(n10826), .B(n15096), .S(n13141), .Z(n10231) );
  NAND2_X1 U12642 ( .A1(n10231), .A2(n6920), .ZN(n10249) );
  INV_X1 U12643 ( .A(n10231), .ZN(n10232) );
  NAND2_X1 U12644 ( .A1(n10232), .A2(n10240), .ZN(n10233) );
  NAND2_X1 U12645 ( .A1(n10249), .A2(n10233), .ZN(n10234) );
  AOI21_X1 U12646 ( .B1(n10236), .B2(n10235), .A(n10234), .ZN(n12733) );
  AND3_X1 U12647 ( .A1(n10236), .A2(n10235), .A3(n10234), .ZN(n10237) );
  OAI21_X1 U12648 ( .B1(n12733), .B2(n10237), .A(n12778), .ZN(n10238) );
  OAI211_X1 U12649 ( .C1(n14994), .C2(n10240), .A(n10239), .B(n10238), .ZN(
        P3_U3187) );
  INV_X1 U12650 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15100) );
  INV_X1 U12651 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15098) );
  XNOR2_X1 U12652 ( .A(n12736), .B(P3_REG1_REG_6__SCAN_IN), .ZN(n12738) );
  OAI21_X1 U12653 ( .B1(n12736), .B2(n15098), .A(n12737), .ZN(n10274) );
  XNOR2_X1 U12654 ( .A(n10274), .B(n10281), .ZN(n10241) );
  AOI21_X1 U12655 ( .B1(n15100), .B2(n10241), .A(n10273), .ZN(n10263) );
  INV_X1 U12656 ( .A(n10281), .ZN(n10254) );
  INV_X1 U12657 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10244) );
  NOR2_X1 U12658 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10242), .ZN(n11072) );
  INV_X1 U12659 ( .A(n11072), .ZN(n10243) );
  OAI21_X1 U12660 ( .B1(n14991), .B2(n10244), .A(n10243), .ZN(n10248) );
  INV_X1 U12661 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11138) );
  INV_X1 U12662 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11151) );
  XNOR2_X1 U12663 ( .A(n12736), .B(n11151), .ZN(n12724) );
  AOI21_X1 U12664 ( .B1(n11138), .B2(n10245), .A(n10284), .ZN(n10246) );
  NOR2_X1 U12665 ( .A1(n10246), .A2(n15008), .ZN(n10247) );
  AOI211_X1 U12666 ( .C1(n12847), .C2(n10254), .A(n10248), .B(n10247), .ZN(
        n10262) );
  INV_X1 U12667 ( .A(n10249), .ZN(n12732) );
  MUX2_X1 U12668 ( .A(n11151), .B(n15098), .S(n13141), .Z(n10250) );
  NAND2_X1 U12669 ( .A1(n10250), .A2(n12736), .ZN(n10259) );
  INV_X1 U12670 ( .A(n10250), .ZN(n10252) );
  NAND2_X1 U12671 ( .A1(n10252), .A2(n10251), .ZN(n10253) );
  AND2_X1 U12672 ( .A1(n10259), .A2(n10253), .ZN(n12731) );
  OAI21_X1 U12673 ( .B1(n12733), .B2(n12732), .A(n12731), .ZN(n12730) );
  MUX2_X1 U12674 ( .A(n11138), .B(n15100), .S(n13141), .Z(n10255) );
  NAND2_X1 U12675 ( .A1(n10255), .A2(n10254), .ZN(n10290) );
  INV_X1 U12676 ( .A(n10255), .ZN(n10256) );
  NAND2_X1 U12677 ( .A1(n10256), .A2(n10281), .ZN(n10257) );
  NAND2_X1 U12678 ( .A1(n10290), .A2(n10257), .ZN(n10258) );
  AND3_X1 U12679 ( .A1(n12730), .A2(n10259), .A3(n10258), .ZN(n10260) );
  OAI21_X1 U12680 ( .B1(n10297), .B2(n10260), .A(n12778), .ZN(n10261) );
  OAI211_X1 U12681 ( .C1(n10263), .C2(n15002), .A(n10262), .B(n10261), .ZN(
        P3_U3189) );
  INV_X1 U12682 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10264) );
  NAND3_X1 U12683 ( .A1(n10266), .A2(n10265), .A3(n10264), .ZN(n10267) );
  OAI21_X1 U12684 ( .B1(n10268), .B2(n10267), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10269) );
  XNOR2_X1 U12685 ( .A(n10269), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14682) );
  INV_X1 U12686 ( .A(n14682), .ZN(n11738) );
  INV_X1 U12687 ( .A(n11628), .ZN(n10271) );
  OAI222_X1 U12688 ( .A1(P1_U3086), .A2(n11738), .B1(n14391), .B2(n10271), 
        .C1(n10270), .C2(n14396), .ZN(P1_U3340) );
  INV_X1 U12689 ( .A(n13364), .ZN(n13375) );
  OAI222_X1 U12690 ( .A1(n13819), .A2(n10272), .B1(n13817), .B2(n10271), .C1(
        n13375), .C2(P2_U3088), .ZN(P2_U3312) );
  NAND2_X1 U12691 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n10407), .ZN(n10275) );
  OAI21_X1 U12692 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n10407), .A(n10275), .ZN(
        n10276) );
  AOI21_X1 U12693 ( .B1(n10277), .B2(n10276), .A(n10406), .ZN(n10302) );
  INV_X1 U12694 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n10279) );
  AND2_X1 U12695 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n11269) );
  INV_X1 U12696 ( .A(n11269), .ZN(n10278) );
  OAI21_X1 U12697 ( .B1(n14991), .B2(n10279), .A(n10278), .ZN(n10289) );
  INV_X1 U12698 ( .A(n10280), .ZN(n10282) );
  NAND2_X1 U12699 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n10407), .ZN(n10285) );
  OAI21_X1 U12700 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n10407), .A(n10285), .ZN(
        n10286) );
  AOI21_X1 U12701 ( .B1(n6610), .B2(n10286), .A(n10394), .ZN(n10287) );
  NOR2_X1 U12702 ( .A1(n10287), .A2(n15008), .ZN(n10288) );
  AOI211_X1 U12703 ( .C1(n12847), .C2(n10291), .A(n10289), .B(n10288), .ZN(
        n10301) );
  INV_X1 U12704 ( .A(n10290), .ZN(n10296) );
  INV_X1 U12705 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11461) );
  INV_X1 U12706 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15102) );
  MUX2_X1 U12707 ( .A(n11461), .B(n15102), .S(n13141), .Z(n10292) );
  NAND2_X1 U12708 ( .A1(n10292), .A2(n10291), .ZN(n10403) );
  INV_X1 U12709 ( .A(n10292), .ZN(n10293) );
  NAND2_X1 U12710 ( .A1(n10293), .A2(n10407), .ZN(n10294) );
  AND2_X1 U12711 ( .A1(n10403), .A2(n10294), .ZN(n10295) );
  OAI21_X1 U12712 ( .B1(n10297), .B2(n10296), .A(n10295), .ZN(n10404) );
  INV_X1 U12713 ( .A(n10404), .ZN(n10299) );
  NOR3_X1 U12714 ( .A1(n10297), .A2(n10296), .A3(n10295), .ZN(n10298) );
  OAI21_X1 U12715 ( .B1(n10299), .B2(n10298), .A(n12778), .ZN(n10300) );
  OAI211_X1 U12716 ( .C1(n10302), .C2(n15002), .A(n10301), .B(n10300), .ZN(
        P3_U3190) );
  XNOR2_X1 U12717 ( .A(n10304), .B(n10303), .ZN(n15035) );
  AND2_X1 U12718 ( .A1(n15023), .A2(n10305), .ZN(n15029) );
  OR2_X1 U12719 ( .A1(n15085), .A2(n15029), .ZN(n15010) );
  XNOR2_X1 U12720 ( .A(n10307), .B(n10306), .ZN(n10308) );
  OAI222_X1 U12721 ( .A1(n12964), .A2(n10309), .B1(n12962), .B2(n10560), .C1(
        n12960), .C2(n10308), .ZN(n15037) );
  INV_X1 U12722 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10311) );
  NAND2_X1 U12723 ( .A1(n10310), .A2(n15065), .ZN(n15033) );
  OAI22_X1 U12724 ( .A1(n15025), .A2(n10311), .B1(n15023), .B2(n15033), .ZN(
        n10312) );
  NOR2_X1 U12725 ( .A1(n15037), .A2(n10312), .ZN(n10313) );
  MUX2_X1 U12726 ( .A(n10314), .B(n10313), .S(n15030), .Z(n10315) );
  OAI21_X1 U12727 ( .B1(n15035), .B2(n11466), .A(n10315), .ZN(P3_U3232) );
  XNOR2_X1 U12728 ( .A(n10316), .B(n10317), .ZN(n15046) );
  INV_X1 U12729 ( .A(n15046), .ZN(n10325) );
  AOI21_X1 U12730 ( .B1(n10318), .B2(n10317), .A(n12960), .ZN(n10321) );
  OAI22_X1 U12731 ( .A1(n10560), .A2(n12964), .B1(n10753), .B2(n12962), .ZN(
        n10319) );
  AOI21_X1 U12732 ( .B1(n10321), .B2(n10320), .A(n10319), .ZN(n15043) );
  MUX2_X1 U12733 ( .A(n10322), .B(n15043), .S(n15030), .Z(n10324) );
  AOI22_X1 U12734 ( .A1(n15016), .A2(n10559), .B1(n15014), .B2(n10569), .ZN(
        n10323) );
  OAI211_X1 U12735 ( .C1(n11466), .C2(n10325), .A(n10324), .B(n10323), .ZN(
        P3_U3230) );
  NAND2_X1 U12736 ( .A1(n10885), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10328) );
  INV_X1 U12737 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10326) );
  MUX2_X1 U12738 ( .A(n10326), .B(P1_REG2_REG_11__SCAN_IN), .S(n10977), .Z(
        n10327) );
  AOI21_X1 U12739 ( .B1(n10329), .B2(n10328), .A(n10327), .ZN(n10549) );
  NAND3_X1 U12740 ( .A1(n10329), .A2(n10328), .A3(n10327), .ZN(n10330) );
  NAND2_X1 U12741 ( .A1(n10330), .A2(n14027), .ZN(n10341) );
  INV_X1 U12742 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10332) );
  MUX2_X1 U12743 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10332), .S(n10977), .Z(
        n10333) );
  OAI21_X1 U12744 ( .B1(n10334), .B2(n10333), .A(n10545), .ZN(n10335) );
  NAND2_X1 U12745 ( .A1(n10335), .A2(n14680), .ZN(n10340) );
  NAND2_X1 U12746 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11724)
         );
  INV_X1 U12747 ( .A(n11724), .ZN(n10338) );
  NOR2_X1 U12748 ( .A1(n14023), .A2(n10336), .ZN(n10337) );
  AOI211_X1 U12749 ( .C1(n13986), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n10338), 
        .B(n10337), .ZN(n10339) );
  OAI211_X1 U12750 ( .C1(n10549), .C2(n10341), .A(n10340), .B(n10339), .ZN(
        P1_U3254) );
  INV_X1 U12751 ( .A(n11802), .ZN(n10452) );
  OAI21_X1 U12752 ( .B1(n10342), .B2(n6597), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10343) );
  XNOR2_X1 U12753 ( .A(n10343), .B(P1_IR_REG_16__SCAN_IN), .ZN(n13989) );
  AOI22_X1 U12754 ( .A1(n13989), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n14389), .ZN(n10344) );
  OAI21_X1 U12755 ( .B1(n10452), .B2(n14391), .A(n10344), .ZN(P1_U3339) );
  INV_X1 U12756 ( .A(n9792), .ZN(n14946) );
  NAND2_X1 U12757 ( .A1(n13642), .A2(n14946), .ZN(n10345) );
  INV_X1 U12758 ( .A(n10346), .ZN(n10354) );
  INV_X1 U12759 ( .A(n10347), .ZN(n10348) );
  MUX2_X1 U12760 ( .A(n10349), .B(n10348), .S(n13642), .Z(n10353) );
  OAI22_X1 U12761 ( .A1(n13589), .A2(n10355), .B1(n10432), .B2(n13639), .ZN(
        n10350) );
  AOI21_X1 U12762 ( .B1(n13646), .B2(n10351), .A(n10350), .ZN(n10352) );
  OAI211_X1 U12763 ( .C1(n13636), .C2(n10354), .A(n10353), .B(n10352), .ZN(
        P2_U3261) );
  NAND2_X1 U12764 ( .A1(n10355), .A2(n10361), .ZN(n10356) );
  XNOR2_X1 U12765 ( .A(n10376), .B(n10364), .ZN(n14934) );
  INV_X1 U12766 ( .A(n10358), .ZN(n10359) );
  NAND2_X1 U12767 ( .A1(n10360), .A2(n10359), .ZN(n10363) );
  NAND2_X1 U12768 ( .A1(n10361), .A2(n10433), .ZN(n10362) );
  XOR2_X1 U12769 ( .A(n10381), .B(n10364), .Z(n10367) );
  NAND2_X1 U12770 ( .A1(n13356), .A2(n13628), .ZN(n10366) );
  NAND2_X1 U12771 ( .A1(n13354), .A2(n13466), .ZN(n10365) );
  AND2_X1 U12772 ( .A1(n10366), .A2(n10365), .ZN(n10576) );
  OAI21_X1 U12773 ( .B1(n10367), .B2(n13603), .A(n10576), .ZN(n14930) );
  INV_X1 U12774 ( .A(n14930), .ZN(n10368) );
  MUX2_X1 U12775 ( .A(n10369), .B(n10368), .S(n13642), .Z(n10374) );
  OR2_X1 U12776 ( .A1(n10371), .A2(n14932), .ZN(n10377) );
  INV_X1 U12777 ( .A(n10377), .ZN(n10370) );
  AOI211_X1 U12778 ( .C1(n14932), .C2(n10371), .A(n13221), .B(n10370), .ZN(
        n14931) );
  INV_X1 U12779 ( .A(n14932), .ZN(n10375) );
  OAI22_X1 U12780 ( .A1(n13589), .A2(n10375), .B1(n13639), .B2(n10579), .ZN(
        n10372) );
  AOI21_X1 U12781 ( .B1(n14931), .B2(n13646), .A(n10372), .ZN(n10373) );
  OAI211_X1 U12782 ( .C1(n13636), .C2(n14934), .A(n10374), .B(n10373), .ZN(
        P2_U3260) );
  INV_X1 U12783 ( .A(n13355), .ZN(n10382) );
  XOR2_X1 U12784 ( .A(n10727), .B(n10726), .Z(n14943) );
  AOI211_X1 U12785 ( .C1(n14938), .C2(n10377), .A(n13221), .B(n10779), .ZN(
        n14937) );
  INV_X1 U12786 ( .A(n14938), .ZN(n10378) );
  OAI22_X1 U12787 ( .A1(n13589), .A2(n10378), .B1(n10719), .B2(n13639), .ZN(
        n10379) );
  AOI21_X1 U12788 ( .B1(n14937), .B2(n13646), .A(n10379), .ZN(n10392) );
  AND2_X1 U12789 ( .A1(n14932), .A2(n10382), .ZN(n10380) );
  OR2_X1 U12790 ( .A1(n10382), .A2(n14932), .ZN(n10383) );
  NAND2_X1 U12791 ( .A1(n10384), .A2(n10726), .ZN(n10385) );
  NAND2_X1 U12792 ( .A1(n10735), .A2(n10385), .ZN(n10389) );
  NAND2_X1 U12793 ( .A1(n13355), .A2(n13628), .ZN(n10387) );
  NAND2_X1 U12794 ( .A1(n13353), .A2(n13466), .ZN(n10386) );
  AND2_X1 U12795 ( .A1(n10387), .A2(n10386), .ZN(n10721) );
  INV_X1 U12796 ( .A(n10721), .ZN(n10388) );
  AOI21_X1 U12797 ( .B1(n10389), .B2(n13625), .A(n10388), .ZN(n14941) );
  MUX2_X1 U12798 ( .A(n10390), .B(n14941), .S(n13642), .Z(n10391) );
  OAI211_X1 U12799 ( .C1(n14943), .C2(n13636), .A(n10392), .B(n10391), .ZN(
        P2_U3259) );
  INV_X1 U12800 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10396) );
  AOI21_X1 U12801 ( .B1(n10396), .B2(n10395), .A(n10683), .ZN(n10416) );
  INV_X1 U12802 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10397) );
  MUX2_X1 U12803 ( .A(n10396), .B(n10397), .S(n13141), .Z(n10398) );
  NAND2_X1 U12804 ( .A1(n10398), .A2(n10697), .ZN(n10686) );
  INV_X1 U12805 ( .A(n10398), .ZN(n10400) );
  NAND2_X1 U12806 ( .A1(n10400), .A2(n10399), .ZN(n10401) );
  NAND2_X1 U12807 ( .A1(n10686), .A2(n10401), .ZN(n10402) );
  AOI21_X1 U12808 ( .B1(n10404), .B2(n10403), .A(n10402), .ZN(n10693) );
  AND3_X1 U12809 ( .A1(n10404), .A2(n10403), .A3(n10402), .ZN(n10405) );
  OAI21_X1 U12810 ( .B1(n10693), .B2(n10405), .A(n12778), .ZN(n10415) );
  XNOR2_X1 U12811 ( .A(n10696), .B(n10697), .ZN(n10408) );
  NOR2_X1 U12812 ( .A1(n10397), .A2(n10408), .ZN(n10698) );
  AOI21_X1 U12813 ( .B1(n10397), .B2(n10408), .A(n10698), .ZN(n10412) );
  NOR2_X1 U12814 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10409), .ZN(n11063) );
  AOI21_X1 U12815 ( .B1(n14987), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11063), .ZN(
        n10411) );
  NAND2_X1 U12816 ( .A1(n12847), .A2(n10697), .ZN(n10410) );
  OAI211_X1 U12817 ( .C1(n10412), .C2(n15002), .A(n10411), .B(n10410), .ZN(
        n10413) );
  INV_X1 U12818 ( .A(n10413), .ZN(n10414) );
  OAI211_X1 U12819 ( .C1(n10416), .C2(n15008), .A(n10415), .B(n10414), .ZN(
        P3_U3191) );
  INV_X1 U12820 ( .A(n10417), .ZN(n10419) );
  NAND2_X1 U12821 ( .A1(n10419), .A2(n10418), .ZN(n10420) );
  XNOR2_X1 U12822 ( .A(n13222), .B(n9108), .ZN(n10422) );
  AND2_X1 U12823 ( .A1(n13357), .A2(n9793), .ZN(n10423) );
  NAND2_X1 U12824 ( .A1(n10422), .A2(n10423), .ZN(n10428) );
  INV_X1 U12825 ( .A(n10422), .ZN(n10426) );
  INV_X1 U12826 ( .A(n10423), .ZN(n10424) );
  NAND2_X1 U12827 ( .A1(n10426), .A2(n10424), .ZN(n10425) );
  NAND2_X1 U12828 ( .A1(n10428), .A2(n10425), .ZN(n10504) );
  INV_X1 U12829 ( .A(n10430), .ZN(n10503) );
  NOR3_X1 U12830 ( .A1(n13329), .A2(n10426), .A3(n7226), .ZN(n10427) );
  AOI21_X1 U12831 ( .B1(n10503), .B2(n13276), .A(n10427), .ZN(n10442) );
  XNOR2_X1 U12832 ( .A(n9794), .B(n10433), .ZN(n10580) );
  NAND2_X1 U12833 ( .A1(n13356), .A2(n9793), .ZN(n10574) );
  XNOR2_X1 U12834 ( .A(n10580), .B(n10574), .ZN(n10441) );
  AND2_X1 U12835 ( .A1(n10441), .A2(n10428), .ZN(n10429) );
  NOR2_X1 U12836 ( .A1(n14816), .A2(n10432), .ZN(n10439) );
  NAND2_X1 U12837 ( .A1(n14812), .A2(n10433), .ZN(n10436) );
  INV_X1 U12838 ( .A(n10434), .ZN(n10435) );
  OAI211_X1 U12839 ( .C1(n10437), .C2(n13282), .A(n10436), .B(n10435), .ZN(
        n10438) );
  AOI211_X1 U12840 ( .C1(n6605), .C2(n13276), .A(n10439), .B(n10438), .ZN(
        n10440) );
  OAI21_X1 U12841 ( .B1(n10442), .B2(n10441), .A(n10440), .ZN(P2_U3202) );
  INV_X1 U12842 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10443) );
  OAI22_X1 U12843 ( .A1(n13642), .A2(n8548), .B1(n10443), .B2(n13639), .ZN(
        n10446) );
  NOR2_X1 U12844 ( .A1(n13659), .A2(n10444), .ZN(n10445) );
  AOI211_X1 U12845 ( .C1(n13655), .C2(n6481), .A(n10446), .B(n10445), .ZN(
        n10450) );
  NAND2_X1 U12846 ( .A1(n10448), .A2(n13642), .ZN(n10449) );
  OAI211_X1 U12847 ( .C1(n13636), .C2(n10451), .A(n10450), .B(n10449), .ZN(
        P2_U3264) );
  INV_X1 U12848 ( .A(n14894), .ZN(n13362) );
  OAI222_X1 U12849 ( .A1(n13819), .A2(n10453), .B1(n13817), .B2(n10452), .C1(
        n13362), .C2(P2_U3088), .ZN(P2_U3311) );
  XNOR2_X1 U12850 ( .A(n10454), .B(n10456), .ZN(n15047) );
  OAI211_X1 U12851 ( .C1(n10457), .C2(n10456), .A(n10455), .B(n13019), .ZN(
        n10460) );
  OAI22_X1 U12852 ( .A1(n11147), .A2(n12962), .B1(n10538), .B2(n12964), .ZN(
        n10458) );
  INV_X1 U12853 ( .A(n10458), .ZN(n10459) );
  AND2_X1 U12854 ( .A1(n10460), .A2(n10459), .ZN(n15048) );
  MUX2_X1 U12855 ( .A(n10461), .B(n15048), .S(n15030), .Z(n10463) );
  AOI22_X1 U12856 ( .A1(n15016), .A2(n15051), .B1(n15014), .B2(n10522), .ZN(
        n10462) );
  OAI211_X1 U12857 ( .C1(n11466), .C2(n15047), .A(n10463), .B(n10462), .ZN(
        P3_U3229) );
  INV_X1 U12858 ( .A(n10464), .ZN(n10473) );
  INV_X1 U12859 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n14837) );
  OAI22_X1 U12860 ( .A1(n13642), .A2(n10465), .B1(n14837), .B2(n13639), .ZN(
        n10468) );
  NOR2_X1 U12861 ( .A1(n13589), .A2(n10466), .ZN(n10467) );
  AOI211_X1 U12862 ( .C1(n10469), .C2(n13646), .A(n10468), .B(n10467), .ZN(
        n10472) );
  NAND2_X1 U12863 ( .A1(n13656), .A2(n10470), .ZN(n10471) );
  OAI211_X1 U12864 ( .C1(n13595), .C2(n10473), .A(n10472), .B(n10471), .ZN(
        P2_U3263) );
  OAI21_X1 U12865 ( .B1(n10475), .B2(n14729), .A(n10474), .ZN(n10476) );
  NOR2_X1 U12866 ( .A1(n10476), .A2(n14294), .ZN(n14727) );
  XNOR2_X1 U12867 ( .A(n10476), .B(n9680), .ZN(n10479) );
  INV_X1 U12868 ( .A(n12471), .ZN(n10478) );
  MUX2_X1 U12869 ( .A(n10479), .B(n10478), .S(n13977), .Z(n10484) );
  OAI21_X1 U12870 ( .B1(n12471), .B2(n10481), .A(n10480), .ZN(n14732) );
  AOI21_X1 U12871 ( .B1(n14732), .B2(n14777), .A(n10482), .ZN(n10483) );
  OAI21_X1 U12872 ( .B1(n10484), .B2(n14710), .A(n10483), .ZN(n14730) );
  AOI21_X1 U12873 ( .B1(n14727), .B2(n14150), .A(n14730), .ZN(n10499) );
  NAND2_X1 U12874 ( .A1(n10486), .A2(n10485), .ZN(n10487) );
  INV_X1 U12875 ( .A(n10488), .ZN(n10490) );
  NAND2_X1 U12876 ( .A1(n10491), .A2(n14609), .ZN(n12464) );
  INV_X1 U12877 ( .A(n12464), .ZN(n10492) );
  NAND2_X1 U12878 ( .A1(n14282), .A2(n10492), .ZN(n10639) );
  INV_X1 U12879 ( .A(n10639), .ZN(n14721) );
  INV_X1 U12880 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10493) );
  OAI22_X1 U12881 ( .A1(n14282), .A2(n10494), .B1(n10493), .B2(n14252), .ZN(
        n10497) );
  INV_X1 U12882 ( .A(n10495), .ZN(n14606) );
  NOR2_X1 U12883 ( .A1(n14258), .A2(n14729), .ZN(n10496) );
  AOI211_X1 U12884 ( .C1(n14721), .C2(n14732), .A(n10497), .B(n10496), .ZN(
        n10498) );
  OAI21_X1 U12885 ( .B1(n10499), .B2(n14724), .A(n10498), .ZN(P1_U3292) );
  INV_X1 U12886 ( .A(n14816), .ZN(n13284) );
  INV_X1 U12887 ( .A(n13282), .ZN(n13298) );
  AOI22_X1 U12888 ( .A1(n13298), .A2(n10500), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10501) );
  OAI21_X1 U12889 ( .B1(n10502), .B2(n13321), .A(n10501), .ZN(n10507) );
  AOI211_X1 U12890 ( .C1(n10505), .C2(n10504), .A(n14808), .B(n10503), .ZN(
        n10506) );
  AOI211_X1 U12891 ( .C1(n13284), .C2(n15241), .A(n10507), .B(n10506), .ZN(
        n10508) );
  INV_X1 U12892 ( .A(n10508), .ZN(P2_U3190) );
  INV_X1 U12893 ( .A(n10509), .ZN(n10517) );
  MUX2_X1 U12894 ( .A(n10510), .B(P1_REG2_REG_3__SCAN_IN), .S(n14724), .Z(
        n10511) );
  INV_X1 U12895 ( .A(n10511), .ZN(n10516) );
  NOR2_X2 U12896 ( .A1(n14102), .A2(n14609), .ZN(n14720) );
  NAND2_X1 U12897 ( .A1(n14720), .A2(n14749), .ZN(n14098) );
  NOR2_X1 U12898 ( .A1(n14098), .A2(n10512), .ZN(n10514) );
  OAI22_X1 U12899 ( .A1(n14258), .A2(n12280), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14252), .ZN(n10513) );
  NOR2_X1 U12900 ( .A1(n10514), .A2(n10513), .ZN(n10515) );
  OAI211_X1 U12901 ( .C1(n10517), .C2(n10639), .A(n10516), .B(n10515), .ZN(
        P1_U3290) );
  INV_X1 U12902 ( .A(n10518), .ZN(n10520) );
  OAI222_X1 U12903 ( .A1(P3_U3151), .A2(n10521), .B1(n6484), .B2(n10520), .C1(
        n10519), .C2(n13143), .ZN(P3_U3275) );
  INV_X1 U12904 ( .A(n10522), .ZN(n10543) );
  XNOR2_X1 U12905 ( .A(n10523), .B(n10559), .ZN(n10530) );
  XNOR2_X1 U12906 ( .A(n10530), .B(n10538), .ZN(n10566) );
  INV_X1 U12907 ( .A(n10566), .ZN(n10527) );
  INV_X1 U12908 ( .A(n10524), .ZN(n10525) );
  NOR2_X1 U12909 ( .A1(n10525), .A2(n12721), .ZN(n10563) );
  INV_X1 U12910 ( .A(n10563), .ZN(n10526) );
  NAND2_X1 U12911 ( .A1(n10527), .A2(n10526), .ZN(n10528) );
  NOR2_X1 U12912 ( .A1(n10529), .A2(n10528), .ZN(n10564) );
  INV_X1 U12913 ( .A(n10530), .ZN(n10531) );
  XNOR2_X1 U12914 ( .A(n12567), .B(n10533), .ZN(n10534) );
  NOR2_X1 U12915 ( .A1(n10534), .A2(n12719), .ZN(n10748) );
  AOI21_X1 U12916 ( .B1(n12719), .B2(n10534), .A(n10748), .ZN(n10535) );
  OAI21_X1 U12917 ( .B1(n10536), .B2(n10535), .A(n10750), .ZN(n10537) );
  NAND2_X1 U12918 ( .A1(n10537), .A2(n12680), .ZN(n10542) );
  OAI22_X1 U12919 ( .A1(n11147), .A2(n12697), .B1(n12652), .B2(n10538), .ZN(
        n10539) );
  AOI211_X1 U12920 ( .C1(n15051), .C2(n6478), .A(n10540), .B(n10539), .ZN(
        n10541) );
  OAI211_X1 U12921 ( .C1(n10543), .C2(n12672), .A(n10542), .B(n10541), .ZN(
        P3_U3170) );
  INV_X1 U12922 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10544) );
  MUX2_X1 U12923 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10544), .S(n11211), .Z(
        n10547) );
  OAI21_X1 U12924 ( .B1(n10547), .B2(n10546), .A(n11000), .ZN(n10548) );
  NAND2_X1 U12925 ( .A1(n10548), .A2(n14680), .ZN(n10557) );
  INV_X1 U12926 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n11279) );
  MUX2_X1 U12927 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n11279), .S(n11211), .Z(
        n10551) );
  AOI21_X1 U12928 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10977), .A(n10549), 
        .ZN(n10550) );
  NAND2_X1 U12929 ( .A1(n10550), .A2(n10551), .ZN(n11003) );
  OAI21_X1 U12930 ( .B1(n10551), .B2(n10550), .A(n11003), .ZN(n10555) );
  NAND2_X1 U12931 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11776)
         );
  NAND2_X1 U12932 ( .A1(n13986), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n10552) );
  OAI211_X1 U12933 ( .C1(n14023), .C2(n10553), .A(n11776), .B(n10552), .ZN(
        n10554) );
  AOI21_X1 U12934 ( .B1(n10555), .B2(n14027), .A(n10554), .ZN(n10556) );
  NAND2_X1 U12935 ( .A1(n10557), .A2(n10556), .ZN(P1_U3255) );
  AOI21_X1 U12936 ( .B1(n6477), .B2(n10559), .A(n10558), .ZN(n10562) );
  OR2_X1 U12937 ( .A1(n12652), .A2(n10560), .ZN(n10561) );
  OAI211_X1 U12938 ( .C1(n10753), .C2(n12697), .A(n10562), .B(n10561), .ZN(
        n10568) );
  OR2_X1 U12939 ( .A1(n10529), .A2(n10563), .ZN(n10565) );
  AOI211_X1 U12940 ( .C1(n10566), .C2(n10565), .A(n12689), .B(n10564), .ZN(
        n10567) );
  AOI211_X1 U12941 ( .C1(n10569), .C2(n12700), .A(n10568), .B(n10567), .ZN(
        n10570) );
  INV_X1 U12942 ( .A(n10570), .ZN(P3_U3158) );
  INV_X1 U12943 ( .A(SI_21_), .ZN(n10572) );
  OAI222_X1 U12944 ( .A1(n6484), .A2(n10573), .B1(n13143), .B2(n10572), .C1(
        P3_U3151), .C2(n10571), .ZN(P3_U3274) );
  INV_X1 U12945 ( .A(n10580), .ZN(n10575) );
  XNOR2_X1 U12946 ( .A(n13222), .B(n14932), .ZN(n10710) );
  NAND2_X1 U12947 ( .A1(n13355), .A2(n9793), .ZN(n10711) );
  XNOR2_X1 U12948 ( .A(n10710), .B(n10711), .ZN(n10581) );
  OR2_X1 U12949 ( .A1(n13282), .A2(n10576), .ZN(n10578) );
  OAI211_X1 U12950 ( .C1(n14816), .C2(n10579), .A(n10578), .B(n10577), .ZN(
        n10584) );
  AOI22_X1 U12951 ( .A1(n13306), .A2(n13356), .B1(n13276), .B2(n10580), .ZN(
        n10582) );
  NOR3_X1 U12952 ( .A1(n6605), .A2(n10582), .A3(n10581), .ZN(n10583) );
  AOI211_X1 U12953 ( .C1(n14932), .C2(n14812), .A(n10584), .B(n10583), .ZN(
        n10585) );
  OAI21_X1 U12954 ( .B1(n10714), .B2(n14808), .A(n10585), .ZN(P2_U3199) );
  NAND2_X1 U12955 ( .A1(n10587), .A2(n12457), .ZN(n10590) );
  AOI22_X1 U12956 ( .A1(n12041), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n12040), 
        .B2(n10588), .ZN(n10589) );
  INV_X2 U12957 ( .A(n12293), .ZN(n13972) );
  INV_X1 U12958 ( .A(n12473), .ZN(n10765) );
  NAND2_X1 U12959 ( .A1(n12292), .A2(n12293), .ZN(n10591) );
  NAND2_X1 U12960 ( .A1(n10592), .A2(n12457), .ZN(n10595) );
  AOI22_X1 U12961 ( .A1(n12041), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12040), 
        .B2(n10593), .ZN(n10594) );
  NAND2_X1 U12962 ( .A1(n10595), .A2(n10594), .ZN(n14716) );
  INV_X4 U12963 ( .A(n12049), .ZN(n12439) );
  NAND2_X1 U12964 ( .A1(n12439), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U12965 ( .A1(n12223), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10600) );
  NAND2_X1 U12966 ( .A1(n10596), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10609) );
  OR2_X1 U12967 ( .A1(n10596), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10597) );
  AND2_X1 U12968 ( .A1(n10609), .A2(n10597), .ZN(n14714) );
  NAND2_X1 U12969 ( .A1(n9937), .A2(n14714), .ZN(n10599) );
  NAND2_X1 U12970 ( .A1(n12441), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10598) );
  NAND4_X1 U12971 ( .A1(n10601), .A2(n10600), .A3(n10599), .A4(n10598), .ZN(
        n13971) );
  XNOR2_X1 U12972 ( .A(n14716), .B(n13971), .ZN(n12474) );
  INV_X1 U12973 ( .A(n12474), .ZN(n14707) );
  NAND2_X1 U12974 ( .A1(n14706), .A2(n14707), .ZN(n10603) );
  OR2_X1 U12975 ( .A1(n14716), .A2(n13971), .ZN(n10602) );
  NAND2_X1 U12976 ( .A1(n10603), .A2(n10602), .ZN(n10830) );
  NAND2_X1 U12977 ( .A1(n10604), .A2(n12457), .ZN(n10607) );
  AOI22_X1 U12978 ( .A1(n12041), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n12040), 
        .B2(n10605), .ZN(n10606) );
  NAND2_X1 U12979 ( .A1(n10607), .A2(n10606), .ZN(n12302) );
  NAND2_X1 U12980 ( .A1(n12440), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10614) );
  NAND2_X1 U12981 ( .A1(n12441), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10613) );
  NAND2_X1 U12982 ( .A1(n10609), .A2(n10608), .ZN(n10610) );
  AND2_X1 U12983 ( .A1(n10624), .A2(n10610), .ZN(n11087) );
  NAND2_X1 U12984 ( .A1(n9937), .A2(n11087), .ZN(n10612) );
  NAND2_X1 U12985 ( .A1(n12439), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10611) );
  NAND4_X1 U12986 ( .A1(n10614), .A2(n10613), .A3(n10612), .A4(n10611), .ZN(
        n13970) );
  INV_X1 U12987 ( .A(n13970), .ZN(n10850) );
  XNOR2_X1 U12988 ( .A(n12302), .B(n10850), .ZN(n12477) );
  XNOR2_X1 U12989 ( .A(n10830), .B(n12477), .ZN(n14755) );
  INV_X1 U12990 ( .A(n14755), .ZN(n10640) );
  NAND2_X1 U12991 ( .A1(n12285), .A2(n13973), .ZN(n10615) );
  NAND2_X1 U12992 ( .A1(n12292), .A2(n13972), .ZN(n10617) );
  OR2_X1 U12993 ( .A1(n12292), .A2(n13972), .ZN(n10618) );
  NAND2_X1 U12994 ( .A1(n14708), .A2(n12474), .ZN(n10622) );
  INV_X1 U12995 ( .A(n13971), .ZN(n10620) );
  NAND2_X1 U12996 ( .A1(n14716), .A2(n10620), .ZN(n10621) );
  NAND2_X1 U12997 ( .A1(n10622), .A2(n10621), .ZN(n10853) );
  XNOR2_X1 U12998 ( .A(n10853), .B(n12477), .ZN(n10632) );
  NAND2_X1 U12999 ( .A1(n13971), .A2(n14064), .ZN(n10631) );
  NAND2_X1 U13000 ( .A1(n12439), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10629) );
  NAND2_X1 U13001 ( .A1(n12440), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10628) );
  NAND2_X1 U13002 ( .A1(n10624), .A2(n10623), .ZN(n10625) );
  NAND2_X1 U13003 ( .A1(n10844), .A2(n10625), .ZN(n11363) );
  INV_X1 U13004 ( .A(n11363), .ZN(n14696) );
  NAND2_X1 U13005 ( .A1(n9937), .A2(n14696), .ZN(n10627) );
  NAND2_X1 U13006 ( .A1(n12441), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10626) );
  NAND4_X1 U13007 ( .A1(n10629), .A2(n10628), .A3(n10627), .A4(n10626), .ZN(
        n13969) );
  NAND2_X1 U13008 ( .A1(n13969), .A2(n6479), .ZN(n10630) );
  AND2_X1 U13009 ( .A1(n10631), .A2(n10630), .ZN(n11090) );
  OAI21_X1 U13010 ( .B1(n10632), .B2(n14710), .A(n11090), .ZN(n10633) );
  AOI21_X1 U13011 ( .B1(n14755), .B2(n14777), .A(n10633), .ZN(n14757) );
  MUX2_X1 U13012 ( .A(n9392), .B(n14757), .S(n14282), .Z(n10638) );
  NOR2_X2 U13013 ( .A1(n14717), .A2(n12302), .ZN(n14701) );
  AND2_X1 U13014 ( .A1(n14717), .A2(n12302), .ZN(n10634) );
  NOR2_X1 U13015 ( .A1(n14701), .A2(n10634), .ZN(n14750) );
  INV_X1 U13016 ( .A(n14098), .ZN(n14280) );
  INV_X1 U13017 ( .A(n12302), .ZN(n14752) );
  INV_X1 U13018 ( .A(n11087), .ZN(n10635) );
  OAI22_X1 U13019 ( .A1(n14752), .A2(n14258), .B1(n14252), .B2(n10635), .ZN(
        n10636) );
  AOI21_X1 U13020 ( .B1(n14750), .B2(n14280), .A(n10636), .ZN(n10637) );
  OAI211_X1 U13021 ( .C1(n10640), .C2(n10639), .A(n10638), .B(n10637), .ZN(
        P1_U3286) );
  XNOR2_X1 U13022 ( .A(n10641), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14004) );
  INV_X1 U13023 ( .A(n14004), .ZN(n14001) );
  INV_X1 U13024 ( .A(n11806), .ZN(n10643) );
  OAI222_X1 U13025 ( .A1(P1_U3086), .A2(n14001), .B1(n14391), .B2(n10643), 
        .C1(n10642), .C2(n14396), .ZN(P1_U3338) );
  INV_X1 U13026 ( .A(n14907), .ZN(n13361) );
  OAI222_X1 U13027 ( .A1(n13819), .A2(n10644), .B1(n13803), .B2(n10643), .C1(
        n13361), .C2(P2_U3088), .ZN(P2_U3310) );
  NAND2_X1 U13028 ( .A1(n13947), .A2(n10807), .ZN(n10646) );
  OAI211_X1 U13029 ( .C1(n10810), .C2(n13949), .A(n10646), .B(n10645), .ZN(
        n10657) );
  OAI22_X1 U13030 ( .A1(n12285), .A2(n12231), .B1(n12286), .B2(n12230), .ZN(
        n10647) );
  XOR2_X1 U13031 ( .A(n12020), .B(n10647), .Z(n10655) );
  INV_X1 U13032 ( .A(n10648), .ZN(n10649) );
  NAND2_X1 U13033 ( .A1(n12287), .A2(n12175), .ZN(n10653) );
  NAND2_X1 U13034 ( .A1(n13973), .A2(n12216), .ZN(n10652) );
  NAND2_X1 U13035 ( .A1(n10653), .A2(n10652), .ZN(n10671) );
  AOI211_X1 U13036 ( .C1(n10655), .C2(n10654), .A(n13955), .B(n10674), .ZN(
        n10656) );
  AOI211_X1 U13037 ( .C1(n13952), .C2(n12287), .A(n10657), .B(n10656), .ZN(
        n10658) );
  INV_X1 U13038 ( .A(n10658), .ZN(P1_U3230) );
  INV_X1 U13039 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10659) );
  MUX2_X1 U13040 ( .A(n10659), .B(P2_REG1_REG_10__SCAN_IN), .S(n11395), .Z(
        n10662) );
  OAI21_X1 U13041 ( .B1(n10664), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10660), .ZN(
        n10661) );
  NOR2_X1 U13042 ( .A1(n10661), .A2(n10662), .ZN(n11394) );
  AOI211_X1 U13043 ( .C1(n10662), .C2(n10661), .A(n14901), .B(n11394), .ZN(
        n10670) );
  OAI21_X1 U13044 ( .B1(n10664), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10663), .ZN(
        n10666) );
  MUX2_X1 U13045 ( .A(n11407), .B(P2_REG2_REG_10__SCAN_IN), .S(n11395), .Z(
        n10665) );
  AOI211_X1 U13046 ( .C1(n10666), .C2(n10665), .A(n14852), .B(n11404), .ZN(
        n10669) );
  AND2_X1 U13047 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11204) );
  AOI21_X1 U13048 ( .B1(n14821), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n11204), 
        .ZN(n10667) );
  OAI21_X1 U13049 ( .B1(n11406), .B2(n14839), .A(n10667), .ZN(n10668) );
  OR3_X1 U13050 ( .A1(n10670), .A2(n10669), .A3(n10668), .ZN(P2_U3224) );
  AND2_X1 U13051 ( .A1(n10672), .A2(n10671), .ZN(n10673) );
  OAI22_X1 U13052 ( .A1(n12292), .A2(n12231), .B1(n12293), .B2(n12230), .ZN(
        n10675) );
  XOR2_X1 U13053 ( .A(n12020), .B(n10675), .Z(n11015) );
  AOI22_X1 U13054 ( .A1(n14736), .A2(n12175), .B1(n12216), .B2(n13972), .ZN(
        n11016) );
  XNOR2_X1 U13055 ( .A(n11015), .B(n11016), .ZN(n10676) );
  XNOR2_X1 U13056 ( .A(n11014), .B(n10676), .ZN(n10681) );
  AOI22_X1 U13057 ( .A1(n14064), .A2(n13973), .B1(n13971), .B2(n6479), .ZN(
        n10767) );
  NAND2_X1 U13058 ( .A1(n13947), .A2(n10772), .ZN(n10678) );
  OAI211_X1 U13059 ( .C1(n10767), .C2(n13949), .A(n10678), .B(n10677), .ZN(
        n10679) );
  AOI21_X1 U13060 ( .B1(n13952), .B2(n14736), .A(n10679), .ZN(n10680) );
  OAI21_X1 U13061 ( .B1(n10681), .B2(n13955), .A(n10680), .ZN(P1_U3227) );
  NOR2_X1 U13062 ( .A1(n10697), .A2(n10682), .ZN(n10684) );
  INV_X1 U13063 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n15020) );
  AOI22_X1 U13064 ( .A1(n10702), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15020), 
        .B2(n11256), .ZN(n10685) );
  AOI21_X1 U13065 ( .B1(n6611), .B2(n10685), .A(n11246), .ZN(n10709) );
  INV_X1 U13066 ( .A(n10686), .ZN(n10692) );
  INV_X1 U13067 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n10687) );
  MUX2_X1 U13068 ( .A(n15020), .B(n10687), .S(n13141), .Z(n10688) );
  NAND2_X1 U13069 ( .A1(n10688), .A2(n10702), .ZN(n11249) );
  INV_X1 U13070 ( .A(n10688), .ZN(n10689) );
  NAND2_X1 U13071 ( .A1(n10689), .A2(n11256), .ZN(n10690) );
  AND2_X1 U13072 ( .A1(n11249), .A2(n10690), .ZN(n10691) );
  OAI21_X1 U13073 ( .B1(n10693), .B2(n10692), .A(n10691), .ZN(n11250) );
  INV_X1 U13074 ( .A(n11250), .ZN(n10695) );
  NOR3_X1 U13075 ( .A1(n10693), .A2(n10692), .A3(n10691), .ZN(n10694) );
  OAI21_X1 U13076 ( .B1(n10695), .B2(n10694), .A(n12778), .ZN(n10708) );
  NOR2_X1 U13077 ( .A1(n10697), .A2(n10696), .ZN(n10699) );
  AOI22_X1 U13078 ( .A1(n10702), .A2(P3_REG1_REG_10__SCAN_IN), .B1(n10687), 
        .B2(n11256), .ZN(n10700) );
  AOI21_X1 U13079 ( .B1(n10701), .B2(n10700), .A(n11255), .ZN(n10705) );
  AND2_X1 U13080 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11368) );
  AOI21_X1 U13081 ( .B1(n14987), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11368), 
        .ZN(n10704) );
  NAND2_X1 U13082 ( .A1(n12847), .A2(n10702), .ZN(n10703) );
  OAI211_X1 U13083 ( .C1(n10705), .C2(n15002), .A(n10704), .B(n10703), .ZN(
        n10706) );
  INV_X1 U13084 ( .A(n10706), .ZN(n10707) );
  OAI211_X1 U13085 ( .C1(n10709), .C2(n15008), .A(n10708), .B(n10707), .ZN(
        P3_U3192) );
  INV_X1 U13086 ( .A(n10710), .ZN(n10712) );
  NAND2_X1 U13087 ( .A1(n10712), .A2(n10711), .ZN(n10713) );
  NAND2_X1 U13088 ( .A1(n10714), .A2(n10713), .ZN(n10940) );
  INV_X1 U13089 ( .A(n10940), .ZN(n10718) );
  XNOR2_X1 U13090 ( .A(n14938), .B(n13222), .ZN(n10795) );
  AND2_X1 U13091 ( .A1(n13354), .A2(n13221), .ZN(n10715) );
  OR2_X1 U13092 ( .A1(n10795), .A2(n10715), .ZN(n10932) );
  INV_X1 U13093 ( .A(n10932), .ZN(n10716) );
  AND2_X1 U13094 ( .A1(n10795), .A2(n10715), .ZN(n10933) );
  NOR2_X1 U13095 ( .A1(n10716), .A2(n10933), .ZN(n10717) );
  NAND2_X1 U13096 ( .A1(n10718), .A2(n10717), .ZN(n10799) );
  OAI211_X1 U13097 ( .C1(n10718), .C2(n10717), .A(n10799), .B(n13276), .ZN(
        n10725) );
  NOR2_X1 U13098 ( .A1(n14816), .A2(n10719), .ZN(n10723) );
  OAI21_X1 U13099 ( .B1(n13282), .B2(n10721), .A(n10720), .ZN(n10722) );
  AOI211_X1 U13100 ( .C1(n14938), .C2(n14812), .A(n10723), .B(n10722), .ZN(
        n10724) );
  NAND2_X1 U13101 ( .A1(n10725), .A2(n10724), .ZN(P2_U3211) );
  OR2_X1 U13102 ( .A1(n14938), .A2(n13354), .ZN(n10728) );
  NAND2_X1 U13103 ( .A1(n10729), .A2(n10728), .ZN(n10777) );
  OR2_X1 U13104 ( .A1(n10804), .A2(n13353), .ZN(n10731) );
  NAND2_X1 U13105 ( .A1(n10732), .A2(n10738), .ZN(n10733) );
  NAND2_X1 U13106 ( .A1(n10951), .A2(n10733), .ZN(n14953) );
  INV_X1 U13107 ( .A(n13353), .ZN(n10929) );
  OR2_X1 U13108 ( .A1(n10804), .A2(n10929), .ZN(n10736) );
  NAND2_X1 U13109 ( .A1(n10804), .A2(n10929), .ZN(n10737) );
  XNOR2_X1 U13110 ( .A(n10956), .B(n10738), .ZN(n10740) );
  OAI22_X1 U13111 ( .A1(n10929), .A2(n13575), .B1(n11202), .B2(n13631), .ZN(
        n10739) );
  AOI21_X1 U13112 ( .B1(n10740), .B2(n13625), .A(n10739), .ZN(n10741) );
  OAI21_X1 U13113 ( .B1(n14953), .B2(n9792), .A(n10741), .ZN(n14956) );
  NAND2_X1 U13114 ( .A1(n14956), .A2(n13642), .ZN(n10747) );
  OAI22_X1 U13115 ( .A1(n13642), .A2(n10742), .B1(n10928), .B2(n13639), .ZN(
        n10745) );
  INV_X1 U13116 ( .A(n10804), .ZN(n14948) );
  NAND2_X1 U13117 ( .A1(n10779), .A2(n14948), .ZN(n10778) );
  INV_X1 U13118 ( .A(n10778), .ZN(n10743) );
  INV_X1 U13119 ( .A(n10954), .ZN(n14955) );
  OAI211_X1 U13120 ( .C1(n10743), .C2(n14955), .A(n13521), .B(n10961), .ZN(
        n14954) );
  NOR2_X1 U13121 ( .A1(n14954), .A2(n13659), .ZN(n10744) );
  AOI211_X1 U13122 ( .C1(n13655), .C2(n10954), .A(n10745), .B(n10744), .ZN(
        n10746) );
  OAI211_X1 U13123 ( .C1(n14953), .C2(n13591), .A(n10747), .B(n10746), .ZN(
        P2_U3257) );
  XNOR2_X1 U13124 ( .A(n12567), .B(n15057), .ZN(n10914) );
  XNOR2_X1 U13125 ( .A(n10914), .B(n12717), .ZN(n10752) );
  INV_X1 U13126 ( .A(n10748), .ZN(n10749) );
  NAND2_X1 U13127 ( .A1(n10750), .A2(n10749), .ZN(n10751) );
  OAI21_X1 U13128 ( .B1(n10752), .B2(n10751), .A(n11049), .ZN(n10760) );
  INV_X1 U13129 ( .A(n10827), .ZN(n10758) );
  OAI22_X1 U13130 ( .A1(n11074), .A2(n12697), .B1(n12652), .B2(n10753), .ZN(
        n10754) );
  INV_X1 U13131 ( .A(n10754), .ZN(n10757) );
  AOI21_X1 U13132 ( .B1(n6478), .B2(n15057), .A(n10755), .ZN(n10756) );
  OAI211_X1 U13133 ( .C1(n12672), .C2(n10758), .A(n10757), .B(n10756), .ZN(
        n10759) );
  AOI21_X1 U13134 ( .B1(n10760), .B2(n12680), .A(n10759), .ZN(n10761) );
  INV_X1 U13135 ( .A(n10761), .ZN(P3_U3167) );
  INV_X1 U13136 ( .A(n10762), .ZN(n10763) );
  XNOR2_X1 U13137 ( .A(n10764), .B(n12473), .ZN(n14738) );
  XNOR2_X1 U13138 ( .A(n10766), .B(n10765), .ZN(n10768) );
  OAI21_X1 U13139 ( .B1(n10768), .B2(n14710), .A(n10767), .ZN(n14733) );
  INV_X1 U13140 ( .A(n14733), .ZN(n10769) );
  MUX2_X1 U13141 ( .A(n9335), .B(n10769), .S(n14282), .Z(n10776) );
  INV_X1 U13142 ( .A(n10770), .ZN(n14718) );
  AOI211_X1 U13143 ( .C1(n14736), .C2(n10771), .A(n14294), .B(n14718), .ZN(
        n14734) );
  INV_X1 U13144 ( .A(n10772), .ZN(n10773) );
  OAI22_X1 U13145 ( .A1(n14258), .A2(n12292), .B1(n14252), .B2(n10773), .ZN(
        n10774) );
  AOI21_X1 U13146 ( .B1(n14734), .B2(n14720), .A(n10774), .ZN(n10775) );
  OAI211_X1 U13147 ( .C1(n14262), .C2(n14738), .A(n10776), .B(n10775), .ZN(
        P1_U3288) );
  XNOR2_X1 U13148 ( .A(n10777), .B(n10782), .ZN(n14952) );
  OAI211_X1 U13149 ( .C1(n10779), .C2(n14948), .A(n10778), .B(n13521), .ZN(
        n14947) );
  INV_X1 U13150 ( .A(n10800), .ZN(n10780) );
  INV_X1 U13151 ( .A(n13639), .ZN(n13654) );
  AOI22_X1 U13152 ( .A1(n13655), .A2(n10804), .B1(n10780), .B2(n13654), .ZN(
        n10781) );
  OAI21_X1 U13153 ( .B1(n14947), .B2(n13659), .A(n10781), .ZN(n10788) );
  XNOR2_X1 U13154 ( .A(n10783), .B(n10782), .ZN(n10786) );
  NAND2_X1 U13155 ( .A1(n13354), .A2(n13628), .ZN(n10785) );
  NAND2_X1 U13156 ( .A1(n13352), .A2(n13466), .ZN(n10784) );
  AND2_X1 U13157 ( .A1(n10785), .A2(n10784), .ZN(n10801) );
  OAI21_X1 U13158 ( .B1(n10786), .B2(n13603), .A(n10801), .ZN(n14949) );
  MUX2_X1 U13159 ( .A(n14949), .B(P2_REG2_REG_7__SCAN_IN), .S(n13595), .Z(
        n10787) );
  AOI211_X1 U13160 ( .C1(n14952), .C2(n13656), .A(n10788), .B(n10787), .ZN(
        n10789) );
  INV_X1 U13161 ( .A(n10789), .ZN(P2_U3258) );
  NOR2_X1 U13162 ( .A1(n13329), .A2(n10790), .ZN(n10796) );
  XNOR2_X1 U13163 ( .A(n10804), .B(n13178), .ZN(n10924) );
  NAND2_X1 U13164 ( .A1(n13353), .A2(n13221), .ZN(n10791) );
  NAND2_X1 U13165 ( .A1(n10924), .A2(n10791), .ZN(n10934) );
  INV_X1 U13166 ( .A(n10924), .ZN(n10793) );
  INV_X1 U13167 ( .A(n10791), .ZN(n10792) );
  NAND2_X1 U13168 ( .A1(n10793), .A2(n10792), .ZN(n10935) );
  NAND2_X1 U13169 ( .A1(n10934), .A2(n10935), .ZN(n10797) );
  AOI21_X1 U13170 ( .B1(n10799), .B2(n10797), .A(n14808), .ZN(n10794) );
  AOI21_X1 U13171 ( .B1(n10796), .B2(n10795), .A(n10794), .ZN(n10806) );
  INV_X1 U13172 ( .A(n10933), .ZN(n10798) );
  AOI21_X1 U13173 ( .B1(n10799), .B2(n10798), .A(n10797), .ZN(n10926) );
  NOR2_X1 U13174 ( .A1(n14816), .A2(n10800), .ZN(n10803) );
  OAI22_X1 U13175 ( .A1(n13282), .A2(n10801), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8657), .ZN(n10802) );
  AOI211_X1 U13176 ( .C1(n10804), .C2(n14812), .A(n10803), .B(n10802), .ZN(
        n10805) );
  OAI21_X1 U13177 ( .B1(n10806), .B2(n10926), .A(n10805), .ZN(P2_U3185) );
  AOI22_X1 U13178 ( .A1(n14715), .A2(n12287), .B1(n10807), .B2(n14713), .ZN(
        n10808) );
  OAI21_X1 U13179 ( .B1(n14270), .B2(n10809), .A(n10808), .ZN(n10814) );
  NAND2_X1 U13180 ( .A1(n10811), .A2(n10810), .ZN(n10812) );
  MUX2_X1 U13181 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10812), .S(n14282), .Z(
        n10813) );
  AOI211_X1 U13182 ( .C1(n14703), .C2(n10815), .A(n10814), .B(n10813), .ZN(
        n10816) );
  INV_X1 U13183 ( .A(n10816), .ZN(P1_U3289) );
  INV_X1 U13184 ( .A(n10817), .ZN(n10820) );
  OAI22_X1 U13185 ( .A1(n10818), .A2(P3_U3151), .B1(SI_22_), .B2(n13143), .ZN(
        n10819) );
  AOI21_X1 U13186 ( .B1(n10820), .B2(n10968), .A(n10819), .ZN(P3_U3273) );
  XOR2_X1 U13187 ( .A(n10821), .B(n10822), .Z(n15053) );
  OAI21_X1 U13188 ( .B1(n10824), .B2(n7979), .A(n10823), .ZN(n10825) );
  AOI222_X1 U13189 ( .A1(n13019), .A2(n10825), .B1(n12719), .B2(n13023), .C1(
        n11134), .C2(n13022), .ZN(n15054) );
  MUX2_X1 U13190 ( .A(n10826), .B(n15054), .S(n15030), .Z(n10829) );
  AOI22_X1 U13191 ( .A1(n15016), .A2(n15057), .B1(n15014), .B2(n10827), .ZN(
        n10828) );
  OAI211_X1 U13192 ( .C1(n11466), .C2(n15053), .A(n10829), .B(n10828), .ZN(
        P3_U3228) );
  NAND2_X1 U13193 ( .A1(n10830), .A2(n12477), .ZN(n10832) );
  OR2_X1 U13194 ( .A1(n12302), .A2(n13970), .ZN(n10831) );
  NAND2_X1 U13195 ( .A1(n10832), .A2(n10831), .ZN(n14698) );
  NAND2_X1 U13196 ( .A1(n10833), .A2(n12457), .ZN(n10836) );
  AOI22_X1 U13197 ( .A1(n12041), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12040), 
        .B2(n10834), .ZN(n10835) );
  NAND2_X1 U13198 ( .A1(n10836), .A2(n10835), .ZN(n14697) );
  XNOR2_X1 U13199 ( .A(n14697), .B(n11350), .ZN(n14699) );
  NAND2_X1 U13200 ( .A1(n14698), .A2(n14699), .ZN(n10838) );
  OR2_X1 U13201 ( .A1(n14697), .A2(n13969), .ZN(n10837) );
  NAND2_X1 U13202 ( .A1(n10838), .A2(n10837), .ZN(n10881) );
  NAND2_X1 U13203 ( .A1(n10839), .A2(n12457), .ZN(n10842) );
  AOI22_X1 U13204 ( .A1(n12041), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n12040), 
        .B2(n10840), .ZN(n10841) );
  NAND2_X1 U13205 ( .A1(n10842), .A2(n10841), .ZN(n12314) );
  NAND2_X1 U13206 ( .A1(n12439), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n10849) );
  NAND2_X1 U13207 ( .A1(n12440), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10848) );
  AND2_X1 U13208 ( .A1(n10844), .A2(n10843), .ZN(n10845) );
  NOR2_X1 U13209 ( .A1(n10901), .A2(n10845), .ZN(n11430) );
  NAND2_X1 U13210 ( .A1(n9937), .A2(n11430), .ZN(n10847) );
  NAND2_X1 U13211 ( .A1(n12441), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10846) );
  NAND4_X1 U13212 ( .A1(n10849), .A2(n10848), .A3(n10847), .A4(n10846), .ZN(
        n13968) );
  XNOR2_X1 U13213 ( .A(n12314), .B(n13968), .ZN(n12479) );
  XNOR2_X1 U13214 ( .A(n10881), .B(n12479), .ZN(n14774) );
  AND2_X1 U13215 ( .A1(n12302), .A2(n10850), .ZN(n10852) );
  OR2_X1 U13216 ( .A1(n12302), .A2(n10850), .ZN(n10851) );
  INV_X1 U13217 ( .A(n14699), .ZN(n10855) );
  NOR2_X1 U13218 ( .A1(n14697), .A2(n11350), .ZN(n10854) );
  OAI21_X1 U13219 ( .B1(n10856), .B2(n12479), .A(n10894), .ZN(n14771) );
  NAND2_X1 U13220 ( .A1(n14282), .A2(n14770), .ZN(n14126) );
  INV_X1 U13221 ( .A(n14126), .ZN(n14284) );
  NAND2_X1 U13222 ( .A1(n14701), .A2(n14760), .ZN(n14700) );
  AOI21_X1 U13223 ( .B1(n14700), .B2(n12314), .A(n14294), .ZN(n10857) );
  NAND2_X1 U13224 ( .A1(n10857), .A2(n10897), .ZN(n14767) );
  NAND2_X1 U13225 ( .A1(n12223), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10862) );
  NAND2_X1 U13226 ( .A1(n12441), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10861) );
  INV_X1 U13227 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10858) );
  XNOR2_X1 U13228 ( .A(n10901), .B(n10858), .ZN(n11532) );
  NAND2_X1 U13229 ( .A1(n9937), .A2(n11532), .ZN(n10860) );
  NAND2_X1 U13230 ( .A1(n12439), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10859) );
  NAND4_X1 U13231 ( .A1(n10862), .A2(n10861), .A3(n10860), .A4(n10859), .ZN(
        n13967) );
  AOI22_X1 U13232 ( .A1(n14064), .A2(n13969), .B1(n13967), .B2(n6479), .ZN(
        n14766) );
  INV_X1 U13233 ( .A(n14766), .ZN(n10863) );
  AOI22_X1 U13234 ( .A1(n10863), .A2(n14282), .B1(n11430), .B2(n14713), .ZN(
        n10864) );
  OAI21_X1 U13235 ( .B1(n10865), .B2(n14282), .A(n10864), .ZN(n10866) );
  AOI21_X1 U13236 ( .B1(n12314), .B2(n14715), .A(n10866), .ZN(n10867) );
  OAI21_X1 U13237 ( .B1(n14767), .B2(n14270), .A(n10867), .ZN(n10868) );
  AOI21_X1 U13238 ( .B1(n14771), .B2(n14284), .A(n10868), .ZN(n10869) );
  OAI21_X1 U13239 ( .B1(n14774), .B2(n14262), .A(n10869), .ZN(P1_U3284) );
  INV_X1 U13240 ( .A(n10870), .ZN(n10879) );
  INV_X1 U13241 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10871) );
  OAI22_X1 U13242 ( .A1(n14282), .A2(n9217), .B1(n10871), .B2(n14252), .ZN(
        n10872) );
  AOI21_X1 U13243 ( .B1(n14715), .B2(n10873), .A(n10872), .ZN(n10874) );
  OAI21_X1 U13244 ( .B1(n14270), .B2(n10875), .A(n10874), .ZN(n10876) );
  AOI21_X1 U13245 ( .B1(n14703), .B2(n10877), .A(n10876), .ZN(n10878) );
  OAI21_X1 U13246 ( .B1(n14724), .B2(n10879), .A(n10878), .ZN(P1_U3291) );
  INV_X1 U13247 ( .A(n12479), .ZN(n10880) );
  NAND2_X1 U13248 ( .A1(n10881), .A2(n10880), .ZN(n10883) );
  OR2_X1 U13249 ( .A1(n12314), .A2(n13968), .ZN(n10882) );
  NAND2_X1 U13250 ( .A1(n10883), .A2(n10882), .ZN(n10973) );
  NAND2_X1 U13251 ( .A1(n10884), .A2(n12457), .ZN(n10887) );
  AOI22_X1 U13252 ( .A1(n12040), .A2(n10885), .B1(n12041), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n10886) );
  INV_X1 U13253 ( .A(n13967), .ZN(n10888) );
  NAND2_X1 U13254 ( .A1(n14778), .A2(n10888), .ZN(n10889) );
  XNOR2_X1 U13255 ( .A(n10973), .B(n12478), .ZN(n14783) );
  INV_X1 U13256 ( .A(n14783), .ZN(n10913) );
  INV_X1 U13257 ( .A(n10894), .ZN(n10891) );
  INV_X1 U13258 ( .A(n13968), .ZN(n10890) );
  AND2_X1 U13259 ( .A1(n12314), .A2(n10890), .ZN(n10892) );
  OAI21_X1 U13260 ( .B1(n10891), .B2(n10892), .A(n12478), .ZN(n10895) );
  NAND3_X1 U13261 ( .A1(n10895), .A2(n14770), .A3(n10981), .ZN(n10896) );
  NAND2_X1 U13262 ( .A1(n13968), .A2(n14064), .ZN(n11528) );
  NAND2_X1 U13263 ( .A1(n10896), .A2(n11528), .ZN(n14781) );
  AOI211_X1 U13264 ( .C1(n14778), .C2(n10897), .A(n14294), .B(n10993), .ZN(
        n10908) );
  NAND2_X1 U13265 ( .A1(n12440), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10906) );
  NAND2_X1 U13266 ( .A1(n12439), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n10905) );
  NAND2_X1 U13267 ( .A1(n10901), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10899) );
  INV_X1 U13268 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10898) );
  NAND2_X1 U13269 ( .A1(n10899), .A2(n10898), .ZN(n10902) );
  AND2_X1 U13270 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n10900) );
  NAND2_X1 U13271 ( .A1(n10901), .A2(n10900), .ZN(n10983) );
  AND2_X1 U13272 ( .A1(n10902), .A2(n10983), .ZN(n11727) );
  NAND2_X1 U13273 ( .A1(n9937), .A2(n11727), .ZN(n10904) );
  NAND2_X1 U13274 ( .A1(n12441), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10903) );
  NAND4_X1 U13275 ( .A1(n10906), .A2(n10905), .A3(n10904), .A4(n10903), .ZN(
        n13966) );
  NAND2_X1 U13276 ( .A1(n13966), .A2(n6479), .ZN(n11529) );
  INV_X1 U13277 ( .A(n11529), .ZN(n10907) );
  NOR2_X1 U13278 ( .A1(n10908), .A2(n10907), .ZN(n14779) );
  AOI22_X1 U13279 ( .A1(n14724), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11532), 
        .B2(n14713), .ZN(n10910) );
  NAND2_X1 U13280 ( .A1(n14778), .A2(n14715), .ZN(n10909) );
  OAI211_X1 U13281 ( .C1(n14779), .C2(n14270), .A(n10910), .B(n10909), .ZN(
        n10911) );
  AOI21_X1 U13282 ( .B1(n14781), .B2(n14282), .A(n10911), .ZN(n10912) );
  OAI21_X1 U13283 ( .B1(n10913), .B2(n14262), .A(n10912), .ZN(P1_U3283) );
  INV_X1 U13284 ( .A(n11049), .ZN(n10916) );
  INV_X1 U13285 ( .A(n10914), .ZN(n10915) );
  NOR2_X1 U13286 ( .A1(n10915), .A2(n12717), .ZN(n11047) );
  NOR2_X1 U13287 ( .A1(n10916), .A2(n11047), .ZN(n10918) );
  XNOR2_X1 U13288 ( .A(n12567), .B(n15064), .ZN(n11050) );
  XNOR2_X1 U13289 ( .A(n11050), .B(n11134), .ZN(n10917) );
  NAND2_X1 U13290 ( .A1(n10918), .A2(n10917), .ZN(n11071) );
  OAI211_X1 U13291 ( .C1(n10918), .C2(n10917), .A(n11071), .B(n12680), .ZN(
        n10923) );
  AND2_X1 U13292 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n12729) );
  AOI21_X1 U13293 ( .B1(n6477), .B2(n15064), .A(n12729), .ZN(n10920) );
  OR2_X1 U13294 ( .A1(n12697), .A2(n11270), .ZN(n10919) );
  OAI211_X1 U13295 ( .C1(n11147), .C2(n12652), .A(n10920), .B(n10919), .ZN(
        n10921) );
  AOI21_X1 U13296 ( .B1(n12700), .B2(n11152), .A(n10921), .ZN(n10922) );
  NAND2_X1 U13297 ( .A1(n10923), .A2(n10922), .ZN(P3_U3179) );
  NOR3_X1 U13298 ( .A1(n13329), .A2(n10929), .A3(n10924), .ZN(n10925) );
  AOI21_X1 U13299 ( .B1(n10926), .B2(n13276), .A(n10925), .ZN(n10945) );
  XNOR2_X1 U13300 ( .A(n10954), .B(n13222), .ZN(n11033) );
  NAND2_X1 U13301 ( .A1(n13352), .A2(n13221), .ZN(n11029) );
  XNOR2_X1 U13302 ( .A(n11033), .B(n11029), .ZN(n10944) );
  OAI22_X1 U13303 ( .A1(n14800), .A2(n11202), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10927), .ZN(n10931) );
  OAI22_X1 U13304 ( .A1(n14801), .A2(n10929), .B1(n10928), .B2(n14816), .ZN(
        n10930) );
  AOI211_X1 U13305 ( .C1(n10954), .C2(n14812), .A(n10931), .B(n10930), .ZN(
        n10943) );
  NAND2_X1 U13306 ( .A1(n10934), .A2(n10932), .ZN(n10939) );
  NAND2_X1 U13307 ( .A1(n10934), .A2(n10933), .ZN(n10936) );
  AND2_X1 U13308 ( .A1(n10936), .A2(n10935), .ZN(n10937) );
  INV_X1 U13309 ( .A(n11037), .ZN(n10941) );
  NAND2_X1 U13310 ( .A1(n10941), .A2(n13276), .ZN(n10942) );
  OAI211_X1 U13311 ( .C1(n10945), .C2(n10944), .A(n10943), .B(n10942), .ZN(
        P2_U3193) );
  NAND2_X1 U13312 ( .A1(n10946), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10947) );
  XNOR2_X1 U13313 ( .A(n10947), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14019) );
  INV_X1 U13314 ( .A(n14019), .ZN(n14012) );
  OAI222_X1 U13315 ( .A1(P1_U3086), .A2(n14012), .B1(n14391), .B2(n12035), 
        .C1(n10948), .C2(n14396), .ZN(P1_U3337) );
  INV_X1 U13316 ( .A(n13385), .ZN(n13370) );
  OAI222_X1 U13317 ( .A1(P2_U3088), .A2(n13370), .B1(n13803), .B2(n12035), 
        .C1(n10949), .C2(n13819), .ZN(P2_U3309) );
  NAND2_X1 U13318 ( .A1(n10954), .A2(n13352), .ZN(n10950) );
  NAND2_X1 U13319 ( .A1(n10951), .A2(n10950), .ZN(n10952) );
  NAND2_X1 U13320 ( .A1(n10952), .A2(n11098), .ZN(n11095) );
  OR2_X1 U13321 ( .A1(n10952), .A2(n11098), .ZN(n10953) );
  NAND2_X1 U13322 ( .A1(n11095), .A2(n10953), .ZN(n14959) );
  INV_X1 U13323 ( .A(n13352), .ZN(n11040) );
  AND2_X1 U13324 ( .A1(n10954), .A2(n11040), .ZN(n10955) );
  XNOR2_X1 U13325 ( .A(n11099), .B(n11098), .ZN(n10958) );
  INV_X1 U13326 ( .A(n13350), .ZN(n11306) );
  OAI22_X1 U13327 ( .A1(n11040), .A2(n13575), .B1(n11306), .B2(n13631), .ZN(
        n10957) );
  AOI21_X1 U13328 ( .B1(n10958), .B2(n13625), .A(n10957), .ZN(n10959) );
  OAI21_X1 U13329 ( .B1(n14959), .B2(n9792), .A(n10959), .ZN(n14962) );
  NAND2_X1 U13330 ( .A1(n14962), .A2(n13642), .ZN(n10967) );
  OAI22_X1 U13331 ( .A1(n13642), .A2(n10960), .B1(n11039), .B2(n13639), .ZN(
        n10965) );
  INV_X1 U13332 ( .A(n11100), .ZN(n14961) );
  INV_X1 U13333 ( .A(n10961), .ZN(n10963) );
  INV_X1 U13334 ( .A(n11106), .ZN(n10962) );
  OAI211_X1 U13335 ( .C1(n14961), .C2(n10963), .A(n10962), .B(n13521), .ZN(
        n14960) );
  NOR2_X1 U13336 ( .A1(n14960), .A2(n13659), .ZN(n10964) );
  AOI211_X1 U13337 ( .C1(n13655), .C2(n11100), .A(n10965), .B(n10964), .ZN(
        n10966) );
  OAI211_X1 U13338 ( .C1(n14959), .C2(n13591), .A(n10967), .B(n10966), .ZN(
        P2_U3256) );
  INV_X1 U13339 ( .A(SI_23_), .ZN(n10972) );
  NAND2_X1 U13340 ( .A1(n10969), .A2(n10968), .ZN(n10971) );
  OAI211_X1 U13341 ( .C1(n10972), .C2(n13143), .A(n10971), .B(n10970), .ZN(
        P3_U3272) );
  NAND2_X1 U13342 ( .A1(n10973), .A2(n12478), .ZN(n10975) );
  OR2_X1 U13343 ( .A1(n14778), .A2(n13967), .ZN(n10974) );
  NAND2_X1 U13344 ( .A1(n10975), .A2(n10974), .ZN(n11208) );
  NAND2_X1 U13345 ( .A1(n10976), .A2(n12457), .ZN(n10979) );
  AOI22_X1 U13346 ( .A1(n12041), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n12040), 
        .B2(n10977), .ZN(n10978) );
  XNOR2_X1 U13347 ( .A(n12320), .B(n13966), .ZN(n12480) );
  INV_X1 U13348 ( .A(n12480), .ZN(n11207) );
  XNOR2_X1 U13349 ( .A(n11208), .B(n11207), .ZN(n14646) );
  INV_X1 U13350 ( .A(n14646), .ZN(n10998) );
  XNOR2_X1 U13351 ( .A(n11227), .B(n12480), .ZN(n10991) );
  NAND2_X1 U13352 ( .A1(n13967), .A2(n14064), .ZN(n10990) );
  NAND2_X1 U13353 ( .A1(n12439), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n10988) );
  NAND2_X1 U13354 ( .A1(n12440), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10987) );
  NAND2_X1 U13355 ( .A1(n10983), .A2(n10982), .ZN(n10984) );
  AND2_X1 U13356 ( .A1(n11221), .A2(n10984), .ZN(n11779) );
  NAND2_X1 U13357 ( .A1(n9937), .A2(n11779), .ZN(n10986) );
  NAND2_X1 U13358 ( .A1(n12441), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10985) );
  NAND4_X1 U13359 ( .A1(n10988), .A2(n10987), .A3(n10986), .A4(n10985), .ZN(
        n13965) );
  NAND2_X1 U13360 ( .A1(n13965), .A2(n6479), .ZN(n10989) );
  AND2_X1 U13361 ( .A1(n10990), .A2(n10989), .ZN(n11725) );
  OAI21_X1 U13362 ( .B1(n10991), .B2(n14710), .A(n11725), .ZN(n14644) );
  INV_X1 U13363 ( .A(n11277), .ZN(n10992) );
  OAI211_X1 U13364 ( .C1(n14643), .C2(n10993), .A(n10992), .B(n14749), .ZN(
        n14642) );
  AOI22_X1 U13365 ( .A1(n14724), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11727), 
        .B2(n14713), .ZN(n10995) );
  NAND2_X1 U13366 ( .A1(n12320), .A2(n14715), .ZN(n10994) );
  OAI211_X1 U13367 ( .C1(n14642), .C2(n14270), .A(n10995), .B(n10994), .ZN(
        n10996) );
  AOI21_X1 U13368 ( .B1(n14644), .B2(n14282), .A(n10996), .ZN(n10997) );
  OAI21_X1 U13369 ( .B1(n10998), .B2(n14262), .A(n10997), .ZN(P1_U3282) );
  INV_X1 U13370 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10999) );
  MUX2_X1 U13371 ( .A(n10999), .B(P1_REG1_REG_13__SCAN_IN), .S(n11217), .Z(
        n11002) );
  OAI21_X1 U13372 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n11211), .A(n11000), 
        .ZN(n11001) );
  NOR2_X1 U13373 ( .A1(n11001), .A2(n11002), .ZN(n11113) );
  AOI211_X1 U13374 ( .C1(n11002), .C2(n11001), .A(n13980), .B(n11113), .ZN(
        n11013) );
  OAI21_X1 U13375 ( .B1(n11211), .B2(P1_REG2_REG_12__SCAN_IN), .A(n11003), 
        .ZN(n11007) );
  INV_X1 U13376 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11004) );
  MUX2_X1 U13377 ( .A(n11004), .B(P1_REG2_REG_13__SCAN_IN), .S(n11217), .Z(
        n11006) );
  INV_X1 U13378 ( .A(n11118), .ZN(n11005) );
  AOI211_X1 U13379 ( .C1(n11007), .C2(n11006), .A(n14686), .B(n11005), .ZN(
        n11012) );
  NAND2_X1 U13380 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n11845)
         );
  INV_X1 U13381 ( .A(n11845), .ZN(n11008) );
  AOI21_X1 U13382 ( .B1(n13986), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n11008), 
        .ZN(n11009) );
  OAI21_X1 U13383 ( .B1(n11010), .B2(n14023), .A(n11009), .ZN(n11011) );
  OR3_X1 U13384 ( .A1(n11013), .A2(n11012), .A3(n11011), .ZN(P1_U3256) );
  NAND2_X1 U13385 ( .A1(n14716), .A2(n12205), .ZN(n11018) );
  NAND2_X1 U13386 ( .A1(n13971), .A2(n12175), .ZN(n11017) );
  NAND2_X1 U13387 ( .A1(n11018), .A2(n11017), .ZN(n11019) );
  XNOR2_X1 U13388 ( .A(n11019), .B(n12172), .ZN(n11081) );
  AND2_X1 U13389 ( .A1(n12216), .A2(n13971), .ZN(n11020) );
  AOI21_X1 U13390 ( .B1(n14716), .B2(n12175), .A(n11020), .ZN(n11082) );
  XNOR2_X1 U13391 ( .A(n11081), .B(n11082), .ZN(n11083) );
  XNOR2_X1 U13392 ( .A(n11084), .B(n11083), .ZN(n11027) );
  OR2_X1 U13393 ( .A1(n12293), .A2(n13917), .ZN(n11022) );
  NAND2_X1 U13394 ( .A1(n13970), .A2(n6479), .ZN(n11021) );
  AND2_X1 U13395 ( .A1(n11022), .A2(n11021), .ZN(n14709) );
  OAI22_X1 U13396 ( .A1(n13949), .A2(n14709), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11023), .ZN(n11024) );
  AOI21_X1 U13397 ( .B1(n14714), .B2(n13947), .A(n11024), .ZN(n11026) );
  NAND2_X1 U13398 ( .A1(n14716), .A2(n13952), .ZN(n11025) );
  OAI211_X1 U13399 ( .C1(n11027), .C2(n13955), .A(n11026), .B(n11025), .ZN(
        P1_U3239) );
  NAND2_X1 U13400 ( .A1(n12718), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n11028) );
  OAI21_X1 U13401 ( .B1(n12877), .B2(n12718), .A(n11028), .ZN(P3_U3519) );
  INV_X1 U13402 ( .A(n11033), .ZN(n11030) );
  NAND2_X1 U13403 ( .A1(n11030), .A2(n11029), .ZN(n11031) );
  XNOR2_X1 U13404 ( .A(n11100), .B(n13222), .ZN(n11194) );
  NAND2_X1 U13405 ( .A1(n13351), .A2(n13221), .ZN(n11195) );
  XNOR2_X1 U13406 ( .A(n11194), .B(n11195), .ZN(n11032) );
  NOR2_X1 U13407 ( .A1(n11198), .A2(n14808), .ZN(n11046) );
  INV_X1 U13408 ( .A(n11032), .ZN(n11036) );
  NAND2_X1 U13409 ( .A1(n11033), .A2(n13276), .ZN(n11034) );
  OAI21_X1 U13410 ( .B1(n11040), .B2(n13329), .A(n11034), .ZN(n11035) );
  NAND3_X1 U13411 ( .A1(n11037), .A2(n11036), .A3(n11035), .ZN(n11044) );
  OAI22_X1 U13412 ( .A1(n14800), .A2(n11306), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11038), .ZN(n11042) );
  OAI22_X1 U13413 ( .A1(n14801), .A2(n11040), .B1(n11039), .B2(n14816), .ZN(
        n11041) );
  NOR2_X1 U13414 ( .A1(n11042), .A2(n11041), .ZN(n11043) );
  OAI211_X1 U13415 ( .C1(n14961), .C2(n13321), .A(n11044), .B(n11043), .ZN(
        n11045) );
  OR2_X1 U13416 ( .A1(n11046), .A2(n11045), .ZN(P2_U3203) );
  XNOR2_X1 U13417 ( .A(n12567), .B(n15080), .ZN(n11372) );
  XNOR2_X1 U13418 ( .A(n11372), .B(n12715), .ZN(n11061) );
  XNOR2_X1 U13419 ( .A(n11132), .B(n12567), .ZN(n11265) );
  AOI211_X1 U13420 ( .C1(n11074), .C2(n11050), .A(n11265), .B(n11047), .ZN(
        n11048) );
  NAND3_X1 U13421 ( .A1(n11049), .A2(n11048), .A3(n11267), .ZN(n11059) );
  INV_X1 U13422 ( .A(n11050), .ZN(n11051) );
  NAND2_X1 U13423 ( .A1(n11051), .A2(n11134), .ZN(n11070) );
  NOR2_X1 U13424 ( .A1(n11052), .A2(n11070), .ZN(n11054) );
  OAI21_X1 U13425 ( .B1(n11052), .B2(n11270), .A(n11265), .ZN(n11053) );
  OAI21_X1 U13426 ( .B1(n11054), .B2(n11265), .A(n11053), .ZN(n11057) );
  INV_X1 U13427 ( .A(n11055), .ZN(n11056) );
  AOI21_X1 U13428 ( .B1(n11061), .B2(n11060), .A(n11375), .ZN(n11067) );
  OAI22_X1 U13429 ( .A1(n11077), .A2(n12652), .B1(n12697), .B2(n11509), .ZN(
        n11062) );
  AOI211_X1 U13430 ( .C1(n11064), .C2(n6477), .A(n11063), .B(n11062), .ZN(
        n11066) );
  NAND2_X1 U13431 ( .A1(n12700), .A2(n11342), .ZN(n11065) );
  OAI211_X1 U13432 ( .C1(n11067), .C2(n12689), .A(n11066), .B(n11065), .ZN(
        P3_U3171) );
  NAND2_X1 U13433 ( .A1(n12718), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n11068) );
  OAI21_X1 U13434 ( .B1(n12572), .B2(n12718), .A(n11068), .ZN(P3_U3520) );
  OAI222_X1 U13435 ( .A1(n11069), .A2(P1_U3086), .B1(n14391), .B2(n12081), 
        .C1(n12082), .C2(n14396), .ZN(P1_U3334) );
  NAND2_X1 U13436 ( .A1(n11071), .A2(n11070), .ZN(n11266) );
  XOR2_X1 U13437 ( .A(n11265), .B(n11266), .Z(n11080) );
  AOI21_X1 U13438 ( .B1(n6478), .B2(n11073), .A(n11072), .ZN(n11076) );
  OR2_X1 U13439 ( .A1(n12652), .A2(n11074), .ZN(n11075) );
  OAI211_X1 U13440 ( .C1(n11077), .C2(n12697), .A(n11076), .B(n11075), .ZN(
        n11078) );
  AOI21_X1 U13441 ( .B1(n12700), .B2(n11137), .A(n11078), .ZN(n11079) );
  OAI21_X1 U13442 ( .B1(n11080), .B2(n12689), .A(n11079), .ZN(P3_U3153) );
  AND2_X1 U13443 ( .A1(n12216), .A2(n13970), .ZN(n11085) );
  AOI21_X1 U13444 ( .B1(n12302), .B2(n12175), .A(n11085), .ZN(n11353) );
  AOI22_X1 U13445 ( .A1(n12302), .A2(n12205), .B1(n12175), .B2(n13970), .ZN(
        n11086) );
  XNOR2_X1 U13446 ( .A(n11086), .B(n12020), .ZN(n11352) );
  XOR2_X1 U13447 ( .A(n11353), .B(n11352), .Z(n11356) );
  XNOR2_X1 U13448 ( .A(n11357), .B(n11356), .ZN(n11093) );
  NAND2_X1 U13449 ( .A1(n13947), .A2(n11087), .ZN(n11089) );
  OAI211_X1 U13450 ( .C1(n11090), .C2(n13949), .A(n11089), .B(n11088), .ZN(
        n11091) );
  AOI21_X1 U13451 ( .B1(n13952), .B2(n12302), .A(n11091), .ZN(n11092) );
  OAI21_X1 U13452 ( .B1(n11093), .B2(n13955), .A(n11092), .ZN(P1_U3213) );
  NAND2_X1 U13453 ( .A1(n11100), .A2(n13351), .ZN(n11094) );
  NAND2_X1 U13454 ( .A1(n11095), .A2(n11094), .ZN(n11096) );
  NAND2_X1 U13455 ( .A1(n11096), .A2(n11157), .ZN(n11156) );
  OR2_X1 U13456 ( .A1(n11096), .A2(n11157), .ZN(n11097) );
  NAND2_X1 U13457 ( .A1(n11156), .A2(n11097), .ZN(n14965) );
  OR2_X1 U13458 ( .A1(n11100), .A2(n11202), .ZN(n11101) );
  XNOR2_X1 U13459 ( .A(n11159), .B(n11157), .ZN(n11104) );
  OAI22_X1 U13460 ( .A1(n11202), .A2(n13575), .B1(n14802), .B2(n13631), .ZN(
        n11103) );
  AOI21_X1 U13461 ( .B1(n11104), .B2(n13625), .A(n11103), .ZN(n11105) );
  OAI21_X1 U13462 ( .B1(n14965), .B2(n9792), .A(n11105), .ZN(n14969) );
  NAND2_X1 U13463 ( .A1(n14969), .A2(n13642), .ZN(n11110) );
  OAI22_X1 U13464 ( .A1(n13642), .A2(n11407), .B1(n11201), .B2(n13639), .ZN(
        n11108) );
  INV_X1 U13465 ( .A(n11189), .ZN(n14968) );
  INV_X1 U13466 ( .A(n11163), .ZN(n11164) );
  OAI211_X1 U13467 ( .C1(n14968), .C2(n11106), .A(n11164), .B(n13521), .ZN(
        n14966) );
  NOR2_X1 U13468 ( .A1(n14966), .A2(n13659), .ZN(n11107) );
  AOI211_X1 U13469 ( .C1(n13655), .C2(n11189), .A(n11108), .B(n11107), .ZN(
        n11109) );
  OAI211_X1 U13470 ( .C1(n14965), .C2(n13591), .A(n11110), .B(n11109), .ZN(
        P2_U3255) );
  OAI222_X1 U13471 ( .A1(n13819), .A2(n11112), .B1(P2_U3088), .B2(n11111), 
        .C1(n13817), .C2(n12081), .ZN(P2_U3306) );
  INV_X1 U13472 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11114) );
  MUX2_X1 U13473 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11114), .S(n11745), .Z(
        n11115) );
  OAI21_X1 U13474 ( .B1(n11116), .B2(n11115), .A(n11736), .ZN(n11128) );
  NAND2_X1 U13475 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n11217), .ZN(n11117) );
  NAND2_X1 U13476 ( .A1(n11118), .A2(n11117), .ZN(n11122) );
  INV_X1 U13477 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11119) );
  MUX2_X1 U13478 ( .A(n11119), .B(P1_REG2_REG_14__SCAN_IN), .S(n11745), .Z(
        n11120) );
  INV_X1 U13479 ( .A(n11120), .ZN(n11121) );
  NAND2_X1 U13480 ( .A1(n11121), .A2(n11122), .ZN(n11746) );
  OAI211_X1 U13481 ( .C1(n11122), .C2(n11121), .A(n14027), .B(n11746), .ZN(
        n11125) );
  NAND2_X1 U13482 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n13832)
         );
  INV_X1 U13483 ( .A(n13832), .ZN(n11123) );
  AOI21_X1 U13484 ( .B1(n13986), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n11123), 
        .ZN(n11124) );
  OAI211_X1 U13485 ( .C1(n14023), .C2(n11126), .A(n11125), .B(n11124), .ZN(
        n11127) );
  AOI21_X1 U13486 ( .B1(n11128), .B2(n14680), .A(n11127), .ZN(n11129) );
  INV_X1 U13487 ( .A(n11129), .ZN(P1_U3257) );
  XNOR2_X1 U13488 ( .A(n11130), .B(n11132), .ZN(n15068) );
  OAI211_X1 U13489 ( .C1(n11133), .C2(n11132), .A(n11131), .B(n13019), .ZN(
        n11136) );
  AOI22_X1 U13490 ( .A1(n13023), .A2(n11134), .B1(n12716), .B2(n13022), .ZN(
        n11135) );
  OAI211_X1 U13491 ( .C1(n15061), .C2(n15068), .A(n11136), .B(n11135), .ZN(
        n15070) );
  AOI21_X1 U13492 ( .B1(n15014), .B2(n11137), .A(n15070), .ZN(n11143) );
  INV_X1 U13493 ( .A(n15068), .ZN(n11141) );
  AND2_X1 U13494 ( .A1(n15030), .A2(n15029), .ZN(n11140) );
  OAI22_X1 U13495 ( .A1(n15067), .A2(n13031), .B1(n15030), .B2(n11138), .ZN(
        n11139) );
  AOI21_X1 U13496 ( .B1(n11141), .B2(n11140), .A(n11139), .ZN(n11142) );
  OAI21_X1 U13497 ( .B1(n11143), .B2(n15032), .A(n11142), .ZN(P3_U3226) );
  XOR2_X1 U13498 ( .A(n11144), .B(n11145), .Z(n15060) );
  AOI21_X1 U13499 ( .B1(n11146), .B2(n11145), .A(n12960), .ZN(n11150) );
  OAI22_X1 U13500 ( .A1(n11270), .A2(n12962), .B1(n11147), .B2(n12964), .ZN(
        n11148) );
  AOI21_X1 U13501 ( .B1(n11150), .B2(n11149), .A(n11148), .ZN(n15059) );
  MUX2_X1 U13502 ( .A(n15059), .B(n11151), .S(n15032), .Z(n11154) );
  AOI22_X1 U13503 ( .A1(n15016), .A2(n15064), .B1(n15014), .B2(n11152), .ZN(
        n11153) );
  OAI211_X1 U13504 ( .C1(n11466), .C2(n15060), .A(n11154), .B(n11153), .ZN(
        P3_U3227) );
  INV_X1 U13505 ( .A(n12065), .ZN(n11323) );
  INV_X1 U13506 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12066) );
  OAI222_X1 U13507 ( .A1(n12257), .A2(P1_U3086), .B1(n14391), .B2(n11323), 
        .C1(n12066), .C2(n14396), .ZN(P1_U3335) );
  XOR2_X1 U13508 ( .A(n11171), .B(n11180), .Z(n11292) );
  INV_X1 U13509 ( .A(n11292), .ZN(n11170) );
  INV_X1 U13510 ( .A(n13348), .ZN(n11621) );
  INV_X1 U13511 ( .A(n11157), .ZN(n11158) );
  NAND2_X1 U13512 ( .A1(n11159), .A2(n11158), .ZN(n11161) );
  OR2_X1 U13513 ( .A1(n11189), .A2(n11306), .ZN(n11160) );
  XOR2_X1 U13514 ( .A(n11171), .B(n11172), .Z(n11162) );
  OAI222_X1 U13515 ( .A1(n13631), .A2(n11621), .B1(n13575), .B2(n11306), .C1(
        n11162), .C2(n13603), .ZN(n11290) );
  NAND2_X1 U13516 ( .A1(n11290), .A2(n13642), .ZN(n11169) );
  INV_X1 U13517 ( .A(n11310), .ZN(n11293) );
  AOI211_X1 U13518 ( .C1(n11310), .C2(n11164), .A(n13221), .B(n6606), .ZN(
        n11291) );
  NOR2_X1 U13519 ( .A1(n11293), .A2(n13589), .ZN(n11167) );
  OAI22_X1 U13520 ( .A1(n13642), .A2(n11165), .B1(n11307), .B2(n13639), .ZN(
        n11166) );
  AOI211_X1 U13521 ( .C1(n11291), .C2(n13646), .A(n11167), .B(n11166), .ZN(
        n11168) );
  OAI211_X1 U13522 ( .C1(n11170), .C2(n13636), .A(n11169), .B(n11168), .ZN(
        P2_U3254) );
  NAND2_X1 U13523 ( .A1(n11310), .A2(n14802), .ZN(n11173) );
  AOI21_X1 U13524 ( .B1(n11175), .B2(n7254), .A(n13603), .ZN(n11177) );
  INV_X1 U13525 ( .A(n13347), .ZN(n14799) );
  OAI22_X1 U13526 ( .A1(n14802), .A2(n13575), .B1(n14799), .B2(n13631), .ZN(
        n11176) );
  AOI21_X1 U13527 ( .B1(n11177), .B2(n11571), .A(n11176), .ZN(n14593) );
  NAND2_X1 U13528 ( .A1(n11293), .A2(n14802), .ZN(n11179) );
  XNOR2_X1 U13529 ( .A(n11565), .B(n7254), .ZN(n14596) );
  NAND2_X1 U13530 ( .A1(n14596), .A2(n13656), .ZN(n11185) );
  OAI22_X1 U13531 ( .A1(n13642), .A2(n11181), .B1(n14815), .B2(n13639), .ZN(
        n11183) );
  INV_X1 U13532 ( .A(n14813), .ZN(n14594) );
  OAI211_X1 U13533 ( .C1(n6606), .C2(n14594), .A(n13521), .B(n11567), .ZN(
        n14592) );
  NOR2_X1 U13534 ( .A1(n14592), .A2(n13659), .ZN(n11182) );
  AOI211_X1 U13535 ( .C1(n13655), .C2(n14813), .A(n11183), .B(n11182), .ZN(
        n11184) );
  OAI211_X1 U13536 ( .C1(n13595), .C2(n14593), .A(n11185), .B(n11184), .ZN(
        P2_U3253) );
  INV_X1 U13537 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11186) );
  INV_X1 U13538 ( .A(n12039), .ZN(n11188) );
  OAI222_X1 U13539 ( .A1(n13819), .A2(n11186), .B1(n13803), .B2(n11188), .C1(
        n13400), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13540 ( .A1(P1_U3086), .A2(n14150), .B1(n14391), .B2(n11188), 
        .C1(n11187), .C2(n14396), .ZN(P1_U3336) );
  XNOR2_X1 U13541 ( .A(n11189), .B(n13222), .ZN(n11301) );
  AND2_X1 U13542 ( .A1(n13350), .A2(n9793), .ZN(n11190) );
  NAND2_X1 U13543 ( .A1(n11301), .A2(n11190), .ZN(n11298) );
  INV_X1 U13544 ( .A(n11301), .ZN(n11192) );
  INV_X1 U13545 ( .A(n11190), .ZN(n11191) );
  NAND2_X1 U13546 ( .A1(n11192), .A2(n11191), .ZN(n11193) );
  AND2_X1 U13547 ( .A1(n11298), .A2(n11193), .ZN(n11200) );
  INV_X1 U13548 ( .A(n11194), .ZN(n11196) );
  NAND2_X1 U13549 ( .A1(n11196), .A2(n11195), .ZN(n11197) );
  OAI211_X1 U13550 ( .C1(n11200), .C2(n11199), .A(n11300), .B(n13276), .ZN(
        n11206) );
  INV_X1 U13551 ( .A(n14800), .ZN(n13318) );
  OAI22_X1 U13552 ( .A1(n14801), .A2(n11202), .B1(n11201), .B2(n14816), .ZN(
        n11203) );
  AOI211_X1 U13553 ( .C1(n13318), .C2(n13349), .A(n11204), .B(n11203), .ZN(
        n11205) );
  OAI211_X1 U13554 ( .C1(n14968), .C2(n13321), .A(n11206), .B(n11205), .ZN(
        P2_U3189) );
  OR2_X1 U13555 ( .A1(n12320), .A2(n13966), .ZN(n11209) );
  NAND2_X1 U13556 ( .A1(n11210), .A2(n12457), .ZN(n11213) );
  AOI22_X1 U13557 ( .A1(n12040), .A2(n11211), .B1(n12041), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n11212) );
  XNOR2_X1 U13558 ( .A(n12329), .B(n13965), .ZN(n12482) );
  NAND2_X1 U13559 ( .A1(n11214), .A2(n12457), .ZN(n11219) );
  NOR2_X1 U13560 ( .A1(n12458), .A2(n11215), .ZN(n11216) );
  AOI21_X1 U13561 ( .B1(n11217), .B2(n12040), .A(n11216), .ZN(n11218) );
  NAND2_X2 U13562 ( .A1(n11219), .A2(n11218), .ZN(n12339) );
  NAND2_X1 U13563 ( .A1(n12223), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11226) );
  NAND2_X1 U13564 ( .A1(n12441), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11225) );
  AND2_X1 U13565 ( .A1(n11221), .A2(n11220), .ZN(n11222) );
  NOR2_X1 U13566 ( .A1(n11232), .A2(n11222), .ZN(n11844) );
  NAND2_X1 U13567 ( .A1(n9937), .A2(n11844), .ZN(n11224) );
  NAND2_X1 U13568 ( .A1(n12439), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11223) );
  NAND4_X1 U13569 ( .A1(n11226), .A2(n11225), .A3(n11224), .A4(n11223), .ZN(
        n13964) );
  INV_X1 U13570 ( .A(n13964), .ZN(n12341) );
  XNOR2_X1 U13571 ( .A(n12339), .B(n12341), .ZN(n12484) );
  XNOR2_X1 U13572 ( .A(n11485), .B(n11475), .ZN(n11470) );
  INV_X1 U13573 ( .A(n13966), .ZN(n11714) );
  OR2_X1 U13574 ( .A1(n12320), .A2(n11714), .ZN(n11228) );
  NAND2_X1 U13575 ( .A1(n11282), .A2(n12482), .ZN(n11231) );
  INV_X1 U13576 ( .A(n13965), .ZN(n11229) );
  OR2_X1 U13577 ( .A1(n12329), .A2(n11229), .ZN(n11230) );
  NAND2_X1 U13578 ( .A1(n11231), .A2(n11230), .ZN(n11476) );
  XNOR2_X1 U13579 ( .A(n11476), .B(n11475), .ZN(n11240) );
  NAND2_X1 U13580 ( .A1(n12223), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11237) );
  NAND2_X1 U13581 ( .A1(n12439), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11236) );
  NOR2_X1 U13582 ( .A1(n11232), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n11233) );
  OR2_X1 U13583 ( .A1(n11491), .A2(n11233), .ZN(n11497) );
  INV_X1 U13584 ( .A(n11497), .ZN(n13834) );
  NAND2_X1 U13585 ( .A1(n9937), .A2(n13834), .ZN(n11235) );
  NAND2_X1 U13586 ( .A1(n12441), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n11234) );
  OR2_X1 U13587 ( .A1(n12010), .A2(n13916), .ZN(n11239) );
  NAND2_X1 U13588 ( .A1(n13965), .A2(n14064), .ZN(n11238) );
  AND2_X1 U13589 ( .A1(n11239), .A2(n11238), .ZN(n11847) );
  OAI21_X1 U13590 ( .B1(n11240), .B2(n14710), .A(n11847), .ZN(n11467) );
  INV_X1 U13591 ( .A(n12339), .ZN(n11243) );
  INV_X1 U13592 ( .A(n12329), .ZN(n11782) );
  INV_X1 U13593 ( .A(n11483), .ZN(n11482) );
  AOI211_X1 U13594 ( .C1(n12339), .C2(n6501), .A(n14294), .B(n11483), .ZN(
        n11468) );
  NAND2_X1 U13595 ( .A1(n11468), .A2(n14720), .ZN(n11242) );
  AOI22_X1 U13596 ( .A1(n14724), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n11844), 
        .B2(n14713), .ZN(n11241) );
  OAI211_X1 U13597 ( .C1(n11243), .C2(n14258), .A(n11242), .B(n11241), .ZN(
        n11244) );
  AOI21_X1 U13598 ( .B1(n11467), .B2(n14282), .A(n11244), .ZN(n11245) );
  OAI21_X1 U13599 ( .B1(n14262), .B2(n11470), .A(n11245), .ZN(P1_U3280) );
  INV_X1 U13600 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11248) );
  AOI21_X1 U13601 ( .B1(n11248), .B2(n11247), .A(n11545), .ZN(n11264) );
  NAND2_X1 U13602 ( .A1(n11250), .A2(n11249), .ZN(n11252) );
  MUX2_X1 U13603 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n13141), .Z(n11551) );
  INV_X1 U13604 ( .A(n11257), .ZN(n11552) );
  XNOR2_X1 U13605 ( .A(n11551), .B(n11552), .ZN(n11251) );
  NAND2_X1 U13606 ( .A1(n11252), .A2(n11251), .ZN(n11556) );
  OAI21_X1 U13607 ( .B1(n11252), .B2(n11251), .A(n11556), .ZN(n11262) );
  INV_X1 U13608 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11253) );
  NOR2_X1 U13609 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11253), .ZN(n11511) );
  AOI21_X1 U13610 ( .B1(n14987), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11511), 
        .ZN(n11254) );
  OAI21_X1 U13611 ( .B1(n14994), .B2(n11257), .A(n11254), .ZN(n11261) );
  INV_X1 U13612 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14582) );
  AOI21_X1 U13613 ( .B1(n14582), .B2(n11258), .A(n11540), .ZN(n11259) );
  NOR2_X1 U13614 ( .A1(n11259), .A2(n15002), .ZN(n11260) );
  AOI211_X1 U13615 ( .C1(n12778), .C2(n11262), .A(n11261), .B(n11260), .ZN(
        n11263) );
  OAI21_X1 U13616 ( .B1(n11264), .B2(n15008), .A(n11263), .ZN(P3_U3193) );
  MUX2_X1 U13617 ( .A(n11266), .B(n7984), .S(n11265), .Z(n11268) );
  XNOR2_X1 U13618 ( .A(n11268), .B(n11267), .ZN(n11275) );
  INV_X1 U13619 ( .A(n12715), .ZN(n11369) );
  AOI21_X1 U13620 ( .B1(n12674), .B2(n11463), .A(n11269), .ZN(n11272) );
  OR2_X1 U13621 ( .A1(n12652), .A2(n11270), .ZN(n11271) );
  OAI211_X1 U13622 ( .C1(n11369), .C2(n12697), .A(n11272), .B(n11271), .ZN(
        n11273) );
  AOI21_X1 U13623 ( .B1(n12700), .B2(n11462), .A(n11273), .ZN(n11274) );
  OAI21_X1 U13624 ( .B1(n11275), .B2(n12689), .A(n11274), .ZN(P3_U3161) );
  XNOR2_X1 U13625 ( .A(n11276), .B(n11283), .ZN(n11325) );
  OAI211_X1 U13626 ( .C1(n11277), .C2(n11782), .A(n14749), .B(n6501), .ZN(
        n11327) );
  INV_X1 U13627 ( .A(n11779), .ZN(n11278) );
  OAI22_X1 U13628 ( .A1(n14282), .A2(n11279), .B1(n11278), .B2(n14252), .ZN(
        n11280) );
  AOI21_X1 U13629 ( .B1(n12329), .B2(n14715), .A(n11280), .ZN(n11281) );
  OAI21_X1 U13630 ( .B1(n11327), .B2(n14270), .A(n11281), .ZN(n11288) );
  XNOR2_X1 U13631 ( .A(n11282), .B(n11283), .ZN(n11284) );
  NAND2_X1 U13632 ( .A1(n11284), .A2(n14770), .ZN(n11328) );
  NAND2_X1 U13633 ( .A1(n13966), .A2(n14064), .ZN(n11286) );
  NAND2_X1 U13634 ( .A1(n13964), .A2(n6479), .ZN(n11285) );
  AND2_X1 U13635 ( .A1(n11286), .A2(n11285), .ZN(n11777) );
  AOI21_X1 U13636 ( .B1(n11328), .B2(n11777), .A(n14724), .ZN(n11287) );
  AOI211_X1 U13637 ( .C1(n11325), .C2(n14703), .A(n11288), .B(n11287), .ZN(
        n11289) );
  INV_X1 U13638 ( .A(n11289), .ZN(P1_U3281) );
  AOI211_X1 U13639 ( .C1(n14951), .C2(n11292), .A(n11291), .B(n11290), .ZN(
        n11297) );
  OAI22_X1 U13640 ( .A1(n11293), .A2(n13794), .B1(n14974), .B2(n8743), .ZN(
        n11294) );
  INV_X1 U13641 ( .A(n11294), .ZN(n11295) );
  OAI21_X1 U13642 ( .B1(n11297), .B2(n14973), .A(n11295), .ZN(P2_U3463) );
  INV_X1 U13643 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U13644 ( .A1(n11310), .A2(n11672), .B1(n14984), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11296) );
  OAI21_X1 U13645 ( .B1(n11297), .B2(n14984), .A(n11296), .ZN(P2_U3510) );
  XNOR2_X1 U13646 ( .A(n11310), .B(n13222), .ZN(n11610) );
  NAND2_X1 U13647 ( .A1(n13349), .A2(n13221), .ZN(n11611) );
  XNOR2_X1 U13648 ( .A(n11610), .B(n11611), .ZN(n11303) );
  AND2_X1 U13649 ( .A1(n11303), .A2(n11298), .ZN(n11299) );
  NAND3_X1 U13650 ( .A1(n11301), .A2(n13306), .A3(n13350), .ZN(n11302) );
  OAI21_X1 U13651 ( .B1(n11300), .B2(n14808), .A(n11302), .ZN(n11305) );
  INV_X1 U13652 ( .A(n11303), .ZN(n11304) );
  NAND2_X1 U13653 ( .A1(n11305), .A2(n11304), .ZN(n11312) );
  NAND2_X1 U13654 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n14860)
         );
  OAI21_X1 U13655 ( .B1(n14801), .B2(n11306), .A(n14860), .ZN(n11309) );
  OAI22_X1 U13656 ( .A1(n14800), .A2(n11621), .B1(n14816), .B2(n11307), .ZN(
        n11308) );
  AOI211_X1 U13657 ( .C1(n11310), .C2(n14812), .A(n11309), .B(n11308), .ZN(
        n11311) );
  OAI211_X1 U13658 ( .C1(n14808), .C2(n11614), .A(n11312), .B(n11311), .ZN(
        P2_U3208) );
  OAI211_X1 U13659 ( .C1(n11314), .C2(n11318), .A(n11313), .B(n13019), .ZN(
        n11316) );
  AOI22_X1 U13660 ( .A1(n13023), .A2(n11505), .B1(n12713), .B2(n13022), .ZN(
        n11315) );
  NAND2_X1 U13661 ( .A1(n11316), .A2(n11315), .ZN(n14578) );
  INV_X1 U13662 ( .A(n14578), .ZN(n11322) );
  XNOR2_X1 U13663 ( .A(n11317), .B(n11318), .ZN(n14580) );
  AOI22_X1 U13664 ( .A1(n15016), .A2(n11510), .B1(n15014), .B2(n11517), .ZN(
        n11319) );
  OAI21_X1 U13665 ( .B1(n11248), .B2(n15030), .A(n11319), .ZN(n11320) );
  AOI21_X1 U13666 ( .B1(n14580), .B2(n13033), .A(n11320), .ZN(n11321) );
  OAI21_X1 U13667 ( .B1(n11322), .B2(n15032), .A(n11321), .ZN(P3_U3222) );
  OAI222_X1 U13668 ( .A1(n13819), .A2(n11324), .B1(P2_U3088), .B2(n6485), .C1(
        n13817), .C2(n11323), .ZN(P2_U3307) );
  NAND2_X1 U13669 ( .A1(n11325), .A2(n14784), .ZN(n11330) );
  INV_X1 U13670 ( .A(n11777), .ZN(n11326) );
  AOI21_X1 U13671 ( .B1(n12329), .B2(n14735), .A(n11326), .ZN(n11329) );
  NAND4_X1 U13672 ( .A1(n11330), .A2(n11329), .A3(n11328), .A4(n11327), .ZN(
        n11332) );
  NAND2_X1 U13673 ( .A1(n11332), .A2(n14798), .ZN(n11331) );
  OAI21_X1 U13674 ( .B1(n14798), .B2(n10544), .A(n11331), .ZN(P1_U3540) );
  INV_X1 U13675 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11334) );
  NAND2_X1 U13676 ( .A1(n11332), .A2(n14748), .ZN(n11333) );
  OAI21_X1 U13677 ( .B1(n14748), .B2(n11334), .A(n11333), .ZN(P1_U3495) );
  XNOR2_X1 U13678 ( .A(n11335), .B(n11338), .ZN(n15082) );
  NAND2_X1 U13679 ( .A1(n11459), .A2(n11458), .ZN(n11457) );
  AND2_X1 U13680 ( .A1(n11457), .A2(n11336), .ZN(n11339) );
  NAND2_X1 U13681 ( .A1(n11457), .A2(n11337), .ZN(n11440) );
  OAI211_X1 U13682 ( .C1(n11339), .C2(n11338), .A(n11440), .B(n13019), .ZN(
        n11341) );
  AOI22_X1 U13683 ( .A1(n12716), .A2(n13023), .B1(n13022), .B2(n11505), .ZN(
        n11340) );
  NAND2_X1 U13684 ( .A1(n11341), .A2(n11340), .ZN(n15083) );
  NAND2_X1 U13685 ( .A1(n15083), .A2(n15030), .ZN(n11346) );
  INV_X1 U13686 ( .A(n11342), .ZN(n11343) );
  OAI22_X1 U13687 ( .A1(n13031), .A2(n15080), .B1(n11343), .B2(n15025), .ZN(
        n11344) );
  AOI21_X1 U13688 ( .B1(P3_REG2_REG_9__SCAN_IN), .B2(n15032), .A(n11344), .ZN(
        n11345) );
  OAI211_X1 U13689 ( .C1(n11466), .C2(n15082), .A(n11346), .B(n11345), .ZN(
        P3_U3224) );
  OAI222_X1 U13690 ( .A1(n13819), .A2(n11349), .B1(P2_U3088), .B2(n11348), 
        .C1(n13817), .C2(n11347), .ZN(P2_U3305) );
  OAI22_X1 U13691 ( .A1(n14760), .A2(n12230), .B1(n11350), .B2(n12228), .ZN(
        n11418) );
  OAI22_X1 U13692 ( .A1(n14760), .A2(n12231), .B1(n11350), .B2(n12230), .ZN(
        n11351) );
  XNOR2_X1 U13693 ( .A(n11351), .B(n12020), .ZN(n11417) );
  XOR2_X1 U13694 ( .A(n11418), .B(n11417), .Z(n11359) );
  INV_X1 U13695 ( .A(n11352), .ZN(n11355) );
  INV_X1 U13696 ( .A(n11353), .ZN(n11354) );
  NAND2_X1 U13697 ( .A1(n11358), .A2(n11359), .ZN(n11425) );
  OAI21_X1 U13698 ( .B1(n11359), .B2(n11358), .A(n11421), .ZN(n11360) );
  NAND2_X1 U13699 ( .A1(n11360), .A2(n13937), .ZN(n11367) );
  NAND2_X1 U13700 ( .A1(n13970), .A2(n14064), .ZN(n11362) );
  NAND2_X1 U13701 ( .A1(n13968), .A2(n6479), .ZN(n11361) );
  NAND2_X1 U13702 ( .A1(n11362), .A2(n11361), .ZN(n14694) );
  NOR2_X1 U13703 ( .A1(n13920), .A2(n11363), .ZN(n11364) );
  AOI211_X1 U13704 ( .C1(n13923), .C2(n14694), .A(n11365), .B(n11364), .ZN(
        n11366) );
  OAI211_X1 U13705 ( .C1(n14760), .C2(n13943), .A(n11367), .B(n11366), .ZN(
        P1_U3221) );
  AOI21_X1 U13706 ( .B1(n6478), .B2(n15017), .A(n11368), .ZN(n11371) );
  OR2_X1 U13707 ( .A1(n12652), .A2(n11369), .ZN(n11370) );
  OAI211_X1 U13708 ( .C1(n11588), .C2(n12697), .A(n11371), .B(n11370), .ZN(
        n11379) );
  XNOR2_X1 U13709 ( .A(n12567), .B(n15017), .ZN(n11504) );
  XNOR2_X1 U13710 ( .A(n11504), .B(n11509), .ZN(n11377) );
  NOR2_X1 U13711 ( .A1(n11372), .A2(n12715), .ZN(n11373) );
  OR2_X1 U13712 ( .A1(n11375), .A2(n11373), .ZN(n11376) );
  AOI211_X1 U13713 ( .C1(n11377), .C2(n11376), .A(n12689), .B(n6609), .ZN(
        n11378) );
  AOI211_X1 U13714 ( .C1(n15015), .C2(n12700), .A(n11379), .B(n11378), .ZN(
        n11380) );
  INV_X1 U13715 ( .A(n11380), .ZN(P3_U3157) );
  OAI211_X1 U13716 ( .C1(n11383), .C2(n11382), .A(n11381), .B(n13019), .ZN(
        n11385) );
  AOI22_X1 U13717 ( .A1(n13023), .A2(n12714), .B1(n12712), .B2(n13022), .ZN(
        n11384) );
  NAND2_X1 U13718 ( .A1(n11385), .A2(n11384), .ZN(n14574) );
  INV_X1 U13719 ( .A(n14574), .ZN(n11393) );
  OAI21_X1 U13720 ( .B1(n11388), .B2(n11387), .A(n11386), .ZN(n14576) );
  NOR2_X1 U13721 ( .A1(n13031), .A2(n14573), .ZN(n11391) );
  INV_X1 U13722 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11547) );
  INV_X1 U13723 ( .A(n11389), .ZN(n11591) );
  OAI22_X1 U13724 ( .A1(n15030), .A2(n11547), .B1(n11591), .B2(n15025), .ZN(
        n11390) );
  AOI211_X1 U13725 ( .C1(n14576), .C2(n13033), .A(n11391), .B(n11390), .ZN(
        n11392) );
  OAI21_X1 U13726 ( .B1(n11393), .B2(n15032), .A(n11392), .ZN(P3_U3221) );
  INV_X1 U13727 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14597) );
  AOI22_X1 U13728 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n14869), .B1(n11410), 
        .B2(n14597), .ZN(n14868) );
  MUX2_X1 U13729 ( .A(n11396), .B(P2_REG1_REG_11__SCAN_IN), .S(n14859), .Z(
        n14855) );
  OAI21_X1 U13730 ( .B1(n14869), .B2(P2_REG1_REG_12__SCAN_IN), .A(n14866), 
        .ZN(n11399) );
  NOR2_X1 U13731 ( .A1(n11412), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n11397) );
  AOI21_X1 U13732 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n11412), .A(n11397), 
        .ZN(n11398) );
  NOR2_X1 U13733 ( .A1(n11399), .A2(n11398), .ZN(n11861) );
  AOI211_X1 U13734 ( .C1(n11399), .C2(n11398), .A(n11861), .B(n14901), .ZN(
        n11403) );
  NOR2_X1 U13735 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8776), .ZN(n11400) );
  AOI21_X1 U13736 ( .B1(n14821), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n11400), 
        .ZN(n11401) );
  OAI21_X1 U13737 ( .B1(n11412), .B2(n14839), .A(n11401), .ZN(n11402) );
  NOR2_X1 U13738 ( .A1(n11403), .A2(n11402), .ZN(n11416) );
  NOR2_X1 U13739 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n14869), .ZN(n11411) );
  NOR2_X1 U13740 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n14859), .ZN(n11409) );
  INV_X1 U13741 ( .A(n11404), .ZN(n11405) );
  OAI21_X1 U13742 ( .B1(n11407), .B2(n11406), .A(n11405), .ZN(n14851) );
  AOI22_X1 U13743 ( .A1(P2_REG2_REG_11__SCAN_IN), .A2(n11408), .B1(n14859), 
        .B2(n11165), .ZN(n14850) );
  NOR2_X1 U13744 ( .A1(n14851), .A2(n14850), .ZN(n14849) );
  AOI22_X1 U13745 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n11410), .B1(n14869), 
        .B2(n11181), .ZN(n14863) );
  NOR2_X1 U13746 ( .A1(n14864), .A2(n14863), .ZN(n14862) );
  AOI22_X1 U13747 ( .A1(n11860), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n13641), 
        .B2(n11412), .ZN(n11413) );
  NAND2_X1 U13748 ( .A1(n11413), .A2(n11414), .ZN(n11851) );
  OAI211_X1 U13749 ( .C1(n11414), .C2(n11413), .A(n14910), .B(n11851), .ZN(
        n11415) );
  NAND2_X1 U13750 ( .A1(n11416), .A2(n11415), .ZN(P2_U3227) );
  INV_X1 U13751 ( .A(n12314), .ZN(n14768) );
  INV_X1 U13752 ( .A(n11417), .ZN(n11420) );
  INV_X1 U13753 ( .A(n11418), .ZN(n11419) );
  NAND2_X1 U13754 ( .A1(n11420), .A2(n11419), .ZN(n11424) );
  AND2_X1 U13755 ( .A1(n11421), .A2(n11424), .ZN(n11427) );
  AND2_X1 U13756 ( .A1(n12216), .A2(n13968), .ZN(n11422) );
  AOI21_X1 U13757 ( .B1(n12314), .B2(n12175), .A(n11422), .ZN(n11521) );
  AOI22_X1 U13758 ( .A1(n12314), .A2(n12205), .B1(n12175), .B2(n13968), .ZN(
        n11423) );
  XNOR2_X1 U13759 ( .A(n11423), .B(n12020), .ZN(n11520) );
  XOR2_X1 U13760 ( .A(n11521), .B(n11520), .Z(n11426) );
  OAI211_X1 U13761 ( .C1(n11427), .C2(n11426), .A(n13937), .B(n11525), .ZN(
        n11432) );
  OAI21_X1 U13762 ( .B1(n13949), .B2(n14766), .A(n11428), .ZN(n11429) );
  AOI21_X1 U13763 ( .B1(n11430), .B2(n13947), .A(n11429), .ZN(n11431) );
  OAI211_X1 U13764 ( .C1(n14768), .C2(n13943), .A(n11432), .B(n11431), .ZN(
        P1_U3231) );
  AOI21_X1 U13765 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n14389), .A(n11433), 
        .ZN(n11434) );
  OAI21_X1 U13766 ( .B1(n12122), .B2(n14391), .A(n11434), .ZN(P1_U3332) );
  NAND2_X1 U13767 ( .A1(n11536), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11435) );
  OAI211_X1 U13768 ( .C1(n12122), .C2(n13803), .A(n11436), .B(n11435), .ZN(
        P2_U3304) );
  INV_X1 U13769 ( .A(n14581), .ZN(n15034) );
  XNOR2_X1 U13770 ( .A(n11437), .B(n11438), .ZN(n15012) );
  NAND2_X1 U13771 ( .A1(n11440), .A2(n11439), .ZN(n11446) );
  NAND2_X1 U13772 ( .A1(n11457), .A2(n11441), .ZN(n11443) );
  AND2_X1 U13773 ( .A1(n11443), .A2(n11442), .ZN(n11444) );
  OAI211_X1 U13774 ( .C1(n11446), .C2(n11445), .A(n11444), .B(n13019), .ZN(
        n11448) );
  AOI22_X1 U13775 ( .A1(n12714), .A2(n13022), .B1(n13023), .B2(n12715), .ZN(
        n11447) );
  AND2_X1 U13776 ( .A1(n11448), .A2(n11447), .ZN(n15011) );
  OAI21_X1 U13777 ( .B1(n15034), .B2(n15012), .A(n15011), .ZN(n11454) );
  INV_X1 U13778 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n11449) );
  OAI22_X1 U13779 ( .A1(n13129), .A2(n11452), .B1(n11449), .B2(n15089), .ZN(
        n11450) );
  AOI21_X1 U13780 ( .B1(n11454), .B2(n15089), .A(n11450), .ZN(n11451) );
  INV_X1 U13781 ( .A(n11451), .ZN(P3_U3420) );
  OAI22_X1 U13782 ( .A1(n13087), .A2(n11452), .B1(n15106), .B2(n10687), .ZN(
        n11453) );
  AOI21_X1 U13783 ( .B1(n11454), .B2(n15106), .A(n11453), .ZN(n11455) );
  INV_X1 U13784 ( .A(n11455), .ZN(P3_U3469) );
  XNOR2_X1 U13785 ( .A(n11456), .B(n11458), .ZN(n15073) );
  OAI21_X1 U13786 ( .B1(n11459), .B2(n11458), .A(n11457), .ZN(n11460) );
  AOI222_X1 U13787 ( .A1(n13019), .A2(n11460), .B1(n12715), .B2(n13022), .C1(
        n7984), .C2(n13023), .ZN(n15074) );
  MUX2_X1 U13788 ( .A(n11461), .B(n15074), .S(n15030), .Z(n11465) );
  AOI22_X1 U13789 ( .A1(n15016), .A2(n11463), .B1(n15014), .B2(n11462), .ZN(
        n11464) );
  OAI211_X1 U13790 ( .C1(n11466), .C2(n15073), .A(n11465), .B(n11464), .ZN(
        P3_U3225) );
  AOI211_X1 U13791 ( .C1(n12339), .C2(n14735), .A(n11468), .B(n11467), .ZN(
        n11469) );
  OAI21_X1 U13792 ( .B1(n14363), .B2(n11470), .A(n11469), .ZN(n11472) );
  NAND2_X1 U13793 ( .A1(n11472), .A2(n14798), .ZN(n11471) );
  OAI21_X1 U13794 ( .B1(n14798), .B2(n10999), .A(n11471), .ZN(P1_U3541) );
  INV_X1 U13795 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11474) );
  NAND2_X1 U13796 ( .A1(n11472), .A2(n14748), .ZN(n11473) );
  OAI21_X1 U13797 ( .B1(n14748), .B2(n11474), .A(n11473), .ZN(P1_U3498) );
  NAND2_X1 U13798 ( .A1(n11476), .A2(n11475), .ZN(n11478) );
  OR2_X1 U13799 ( .A1(n12339), .A2(n12341), .ZN(n11477) );
  NAND2_X1 U13800 ( .A1(n11478), .A2(n11477), .ZN(n11627) );
  NAND2_X1 U13801 ( .A1(n11479), .A2(n12457), .ZN(n11481) );
  AOI22_X1 U13802 ( .A1(n11745), .A2(n12040), .B1(n12041), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11480) );
  OR2_X1 U13803 ( .A1(n12008), .A2(n12010), .ZN(n12343) );
  NAND2_X1 U13804 ( .A1(n12008), .A2(n12010), .ZN(n12333) );
  NAND2_X1 U13805 ( .A1(n12343), .A2(n12333), .ZN(n12485) );
  XNOR2_X1 U13806 ( .A(n11627), .B(n12485), .ZN(n14641) );
  AOI21_X1 U13807 ( .B1(n12008), .B2(n11482), .A(n14294), .ZN(n11484) );
  NAND2_X1 U13808 ( .A1(n11484), .A2(n11824), .ZN(n14635) );
  NAND2_X1 U13809 ( .A1(n11485), .A2(n12484), .ZN(n11487) );
  OR2_X1 U13810 ( .A1(n12339), .A2(n13964), .ZN(n11486) );
  INV_X1 U13811 ( .A(n12485), .ZN(n11490) );
  NAND2_X1 U13812 ( .A1(n11489), .A2(n11490), .ZN(n14637) );
  NAND3_X1 U13813 ( .A1(n14638), .A2(n14637), .A3(n14703), .ZN(n11501) );
  NAND2_X1 U13814 ( .A1(n12440), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11496) );
  OR2_X1 U13815 ( .A1(n11491), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n11492) );
  AND2_X1 U13816 ( .A1(n11634), .A2(n11492), .ZN(n13946) );
  NAND2_X1 U13817 ( .A1(n9937), .A2(n13946), .ZN(n11495) );
  NAND2_X1 U13818 ( .A1(n12441), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11494) );
  NAND2_X1 U13819 ( .A1(n12439), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11493) );
  AND4_X1 U13820 ( .A1(n11496), .A2(n11495), .A3(n11494), .A4(n11493), .ZN(
        n11631) );
  INV_X1 U13821 ( .A(n11631), .ZN(n13962) );
  AOI22_X1 U13822 ( .A1(n13962), .A2(n6479), .B1(n14064), .B2(n13964), .ZN(
        n14634) );
  OAI22_X1 U13823 ( .A1(n14634), .A2(n14724), .B1(n11497), .B2(n14252), .ZN(
        n11499) );
  INV_X1 U13824 ( .A(n12008), .ZN(n14636) );
  NOR2_X1 U13825 ( .A1(n14636), .A2(n14258), .ZN(n11498) );
  AOI211_X1 U13826 ( .C1(n14724), .C2(P1_REG2_REG_14__SCAN_IN), .A(n11499), 
        .B(n11498), .ZN(n11500) );
  OAI211_X1 U13827 ( .C1(n14635), .C2(n14270), .A(n11501), .B(n11500), .ZN(
        n11502) );
  AOI21_X1 U13828 ( .B1(n14284), .B2(n14641), .A(n11502), .ZN(n11503) );
  INV_X1 U13829 ( .A(n11503), .ZN(P1_U3279) );
  INV_X1 U13830 ( .A(n11504), .ZN(n11506) );
  NAND2_X1 U13831 ( .A1(n11506), .A2(n11505), .ZN(n11507) );
  XNOR2_X1 U13832 ( .A(n14577), .B(n12567), .ZN(n11583) );
  INV_X1 U13833 ( .A(n11583), .ZN(n11508) );
  XNOR2_X1 U13834 ( .A(n11581), .B(n12714), .ZN(n11519) );
  OR2_X1 U13835 ( .A1(n12652), .A2(n11509), .ZN(n11515) );
  OR2_X1 U13836 ( .A1(n12697), .A2(n11700), .ZN(n11514) );
  NAND2_X1 U13837 ( .A1(n12674), .A2(n11510), .ZN(n11513) );
  INV_X1 U13838 ( .A(n11511), .ZN(n11512) );
  NAND4_X1 U13839 ( .A1(n11515), .A2(n11514), .A3(n11513), .A4(n11512), .ZN(
        n11516) );
  AOI21_X1 U13840 ( .B1(n12700), .B2(n11517), .A(n11516), .ZN(n11518) );
  OAI21_X1 U13841 ( .B1(n11519), .B2(n12689), .A(n11518), .ZN(P3_U3176) );
  INV_X1 U13842 ( .A(n11520), .ZN(n11523) );
  AND2_X1 U13843 ( .A1(n12216), .A2(n13967), .ZN(n11526) );
  AOI21_X1 U13844 ( .B1(n14778), .B2(n12175), .A(n11526), .ZN(n11717) );
  AOI22_X1 U13845 ( .A1(n14778), .A2(n12205), .B1(n12175), .B2(n13967), .ZN(
        n11527) );
  XNOR2_X1 U13846 ( .A(n11527), .B(n12020), .ZN(n11716) );
  XOR2_X1 U13847 ( .A(n11717), .B(n11716), .Z(n11720) );
  XNOR2_X1 U13848 ( .A(n11721), .B(n11720), .ZN(n11535) );
  AOI21_X1 U13849 ( .B1(n11529), .B2(n11528), .A(n13949), .ZN(n11530) );
  AOI211_X1 U13850 ( .C1(n11532), .C2(n13947), .A(n11531), .B(n11530), .ZN(
        n11534) );
  NAND2_X1 U13851 ( .A1(n14778), .A2(n13952), .ZN(n11533) );
  OAI211_X1 U13852 ( .C1(n11535), .C2(n13955), .A(n11534), .B(n11533), .ZN(
        P1_U3217) );
  AOI22_X1 U13853 ( .A1(n11537), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n11536), .ZN(n11538) );
  OAI21_X1 U13854 ( .B1(n12142), .B2(n13803), .A(n11538), .ZN(P2_U3303) );
  NOR2_X1 U13855 ( .A1(n11552), .A2(n11539), .ZN(n11541) );
  INV_X1 U13856 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n11554) );
  MUX2_X1 U13857 ( .A(n11554), .B(P3_REG1_REG_12__SCAN_IN), .S(n11921), .Z(
        n11542) );
  AOI21_X1 U13858 ( .B1(n11543), .B2(n11542), .A(n11916), .ZN(n11564) );
  NOR2_X1 U13859 ( .A1(n11552), .A2(n11544), .ZN(n11546) );
  INV_X1 U13860 ( .A(n11921), .ZN(n11927) );
  AOI22_X1 U13861 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11927), .B1(n11921), 
        .B2(n11547), .ZN(n11548) );
  AOI21_X1 U13862 ( .B1(n11549), .B2(n11548), .A(n11920), .ZN(n11561) );
  AND2_X1 U13863 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n11587) );
  NOR2_X1 U13864 ( .A1(n14994), .A2(n11921), .ZN(n11550) );
  AOI211_X1 U13865 ( .C1(n14987), .C2(P3_ADDR_REG_12__SCAN_IN), .A(n11587), 
        .B(n11550), .ZN(n11560) );
  INV_X1 U13866 ( .A(n11551), .ZN(n11553) );
  NAND2_X1 U13867 ( .A1(n11553), .A2(n11552), .ZN(n11555) );
  AND2_X1 U13868 ( .A1(n11556), .A2(n11555), .ZN(n11558) );
  MUX2_X1 U13869 ( .A(n11547), .B(n11554), .S(n13141), .Z(n11926) );
  XNOR2_X1 U13870 ( .A(n11926), .B(n11921), .ZN(n11557) );
  NAND3_X1 U13871 ( .A1(n11556), .A2(n11555), .A3(n11557), .ZN(n11925) );
  OAI211_X1 U13872 ( .C1(n11558), .C2(n11557), .A(n12778), .B(n11925), .ZN(
        n11559) );
  OAI211_X1 U13873 ( .C1(n11561), .C2(n15008), .A(n11560), .B(n11559), .ZN(
        n11562) );
  INV_X1 U13874 ( .A(n11562), .ZN(n11563) );
  OAI21_X1 U13875 ( .B1(n11564), .B2(n15002), .A(n11563), .ZN(P3_U3194) );
  XOR2_X1 U13876 ( .A(n11657), .B(n11651), .Z(n13638) );
  NAND2_X1 U13877 ( .A1(n11567), .A2(n13644), .ZN(n11568) );
  NAND2_X1 U13878 ( .A1(n11568), .A2(n13521), .ZN(n11569) );
  NOR2_X1 U13879 ( .A1(n11658), .A2(n11569), .ZN(n13647) );
  OR2_X1 U13880 ( .A1(n14813), .A2(n11621), .ZN(n11570) );
  NAND2_X1 U13881 ( .A1(n11571), .A2(n11570), .ZN(n11652) );
  XNOR2_X1 U13882 ( .A(n11652), .B(n11651), .ZN(n11572) );
  OAI222_X1 U13883 ( .A1(n13631), .A2(n11787), .B1(n13575), .B2(n11621), .C1(
        n11572), .C2(n13603), .ZN(n13645) );
  AOI211_X1 U13884 ( .C1(n13638), .C2(n14951), .A(n13647), .B(n13645), .ZN(
        n11576) );
  AOI22_X1 U13885 ( .A1(n13644), .A2(n11672), .B1(n14984), .B2(
        P2_REG1_REG_13__SCAN_IN), .ZN(n11573) );
  OAI21_X1 U13886 ( .B1(n11576), .B2(n14984), .A(n11573), .ZN(P2_U3512) );
  OAI22_X1 U13887 ( .A1(n6771), .A2(n13794), .B1(n14974), .B2(n8780), .ZN(
        n11574) );
  INV_X1 U13888 ( .A(n11574), .ZN(n11575) );
  OAI21_X1 U13889 ( .B1(n11576), .B2(n14973), .A(n11575), .ZN(P2_U3469) );
  INV_X1 U13890 ( .A(n11577), .ZN(n11578) );
  OAI222_X1 U13891 ( .A1(n13143), .A2(n11580), .B1(P3_U3151), .B2(n11579), 
        .C1(n6484), .C2(n11578), .ZN(P3_U3270) );
  NAND2_X1 U13892 ( .A1(n11581), .A2(n12714), .ZN(n11585) );
  NAND2_X1 U13893 ( .A1(n11582), .A2(n11583), .ZN(n11584) );
  XOR2_X1 U13894 ( .A(n12567), .B(n14573), .Z(n11701) );
  XNOR2_X1 U13895 ( .A(n11701), .B(n12713), .ZN(n11586) );
  XNOR2_X1 U13896 ( .A(n11704), .B(n11586), .ZN(n11595) );
  INV_X1 U13897 ( .A(n14573), .ZN(n11593) );
  AOI21_X1 U13898 ( .B1(n12649), .B2(n12712), .A(n11587), .ZN(n11590) );
  OR2_X1 U13899 ( .A1(n12652), .A2(n11588), .ZN(n11589) );
  OAI211_X1 U13900 ( .C1(n12672), .C2(n11591), .A(n11590), .B(n11589), .ZN(
        n11592) );
  AOI21_X1 U13901 ( .B1(n11593), .B2(n6478), .A(n11592), .ZN(n11594) );
  OAI21_X1 U13902 ( .B1(n11595), .B2(n12689), .A(n11594), .ZN(P3_U3164) );
  INV_X1 U13903 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12143) );
  OAI222_X1 U13904 ( .A1(n11596), .A2(P1_U3086), .B1(n14391), .B2(n12142), 
        .C1(n12143), .C2(n14396), .ZN(P1_U3331) );
  XNOR2_X1 U13905 ( .A(n11597), .B(n11598), .ZN(n11599) );
  OAI222_X1 U13906 ( .A1(n12964), .A2(n11700), .B1(n12962), .B2(n12526), .C1(
        n11599), .C2(n12960), .ZN(n14570) );
  INV_X1 U13907 ( .A(n14570), .ZN(n11605) );
  XNOR2_X1 U13908 ( .A(n11601), .B(n11600), .ZN(n14572) );
  AOI22_X1 U13909 ( .A1(n15032), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15014), 
        .B2(n11706), .ZN(n11602) );
  OAI21_X1 U13910 ( .B1(n14569), .B2(n13031), .A(n11602), .ZN(n11603) );
  AOI21_X1 U13911 ( .B1(n14572), .B2(n13033), .A(n11603), .ZN(n11604) );
  OAI21_X1 U13912 ( .B1(n11605), .B2(n15032), .A(n11604), .ZN(P3_U3220) );
  XNOR2_X1 U13913 ( .A(n13644), .B(n13222), .ZN(n11688) );
  AND2_X1 U13914 ( .A1(n13347), .A2(n13221), .ZN(n11606) );
  NAND2_X1 U13915 ( .A1(n11688), .A2(n11606), .ZN(n11685) );
  INV_X1 U13916 ( .A(n11688), .ZN(n11608) );
  INV_X1 U13917 ( .A(n11606), .ZN(n11607) );
  NAND2_X1 U13918 ( .A1(n11608), .A2(n11607), .ZN(n11609) );
  AND2_X1 U13919 ( .A1(n11685), .A2(n11609), .ZN(n11620) );
  INV_X1 U13920 ( .A(n11610), .ZN(n11612) );
  NAND2_X1 U13921 ( .A1(n11612), .A2(n11611), .ZN(n11613) );
  XNOR2_X1 U13922 ( .A(n14813), .B(n13178), .ZN(n11615) );
  NAND2_X1 U13923 ( .A1(n13348), .A2(n13221), .ZN(n11616) );
  AND2_X1 U13924 ( .A1(n11615), .A2(n11616), .ZN(n14809) );
  INV_X1 U13925 ( .A(n11615), .ZN(n11618) );
  INV_X1 U13926 ( .A(n11616), .ZN(n11617) );
  NAND2_X1 U13927 ( .A1(n11618), .A2(n11617), .ZN(n14805) );
  OAI211_X1 U13928 ( .C1(n11620), .C2(n11619), .A(n11687), .B(n13276), .ZN(
        n11625) );
  OAI22_X1 U13929 ( .A1(n14800), .A2(n11787), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8776), .ZN(n11623) );
  OAI22_X1 U13930 ( .A1(n14801), .A2(n11621), .B1(n13640), .B2(n14816), .ZN(
        n11622) );
  AOI211_X1 U13931 ( .C1(n13644), .C2(n14812), .A(n11623), .B(n11622), .ZN(
        n11624) );
  NAND2_X1 U13932 ( .A1(n11625), .A2(n11624), .ZN(P2_U3206) );
  INV_X1 U13933 ( .A(n12343), .ZN(n11626) );
  NAND2_X1 U13934 ( .A1(n11628), .A2(n12457), .ZN(n11630) );
  AOI22_X1 U13935 ( .A1(n14682), .A2(n12040), .B1(n12041), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n11629) );
  NAND2_X1 U13936 ( .A1(n13953), .A2(n11631), .ZN(n12349) );
  NAND2_X1 U13937 ( .A1(n12344), .A2(n12349), .ZN(n12486) );
  AOI21_X1 U13938 ( .B1(n11632), .B2(n12486), .A(n14710), .ZN(n11643) );
  OR2_X1 U13939 ( .A1(n12010), .A2(n13917), .ZN(n11641) );
  INV_X1 U13940 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n11633) );
  NAND2_X1 U13941 ( .A1(n11634), .A2(n11633), .ZN(n11635) );
  NAND2_X1 U13942 ( .A1(n11810), .A2(n11635), .ZN(n14604) );
  NAND2_X1 U13943 ( .A1(n12441), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11637) );
  NAND2_X1 U13944 ( .A1(n12439), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11636) );
  AND2_X1 U13945 ( .A1(n11637), .A2(n11636), .ZN(n11639) );
  NAND2_X1 U13946 ( .A1(n12440), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11638) );
  OAI211_X1 U13947 ( .C1(n14604), .C2(n12092), .A(n11639), .B(n11638), .ZN(
        n13961) );
  NAND2_X1 U13948 ( .A1(n13961), .A2(n6479), .ZN(n11640) );
  AND2_X1 U13949 ( .A1(n11641), .A2(n11640), .ZN(n13950) );
  INV_X1 U13950 ( .A(n13950), .ZN(n11642) );
  AOI21_X1 U13951 ( .B1(n11643), .B2(n11801), .A(n11642), .ZN(n14630) );
  INV_X1 U13952 ( .A(n12010), .ZN(n13963) );
  NAND2_X1 U13953 ( .A1(n12008), .A2(n13963), .ZN(n11644) );
  OAI21_X1 U13954 ( .B1(n6603), .B2(n12486), .A(n11821), .ZN(n14633) );
  NAND2_X1 U13955 ( .A1(n14633), .A2(n14703), .ZN(n11650) );
  XOR2_X1 U13956 ( .A(n11824), .B(n13953), .Z(n11645) );
  NAND2_X1 U13957 ( .A1(n11645), .A2(n14749), .ZN(n14629) );
  INV_X1 U13958 ( .A(n14629), .ZN(n11648) );
  INV_X1 U13959 ( .A(n13953), .ZN(n14631) );
  AOI22_X1 U13960 ( .A1(n14724), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13946), 
        .B2(n14713), .ZN(n11646) );
  OAI21_X1 U13961 ( .B1(n14631), .B2(n14258), .A(n11646), .ZN(n11647) );
  AOI21_X1 U13962 ( .B1(n11648), .B2(n14720), .A(n11647), .ZN(n11649) );
  OAI211_X1 U13963 ( .C1(n14724), .C2(n14630), .A(n11650), .B(n11649), .ZN(
        P1_U3278) );
  NAND2_X1 U13964 ( .A1(n11652), .A2(n11651), .ZN(n11654) );
  OR2_X1 U13965 ( .A1(n13644), .A2(n14799), .ZN(n11653) );
  XNOR2_X1 U13966 ( .A(n11784), .B(n11789), .ZN(n11655) );
  AOI22_X1 U13967 ( .A1(n13466), .A2(n13629), .B1(n13347), .B2(n13628), .ZN(
        n11694) );
  OAI21_X1 U13968 ( .B1(n11655), .B2(n13603), .A(n11694), .ZN(n11666) );
  INV_X1 U13969 ( .A(n11666), .ZN(n11665) );
  XOR2_X1 U13970 ( .A(n11789), .B(n11790), .Z(n11668) );
  NAND2_X1 U13971 ( .A1(n11668), .A2(n13656), .ZN(n11664) );
  INV_X1 U13972 ( .A(n11793), .ZN(n11659) );
  AOI211_X1 U13973 ( .C1(n11697), .C2(n6773), .A(n13221), .B(n11659), .ZN(
        n11667) );
  NOR2_X1 U13974 ( .A1(n11788), .A2(n13589), .ZN(n11662) );
  OAI22_X1 U13975 ( .A1(n13642), .A2(n11660), .B1(n11693), .B2(n13639), .ZN(
        n11661) );
  AOI211_X1 U13976 ( .C1(n11667), .C2(n13646), .A(n11662), .B(n11661), .ZN(
        n11663) );
  OAI211_X1 U13977 ( .C1(n13595), .C2(n11665), .A(n11664), .B(n11663), .ZN(
        P2_U3251) );
  AOI211_X1 U13978 ( .C1(n11668), .C2(n14951), .A(n11667), .B(n11666), .ZN(
        n11674) );
  INV_X1 U13979 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11669) );
  OAI22_X1 U13980 ( .A1(n11788), .A2(n13794), .B1(n14974), .B2(n11669), .ZN(
        n11670) );
  INV_X1 U13981 ( .A(n11670), .ZN(n11671) );
  OAI21_X1 U13982 ( .B1(n11674), .B2(n14973), .A(n11671), .ZN(P2_U3472) );
  AOI22_X1 U13983 ( .A1(n11697), .A2(n11672), .B1(n14984), .B2(
        P2_REG1_REG_14__SCAN_IN), .ZN(n11673) );
  OAI21_X1 U13984 ( .B1(n11674), .B2(n14984), .A(n11673), .ZN(P2_U3513) );
  XNOR2_X1 U13985 ( .A(n11675), .B(n11678), .ZN(n11676) );
  OAI222_X1 U13986 ( .A1(n12962), .A2(n12625), .B1(n12964), .B2(n11677), .C1(
        n11676), .C2(n12960), .ZN(n11831) );
  INV_X1 U13987 ( .A(n11831), .ZN(n11684) );
  OAI21_X1 U13988 ( .B1(n11680), .B2(n7729), .A(n11679), .ZN(n11832) );
  AOI22_X1 U13989 ( .A1(n15032), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15014), 
        .B2(n11875), .ZN(n11681) );
  OAI21_X1 U13990 ( .B1(n11874), .B2(n13031), .A(n11681), .ZN(n11682) );
  AOI21_X1 U13991 ( .B1(n11832), .B2(n13033), .A(n11682), .ZN(n11683) );
  OAI21_X1 U13992 ( .B1(n11684), .B2(n15032), .A(n11683), .ZN(P3_U3219) );
  XNOR2_X1 U13993 ( .A(n11788), .B(n13222), .ZN(n11894) );
  NOR2_X1 U13994 ( .A1(n11787), .A2(n13521), .ZN(n11892) );
  XNOR2_X1 U13995 ( .A(n11894), .B(n11892), .ZN(n11690) );
  NAND3_X1 U13996 ( .A1(n11688), .A2(n13306), .A3(n13347), .ZN(n11689) );
  OAI21_X1 U13997 ( .B1(n11687), .B2(n14808), .A(n11689), .ZN(n11692) );
  INV_X1 U13998 ( .A(n11690), .ZN(n11691) );
  NAND2_X1 U13999 ( .A1(n11692), .A2(n11691), .ZN(n11699) );
  NOR2_X1 U14000 ( .A1(n14816), .A2(n11693), .ZN(n11696) );
  OAI22_X1 U14001 ( .A1(n13282), .A2(n11694), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14875), .ZN(n11695) );
  AOI211_X1 U14002 ( .C1(n11697), .C2(n14812), .A(n11696), .B(n11695), .ZN(
        n11698) );
  OAI211_X1 U14003 ( .C1(n11896), .C2(n14808), .A(n11699), .B(n11698), .ZN(
        P2_U3187) );
  NOR2_X1 U14004 ( .A1(n11701), .A2(n11700), .ZN(n11703) );
  NAND2_X1 U14005 ( .A1(n11701), .A2(n11700), .ZN(n11702) );
  XNOR2_X1 U14006 ( .A(n14569), .B(n12567), .ZN(n11872) );
  XNOR2_X1 U14007 ( .A(n11872), .B(n12712), .ZN(n11705) );
  XNOR2_X1 U14008 ( .A(n6622), .B(n11705), .ZN(n11713) );
  NAND2_X1 U14009 ( .A1(n12700), .A2(n11706), .ZN(n11709) );
  INV_X1 U14010 ( .A(n12652), .ZN(n12695) );
  NOR2_X1 U14011 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11707), .ZN(n15006) );
  AOI21_X1 U14012 ( .B1(n12695), .B2(n12713), .A(n15006), .ZN(n11708) );
  OAI211_X1 U14013 ( .C1(n12526), .C2(n12697), .A(n11709), .B(n11708), .ZN(
        n11710) );
  AOI21_X1 U14014 ( .B1(n11711), .B2(n12674), .A(n11710), .ZN(n11712) );
  OAI21_X1 U14015 ( .B1(n11713), .B2(n12689), .A(n11712), .ZN(P3_U3174) );
  OAI22_X1 U14016 ( .A1(n14643), .A2(n12230), .B1(n11714), .B2(n12228), .ZN(
        n11765) );
  OAI22_X1 U14017 ( .A1(n14643), .A2(n12231), .B1(n11714), .B2(n12230), .ZN(
        n11715) );
  XNOR2_X1 U14018 ( .A(n11715), .B(n12020), .ZN(n11764) );
  XOR2_X1 U14019 ( .A(n11765), .B(n11764), .Z(n11722) );
  INV_X1 U14020 ( .A(n11716), .ZN(n11719) );
  INV_X1 U14021 ( .A(n11717), .ZN(n11718) );
  OAI21_X1 U14022 ( .B1(n11722), .B2(n6604), .A(n11773), .ZN(n11723) );
  NAND2_X1 U14023 ( .A1(n11723), .A2(n13937), .ZN(n11729) );
  OAI21_X1 U14024 ( .B1(n13949), .B2(n11725), .A(n11724), .ZN(n11726) );
  AOI21_X1 U14025 ( .B1(n11727), .B2(n13947), .A(n11726), .ZN(n11728) );
  OAI211_X1 U14026 ( .C1(n14643), .C2(n13943), .A(n11729), .B(n11728), .ZN(
        P1_U3236) );
  INV_X1 U14027 ( .A(n12162), .ZN(n11733) );
  OAI222_X1 U14028 ( .A1(n13819), .A2(n11731), .B1(n13803), .B2(n11733), .C1(
        n11730), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U14029 ( .A(n11732), .ZN(n11734) );
  OAI222_X1 U14030 ( .A1(P1_U3086), .A2(n11734), .B1(n14391), .B2(n11733), 
        .C1(n15118), .C2(n14396), .ZN(P1_U3330) );
  INV_X1 U14031 ( .A(n14023), .ZN(n14683) );
  INV_X1 U14032 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n11735) );
  NAND2_X1 U14033 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13876)
         );
  OAI21_X1 U14034 ( .B1(n14691), .B2(n11735), .A(n13876), .ZN(n11744) );
  NAND2_X1 U14035 ( .A1(n11738), .A2(n11737), .ZN(n11739) );
  INV_X1 U14036 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14678) );
  NAND2_X1 U14037 ( .A1(n14679), .A2(n14678), .ZN(n14677) );
  NAND2_X1 U14038 ( .A1(n11739), .A2(n14677), .ZN(n11742) );
  INV_X1 U14039 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n11740) );
  MUX2_X1 U14040 ( .A(n11740), .B(P1_REG1_REG_16__SCAN_IN), .S(n13989), .Z(
        n11741) );
  NOR2_X1 U14041 ( .A1(n11741), .A2(n11742), .ZN(n13978) );
  AOI211_X1 U14042 ( .C1(n11742), .C2(n11741), .A(n13978), .B(n13980), .ZN(
        n11743) );
  AOI211_X1 U14043 ( .C1(n14683), .C2(n13989), .A(n11744), .B(n11743), .ZN(
        n11754) );
  NAND2_X1 U14044 ( .A1(n11745), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11747) );
  NAND2_X1 U14045 ( .A1(n11747), .A2(n11746), .ZN(n11748) );
  NOR2_X1 U14046 ( .A1(n14682), .A2(n11748), .ZN(n11749) );
  XNOR2_X1 U14047 ( .A(n14682), .B(n11748), .ZN(n14676) );
  NOR2_X1 U14048 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14676), .ZN(n14675) );
  NOR2_X1 U14049 ( .A1(n11749), .A2(n14675), .ZN(n11752) );
  INV_X1 U14050 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11750) );
  MUX2_X1 U14051 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n11750), .S(n13989), .Z(
        n11751) );
  NAND2_X1 U14052 ( .A1(n11751), .A2(n11752), .ZN(n13990) );
  OAI211_X1 U14053 ( .C1(n11752), .C2(n11751), .A(n14027), .B(n13990), .ZN(
        n11753) );
  NAND2_X1 U14054 ( .A1(n11754), .A2(n11753), .ZN(P1_U3259) );
  XNOR2_X1 U14055 ( .A(n11756), .B(n11755), .ZN(n11757) );
  OAI222_X1 U14056 ( .A1(n12962), .A2(n12698), .B1(n12964), .B2(n12526), .C1(
        n11757), .C2(n12960), .ZN(n11910) );
  INV_X1 U14057 ( .A(n11910), .ZN(n11763) );
  XNOR2_X1 U14058 ( .A(n11759), .B(n11758), .ZN(n11911) );
  INV_X1 U14059 ( .A(n12529), .ZN(n12705) );
  AOI22_X1 U14060 ( .A1(n15032), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15014), 
        .B2(n12701), .ZN(n11760) );
  OAI21_X1 U14061 ( .B1(n12705), .B2(n13031), .A(n11760), .ZN(n11761) );
  AOI21_X1 U14062 ( .B1(n11911), .B2(n13033), .A(n11761), .ZN(n11762) );
  OAI21_X1 U14063 ( .B1(n11763), .B2(n15032), .A(n11762), .ZN(P3_U3218) );
  INV_X1 U14064 ( .A(n11764), .ZN(n11767) );
  INV_X1 U14065 ( .A(n11765), .ZN(n11766) );
  NAND2_X1 U14066 ( .A1(n11767), .A2(n11766), .ZN(n11772) );
  AND2_X1 U14067 ( .A1(n11773), .A2(n11772), .ZN(n11775) );
  NAND2_X1 U14068 ( .A1(n12329), .A2(n12205), .ZN(n11769) );
  NAND2_X1 U14069 ( .A1(n13965), .A2(n12175), .ZN(n11768) );
  NAND2_X1 U14070 ( .A1(n11769), .A2(n11768), .ZN(n11770) );
  XNOR2_X1 U14071 ( .A(n11770), .B(n12020), .ZN(n11838) );
  AND2_X1 U14072 ( .A1(n12216), .A2(n13965), .ZN(n11771) );
  AOI21_X1 U14073 ( .B1(n12329), .B2(n12175), .A(n11771), .ZN(n11839) );
  XNOR2_X1 U14074 ( .A(n11838), .B(n11839), .ZN(n11774) );
  NAND3_X1 U14075 ( .A1(n11773), .A2(n11774), .A3(n11772), .ZN(n11841) );
  OAI211_X1 U14076 ( .C1(n11775), .C2(n11774), .A(n13937), .B(n11841), .ZN(
        n11781) );
  OAI21_X1 U14077 ( .B1(n13949), .B2(n11777), .A(n11776), .ZN(n11778) );
  AOI21_X1 U14078 ( .B1(n11779), .B2(n13947), .A(n11778), .ZN(n11780) );
  OAI211_X1 U14079 ( .C1(n11782), .C2(n13943), .A(n11781), .B(n11780), .ZN(
        P1_U3224) );
  AND2_X1 U14080 ( .A1(n11788), .A2(n13346), .ZN(n11783) );
  XNOR2_X1 U14081 ( .A(n11948), .B(n11792), .ZN(n11786) );
  NAND2_X1 U14082 ( .A1(n13345), .A2(n13466), .ZN(n11785) );
  OAI21_X1 U14083 ( .B1(n11787), .B2(n13575), .A(n11785), .ZN(n11899) );
  AOI21_X1 U14084 ( .B1(n11786), .B2(n13625), .A(n11899), .ZN(n13750) );
  AOI21_X1 U14085 ( .B1(n11792), .B2(n11791), .A(n11977), .ZN(n13752) );
  INV_X1 U14086 ( .A(n13752), .ZN(n11799) );
  AOI21_X1 U14087 ( .B1(n11976), .B2(n11793), .A(n9793), .ZN(n11794) );
  INV_X1 U14088 ( .A(n11993), .ZN(n13619) );
  NAND2_X1 U14089 ( .A1(n11794), .A2(n13619), .ZN(n13749) );
  OAI22_X1 U14090 ( .A1(n13642), .A2(n11795), .B1(n11901), .B2(n13639), .ZN(
        n11796) );
  AOI21_X1 U14091 ( .B1(n11976), .B2(n13655), .A(n11796), .ZN(n11797) );
  OAI21_X1 U14092 ( .B1(n13749), .B2(n13659), .A(n11797), .ZN(n11798) );
  AOI21_X1 U14093 ( .B1(n11799), .B2(n13656), .A(n11798), .ZN(n11800) );
  OAI21_X1 U14094 ( .B1(n13595), .B2(n13750), .A(n11800), .ZN(P2_U3250) );
  NAND2_X1 U14095 ( .A1(n11802), .A2(n12457), .ZN(n11804) );
  AOI22_X1 U14096 ( .A1(n12041), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12040), 
        .B2(n13989), .ZN(n11803) );
  XNOR2_X1 U14097 ( .A(n14607), .B(n13961), .ZN(n12487) );
  INV_X1 U14098 ( .A(n13961), .ZN(n12352) );
  NAND2_X1 U14099 ( .A1(n14607), .A2(n12352), .ZN(n11805) );
  NAND2_X1 U14100 ( .A1(n14610), .A2(n11805), .ZN(n14050) );
  NAND2_X1 U14101 ( .A1(n11806), .A2(n12457), .ZN(n11808) );
  AOI22_X1 U14102 ( .A1(n12041), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n12040), 
        .B2(n14004), .ZN(n11807) );
  INV_X1 U14103 ( .A(n14619), .ZN(n12366) );
  INV_X1 U14104 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11809) );
  AND2_X1 U14105 ( .A1(n11810), .A2(n11809), .ZN(n11811) );
  OR2_X1 U14106 ( .A1(n11811), .A2(n11814), .ZN(n13886) );
  AOI22_X1 U14107 ( .A1(n12439), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n12440), 
        .B2(P1_REG2_REG_17__SCAN_IN), .ZN(n11813) );
  NAND2_X1 U14108 ( .A1(n12441), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11812) );
  OAI211_X1 U14109 ( .C1(n13886), .C2(n12092), .A(n11813), .B(n11812), .ZN(
        n14047) );
  XNOR2_X1 U14110 ( .A(n12366), .B(n14047), .ZN(n12488) );
  XNOR2_X1 U14111 ( .A(n14050), .B(n14049), .ZN(n11820) );
  NAND2_X1 U14112 ( .A1(n11814), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n12045) );
  OR2_X1 U14113 ( .A1(n11814), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11815) );
  AND2_X1 U14114 ( .A1(n12045), .A2(n11815), .ZN(n14266) );
  NAND2_X1 U14115 ( .A1(n14266), .A2(n9937), .ZN(n11818) );
  AOI22_X1 U14116 ( .A1(n12439), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n12223), 
        .B2(P1_REG2_REG_18__SCAN_IN), .ZN(n11817) );
  NAND2_X1 U14117 ( .A1(n12441), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11816) );
  AND3_X1 U14118 ( .A1(n11818), .A2(n11817), .A3(n11816), .ZN(n13851) );
  OAI22_X1 U14119 ( .A1(n13851), .A2(n13916), .B1(n12352), .B2(n13917), .ZN(
        n13888) );
  INV_X1 U14120 ( .A(n13888), .ZN(n11819) );
  OAI21_X1 U14121 ( .B1(n11820), .B2(n14710), .A(n11819), .ZN(n14620) );
  INV_X1 U14122 ( .A(n14620), .ZN(n11830) );
  NAND2_X1 U14123 ( .A1(n14599), .A2(n14613), .ZN(n11823) );
  OR2_X1 U14124 ( .A1(n14607), .A2(n13961), .ZN(n11822) );
  XNOR2_X1 U14125 ( .A(n14069), .B(n14049), .ZN(n14622) );
  OR2_X1 U14126 ( .A1(n13953), .A2(n11824), .ZN(n14600) );
  AND2_X1 U14127 ( .A1(n14601), .A2(n14619), .ZN(n14265) );
  NOR2_X1 U14128 ( .A1(n14619), .A2(n14601), .ZN(n11825) );
  OR3_X1 U14129 ( .A1(n14265), .A2(n11825), .A3(n14294), .ZN(n14618) );
  INV_X1 U14130 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13987) );
  OAI22_X1 U14131 ( .A1(n14282), .A2(n13987), .B1(n13886), .B2(n14252), .ZN(
        n11826) );
  AOI21_X1 U14132 ( .B1(n12366), .B2(n14715), .A(n11826), .ZN(n11827) );
  OAI21_X1 U14133 ( .B1(n14618), .B2(n14270), .A(n11827), .ZN(n11828) );
  AOI21_X1 U14134 ( .B1(n14622), .B2(n14703), .A(n11828), .ZN(n11829) );
  OAI21_X1 U14135 ( .B1(n11830), .B2(n14724), .A(n11829), .ZN(P1_U3276) );
  INV_X1 U14136 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n11833) );
  AOI21_X1 U14137 ( .B1(n14581), .B2(n11832), .A(n11831), .ZN(n11835) );
  MUX2_X1 U14138 ( .A(n11833), .B(n11835), .S(n15106), .Z(n11834) );
  OAI21_X1 U14139 ( .B1(n11874), .B2(n13087), .A(n11834), .ZN(P3_U3473) );
  INV_X1 U14140 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n11836) );
  MUX2_X1 U14141 ( .A(n11836), .B(n11835), .S(n15089), .Z(n11837) );
  OAI21_X1 U14142 ( .B1(n11874), .B2(n13129), .A(n11837), .ZN(P3_U3432) );
  INV_X1 U14143 ( .A(n11838), .ZN(n11840) );
  NAND2_X1 U14144 ( .A1(n11841), .A2(n7440), .ZN(n12007) );
  AND2_X1 U14145 ( .A1(n12216), .A2(n13964), .ZN(n11842) );
  AOI21_X1 U14146 ( .B1(n12339), .B2(n12175), .A(n11842), .ZN(n12003) );
  AOI22_X1 U14147 ( .A1(n12339), .A2(n12205), .B1(n12175), .B2(n13964), .ZN(
        n11843) );
  XNOR2_X1 U14148 ( .A(n11843), .B(n12020), .ZN(n12002) );
  XOR2_X1 U14149 ( .A(n12003), .B(n12002), .Z(n12006) );
  XNOR2_X1 U14150 ( .A(n12007), .B(n12006), .ZN(n11850) );
  NAND2_X1 U14151 ( .A1(n13947), .A2(n11844), .ZN(n11846) );
  OAI211_X1 U14152 ( .C1(n11847), .C2(n13949), .A(n11846), .B(n11845), .ZN(
        n11848) );
  AOI21_X1 U14153 ( .B1(n12339), .B2(n13952), .A(n11848), .ZN(n11849) );
  OAI21_X1 U14154 ( .B1(n11850), .B2(n13955), .A(n11849), .ZN(P1_U3234) );
  INV_X1 U14155 ( .A(n11851), .ZN(n11852) );
  OR2_X1 U14156 ( .A1(n11853), .A2(n11854), .ZN(n11855) );
  XNOR2_X1 U14157 ( .A(n11854), .B(n14882), .ZN(n14884) );
  NAND2_X1 U14158 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n14884), .ZN(n14883) );
  NAND2_X1 U14159 ( .A1(n11855), .A2(n14883), .ZN(n13363) );
  XNOR2_X1 U14160 ( .A(n13375), .B(n13363), .ZN(n11856) );
  NAND2_X1 U14161 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n11856), .ZN(n13365) );
  OAI211_X1 U14162 ( .C1(n11856), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14910), 
        .B(n13365), .ZN(n11870) );
  OR2_X1 U14163 ( .A1(n14882), .A2(n11857), .ZN(n11859) );
  NAND2_X1 U14164 ( .A1(n14882), .A2(n11857), .ZN(n11858) );
  NAND2_X1 U14165 ( .A1(n11859), .A2(n11858), .ZN(n14878) );
  NAND2_X1 U14166 ( .A1(n14882), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n11862) );
  XNOR2_X1 U14167 ( .A(n13376), .B(n13375), .ZN(n11863) );
  NOR2_X1 U14168 ( .A1(n15131), .A2(n11863), .ZN(n13377) );
  AOI211_X1 U14169 ( .C1(n11863), .C2(n15131), .A(n13377), .B(n14901), .ZN(
        n11868) );
  NOR2_X1 U14170 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11864), .ZN(n11865) );
  AOI21_X1 U14171 ( .B1(n14821), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n11865), 
        .ZN(n11866) );
  OAI21_X1 U14172 ( .B1(n13375), .B2(n14839), .A(n11866), .ZN(n11867) );
  NOR2_X1 U14173 ( .A1(n11868), .A2(n11867), .ZN(n11869) );
  NAND2_X1 U14174 ( .A1(n11870), .A2(n11869), .ZN(P2_U3229) );
  NAND2_X1 U14175 ( .A1(n11872), .A2(n12712), .ZN(n11873) );
  XNOR2_X1 U14176 ( .A(n11874), .B(n12567), .ZN(n12525) );
  XNOR2_X1 U14177 ( .A(n12525), .B(n12526), .ZN(n12523) );
  XNOR2_X1 U14178 ( .A(n12524), .B(n12523), .ZN(n11881) );
  NAND2_X1 U14179 ( .A1(n12700), .A2(n11875), .ZN(n11877) );
  AND2_X1 U14180 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n11933) );
  AOI21_X1 U14181 ( .B1(n12695), .B2(n12712), .A(n11933), .ZN(n11876) );
  OAI211_X1 U14182 ( .C1(n12625), .C2(n12697), .A(n11877), .B(n11876), .ZN(
        n11878) );
  AOI21_X1 U14183 ( .B1(n11879), .B2(n6477), .A(n11878), .ZN(n11880) );
  OAI21_X1 U14184 ( .B1(n11881), .B2(n12689), .A(n11880), .ZN(P3_U3155) );
  OAI211_X1 U14185 ( .C1(n11882), .C2(n7998), .A(n13019), .B(n13017), .ZN(
        n11884) );
  AOI22_X1 U14186 ( .A1(n13004), .A2(n13022), .B1(n13023), .B2(n12710), .ZN(
        n11883) );
  NAND2_X1 U14187 ( .A1(n11884), .A2(n11883), .ZN(n13083) );
  INV_X1 U14188 ( .A(n13083), .ZN(n11891) );
  OAI21_X1 U14189 ( .B1(n11887), .B2(n11886), .A(n11885), .ZN(n13084) );
  INV_X1 U14190 ( .A(n12627), .ZN(n13130) );
  AOI22_X1 U14191 ( .A1(n15032), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15014), 
        .B2(n12622), .ZN(n11888) );
  OAI21_X1 U14192 ( .B1(n13130), .B2(n13031), .A(n11888), .ZN(n11889) );
  AOI21_X1 U14193 ( .B1(n13084), .B2(n13033), .A(n11889), .ZN(n11890) );
  OAI21_X1 U14194 ( .B1(n11891), .B2(n15032), .A(n11890), .ZN(P3_U3217) );
  INV_X1 U14195 ( .A(n11892), .ZN(n11893) );
  NAND2_X1 U14196 ( .A1(n11894), .A2(n11893), .ZN(n11895) );
  XNOR2_X1 U14197 ( .A(n11976), .B(n13222), .ZN(n13146) );
  AOI22_X1 U14198 ( .A1(n11898), .A2(n13276), .B1(n13306), .B2(n13629), .ZN(
        n11905) );
  AND2_X1 U14199 ( .A1(n13629), .A2(n9793), .ZN(n11897) );
  INV_X1 U14200 ( .A(n13149), .ZN(n11904) );
  AOI22_X1 U14201 ( .A1(n13298), .A2(n11899), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11900) );
  OAI21_X1 U14202 ( .B1(n11901), .B2(n14816), .A(n11900), .ZN(n11902) );
  AOI21_X1 U14203 ( .B1(n11976), .B2(n14812), .A(n11902), .ZN(n11903) );
  OAI21_X1 U14204 ( .B1(n11905), .B2(n11904), .A(n11903), .ZN(P2_U3213) );
  INV_X1 U14205 ( .A(n12183), .ZN(n11907) );
  OAI222_X1 U14206 ( .A1(n11906), .A2(P1_U3086), .B1(n14391), .B2(n11907), 
        .C1(n12184), .C2(n14396), .ZN(P1_U3329) );
  OAI222_X1 U14207 ( .A1(n13819), .A2(n11909), .B1(P2_U3088), .B2(n11908), 
        .C1(n11907), .C2(n13817), .ZN(P2_U3301) );
  INV_X1 U14208 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n11912) );
  AOI21_X1 U14209 ( .B1(n11911), .B2(n14581), .A(n11910), .ZN(n11914) );
  MUX2_X1 U14210 ( .A(n11912), .B(n11914), .S(n15089), .Z(n11913) );
  OAI21_X1 U14211 ( .B1(n12705), .B2(n13129), .A(n11913), .ZN(P3_U3435) );
  INV_X1 U14212 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14552) );
  MUX2_X1 U14213 ( .A(n14552), .B(n11914), .S(n15106), .Z(n11915) );
  OAI21_X1 U14214 ( .B1(n12705), .B2(n13087), .A(n11915), .ZN(P3_U3474) );
  NOR2_X1 U14215 ( .A1(n11922), .A2(n11917), .ZN(n11918) );
  INV_X1 U14216 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n15259) );
  NAND2_X1 U14217 ( .A1(n12752), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12753) );
  OAI21_X1 U14218 ( .B1(P3_REG1_REG_14__SCAN_IN), .B2(n12752), .A(n12753), 
        .ZN(n11929) );
  AOI21_X1 U14219 ( .B1(n11919), .B2(n11929), .A(n12746), .ZN(n11939) );
  NOR2_X1 U14220 ( .A1(n11922), .A2(n11923), .ZN(n11924) );
  INV_X1 U14221 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14990) );
  XNOR2_X1 U14222 ( .A(n12752), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12766) );
  XNOR2_X1 U14223 ( .A(n12767), .B(n12766), .ZN(n11937) );
  OAI21_X1 U14224 ( .B1(n11927), .B2(n11926), .A(n11925), .ZN(n14998) );
  MUX2_X1 U14225 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n13141), .Z(n11928) );
  XNOR2_X1 U14226 ( .A(n11928), .B(n14993), .ZN(n14999) );
  NOR2_X1 U14227 ( .A1(n11928), .A2(n14993), .ZN(n11931) );
  MUX2_X1 U14228 ( .A(n12766), .B(n11929), .S(n13141), .Z(n11930) );
  OAI21_X1 U14229 ( .B1(n14997), .B2(n11931), .A(n11930), .ZN(n11932) );
  NAND3_X1 U14230 ( .A1(n11932), .A2(n12778), .A3(n12755), .ZN(n11935) );
  AOI21_X1 U14231 ( .B1(n14987), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n11933), 
        .ZN(n11934) );
  OAI211_X1 U14232 ( .C1(n14994), .C2(n12752), .A(n11935), .B(n11934), .ZN(
        n11936) );
  AOI21_X1 U14233 ( .B1(n11937), .B2(n12820), .A(n11936), .ZN(n11938) );
  OAI21_X1 U14234 ( .B1(n11939), .B2(n15002), .A(n11938), .ZN(P3_U3196) );
  INV_X1 U14235 ( .A(n11940), .ZN(n11942) );
  INV_X1 U14236 ( .A(SI_30_), .ZN(n11941) );
  OAI222_X1 U14237 ( .A1(P3_U3151), .A2(n11943), .B1(n6484), .B2(n11942), .C1(
        n11941), .C2(n13143), .ZN(P3_U3265) );
  INV_X1 U14238 ( .A(n13811), .ZN(n11944) );
  OR2_X1 U14239 ( .A1(n11976), .A2(n13258), .ZN(n11946) );
  NOR2_X1 U14240 ( .A1(n13744), .A2(n13269), .ZN(n13601) );
  NOR2_X1 U14241 ( .A1(n13600), .A2(n13601), .ZN(n11949) );
  NOR2_X1 U14242 ( .A1(n13590), .A2(n13344), .ZN(n11951) );
  INV_X1 U14243 ( .A(n13343), .ZN(n13576) );
  NAND2_X1 U14244 ( .A1(n13546), .A2(n13549), .ZN(n11955) );
  NAND2_X1 U14245 ( .A1(n13724), .A2(n13300), .ZN(n11954) );
  NAND2_X1 U14246 ( .A1(n11955), .A2(n11954), .ZN(n13536) );
  INV_X1 U14247 ( .A(n13341), .ZN(n13517) );
  AND2_X1 U14248 ( .A1(n13539), .A2(n13517), .ZN(n11957) );
  OR2_X1 U14249 ( .A1(n13539), .A2(n13517), .ZN(n11956) );
  NAND2_X1 U14250 ( .A1(n13515), .A2(n13520), .ZN(n11961) );
  OR2_X1 U14251 ( .A1(n13526), .A2(n11959), .ZN(n11960) );
  NAND2_X1 U14252 ( .A1(n11961), .A2(n11960), .ZN(n13502) );
  NAND2_X1 U14253 ( .A1(n13502), .A2(n13509), .ZN(n11963) );
  INV_X1 U14254 ( .A(n13339), .ZN(n13518) );
  OR2_X1 U14255 ( .A1(n13507), .A2(n13518), .ZN(n11962) );
  NAND2_X1 U14256 ( .A1(n13455), .A2(n11967), .ZN(n13432) );
  INV_X1 U14257 ( .A(n13415), .ZN(n13424) );
  OR2_X1 U14258 ( .A1(n13769), .A2(n13459), .ZN(n13425) );
  NAND3_X1 U14259 ( .A1(n13433), .A2(n13424), .A3(n13425), .ZN(n13423) );
  NAND2_X1 U14260 ( .A1(n13423), .A2(n11968), .ZN(n11970) );
  INV_X1 U14261 ( .A(P2_B_REG_SCAN_IN), .ZN(n11971) );
  NOR2_X1 U14262 ( .A1(n13816), .A2(n11971), .ZN(n11972) );
  NOR2_X1 U14263 ( .A1(n13631), .A2(n11972), .ZN(n13405) );
  INV_X1 U14264 ( .A(n13700), .ZN(n13288) );
  INV_X1 U14265 ( .A(n11976), .ZN(n13795) );
  INV_X1 U14266 ( .A(n13600), .ZN(n11979) );
  INV_X1 U14267 ( .A(n13608), .ZN(n13789) );
  AOI21_X1 U14268 ( .B1(n13263), .B2(n13590), .A(n13577), .ZN(n13561) );
  INV_X1 U14269 ( .A(n11980), .ZN(n11982) );
  NOR2_X1 U14270 ( .A1(n13724), .A2(n13342), .ZN(n11984) );
  INV_X1 U14271 ( .A(n13724), .ZN(n11983) );
  INV_X1 U14272 ( .A(n13509), .ZN(n11986) );
  NOR2_X1 U14273 ( .A1(n13507), .A2(n13339), .ZN(n11985) );
  AOI21_X1 U14274 ( .B1(n13510), .B2(n11986), .A(n11985), .ZN(n13496) );
  NAND2_X1 U14275 ( .A1(n13773), .A2(n13279), .ZN(n11987) );
  NOR2_X1 U14276 ( .A1(n13688), .A2(n13467), .ZN(n11988) );
  INV_X1 U14277 ( .A(n13688), .ZN(n13454) );
  NAND2_X1 U14278 ( .A1(n13416), .A2(n13415), .ZN(n11989) );
  NAND2_X1 U14279 ( .A1(n11989), .A2(n7428), .ZN(n11991) );
  XNOR2_X1 U14280 ( .A(n11991), .B(n11990), .ZN(n13671) );
  NOR2_X1 U14281 ( .A1(n13608), .A2(n13620), .ZN(n13611) );
  NAND2_X1 U14282 ( .A1(n13590), .A2(n13611), .ZN(n13583) );
  NAND2_X1 U14283 ( .A1(n11994), .A2(n13417), .ZN(n13408) );
  OAI211_X1 U14284 ( .C1(n11994), .C2(n13417), .A(n13521), .B(n13408), .ZN(
        n13674) );
  OAI22_X1 U14285 ( .A1(n13642), .A2(n11996), .B1(n11995), .B2(n13639), .ZN(
        n11997) );
  AOI21_X1 U14286 ( .B1(n13672), .B2(n13655), .A(n11997), .ZN(n11998) );
  OAI21_X1 U14287 ( .B1(n13674), .B2(n13659), .A(n11998), .ZN(n11999) );
  AOI21_X1 U14288 ( .B1(n13671), .B2(n13656), .A(n11999), .ZN(n12000) );
  OAI21_X1 U14289 ( .B1(n13676), .B2(n13595), .A(n12000), .ZN(P2_U3236) );
  INV_X1 U14290 ( .A(n12431), .ZN(n13806) );
  OAI222_X1 U14291 ( .A1(n14391), .A2(n13806), .B1(n12001), .B2(P1_U3086), 
        .C1(n12432), .C2(n14396), .ZN(P1_U3325) );
  INV_X1 U14292 ( .A(n12002), .ZN(n12005) );
  INV_X1 U14293 ( .A(n12003), .ZN(n12004) );
  AOI22_X1 U14294 ( .A1(n12008), .A2(n12205), .B1(n12175), .B2(n13963), .ZN(
        n12009) );
  XOR2_X1 U14295 ( .A(n12020), .B(n12009), .Z(n12012) );
  OAI22_X1 U14296 ( .A1(n14636), .A2(n12230), .B1(n12010), .B2(n12228), .ZN(
        n12011) );
  NOR2_X1 U14297 ( .A1(n12012), .A2(n12011), .ZN(n12013) );
  AOI21_X1 U14298 ( .B1(n12012), .B2(n12011), .A(n12013), .ZN(n13830) );
  NAND2_X1 U14299 ( .A1(n13829), .A2(n13830), .ZN(n13828) );
  INV_X1 U14300 ( .A(n12013), .ZN(n12014) );
  AOI22_X1 U14301 ( .A1(n13953), .A2(n12205), .B1(n12175), .B2(n13962), .ZN(
        n12015) );
  XNOR2_X1 U14302 ( .A(n12015), .B(n12020), .ZN(n12017) );
  AOI22_X1 U14303 ( .A1(n13953), .A2(n12175), .B1(n12216), .B2(n13962), .ZN(
        n13945) );
  NAND2_X1 U14304 ( .A1(n14607), .A2(n12205), .ZN(n12019) );
  NAND2_X1 U14305 ( .A1(n13961), .A2(n12175), .ZN(n12018) );
  NAND2_X1 U14306 ( .A1(n12019), .A2(n12018), .ZN(n12021) );
  INV_X1 U14307 ( .A(n12020), .ZN(n12172) );
  XNOR2_X1 U14308 ( .A(n12021), .B(n12172), .ZN(n12024) );
  AND2_X1 U14309 ( .A1(n13961), .A2(n12216), .ZN(n12022) );
  AOI21_X1 U14310 ( .B1(n14607), .B2(n12175), .A(n12022), .ZN(n12023) );
  NAND2_X1 U14311 ( .A1(n12024), .A2(n12023), .ZN(n12025) );
  OAI21_X1 U14312 ( .B1(n12024), .B2(n12023), .A(n12025), .ZN(n13875) );
  INV_X1 U14313 ( .A(n12025), .ZN(n13883) );
  INV_X1 U14314 ( .A(n14047), .ZN(n14067) );
  OAI22_X1 U14315 ( .A1(n14619), .A2(n12231), .B1(n14067), .B2(n12230), .ZN(
        n12026) );
  XNOR2_X1 U14316 ( .A(n12026), .B(n12172), .ZN(n12029) );
  OR2_X1 U14317 ( .A1(n14619), .A2(n12230), .ZN(n12028) );
  NAND2_X1 U14318 ( .A1(n14047), .A2(n12216), .ZN(n12027) );
  AND2_X1 U14319 ( .A1(n12028), .A2(n12027), .ZN(n12030) );
  NAND2_X1 U14320 ( .A1(n12029), .A2(n12030), .ZN(n12034) );
  INV_X1 U14321 ( .A(n12029), .ZN(n12032) );
  INV_X1 U14322 ( .A(n12030), .ZN(n12031) );
  NAND2_X1 U14323 ( .A1(n12032), .A2(n12031), .ZN(n12033) );
  AND2_X1 U14324 ( .A1(n12034), .A2(n12033), .ZN(n13882) );
  NAND2_X1 U14325 ( .A1(n13881), .A2(n12034), .ZN(n13927) );
  AOI22_X1 U14326 ( .A1(n12041), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n12040), 
        .B2(n14019), .ZN(n12036) );
  OAI22_X1 U14327 ( .A1(n14366), .A2(n12230), .B1(n13851), .B2(n12228), .ZN(
        n12058) );
  OAI22_X1 U14328 ( .A1(n14366), .A2(n12231), .B1(n13851), .B2(n12230), .ZN(
        n12038) );
  XNOR2_X1 U14329 ( .A(n12038), .B(n12020), .ZN(n12057) );
  XOR2_X1 U14330 ( .A(n12058), .B(n12057), .Z(n13928) );
  NAND2_X1 U14331 ( .A1(n12039), .A2(n12457), .ZN(n12043) );
  AOI22_X1 U14332 ( .A1(n12041), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14609), 
        .B2(n12040), .ZN(n12042) );
  NAND2_X2 U14333 ( .A1(n12043), .A2(n12042), .ZN(n12379) );
  NAND2_X1 U14334 ( .A1(n12379), .A2(n12205), .ZN(n12054) );
  INV_X1 U14335 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n12044) );
  NAND2_X1 U14336 ( .A1(n12045), .A2(n12044), .ZN(n12046) );
  NAND2_X1 U14337 ( .A1(n12069), .A2(n12046), .ZN(n14253) );
  OR2_X1 U14338 ( .A1(n14253), .A2(n12092), .ZN(n12052) );
  INV_X1 U14339 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14016) );
  NAND2_X1 U14340 ( .A1(n12440), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n12048) );
  NAND2_X1 U14341 ( .A1(n12441), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n12047) );
  OAI211_X1 U14342 ( .C1(n12049), .C2(n14016), .A(n12048), .B(n12047), .ZN(
        n12050) );
  INV_X1 U14343 ( .A(n12050), .ZN(n12051) );
  AND2_X1 U14344 ( .A1(n12052), .A2(n12051), .ZN(n12378) );
  INV_X1 U14345 ( .A(n12378), .ZN(n14074) );
  NAND2_X1 U14346 ( .A1(n14074), .A2(n12175), .ZN(n12053) );
  NAND2_X1 U14347 ( .A1(n12054), .A2(n12053), .ZN(n12055) );
  XNOR2_X1 U14348 ( .A(n12055), .B(n12020), .ZN(n12062) );
  NOR2_X1 U14349 ( .A1(n12378), .A2(n12228), .ZN(n12056) );
  AOI21_X1 U14350 ( .B1(n12379), .B2(n12175), .A(n12056), .ZN(n12063) );
  XNOR2_X1 U14351 ( .A(n12062), .B(n12063), .ZN(n13849) );
  INV_X1 U14352 ( .A(n12057), .ZN(n12060) );
  INV_X1 U14353 ( .A(n12058), .ZN(n12059) );
  NAND2_X1 U14354 ( .A1(n12060), .A2(n12059), .ZN(n13847) );
  NAND2_X1 U14355 ( .A1(n13926), .A2(n12061), .ZN(n13848) );
  INV_X1 U14356 ( .A(n12062), .ZN(n12064) );
  NAND2_X1 U14357 ( .A1(n12065), .A2(n12457), .ZN(n12068) );
  OR2_X1 U14358 ( .A1(n12458), .A2(n12066), .ZN(n12067) );
  INV_X1 U14359 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13907) );
  NAND2_X1 U14360 ( .A1(n12069), .A2(n13907), .ZN(n12070) );
  NAND2_X1 U14361 ( .A1(n12085), .A2(n12070), .ZN(n14238) );
  INV_X1 U14362 ( .A(n14238), .ZN(n12071) );
  NAND2_X1 U14363 ( .A1(n12071), .A2(n9937), .ZN(n12077) );
  INV_X1 U14364 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n12074) );
  INV_X1 U14365 ( .A(n12441), .ZN(n12438) );
  NAND2_X1 U14366 ( .A1(n12439), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n12073) );
  NAND2_X1 U14367 ( .A1(n12440), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n12072) );
  OAI211_X1 U14368 ( .C1(n12074), .C2(n12438), .A(n12073), .B(n12072), .ZN(
        n12075) );
  INV_X1 U14369 ( .A(n12075), .ZN(n12076) );
  OAI22_X1 U14370 ( .A1(n14241), .A2(n12230), .B1(n14077), .B2(n12228), .ZN(
        n12080) );
  OAI22_X1 U14371 ( .A1(n14241), .A2(n12231), .B1(n14077), .B2(n12230), .ZN(
        n12078) );
  XNOR2_X1 U14372 ( .A(n12078), .B(n12020), .ZN(n12079) );
  XOR2_X1 U14373 ( .A(n12080), .B(n12079), .Z(n13902) );
  OR2_X1 U14374 ( .A1(n12081), .A2(n12141), .ZN(n12084) );
  OR2_X1 U14375 ( .A1(n12458), .A2(n12082), .ZN(n12083) );
  NAND2_X1 U14376 ( .A1(n14346), .A2(n12205), .ZN(n12094) );
  INV_X1 U14377 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13859) );
  AND2_X1 U14378 ( .A1(n12085), .A2(n13859), .ZN(n12086) );
  OR2_X1 U14379 ( .A1(n12086), .A2(n12104), .ZN(n14224) );
  INV_X1 U14380 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n12089) );
  NAND2_X1 U14381 ( .A1(n12440), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n12088) );
  NAND2_X1 U14382 ( .A1(n12439), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n12087) );
  OAI211_X1 U14383 ( .C1(n12438), .C2(n12089), .A(n12088), .B(n12087), .ZN(
        n12090) );
  INV_X1 U14384 ( .A(n12090), .ZN(n12091) );
  NAND2_X1 U14385 ( .A1(n14079), .A2(n12175), .ZN(n12093) );
  NAND2_X1 U14386 ( .A1(n12094), .A2(n12093), .ZN(n12095) );
  XNOR2_X1 U14387 ( .A(n12095), .B(n12020), .ZN(n12099) );
  NAND2_X1 U14388 ( .A1(n14346), .A2(n12175), .ZN(n12097) );
  NAND2_X1 U14389 ( .A1(n14079), .A2(n12216), .ZN(n12096) );
  NAND2_X1 U14390 ( .A1(n12097), .A2(n12096), .ZN(n12098) );
  NOR2_X1 U14391 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  AOI21_X1 U14392 ( .B1(n12099), .B2(n12098), .A(n12100), .ZN(n13855) );
  INV_X1 U14393 ( .A(n12100), .ZN(n13912) );
  OR2_X1 U14394 ( .A1(n12102), .A2(n12101), .ZN(n12103) );
  XNOR2_X1 U14395 ( .A(n12103), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14399) );
  NAND2_X1 U14396 ( .A1(n14339), .A2(n12205), .ZN(n12113) );
  OR2_X1 U14397 ( .A1(n12104), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n12105) );
  NAND2_X1 U14398 ( .A1(n12104), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n12127) );
  AND2_X1 U14399 ( .A1(n12105), .A2(n12127), .ZN(n14211) );
  NAND2_X1 U14400 ( .A1(n14211), .A2(n9937), .ZN(n12111) );
  INV_X1 U14401 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n12108) );
  NAND2_X1 U14402 ( .A1(n12439), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n12107) );
  NAND2_X1 U14403 ( .A1(n12440), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n12106) );
  OAI211_X1 U14404 ( .C1(n12108), .C2(n12438), .A(n12107), .B(n12106), .ZN(
        n12109) );
  INV_X1 U14405 ( .A(n12109), .ZN(n12110) );
  NAND2_X1 U14406 ( .A1(n12111), .A2(n12110), .ZN(n14082) );
  NAND2_X1 U14407 ( .A1(n14082), .A2(n12175), .ZN(n12112) );
  NAND2_X1 U14408 ( .A1(n12113), .A2(n12112), .ZN(n12114) );
  XNOR2_X1 U14409 ( .A(n12114), .B(n12172), .ZN(n12116) );
  AND2_X1 U14410 ( .A1(n14082), .A2(n12216), .ZN(n12115) );
  AOI21_X1 U14411 ( .B1(n14339), .B2(n12175), .A(n12115), .ZN(n12117) );
  NAND2_X1 U14412 ( .A1(n12116), .A2(n12117), .ZN(n12121) );
  INV_X1 U14413 ( .A(n12116), .ZN(n12119) );
  INV_X1 U14414 ( .A(n12117), .ZN(n12118) );
  NAND2_X1 U14415 ( .A1(n12119), .A2(n12118), .ZN(n12120) );
  NAND2_X1 U14416 ( .A1(n12121), .A2(n12120), .ZN(n13911) );
  INV_X1 U14417 ( .A(n12121), .ZN(n13839) );
  OR2_X1 U14418 ( .A1(n12122), .A2(n12141), .ZN(n12125) );
  INV_X1 U14419 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12123) );
  OR2_X1 U14420 ( .A1(n12458), .A2(n12123), .ZN(n12124) );
  NAND2_X1 U14421 ( .A1(n14332), .A2(n12205), .ZN(n12133) );
  NAND2_X1 U14422 ( .A1(n12439), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n12131) );
  NAND2_X1 U14423 ( .A1(n12223), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n12130) );
  INV_X1 U14424 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13842) );
  INV_X1 U14425 ( .A(n12127), .ZN(n12126) );
  NAND2_X1 U14426 ( .A1(n12126), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n12147) );
  AOI21_X1 U14427 ( .B1(n13842), .B2(n12127), .A(n12146), .ZN(n13841) );
  NAND2_X1 U14428 ( .A1(n9937), .A2(n13841), .ZN(n12129) );
  NAND2_X1 U14429 ( .A1(n12441), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n12128) );
  NAND4_X1 U14430 ( .A1(n12131), .A2(n12130), .A3(n12129), .A4(n12128), .ZN(
        n14084) );
  NAND2_X1 U14431 ( .A1(n14084), .A2(n12175), .ZN(n12132) );
  NAND2_X1 U14432 ( .A1(n12133), .A2(n12132), .ZN(n12134) );
  XNOR2_X1 U14433 ( .A(n12134), .B(n12172), .ZN(n12136) );
  AND2_X1 U14434 ( .A1(n12216), .A2(n14084), .ZN(n12135) );
  AOI21_X1 U14435 ( .B1(n14332), .B2(n12175), .A(n12135), .ZN(n12137) );
  NAND2_X1 U14436 ( .A1(n12136), .A2(n12137), .ZN(n13891) );
  INV_X1 U14437 ( .A(n12136), .ZN(n12139) );
  INV_X1 U14438 ( .A(n12137), .ZN(n12138) );
  NAND2_X1 U14439 ( .A1(n12139), .A2(n12138), .ZN(n12140) );
  AND2_X1 U14440 ( .A1(n13891), .A2(n12140), .ZN(n13838) );
  NAND2_X1 U14441 ( .A1(n13837), .A2(n13891), .ZN(n12161) );
  OR2_X1 U14442 ( .A1(n12142), .A2(n12141), .ZN(n12145) );
  OR2_X1 U14443 ( .A1(n12458), .A2(n12143), .ZN(n12144) );
  NAND2_X2 U14444 ( .A1(n12145), .A2(n12144), .ZN(n14327) );
  NAND2_X1 U14445 ( .A1(n14327), .A2(n12205), .ZN(n12153) );
  NAND2_X1 U14446 ( .A1(n12439), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U14447 ( .A1(n12440), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n12150) );
  INV_X1 U14448 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13897) );
  AOI21_X1 U14449 ( .B1(n13897), .B2(n12147), .A(n12187), .ZN(n14185) );
  NAND2_X1 U14450 ( .A1(n9937), .A2(n14185), .ZN(n12149) );
  NAND2_X1 U14451 ( .A1(n12441), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n12148) );
  NAND4_X1 U14452 ( .A1(n12151), .A2(n12150), .A3(n12149), .A4(n12148), .ZN(
        n14086) );
  NAND2_X1 U14453 ( .A1(n14086), .A2(n12175), .ZN(n12152) );
  NAND2_X1 U14454 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  XNOR2_X1 U14455 ( .A(n12154), .B(n12172), .ZN(n12156) );
  AND2_X1 U14456 ( .A1(n12216), .A2(n14086), .ZN(n12155) );
  AOI21_X1 U14457 ( .B1(n14327), .B2(n12175), .A(n12155), .ZN(n12157) );
  NAND2_X1 U14458 ( .A1(n12156), .A2(n12157), .ZN(n13864) );
  INV_X1 U14459 ( .A(n12156), .ZN(n12159) );
  INV_X1 U14460 ( .A(n12157), .ZN(n12158) );
  NAND2_X1 U14461 ( .A1(n12159), .A2(n12158), .ZN(n12160) );
  NAND2_X1 U14462 ( .A1(n12161), .A2(n13892), .ZN(n13863) );
  NAND2_X1 U14463 ( .A1(n13863), .A2(n13864), .ZN(n12181) );
  NAND2_X1 U14464 ( .A1(n12162), .A2(n12457), .ZN(n12164) );
  OR2_X1 U14465 ( .A1(n12458), .A2(n15118), .ZN(n12163) );
  NAND2_X1 U14466 ( .A1(n14320), .A2(n12205), .ZN(n12171) );
  NAND2_X1 U14467 ( .A1(n12439), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12169) );
  NAND2_X1 U14468 ( .A1(n12223), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n12168) );
  XNOR2_X1 U14469 ( .A(P1_REG3_REG_25__SCAN_IN), .B(n12165), .ZN(n14169) );
  NAND2_X1 U14470 ( .A1(n9937), .A2(n14169), .ZN(n12167) );
  NAND2_X1 U14471 ( .A1(n12441), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n12166) );
  NAND4_X1 U14472 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n13960) );
  NAND2_X1 U14473 ( .A1(n13960), .A2(n12175), .ZN(n12170) );
  NAND2_X1 U14474 ( .A1(n12171), .A2(n12170), .ZN(n12173) );
  XNOR2_X1 U14475 ( .A(n12173), .B(n12172), .ZN(n12176) );
  AND2_X1 U14476 ( .A1(n12216), .A2(n13960), .ZN(n12174) );
  AOI21_X1 U14477 ( .B1(n14320), .B2(n12175), .A(n12174), .ZN(n12177) );
  NAND2_X1 U14478 ( .A1(n12176), .A2(n12177), .ZN(n12182) );
  INV_X1 U14479 ( .A(n12176), .ZN(n12179) );
  INV_X1 U14480 ( .A(n12177), .ZN(n12178) );
  NAND2_X1 U14481 ( .A1(n12179), .A2(n12178), .ZN(n12180) );
  NAND2_X1 U14482 ( .A1(n12181), .A2(n13865), .ZN(n13867) );
  NAND2_X1 U14483 ( .A1(n12183), .A2(n12457), .ZN(n12186) );
  OR2_X1 U14484 ( .A1(n12458), .A2(n12184), .ZN(n12185) );
  NAND2_X1 U14485 ( .A1(n14315), .A2(n12205), .ZN(n12195) );
  NAND2_X1 U14486 ( .A1(n12439), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12193) );
  NAND2_X1 U14487 ( .A1(n12440), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n12192) );
  NAND3_X1 U14488 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(P1_REG3_REG_26__SCAN_IN), 
        .A3(n12187), .ZN(n12207) );
  INV_X1 U14489 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13939) );
  NAND2_X1 U14490 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n12187), .ZN(n12188) );
  NAND2_X1 U14491 ( .A1(n13939), .A2(n12188), .ZN(n12189) );
  AND2_X1 U14492 ( .A1(n12207), .A2(n12189), .ZN(n14154) );
  NAND2_X1 U14493 ( .A1(n9937), .A2(n14154), .ZN(n12191) );
  NAND2_X1 U14494 ( .A1(n12441), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n12190) );
  NAND4_X1 U14495 ( .A1(n12193), .A2(n12192), .A3(n12191), .A4(n12190), .ZN(
        n14060) );
  NAND2_X1 U14496 ( .A1(n14060), .A2(n12175), .ZN(n12194) );
  NAND2_X1 U14497 ( .A1(n12195), .A2(n12194), .ZN(n12196) );
  XNOR2_X1 U14498 ( .A(n12196), .B(n12020), .ZN(n12200) );
  NAND2_X1 U14499 ( .A1(n14315), .A2(n12175), .ZN(n12198) );
  NAND2_X1 U14500 ( .A1(n14060), .A2(n12216), .ZN(n12197) );
  NAND2_X1 U14501 ( .A1(n12198), .A2(n12197), .ZN(n12199) );
  NOR2_X1 U14502 ( .A1(n12200), .A2(n12199), .ZN(n12201) );
  AOI21_X1 U14503 ( .B1(n12200), .B2(n12199), .A(n12201), .ZN(n13936) );
  INV_X1 U14504 ( .A(n12201), .ZN(n12202) );
  NAND2_X1 U14505 ( .A1(n13815), .A2(n12457), .ZN(n12204) );
  OR2_X1 U14506 ( .A1(n12458), .A2(n15230), .ZN(n12203) );
  NAND2_X1 U14507 ( .A1(n14310), .A2(n12205), .ZN(n12214) );
  NAND2_X1 U14508 ( .A1(n12439), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U14509 ( .A1(n12223), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n12211) );
  INV_X1 U14510 ( .A(n12207), .ZN(n12206) );
  NAND2_X1 U14511 ( .A1(n12206), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n12236) );
  INV_X1 U14512 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n15112) );
  NAND2_X1 U14513 ( .A1(n12207), .A2(n15112), .ZN(n12208) );
  NAND2_X1 U14514 ( .A1(n9937), .A2(n14136), .ZN(n12210) );
  NAND2_X1 U14515 ( .A1(n12441), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n12209) );
  NAND4_X1 U14516 ( .A1(n12212), .A2(n12211), .A3(n12210), .A4(n12209), .ZN(
        n13959) );
  NAND2_X1 U14517 ( .A1(n13959), .A2(n12175), .ZN(n12213) );
  NAND2_X1 U14518 ( .A1(n12214), .A2(n12213), .ZN(n12215) );
  XNOR2_X1 U14519 ( .A(n12215), .B(n12020), .ZN(n12220) );
  NAND2_X1 U14520 ( .A1(n14310), .A2(n12175), .ZN(n12218) );
  NAND2_X1 U14521 ( .A1(n13959), .A2(n12216), .ZN(n12217) );
  NAND2_X1 U14522 ( .A1(n12218), .A2(n12217), .ZN(n12219) );
  NOR2_X1 U14523 ( .A1(n12220), .A2(n12219), .ZN(n12221) );
  AOI21_X1 U14524 ( .B1(n12220), .B2(n12219), .A(n12221), .ZN(n13824) );
  OR2_X1 U14525 ( .A1(n12458), .A2(n15143), .ZN(n12222) );
  NAND2_X1 U14526 ( .A1(n12439), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n12227) );
  NAND2_X1 U14527 ( .A1(n12223), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n12226) );
  XNOR2_X1 U14528 ( .A(n12236), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n12235) );
  NAND2_X1 U14529 ( .A1(n9937), .A2(n12235), .ZN(n12225) );
  NAND2_X1 U14530 ( .A1(n12441), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n12224) );
  OAI22_X1 U14531 ( .A1(n14303), .A2(n12230), .B1(n14061), .B2(n12228), .ZN(
        n12229) );
  XNOR2_X1 U14532 ( .A(n12229), .B(n12020), .ZN(n12233) );
  OAI22_X1 U14533 ( .A1(n14303), .A2(n12231), .B1(n14061), .B2(n12230), .ZN(
        n12232) );
  XNOR2_X1 U14534 ( .A(n12233), .B(n12232), .ZN(n12234) );
  INV_X1 U14535 ( .A(n12235), .ZN(n14120) );
  INV_X1 U14536 ( .A(n13959), .ZN(n14090) );
  NAND2_X1 U14537 ( .A1(n12439), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12241) );
  NAND2_X1 U14538 ( .A1(n12440), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12240) );
  INV_X1 U14539 ( .A(n12236), .ZN(n12237) );
  AND2_X1 U14540 ( .A1(n12237), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14103) );
  NAND2_X1 U14541 ( .A1(n9937), .A2(n14103), .ZN(n12239) );
  NAND2_X1 U14542 ( .A1(n12441), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n12238) );
  NAND4_X1 U14543 ( .A1(n12241), .A2(n12240), .A3(n12239), .A4(n12238), .ZN(
        n13958) );
  INV_X1 U14544 ( .A(n13958), .ZN(n12242) );
  OAI22_X1 U14545 ( .A1(n14090), .A2(n13917), .B1(n12242), .B2(n13916), .ZN(
        n14119) );
  AOI22_X1 U14546 ( .A1(n14119), .A2(n13923), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n12243) );
  OAI21_X1 U14547 ( .B1(n13920), .B2(n14120), .A(n12243), .ZN(n12244) );
  AOI21_X1 U14548 ( .B1(n14062), .B2(n13952), .A(n12244), .ZN(n12245) );
  OAI21_X1 U14549 ( .B1(n12246), .B2(n13955), .A(n12245), .ZN(P1_U3220) );
  INV_X1 U14550 ( .A(n12247), .ZN(n12249) );
  INV_X1 U14551 ( .A(SI_24_), .ZN(n12248) );
  OAI222_X1 U14552 ( .A1(n6484), .A2(n12249), .B1(n13143), .B2(n12248), .C1(
        P3_U3151), .C2(n8032), .ZN(P3_U3271) );
  INV_X1 U14553 ( .A(n12250), .ZN(n12253) );
  OAI222_X1 U14554 ( .A1(n6484), .A2(n12253), .B1(n13143), .B2(n12252), .C1(
        P3_U3151), .C2(n12251), .ZN(P3_U3269) );
  NAND2_X1 U14555 ( .A1(n12445), .A2(n12447), .ZN(n12258) );
  AOI21_X1 U14556 ( .B1(n12263), .B2(n12262), .A(n12261), .ZN(n12264) );
  MUX2_X1 U14557 ( .A(n12265), .B(n12264), .S(n12449), .Z(n12266) );
  OAI21_X1 U14558 ( .B1(n7454), .B2(n7453), .A(n12266), .ZN(n12284) );
  INV_X1 U14559 ( .A(n12277), .ZN(n12267) );
  NAND3_X1 U14560 ( .A1(n12279), .A2(n12451), .A3(n12267), .ZN(n12274) );
  NAND3_X1 U14561 ( .A1(n6483), .A2(n12269), .A3(n12268), .ZN(n12273) );
  INV_X1 U14562 ( .A(n12270), .ZN(n12271) );
  NAND3_X1 U14563 ( .A1(n12279), .A2(n12271), .A3(n6483), .ZN(n12272) );
  NAND3_X1 U14564 ( .A1(n12274), .A2(n12273), .A3(n12272), .ZN(n12276) );
  INV_X1 U14565 ( .A(n12472), .ZN(n12275) );
  INV_X1 U14566 ( .A(n12259), .ZN(n12278) );
  NAND4_X1 U14567 ( .A1(n12279), .A2(n12278), .A3(n6483), .A4(n12277), .ZN(
        n12282) );
  NAND3_X1 U14568 ( .A1(n12451), .A2(n12280), .A3(n13974), .ZN(n12281) );
  NAND3_X1 U14569 ( .A1(n12284), .A2(n12283), .A3(n7452), .ZN(n12291) );
  OAI21_X1 U14570 ( .B1(n12467), .B2(n12286), .A(n12285), .ZN(n12289) );
  OAI21_X1 U14571 ( .B1(n6483), .B2(n13973), .A(n12287), .ZN(n12288) );
  NAND2_X1 U14572 ( .A1(n12289), .A2(n12288), .ZN(n12290) );
  NAND2_X1 U14573 ( .A1(n12291), .A2(n12290), .ZN(n12296) );
  MUX2_X1 U14574 ( .A(n12293), .B(n12292), .S(n6483), .Z(n12295) );
  MUX2_X1 U14575 ( .A(n13972), .B(n14736), .S(n12451), .Z(n12294) );
  OAI21_X1 U14576 ( .B1(n12296), .B2(n12295), .A(n12294), .ZN(n12298) );
  NAND2_X1 U14577 ( .A1(n12296), .A2(n12295), .ZN(n12297) );
  MUX2_X1 U14578 ( .A(n13971), .B(n14716), .S(n12451), .Z(n12300) );
  MUX2_X1 U14579 ( .A(n13971), .B(n14716), .S(n6483), .Z(n12299) );
  INV_X1 U14580 ( .A(n12300), .ZN(n12301) );
  MUX2_X1 U14581 ( .A(n13970), .B(n12302), .S(n6483), .Z(n12306) );
  NAND2_X1 U14582 ( .A1(n12305), .A2(n12306), .ZN(n12304) );
  MUX2_X1 U14583 ( .A(n13970), .B(n12302), .S(n12451), .Z(n12303) );
  NAND2_X1 U14584 ( .A1(n12304), .A2(n12303), .ZN(n12310) );
  INV_X1 U14585 ( .A(n12305), .ZN(n12308) );
  INV_X1 U14586 ( .A(n12306), .ZN(n12307) );
  NAND2_X1 U14587 ( .A1(n12308), .A2(n12307), .ZN(n12309) );
  NAND2_X1 U14588 ( .A1(n12310), .A2(n12309), .ZN(n12312) );
  MUX2_X1 U14589 ( .A(n13969), .B(n14697), .S(n12451), .Z(n12313) );
  MUX2_X1 U14590 ( .A(n13969), .B(n14697), .S(n6483), .Z(n12311) );
  MUX2_X1 U14591 ( .A(n13968), .B(n12314), .S(n6483), .Z(n12316) );
  MUX2_X1 U14592 ( .A(n13968), .B(n12314), .S(n12451), .Z(n12315) );
  MUX2_X1 U14593 ( .A(n13967), .B(n14778), .S(n12451), .Z(n12319) );
  MUX2_X1 U14594 ( .A(n13967), .B(n14778), .S(n6483), .Z(n12317) );
  MUX2_X1 U14595 ( .A(n13966), .B(n12320), .S(n6483), .Z(n12324) );
  MUX2_X1 U14596 ( .A(n13966), .B(n12320), .S(n12451), .Z(n12321) );
  NAND2_X1 U14597 ( .A1(n12322), .A2(n12321), .ZN(n12328) );
  INV_X1 U14598 ( .A(n12323), .ZN(n12326) );
  INV_X1 U14599 ( .A(n12324), .ZN(n12325) );
  NAND2_X1 U14600 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  MUX2_X1 U14601 ( .A(n13965), .B(n12329), .S(n12451), .Z(n12331) );
  MUX2_X1 U14602 ( .A(n13965), .B(n12329), .S(n6483), .Z(n12330) );
  INV_X1 U14603 ( .A(n12331), .ZN(n12332) );
  MUX2_X1 U14604 ( .A(n13964), .B(n12339), .S(n6483), .Z(n12337) );
  OR2_X1 U14605 ( .A1(n12485), .A2(n12337), .ZN(n12335) );
  AND2_X1 U14606 ( .A1(n12349), .A2(n12333), .ZN(n12334) );
  NAND2_X1 U14607 ( .A1(n12336), .A2(n12344), .ZN(n12348) );
  NAND2_X1 U14608 ( .A1(n12344), .A2(n12339), .ZN(n12340) );
  MUX2_X1 U14609 ( .A(n12341), .B(n12340), .S(n12451), .Z(n12342) );
  NOR2_X1 U14610 ( .A1(n12342), .A2(n12485), .ZN(n12346) );
  AOI21_X1 U14611 ( .B1(n12344), .B2(n12343), .A(n12467), .ZN(n12345) );
  NAND2_X1 U14612 ( .A1(n12348), .A2(n12347), .ZN(n12351) );
  OR2_X1 U14613 ( .A1(n12349), .A2(n12451), .ZN(n12350) );
  NAND2_X1 U14614 ( .A1(n12351), .A2(n12350), .ZN(n12360) );
  MUX2_X1 U14615 ( .A(n13961), .B(n14607), .S(n6483), .Z(n12370) );
  AND2_X1 U14616 ( .A1(n12352), .A2(n6483), .ZN(n12369) );
  AOI21_X1 U14617 ( .B1(n12370), .B2(n14047), .A(n12369), .ZN(n12358) );
  INV_X1 U14618 ( .A(n14607), .ZN(n14625) );
  AND2_X1 U14619 ( .A1(n14047), .A2(n12451), .ZN(n12362) );
  INV_X1 U14620 ( .A(n12369), .ZN(n12353) );
  NOR2_X1 U14621 ( .A1(n14047), .A2(n12353), .ZN(n12354) );
  AOI21_X1 U14622 ( .B1(n14625), .B2(n12362), .A(n12354), .ZN(n12364) );
  NAND2_X1 U14623 ( .A1(n12370), .A2(n14067), .ZN(n12355) );
  OR2_X1 U14624 ( .A1(n14607), .A2(n6483), .ZN(n12361) );
  NAND2_X1 U14625 ( .A1(n12355), .A2(n12361), .ZN(n12356) );
  NAND2_X1 U14626 ( .A1(n12356), .A2(n14619), .ZN(n12357) );
  OAI211_X1 U14627 ( .C1(n12358), .C2(n14619), .A(n12364), .B(n12357), .ZN(
        n12359) );
  NAND2_X1 U14628 ( .A1(n12360), .A2(n12359), .ZN(n12376) );
  INV_X1 U14629 ( .A(n12361), .ZN(n12363) );
  AOI21_X1 U14630 ( .B1(n12370), .B2(n12363), .A(n12362), .ZN(n12367) );
  INV_X1 U14631 ( .A(n12370), .ZN(n12365) );
  OAI22_X1 U14632 ( .A1(n12367), .A2(n12366), .B1(n12365), .B2(n12364), .ZN(
        n12368) );
  INV_X1 U14633 ( .A(n12368), .ZN(n12375) );
  NAND2_X1 U14634 ( .A1(n12370), .A2(n12369), .ZN(n12372) );
  OR2_X1 U14635 ( .A1(n14047), .A2(n12451), .ZN(n12371) );
  AOI21_X1 U14636 ( .B1(n12372), .B2(n12371), .A(n14619), .ZN(n12373) );
  INV_X1 U14637 ( .A(n12373), .ZN(n12374) );
  INV_X1 U14638 ( .A(n13851), .ZN(n14051) );
  OR2_X1 U14639 ( .A1(n14267), .A2(n14051), .ZN(n14071) );
  MUX2_X1 U14640 ( .A(n13851), .B(n14366), .S(n12467), .Z(n12377) );
  AND2_X1 U14641 ( .A1(n14267), .A2(n14051), .ZN(n14070) );
  OR2_X1 U14642 ( .A1(n12379), .A2(n12378), .ZN(n12380) );
  NAND2_X1 U14643 ( .A1(n12379), .A2(n12378), .ZN(n14053) );
  MUX2_X1 U14644 ( .A(n14053), .B(n12380), .S(n6483), .Z(n12381) );
  MUX2_X1 U14645 ( .A(n14077), .B(n14241), .S(n6483), .Z(n12383) );
  MUX2_X1 U14646 ( .A(n14054), .B(n14351), .S(n12467), .Z(n12382) );
  OAI21_X1 U14647 ( .B1(n12384), .B2(n12383), .A(n12382), .ZN(n12386) );
  NAND2_X1 U14648 ( .A1(n12384), .A2(n12383), .ZN(n12385) );
  MUX2_X1 U14649 ( .A(n14079), .B(n14346), .S(n12467), .Z(n12388) );
  MUX2_X1 U14650 ( .A(n14079), .B(n14346), .S(n6483), .Z(n12387) );
  INV_X1 U14651 ( .A(n12388), .ZN(n12389) );
  MUX2_X1 U14652 ( .A(n14082), .B(n14339), .S(n6483), .Z(n12393) );
  NAND2_X1 U14653 ( .A1(n12392), .A2(n12393), .ZN(n12391) );
  MUX2_X1 U14654 ( .A(n14082), .B(n14339), .S(n12467), .Z(n12390) );
  NAND2_X1 U14655 ( .A1(n12391), .A2(n12390), .ZN(n12397) );
  INV_X1 U14656 ( .A(n12392), .ZN(n12395) );
  INV_X1 U14657 ( .A(n12393), .ZN(n12394) );
  NAND2_X1 U14658 ( .A1(n12395), .A2(n12394), .ZN(n12396) );
  MUX2_X1 U14659 ( .A(n14084), .B(n14332), .S(n12467), .Z(n12399) );
  MUX2_X1 U14660 ( .A(n14084), .B(n14332), .S(n6483), .Z(n12398) );
  MUX2_X1 U14661 ( .A(n14086), .B(n14327), .S(n6483), .Z(n12401) );
  MUX2_X1 U14662 ( .A(n14086), .B(n14327), .S(n12467), .Z(n12400) );
  INV_X1 U14663 ( .A(n12401), .ZN(n12402) );
  MUX2_X1 U14664 ( .A(n13960), .B(n14320), .S(n12467), .Z(n12405) );
  MUX2_X1 U14665 ( .A(n13960), .B(n14320), .S(n6483), .Z(n12403) );
  INV_X1 U14666 ( .A(n12405), .ZN(n12406) );
  MUX2_X1 U14667 ( .A(n14315), .B(n14060), .S(n12467), .Z(n12410) );
  MUX2_X1 U14668 ( .A(n14060), .B(n14315), .S(n12467), .Z(n12407) );
  INV_X1 U14669 ( .A(n12409), .ZN(n12412) );
  INV_X1 U14670 ( .A(n12410), .ZN(n12411) );
  MUX2_X1 U14671 ( .A(n13959), .B(n14310), .S(n12467), .Z(n12414) );
  NAND2_X1 U14672 ( .A1(n12413), .A2(n12414), .ZN(n12417) );
  MUX2_X1 U14673 ( .A(n13959), .B(n14310), .S(n6483), .Z(n12416) );
  INV_X1 U14674 ( .A(n12414), .ZN(n12415) );
  MUX2_X1 U14675 ( .A(n14061), .B(n14303), .S(n6483), .Z(n12419) );
  MUX2_X1 U14676 ( .A(n14065), .B(n14062), .S(n12467), .Z(n12418) );
  OAI21_X1 U14677 ( .B1(n12420), .B2(n12419), .A(n12418), .ZN(n12422) );
  NAND2_X1 U14678 ( .A1(n12420), .A2(n12419), .ZN(n12421) );
  NAND2_X1 U14679 ( .A1(n12422), .A2(n12421), .ZN(n12427) );
  NAND2_X1 U14680 ( .A1(n13807), .A2(n12457), .ZN(n12424) );
  OR2_X1 U14681 ( .A1(n12458), .A2(n14393), .ZN(n12423) );
  MUX2_X1 U14682 ( .A(n13958), .B(n14297), .S(n12467), .Z(n12428) );
  NAND2_X1 U14683 ( .A1(n12427), .A2(n12428), .ZN(n12426) );
  MUX2_X1 U14684 ( .A(n14297), .B(n13958), .S(n12467), .Z(n12425) );
  INV_X1 U14685 ( .A(n12427), .ZN(n12430) );
  INV_X1 U14686 ( .A(n12428), .ZN(n12429) );
  NAND2_X1 U14687 ( .A1(n12431), .A2(n12457), .ZN(n12434) );
  OR2_X1 U14688 ( .A1(n12458), .A2(n12432), .ZN(n12433) );
  INV_X1 U14689 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n12437) );
  NAND2_X1 U14690 ( .A1(n12440), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n12436) );
  NAND2_X1 U14691 ( .A1(n12439), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n12435) );
  OAI211_X1 U14692 ( .C1(n12438), .C2(n12437), .A(n12436), .B(n12435), .ZN(
        n14099) );
  NAND2_X1 U14693 ( .A1(n12439), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n12444) );
  NAND2_X1 U14694 ( .A1(n12440), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n12443) );
  NAND2_X1 U14695 ( .A1(n12441), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12442) );
  AND3_X1 U14696 ( .A1(n12444), .A2(n12443), .A3(n12442), .ZN(n14038) );
  INV_X1 U14697 ( .A(n12445), .ZN(n12446) );
  OAI22_X1 U14698 ( .A1(n6483), .A2(n14038), .B1(n12447), .B2(n12446), .ZN(
        n12448) );
  AOI22_X1 U14699 ( .A1(n14034), .A2(n12449), .B1(n14099), .B2(n12448), .ZN(
        n12453) );
  OAI21_X1 U14700 ( .B1(n13957), .B2(n12450), .A(n14099), .ZN(n12452) );
  MUX2_X1 U14701 ( .A(n12452), .B(n14293), .S(n12451), .Z(n12455) );
  INV_X1 U14702 ( .A(n12511), .ZN(n12466) );
  NAND2_X1 U14703 ( .A1(n13796), .A2(n12457), .ZN(n12460) );
  OR2_X1 U14704 ( .A1(n12458), .A2(n9352), .ZN(n12459) );
  XOR2_X1 U14705 ( .A(n13957), .B(n14035), .Z(n12497) );
  NAND2_X1 U14706 ( .A1(n12462), .A2(n12461), .ZN(n12463) );
  NAND2_X1 U14707 ( .A1(n12464), .A2(n12463), .ZN(n12504) );
  NOR2_X1 U14708 ( .A1(n12497), .A2(n12504), .ZN(n12465) );
  NAND2_X1 U14709 ( .A1(n12466), .A2(n12465), .ZN(n12513) );
  NOR2_X1 U14710 ( .A1(n14035), .A2(n12467), .ZN(n12503) );
  NAND2_X1 U14711 ( .A1(n12504), .A2(n12508), .ZN(n12499) );
  NAND2_X1 U14712 ( .A1(n14035), .A2(n12467), .ZN(n12501) );
  NOR2_X1 U14713 ( .A1(n12501), .A2(n13957), .ZN(n12468) );
  AOI211_X1 U14714 ( .C1(n12503), .C2(n13957), .A(n12499), .B(n12468), .ZN(
        n12469) );
  XOR2_X1 U14715 ( .A(n14099), .B(n14034), .Z(n12496) );
  XNOR2_X1 U14716 ( .A(n14297), .B(n13958), .ZN(n14093) );
  INV_X1 U14717 ( .A(n14060), .ZN(n14089) );
  XNOR2_X1 U14718 ( .A(n14315), .B(n14089), .ZN(n14152) );
  INV_X1 U14719 ( .A(n13960), .ZN(n14087) );
  XNOR2_X1 U14720 ( .A(n14320), .B(n14087), .ZN(n14173) );
  INV_X1 U14721 ( .A(n14086), .ZN(n14059) );
  XNOR2_X1 U14722 ( .A(n14327), .B(n14059), .ZN(n14058) );
  XNOR2_X1 U14723 ( .A(n14332), .B(n14084), .ZN(n14199) );
  INV_X1 U14724 ( .A(n14082), .ZN(n13858) );
  XNOR2_X1 U14725 ( .A(n7153), .B(n13858), .ZN(n14206) );
  INV_X1 U14726 ( .A(n14079), .ZN(n13918) );
  XNOR2_X1 U14727 ( .A(n14346), .B(n13918), .ZN(n14220) );
  INV_X1 U14728 ( .A(n14249), .ZN(n14073) );
  NOR4_X1 U14729 ( .A1(n9878), .A2(n12471), .A3(n14283), .A4(n12470), .ZN(
        n12475) );
  NAND4_X1 U14730 ( .A1(n12475), .A2(n12474), .A3(n12473), .A4(n12472), .ZN(
        n12476) );
  NOR4_X1 U14731 ( .A1(n12478), .A2(n12477), .A3(n14699), .A4(n12476), .ZN(
        n12481) );
  NAND4_X1 U14732 ( .A1(n12482), .A2(n12481), .A3(n12480), .A4(n12479), .ZN(
        n12483) );
  NOR4_X1 U14733 ( .A1(n12486), .A2(n12485), .A3(n12484), .A4(n12483), .ZN(
        n12489) );
  NAND4_X1 U14734 ( .A1(n14272), .A2(n12489), .A3(n12488), .A4(n12487), .ZN(
        n12490) );
  NOR3_X1 U14735 ( .A1(n14220), .A2(n14073), .A3(n12490), .ZN(n12491) );
  XNOR2_X1 U14736 ( .A(n14351), .B(n14054), .ZN(n14243) );
  NAND4_X1 U14737 ( .A1(n14199), .A2(n14206), .A3(n12491), .A4(n14243), .ZN(
        n12492) );
  NOR4_X1 U14738 ( .A1(n14152), .A2(n14173), .A3(n14058), .A4(n12492), .ZN(
        n12494) );
  NAND2_X1 U14739 ( .A1(n14062), .A2(n14065), .ZN(n14092) );
  OR2_X1 U14740 ( .A1(n14062), .A2(n14065), .ZN(n12493) );
  NAND2_X1 U14741 ( .A1(n14092), .A2(n12493), .ZN(n14112) );
  NAND4_X1 U14742 ( .A1(n14093), .A2(n12494), .A3(n14112), .A4(n14133), .ZN(
        n12495) );
  NOR3_X1 U14743 ( .A1(n12497), .A2(n12496), .A3(n12495), .ZN(n12498) );
  XNOR2_X1 U14744 ( .A(n12498), .B(n14609), .ZN(n12509) );
  NOR3_X1 U14745 ( .A1(n14290), .A2(n13957), .A3(n12499), .ZN(n12502) );
  NOR3_X1 U14746 ( .A1(n12501), .A2(n13957), .A3(n12504), .ZN(n12500) );
  AOI21_X1 U14747 ( .B1(n12502), .B2(n12501), .A(n12500), .ZN(n12507) );
  XOR2_X1 U14748 ( .A(n12504), .B(n12503), .Z(n12505) );
  NAND4_X1 U14749 ( .A1(n12505), .A2(n14290), .A3(n13957), .A4(n12508), .ZN(
        n12506) );
  OAI211_X1 U14750 ( .C1(n12509), .C2(n12508), .A(n12507), .B(n12506), .ZN(
        n12510) );
  AOI21_X1 U14751 ( .B1(n12511), .B2(n12469), .A(n12510), .ZN(n12512) );
  NOR3_X1 U14752 ( .A1(n12514), .A2(n14398), .A3(n13917), .ZN(n12516) );
  OAI21_X1 U14753 ( .B1(n12517), .B2(n12254), .A(P1_B_REG_SCAN_IN), .ZN(n12515) );
  OAI22_X1 U14754 ( .A1(n12518), .A2(n12517), .B1(n12516), .B2(n12515), .ZN(
        P1_U3242) );
  INV_X1 U14755 ( .A(n12519), .ZN(n12520) );
  OAI222_X1 U14756 ( .A1(n13143), .A2(n12522), .B1(P3_U3151), .B2(n12521), 
        .C1(n6484), .C2(n12520), .ZN(P3_U3267) );
  NAND2_X1 U14757 ( .A1(n12525), .A2(n12711), .ZN(n12527) );
  NAND2_X1 U14758 ( .A1(n12528), .A2(n12527), .ZN(n12686) );
  XNOR2_X1 U14759 ( .A(n12529), .B(n12567), .ZN(n12530) );
  NAND2_X1 U14760 ( .A1(n12530), .A2(n12625), .ZN(n12687) );
  INV_X1 U14761 ( .A(n12530), .ZN(n12531) );
  NAND2_X1 U14762 ( .A1(n12531), .A2(n12710), .ZN(n12688) );
  XOR2_X1 U14763 ( .A(n12567), .B(n12627), .Z(n12619) );
  XNOR2_X1 U14764 ( .A(n13028), .B(n12567), .ZN(n12532) );
  XNOR2_X1 U14765 ( .A(n12532), .B(n13004), .ZN(n12630) );
  NAND2_X1 U14766 ( .A1(n12631), .A2(n12630), .ZN(n12535) );
  INV_X1 U14767 ( .A(n12532), .ZN(n12533) );
  NAND2_X1 U14768 ( .A1(n12533), .A2(n13004), .ZN(n12534) );
  NAND2_X1 U14769 ( .A1(n12535), .A2(n12534), .ZN(n12665) );
  XNOR2_X1 U14770 ( .A(n13074), .B(n12567), .ZN(n12536) );
  XNOR2_X1 U14771 ( .A(n12536), .B(n13021), .ZN(n12667) );
  NOR2_X1 U14772 ( .A1(n12536), .A2(n12593), .ZN(n12537) );
  XNOR2_X1 U14773 ( .A(n13120), .B(n12567), .ZN(n12538) );
  XNOR2_X1 U14774 ( .A(n12538), .B(n13005), .ZN(n12590) );
  XNOR2_X1 U14775 ( .A(n12983), .B(n12567), .ZN(n12539) );
  XNOR2_X1 U14776 ( .A(n12539), .B(n12990), .ZN(n12647) );
  INV_X1 U14777 ( .A(n12539), .ZN(n12540) );
  XNOR2_X1 U14778 ( .A(n12605), .B(n12567), .ZN(n12541) );
  NAND2_X1 U14779 ( .A1(n12541), .A2(n12950), .ZN(n12542) );
  OAI21_X1 U14780 ( .B1(n12541), .B2(n12950), .A(n12542), .ZN(n12601) );
  XNOR2_X1 U14781 ( .A(n12662), .B(n12567), .ZN(n12544) );
  INV_X1 U14782 ( .A(n12544), .ZN(n12543) );
  INV_X1 U14783 ( .A(n12551), .ZN(n12549) );
  XNOR2_X1 U14784 ( .A(n12940), .B(n12567), .ZN(n12550) );
  INV_X1 U14785 ( .A(n12550), .ZN(n12548) );
  NAND2_X1 U14786 ( .A1(n12549), .A2(n12548), .ZN(n12552) );
  NAND2_X1 U14787 ( .A1(n12551), .A2(n12550), .ZN(n12638) );
  XNOR2_X1 U14788 ( .A(n13100), .B(n10532), .ZN(n12553) );
  NAND2_X1 U14789 ( .A1(n12553), .A2(n12586), .ZN(n12609) );
  INV_X1 U14790 ( .A(n12553), .ZN(n12554) );
  NAND2_X1 U14791 ( .A1(n12554), .A2(n12935), .ZN(n12555) );
  NAND2_X1 U14792 ( .A1(n12556), .A2(n12639), .ZN(n12608) );
  NAND2_X1 U14793 ( .A1(n12608), .A2(n12609), .ZN(n12560) );
  XNOR2_X1 U14794 ( .A(n13096), .B(n10532), .ZN(n12557) );
  NAND2_X1 U14795 ( .A1(n12557), .A2(n12890), .ZN(n12561) );
  INV_X1 U14796 ( .A(n12557), .ZN(n12558) );
  NAND2_X1 U14797 ( .A1(n12558), .A2(n12920), .ZN(n12559) );
  NAND2_X1 U14798 ( .A1(n12560), .A2(n12610), .ZN(n12612) );
  XNOR2_X1 U14799 ( .A(n12896), .B(n10532), .ZN(n12562) );
  NOR2_X1 U14800 ( .A1(n12562), .A2(n12906), .ZN(n12563) );
  AOI21_X1 U14801 ( .B1(n12562), .B2(n12906), .A(n12563), .ZN(n12679) );
  INV_X1 U14802 ( .A(n12563), .ZN(n12564) );
  XNOR2_X1 U14803 ( .A(n13036), .B(n10532), .ZN(n12565) );
  NOR2_X1 U14804 ( .A1(n12565), .A2(n12708), .ZN(n12566) );
  AOI21_X1 U14805 ( .B1(n12565), .B2(n12708), .A(n12566), .ZN(n12578) );
  XNOR2_X1 U14806 ( .A(n12568), .B(n12567), .ZN(n12569) );
  INV_X1 U14807 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n12570) );
  OAI22_X1 U14808 ( .A1(n12891), .A2(n12652), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12570), .ZN(n12574) );
  INV_X1 U14809 ( .A(n12868), .ZN(n12571) );
  OAI22_X1 U14810 ( .A1(n12572), .A2(n12697), .B1(n12571), .B2(n12672), .ZN(
        n12573) );
  AOI211_X1 U14811 ( .C1(n12575), .C2(n12674), .A(n12574), .B(n12573), .ZN(
        n12576) );
  OAI21_X1 U14812 ( .B1(n12577), .B2(n12689), .A(n12576), .ZN(P3_U3160) );
  INV_X1 U14813 ( .A(n12674), .ZN(n12704) );
  OAI22_X1 U14814 ( .A1(n12878), .A2(n12652), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12579), .ZN(n12581) );
  NOR2_X1 U14815 ( .A1(n12877), .A2(n12697), .ZN(n12580) );
  AOI211_X1 U14816 ( .C1(n12883), .C2(n12700), .A(n12581), .B(n12580), .ZN(
        n12582) );
  AOI21_X1 U14817 ( .B1(n12709), .B2(n12583), .A(n6487), .ZN(n12589) );
  AOI22_X1 U14818 ( .A1(n12695), .A2(n12934), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12585) );
  NAND2_X1 U14819 ( .A1(n12700), .A2(n12941), .ZN(n12584) );
  OAI211_X1 U14820 ( .C1(n12586), .C2(n12697), .A(n12585), .B(n12584), .ZN(
        n12587) );
  AOI21_X1 U14821 ( .B1(n12940), .B2(n6478), .A(n12587), .ZN(n12588) );
  OAI21_X1 U14822 ( .B1(n12589), .B2(n12689), .A(n12588), .ZN(P3_U3156) );
  XNOR2_X1 U14823 ( .A(n12591), .B(n12590), .ZN(n12597) );
  NAND2_X1 U14824 ( .A1(n12649), .A2(n12990), .ZN(n12592) );
  NAND2_X1 U14825 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12835)
         );
  OAI211_X1 U14826 ( .C1(n12593), .C2(n12652), .A(n12592), .B(n12835), .ZN(
        n12595) );
  NOR2_X1 U14827 ( .A1(n13120), .A2(n12704), .ZN(n12594) );
  AOI211_X1 U14828 ( .C1(n12995), .C2(n12700), .A(n12595), .B(n12594), .ZN(
        n12596) );
  OAI21_X1 U14829 ( .B1(n12597), .B2(n12689), .A(n12596), .ZN(P3_U3159) );
  AOI21_X1 U14830 ( .B1(n12601), .B2(n12600), .A(n12599), .ZN(n12607) );
  NAND2_X1 U14831 ( .A1(n12700), .A2(n12967), .ZN(n12603) );
  AOI22_X1 U14832 ( .A1(n12695), .A2(n12990), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12602) );
  OAI211_X1 U14833 ( .C1(n12961), .C2(n12697), .A(n12603), .B(n12602), .ZN(
        n12604) );
  AOI21_X1 U14834 ( .B1(n12605), .B2(n12674), .A(n12604), .ZN(n12606) );
  OAI21_X1 U14835 ( .B1(n12607), .B2(n12689), .A(n12606), .ZN(P3_U3163) );
  INV_X1 U14836 ( .A(n12608), .ZN(n12641) );
  INV_X1 U14837 ( .A(n12609), .ZN(n12611) );
  NOR3_X1 U14838 ( .A1(n12641), .A2(n12611), .A3(n12610), .ZN(n12614) );
  INV_X1 U14839 ( .A(n12612), .ZN(n12613) );
  OAI21_X1 U14840 ( .B1(n12614), .B2(n12613), .A(n12680), .ZN(n12618) );
  AOI22_X1 U14841 ( .A1(n12935), .A2(n12695), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12615) );
  OAI21_X1 U14842 ( .B1(n12878), .B2(n12697), .A(n12615), .ZN(n12616) );
  AOI21_X1 U14843 ( .B1(n12912), .B2(n12700), .A(n12616), .ZN(n12617) );
  OAI211_X1 U14844 ( .C1(n13096), .C2(n12704), .A(n12618), .B(n12617), .ZN(
        P3_U3165) );
  XNOR2_X1 U14845 ( .A(n12619), .B(n12698), .ZN(n12620) );
  XNOR2_X1 U14846 ( .A(n12621), .B(n12620), .ZN(n12629) );
  NAND2_X1 U14847 ( .A1(n12700), .A2(n12622), .ZN(n12624) );
  AND2_X1 U14848 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12763) );
  AOI21_X1 U14849 ( .B1(n12649), .B2(n13004), .A(n12763), .ZN(n12623) );
  OAI211_X1 U14850 ( .C1(n12625), .C2(n12652), .A(n12624), .B(n12623), .ZN(
        n12626) );
  AOI21_X1 U14851 ( .B1(n12627), .B2(n6477), .A(n12626), .ZN(n12628) );
  OAI21_X1 U14852 ( .B1(n12629), .B2(n12689), .A(n12628), .ZN(P3_U3166) );
  XNOR2_X1 U14853 ( .A(n12631), .B(n12630), .ZN(n12637) );
  NAND2_X1 U14854 ( .A1(n12700), .A2(n13029), .ZN(n12634) );
  NOR2_X1 U14855 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12632), .ZN(n12787) );
  AOI21_X1 U14856 ( .B1(n12649), .B2(n13021), .A(n12787), .ZN(n12633) );
  OAI211_X1 U14857 ( .C1(n12698), .C2(n12652), .A(n12634), .B(n12633), .ZN(
        n12635) );
  AOI21_X1 U14858 ( .B1(n13028), .B2(n6478), .A(n12635), .ZN(n12636) );
  OAI21_X1 U14859 ( .B1(n12637), .B2(n12689), .A(n12636), .ZN(P3_U3168) );
  INV_X1 U14860 ( .A(n12638), .ZN(n12640) );
  NOR3_X1 U14861 ( .A1(n6487), .A2(n12640), .A3(n12639), .ZN(n12642) );
  OAI21_X1 U14862 ( .B1(n12642), .B2(n12641), .A(n12680), .ZN(n12646) );
  AOI22_X1 U14863 ( .A1(n12920), .A2(n12649), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12643) );
  OAI21_X1 U14864 ( .B1(n12949), .B2(n12652), .A(n12643), .ZN(n12644) );
  AOI21_X1 U14865 ( .B1(n12927), .B2(n12700), .A(n12644), .ZN(n12645) );
  OAI211_X1 U14866 ( .C1(n13100), .C2(n12704), .A(n12646), .B(n12645), .ZN(
        P3_U3169) );
  XNOR2_X1 U14867 ( .A(n12648), .B(n12647), .ZN(n12655) );
  NAND2_X1 U14868 ( .A1(n12700), .A2(n12984), .ZN(n12651) );
  AOI22_X1 U14869 ( .A1(n12649), .A2(n12976), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12650) );
  OAI211_X1 U14870 ( .C1(n12669), .C2(n12652), .A(n12651), .B(n12650), .ZN(
        n12653) );
  AOI21_X1 U14871 ( .B1(n12983), .B2(n12674), .A(n12653), .ZN(n12654) );
  OAI21_X1 U14872 ( .B1(n12655), .B2(n12689), .A(n12654), .ZN(P3_U3173) );
  INV_X1 U14873 ( .A(n12657), .ZN(n12658) );
  AOI21_X1 U14874 ( .B1(n12934), .B2(n12656), .A(n12658), .ZN(n12664) );
  NAND2_X1 U14875 ( .A1(n12700), .A2(n12953), .ZN(n12660) );
  AOI22_X1 U14876 ( .A1(n12695), .A2(n12976), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12659) );
  OAI211_X1 U14877 ( .C1(n12949), .C2(n12697), .A(n12660), .B(n12659), .ZN(
        n12661) );
  AOI21_X1 U14878 ( .B1(n12662), .B2(n6477), .A(n12661), .ZN(n12663) );
  OAI21_X1 U14879 ( .B1(n12664), .B2(n12689), .A(n12663), .ZN(P3_U3175) );
  XNOR2_X1 U14880 ( .A(n12666), .B(n12667), .ZN(n12676) );
  INV_X1 U14881 ( .A(n12668), .ZN(n13008) );
  NAND2_X1 U14882 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12821)
         );
  OAI21_X1 U14883 ( .B1(n12697), .B2(n12669), .A(n12821), .ZN(n12670) );
  AOI21_X1 U14884 ( .B1(n12695), .B2(n13004), .A(n12670), .ZN(n12671) );
  OAI21_X1 U14885 ( .B1(n13008), .B2(n12672), .A(n12671), .ZN(n12673) );
  AOI21_X1 U14886 ( .B1(n13074), .B2(n6478), .A(n12673), .ZN(n12675) );
  OAI21_X1 U14887 ( .B1(n12676), .B2(n12689), .A(n12675), .ZN(P3_U3178) );
  OAI21_X1 U14888 ( .B1(n12679), .B2(n12678), .A(n12677), .ZN(n12681) );
  NAND2_X1 U14889 ( .A1(n12681), .A2(n12680), .ZN(n12685) );
  AOI22_X1 U14890 ( .A1(n12920), .A2(n12695), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12682) );
  OAI21_X1 U14891 ( .B1(n12891), .B2(n12697), .A(n12682), .ZN(n12683) );
  AOI21_X1 U14892 ( .B1(n12892), .B2(n12700), .A(n12683), .ZN(n12684) );
  OAI211_X1 U14893 ( .C1(n13092), .C2(n12704), .A(n12685), .B(n12684), .ZN(
        P3_U3180) );
  INV_X1 U14894 ( .A(n12688), .ZN(n12693) );
  AOI21_X1 U14895 ( .B1(n12688), .B2(n12687), .A(n12686), .ZN(n12690) );
  NOR2_X1 U14896 ( .A1(n12690), .A2(n12689), .ZN(n12691) );
  OAI21_X1 U14897 ( .B1(n12693), .B2(n12692), .A(n12691), .ZN(n12703) );
  NOR2_X1 U14898 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12694), .ZN(n14560) );
  AOI21_X1 U14899 ( .B1(n12695), .B2(n12711), .A(n14560), .ZN(n12696) );
  OAI21_X1 U14900 ( .B1(n12698), .B2(n12697), .A(n12696), .ZN(n12699) );
  AOI21_X1 U14901 ( .B1(n12701), .B2(n12700), .A(n12699), .ZN(n12702) );
  OAI211_X1 U14902 ( .C1(n12705), .C2(n12704), .A(n12703), .B(n12702), .ZN(
        P3_U3181) );
  MUX2_X1 U14903 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12706), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14904 ( .A(n12707), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12718), .Z(
        P3_U3521) );
  MUX2_X1 U14905 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12708), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14906 ( .A(n12906), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12718), .Z(
        P3_U3517) );
  MUX2_X1 U14907 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12920), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14908 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12935), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14909 ( .A(n12709), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12718), .Z(
        P3_U3514) );
  MUX2_X1 U14910 ( .A(n12934), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12718), .Z(
        P3_U3513) );
  MUX2_X1 U14911 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12990), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14912 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n13005), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14913 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n13021), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14914 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n13004), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14915 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n13024), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14916 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12710), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14917 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12711), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14918 ( .A(n12712), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12718), .Z(
        P3_U3504) );
  MUX2_X1 U14919 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12713), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14920 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12714), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14921 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12715), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14922 ( .A(n12716), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12718), .Z(
        P3_U3499) );
  MUX2_X1 U14923 ( .A(n7984), .B(P3_DATAO_REG_7__SCAN_IN), .S(n12718), .Z(
        P3_U3498) );
  MUX2_X1 U14924 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12717), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14925 ( .A(n12719), .B(P3_DATAO_REG_4__SCAN_IN), .S(n12718), .Z(
        P3_U3495) );
  MUX2_X1 U14926 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12720), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14927 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12721), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14928 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n12722), .S(P3_U3897), .Z(
        P3_U3491) );
  INV_X1 U14929 ( .A(n12723), .ZN(n12727) );
  NAND3_X1 U14930 ( .A1(n12725), .A2(n12724), .A3(n6504), .ZN(n12726) );
  AOI21_X1 U14931 ( .B1(n12727), .B2(n12726), .A(n15008), .ZN(n12728) );
  AOI211_X1 U14932 ( .C1(n14987), .C2(P3_ADDR_REG_6__SCAN_IN), .A(n12729), .B(
        n12728), .ZN(n12745) );
  INV_X1 U14933 ( .A(n12730), .ZN(n12735) );
  NOR3_X1 U14934 ( .A1(n12733), .A2(n12732), .A3(n12731), .ZN(n12734) );
  OAI21_X1 U14935 ( .B1(n12735), .B2(n12734), .A(n12778), .ZN(n12744) );
  NAND2_X1 U14936 ( .A1(n12847), .A2(n12736), .ZN(n12743) );
  INV_X1 U14937 ( .A(n12737), .ZN(n12741) );
  NOR3_X1 U14938 ( .A1(n12739), .A2(n6917), .A3(n12738), .ZN(n12740) );
  OAI21_X1 U14939 ( .B1(n12741), .B2(n12740), .A(n12811), .ZN(n12742) );
  NAND4_X1 U14940 ( .A1(n12745), .A2(n12744), .A3(n12743), .A4(n12742), .ZN(
        P3_U3188) );
  NOR2_X1 U14941 ( .A1(n12769), .A2(n12747), .ZN(n12748) );
  XNOR2_X1 U14942 ( .A(n12747), .B(n12769), .ZN(n14551) );
  NAND2_X1 U14943 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n12783), .ZN(n12749) );
  OAI21_X1 U14944 ( .B1(P3_REG1_REG_16__SCAN_IN), .B2(n12783), .A(n12749), 
        .ZN(n12750) );
  AOI21_X1 U14945 ( .B1(n12751), .B2(n12750), .A(n12781), .ZN(n12780) );
  NAND2_X1 U14946 ( .A1(n12752), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12765) );
  MUX2_X1 U14947 ( .A(n12765), .B(n12753), .S(n13141), .Z(n12754) );
  INV_X1 U14948 ( .A(n12756), .ZN(n12757) );
  MUX2_X1 U14949 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n13141), .Z(n14555) );
  NOR2_X1 U14950 ( .A1(n14554), .A2(n14555), .ZN(n14553) );
  AOI21_X1 U14951 ( .B1(n12757), .B2(n12769), .A(n14553), .ZN(n12792) );
  INV_X1 U14952 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12758) );
  INV_X1 U14953 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13085) );
  MUX2_X1 U14954 ( .A(n12758), .B(n13085), .S(n13141), .Z(n12760) );
  NOR2_X1 U14955 ( .A1(n12760), .A2(n12759), .ZN(n12791) );
  INV_X1 U14956 ( .A(n12791), .ZN(n12761) );
  NAND2_X1 U14957 ( .A1(n12760), .A2(n12759), .ZN(n12790) );
  NAND2_X1 U14958 ( .A1(n12761), .A2(n12790), .ZN(n12762) );
  XNOR2_X1 U14959 ( .A(n12792), .B(n12762), .ZN(n12777) );
  AOI21_X1 U14960 ( .B1(n14987), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n12763), 
        .ZN(n12764) );
  OAI21_X1 U14961 ( .B1(n14994), .B2(n12783), .A(n12764), .ZN(n12776) );
  INV_X1 U14962 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14548) );
  NOR2_X2 U14963 ( .A1(n14547), .A2(n14548), .ZN(n14546) );
  NOR2_X1 U14964 ( .A1(n12769), .A2(n12768), .ZN(n12770) );
  NAND2_X1 U14965 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12783), .ZN(n12771) );
  OAI21_X1 U14966 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12783), .A(n12771), 
        .ZN(n12772) );
  AOI21_X1 U14967 ( .B1(n12773), .B2(n12772), .A(n6537), .ZN(n12774) );
  NOR2_X1 U14968 ( .A1(n12774), .A2(n15008), .ZN(n12775) );
  AOI211_X1 U14969 ( .C1(n12778), .C2(n12777), .A(n12776), .B(n12775), .ZN(
        n12779) );
  OAI21_X1 U14970 ( .B1(n12780), .B2(n15002), .A(n12779), .ZN(P3_U3198) );
  INV_X1 U14971 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13081) );
  AOI21_X1 U14972 ( .B1(n13081), .B2(n12782), .A(n12804), .ZN(n12798) );
  INV_X1 U14973 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12785) );
  AOI21_X1 U14974 ( .B1(n12786), .B2(n12785), .A(n12784), .ZN(n12789) );
  AOI21_X1 U14975 ( .B1(n14987), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12787), 
        .ZN(n12788) );
  OAI21_X1 U14976 ( .B1(n12789), .B2(n15008), .A(n12788), .ZN(n12796) );
  MUX2_X1 U14977 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n13141), .Z(n12801) );
  XOR2_X1 U14978 ( .A(n12813), .B(n12801), .Z(n12794) );
  NOR2_X1 U14979 ( .A1(n12793), .A2(n12794), .ZN(n12799) );
  AOI211_X1 U14980 ( .C1(n12794), .C2(n12793), .A(n15000), .B(n12799), .ZN(
        n12795) );
  AOI211_X1 U14981 ( .C1(n12847), .C2(n12813), .A(n12796), .B(n12795), .ZN(
        n12797) );
  OAI21_X1 U14982 ( .B1(n12798), .B2(n15002), .A(n12797), .ZN(P3_U3199) );
  MUX2_X1 U14983 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n13141), .Z(n12803) );
  AOI21_X1 U14984 ( .B1(n12801), .B2(n12800), .A(n12799), .ZN(n12842) );
  XNOR2_X1 U14985 ( .A(n12842), .B(n12841), .ZN(n12802) );
  NOR2_X1 U14986 ( .A1(n12802), .A2(n12803), .ZN(n12840) );
  AOI21_X1 U14987 ( .B1(n12803), .B2(n12802), .A(n12840), .ZN(n12826) );
  OR2_X1 U14988 ( .A1(n12805), .A2(n12813), .ZN(n12809) );
  INV_X1 U14989 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12806) );
  OR2_X1 U14990 ( .A1(n12841), .A2(n12806), .ZN(n12827) );
  NAND2_X1 U14991 ( .A1(n12841), .A2(n12806), .ZN(n12807) );
  NAND2_X1 U14992 ( .A1(n12827), .A2(n12807), .ZN(n12808) );
  AND3_X1 U14993 ( .A1(n12810), .A2(n12809), .A3(n12808), .ZN(n12812) );
  OAI21_X1 U14994 ( .B1(n12829), .B2(n12812), .A(n12811), .ZN(n12825) );
  INV_X1 U14995 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14540) );
  INV_X1 U14996 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13009) );
  NOR2_X1 U14997 ( .A1(n12841), .A2(n13009), .ZN(n12830) );
  AOI21_X1 U14998 ( .B1(n12841), .B2(n13009), .A(n12830), .ZN(n12818) );
  OAI21_X1 U14999 ( .B1(n12818), .B2(n12817), .A(n12832), .ZN(n12819) );
  NAND2_X1 U15000 ( .A1(n12820), .A2(n12819), .ZN(n12822) );
  OAI211_X1 U15001 ( .C1(n14991), .C2(n14540), .A(n12822), .B(n12821), .ZN(
        n12823) );
  AOI21_X1 U15002 ( .B1(n12841), .B2(n12847), .A(n12823), .ZN(n12824) );
  OAI211_X1 U15003 ( .C1(n12826), .C2(n15000), .A(n12825), .B(n12824), .ZN(
        P3_U3200) );
  XNOR2_X1 U15004 ( .A(n12833), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12839) );
  INV_X1 U15005 ( .A(n12827), .ZN(n12828) );
  INV_X1 U15006 ( .A(n12830), .ZN(n12831) );
  XNOR2_X1 U15007 ( .A(n12833), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12838) );
  NAND2_X1 U15008 ( .A1(n14987), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12834) );
  OAI211_X1 U15009 ( .C1(n15008), .C2(n12836), .A(n12835), .B(n12834), .ZN(
        n12846) );
  MUX2_X1 U15010 ( .A(n12839), .B(n12838), .S(n12837), .Z(n12843) );
  NOR2_X1 U15011 ( .A1(n12844), .A2(n15000), .ZN(n12845) );
  AOI211_X1 U15012 ( .C1(n12848), .C2(n12847), .A(n12846), .B(n12845), .ZN(
        n12849) );
  OAI21_X1 U15013 ( .B1(n12850), .B2(n15002), .A(n12849), .ZN(P3_U3201) );
  INV_X1 U15014 ( .A(n8130), .ZN(n12855) );
  NAND2_X1 U15015 ( .A1(n12853), .A2(n15014), .ZN(n12861) );
  OAI21_X1 U15016 ( .B1(n15032), .B2(n14563), .A(n12861), .ZN(n12856) );
  AOI21_X1 U15017 ( .B1(n15032), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12856), 
        .ZN(n12854) );
  OAI21_X1 U15018 ( .B1(n12855), .B2(n13031), .A(n12854), .ZN(P3_U3202) );
  AOI21_X1 U15019 ( .B1(n15032), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12856), 
        .ZN(n12857) );
  OAI21_X1 U15020 ( .B1(n12858), .B2(n13031), .A(n12857), .ZN(P3_U3203) );
  INV_X1 U15021 ( .A(n12859), .ZN(n12866) );
  NAND2_X1 U15022 ( .A1(n15032), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n12860) );
  OAI211_X1 U15023 ( .C1(n12862), .C2(n13031), .A(n12861), .B(n12860), .ZN(
        n12863) );
  AOI21_X1 U15024 ( .B1(n12864), .B2(n13033), .A(n12863), .ZN(n12865) );
  OAI21_X1 U15025 ( .B1(n12866), .B2(n15032), .A(n12865), .ZN(P3_U3204) );
  INV_X1 U15026 ( .A(n12867), .ZN(n12874) );
  AOI22_X1 U15027 ( .A1(n12868), .A2(n15014), .B1(n15032), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12869) );
  OAI21_X1 U15028 ( .B1(n12870), .B2(n13031), .A(n12869), .ZN(n12871) );
  AOI21_X1 U15029 ( .B1(n12872), .B2(n13033), .A(n12871), .ZN(n12873) );
  OAI21_X1 U15030 ( .B1(n12874), .B2(n15032), .A(n12873), .ZN(P3_U3205) );
  INV_X1 U15031 ( .A(n12879), .ZN(n13039) );
  OAI21_X1 U15032 ( .B1(n12882), .B2(n12881), .A(n12880), .ZN(n13037) );
  AOI22_X1 U15033 ( .A1(n12883), .A2(n15014), .B1(n15032), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12884) );
  OAI21_X1 U15034 ( .B1(n12885), .B2(n13031), .A(n12884), .ZN(n12886) );
  AOI21_X1 U15035 ( .B1(n13037), .B2(n13033), .A(n12886), .ZN(n12887) );
  OAI21_X1 U15036 ( .B1(n13039), .B2(n15032), .A(n12887), .ZN(P3_U3206) );
  XNOR2_X1 U15037 ( .A(n12888), .B(n12897), .ZN(n12889) );
  OAI222_X1 U15038 ( .A1(n12962), .A2(n12891), .B1(n12964), .B2(n12890), .C1(
        n12889), .C2(n12960), .ZN(n13040) );
  INV_X1 U15039 ( .A(n13040), .ZN(n12902) );
  NAND2_X1 U15040 ( .A1(n12892), .A2(n15014), .ZN(n12893) );
  OAI21_X1 U15041 ( .B1(n15030), .B2(n12894), .A(n12893), .ZN(n12895) );
  AOI21_X1 U15042 ( .B1(n12896), .B2(n15016), .A(n12895), .ZN(n12901) );
  NAND2_X1 U15043 ( .A1(n12898), .A2(n12897), .ZN(n12899) );
  NAND2_X1 U15044 ( .A1(n13041), .A2(n13033), .ZN(n12900) );
  OAI211_X1 U15045 ( .C1(n12902), .C2(n15032), .A(n12901), .B(n12900), .ZN(
        P3_U3207) );
  OAI211_X1 U15046 ( .C1(n12905), .C2(n12904), .A(n12903), .B(n13019), .ZN(
        n12908) );
  AOI22_X1 U15047 ( .A1(n12906), .A2(n13022), .B1(n13023), .B2(n12935), .ZN(
        n12907) );
  NAND2_X1 U15048 ( .A1(n12908), .A2(n12907), .ZN(n13044) );
  INV_X1 U15049 ( .A(n13044), .ZN(n12916) );
  OAI21_X1 U15050 ( .B1(n12911), .B2(n12910), .A(n12909), .ZN(n13045) );
  AOI22_X1 U15051 ( .A1(n12912), .A2(n15014), .B1(n15032), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12913) );
  OAI21_X1 U15052 ( .B1(n13096), .B2(n13031), .A(n12913), .ZN(n12914) );
  AOI21_X1 U15053 ( .B1(n13045), .B2(n13033), .A(n12914), .ZN(n12915) );
  OAI21_X1 U15054 ( .B1(n12916), .B2(n15032), .A(n12915), .ZN(P3_U3208) );
  OAI211_X1 U15055 ( .C1(n12918), .C2(n12924), .A(n12917), .B(n13019), .ZN(
        n12922) );
  NOR2_X1 U15056 ( .A1(n12949), .A2(n12964), .ZN(n12919) );
  AOI21_X1 U15057 ( .B1(n12920), .B2(n13022), .A(n12919), .ZN(n12921) );
  NAND2_X1 U15058 ( .A1(n12922), .A2(n12921), .ZN(n13050) );
  INV_X1 U15059 ( .A(n13050), .ZN(n12931) );
  NAND2_X1 U15060 ( .A1(n12923), .A2(n12924), .ZN(n12925) );
  NAND2_X1 U15061 ( .A1(n12926), .A2(n12925), .ZN(n13048) );
  AOI22_X1 U15062 ( .A1(n15032), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n12927), 
        .B2(n15014), .ZN(n12928) );
  OAI21_X1 U15063 ( .B1(n13100), .B2(n13031), .A(n12928), .ZN(n12929) );
  AOI21_X1 U15064 ( .B1(n13048), .B2(n13033), .A(n12929), .ZN(n12930) );
  OAI21_X1 U15065 ( .B1(n12931), .B2(n15032), .A(n12930), .ZN(P3_U3209) );
  OAI211_X1 U15066 ( .C1(n12933), .C2(n12939), .A(n12932), .B(n13019), .ZN(
        n12937) );
  AOI22_X1 U15067 ( .A1(n12935), .A2(n13022), .B1(n13023), .B2(n12934), .ZN(
        n12936) );
  NAND2_X1 U15068 ( .A1(n12937), .A2(n12936), .ZN(n13053) );
  INV_X1 U15069 ( .A(n13053), .ZN(n12945) );
  XNOR2_X1 U15070 ( .A(n12938), .B(n12939), .ZN(n13054) );
  INV_X1 U15071 ( .A(n12940), .ZN(n13104) );
  AOI22_X1 U15072 ( .A1(n15032), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15014), 
        .B2(n12941), .ZN(n12942) );
  OAI21_X1 U15073 ( .B1(n13104), .B2(n13031), .A(n12942), .ZN(n12943) );
  AOI21_X1 U15074 ( .B1(n13054), .B2(n13033), .A(n12943), .ZN(n12944) );
  OAI21_X1 U15075 ( .B1(n12945), .B2(n15032), .A(n12944), .ZN(P3_U3210) );
  XNOR2_X1 U15076 ( .A(n12947), .B(n12946), .ZN(n12948) );
  OAI222_X1 U15077 ( .A1(n12964), .A2(n12950), .B1(n12962), .B2(n12949), .C1(
        n12960), .C2(n12948), .ZN(n13057) );
  INV_X1 U15078 ( .A(n13057), .ZN(n12957) );
  XNOR2_X1 U15079 ( .A(n12951), .B(n12952), .ZN(n13058) );
  AOI22_X1 U15080 ( .A1(n15032), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15014), 
        .B2(n12953), .ZN(n12954) );
  OAI21_X1 U15081 ( .B1(n13108), .B2(n13031), .A(n12954), .ZN(n12955) );
  AOI21_X1 U15082 ( .B1(n13058), .B2(n13033), .A(n12955), .ZN(n12956) );
  OAI21_X1 U15083 ( .B1(n12957), .B2(n15032), .A(n12956), .ZN(P3_U3211) );
  XOR2_X1 U15084 ( .A(n12966), .B(n12958), .Z(n12959) );
  OAI222_X1 U15085 ( .A1(n12964), .A2(n12963), .B1(n12962), .B2(n12961), .C1(
        n12960), .C2(n12959), .ZN(n13061) );
  INV_X1 U15086 ( .A(n13061), .ZN(n12971) );
  XOR2_X1 U15087 ( .A(n12965), .B(n12966), .Z(n13062) );
  AOI22_X1 U15088 ( .A1(n15032), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15014), 
        .B2(n12967), .ZN(n12968) );
  OAI21_X1 U15089 ( .B1(n13112), .B2(n13031), .A(n12968), .ZN(n12969) );
  AOI21_X1 U15090 ( .B1(n13062), .B2(n13033), .A(n12969), .ZN(n12970) );
  OAI21_X1 U15091 ( .B1(n12971), .B2(n15032), .A(n12970), .ZN(P3_U3212) );
  NAND2_X1 U15092 ( .A1(n12972), .A2(n12973), .ZN(n12975) );
  NAND2_X1 U15093 ( .A1(n12975), .A2(n12982), .ZN(n12974) );
  OAI211_X1 U15094 ( .C1(n12975), .C2(n12982), .A(n12974), .B(n13019), .ZN(
        n12978) );
  AOI22_X1 U15095 ( .A1(n12976), .A2(n13022), .B1(n13023), .B2(n13005), .ZN(
        n12977) );
  NAND2_X1 U15096 ( .A1(n12978), .A2(n12977), .ZN(n13065) );
  INV_X1 U15097 ( .A(n13065), .ZN(n12988) );
  INV_X1 U15098 ( .A(n12979), .ZN(n12980) );
  AOI21_X1 U15099 ( .B1(n12982), .B2(n12981), .A(n12980), .ZN(n13066) );
  INV_X1 U15100 ( .A(n12983), .ZN(n13116) );
  AOI22_X1 U15101 ( .A1(n15032), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15014), 
        .B2(n12984), .ZN(n12985) );
  OAI21_X1 U15102 ( .B1(n13116), .B2(n13031), .A(n12985), .ZN(n12986) );
  AOI21_X1 U15103 ( .B1(n13066), .B2(n13033), .A(n12986), .ZN(n12987) );
  OAI21_X1 U15104 ( .B1(n12988), .B2(n15032), .A(n12987), .ZN(P3_U3213) );
  OAI211_X1 U15105 ( .C1(n12989), .C2(n8004), .A(n12972), .B(n13019), .ZN(
        n12992) );
  AOI22_X1 U15106 ( .A1(n12990), .A2(n13022), .B1(n13023), .B2(n13021), .ZN(
        n12991) );
  NAND2_X1 U15107 ( .A1(n12992), .A2(n12991), .ZN(n13069) );
  INV_X1 U15108 ( .A(n13069), .ZN(n12999) );
  XOR2_X1 U15109 ( .A(n12994), .B(n12993), .Z(n13070) );
  AOI22_X1 U15110 ( .A1(n15032), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15014), 
        .B2(n12995), .ZN(n12996) );
  OAI21_X1 U15111 ( .B1(n13120), .B2(n13031), .A(n12996), .ZN(n12997) );
  AOI21_X1 U15112 ( .B1(n13070), .B2(n13033), .A(n12997), .ZN(n12998) );
  OAI21_X1 U15113 ( .B1(n12999), .B2(n15032), .A(n12998), .ZN(P3_U3214) );
  NAND2_X1 U15114 ( .A1(n13001), .A2(n13000), .ZN(n13002) );
  NAND2_X1 U15115 ( .A1(n6598), .A2(n13002), .ZN(n13003) );
  NAND2_X1 U15116 ( .A1(n13003), .A2(n13019), .ZN(n13007) );
  AOI22_X1 U15117 ( .A1(n13022), .A2(n13005), .B1(n13004), .B2(n13023), .ZN(
        n13006) );
  NAND2_X1 U15118 ( .A1(n13007), .A2(n13006), .ZN(n13078) );
  INV_X1 U15119 ( .A(n13078), .ZN(n13015) );
  OAI22_X1 U15120 ( .A1(n15030), .A2(n13009), .B1(n13008), .B2(n15025), .ZN(
        n13010) );
  AOI21_X1 U15121 ( .B1(n13074), .B2(n15016), .A(n13010), .ZN(n13014) );
  NAND2_X1 U15122 ( .A1(n13012), .A2(n13011), .ZN(n13072) );
  NAND3_X1 U15123 ( .A1(n13073), .A2(n13072), .A3(n13033), .ZN(n13013) );
  OAI211_X1 U15124 ( .C1(n13015), .C2(n15032), .A(n13014), .B(n13013), .ZN(
        P3_U3215) );
  NAND3_X1 U15125 ( .A1(n13017), .A2(n6884), .A3(n13016), .ZN(n13018) );
  NAND3_X1 U15126 ( .A1(n13020), .A2(n13019), .A3(n13018), .ZN(n13026) );
  AOI22_X1 U15127 ( .A1(n13024), .A2(n13023), .B1(n13022), .B2(n13021), .ZN(
        n13025) );
  NAND2_X1 U15128 ( .A1(n13026), .A2(n13025), .ZN(n13079) );
  INV_X1 U15129 ( .A(n13079), .ZN(n13035) );
  XNOR2_X1 U15130 ( .A(n13027), .B(n6884), .ZN(n13080) );
  INV_X1 U15131 ( .A(n13028), .ZN(n13125) );
  AOI22_X1 U15132 ( .A1(n15032), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15014), 
        .B2(n13029), .ZN(n13030) );
  OAI21_X1 U15133 ( .B1(n13125), .B2(n13031), .A(n13030), .ZN(n13032) );
  AOI21_X1 U15134 ( .B1(n13080), .B2(n13033), .A(n13032), .ZN(n13034) );
  OAI21_X1 U15135 ( .B1(n13035), .B2(n15032), .A(n13034), .ZN(P3_U3216) );
  AOI22_X1 U15136 ( .A1(n13037), .A2(n14581), .B1(n15065), .B2(n13036), .ZN(
        n13038) );
  NAND2_X1 U15137 ( .A1(n13039), .A2(n13038), .ZN(n13088) );
  MUX2_X1 U15138 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13088), .S(n15106), .Z(
        P3_U3486) );
  INV_X1 U15139 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13042) );
  AOI21_X1 U15140 ( .B1(n13041), .B2(n14581), .A(n13040), .ZN(n13089) );
  MUX2_X1 U15141 ( .A(n13042), .B(n13089), .S(n15106), .Z(n13043) );
  OAI21_X1 U15142 ( .B1(n13092), .B2(n13087), .A(n13043), .ZN(P3_U3485) );
  INV_X1 U15143 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13046) );
  AOI21_X1 U15144 ( .B1(n14581), .B2(n13045), .A(n13044), .ZN(n13093) );
  MUX2_X1 U15145 ( .A(n13046), .B(n13093), .S(n15106), .Z(n13047) );
  OAI21_X1 U15146 ( .B1(n13096), .B2(n13087), .A(n13047), .ZN(P3_U3484) );
  AND2_X1 U15147 ( .A1(n13048), .A2(n14581), .ZN(n13049) );
  MUX2_X1 U15148 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13097), .S(n15106), .Z(
        n13051) );
  INV_X1 U15149 ( .A(n13051), .ZN(n13052) );
  OAI21_X1 U15150 ( .B1(n13100), .B2(n13087), .A(n13052), .ZN(P3_U3483) );
  INV_X1 U15151 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13055) );
  AOI21_X1 U15152 ( .B1(n13054), .B2(n14581), .A(n13053), .ZN(n13101) );
  MUX2_X1 U15153 ( .A(n13055), .B(n13101), .S(n15106), .Z(n13056) );
  OAI21_X1 U15154 ( .B1(n13104), .B2(n13087), .A(n13056), .ZN(P3_U3482) );
  INV_X1 U15155 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13059) );
  AOI21_X1 U15156 ( .B1(n14581), .B2(n13058), .A(n13057), .ZN(n13105) );
  MUX2_X1 U15157 ( .A(n13059), .B(n13105), .S(n15106), .Z(n13060) );
  OAI21_X1 U15158 ( .B1(n13108), .B2(n13087), .A(n13060), .ZN(P3_U3481) );
  INV_X1 U15159 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13063) );
  AOI21_X1 U15160 ( .B1(n13062), .B2(n14581), .A(n13061), .ZN(n13109) );
  MUX2_X1 U15161 ( .A(n13063), .B(n13109), .S(n15106), .Z(n13064) );
  OAI21_X1 U15162 ( .B1(n13112), .B2(n13087), .A(n13064), .ZN(P3_U3480) );
  INV_X1 U15163 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13067) );
  AOI21_X1 U15164 ( .B1(n13066), .B2(n14581), .A(n13065), .ZN(n13113) );
  MUX2_X1 U15165 ( .A(n13067), .B(n13113), .S(n15106), .Z(n13068) );
  OAI21_X1 U15166 ( .B1(n13116), .B2(n13087), .A(n13068), .ZN(P3_U3479) );
  INV_X1 U15167 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n15273) );
  AOI21_X1 U15168 ( .B1(n14581), .B2(n13070), .A(n13069), .ZN(n13117) );
  MUX2_X1 U15169 ( .A(n15273), .B(n13117), .S(n15106), .Z(n13071) );
  OAI21_X1 U15170 ( .B1(n13087), .B2(n13120), .A(n13071), .ZN(P3_U3478) );
  NAND3_X1 U15171 ( .A1(n13073), .A2(n13072), .A3(n14581), .ZN(n13076) );
  NAND2_X1 U15172 ( .A1(n13074), .A2(n15065), .ZN(n13075) );
  NAND2_X1 U15173 ( .A1(n13076), .A2(n13075), .ZN(n13077) );
  MUX2_X1 U15174 ( .A(n13121), .B(P3_REG1_REG_18__SCAN_IN), .S(n15104), .Z(
        P3_U3477) );
  AOI21_X1 U15175 ( .B1(n13080), .B2(n14581), .A(n13079), .ZN(n13122) );
  MUX2_X1 U15176 ( .A(n13081), .B(n13122), .S(n15106), .Z(n13082) );
  OAI21_X1 U15177 ( .B1(n13125), .B2(n13087), .A(n13082), .ZN(P3_U3476) );
  AOI21_X1 U15178 ( .B1(n14581), .B2(n13084), .A(n13083), .ZN(n13126) );
  MUX2_X1 U15179 ( .A(n13085), .B(n13126), .S(n15106), .Z(n13086) );
  OAI21_X1 U15180 ( .B1(n13130), .B2(n13087), .A(n13086), .ZN(P3_U3475) );
  MUX2_X1 U15181 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n13088), .S(n15089), .Z(
        P3_U3454) );
  INV_X1 U15182 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13090) );
  MUX2_X1 U15183 ( .A(n13090), .B(n13089), .S(n15089), .Z(n13091) );
  OAI21_X1 U15184 ( .B1(n13092), .B2(n13129), .A(n13091), .ZN(P3_U3453) );
  INV_X1 U15185 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13094) );
  MUX2_X1 U15186 ( .A(n13094), .B(n13093), .S(n15089), .Z(n13095) );
  OAI21_X1 U15187 ( .B1(n13096), .B2(n13129), .A(n13095), .ZN(P3_U3452) );
  MUX2_X1 U15188 ( .A(n13097), .B(P3_REG0_REG_24__SCAN_IN), .S(n15087), .Z(
        n13098) );
  INV_X1 U15189 ( .A(n13098), .ZN(n13099) );
  OAI21_X1 U15190 ( .B1(n13100), .B2(n13129), .A(n13099), .ZN(P3_U3451) );
  INV_X1 U15191 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13102) );
  MUX2_X1 U15192 ( .A(n13102), .B(n13101), .S(n15089), .Z(n13103) );
  OAI21_X1 U15193 ( .B1(n13104), .B2(n13129), .A(n13103), .ZN(P3_U3450) );
  INV_X1 U15194 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13106) );
  MUX2_X1 U15195 ( .A(n13106), .B(n13105), .S(n15089), .Z(n13107) );
  OAI21_X1 U15196 ( .B1(n13108), .B2(n13129), .A(n13107), .ZN(P3_U3449) );
  INV_X1 U15197 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13110) );
  MUX2_X1 U15198 ( .A(n13110), .B(n13109), .S(n15089), .Z(n13111) );
  OAI21_X1 U15199 ( .B1(n13112), .B2(n13129), .A(n13111), .ZN(P3_U3448) );
  INV_X1 U15200 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13114) );
  MUX2_X1 U15201 ( .A(n13114), .B(n13113), .S(n15089), .Z(n13115) );
  OAI21_X1 U15202 ( .B1(n13116), .B2(n13129), .A(n13115), .ZN(P3_U3447) );
  INV_X1 U15203 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13118) );
  MUX2_X1 U15204 ( .A(n13118), .B(n13117), .S(n15089), .Z(n13119) );
  OAI21_X1 U15205 ( .B1(n13129), .B2(n13120), .A(n13119), .ZN(P3_U3446) );
  MUX2_X1 U15206 ( .A(n13121), .B(P3_REG0_REG_18__SCAN_IN), .S(n15087), .Z(
        P3_U3444) );
  INV_X1 U15207 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13123) );
  MUX2_X1 U15208 ( .A(n13123), .B(n13122), .S(n15089), .Z(n13124) );
  OAI21_X1 U15209 ( .B1(n13125), .B2(n13129), .A(n13124), .ZN(P3_U3441) );
  INV_X1 U15210 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13127) );
  MUX2_X1 U15211 ( .A(n13127), .B(n13126), .S(n15089), .Z(n13128) );
  OAI21_X1 U15212 ( .B1(n13130), .B2(n13129), .A(n13128), .ZN(P3_U3438) );
  MUX2_X1 U15213 ( .A(P3_D_REG_0__SCAN_IN), .B(n13132), .S(n13131), .Z(
        P3_U3376) );
  INV_X1 U15214 ( .A(n13143), .ZN(n13134) );
  NOR4_X1 U15215 ( .A1(n7480), .A2(P3_IR_REG_30__SCAN_IN), .A3(n7083), .A4(
        P3_U3151), .ZN(n13133) );
  AOI21_X1 U15216 ( .B1(n13134), .B2(SI_31_), .A(n13133), .ZN(n13135) );
  OAI21_X1 U15217 ( .B1(n6590), .B2(n6484), .A(n13135), .ZN(P3_U3264) );
  INV_X1 U15218 ( .A(n13136), .ZN(n13138) );
  OAI222_X1 U15219 ( .A1(n13143), .A2(n13139), .B1(n6484), .B2(n13138), .C1(
        n13137), .C2(P3_U3151), .ZN(P3_U3266) );
  INV_X1 U15220 ( .A(n13140), .ZN(n13144) );
  INV_X1 U15221 ( .A(SI_27_), .ZN(n13142) );
  OAI222_X1 U15222 ( .A1(n6484), .A2(n13144), .B1(n13143), .B2(n13142), .C1(
        P3_U3151), .C2(n13141), .ZN(P3_U3268) );
  MUX2_X1 U15223 ( .A(n13145), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  INV_X1 U15224 ( .A(n13146), .ZN(n13147) );
  XNOR2_X1 U15225 ( .A(n13744), .B(n13178), .ZN(n13270) );
  NAND2_X1 U15226 ( .A1(n13345), .A2(n13221), .ZN(n13150) );
  XNOR2_X1 U15227 ( .A(n13270), .B(n13150), .ZN(n13257) );
  NAND2_X1 U15228 ( .A1(n13270), .A2(n13150), .ZN(n13151) );
  NAND2_X1 U15229 ( .A1(n13254), .A2(n13151), .ZN(n13152) );
  XNOR2_X1 U15230 ( .A(n13608), .B(n13178), .ZN(n13155) );
  NOR2_X1 U15231 ( .A1(n13632), .A2(n13521), .ZN(n13153) );
  XNOR2_X1 U15232 ( .A(n13155), .B(n13153), .ZN(n13268) );
  INV_X1 U15233 ( .A(n13153), .ZN(n13154) );
  NAND2_X1 U15234 ( .A1(n13155), .A2(n13154), .ZN(n13156) );
  XNOR2_X1 U15235 ( .A(n13590), .B(n13178), .ZN(n13209) );
  NOR2_X1 U15236 ( .A1(n13263), .A2(n13521), .ZN(n13157) );
  NAND2_X1 U15237 ( .A1(n13209), .A2(n13157), .ZN(n13161) );
  INV_X1 U15238 ( .A(n13209), .ZN(n13159) );
  INV_X1 U15239 ( .A(n13157), .ZN(n13158) );
  NAND2_X1 U15240 ( .A1(n13159), .A2(n13158), .ZN(n13160) );
  NAND2_X1 U15241 ( .A1(n13161), .A2(n13160), .ZN(n13314) );
  NAND2_X1 U15242 ( .A1(n13343), .A2(n13221), .ZN(n13164) );
  XNOR2_X1 U15243 ( .A(n13163), .B(n13164), .ZN(n13211) );
  AND2_X1 U15244 ( .A1(n13211), .A2(n13161), .ZN(n13162) );
  INV_X1 U15245 ( .A(n13163), .ZN(n13165) );
  XNOR2_X1 U15246 ( .A(n13724), .B(n13178), .ZN(n13166) );
  NAND2_X1 U15247 ( .A1(n13342), .A2(n13221), .ZN(n13167) );
  INV_X1 U15248 ( .A(n13166), .ZN(n13294) );
  INV_X1 U15249 ( .A(n13167), .ZN(n13168) );
  NAND2_X1 U15250 ( .A1(n13294), .A2(n13168), .ZN(n13291) );
  XNOR2_X1 U15251 ( .A(n13539), .B(n13222), .ZN(n13171) );
  NAND2_X1 U15252 ( .A1(n13341), .A2(n13221), .ZN(n13169) );
  XNOR2_X1 U15253 ( .A(n13171), .B(n13169), .ZN(n13235) );
  INV_X1 U15254 ( .A(n13169), .ZN(n13170) );
  XNOR2_X1 U15255 ( .A(n13526), .B(n13222), .ZN(n13172) );
  AND2_X1 U15256 ( .A1(n13340), .A2(n9793), .ZN(n13305) );
  XNOR2_X1 U15257 ( .A(n13507), .B(n13222), .ZN(n13173) );
  NAND2_X1 U15258 ( .A1(n13339), .A2(n13221), .ZN(n13198) );
  INV_X1 U15259 ( .A(n13173), .ZN(n13175) );
  AOI22_X1 U15260 ( .A1(n13199), .A2(n13198), .B1(n13175), .B2(n13174), .ZN(
        n13278) );
  XNOR2_X1 U15261 ( .A(n13700), .B(n13178), .ZN(n13244) );
  NAND2_X1 U15262 ( .A1(n13468), .A2(n13221), .ZN(n13176) );
  NOR2_X1 U15263 ( .A1(n13244), .A2(n13176), .ZN(n13177) );
  AOI21_X1 U15264 ( .B1(n13244), .B2(n13176), .A(n13177), .ZN(n13277) );
  NAND2_X1 U15265 ( .A1(n13278), .A2(n13277), .ZN(n13242) );
  INV_X1 U15266 ( .A(n13177), .ZN(n13183) );
  XNOR2_X1 U15267 ( .A(n13773), .B(n13178), .ZN(n13179) );
  NOR2_X1 U15268 ( .A1(n13279), .A2(n13521), .ZN(n13180) );
  NAND2_X1 U15269 ( .A1(n13179), .A2(n13180), .ZN(n13184) );
  INV_X1 U15270 ( .A(n13179), .ZN(n13330) );
  INV_X1 U15271 ( .A(n13180), .ZN(n13181) );
  NAND2_X1 U15272 ( .A1(n13330), .A2(n13181), .ZN(n13182) );
  NAND2_X1 U15273 ( .A1(n13184), .A2(n13182), .ZN(n13243) );
  NAND2_X1 U15274 ( .A1(n13467), .A2(n13221), .ZN(n13187) );
  XNOR2_X1 U15275 ( .A(n13688), .B(n13222), .ZN(n13186) );
  XOR2_X1 U15276 ( .A(n13187), .B(n13186), .Z(n13328) );
  INV_X1 U15277 ( .A(n13184), .ZN(n13185) );
  INV_X1 U15278 ( .A(n13186), .ZN(n13188) );
  NAND2_X1 U15279 ( .A1(n13188), .A2(n13187), .ZN(n13189) );
  XNOR2_X1 U15280 ( .A(n13769), .B(n13222), .ZN(n13191) );
  OR2_X1 U15281 ( .A1(n13325), .A2(n13521), .ZN(n13190) );
  NOR2_X1 U15282 ( .A1(n13191), .A2(n13190), .ZN(n13219) );
  AOI21_X1 U15283 ( .B1(n13191), .B2(n13190), .A(n13219), .ZN(n13192) );
  OAI211_X1 U15284 ( .C1(n13193), .C2(n13192), .A(n13220), .B(n13276), .ZN(
        n13197) );
  NOR2_X1 U15285 ( .A1(n14800), .A2(n13436), .ZN(n13195) );
  OAI22_X1 U15286 ( .A1(n14801), .A2(n13437), .B1(n13442), .B2(n14816), .ZN(
        n13194) );
  AOI211_X1 U15287 ( .C1(P2_REG3_REG_27__SCAN_IN), .C2(P2_U3088), .A(n13195), 
        .B(n13194), .ZN(n13196) );
  OAI211_X1 U15288 ( .C1(n13769), .C2(n13321), .A(n13197), .B(n13196), .ZN(
        P2_U3186) );
  NAND2_X1 U15289 ( .A1(n13306), .A2(n13339), .ZN(n13201) );
  NAND2_X1 U15290 ( .A1(n13276), .A2(n13198), .ZN(n13200) );
  MUX2_X1 U15291 ( .A(n13201), .B(n13200), .S(n13199), .Z(n13207) );
  NAND2_X1 U15292 ( .A1(n13340), .A2(n13628), .ZN(n13203) );
  NAND2_X1 U15293 ( .A1(n13468), .A2(n13466), .ZN(n13202) );
  NAND2_X1 U15294 ( .A1(n13203), .A2(n13202), .ZN(n13706) );
  AOI22_X1 U15295 ( .A1(n13298), .A2(n13706), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13204) );
  OAI21_X1 U15296 ( .B1(n13501), .B2(n14816), .A(n13204), .ZN(n13205) );
  AOI21_X1 U15297 ( .B1(n13507), .B2(n14812), .A(n13205), .ZN(n13206) );
  NAND2_X1 U15298 ( .A1(n13207), .A2(n13206), .ZN(P2_U3188) );
  NAND3_X1 U15299 ( .A1(n13209), .A2(n13306), .A3(n13344), .ZN(n13210) );
  OAI21_X1 U15300 ( .B1(n13208), .B2(n14808), .A(n13210), .ZN(n13213) );
  INV_X1 U15301 ( .A(n13211), .ZN(n13212) );
  NAND2_X1 U15302 ( .A1(n13213), .A2(n13212), .ZN(n13217) );
  NOR2_X1 U15303 ( .A1(n14816), .A2(n13567), .ZN(n13215) );
  AOI22_X1 U15304 ( .A1(n13342), .A2(n13466), .B1(n13628), .B2(n13344), .ZN(
        n13564) );
  NAND2_X1 U15305 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13402)
         );
  OAI21_X1 U15306 ( .B1(n13282), .B2(n13564), .A(n13402), .ZN(n13214) );
  OAI211_X1 U15307 ( .C1(n14808), .C2(n13218), .A(n13217), .B(n13216), .ZN(
        P2_U3191) );
  NAND2_X1 U15308 ( .A1(n13338), .A2(n13221), .ZN(n13223) );
  XOR2_X1 U15309 ( .A(n13223), .B(n13222), .Z(n13224) );
  XNOR2_X1 U15310 ( .A(n13418), .B(n13224), .ZN(n13225) );
  XNOR2_X1 U15311 ( .A(n13226), .B(n13225), .ZN(n13232) );
  OAI22_X1 U15312 ( .A1(n14801), .A2(n13325), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13227), .ZN(n13230) );
  OAI22_X1 U15313 ( .A1(n14800), .A2(n13228), .B1(n13419), .B2(n14816), .ZN(
        n13229) );
  AOI211_X1 U15314 ( .C1(n13680), .C2(n14812), .A(n13230), .B(n13229), .ZN(
        n13231) );
  OAI21_X1 U15315 ( .B1(n13232), .B2(n14808), .A(n13231), .ZN(P2_U3192) );
  INV_X1 U15316 ( .A(n13539), .ZN(n13782) );
  OAI211_X1 U15317 ( .C1(n13233), .C2(n13235), .A(n13234), .B(n13276), .ZN(
        n13241) );
  INV_X1 U15318 ( .A(n13532), .ZN(n13239) );
  AND2_X1 U15319 ( .A1(n13340), .A2(n13466), .ZN(n13236) );
  AOI21_X1 U15320 ( .B1(n13342), .B2(n13628), .A(n13236), .ZN(n13537) );
  OAI22_X1 U15321 ( .A1(n13282), .A2(n13537), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13237), .ZN(n13238) );
  AOI21_X1 U15322 ( .B1(n13239), .B2(n13284), .A(n13238), .ZN(n13240) );
  OAI211_X1 U15323 ( .C1(n13782), .C2(n13321), .A(n13241), .B(n13240), .ZN(
        P2_U3195) );
  AOI21_X1 U15324 ( .B1(n13242), .B2(n13243), .A(n14808), .ZN(n13246) );
  NOR3_X1 U15325 ( .A1(n13244), .A2(n13249), .A3(n13329), .ZN(n13245) );
  NOR2_X1 U15326 ( .A1(n13246), .A2(n13245), .ZN(n13253) );
  OAI22_X1 U15327 ( .A1(n14800), .A2(n13437), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13248), .ZN(n13251) );
  OAI22_X1 U15328 ( .A1(n14801), .A2(n13249), .B1(n14816), .B2(n13476), .ZN(
        n13250) );
  AOI211_X1 U15329 ( .C1(n13475), .C2(n14812), .A(n13251), .B(n13250), .ZN(
        n13252) );
  OAI21_X1 U15330 ( .B1(n13253), .B2(n13247), .A(n13252), .ZN(P2_U3197) );
  INV_X1 U15331 ( .A(n13254), .ZN(n13255) );
  AOI21_X1 U15332 ( .B1(n13257), .B2(n13256), .A(n13255), .ZN(n13262) );
  NAND2_X1 U15333 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14888)
         );
  OAI21_X1 U15334 ( .B1(n14800), .B2(n13632), .A(n14888), .ZN(n13260) );
  OAI22_X1 U15335 ( .A1(n14801), .A2(n13258), .B1(n13616), .B2(n14816), .ZN(
        n13259) );
  AOI211_X1 U15336 ( .C1(n13744), .C2(n14812), .A(n13260), .B(n13259), .ZN(
        n13261) );
  OAI21_X1 U15337 ( .B1(n13262), .B2(n14808), .A(n13261), .ZN(P2_U3198) );
  OR2_X1 U15338 ( .A1(n13263), .A2(n13631), .ZN(n13265) );
  NAND2_X1 U15339 ( .A1(n13345), .A2(n13628), .ZN(n13264) );
  NAND2_X1 U15340 ( .A1(n13265), .A2(n13264), .ZN(n13606) );
  AOI22_X1 U15341 ( .A1(n13298), .A2(n13606), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13266) );
  OAI21_X1 U15342 ( .B1(n13597), .B2(n14816), .A(n13266), .ZN(n13267) );
  AOI21_X1 U15343 ( .B1(n13608), .B2(n14812), .A(n13267), .ZN(n13274) );
  INV_X1 U15344 ( .A(n13268), .ZN(n13272) );
  OAI22_X1 U15345 ( .A1(n13270), .A2(n14808), .B1(n13269), .B2(n13329), .ZN(
        n13271) );
  NAND3_X1 U15346 ( .A1(n13254), .A2(n13272), .A3(n13271), .ZN(n13273) );
  OAI211_X1 U15347 ( .C1(n13275), .C2(n14808), .A(n13274), .B(n13273), .ZN(
        P2_U3200) );
  OAI211_X1 U15348 ( .C1(n13278), .C2(n13277), .A(n13242), .B(n13276), .ZN(
        n13287) );
  INV_X1 U15349 ( .A(n13487), .ZN(n13285) );
  OR2_X1 U15350 ( .A1(n13279), .A2(n13631), .ZN(n13281) );
  NAND2_X1 U15351 ( .A1(n13339), .A2(n13628), .ZN(n13280) );
  NAND2_X1 U15352 ( .A1(n13281), .A2(n13280), .ZN(n13699) );
  INV_X1 U15353 ( .A(n13699), .ZN(n13486) );
  OAI22_X1 U15354 ( .A1(n13282), .A2(n13486), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15141), .ZN(n13283) );
  AOI21_X1 U15355 ( .B1(n13285), .B2(n13284), .A(n13283), .ZN(n13286) );
  OAI211_X1 U15356 ( .C1(n13288), .C2(n13321), .A(n13287), .B(n13286), .ZN(
        P2_U3201) );
  INV_X1 U15357 ( .A(n13233), .ZN(n13295) );
  INV_X1 U15358 ( .A(n13289), .ZN(n13292) );
  AOI21_X1 U15359 ( .B1(n13292), .B2(n13291), .A(n13290), .ZN(n13293) );
  AOI21_X1 U15360 ( .B1(n13295), .B2(n13294), .A(n13293), .ZN(n13304) );
  NAND2_X1 U15361 ( .A1(n13341), .A2(n13466), .ZN(n13297) );
  NAND2_X1 U15362 ( .A1(n13343), .A2(n13628), .ZN(n13296) );
  NAND2_X1 U15363 ( .A1(n13297), .A2(n13296), .ZN(n13547) );
  AOI22_X1 U15364 ( .A1(n13298), .A2(n13547), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13299) );
  OAI21_X1 U15365 ( .B1(n13551), .B2(n14816), .A(n13299), .ZN(n13302) );
  NOR3_X1 U15366 ( .A1(n13233), .A2(n13300), .A3(n13329), .ZN(n13301) );
  AOI211_X1 U15367 ( .C1(n13724), .C2(n14812), .A(n13302), .B(n13301), .ZN(
        n13303) );
  OAI21_X1 U15368 ( .B1(n13304), .B2(n14808), .A(n13303), .ZN(P2_U3205) );
  OR2_X1 U15369 ( .A1(n14808), .A2(n13305), .ZN(n13309) );
  NAND2_X1 U15370 ( .A1(n13306), .A2(n13340), .ZN(n13308) );
  MUX2_X1 U15371 ( .A(n13309), .B(n13308), .S(n13307), .Z(n13313) );
  NOR2_X1 U15372 ( .A1(n14801), .A2(n13517), .ZN(n13311) );
  OAI22_X1 U15373 ( .A1(n14800), .A2(n13518), .B1(n14816), .B2(n13523), .ZN(
        n13310) );
  AOI211_X1 U15374 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3088), .A(n13311), 
        .B(n13310), .ZN(n13312) );
  OAI211_X1 U15375 ( .C1(n13713), .C2(n13321), .A(n13313), .B(n13312), .ZN(
        P2_U3207) );
  AOI21_X1 U15376 ( .B1(n13315), .B2(n13314), .A(n14808), .ZN(n13316) );
  NAND2_X1 U15377 ( .A1(n13316), .A2(n13208), .ZN(n13320) );
  AND2_X1 U15378 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13374) );
  OAI22_X1 U15379 ( .A1(n14801), .A2(n13632), .B1(n14816), .B2(n13586), .ZN(
        n13317) );
  AOI211_X1 U15380 ( .C1(n13318), .C2(n13343), .A(n13374), .B(n13317), .ZN(
        n13319) );
  OAI211_X1 U15381 ( .C1(n13590), .C2(n13321), .A(n13320), .B(n13319), .ZN(
        P2_U3210) );
  AOI21_X1 U15382 ( .B1(n13328), .B2(n13247), .A(n13323), .ZN(n13336) );
  NOR2_X1 U15383 ( .A1(n14816), .A2(n13451), .ZN(n13327) );
  OAI22_X1 U15384 ( .A1(n14800), .A2(n13325), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13324), .ZN(n13326) );
  AOI211_X1 U15385 ( .C1(n13688), .C2(n14812), .A(n13327), .B(n13326), .ZN(
        n13335) );
  INV_X1 U15386 ( .A(n13328), .ZN(n13331) );
  NOR3_X1 U15387 ( .A1(n13331), .A2(n13330), .A3(n13329), .ZN(n13333) );
  INV_X1 U15388 ( .A(n14801), .ZN(n13332) );
  OAI21_X1 U15389 ( .B1(n13333), .B2(n13332), .A(n13458), .ZN(n13334) );
  OAI211_X1 U15390 ( .C1(n13336), .C2(n14808), .A(n13335), .B(n13334), .ZN(
        P2_U3212) );
  MUX2_X1 U15391 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13337), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U15392 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13426), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15393 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13338), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15394 ( .A(n13459), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13360), .Z(
        P2_U3558) );
  MUX2_X1 U15395 ( .A(n13467), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13360), .Z(
        P2_U3557) );
  MUX2_X1 U15396 ( .A(n13458), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13360), .Z(
        P2_U3556) );
  MUX2_X1 U15397 ( .A(n13468), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13360), .Z(
        P2_U3555) );
  MUX2_X1 U15398 ( .A(n13339), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13360), .Z(
        P2_U3554) );
  MUX2_X1 U15399 ( .A(n13340), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13360), .Z(
        P2_U3553) );
  MUX2_X1 U15400 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13341), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U15401 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13342), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15402 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13343), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U15403 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13344), .S(P2_U3947), .Z(
        P2_U3549) );
  MUX2_X1 U15404 ( .A(n13345), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13360), .Z(
        P2_U3547) );
  MUX2_X1 U15405 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13629), .S(P2_U3947), .Z(
        P2_U3546) );
  MUX2_X1 U15406 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13346), .S(P2_U3947), .Z(
        P2_U3545) );
  MUX2_X1 U15407 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13347), .S(P2_U3947), .Z(
        P2_U3544) );
  MUX2_X1 U15408 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13348), .S(P2_U3947), .Z(
        P2_U3543) );
  MUX2_X1 U15409 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13349), .S(P2_U3947), .Z(
        P2_U3542) );
  MUX2_X1 U15410 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13350), .S(P2_U3947), .Z(
        P2_U3541) );
  MUX2_X1 U15411 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13351), .S(P2_U3947), .Z(
        P2_U3540) );
  MUX2_X1 U15412 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13352), .S(P2_U3947), .Z(
        P2_U3539) );
  MUX2_X1 U15413 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13353), .S(P2_U3947), .Z(
        P2_U3538) );
  MUX2_X1 U15414 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13354), .S(P2_U3947), .Z(
        P2_U3537) );
  MUX2_X1 U15415 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13355), .S(P2_U3947), .Z(
        P2_U3536) );
  MUX2_X1 U15416 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13356), .S(P2_U3947), .Z(
        P2_U3535) );
  MUX2_X1 U15417 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13357), .S(P2_U3947), .Z(
        P2_U3534) );
  MUX2_X1 U15418 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13358), .S(P2_U3947), .Z(
        P2_U3533) );
  MUX2_X1 U15419 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13359), .S(P2_U3947), .Z(
        P2_U3532) );
  AOI22_X1 U15420 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n14907), .B1(n13361), 
        .B2(n13598), .ZN(n14912) );
  NAND2_X1 U15421 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n14894), .ZN(n13367) );
  AOI22_X1 U15422 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n14894), .B1(n13362), 
        .B2(n13617), .ZN(n14897) );
  NAND2_X1 U15423 ( .A1(n13364), .A2(n13363), .ZN(n13366) );
  NAND2_X1 U15424 ( .A1(n13366), .A2(n13365), .ZN(n14896) );
  NAND2_X1 U15425 ( .A1(n14897), .A2(n14896), .ZN(n14895) );
  NAND2_X1 U15426 ( .A1(n13367), .A2(n14895), .ZN(n14911) );
  NAND2_X1 U15427 ( .A1(n14912), .A2(n14911), .ZN(n14909) );
  NAND2_X1 U15428 ( .A1(n14907), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13368) );
  INV_X1 U15429 ( .A(n13391), .ZN(n13369) );
  OAI21_X1 U15430 ( .B1(n13371), .B2(n13370), .A(n13369), .ZN(n13372) );
  AOI21_X1 U15431 ( .B1(n13372), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13390), 
        .ZN(n13373) );
  OR2_X1 U15432 ( .A1(n13373), .A2(n14852), .ZN(n13389) );
  AOI21_X1 U15433 ( .B1(n14821), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n13374), 
        .ZN(n13388) );
  NAND2_X1 U15434 ( .A1(n14907), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n13380) );
  NOR2_X1 U15435 ( .A1(n13376), .A2(n13375), .ZN(n13378) );
  NOR2_X1 U15436 ( .A1(n13378), .A2(n13377), .ZN(n14891) );
  XNOR2_X1 U15437 ( .A(n14894), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14890) );
  NOR2_X1 U15438 ( .A1(n14891), .A2(n14890), .ZN(n14889) );
  AOI21_X1 U15439 ( .B1(n14894), .B2(P2_REG1_REG_16__SCAN_IN), .A(n14889), 
        .ZN(n14904) );
  XNOR2_X1 U15440 ( .A(n14907), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14903) );
  NOR2_X1 U15441 ( .A1(n14904), .A2(n14903), .ZN(n14902) );
  INV_X1 U15442 ( .A(n14902), .ZN(n13379) );
  NAND2_X1 U15443 ( .A1(n13380), .A2(n13379), .ZN(n13381) );
  AND2_X1 U15444 ( .A1(n13385), .A2(n13381), .ZN(n13393) );
  NOR2_X1 U15445 ( .A1(n13385), .A2(n13381), .ZN(n13382) );
  NOR2_X1 U15446 ( .A1(n13393), .A2(n13382), .ZN(n13384) );
  INV_X1 U15447 ( .A(n13394), .ZN(n13383) );
  OAI211_X1 U15448 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13384), .A(n14876), 
        .B(n13383), .ZN(n13387) );
  INV_X1 U15449 ( .A(n14839), .ZN(n14908) );
  NAND2_X1 U15450 ( .A1(n14908), .A2(n13385), .ZN(n13386) );
  NAND4_X1 U15451 ( .A1(n13389), .A2(n13388), .A3(n13387), .A4(n13386), .ZN(
        P2_U3232) );
  INV_X1 U15452 ( .A(n14821), .ZN(n14916) );
  XOR2_X1 U15453 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13392), .Z(n13399) );
  INV_X1 U15454 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13395) );
  NAND2_X1 U15455 ( .A1(n13396), .A2(n14876), .ZN(n13397) );
  AOI22_X1 U15456 ( .A1(n13399), .A2(n14910), .B1(n14876), .B2(n13398), .ZN(
        n13401) );
  NAND2_X1 U15457 ( .A1(n13405), .A2(n13404), .ZN(n13667) );
  NOR2_X1 U15458 ( .A1(n13595), .A2(n13667), .ZN(n13413) );
  NOR2_X1 U15459 ( .A1(n13759), .A2(n13589), .ZN(n13406) );
  AOI211_X1 U15460 ( .C1(n13595), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13413), 
        .B(n13406), .ZN(n13407) );
  OAI21_X1 U15461 ( .B1(n13664), .B2(n13659), .A(n13407), .ZN(P2_U3234) );
  NAND2_X1 U15462 ( .A1(n13411), .A2(n13408), .ZN(n13409) );
  NAND3_X1 U15463 ( .A1(n13410), .A2(n13521), .A3(n13409), .ZN(n13668) );
  INV_X1 U15464 ( .A(n13411), .ZN(n13763) );
  NOR2_X1 U15465 ( .A1(n13763), .A2(n13589), .ZN(n13412) );
  AOI211_X1 U15466 ( .C1(n13595), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13413), 
        .B(n13412), .ZN(n13414) );
  OAI21_X1 U15467 ( .B1(n13659), .B2(n13668), .A(n13414), .ZN(P2_U3235) );
  XNOR2_X1 U15468 ( .A(n13416), .B(n13415), .ZN(n13681) );
  AOI211_X1 U15469 ( .C1(n13680), .C2(n6763), .A(n13221), .B(n13417), .ZN(
        n13679) );
  NOR2_X1 U15470 ( .A1(n13418), .A2(n13589), .ZN(n13422) );
  OAI22_X1 U15471 ( .A1(n13642), .A2(n13420), .B1(n13419), .B2(n13639), .ZN(
        n13421) );
  AOI211_X1 U15472 ( .C1(n13679), .C2(n13646), .A(n13422), .B(n13421), .ZN(
        n13431) );
  NAND2_X1 U15473 ( .A1(n13423), .A2(n13625), .ZN(n13429) );
  AOI21_X1 U15474 ( .B1(n13433), .B2(n13425), .A(n13424), .ZN(n13428) );
  AOI22_X1 U15475 ( .A1(n13466), .A2(n13426), .B1(n13459), .B2(n13628), .ZN(
        n13427) );
  OAI21_X1 U15476 ( .B1(n13429), .B2(n13428), .A(n13427), .ZN(n13678) );
  NAND2_X1 U15477 ( .A1(n13678), .A2(n13642), .ZN(n13430) );
  OAI211_X1 U15478 ( .C1(n13681), .C2(n13636), .A(n13431), .B(n13430), .ZN(
        P2_U3237) );
  INV_X1 U15479 ( .A(n13432), .ZN(n13435) );
  INV_X1 U15480 ( .A(n13682), .ZN(n13448) );
  XNOR2_X1 U15481 ( .A(n13439), .B(n13438), .ZN(n13684) );
  NAND2_X1 U15482 ( .A1(n13684), .A2(n13656), .ZN(n13447) );
  INV_X1 U15483 ( .A(n13450), .ZN(n13441) );
  AOI211_X1 U15484 ( .C1(n6764), .C2(n13441), .A(n13221), .B(n13440), .ZN(
        n13683) );
  NOR2_X1 U15485 ( .A1(n13769), .A2(n13589), .ZN(n13445) );
  OAI22_X1 U15486 ( .A1(n13642), .A2(n13443), .B1(n13442), .B2(n13639), .ZN(
        n13444) );
  AOI211_X1 U15487 ( .C1(n13683), .C2(n13646), .A(n13445), .B(n13444), .ZN(
        n13446) );
  OAI211_X1 U15488 ( .C1(n13595), .C2(n13448), .A(n13447), .B(n13446), .ZN(
        P2_U3238) );
  XNOR2_X1 U15489 ( .A(n13449), .B(n13457), .ZN(n13691) );
  AOI211_X1 U15490 ( .C1(n13688), .C2(n13472), .A(n13221), .B(n13450), .ZN(
        n13687) );
  INV_X1 U15491 ( .A(n13451), .ZN(n13452) );
  AOI22_X1 U15492 ( .A1(n13595), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n13452), 
        .B2(n13654), .ZN(n13453) );
  OAI21_X1 U15493 ( .B1(n13454), .B2(n13589), .A(n13453), .ZN(n13462) );
  OAI21_X1 U15494 ( .B1(n13457), .B2(n13456), .A(n13455), .ZN(n13460) );
  AOI222_X1 U15495 ( .A1(n13625), .A2(n13460), .B1(n13459), .B2(n13466), .C1(
        n13458), .C2(n13628), .ZN(n13690) );
  NOR2_X1 U15496 ( .A1(n13690), .A2(n13595), .ZN(n13461) );
  AOI211_X1 U15497 ( .C1(n13687), .C2(n13646), .A(n13462), .B(n13461), .ZN(
        n13463) );
  OAI21_X1 U15498 ( .B1(n13691), .B2(n13636), .A(n13463), .ZN(P2_U3239) );
  OAI21_X1 U15499 ( .B1(n13470), .B2(n13465), .A(n13464), .ZN(n13469) );
  XNOR2_X1 U15500 ( .A(n13471), .B(n13470), .ZN(n13695) );
  NAND2_X1 U15501 ( .A1(n13695), .A2(n13656), .ZN(n13481) );
  INV_X1 U15502 ( .A(n13490), .ZN(n13474) );
  INV_X1 U15503 ( .A(n13472), .ZN(n13473) );
  AOI211_X1 U15504 ( .C1(n13475), .C2(n13474), .A(n13221), .B(n13473), .ZN(
        n13694) );
  NOR2_X1 U15505 ( .A1(n13773), .A2(n13589), .ZN(n13479) );
  OAI22_X1 U15506 ( .A1(n13642), .A2(n13477), .B1(n13476), .B2(n13639), .ZN(
        n13478) );
  AOI211_X1 U15507 ( .C1(n13694), .C2(n13646), .A(n13479), .B(n13478), .ZN(
        n13480) );
  OAI211_X1 U15508 ( .C1(n13595), .C2(n13692), .A(n13481), .B(n13480), .ZN(
        P2_U3240) );
  NAND2_X1 U15509 ( .A1(n13482), .A2(n13495), .ZN(n13483) );
  NAND2_X1 U15510 ( .A1(n13484), .A2(n13483), .ZN(n13485) );
  NAND2_X1 U15511 ( .A1(n13485), .A2(n13625), .ZN(n13702) );
  OAI211_X1 U15512 ( .C1(n13639), .C2(n13487), .A(n13702), .B(n13486), .ZN(
        n13499) );
  NAND2_X1 U15513 ( .A1(n13700), .A2(n13505), .ZN(n13488) );
  NAND2_X1 U15514 ( .A1(n13488), .A2(n13521), .ZN(n13489) );
  OR2_X1 U15515 ( .A1(n13490), .A2(n13489), .ZN(n13701) );
  NOR2_X1 U15516 ( .A1(n13642), .A2(n13491), .ZN(n13492) );
  AOI21_X1 U15517 ( .B1(n13700), .B2(n13655), .A(n13492), .ZN(n13493) );
  OAI21_X1 U15518 ( .B1(n13701), .B2(n13659), .A(n13493), .ZN(n13498) );
  OAI21_X1 U15519 ( .B1(n13496), .B2(n13495), .A(n13494), .ZN(n13698) );
  NOR2_X1 U15520 ( .A1(n13698), .A2(n13636), .ZN(n13497) );
  AOI211_X1 U15521 ( .C1(n13642), .C2(n13499), .A(n13498), .B(n13497), .ZN(
        n13500) );
  INV_X1 U15522 ( .A(n13500), .ZN(P2_U3241) );
  INV_X1 U15523 ( .A(n13501), .ZN(n13504) );
  XNOR2_X1 U15524 ( .A(n13502), .B(n13509), .ZN(n13503) );
  NOR2_X1 U15525 ( .A1(n13503), .A2(n13603), .ZN(n13708) );
  AOI211_X1 U15526 ( .C1(n13654), .C2(n13504), .A(n13706), .B(n13708), .ZN(
        n13514) );
  INV_X1 U15527 ( .A(n13505), .ZN(n13506) );
  AOI211_X1 U15528 ( .C1(n13507), .C2(n13522), .A(n13221), .B(n13506), .ZN(
        n13707) );
  OAI22_X1 U15529 ( .A1(n6766), .A2(n13589), .B1(n13508), .B2(n13642), .ZN(
        n13512) );
  XNOR2_X1 U15530 ( .A(n13510), .B(n13509), .ZN(n13705) );
  NOR2_X1 U15531 ( .A1(n13705), .A2(n13636), .ZN(n13511) );
  AOI211_X1 U15532 ( .C1(n13707), .C2(n13646), .A(n13512), .B(n13511), .ZN(
        n13513) );
  OAI21_X1 U15533 ( .B1(n13595), .B2(n13514), .A(n13513), .ZN(P2_U3242) );
  XNOR2_X1 U15534 ( .A(n13515), .B(n13520), .ZN(n13516) );
  OAI222_X1 U15535 ( .A1(n13631), .A2(n13518), .B1(n13575), .B2(n13517), .C1(
        n13516), .C2(n13603), .ZN(n13715) );
  INV_X1 U15536 ( .A(n13715), .ZN(n13530) );
  AOI21_X1 U15537 ( .B1(n13520), .B2(n13519), .A(n6547), .ZN(n13716) );
  OAI211_X1 U15538 ( .C1(n6508), .C2(n13713), .A(n13522), .B(n13521), .ZN(
        n13712) );
  OAI22_X1 U15539 ( .A1(n13642), .A2(n13524), .B1(n13523), .B2(n13639), .ZN(
        n13525) );
  AOI21_X1 U15540 ( .B1(n13526), .B2(n13655), .A(n13525), .ZN(n13527) );
  OAI21_X1 U15541 ( .B1(n13712), .B2(n13659), .A(n13527), .ZN(n13528) );
  AOI21_X1 U15542 ( .B1(n13716), .B2(n13656), .A(n13528), .ZN(n13529) );
  OAI21_X1 U15543 ( .B1(n13595), .B2(n13530), .A(n13529), .ZN(P2_U3243) );
  XNOR2_X1 U15544 ( .A(n13531), .B(n13535), .ZN(n13720) );
  NAND2_X1 U15545 ( .A1(n13720), .A2(n13656), .ZN(n13545) );
  INV_X1 U15546 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13533) );
  OAI22_X1 U15547 ( .A1(n13642), .A2(n13533), .B1(n13532), .B2(n13639), .ZN(
        n13534) );
  AOI21_X1 U15548 ( .B1(n13539), .B2(n13655), .A(n13534), .ZN(n13544) );
  XOR2_X1 U15549 ( .A(n13536), .B(n13535), .Z(n13538) );
  OAI21_X1 U15550 ( .B1(n13538), .B2(n13603), .A(n13537), .ZN(n13718) );
  NAND2_X1 U15551 ( .A1(n13718), .A2(n13642), .ZN(n13543) );
  NAND2_X1 U15552 ( .A1(n13555), .A2(n13539), .ZN(n13540) );
  NAND2_X1 U15553 ( .A1(n13540), .A2(n13521), .ZN(n13541) );
  NOR2_X1 U15554 ( .A1(n6508), .A2(n13541), .ZN(n13719) );
  NAND2_X1 U15555 ( .A1(n13719), .A2(n13646), .ZN(n13542) );
  NAND4_X1 U15556 ( .A1(n13545), .A2(n13544), .A3(n13543), .A4(n13542), .ZN(
        P2_U3244) );
  XNOR2_X1 U15557 ( .A(n13546), .B(n13549), .ZN(n13548) );
  AOI21_X1 U15558 ( .B1(n13548), .B2(n13625), .A(n13547), .ZN(n13726) );
  XNOR2_X1 U15559 ( .A(n13550), .B(n13549), .ZN(n13727) );
  INV_X1 U15560 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13552) );
  OAI22_X1 U15561 ( .A1(n13642), .A2(n13552), .B1(n13551), .B2(n13639), .ZN(
        n13553) );
  AOI21_X1 U15562 ( .B1(n13724), .B2(n13655), .A(n13553), .ZN(n13558) );
  INV_X1 U15563 ( .A(n13554), .ZN(n13566) );
  AOI21_X1 U15564 ( .B1(n13566), .B2(n13724), .A(n9793), .ZN(n13556) );
  AND2_X1 U15565 ( .A1(n13556), .A2(n13555), .ZN(n13723) );
  NAND2_X1 U15566 ( .A1(n13723), .A2(n13646), .ZN(n13557) );
  OAI211_X1 U15567 ( .C1(n13727), .C2(n13636), .A(n13558), .B(n13557), .ZN(
        n13559) );
  INV_X1 U15568 ( .A(n13559), .ZN(n13560) );
  OAI21_X1 U15569 ( .B1(n13595), .B2(n13726), .A(n13560), .ZN(P2_U3245) );
  XOR2_X1 U15570 ( .A(n13562), .B(n13561), .Z(n13731) );
  XNOR2_X1 U15571 ( .A(n13563), .B(n13562), .ZN(n13565) );
  OAI21_X1 U15572 ( .B1(n13565), .B2(n13603), .A(n13564), .ZN(n13728) );
  NAND2_X1 U15573 ( .A1(n13729), .A2(n13646), .ZN(n13570) );
  INV_X1 U15574 ( .A(n13567), .ZN(n13568) );
  AOI22_X1 U15575 ( .A1(n13595), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13568), 
        .B2(n13654), .ZN(n13569) );
  OAI211_X1 U15576 ( .C1(n13571), .C2(n13589), .A(n13570), .B(n13569), .ZN(
        n13572) );
  AOI21_X1 U15577 ( .B1(n13642), .B2(n13728), .A(n13572), .ZN(n13573) );
  OAI21_X1 U15578 ( .B1(n13731), .B2(n13636), .A(n13573), .ZN(P2_U3246) );
  XNOR2_X1 U15579 ( .A(n13574), .B(n13579), .ZN(n13582) );
  OAI22_X1 U15580 ( .A1(n13576), .A2(n13631), .B1(n13632), .B2(n13575), .ZN(
        n13581) );
  AOI21_X1 U15581 ( .B1(n13579), .B2(n13578), .A(n13577), .ZN(n13736) );
  NOR2_X1 U15582 ( .A1(n13736), .A2(n9792), .ZN(n13580) );
  AOI211_X1 U15583 ( .C1(n13625), .C2(n13582), .A(n13581), .B(n13580), .ZN(
        n13735) );
  INV_X1 U15584 ( .A(n13611), .ZN(n13585) );
  INV_X1 U15585 ( .A(n13583), .ZN(n13584) );
  AOI211_X1 U15586 ( .C1(n13733), .C2(n13585), .A(n13221), .B(n13584), .ZN(
        n13732) );
  INV_X1 U15587 ( .A(n13586), .ZN(n13587) );
  AOI22_X1 U15588 ( .A1(n13595), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13587), 
        .B2(n13654), .ZN(n13588) );
  OAI21_X1 U15589 ( .B1(n13590), .B2(n13589), .A(n13588), .ZN(n13593) );
  NOR2_X1 U15590 ( .A1(n13736), .A2(n13591), .ZN(n13592) );
  AOI211_X1 U15591 ( .C1(n13732), .C2(n13646), .A(n13593), .B(n13592), .ZN(
        n13594) );
  OAI21_X1 U15592 ( .B1(n13735), .B2(n13595), .A(n13594), .ZN(P2_U3247) );
  XNOR2_X1 U15593 ( .A(n13596), .B(n13600), .ZN(n13739) );
  NAND2_X1 U15594 ( .A1(n13739), .A2(n13656), .ZN(n13615) );
  OAI22_X1 U15595 ( .A1(n13642), .A2(n13598), .B1(n13597), .B2(n13639), .ZN(
        n13599) );
  AOI21_X1 U15596 ( .B1(n13608), .B2(n13655), .A(n13599), .ZN(n13614) );
  INV_X1 U15597 ( .A(n13624), .ZN(n13602) );
  OAI21_X1 U15598 ( .B1(n13602), .B2(n13601), .A(n13600), .ZN(n13605) );
  AOI21_X1 U15599 ( .B1(n13605), .B2(n13604), .A(n13603), .ZN(n13607) );
  NAND2_X1 U15600 ( .A1(n13737), .A2(n13642), .ZN(n13613) );
  NAND2_X1 U15601 ( .A1(n13608), .A2(n13620), .ZN(n13609) );
  NAND2_X1 U15602 ( .A1(n13609), .A2(n13521), .ZN(n13610) );
  NOR2_X1 U15603 ( .A1(n13611), .A2(n13610), .ZN(n13738) );
  NAND2_X1 U15604 ( .A1(n13738), .A2(n13646), .ZN(n13612) );
  NAND4_X1 U15605 ( .A1(n13615), .A2(n13614), .A3(n13613), .A4(n13612), .ZN(
        P2_U3248) );
  XNOR2_X1 U15606 ( .A(n6588), .B(n13626), .ZN(n13742) );
  INV_X1 U15607 ( .A(n13742), .ZN(n13637) );
  OAI22_X1 U15608 ( .A1(n13642), .A2(n13617), .B1(n13616), .B2(n13639), .ZN(
        n13623) );
  AOI21_X1 U15609 ( .B1(n13744), .B2(n13619), .A(n9793), .ZN(n13621) );
  NAND2_X1 U15610 ( .A1(n13621), .A2(n13620), .ZN(n13745) );
  NOR2_X1 U15611 ( .A1(n13745), .A2(n13659), .ZN(n13622) );
  AOI211_X1 U15612 ( .C1(n13655), .C2(n13744), .A(n13623), .B(n13622), .ZN(
        n13635) );
  OAI211_X1 U15613 ( .C1(n13627), .C2(n13626), .A(n13625), .B(n13624), .ZN(
        n13746) );
  INV_X1 U15614 ( .A(n13746), .ZN(n13633) );
  NAND2_X1 U15615 ( .A1(n13629), .A2(n13628), .ZN(n13630) );
  OAI21_X1 U15616 ( .B1(n13632), .B2(n13631), .A(n13630), .ZN(n13743) );
  OAI21_X1 U15617 ( .B1(n13633), .B2(n13743), .A(n13642), .ZN(n13634) );
  OAI211_X1 U15618 ( .C1(n13637), .C2(n13636), .A(n13635), .B(n13634), .ZN(
        P2_U3249) );
  NAND2_X1 U15619 ( .A1(n13638), .A2(n13656), .ZN(n13651) );
  OAI22_X1 U15620 ( .A1(n13642), .A2(n13641), .B1(n13640), .B2(n13639), .ZN(
        n13643) );
  AOI21_X1 U15621 ( .B1(n13644), .B2(n13655), .A(n13643), .ZN(n13650) );
  NAND2_X1 U15622 ( .A1(n13645), .A2(n13642), .ZN(n13649) );
  NAND2_X1 U15623 ( .A1(n13647), .A2(n13646), .ZN(n13648) );
  NAND4_X1 U15624 ( .A1(n13651), .A2(n13650), .A3(n13649), .A4(n13648), .ZN(
        P2_U3252) );
  MUX2_X1 U15625 ( .A(n13653), .B(n13652), .S(n13642), .Z(n13663) );
  AOI22_X1 U15626 ( .A1(n13655), .A2(n9108), .B1(n15241), .B2(n13654), .ZN(
        n13662) );
  NAND2_X1 U15627 ( .A1(n13657), .A2(n13656), .ZN(n13661) );
  OR2_X1 U15628 ( .A1(n13659), .A2(n13658), .ZN(n13660) );
  NAND4_X1 U15629 ( .A1(n13663), .A2(n13662), .A3(n13661), .A4(n13660), .ZN(
        P2_U3262) );
  INV_X1 U15630 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13665) );
  MUX2_X1 U15631 ( .A(n13665), .B(n13756), .S(n14986), .Z(n13666) );
  OAI21_X1 U15632 ( .B1(n13759), .B2(n13755), .A(n13666), .ZN(P2_U3530) );
  INV_X1 U15633 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13669) );
  AND2_X1 U15634 ( .A1(n13668), .A2(n13667), .ZN(n13760) );
  MUX2_X1 U15635 ( .A(n13669), .B(n13760), .S(n14986), .Z(n13670) );
  OAI21_X1 U15636 ( .B1(n13763), .B2(n13755), .A(n13670), .ZN(P2_U3529) );
  NAND2_X1 U15637 ( .A1(n13671), .A2(n14951), .ZN(n13677) );
  NAND2_X1 U15638 ( .A1(n13672), .A2(n14939), .ZN(n13673) );
  MUX2_X1 U15639 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13764), .S(n14986), .Z(
        P2_U3528) );
  MUX2_X1 U15640 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13765), .S(n14986), .Z(
        P2_U3527) );
  MUX2_X1 U15641 ( .A(n13685), .B(n13766), .S(n14986), .Z(n13686) );
  OAI21_X1 U15642 ( .B1(n13769), .B2(n13755), .A(n13686), .ZN(P2_U3526) );
  AOI21_X1 U15643 ( .B1(n14939), .B2(n13688), .A(n13687), .ZN(n13689) );
  OAI211_X1 U15644 ( .C1(n13691), .C2(n13751), .A(n13690), .B(n13689), .ZN(
        n13770) );
  MUX2_X1 U15645 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13770), .S(n14986), .Z(
        P2_U3525) );
  INV_X1 U15646 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13696) );
  INV_X1 U15647 ( .A(n13692), .ZN(n13693) );
  MUX2_X1 U15648 ( .A(n13696), .B(n13771), .S(n14986), .Z(n13697) );
  OAI21_X1 U15649 ( .B1(n13773), .B2(n13755), .A(n13697), .ZN(P2_U3524) );
  OR2_X1 U15650 ( .A1(n13698), .A2(n13751), .ZN(n13704) );
  AOI21_X1 U15651 ( .B1(n13700), .B2(n14939), .A(n13699), .ZN(n13703) );
  NAND4_X1 U15652 ( .A1(n13704), .A2(n13703), .A3(n13702), .A4(n13701), .ZN(
        n13774) );
  MUX2_X1 U15653 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13774), .S(n14986), .Z(
        P2_U3523) );
  INV_X1 U15654 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n13710) );
  NOR2_X1 U15655 ( .A1(n13705), .A2(n13751), .ZN(n13709) );
  NOR4_X1 U15656 ( .A1(n13709), .A2(n13708), .A3(n13707), .A4(n13706), .ZN(
        n13775) );
  MUX2_X1 U15657 ( .A(n13710), .B(n13775), .S(n14986), .Z(n13711) );
  OAI21_X1 U15658 ( .B1(n6766), .B2(n13755), .A(n13711), .ZN(P2_U3522) );
  OAI21_X1 U15659 ( .B1(n13713), .B2(n14967), .A(n13712), .ZN(n13714) );
  AOI211_X1 U15660 ( .C1(n13716), .C2(n14951), .A(n13715), .B(n13714), .ZN(
        n13717) );
  INV_X1 U15661 ( .A(n13717), .ZN(n13778) );
  MUX2_X1 U15662 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13778), .S(n14986), .Z(
        P2_U3521) );
  INV_X1 U15663 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13721) );
  AOI211_X1 U15664 ( .C1(n13720), .C2(n14951), .A(n13719), .B(n13718), .ZN(
        n13779) );
  MUX2_X1 U15665 ( .A(n13721), .B(n13779), .S(n14986), .Z(n13722) );
  OAI21_X1 U15666 ( .B1(n13782), .B2(n13755), .A(n13722), .ZN(P2_U3520) );
  AOI21_X1 U15667 ( .B1(n14939), .B2(n13724), .A(n13723), .ZN(n13725) );
  OAI211_X1 U15668 ( .C1(n13727), .C2(n13751), .A(n13726), .B(n13725), .ZN(
        n13783) );
  MUX2_X1 U15669 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13783), .S(n14986), .Z(
        P2_U3519) );
  OAI21_X1 U15670 ( .B1(n13731), .B2(n13751), .A(n13730), .ZN(n13784) );
  MUX2_X1 U15671 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13784), .S(n14986), .Z(
        P2_U3518) );
  AOI21_X1 U15672 ( .B1(n14939), .B2(n13733), .A(n13732), .ZN(n13734) );
  OAI211_X1 U15673 ( .C1(n13736), .C2(n14942), .A(n13735), .B(n13734), .ZN(
        n13785) );
  MUX2_X1 U15674 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13785), .S(n14986), .Z(
        P2_U3517) );
  INV_X1 U15675 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13740) );
  AOI211_X1 U15676 ( .C1(n13739), .C2(n14951), .A(n13738), .B(n13737), .ZN(
        n13786) );
  MUX2_X1 U15677 ( .A(n13740), .B(n13786), .S(n14986), .Z(n13741) );
  OAI21_X1 U15678 ( .B1(n13789), .B2(n13755), .A(n13741), .ZN(P2_U3516) );
  NAND2_X1 U15679 ( .A1(n13742), .A2(n14951), .ZN(n13748) );
  AOI21_X1 U15680 ( .B1(n13744), .B2(n14939), .A(n13743), .ZN(n13747) );
  NAND4_X1 U15681 ( .A1(n13748), .A2(n13747), .A3(n13746), .A4(n13745), .ZN(
        n13790) );
  MUX2_X1 U15682 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13790), .S(n14986), .Z(
        P2_U3515) );
  OAI211_X1 U15683 ( .C1(n13752), .C2(n13751), .A(n13750), .B(n13749), .ZN(
        n13753) );
  INV_X1 U15684 ( .A(n13753), .ZN(n13791) );
  MUX2_X1 U15685 ( .A(n15131), .B(n13791), .S(n14986), .Z(n13754) );
  OAI21_X1 U15686 ( .B1(n13795), .B2(n13755), .A(n13754), .ZN(P2_U3514) );
  MUX2_X1 U15687 ( .A(n13757), .B(n13756), .S(n14974), .Z(n13758) );
  OAI21_X1 U15688 ( .B1(n13759), .B2(n13794), .A(n13758), .ZN(P2_U3498) );
  MUX2_X1 U15689 ( .A(n13761), .B(n13760), .S(n14974), .Z(n13762) );
  OAI21_X1 U15690 ( .B1(n13763), .B2(n13794), .A(n13762), .ZN(P2_U3497) );
  MUX2_X1 U15691 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13764), .S(n14974), .Z(
        P2_U3496) );
  MUX2_X1 U15692 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13765), .S(n14974), .Z(
        P2_U3495) );
  INV_X1 U15693 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13767) );
  MUX2_X1 U15694 ( .A(n13767), .B(n13766), .S(n14974), .Z(n13768) );
  OAI21_X1 U15695 ( .B1(n13769), .B2(n13794), .A(n13768), .ZN(P2_U3494) );
  MUX2_X1 U15696 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13770), .S(n14974), .Z(
        P2_U3493) );
  MUX2_X1 U15697 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13774), .S(n14974), .Z(
        P2_U3491) );
  MUX2_X1 U15698 ( .A(n13776), .B(n13775), .S(n14974), .Z(n13777) );
  OAI21_X1 U15699 ( .B1(n6766), .B2(n13794), .A(n13777), .ZN(P2_U3490) );
  MUX2_X1 U15700 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13778), .S(n14974), .Z(
        P2_U3489) );
  MUX2_X1 U15701 ( .A(n13780), .B(n13779), .S(n14974), .Z(n13781) );
  OAI21_X1 U15702 ( .B1(n13782), .B2(n13794), .A(n13781), .ZN(P2_U3488) );
  MUX2_X1 U15703 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13783), .S(n14974), .Z(
        P2_U3487) );
  MUX2_X1 U15704 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13784), .S(n14974), .Z(
        P2_U3486) );
  MUX2_X1 U15705 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13785), .S(n14974), .Z(
        P2_U3484) );
  MUX2_X1 U15706 ( .A(n13787), .B(n13786), .S(n14974), .Z(n13788) );
  OAI21_X1 U15707 ( .B1(n13789), .B2(n13794), .A(n13788), .ZN(P2_U3481) );
  MUX2_X1 U15708 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13790), .S(n14974), .Z(
        P2_U3478) );
  MUX2_X1 U15709 ( .A(n13792), .B(n13791), .S(n14974), .Z(n13793) );
  OAI21_X1 U15710 ( .B1(n13795), .B2(n13794), .A(n13793), .ZN(P2_U3475) );
  INV_X1 U15711 ( .A(n13796), .ZN(n14392) );
  INV_X1 U15712 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13797) );
  NAND3_X1 U15713 ( .A1(n13797), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13800) );
  OAI22_X1 U15714 ( .A1(n7418), .A2(n13800), .B1(n13799), .B2(n13798), .ZN(
        n13801) );
  INV_X1 U15715 ( .A(n13801), .ZN(n13802) );
  OAI21_X1 U15716 ( .B1(n14392), .B2(n13803), .A(n13802), .ZN(P2_U3296) );
  OAI222_X1 U15717 ( .A1(n13817), .A2(n13806), .B1(P2_U3088), .B2(n13804), 
        .C1(n13805), .C2(n13819), .ZN(P2_U3297) );
  INV_X1 U15718 ( .A(n13807), .ZN(n14395) );
  OAI222_X1 U15719 ( .A1(n13817), .A2(n14395), .B1(P2_U3088), .B2(n13809), 
        .C1(n13808), .C2(n13819), .ZN(P2_U3298) );
  NAND2_X1 U15720 ( .A1(n13811), .A2(n13810), .ZN(n13813) );
  OAI211_X1 U15721 ( .C1(n13819), .C2(n13814), .A(n13813), .B(n13812), .ZN(
        P2_U3299) );
  INV_X1 U15722 ( .A(n13815), .ZN(n14397) );
  OAI222_X1 U15723 ( .A1(n13819), .A2(n13818), .B1(n13817), .B2(n14397), .C1(
        P2_U3088), .C2(n13816), .ZN(P2_U3300) );
  INV_X1 U15724 ( .A(n13820), .ZN(n13821) );
  MUX2_X1 U15725 ( .A(n13821), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  INV_X1 U15726 ( .A(n14310), .ZN(n14091) );
  OAI21_X1 U15727 ( .B1(n13824), .B2(n13823), .A(n13822), .ZN(n13825) );
  AOI22_X1 U15728 ( .A1(n14065), .A2(n6479), .B1(n14064), .B2(n14060), .ZN(
        n14128) );
  OAI22_X1 U15729 ( .A1(n14128), .A2(n13949), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15112), .ZN(n13826) );
  AOI21_X1 U15730 ( .B1(n14136), .B2(n13947), .A(n13826), .ZN(n13827) );
  OAI21_X1 U15731 ( .B1(n13830), .B2(n13829), .A(n13828), .ZN(n13831) );
  NAND2_X1 U15732 ( .A1(n13831), .A2(n13937), .ZN(n13836) );
  OAI21_X1 U15733 ( .B1(n14634), .B2(n13949), .A(n13832), .ZN(n13833) );
  AOI21_X1 U15734 ( .B1(n13834), .B2(n13947), .A(n13833), .ZN(n13835) );
  OAI211_X1 U15735 ( .C1(n14636), .C2(n13943), .A(n13836), .B(n13835), .ZN(
        P1_U3215) );
  INV_X1 U15736 ( .A(n14332), .ZN(n13846) );
  INV_X1 U15737 ( .A(n13837), .ZN(n13894) );
  NOR3_X1 U15738 ( .A1(n13915), .A2(n13839), .A3(n13838), .ZN(n13840) );
  OAI21_X1 U15739 ( .B1(n13894), .B2(n13840), .A(n13937), .ZN(n13845) );
  OAI22_X1 U15740 ( .A1(n13858), .A2(n13917), .B1(n14059), .B2(n13916), .ZN(
        n14193) );
  INV_X1 U15741 ( .A(n13841), .ZN(n14198) );
  OAI22_X1 U15742 ( .A1(n13920), .A2(n14198), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13842), .ZN(n13843) );
  AOI21_X1 U15743 ( .B1(n14193), .B2(n13923), .A(n13843), .ZN(n13844) );
  OAI211_X1 U15744 ( .C1(n13846), .C2(n13943), .A(n13845), .B(n13844), .ZN(
        P1_U3216) );
  INV_X1 U15745 ( .A(n12379), .ZN(n14259) );
  AND2_X1 U15746 ( .A1(n13926), .A2(n13847), .ZN(n13850) );
  OAI211_X1 U15747 ( .C1(n13850), .C2(n13849), .A(n13937), .B(n13848), .ZN(
        n13854) );
  OAI22_X1 U15748 ( .A1(n14077), .A2(n13916), .B1(n13851), .B2(n13917), .ZN(
        n14358) );
  NAND2_X1 U15749 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14031)
         );
  OAI21_X1 U15750 ( .B1(n13920), .B2(n14253), .A(n14031), .ZN(n13852) );
  AOI21_X1 U15751 ( .B1(n14358), .B2(n13923), .A(n13852), .ZN(n13853) );
  OAI211_X1 U15752 ( .C1(n14259), .C2(n13943), .A(n13854), .B(n13853), .ZN(
        P1_U3219) );
  INV_X1 U15753 ( .A(n14346), .ZN(n14228) );
  OAI21_X1 U15754 ( .B1(n13856), .B2(n13855), .A(n13913), .ZN(n13857) );
  NAND2_X1 U15755 ( .A1(n13857), .A2(n13937), .ZN(n13862) );
  OAI22_X1 U15756 ( .A1(n13858), .A2(n13916), .B1(n14077), .B2(n13917), .ZN(
        n14345) );
  OAI22_X1 U15757 ( .A1(n14224), .A2(n13920), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13859), .ZN(n13860) );
  AOI21_X1 U15758 ( .B1(n14345), .B2(n13923), .A(n13860), .ZN(n13861) );
  OAI211_X1 U15759 ( .C1(n14228), .C2(n13943), .A(n13862), .B(n13861), .ZN(
        P1_U3223) );
  INV_X1 U15760 ( .A(n14320), .ZN(n14088) );
  INV_X1 U15761 ( .A(n13863), .ZN(n13895) );
  INV_X1 U15762 ( .A(n13864), .ZN(n13866) );
  NOR3_X1 U15763 ( .A1(n13895), .A2(n13866), .A3(n13865), .ZN(n13869) );
  INV_X1 U15764 ( .A(n13867), .ZN(n13868) );
  OAI21_X1 U15765 ( .B1(n13869), .B2(n13868), .A(n13937), .ZN(n13873) );
  AOI22_X1 U15766 ( .A1(n14064), .A2(n14086), .B1(n14060), .B2(n6479), .ZN(
        n14163) );
  INV_X1 U15767 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13870) );
  OAI22_X1 U15768 ( .A1(n13949), .A2(n14163), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13870), .ZN(n13871) );
  AOI21_X1 U15769 ( .B1(n14169), .B2(n13947), .A(n13871), .ZN(n13872) );
  OAI211_X1 U15770 ( .C1(n14088), .C2(n13943), .A(n13873), .B(n13872), .ZN(
        P1_U3225) );
  AOI21_X1 U15771 ( .B1(n13875), .B2(n13874), .A(n6527), .ZN(n13880) );
  NOR2_X1 U15772 ( .A1(n13920), .A2(n14604), .ZN(n13878) );
  AOI22_X1 U15773 ( .A1(n14047), .A2(n6479), .B1(n13962), .B2(n14064), .ZN(
        n14614) );
  OAI21_X1 U15774 ( .B1(n14614), .B2(n13949), .A(n13876), .ZN(n13877) );
  AOI211_X1 U15775 ( .C1(n14607), .C2(n13952), .A(n13878), .B(n13877), .ZN(
        n13879) );
  OAI21_X1 U15776 ( .B1(n13880), .B2(n13955), .A(n13879), .ZN(P1_U3226) );
  INV_X1 U15777 ( .A(n13881), .ZN(n13885) );
  NOR3_X1 U15778 ( .A1(n6527), .A2(n13883), .A3(n13882), .ZN(n13884) );
  OAI21_X1 U15779 ( .B1(n13885), .B2(n13884), .A(n13937), .ZN(n13890) );
  AND2_X1 U15780 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13985) );
  NOR2_X1 U15781 ( .A1(n13920), .A2(n13886), .ZN(n13887) );
  AOI211_X1 U15782 ( .C1(n13923), .C2(n13888), .A(n13985), .B(n13887), .ZN(
        n13889) );
  OAI211_X1 U15783 ( .C1(n14619), .C2(n13943), .A(n13890), .B(n13889), .ZN(
        P1_U3228) );
  INV_X1 U15784 ( .A(n14327), .ZN(n14188) );
  INV_X1 U15785 ( .A(n13891), .ZN(n13893) );
  NOR3_X1 U15786 ( .A1(n13894), .A2(n13893), .A3(n13892), .ZN(n13896) );
  OAI21_X1 U15787 ( .B1(n13896), .B2(n13895), .A(n13937), .ZN(n13900) );
  AOI22_X1 U15788 ( .A1(n14064), .A2(n14084), .B1(n13960), .B2(n6479), .ZN(
        n14179) );
  OAI22_X1 U15789 ( .A1(n13949), .A2(n14179), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13897), .ZN(n13898) );
  AOI21_X1 U15790 ( .B1(n14185), .B2(n13947), .A(n13898), .ZN(n13899) );
  OAI211_X1 U15791 ( .C1(n14188), .C2(n13943), .A(n13900), .B(n13899), .ZN(
        P1_U3229) );
  XOR2_X1 U15792 ( .A(n13901), .B(n13902), .Z(n13903) );
  NAND2_X1 U15793 ( .A1(n13903), .A2(n13937), .ZN(n13910) );
  NAND2_X1 U15794 ( .A1(n14079), .A2(n6479), .ZN(n13906) );
  NAND2_X1 U15795 ( .A1(n14074), .A2(n14064), .ZN(n13905) );
  NAND2_X1 U15796 ( .A1(n13906), .A2(n13905), .ZN(n14234) );
  OAI22_X1 U15797 ( .A1(n13920), .A2(n14238), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13907), .ZN(n13908) );
  AOI21_X1 U15798 ( .B1(n14234), .B2(n13923), .A(n13908), .ZN(n13909) );
  OAI211_X1 U15799 ( .C1(n14241), .C2(n13943), .A(n13910), .B(n13909), .ZN(
        P1_U3233) );
  AND3_X1 U15800 ( .A1(n13913), .A2(n13912), .A3(n13911), .ZN(n13914) );
  OAI21_X1 U15801 ( .B1(n13915), .B2(n13914), .A(n13937), .ZN(n13925) );
  INV_X1 U15802 ( .A(n14084), .ZN(n14057) );
  OAI22_X1 U15803 ( .A1(n13918), .A2(n13917), .B1(n14057), .B2(n13916), .ZN(
        n14338) );
  INV_X1 U15804 ( .A(n14211), .ZN(n13921) );
  INV_X1 U15805 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13919) );
  OAI22_X1 U15806 ( .A1(n13921), .A2(n13920), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13919), .ZN(n13922) );
  AOI21_X1 U15807 ( .B1(n14338), .B2(n13923), .A(n13922), .ZN(n13924) );
  OAI211_X1 U15808 ( .C1(n13943), .C2(n7153), .A(n13925), .B(n13924), .ZN(
        P1_U3235) );
  OAI21_X1 U15809 ( .B1(n13928), .B2(n13927), .A(n13926), .ZN(n13929) );
  NAND2_X1 U15810 ( .A1(n13929), .A2(n13937), .ZN(n13933) );
  AND2_X1 U15811 ( .A1(n14047), .A2(n14064), .ZN(n13930) );
  AOI21_X1 U15812 ( .B1(n14074), .B2(n6479), .A(n13930), .ZN(n14364) );
  NAND2_X1 U15813 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13997)
         );
  OAI21_X1 U15814 ( .B1(n14364), .B2(n13949), .A(n13997), .ZN(n13931) );
  AOI21_X1 U15815 ( .B1(n14266), .B2(n13947), .A(n13931), .ZN(n13932) );
  OAI211_X1 U15816 ( .C1(n14366), .C2(n13943), .A(n13933), .B(n13932), .ZN(
        P1_U3238) );
  OAI21_X1 U15817 ( .B1(n13936), .B2(n13935), .A(n13934), .ZN(n13938) );
  NAND2_X1 U15818 ( .A1(n13938), .A2(n13937), .ZN(n13942) );
  AOI22_X1 U15819 ( .A1(n14064), .A2(n13960), .B1(n13959), .B2(n6479), .ZN(
        n14146) );
  OAI22_X1 U15820 ( .A1(n13949), .A2(n14146), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13939), .ZN(n13940) );
  AOI21_X1 U15821 ( .B1(n14154), .B2(n13947), .A(n13940), .ZN(n13941) );
  OAI211_X1 U15822 ( .C1(n14156), .C2(n13943), .A(n13942), .B(n13941), .ZN(
        P1_U3240) );
  XNOR2_X1 U15823 ( .A(n13944), .B(n13945), .ZN(n13956) );
  NAND2_X1 U15824 ( .A1(n13947), .A2(n13946), .ZN(n13948) );
  NAND2_X1 U15825 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14689)
         );
  OAI211_X1 U15826 ( .C1(n13950), .C2(n13949), .A(n13948), .B(n14689), .ZN(
        n13951) );
  AOI21_X1 U15827 ( .B1(n13953), .B2(n13952), .A(n13951), .ZN(n13954) );
  OAI21_X1 U15828 ( .B1(n13956), .B2(n13955), .A(n13954), .ZN(P1_U3241) );
  MUX2_X1 U15829 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13957), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15830 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14099), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15831 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13958), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15832 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14065), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15833 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13959), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15834 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14060), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15835 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13960), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15836 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14086), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15837 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14084), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15838 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14082), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15839 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14079), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15840 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14054), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15841 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14074), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15842 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14051), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15843 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14047), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15844 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13961), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15845 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13962), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15846 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13963), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15847 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13964), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15848 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13965), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15849 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13966), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15850 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13967), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15851 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13968), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15852 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13969), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15853 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13970), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15854 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13971), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15855 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13972), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15856 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13973), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15857 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13974), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15858 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13975), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15859 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13976), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15860 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n13977), .S(P1_U4016), .Z(
        P1_U3560) );
  INV_X1 U15861 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14623) );
  NOR2_X1 U15862 ( .A1(n14004), .A2(n14623), .ZN(n13979) );
  AOI21_X1 U15863 ( .B1(n14004), .B2(n14623), .A(n13979), .ZN(n13981) );
  AOI211_X1 U15864 ( .C1(n13982), .C2(n13981), .A(n14003), .B(n13980), .ZN(
        n13983) );
  INV_X1 U15865 ( .A(n13983), .ZN(n13996) );
  NOR2_X1 U15866 ( .A1(n14023), .A2(n14001), .ZN(n13984) );
  AOI211_X1 U15867 ( .C1(n13986), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n13985), 
        .B(n13984), .ZN(n13995) );
  NOR2_X1 U15868 ( .A1(n14001), .A2(n13987), .ZN(n13988) );
  AOI21_X1 U15869 ( .B1(n13987), .B2(n14001), .A(n13988), .ZN(n13993) );
  INV_X1 U15870 ( .A(n13989), .ZN(n13991) );
  OAI21_X1 U15871 ( .B1(n13991), .B2(n11750), .A(n13990), .ZN(n13992) );
  NAND2_X1 U15872 ( .A1(n13993), .A2(n13992), .ZN(n14000) );
  OAI211_X1 U15873 ( .C1(n13993), .C2(n13992), .A(n14027), .B(n14000), .ZN(
        n13994) );
  NAND3_X1 U15874 ( .A1(n13996), .A2(n13995), .A3(n13994), .ZN(P1_U3260) );
  INV_X1 U15875 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n13998) );
  OAI21_X1 U15876 ( .B1(n14691), .B2(n13998), .A(n13997), .ZN(n13999) );
  AOI21_X1 U15877 ( .B1(n14683), .B2(n14019), .A(n13999), .ZN(n14011) );
  OAI21_X1 U15878 ( .B1(n13987), .B2(n14001), .A(n14000), .ZN(n14018) );
  XNOR2_X1 U15879 ( .A(n14012), .B(n14018), .ZN(n14002) );
  NAND2_X1 U15880 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14002), .ZN(n14021) );
  OAI211_X1 U15881 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14002), .A(n14027), 
        .B(n14021), .ZN(n14010) );
  INV_X1 U15882 ( .A(n14005), .ZN(n14008) );
  INV_X1 U15883 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14006) );
  NOR2_X1 U15884 ( .A1(n14006), .A2(n14005), .ZN(n14015) );
  INV_X1 U15885 ( .A(n14015), .ZN(n14007) );
  OAI211_X1 U15886 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n14008), .A(n14680), 
        .B(n14007), .ZN(n14009) );
  NAND3_X1 U15887 ( .A1(n14011), .A2(n14010), .A3(n14009), .ZN(P1_U3261) );
  NOR2_X1 U15888 ( .A1(n14013), .A2(n14012), .ZN(n14014) );
  NOR2_X1 U15889 ( .A1(n14015), .A2(n14014), .ZN(n14017) );
  XOR2_X1 U15890 ( .A(n14017), .B(n14016), .Z(n14028) );
  INV_X1 U15891 ( .A(n14028), .ZN(n14025) );
  NAND2_X1 U15892 ( .A1(n14019), .A2(n14018), .ZN(n14020) );
  NAND2_X1 U15893 ( .A1(n14021), .A2(n14020), .ZN(n14022) );
  XOR2_X1 U15894 ( .A(n14022), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14026) );
  OAI21_X1 U15895 ( .B1(n14026), .B2(n14686), .A(n14023), .ZN(n14024) );
  AOI21_X1 U15896 ( .B1(n14025), .B2(n14680), .A(n14024), .ZN(n14030) );
  AOI22_X1 U15897 ( .A1(n14028), .A2(n14680), .B1(n14027), .B2(n14026), .ZN(
        n14029) );
  MUX2_X1 U15898 ( .A(n14030), .B(n14029), .S(n14150), .Z(n14032) );
  OAI211_X1 U15899 ( .C1(n14033), .C2(n14691), .A(n14032), .B(n14031), .ZN(
        P1_U3262) );
  NAND2_X1 U15900 ( .A1(n14251), .A2(n14241), .ZN(n14223) );
  NAND2_X1 U15901 ( .A1(n14303), .A2(n14135), .ZN(n14118) );
  OR2_X2 U15902 ( .A1(n14297), .A2(n14118), .ZN(n14096) );
  XNOR2_X1 U15903 ( .A(n14041), .B(n14035), .ZN(n14036) );
  NAND2_X1 U15904 ( .A1(n14036), .A2(n14749), .ZN(n14289) );
  OAI21_X1 U15905 ( .B1(n14398), .B2(n14037), .A(n6479), .ZN(n14100) );
  OR2_X1 U15906 ( .A1(n14038), .A2(n14100), .ZN(n14291) );
  NOR2_X1 U15907 ( .A1(n14724), .A2(n14291), .ZN(n14045) );
  NOR2_X1 U15908 ( .A1(n14290), .A2(n14258), .ZN(n14039) );
  AOI211_X1 U15909 ( .C1(n14724), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14045), 
        .B(n14039), .ZN(n14040) );
  OAI21_X1 U15910 ( .B1(n14289), .B2(n14270), .A(n14040), .ZN(P1_U3263) );
  INV_X1 U15911 ( .A(n14096), .ZN(n14043) );
  INV_X1 U15912 ( .A(n14041), .ZN(n14042) );
  NOR2_X1 U15913 ( .A1(n14293), .A2(n14258), .ZN(n14044) );
  AOI211_X1 U15914 ( .C1(n14724), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14045), 
        .B(n14044), .ZN(n14046) );
  OAI21_X1 U15915 ( .B1(n14270), .B2(n14292), .A(n14046), .ZN(P1_U3264) );
  NAND2_X1 U15916 ( .A1(n14619), .A2(n14047), .ZN(n14048) );
  OAI21_X1 U15917 ( .B1(n14059), .B2(n14327), .A(n14177), .ZN(n14162) );
  NOR2_X1 U15918 ( .A1(n14162), .A2(n14173), .ZN(n14161) );
  NAND2_X1 U15919 ( .A1(n14062), .A2(n14061), .ZN(n14063) );
  AND2_X1 U15920 ( .A1(n14619), .A2(n14067), .ZN(n14068) );
  OAI22_X1 U15921 ( .A1(n14069), .A2(n14068), .B1(n14619), .B2(n14067), .ZN(
        n14263) );
  OR2_X1 U15922 ( .A1(n12379), .A2(n14074), .ZN(n14075) );
  OR2_X1 U15923 ( .A1(n14241), .A2(n14077), .ZN(n14078) );
  NAND2_X1 U15924 ( .A1(n14353), .A2(n14078), .ZN(n14219) );
  OR2_X1 U15925 ( .A1(n14346), .A2(n14079), .ZN(n14080) );
  INV_X1 U15926 ( .A(n14206), .ZN(n14081) );
  NAND2_X1 U15927 ( .A1(n14332), .A2(n14084), .ZN(n14085) );
  NAND2_X1 U15928 ( .A1(n14321), .A2(n7431), .ZN(n14153) );
  NAND2_X1 U15929 ( .A1(n14153), .A2(n14152), .ZN(n14151) );
  INV_X1 U15930 ( .A(n14112), .ZN(n14114) );
  NAND2_X1 U15931 ( .A1(n14117), .A2(n14092), .ZN(n14095) );
  INV_X1 U15932 ( .A(n14093), .ZN(n14094) );
  INV_X1 U15933 ( .A(n14299), .ZN(n14110) );
  INV_X1 U15934 ( .A(n14297), .ZN(n14107) );
  INV_X1 U15935 ( .A(n14118), .ZN(n14097) );
  NOR2_X1 U15936 ( .A1(n14295), .A2(n14098), .ZN(n14109) );
  INV_X1 U15937 ( .A(n14099), .ZN(n14101) );
  NOR2_X1 U15938 ( .A1(n14101), .A2(n14100), .ZN(n14296) );
  INV_X1 U15939 ( .A(n14102), .ZN(n14104) );
  AOI22_X1 U15940 ( .A1(n14296), .A2(n14104), .B1(n14713), .B2(n14103), .ZN(
        n14106) );
  NAND2_X1 U15941 ( .A1(n14724), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n14105) );
  OAI211_X1 U15942 ( .C1(n14107), .C2(n14258), .A(n14106), .B(n14105), .ZN(
        n14108) );
  AOI211_X1 U15943 ( .C1(n14110), .C2(n14703), .A(n14109), .B(n14108), .ZN(
        n14111) );
  OAI21_X1 U15944 ( .B1(n14298), .B2(n14724), .A(n14111), .ZN(P1_U3356) );
  OAI211_X1 U15945 ( .C1(n14303), .C2(n14135), .A(n14749), .B(n14118), .ZN(
        n14302) );
  INV_X1 U15946 ( .A(n14119), .ZN(n14301) );
  OAI22_X1 U15947 ( .A1(n14301), .A2(n14724), .B1(n14120), .B2(n14252), .ZN(
        n14122) );
  NOR2_X1 U15948 ( .A1(n14303), .A2(n14258), .ZN(n14121) );
  AOI211_X1 U15949 ( .C1(n14724), .C2(P1_REG2_REG_28__SCAN_IN), .A(n14122), 
        .B(n14121), .ZN(n14123) );
  OAI21_X1 U15950 ( .B1(n14302), .B2(n14270), .A(n14123), .ZN(n14124) );
  AOI21_X1 U15951 ( .B1(n7445), .B2(n14703), .A(n14124), .ZN(n14125) );
  OAI21_X1 U15952 ( .B1(n14300), .B2(n14126), .A(n14125), .ZN(P1_U3265) );
  XNOR2_X1 U15953 ( .A(n14127), .B(n14133), .ZN(n14130) );
  INV_X1 U15954 ( .A(n14128), .ZN(n14129) );
  AOI21_X1 U15955 ( .B1(n14133), .B2(n14132), .A(n14131), .ZN(n14313) );
  INV_X1 U15956 ( .A(n14313), .ZN(n14140) );
  AND2_X1 U15957 ( .A1(n14310), .A2(n14142), .ZN(n14134) );
  OR3_X1 U15958 ( .A1(n14135), .A2(n14134), .A3(n14294), .ZN(n14308) );
  AOI22_X1 U15959 ( .A1(n14724), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14136), 
        .B2(n14713), .ZN(n14138) );
  NAND2_X1 U15960 ( .A1(n14310), .A2(n14715), .ZN(n14137) );
  OAI211_X1 U15961 ( .C1(n14308), .C2(n14270), .A(n14138), .B(n14137), .ZN(
        n14139) );
  AOI21_X1 U15962 ( .B1(n14140), .B2(n14703), .A(n14139), .ZN(n14141) );
  OAI21_X1 U15963 ( .B1(n14312), .B2(n14724), .A(n14141), .ZN(P1_U3266) );
  INV_X1 U15964 ( .A(n14168), .ZN(n14144) );
  INV_X1 U15965 ( .A(n14142), .ZN(n14143) );
  AOI211_X1 U15966 ( .C1(n14315), .C2(n14144), .A(n14294), .B(n14143), .ZN(
        n14314) );
  XNOR2_X1 U15967 ( .A(n14145), .B(n14152), .ZN(n14148) );
  INV_X1 U15968 ( .A(n14146), .ZN(n14147) );
  AOI21_X1 U15969 ( .B1(n14148), .B2(n14770), .A(n14147), .ZN(n14317) );
  INV_X1 U15970 ( .A(n14317), .ZN(n14149) );
  AOI21_X1 U15971 ( .B1(n14314), .B2(n14150), .A(n14149), .ZN(n14160) );
  OAI21_X1 U15972 ( .B1(n14153), .B2(n14152), .A(n14151), .ZN(n14318) );
  INV_X1 U15973 ( .A(n14318), .ZN(n14158) );
  AOI22_X1 U15974 ( .A1(n14724), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14154), 
        .B2(n14713), .ZN(n14155) );
  OAI21_X1 U15975 ( .B1(n14156), .B2(n14258), .A(n14155), .ZN(n14157) );
  AOI21_X1 U15976 ( .B1(n14158), .B2(n14703), .A(n14157), .ZN(n14159) );
  OAI21_X1 U15977 ( .B1(n14160), .B2(n14724), .A(n14159), .ZN(P1_U3267) );
  AOI21_X1 U15978 ( .B1(n14173), .B2(n14162), .A(n14161), .ZN(n14164) );
  OAI21_X1 U15979 ( .B1(n14164), .B2(n14710), .A(n14163), .ZN(n14165) );
  INV_X1 U15980 ( .A(n14165), .ZN(n14325) );
  NAND2_X1 U15981 ( .A1(n14320), .A2(n6507), .ZN(n14166) );
  NAND2_X1 U15982 ( .A1(n14166), .A2(n14749), .ZN(n14167) );
  NOR2_X1 U15983 ( .A1(n14168), .A2(n14167), .ZN(n14319) );
  NAND2_X1 U15984 ( .A1(n14320), .A2(n14715), .ZN(n14171) );
  AOI22_X1 U15985 ( .A1(n14724), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n14713), 
        .B2(n14169), .ZN(n14170) );
  NAND2_X1 U15986 ( .A1(n14171), .A2(n14170), .ZN(n14172) );
  AOI21_X1 U15987 ( .B1(n14319), .B2(n14720), .A(n14172), .ZN(n14176) );
  OR2_X1 U15988 ( .A1(n14174), .A2(n14173), .ZN(n14322) );
  NAND3_X1 U15989 ( .A1(n14322), .A2(n14321), .A3(n14703), .ZN(n14175) );
  OAI211_X1 U15990 ( .C1(n14325), .C2(n14724), .A(n14176), .B(n14175), .ZN(
        P1_U3268) );
  OAI211_X1 U15991 ( .C1(n14178), .C2(n14183), .A(n14177), .B(n14770), .ZN(
        n14180) );
  AOI21_X1 U15992 ( .B1(n14183), .B2(n14182), .A(n14181), .ZN(n14330) );
  INV_X1 U15993 ( .A(n14330), .ZN(n14190) );
  AOI21_X1 U15994 ( .B1(n14327), .B2(n6502), .A(n14294), .ZN(n14184) );
  AND2_X1 U15995 ( .A1(n14184), .A2(n6507), .ZN(n14326) );
  NAND2_X1 U15996 ( .A1(n14326), .A2(n14720), .ZN(n14187) );
  AOI22_X1 U15997 ( .A1(n14724), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14185), 
        .B2(n14713), .ZN(n14186) );
  OAI211_X1 U15998 ( .C1(n14188), .C2(n14258), .A(n14187), .B(n14186), .ZN(
        n14189) );
  AOI21_X1 U15999 ( .B1(n14190), .B2(n14703), .A(n14189), .ZN(n14191) );
  OAI21_X1 U16000 ( .B1(n14329), .B2(n14724), .A(n14191), .ZN(P1_U3269) );
  XNOR2_X1 U16001 ( .A(n14192), .B(n14199), .ZN(n14194) );
  AOI21_X1 U16002 ( .B1(n14194), .B2(n14770), .A(n14193), .ZN(n14334) );
  AOI21_X1 U16003 ( .B1(n14209), .B2(n14332), .A(n14294), .ZN(n14195) );
  AND2_X1 U16004 ( .A1(n14195), .A2(n6502), .ZN(n14331) );
  NAND2_X1 U16005 ( .A1(n14332), .A2(n14715), .ZN(n14197) );
  NAND2_X1 U16006 ( .A1(n14724), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n14196) );
  OAI211_X1 U16007 ( .C1(n14252), .C2(n14198), .A(n14197), .B(n14196), .ZN(
        n14202) );
  OAI21_X1 U16008 ( .B1(n7424), .B2(n14083), .A(n14200), .ZN(n14335) );
  NOR2_X1 U16009 ( .A1(n14335), .A2(n14262), .ZN(n14201) );
  AOI211_X1 U16010 ( .C1(n14331), .C2(n14720), .A(n14202), .B(n14201), .ZN(
        n14203) );
  OAI21_X1 U16011 ( .B1(n14334), .B2(n14724), .A(n14203), .ZN(P1_U3270) );
  XNOR2_X1 U16012 ( .A(n14204), .B(n14206), .ZN(n14342) );
  OAI21_X1 U16013 ( .B1(n14207), .B2(n14206), .A(n14205), .ZN(n14336) );
  NAND2_X1 U16014 ( .A1(n14336), .A2(n14284), .ZN(n14216) );
  INV_X1 U16015 ( .A(n14209), .ZN(n14210) );
  AOI211_X1 U16016 ( .C1(n14339), .C2(n14222), .A(n14294), .B(n14210), .ZN(
        n14337) );
  AOI22_X1 U16017 ( .A1(n14211), .A2(n14713), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n14724), .ZN(n14213) );
  NAND2_X1 U16018 ( .A1(n14338), .A2(n14282), .ZN(n14212) );
  OAI211_X1 U16019 ( .C1(n7153), .C2(n14258), .A(n14213), .B(n14212), .ZN(
        n14214) );
  AOI21_X1 U16020 ( .B1(n14337), .B2(n14720), .A(n14214), .ZN(n14215) );
  OAI211_X1 U16021 ( .C1(n14342), .C2(n14262), .A(n14216), .B(n14215), .ZN(
        P1_U3271) );
  INV_X1 U16022 ( .A(n14217), .ZN(n14218) );
  AOI21_X1 U16023 ( .B1(n7139), .B2(n14219), .A(n14218), .ZN(n14349) );
  AOI21_X1 U16024 ( .B1(n14221), .B2(n14220), .A(n6551), .ZN(n14343) );
  NAND2_X1 U16025 ( .A1(n14343), .A2(n14284), .ZN(n14231) );
  AOI211_X1 U16026 ( .C1(n14346), .C2(n14223), .A(n14294), .B(n14208), .ZN(
        n14344) );
  INV_X1 U16027 ( .A(n14224), .ZN(n14225) );
  AOI22_X1 U16028 ( .A1(n14225), .A2(n14713), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n14724), .ZN(n14227) );
  NAND2_X1 U16029 ( .A1(n14345), .A2(n14282), .ZN(n14226) );
  OAI211_X1 U16030 ( .C1(n14228), .C2(n14258), .A(n14227), .B(n14226), .ZN(
        n14229) );
  AOI21_X1 U16031 ( .B1(n14344), .B2(n14720), .A(n14229), .ZN(n14230) );
  OAI211_X1 U16032 ( .C1(n14349), .C2(n14262), .A(n14231), .B(n14230), .ZN(
        P1_U3272) );
  AOI211_X1 U16033 ( .C1(n14076), .C2(n14233), .A(n14710), .B(n14232), .ZN(
        n14235) );
  NOR2_X1 U16034 ( .A1(n14235), .A2(n14234), .ZN(n14356) );
  XNOR2_X1 U16035 ( .A(n14251), .B(n14351), .ZN(n14236) );
  AND2_X1 U16036 ( .A1(n14236), .A2(n14749), .ZN(n14350) );
  INV_X1 U16037 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14237) );
  OAI22_X1 U16038 ( .A1(n14238), .A2(n14252), .B1(n14282), .B2(n14237), .ZN(
        n14239) );
  INV_X1 U16039 ( .A(n14239), .ZN(n14240) );
  OAI21_X1 U16040 ( .B1(n14241), .B2(n14258), .A(n14240), .ZN(n14242) );
  AOI21_X1 U16041 ( .B1(n14350), .B2(n14720), .A(n14242), .ZN(n14246) );
  NAND2_X1 U16042 ( .A1(n14244), .A2(n14243), .ZN(n14352) );
  NAND3_X1 U16043 ( .A1(n14353), .A2(n14352), .A3(n14703), .ZN(n14245) );
  OAI211_X1 U16044 ( .C1(n14356), .C2(n14724), .A(n14246), .B(n14245), .ZN(
        P1_U3273) );
  XNOR2_X1 U16045 ( .A(n14249), .B(n14247), .ZN(n14362) );
  OAI21_X1 U16046 ( .B1(n14250), .B2(n14249), .A(n14248), .ZN(n14359) );
  AOI211_X1 U16047 ( .C1(n12379), .C2(n14264), .A(n14294), .B(n14251), .ZN(
        n14357) );
  NAND2_X1 U16048 ( .A1(n14357), .A2(n14720), .ZN(n14257) );
  INV_X1 U16049 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14254) );
  OAI22_X1 U16050 ( .A1(n14282), .A2(n14254), .B1(n14253), .B2(n14252), .ZN(
        n14255) );
  AOI21_X1 U16051 ( .B1(n14358), .B2(n14282), .A(n14255), .ZN(n14256) );
  OAI211_X1 U16052 ( .C1(n14259), .C2(n14258), .A(n14257), .B(n14256), .ZN(
        n14260) );
  AOI21_X1 U16053 ( .B1(n14284), .B2(n14359), .A(n14260), .ZN(n14261) );
  OAI21_X1 U16054 ( .B1(n14362), .B2(n14262), .A(n14261), .ZN(P1_U3274) );
  XNOR2_X1 U16055 ( .A(n14263), .B(n14272), .ZN(n14370) );
  OAI211_X1 U16056 ( .C1(n14366), .C2(n14265), .A(n14749), .B(n14264), .ZN(
        n14365) );
  AOI22_X1 U16057 ( .A1(n14724), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14266), 
        .B2(n14713), .ZN(n14269) );
  NAND2_X1 U16058 ( .A1(n14267), .A2(n14715), .ZN(n14268) );
  OAI211_X1 U16059 ( .C1(n14365), .C2(n14270), .A(n14269), .B(n14268), .ZN(
        n14277) );
  NOR2_X1 U16060 ( .A1(n14273), .A2(n14272), .ZN(n14274) );
  AOI21_X1 U16061 ( .B1(n14367), .B2(n14364), .A(n14724), .ZN(n14276) );
  AOI211_X1 U16062 ( .C1(n14703), .C2(n14370), .A(n14277), .B(n14276), .ZN(
        n14278) );
  INV_X1 U16063 ( .A(n14278), .ZN(P1_U3275) );
  OAI21_X1 U16064 ( .B1(n14280), .B2(n14715), .A(n14279), .ZN(n14288) );
  AOI22_X1 U16065 ( .A1(n14282), .A2(n14281), .B1(n14713), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n14287) );
  OAI21_X1 U16066 ( .B1(n14284), .B2(n14703), .A(n14283), .ZN(n14286) );
  NAND2_X1 U16067 ( .A1(n14724), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n14285) );
  NAND4_X1 U16068 ( .A1(n14288), .A2(n14287), .A3(n14286), .A4(n14285), .ZN(
        P1_U3293) );
  OAI211_X1 U16069 ( .C1(n14290), .C2(n14780), .A(n14289), .B(n14291), .ZN(
        n14372) );
  MUX2_X1 U16070 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14372), .S(n14798), .Z(
        P1_U3559) );
  MUX2_X1 U16071 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14373), .S(n14798), .Z(
        P1_U3558) );
  MUX2_X1 U16072 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14374), .S(n14798), .Z(
        P1_U3557) );
  OAI211_X1 U16073 ( .C1(n14303), .C2(n14780), .A(n14302), .B(n14301), .ZN(
        n14304) );
  NAND2_X1 U16074 ( .A1(n14307), .A2(n7429), .ZN(n14375) );
  MUX2_X1 U16075 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14375), .S(n14798), .Z(
        P1_U3556) );
  INV_X1 U16076 ( .A(n14308), .ZN(n14309) );
  AOI21_X1 U16077 ( .B1(n14310), .B2(n14735), .A(n14309), .ZN(n14311) );
  OAI211_X1 U16078 ( .C1(n14363), .C2(n14313), .A(n14312), .B(n14311), .ZN(
        n14376) );
  MUX2_X1 U16079 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14376), .S(n14798), .Z(
        P1_U3555) );
  AOI21_X1 U16080 ( .B1(n14315), .B2(n14735), .A(n14314), .ZN(n14316) );
  OAI211_X1 U16081 ( .C1(n14363), .C2(n14318), .A(n14317), .B(n14316), .ZN(
        n14377) );
  MUX2_X1 U16082 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14377), .S(n14798), .Z(
        P1_U3554) );
  AOI21_X1 U16083 ( .B1(n14320), .B2(n14735), .A(n14319), .ZN(n14324) );
  NAND3_X1 U16084 ( .A1(n14322), .A2(n14784), .A3(n14321), .ZN(n14323) );
  NAND3_X1 U16085 ( .A1(n14325), .A2(n14324), .A3(n14323), .ZN(n14378) );
  MUX2_X1 U16086 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14378), .S(n14798), .Z(
        P1_U3553) );
  AOI21_X1 U16087 ( .B1(n14327), .B2(n14735), .A(n14326), .ZN(n14328) );
  OAI211_X1 U16088 ( .C1(n14363), .C2(n14330), .A(n14329), .B(n14328), .ZN(
        n14379) );
  MUX2_X1 U16089 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14379), .S(n14798), .Z(
        P1_U3552) );
  AOI21_X1 U16090 ( .B1(n14332), .B2(n14735), .A(n14331), .ZN(n14333) );
  OAI211_X1 U16091 ( .C1(n14363), .C2(n14335), .A(n14334), .B(n14333), .ZN(
        n14380) );
  MUX2_X1 U16092 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14380), .S(n14798), .Z(
        P1_U3551) );
  NAND2_X1 U16093 ( .A1(n14336), .A2(n14770), .ZN(n14341) );
  AOI211_X1 U16094 ( .C1(n14339), .C2(n14735), .A(n14338), .B(n14337), .ZN(
        n14340) );
  OAI211_X1 U16095 ( .C1(n14363), .C2(n14342), .A(n14341), .B(n14340), .ZN(
        n14381) );
  MUX2_X1 U16096 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14381), .S(n14798), .Z(
        P1_U3550) );
  NAND2_X1 U16097 ( .A1(n14343), .A2(n14770), .ZN(n14348) );
  AOI211_X1 U16098 ( .C1(n14346), .C2(n14735), .A(n14345), .B(n14344), .ZN(
        n14347) );
  OAI211_X1 U16099 ( .C1(n14363), .C2(n14349), .A(n14348), .B(n14347), .ZN(
        n14382) );
  MUX2_X1 U16100 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14382), .S(n14798), .Z(
        P1_U3549) );
  AOI21_X1 U16101 ( .B1(n14351), .B2(n14735), .A(n14350), .ZN(n14355) );
  NAND3_X1 U16102 ( .A1(n14353), .A2(n14352), .A3(n14784), .ZN(n14354) );
  NAND3_X1 U16103 ( .A1(n14356), .A2(n14355), .A3(n14354), .ZN(n14383) );
  MUX2_X1 U16104 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14383), .S(n14798), .Z(
        P1_U3548) );
  AOI211_X1 U16105 ( .C1(n12379), .C2(n14735), .A(n14358), .B(n14357), .ZN(
        n14361) );
  NAND2_X1 U16106 ( .A1(n14359), .A2(n14770), .ZN(n14360) );
  OAI211_X1 U16107 ( .C1(n14363), .C2(n14362), .A(n14361), .B(n14360), .ZN(
        n14384) );
  MUX2_X1 U16108 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14384), .S(n14798), .Z(
        P1_U3547) );
  OAI211_X1 U16109 ( .C1(n14366), .C2(n14780), .A(n14365), .B(n14364), .ZN(
        n14369) );
  INV_X1 U16110 ( .A(n14367), .ZN(n14368) );
  AOI211_X1 U16111 ( .C1(n14784), .C2(n14370), .A(n14369), .B(n14368), .ZN(
        n14371) );
  INV_X1 U16112 ( .A(n14371), .ZN(n14385) );
  MUX2_X1 U16113 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14385), .S(n14798), .Z(
        P1_U3546) );
  MUX2_X1 U16114 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14372), .S(n14748), .Z(
        P1_U3527) );
  MUX2_X1 U16115 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14373), .S(n14748), .Z(
        P1_U3526) );
  MUX2_X1 U16116 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14374), .S(n14748), .Z(
        P1_U3525) );
  MUX2_X1 U16117 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14375), .S(n14748), .Z(
        P1_U3524) );
  MUX2_X1 U16118 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14376), .S(n14748), .Z(
        P1_U3523) );
  MUX2_X1 U16119 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14377), .S(n14748), .Z(
        P1_U3522) );
  MUX2_X1 U16120 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14378), .S(n14748), .Z(
        P1_U3521) );
  MUX2_X1 U16121 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14379), .S(n14748), .Z(
        P1_U3520) );
  MUX2_X1 U16122 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14380), .S(n14748), .Z(
        P1_U3519) );
  MUX2_X1 U16123 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14381), .S(n14748), .Z(
        P1_U3518) );
  MUX2_X1 U16124 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14382), .S(n14748), .Z(
        P1_U3517) );
  MUX2_X1 U16125 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14383), .S(n14748), .Z(
        P1_U3516) );
  MUX2_X1 U16126 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14384), .S(n14748), .Z(
        P1_U3515) );
  MUX2_X1 U16127 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14385), .S(n14748), .Z(
        P1_U3513) );
  NOR4_X1 U16128 ( .A1(n14387), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n14386), .ZN(n14388) );
  AOI21_X1 U16129 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n14389), .A(n14388), 
        .ZN(n14390) );
  OAI21_X1 U16130 ( .B1(n14392), .B2(n14391), .A(n14390), .ZN(P1_U3324) );
  OAI222_X1 U16131 ( .A1(n14391), .A2(n14395), .B1(n14394), .B2(P1_U3086), 
        .C1(n14393), .C2(n14396), .ZN(P1_U3326) );
  OAI222_X1 U16132 ( .A1(n14398), .A2(P1_U3086), .B1(n14391), .B2(n14397), 
        .C1(n15230), .C2(n14396), .ZN(P1_U3328) );
  MUX2_X1 U16133 ( .A(n12254), .B(n14399), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16134 ( .A(n14400), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16135 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14441) );
  INV_X1 U16136 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14692) );
  INV_X1 U16137 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14433) );
  XOR2_X1 U16138 ( .A(n14433), .B(P1_ADDR_REG_14__SCAN_IN), .Z(n14511) );
  INV_X1 U16139 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14992) );
  INV_X1 U16140 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14430) );
  INV_X1 U16141 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14450) );
  NOR2_X1 U16142 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n14450), .ZN(n14428) );
  INV_X1 U16143 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14424) );
  XOR2_X1 U16144 ( .A(n14424), .B(P3_ADDR_REG_9__SCAN_IN), .Z(n14490) );
  NOR2_X2 U16145 ( .A1(n14461), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n14460) );
  INV_X1 U16146 ( .A(n14460), .ZN(n14401) );
  XNOR2_X1 U16147 ( .A(n14403), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n14457) );
  INV_X1 U16148 ( .A(n14457), .ZN(n14405) );
  NOR2_X1 U16149 ( .A1(n14408), .A2(n14407), .ZN(n14410) );
  NOR2_X1 U16150 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n14467), .ZN(n14409) );
  NOR2_X1 U16151 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n14455), .ZN(n14413) );
  NOR2_X1 U16152 ( .A1(n14411), .A2(n6865), .ZN(n14412) );
  INV_X1 U16153 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14414) );
  NOR2_X1 U16154 ( .A1(n14415), .A2(n14414), .ZN(n14417) );
  AND2_X1 U16155 ( .A1(n14476), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n14418) );
  NOR2_X1 U16156 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14419), .ZN(n14421) );
  XNOR2_X1 U16157 ( .A(n14419), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14481) );
  INV_X1 U16158 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14482) );
  XOR2_X1 U16159 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Z(
        n14453) );
  NAND2_X1 U16160 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14425), .ZN(n14497) );
  NAND2_X1 U16161 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n14497), .ZN(n14426) );
  INV_X1 U16162 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14427) );
  XNOR2_X1 U16163 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n14430), .ZN(n14448) );
  AND2_X1 U16164 ( .A1(n14992), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14431) );
  NAND2_X1 U16165 ( .A1(n14511), .A2(n14510), .ZN(n14432) );
  INV_X1 U16166 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14549) );
  NAND2_X1 U16167 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14549), .ZN(n14434) );
  AOI22_X1 U16168 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14692), .B1(n14444), 
        .B2(n14434), .ZN(n14443) );
  OR2_X1 U16169 ( .A1(n14441), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n14435) );
  AOI22_X1 U16170 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14441), .B1(n14443), 
        .B2(n14435), .ZN(n14436) );
  INV_X1 U16171 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14437) );
  NAND2_X1 U16172 ( .A1(n14436), .A2(n14437), .ZN(n14439) );
  XOR2_X1 U16173 ( .A(n14437), .B(n14436), .Z(n14514) );
  NAND2_X1 U16174 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14514), .ZN(n14438) );
  NAND2_X1 U16175 ( .A1(n14439), .A2(n14438), .ZN(n14537) );
  NOR2_X1 U16176 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14540), .ZN(n14440) );
  AOI21_X1 U16177 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14540), .A(n14440), 
        .ZN(n14538) );
  XNOR2_X1 U16178 ( .A(n14537), .B(n14538), .ZN(n14533) );
  INV_X1 U16179 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14915) );
  XNOR2_X1 U16180 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(n14441), .ZN(n14442) );
  XNOR2_X1 U16181 ( .A(n14443), .B(n14442), .ZN(n14673) );
  XOR2_X1 U16182 ( .A(n14692), .B(P3_ADDR_REG_15__SCAN_IN), .Z(n14445) );
  XNOR2_X1 U16183 ( .A(n14445), .B(n14444), .ZN(n14668) );
  INV_X1 U16184 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14887) );
  XNOR2_X1 U16185 ( .A(n14992), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n14446) );
  XNOR2_X1 U16186 ( .A(n14447), .B(n14446), .ZN(n14659) );
  XNOR2_X1 U16187 ( .A(n14449), .B(n14448), .ZN(n14504) );
  XOR2_X1 U16188 ( .A(n14450), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n14452) );
  XNOR2_X1 U16189 ( .A(n14452), .B(n14451), .ZN(n14503) );
  INV_X1 U16190 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14501) );
  XOR2_X1 U16191 ( .A(n14454), .B(n14453), .Z(n14486) );
  NAND2_X1 U16192 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14456), .ZN(n14470) );
  INV_X1 U16193 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14848) );
  XNOR2_X1 U16194 ( .A(n14458), .B(n14457), .ZN(n14466) );
  XOR2_X1 U16195 ( .A(n14460), .B(n14459), .Z(n14462) );
  NAND2_X1 U16196 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14462), .ZN(n14464) );
  AOI21_X1 U16197 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14461), .A(n14460), .ZN(
        n15301) );
  INV_X1 U16198 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15300) );
  NOR2_X1 U16199 ( .A1(n15301), .A2(n15300), .ZN(n15310) );
  NAND2_X1 U16200 ( .A1(n14464), .A2(n14463), .ZN(n14465) );
  NAND2_X1 U16201 ( .A1(n14466), .A2(n14465), .ZN(n14518) );
  NOR2_X1 U16202 ( .A1(n14466), .A2(n14465), .ZN(n14519) );
  INV_X1 U16203 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n15145) );
  XOR2_X1 U16204 ( .A(n15145), .B(n14467), .Z(n15306) );
  NOR2_X1 U16205 ( .A1(n15305), .A2(n15306), .ZN(n14468) );
  INV_X1 U16206 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15307) );
  NAND2_X1 U16207 ( .A1(n15305), .A2(n15306), .ZN(n15304) );
  OAI21_X1 U16208 ( .B1(n14468), .B2(n15307), .A(n15304), .ZN(n15297) );
  NAND2_X1 U16209 ( .A1(n15298), .A2(n15297), .ZN(n14469) );
  NAND2_X1 U16210 ( .A1(n14475), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14480) );
  INV_X1 U16211 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14474) );
  XOR2_X1 U16212 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n14476), .Z(n14478) );
  XOR2_X1 U16213 ( .A(n14478), .B(n14477), .Z(n14521) );
  NAND2_X1 U16214 ( .A1(n14522), .A2(n14521), .ZN(n14479) );
  XOR2_X1 U16215 ( .A(n14482), .B(n14481), .Z(n15303) );
  NAND2_X1 U16216 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14483), .ZN(n14484) );
  XNOR2_X1 U16217 ( .A(n14486), .B(n14485), .ZN(n14523) );
  NOR2_X1 U16218 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n14523), .ZN(n14488) );
  NOR2_X1 U16219 ( .A1(n14486), .A2(n14485), .ZN(n14487) );
  NOR2_X2 U16220 ( .A1(n14488), .A2(n14487), .ZN(n14493) );
  XNOR2_X1 U16221 ( .A(n14490), .B(n14489), .ZN(n14491) );
  NAND2_X1 U16222 ( .A1(n14493), .A2(n14491), .ZN(n14495) );
  NAND2_X1 U16223 ( .A1(n14524), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n14494) );
  NAND2_X1 U16224 ( .A1(n14495), .A2(n14494), .ZN(n14526) );
  INV_X1 U16225 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14499) );
  NAND2_X1 U16226 ( .A1(n14497), .A2(n14496), .ZN(n14498) );
  XNOR2_X1 U16227 ( .A(n14499), .B(n14498), .ZN(n14527) );
  NAND2_X1 U16228 ( .A1(n14526), .A2(n14527), .ZN(n14500) );
  NOR2_X1 U16229 ( .A1(n14526), .A2(n14527), .ZN(n14525) );
  AOI21_X2 U16230 ( .B1(n14501), .B2(n14500), .A(n14525), .ZN(n14502) );
  NAND2_X1 U16231 ( .A1(n14503), .A2(n14502), .ZN(n15294) );
  INV_X1 U16232 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n15291) );
  NOR2_X1 U16233 ( .A1(n14503), .A2(n14502), .ZN(n15292) );
  AOI21_X2 U16234 ( .B1(n15294), .B2(n15291), .A(n15292), .ZN(n14505) );
  INV_X1 U16235 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14506) );
  NAND2_X1 U16236 ( .A1(n14507), .A2(n14506), .ZN(n14508) );
  XNOR2_X1 U16237 ( .A(n14511), .B(n14510), .ZN(n14663) );
  INV_X1 U16238 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14669) );
  NAND2_X1 U16239 ( .A1(n14668), .A2(n14667), .ZN(n14666) );
  OAI21_X2 U16240 ( .B1(n14512), .B2(n14669), .A(n14666), .ZN(n14672) );
  NAND2_X1 U16241 ( .A1(n14673), .A2(n14672), .ZN(n14513) );
  INV_X1 U16242 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14900) );
  XNOR2_X1 U16243 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14514), .ZN(n14529) );
  XNOR2_X1 U16244 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14532), .ZN(SUB_1596_U62)
         );
  INV_X1 U16245 ( .A(P2_WR_REG_SCAN_IN), .ZN(n14516) );
  INV_X1 U16246 ( .A(P1_WR_REG_SCAN_IN), .ZN(n14515) );
  INV_X1 U16247 ( .A(P3_WR_REG_SCAN_IN), .ZN(n15231) );
  OAI221_X1 U16248 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .C1(
        n14516), .C2(n14515), .A(n15231), .ZN(U28) );
  AOI21_X1 U16249 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14517) );
  OAI21_X1 U16250 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14517), 
        .ZN(U29) );
  INV_X1 U16251 ( .A(n14518), .ZN(n14520) );
  AOI222_X1 U16252 ( .A1(n14848), .A2(n14520), .B1(n14848), .B2(n14519), .C1(
        n15305), .C2(n14518), .ZN(SUB_1596_U61) );
  XOR2_X1 U16253 ( .A(n14522), .B(n14521), .Z(SUB_1596_U57) );
  XNOR2_X1 U16254 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14523), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16255 ( .A(n14524), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  AOI21_X1 U16256 ( .B1(n14527), .B2(n14526), .A(n14525), .ZN(n14528) );
  XOR2_X1 U16257 ( .A(n14528), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  AOI21_X1 U16258 ( .B1(n14530), .B2(n14529), .A(n6577), .ZN(n14531) );
  XOR2_X1 U16259 ( .A(n14531), .B(P2_ADDR_REG_17__SCAN_IN), .Z(SUB_1596_U63)
         );
  NOR2_X1 U16260 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n14532), .ZN(n14536) );
  NOR2_X1 U16261 ( .A1(n14534), .A2(n14533), .ZN(n14535) );
  NOR2_X1 U16262 ( .A1(n14536), .A2(n14535), .ZN(n14545) );
  NAND2_X1 U16263 ( .A1(n14538), .A2(n14537), .ZN(n14539) );
  OAI21_X1 U16264 ( .B1(n14540), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14539), 
        .ZN(n14543) );
  XNOR2_X1 U16265 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14541) );
  XNOR2_X1 U16266 ( .A(n14541), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n14542) );
  XNOR2_X1 U16267 ( .A(n14543), .B(n14542), .ZN(n14544) );
  XNOR2_X1 U16268 ( .A(n14545), .B(n14544), .ZN(SUB_1596_U4) );
  AOI21_X1 U16269 ( .B1(n14548), .B2(n14547), .A(n14546), .ZN(n14562) );
  OAI22_X1 U16270 ( .A1(n14994), .A2(n6687), .B1(n14549), .B2(n14991), .ZN(
        n14559) );
  AOI21_X1 U16271 ( .B1(n14552), .B2(n14551), .A(n14550), .ZN(n14557) );
  AOI21_X1 U16272 ( .B1(n14555), .B2(n14554), .A(n14553), .ZN(n14556) );
  OAI22_X1 U16273 ( .A1(n14557), .A2(n15002), .B1(n14556), .B2(n15000), .ZN(
        n14558) );
  NOR3_X1 U16274 ( .A1(n14560), .A2(n14559), .A3(n14558), .ZN(n14561) );
  OAI21_X1 U16275 ( .B1(n14562), .B2(n15008), .A(n14561), .ZN(P3_U3197) );
  AOI21_X1 U16276 ( .B1(n8130), .B2(n15065), .A(n14565), .ZN(n14584) );
  INV_X1 U16277 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14564) );
  AOI22_X1 U16278 ( .A1(n15106), .A2(n14584), .B1(n14564), .B2(n15104), .ZN(
        P3_U3490) );
  AOI21_X1 U16279 ( .B1(n14566), .B2(n15065), .A(n14565), .ZN(n14586) );
  INV_X1 U16280 ( .A(n14586), .ZN(n14567) );
  OAI22_X1 U16281 ( .A1(n15104), .A2(n14567), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n15106), .ZN(n14568) );
  INV_X1 U16282 ( .A(n14568), .ZN(P3_U3489) );
  NOR2_X1 U16283 ( .A1(n14569), .A2(n15079), .ZN(n14571) );
  AOI211_X1 U16284 ( .C1(n14572), .C2(n14581), .A(n14571), .B(n14570), .ZN(
        n14588) );
  AOI22_X1 U16285 ( .A1(n15106), .A2(n14588), .B1(n15259), .B2(n15104), .ZN(
        P3_U3472) );
  NOR2_X1 U16286 ( .A1(n14573), .A2(n15079), .ZN(n14575) );
  AOI211_X1 U16287 ( .C1(n14581), .C2(n14576), .A(n14575), .B(n14574), .ZN(
        n14589) );
  AOI22_X1 U16288 ( .A1(n15106), .A2(n14589), .B1(n11554), .B2(n15104), .ZN(
        P3_U3471) );
  NOR2_X1 U16289 ( .A1(n14577), .A2(n15079), .ZN(n14579) );
  AOI211_X1 U16290 ( .C1(n14581), .C2(n14580), .A(n14579), .B(n14578), .ZN(
        n14591) );
  AOI22_X1 U16291 ( .A1(n15106), .A2(n14591), .B1(n14582), .B2(n15104), .ZN(
        P3_U3470) );
  INV_X1 U16292 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14583) );
  AOI22_X1 U16293 ( .A1(n15089), .A2(n14584), .B1(n14583), .B2(n15087), .ZN(
        P3_U3458) );
  AOI22_X1 U16294 ( .A1(n15089), .A2(n14586), .B1(n14585), .B2(n15087), .ZN(
        P3_U3457) );
  INV_X1 U16295 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14587) );
  AOI22_X1 U16296 ( .A1(n15089), .A2(n14588), .B1(n14587), .B2(n15087), .ZN(
        P3_U3429) );
  INV_X1 U16297 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n15128) );
  AOI22_X1 U16298 ( .A1(n15089), .A2(n14589), .B1(n15128), .B2(n15087), .ZN(
        P3_U3426) );
  INV_X1 U16299 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14590) );
  AOI22_X1 U16300 ( .A1(n15089), .A2(n14591), .B1(n14590), .B2(n15087), .ZN(
        P3_U3423) );
  OAI211_X1 U16301 ( .C1(n14594), .C2(n14967), .A(n14593), .B(n14592), .ZN(
        n14595) );
  AOI21_X1 U16302 ( .B1(n14951), .B2(n14596), .A(n14595), .ZN(n14598) );
  AOI22_X1 U16303 ( .A1(n14986), .A2(n14598), .B1(n14597), .B2(n14984), .ZN(
        P2_U3511) );
  AOI22_X1 U16304 ( .A1(n14974), .A2(n14598), .B1(n8759), .B2(n14973), .ZN(
        P2_U3466) );
  XNOR2_X1 U16305 ( .A(n14599), .B(n14613), .ZN(n14628) );
  INV_X1 U16306 ( .A(n14600), .ZN(n14603) );
  INV_X1 U16307 ( .A(n14601), .ZN(n14602) );
  OAI211_X1 U16308 ( .C1(n14625), .C2(n14603), .A(n14602), .B(n14749), .ZN(
        n14624) );
  INV_X1 U16309 ( .A(n14604), .ZN(n14605) );
  AOI22_X1 U16310 ( .A1(n14607), .A2(n14606), .B1(n14605), .B2(n14713), .ZN(
        n14608) );
  OAI21_X1 U16311 ( .B1(n14624), .B2(n14609), .A(n14608), .ZN(n14616) );
  INV_X1 U16312 ( .A(n14610), .ZN(n14611) );
  AOI21_X1 U16313 ( .B1(n14613), .B2(n14612), .A(n14611), .ZN(n14615) );
  OAI21_X1 U16314 ( .B1(n14615), .B2(n14710), .A(n14614), .ZN(n14626) );
  AOI211_X1 U16315 ( .C1(n14703), .C2(n14628), .A(n14616), .B(n14626), .ZN(
        n14617) );
  AOI22_X1 U16316 ( .A1(n14724), .A2(n11750), .B1(n14617), .B2(n14282), .ZN(
        P1_U3277) );
  OAI21_X1 U16317 ( .B1(n14619), .B2(n14780), .A(n14618), .ZN(n14621) );
  AOI211_X1 U16318 ( .C1(n14622), .C2(n14784), .A(n14621), .B(n14620), .ZN(
        n14648) );
  AOI22_X1 U16319 ( .A1(n14798), .A2(n14648), .B1(n14623), .B2(n14796), .ZN(
        P1_U3545) );
  OAI21_X1 U16320 ( .B1(n14625), .B2(n14780), .A(n14624), .ZN(n14627) );
  AOI211_X1 U16321 ( .C1(n14628), .C2(n14784), .A(n14627), .B(n14626), .ZN(
        n14650) );
  AOI22_X1 U16322 ( .A1(n14798), .A2(n14650), .B1(n11740), .B2(n14796), .ZN(
        P1_U3544) );
  OAI211_X1 U16323 ( .C1(n14631), .C2(n14780), .A(n14630), .B(n14629), .ZN(
        n14632) );
  AOI21_X1 U16324 ( .B1(n14784), .B2(n14633), .A(n14632), .ZN(n14652) );
  AOI22_X1 U16325 ( .A1(n14798), .A2(n14652), .B1(n14678), .B2(n14796), .ZN(
        P1_U3543) );
  OAI211_X1 U16326 ( .C1(n14636), .C2(n14780), .A(n14635), .B(n14634), .ZN(
        n14640) );
  AND3_X1 U16327 ( .A1(n14638), .A2(n14784), .A3(n14637), .ZN(n14639) );
  AOI211_X1 U16328 ( .C1(n14770), .C2(n14641), .A(n14640), .B(n14639), .ZN(
        n14654) );
  AOI22_X1 U16329 ( .A1(n14798), .A2(n14654), .B1(n11114), .B2(n14796), .ZN(
        P1_U3542) );
  OAI21_X1 U16330 ( .B1(n14643), .B2(n14780), .A(n14642), .ZN(n14645) );
  AOI211_X1 U16331 ( .C1(n14646), .C2(n14784), .A(n14645), .B(n14644), .ZN(
        n14656) );
  AOI22_X1 U16332 ( .A1(n14798), .A2(n14656), .B1(n10332), .B2(n14796), .ZN(
        P1_U3539) );
  INV_X1 U16333 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14647) );
  AOI22_X1 U16334 ( .A1(n14748), .A2(n14648), .B1(n14647), .B2(n14785), .ZN(
        P1_U3510) );
  INV_X1 U16335 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14649) );
  AOI22_X1 U16336 ( .A1(n14748), .A2(n14650), .B1(n14649), .B2(n14785), .ZN(
        P1_U3507) );
  INV_X1 U16337 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14651) );
  AOI22_X1 U16338 ( .A1(n14748), .A2(n14652), .B1(n14651), .B2(n14785), .ZN(
        P1_U3504) );
  INV_X1 U16339 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14653) );
  AOI22_X1 U16340 ( .A1(n14748), .A2(n14654), .B1(n14653), .B2(n14785), .ZN(
        P1_U3501) );
  INV_X1 U16341 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14655) );
  AOI22_X1 U16342 ( .A1(n14748), .A2(n14656), .B1(n14655), .B2(n14785), .ZN(
        P1_U3492) );
  INV_X1 U16343 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14874) );
  XOR2_X1 U16344 ( .A(n14874), .B(n14657), .Z(SUB_1596_U68) );
  AOI21_X1 U16345 ( .B1(n14660), .B2(n14659), .A(n14658), .ZN(n14661) );
  XOR2_X1 U16346 ( .A(n14661), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16347 ( .B1(n14664), .B2(n14663), .A(n14662), .ZN(n14665) );
  XOR2_X1 U16348 ( .A(n14665), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  OAI21_X1 U16349 ( .B1(n14668), .B2(n14667), .A(n14666), .ZN(n14670) );
  XOR2_X1 U16350 ( .A(n14670), .B(n14669), .Z(SUB_1596_U65) );
  AOI21_X1 U16351 ( .B1(n14673), .B2(n14672), .A(n14671), .ZN(n14674) );
  XOR2_X1 U16352 ( .A(n14674), .B(P2_ADDR_REG_16__SCAN_IN), .Z(SUB_1596_U64)
         );
  AOI21_X1 U16353 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14676), .A(n14675), 
        .ZN(n14687) );
  OAI21_X1 U16354 ( .B1(n14679), .B2(n14678), .A(n14677), .ZN(n14681) );
  NAND2_X1 U16355 ( .A1(n14681), .A2(n14680), .ZN(n14685) );
  NAND2_X1 U16356 ( .A1(n14683), .A2(n14682), .ZN(n14684) );
  OAI211_X1 U16357 ( .C1(n14687), .C2(n14686), .A(n14685), .B(n14684), .ZN(
        n14688) );
  INV_X1 U16358 ( .A(n14688), .ZN(n14690) );
  OAI211_X1 U16359 ( .C1(n14692), .C2(n14691), .A(n14690), .B(n14689), .ZN(
        P1_U3258) );
  XNOR2_X1 U16360 ( .A(n14693), .B(n14699), .ZN(n14695) );
  AOI21_X1 U16361 ( .B1(n14695), .B2(n14770), .A(n14694), .ZN(n14761) );
  AOI222_X1 U16362 ( .A1(n14697), .A2(n14715), .B1(n14696), .B2(n14713), .C1(
        P1_REG2_REG_8__SCAN_IN), .C2(n14724), .ZN(n14705) );
  XNOR2_X1 U16363 ( .A(n14698), .B(n14699), .ZN(n14764) );
  OAI211_X1 U16364 ( .C1(n14701), .C2(n14760), .A(n14749), .B(n14700), .ZN(
        n14759) );
  INV_X1 U16365 ( .A(n14759), .ZN(n14702) );
  AOI22_X1 U16366 ( .A1(n14764), .A2(n14703), .B1(n14720), .B2(n14702), .ZN(
        n14704) );
  OAI211_X1 U16367 ( .C1(n14724), .C2(n14761), .A(n14705), .B(n14704), .ZN(
        P1_U3285) );
  XNOR2_X1 U16368 ( .A(n14706), .B(n14707), .ZN(n14746) );
  XNOR2_X1 U16369 ( .A(n14708), .B(n14707), .ZN(n14711) );
  OAI21_X1 U16370 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(n14712) );
  AOI21_X1 U16371 ( .B1(n14746), .B2(n14777), .A(n14712), .ZN(n14743) );
  AOI222_X1 U16372 ( .A1(n14716), .A2(n14715), .B1(n14714), .B2(n14713), .C1(
        P1_REG2_REG_6__SCAN_IN), .C2(n14724), .ZN(n14723) );
  OAI211_X1 U16373 ( .C1(n14718), .C2(n6867), .A(n14749), .B(n14717), .ZN(
        n14742) );
  INV_X1 U16374 ( .A(n14742), .ZN(n14719) );
  AOI22_X1 U16375 ( .A1(n14746), .A2(n14721), .B1(n14720), .B2(n14719), .ZN(
        n14722) );
  OAI211_X1 U16376 ( .C1(n14724), .C2(n14743), .A(n14723), .B(n14722), .ZN(
        P1_U3287) );
  INV_X1 U16377 ( .A(n14726), .ZN(n14725) );
  INV_X1 U16378 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n15263) );
  NOR2_X1 U16379 ( .A1(n14725), .A2(n15263), .ZN(P1_U3294) );
  AND2_X1 U16380 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14726), .ZN(P1_U3295) );
  AND2_X1 U16381 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14726), .ZN(P1_U3296) );
  AND2_X1 U16382 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14726), .ZN(P1_U3297) );
  AND2_X1 U16383 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14726), .ZN(P1_U3298) );
  AND2_X1 U16384 ( .A1(n14726), .A2(P1_D_REG_26__SCAN_IN), .ZN(P1_U3299) );
  AND2_X1 U16385 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14726), .ZN(P1_U3300) );
  AND2_X1 U16386 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14726), .ZN(P1_U3301) );
  AND2_X1 U16387 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14726), .ZN(P1_U3302) );
  AND2_X1 U16388 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14726), .ZN(P1_U3303) );
  AND2_X1 U16389 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14726), .ZN(P1_U3304) );
  AND2_X1 U16390 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14726), .ZN(P1_U3305) );
  AND2_X1 U16391 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14726), .ZN(P1_U3306) );
  AND2_X1 U16392 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14726), .ZN(P1_U3307) );
  AND2_X1 U16393 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14726), .ZN(P1_U3308) );
  AND2_X1 U16394 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14726), .ZN(P1_U3309) );
  AND2_X1 U16395 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14726), .ZN(P1_U3310) );
  AND2_X1 U16396 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14726), .ZN(P1_U3311) );
  AND2_X1 U16397 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14726), .ZN(P1_U3312) );
  AND2_X1 U16398 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14726), .ZN(P1_U3313) );
  AND2_X1 U16399 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14726), .ZN(P1_U3314) );
  AND2_X1 U16400 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14726), .ZN(P1_U3315) );
  INV_X1 U16401 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n15237) );
  NOR2_X1 U16402 ( .A1(n14725), .A2(n15237), .ZN(P1_U3316) );
  AND2_X1 U16403 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14726), .ZN(P1_U3317) );
  AND2_X1 U16404 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14726), .ZN(P1_U3318) );
  AND2_X1 U16405 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14726), .ZN(P1_U3319) );
  AND2_X1 U16406 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14726), .ZN(P1_U3320) );
  INV_X1 U16407 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n15132) );
  NOR2_X1 U16408 ( .A1(n14725), .A2(n15132), .ZN(P1_U3321) );
  AND2_X1 U16409 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14726), .ZN(P1_U3322) );
  AND2_X1 U16410 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14726), .ZN(P1_U3323) );
  INV_X1 U16411 ( .A(n14727), .ZN(n14728) );
  OAI21_X1 U16412 ( .B1(n14729), .B2(n14780), .A(n14728), .ZN(n14731) );
  AOI211_X1 U16413 ( .C1(n14754), .C2(n14732), .A(n14731), .B(n14730), .ZN(
        n14788) );
  INV_X1 U16414 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n15274) );
  AOI22_X1 U16415 ( .A1(n14748), .A2(n14788), .B1(n15274), .B2(n14785), .ZN(
        P1_U3462) );
  INV_X1 U16416 ( .A(n14738), .ZN(n14740) );
  AOI211_X1 U16417 ( .C1(n14736), .C2(n14735), .A(n14734), .B(n14733), .ZN(
        n14737) );
  OAI21_X1 U16418 ( .B1(n14773), .B2(n14738), .A(n14737), .ZN(n14739) );
  AOI21_X1 U16419 ( .B1(n14777), .B2(n14740), .A(n14739), .ZN(n14790) );
  INV_X1 U16420 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14741) );
  AOI22_X1 U16421 ( .A1(n14748), .A2(n14790), .B1(n14741), .B2(n14785), .ZN(
        P1_U3474) );
  OAI21_X1 U16422 ( .B1(n6867), .B2(n14780), .A(n14742), .ZN(n14745) );
  INV_X1 U16423 ( .A(n14743), .ZN(n14744) );
  AOI211_X1 U16424 ( .C1(n14754), .C2(n14746), .A(n14745), .B(n14744), .ZN(
        n14792) );
  INV_X1 U16425 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14747) );
  AOI22_X1 U16426 ( .A1(n14748), .A2(n14792), .B1(n14747), .B2(n14785), .ZN(
        P1_U3477) );
  NAND2_X1 U16427 ( .A1(n14750), .A2(n14749), .ZN(n14751) );
  OAI21_X1 U16428 ( .B1(n14752), .B2(n14780), .A(n14751), .ZN(n14753) );
  AOI21_X1 U16429 ( .B1(n14755), .B2(n14754), .A(n14753), .ZN(n14756) );
  AND2_X1 U16430 ( .A1(n14757), .A2(n14756), .ZN(n14793) );
  INV_X1 U16431 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14758) );
  AOI22_X1 U16432 ( .A1(n14748), .A2(n14793), .B1(n14758), .B2(n14785), .ZN(
        P1_U3480) );
  OAI21_X1 U16433 ( .B1(n14760), .B2(n14780), .A(n14759), .ZN(n14763) );
  INV_X1 U16434 ( .A(n14761), .ZN(n14762) );
  AOI211_X1 U16435 ( .C1(n14764), .C2(n14784), .A(n14763), .B(n14762), .ZN(
        n14794) );
  INV_X1 U16436 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14765) );
  AOI22_X1 U16437 ( .A1(n14748), .A2(n14794), .B1(n14765), .B2(n14785), .ZN(
        P1_U3483) );
  INV_X1 U16438 ( .A(n14774), .ZN(n14776) );
  OAI211_X1 U16439 ( .C1(n14768), .C2(n14780), .A(n14767), .B(n14766), .ZN(
        n14769) );
  AOI21_X1 U16440 ( .B1(n14771), .B2(n14770), .A(n14769), .ZN(n14772) );
  OAI21_X1 U16441 ( .B1(n14774), .B2(n14773), .A(n14772), .ZN(n14775) );
  AOI21_X1 U16442 ( .B1(n14777), .B2(n14776), .A(n14775), .ZN(n14795) );
  INV_X1 U16443 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15271) );
  AOI22_X1 U16444 ( .A1(n14748), .A2(n14795), .B1(n15271), .B2(n14785), .ZN(
        P1_U3486) );
  OAI21_X1 U16445 ( .B1(n6872), .B2(n14780), .A(n14779), .ZN(n14782) );
  AOI211_X1 U16446 ( .C1(n14784), .C2(n14783), .A(n14782), .B(n14781), .ZN(
        n14797) );
  INV_X1 U16447 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14786) );
  AOI22_X1 U16448 ( .A1(n14748), .A2(n14797), .B1(n14786), .B2(n14785), .ZN(
        P1_U3489) );
  AOI22_X1 U16449 ( .A1(n14798), .A2(n14788), .B1(n14787), .B2(n14796), .ZN(
        P1_U3529) );
  INV_X1 U16450 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14789) );
  AOI22_X1 U16451 ( .A1(n14798), .A2(n14790), .B1(n14789), .B2(n14796), .ZN(
        P1_U3533) );
  INV_X1 U16452 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14791) );
  AOI22_X1 U16453 ( .A1(n14798), .A2(n14792), .B1(n14791), .B2(n14796), .ZN(
        P1_U3534) );
  AOI22_X1 U16454 ( .A1(n14798), .A2(n14793), .B1(n9387), .B2(n14796), .ZN(
        P1_U3535) );
  AOI22_X1 U16455 ( .A1(n14798), .A2(n14794), .B1(n9476), .B2(n14796), .ZN(
        P1_U3536) );
  AOI22_X1 U16456 ( .A1(n14798), .A2(n14795), .B1(n9666), .B2(n14796), .ZN(
        P1_U3537) );
  AOI22_X1 U16457 ( .A1(n14798), .A2(n14797), .B1(n9979), .B2(n14796), .ZN(
        P1_U3538) );
  NOR2_X1 U16458 ( .A1(n14821), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI22_X1 U16459 ( .A1(n14802), .A2(n14801), .B1(n14800), .B2(n14799), .ZN(
        n14811) );
  INV_X1 U16460 ( .A(n14804), .ZN(n14806) );
  MUX2_X1 U16461 ( .A(n14803), .B(n14806), .S(n14805), .Z(n14807) );
  AOI211_X1 U16462 ( .C1(n14809), .C2(n14803), .A(n14808), .B(n14807), .ZN(
        n14810) );
  AOI211_X1 U16463 ( .C1(n14813), .C2(n14812), .A(n14811), .B(n14810), .ZN(
        n14814) );
  NAND2_X1 U16464 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n14872)
         );
  OAI211_X1 U16465 ( .C1(n14816), .C2(n14815), .A(n14814), .B(n14872), .ZN(
        P2_U3196) );
  AOI22_X1 U16466 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n14910), .B1(n14876), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n14820) );
  AOI22_X1 U16467 ( .A1(n14821), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14819) );
  OAI22_X1 U16468 ( .A1(n14852), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n14901), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n14817) );
  OAI21_X1 U16469 ( .B1(n14908), .B2(n14817), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14818) );
  OAI211_X1 U16470 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14820), .A(n14819), .B(
        n14818), .ZN(P2_U3214) );
  AOI22_X1 U16471 ( .A1(n14821), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14833) );
  XNOR2_X1 U16472 ( .A(n14823), .B(n14822), .ZN(n14825) );
  AOI22_X1 U16473 ( .A1(n14876), .A2(n14825), .B1(n6482), .B2(n14908), .ZN(
        n14832) );
  AND2_X1 U16474 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n14830) );
  INV_X1 U16475 ( .A(n14826), .ZN(n14829) );
  INV_X1 U16476 ( .A(n14827), .ZN(n14828) );
  OAI211_X1 U16477 ( .C1(n14830), .C2(n14829), .A(n14910), .B(n14828), .ZN(
        n14831) );
  NAND3_X1 U16478 ( .A1(n14833), .A2(n14832), .A3(n14831), .ZN(P2_U3215) );
  AOI211_X1 U16479 ( .C1(n14836), .C2(n14835), .A(n14834), .B(n14901), .ZN(
        n14841) );
  OAI22_X1 U16480 ( .A1(n14839), .A2(n14838), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14837), .ZN(n14840) );
  NOR2_X1 U16481 ( .A1(n14841), .A2(n14840), .ZN(n14847) );
  AOI211_X1 U16482 ( .C1(n14844), .C2(n14843), .A(n14842), .B(n14852), .ZN(
        n14845) );
  INV_X1 U16483 ( .A(n14845), .ZN(n14846) );
  OAI211_X1 U16484 ( .C1(n14916), .C2(n14848), .A(n14847), .B(n14846), .ZN(
        P2_U3216) );
  AOI21_X1 U16485 ( .B1(n14851), .B2(n14850), .A(n14849), .ZN(n14853) );
  NOR2_X1 U16486 ( .A1(n14853), .A2(n14852), .ZN(n14858) );
  AOI211_X1 U16487 ( .C1(n14856), .C2(n14855), .A(n14901), .B(n14854), .ZN(
        n14857) );
  AOI211_X1 U16488 ( .C1(n14908), .C2(n14859), .A(n14858), .B(n14857), .ZN(
        n14861) );
  OAI211_X1 U16489 ( .C1(n15291), .C2(n14916), .A(n14861), .B(n14860), .ZN(
        P2_U3225) );
  AOI21_X1 U16490 ( .B1(n14864), .B2(n14863), .A(n14862), .ZN(n14865) );
  INV_X1 U16491 ( .A(n14865), .ZN(n14871) );
  OAI21_X1 U16492 ( .B1(n14868), .B2(n14867), .A(n14866), .ZN(n14870) );
  AOI222_X1 U16493 ( .A1(n14871), .A2(n14910), .B1(n14876), .B2(n14870), .C1(
        n14869), .C2(n14908), .ZN(n14873) );
  OAI211_X1 U16494 ( .C1(n14874), .C2(n14916), .A(n14873), .B(n14872), .ZN(
        P2_U3226) );
  NOR2_X1 U16495 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14875), .ZN(n14881) );
  OAI211_X1 U16496 ( .C1(n14878), .C2(n14877), .A(n14876), .B(n6593), .ZN(
        n14879) );
  INV_X1 U16497 ( .A(n14879), .ZN(n14880) );
  AOI211_X1 U16498 ( .C1(n14908), .C2(n14882), .A(n14881), .B(n14880), .ZN(
        n14886) );
  OAI211_X1 U16499 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n14884), .A(n14910), 
        .B(n14883), .ZN(n14885) );
  OAI211_X1 U16500 ( .C1(n14916), .C2(n14887), .A(n14886), .B(n14885), .ZN(
        P2_U3228) );
  INV_X1 U16501 ( .A(n14888), .ZN(n14893) );
  AOI211_X1 U16502 ( .C1(n14891), .C2(n14890), .A(n14889), .B(n14901), .ZN(
        n14892) );
  AOI211_X1 U16503 ( .C1(n14894), .C2(n14908), .A(n14893), .B(n14892), .ZN(
        n14899) );
  OAI211_X1 U16504 ( .C1(n14897), .C2(n14896), .A(n14910), .B(n14895), .ZN(
        n14898) );
  OAI211_X1 U16505 ( .C1(n14916), .C2(n14900), .A(n14899), .B(n14898), .ZN(
        P2_U3230) );
  NOR2_X1 U16506 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15265), .ZN(n14906) );
  AOI211_X1 U16507 ( .C1(n14904), .C2(n14903), .A(n14902), .B(n14901), .ZN(
        n14905) );
  AOI211_X1 U16508 ( .C1(n14908), .C2(n14907), .A(n14906), .B(n14905), .ZN(
        n14914) );
  OAI211_X1 U16509 ( .C1(n14912), .C2(n14911), .A(n14910), .B(n14909), .ZN(
        n14913) );
  OAI211_X1 U16510 ( .C1(n14916), .C2(n14915), .A(n14914), .B(n14913), .ZN(
        P2_U3231) );
  NOR2_X1 U16511 ( .A1(n14922), .A2(n14917), .ZN(n14918) );
  AND2_X1 U16512 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14919), .ZN(P2_U3266) );
  AND2_X1 U16513 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14919), .ZN(P2_U3267) );
  INV_X1 U16514 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15256) );
  NOR2_X1 U16515 ( .A1(n14918), .A2(n15256), .ZN(P2_U3268) );
  AND2_X1 U16516 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14919), .ZN(P2_U3269) );
  AND2_X1 U16517 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14919), .ZN(P2_U3270) );
  AND2_X1 U16518 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14919), .ZN(P2_U3271) );
  AND2_X1 U16519 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14919), .ZN(P2_U3272) );
  AND2_X1 U16520 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14919), .ZN(P2_U3273) );
  AND2_X1 U16521 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14919), .ZN(P2_U3274) );
  AND2_X1 U16522 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14919), .ZN(P2_U3275) );
  AND2_X1 U16523 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14919), .ZN(P2_U3276) );
  AND2_X1 U16524 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14919), .ZN(P2_U3277) );
  AND2_X1 U16525 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14919), .ZN(P2_U3278) );
  AND2_X1 U16526 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14919), .ZN(P2_U3279) );
  AND2_X1 U16527 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14919), .ZN(P2_U3280) );
  AND2_X1 U16528 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14919), .ZN(P2_U3281) );
  AND2_X1 U16529 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14919), .ZN(P2_U3282) );
  AND2_X1 U16530 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14919), .ZN(P2_U3283) );
  AND2_X1 U16531 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14919), .ZN(P2_U3284) );
  AND2_X1 U16532 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14919), .ZN(P2_U3285) );
  AND2_X1 U16533 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14919), .ZN(P2_U3286) );
  AND2_X1 U16534 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14919), .ZN(P2_U3287) );
  AND2_X1 U16535 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14919), .ZN(P2_U3288) );
  AND2_X1 U16536 ( .A1(n14919), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3289) );
  AND2_X1 U16537 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14919), .ZN(P2_U3290) );
  AND2_X1 U16538 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14919), .ZN(P2_U3291) );
  AND2_X1 U16539 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14919), .ZN(P2_U3292) );
  AND2_X1 U16540 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14919), .ZN(P2_U3293) );
  AND2_X1 U16541 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14919), .ZN(P2_U3294) );
  AND2_X1 U16542 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14919), .ZN(P2_U3295) );
  OAI21_X1 U16543 ( .B1(n14925), .B2(n14921), .A(n14920), .ZN(P2_U3416) );
  AOI22_X1 U16544 ( .A1(n14925), .A2(n14924), .B1(n14923), .B2(n14922), .ZN(
        P2_U3417) );
  OAI211_X1 U16545 ( .C1(n14928), .C2(n14942), .A(n14927), .B(n14926), .ZN(
        n14975) );
  OAI22_X1 U16546 ( .A1(n14973), .A2(n14975), .B1(P2_REG0_REG_0__SCAN_IN), 
        .B2(n14974), .ZN(n14929) );
  INV_X1 U16547 ( .A(n14929), .ZN(P2_U3430) );
  INV_X1 U16548 ( .A(n14934), .ZN(n14936) );
  AOI211_X1 U16549 ( .C1(n14939), .C2(n14932), .A(n14931), .B(n14930), .ZN(
        n14933) );
  OAI21_X1 U16550 ( .B1(n14942), .B2(n14934), .A(n14933), .ZN(n14935) );
  AOI21_X1 U16551 ( .B1(n14946), .B2(n14936), .A(n14935), .ZN(n14977) );
  AOI22_X1 U16552 ( .A1(n14974), .A2(n14977), .B1(n8627), .B2(n14973), .ZN(
        P2_U3445) );
  INV_X1 U16553 ( .A(n14943), .ZN(n14945) );
  AOI21_X1 U16554 ( .B1(n14939), .B2(n14938), .A(n14937), .ZN(n14940) );
  OAI211_X1 U16555 ( .C1(n14943), .C2(n14942), .A(n14941), .B(n14940), .ZN(
        n14944) );
  AOI21_X1 U16556 ( .B1(n14946), .B2(n14945), .A(n14944), .ZN(n14979) );
  AOI22_X1 U16557 ( .A1(n14974), .A2(n14979), .B1(n8635), .B2(n14973), .ZN(
        P2_U3448) );
  OAI21_X1 U16558 ( .B1(n14948), .B2(n14967), .A(n14947), .ZN(n14950) );
  AOI211_X1 U16559 ( .C1(n14952), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        n14981) );
  AOI22_X1 U16560 ( .A1(n14974), .A2(n14981), .B1(n8662), .B2(n14973), .ZN(
        P2_U3451) );
  INV_X1 U16561 ( .A(n14953), .ZN(n14958) );
  OAI21_X1 U16562 ( .B1(n14955), .B2(n14967), .A(n14954), .ZN(n14957) );
  AOI211_X1 U16563 ( .C1(n14972), .C2(n14958), .A(n14957), .B(n14956), .ZN(
        n14982) );
  AOI22_X1 U16564 ( .A1(n14974), .A2(n14982), .B1(n8680), .B2(n14973), .ZN(
        P2_U3454) );
  INV_X1 U16565 ( .A(n14959), .ZN(n14964) );
  OAI21_X1 U16566 ( .B1(n14961), .B2(n14967), .A(n14960), .ZN(n14963) );
  AOI211_X1 U16567 ( .C1(n14972), .C2(n14964), .A(n14963), .B(n14962), .ZN(
        n14983) );
  AOI22_X1 U16568 ( .A1(n14974), .A2(n14983), .B1(n8702), .B2(n14973), .ZN(
        P2_U3457) );
  INV_X1 U16569 ( .A(n14965), .ZN(n14971) );
  OAI21_X1 U16570 ( .B1(n14968), .B2(n14967), .A(n14966), .ZN(n14970) );
  AOI211_X1 U16571 ( .C1(n14972), .C2(n14971), .A(n14970), .B(n14969), .ZN(
        n14985) );
  AOI22_X1 U16572 ( .A1(n14974), .A2(n14985), .B1(n8719), .B2(n14973), .ZN(
        P2_U3460) );
  OAI22_X1 U16573 ( .A1(n14984), .A2(n14975), .B1(P2_REG1_REG_0__SCAN_IN), 
        .B2(n14986), .ZN(n14976) );
  INV_X1 U16574 ( .A(n14976), .ZN(P2_U3499) );
  AOI22_X1 U16575 ( .A1(n14986), .A2(n14977), .B1(n9454), .B2(n14984), .ZN(
        P2_U3504) );
  INV_X1 U16576 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14978) );
  AOI22_X1 U16577 ( .A1(n14986), .A2(n14979), .B1(n14978), .B2(n14984), .ZN(
        P2_U3505) );
  INV_X1 U16578 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n14980) );
  AOI22_X1 U16579 ( .A1(n14986), .A2(n14981), .B1(n14980), .B2(n14984), .ZN(
        P2_U3506) );
  AOI22_X1 U16580 ( .A1(n14986), .A2(n14982), .B1(n9847), .B2(n14984), .ZN(
        P2_U3507) );
  AOI22_X1 U16581 ( .A1(n14986), .A2(n14983), .B1(n10121), .B2(n14984), .ZN(
        P2_U3508) );
  AOI22_X1 U16582 ( .A1(n14986), .A2(n14985), .B1(n10659), .B2(n14984), .ZN(
        P2_U3509) );
  NOR2_X1 U16583 ( .A1(P3_U3897), .A2(n14987), .ZN(P3_U3150) );
  AOI21_X1 U16584 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n15009) );
  OAI22_X1 U16585 ( .A1(n14994), .A2(n14993), .B1(n14992), .B2(n14991), .ZN(
        n15005) );
  AOI21_X1 U16586 ( .B1(n15259), .B2(n14996), .A(n14995), .ZN(n15003) );
  AOI21_X1 U16587 ( .B1(n14999), .B2(n14998), .A(n14997), .ZN(n15001) );
  OAI22_X1 U16588 ( .A1(n15003), .A2(n15002), .B1(n15001), .B2(n15000), .ZN(
        n15004) );
  NOR3_X1 U16589 ( .A1(n15006), .A2(n15005), .A3(n15004), .ZN(n15007) );
  OAI21_X1 U16590 ( .B1(n15009), .B2(n15008), .A(n15007), .ZN(P3_U3195) );
  INV_X1 U16591 ( .A(n15010), .ZN(n15013) );
  OAI21_X1 U16592 ( .B1(n15013), .B2(n15012), .A(n15011), .ZN(n15018) );
  AOI222_X1 U16593 ( .A1(n15018), .A2(n15030), .B1(n15017), .B2(n15016), .C1(
        n15015), .C2(n15014), .ZN(n15019) );
  OAI21_X1 U16594 ( .B1(n15030), .B2(n15020), .A(n15019), .ZN(P3_U3223) );
  INV_X1 U16595 ( .A(n15021), .ZN(n15028) );
  OAI22_X1 U16596 ( .A1(n15025), .A2(n15024), .B1(n15023), .B2(n15022), .ZN(
        n15027) );
  AOI211_X1 U16597 ( .C1(n15029), .C2(n15028), .A(n15027), .B(n15026), .ZN(
        n15031) );
  AOI22_X1 U16598 ( .A1(n15032), .A2(n10163), .B1(n15031), .B2(n15030), .ZN(
        P3_U3231) );
  OAI21_X1 U16599 ( .B1(n15035), .B2(n15034), .A(n15033), .ZN(n15036) );
  NOR2_X1 U16600 ( .A1(n15037), .A2(n15036), .ZN(n15091) );
  INV_X1 U16601 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n15038) );
  AOI22_X1 U16602 ( .A1(n15089), .A2(n15091), .B1(n15038), .B2(n15087), .ZN(
        P3_U3393) );
  INV_X1 U16603 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15039) );
  AOI22_X1 U16604 ( .A1(n15089), .A2(n15040), .B1(n15039), .B2(n15087), .ZN(
        P3_U3396) );
  NAND2_X1 U16605 ( .A1(n15046), .A2(n15041), .ZN(n15042) );
  OAI211_X1 U16606 ( .C1(n15079), .C2(n15044), .A(n15043), .B(n15042), .ZN(
        n15045) );
  AOI21_X1 U16607 ( .B1(n15046), .B2(n15085), .A(n15045), .ZN(n15093) );
  AOI22_X1 U16608 ( .A1(n15089), .A2(n15093), .B1(n7551), .B2(n15087), .ZN(
        P3_U3399) );
  AOI21_X1 U16609 ( .B1(n15061), .B2(n15081), .A(n15047), .ZN(n15050) );
  INV_X1 U16610 ( .A(n15048), .ZN(n15049) );
  AOI211_X1 U16611 ( .C1(n15051), .C2(n15065), .A(n15050), .B(n15049), .ZN(
        n15095) );
  INV_X1 U16612 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15052) );
  AOI22_X1 U16613 ( .A1(n15089), .A2(n15095), .B1(n15052), .B2(n15087), .ZN(
        P3_U3402) );
  AOI21_X1 U16614 ( .B1(n15061), .B2(n15081), .A(n15053), .ZN(n15056) );
  INV_X1 U16615 ( .A(n15054), .ZN(n15055) );
  AOI211_X1 U16616 ( .C1(n15057), .C2(n15065), .A(n15056), .B(n15055), .ZN(
        n15097) );
  INV_X1 U16617 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U16618 ( .A1(n15089), .A2(n15097), .B1(n15058), .B2(n15087), .ZN(
        P3_U3405) );
  INV_X1 U16619 ( .A(n15059), .ZN(n15063) );
  AOI21_X1 U16620 ( .B1(n15061), .B2(n15081), .A(n15060), .ZN(n15062) );
  AOI211_X1 U16621 ( .C1(n15065), .C2(n15064), .A(n15063), .B(n15062), .ZN(
        n15099) );
  INV_X1 U16622 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15066) );
  AOI22_X1 U16623 ( .A1(n15089), .A2(n15099), .B1(n15066), .B2(n15087), .ZN(
        P3_U3408) );
  OAI22_X1 U16624 ( .A1(n15068), .A2(n15081), .B1(n15067), .B2(n15079), .ZN(
        n15069) );
  NOR2_X1 U16625 ( .A1(n15070), .A2(n15069), .ZN(n15101) );
  INV_X1 U16626 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15071) );
  AOI22_X1 U16627 ( .A1(n15089), .A2(n15101), .B1(n15071), .B2(n15087), .ZN(
        P3_U3411) );
  INV_X1 U16628 ( .A(n15073), .ZN(n15077) );
  OAI22_X1 U16629 ( .A1(n15073), .A2(n15081), .B1(n15072), .B2(n15079), .ZN(
        n15076) );
  INV_X1 U16630 ( .A(n15074), .ZN(n15075) );
  AOI211_X1 U16631 ( .C1(n15077), .C2(n15085), .A(n15076), .B(n15075), .ZN(
        n15103) );
  INV_X1 U16632 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15078) );
  AOI22_X1 U16633 ( .A1(n15089), .A2(n15103), .B1(n15078), .B2(n15087), .ZN(
        P3_U3414) );
  INV_X1 U16634 ( .A(n15082), .ZN(n15086) );
  OAI22_X1 U16635 ( .A1(n15082), .A2(n15081), .B1(n15080), .B2(n15079), .ZN(
        n15084) );
  AOI211_X1 U16636 ( .C1(n15086), .C2(n15085), .A(n15084), .B(n15083), .ZN(
        n15105) );
  INV_X1 U16637 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15088) );
  AOI22_X1 U16638 ( .A1(n15089), .A2(n15105), .B1(n15088), .B2(n15087), .ZN(
        P3_U3417) );
  AOI22_X1 U16639 ( .A1(n15106), .A2(n15091), .B1(n15090), .B2(n15104), .ZN(
        P3_U3460) );
  AOI22_X1 U16640 ( .A1(n15106), .A2(n15093), .B1(n15092), .B2(n15104), .ZN(
        P3_U3462) );
  AOI22_X1 U16641 ( .A1(n15106), .A2(n15095), .B1(n15094), .B2(n15104), .ZN(
        P3_U3463) );
  AOI22_X1 U16642 ( .A1(n15106), .A2(n15097), .B1(n15096), .B2(n15104), .ZN(
        P3_U3464) );
  AOI22_X1 U16643 ( .A1(n15106), .A2(n15099), .B1(n15098), .B2(n15104), .ZN(
        P3_U3465) );
  AOI22_X1 U16644 ( .A1(n15106), .A2(n15101), .B1(n15100), .B2(n15104), .ZN(
        P3_U3466) );
  AOI22_X1 U16645 ( .A1(n15106), .A2(n15103), .B1(n15102), .B2(n15104), .ZN(
        P3_U3467) );
  AOI22_X1 U16646 ( .A1(n15106), .A2(n15105), .B1(n10397), .B2(n15104), .ZN(
        P3_U3468) );
  AOI22_X1 U16647 ( .A1(n7422), .A2(keyinput122), .B1(keyinput79), .B2(n8549), 
        .ZN(n15107) );
  OAI221_X1 U16648 ( .B1(n7422), .B2(keyinput122), .C1(n8549), .C2(keyinput79), 
        .A(n15107), .ZN(n15116) );
  AOI22_X1 U16649 ( .A1(n11996), .A2(keyinput116), .B1(n15109), .B2(
        keyinput111), .ZN(n15108) );
  OAI221_X1 U16650 ( .B1(n11996), .B2(keyinput116), .C1(n15109), .C2(
        keyinput111), .A(n15108), .ZN(n15115) );
  AOI22_X1 U16651 ( .A1(n15231), .A2(keyinput71), .B1(keyinput109), .B2(n15249), .ZN(n15110) );
  OAI221_X1 U16652 ( .B1(n15231), .B2(keyinput71), .C1(n15249), .C2(
        keyinput109), .A(n15110), .ZN(n15114) );
  AOI22_X1 U16653 ( .A1(n15238), .A2(keyinput85), .B1(keyinput73), .B2(n15112), 
        .ZN(n15111) );
  OAI221_X1 U16654 ( .B1(n15238), .B2(keyinput85), .C1(n15112), .C2(keyinput73), .A(n15111), .ZN(n15113) );
  NOR4_X1 U16655 ( .A1(n15116), .A2(n15115), .A3(n15114), .A4(n15113), .ZN(
        n15156) );
  AOI22_X1 U16656 ( .A1(n15118), .A2(keyinput76), .B1(keyinput81), .B2(n15241), 
        .ZN(n15117) );
  OAI221_X1 U16657 ( .B1(n15118), .B2(keyinput76), .C1(n15241), .C2(keyinput81), .A(n15117), .ZN(n15126) );
  AOI22_X1 U16658 ( .A1(P1_REG1_REG_1__SCAN_IN), .A2(keyinput127), .B1(
        P1_D_REG_9__SCAN_IN), .B2(keyinput100), .ZN(n15119) );
  OAI221_X1 U16659 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(keyinput127), .C1(
        P1_D_REG_9__SCAN_IN), .C2(keyinput100), .A(n15119), .ZN(n15125) );
  XNOR2_X1 U16660 ( .A(P3_REG3_REG_9__SCAN_IN), .B(keyinput126), .ZN(n15123)
         );
  XNOR2_X1 U16661 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput72), .ZN(n15122) );
  XNOR2_X1 U16662 ( .A(P3_IR_REG_28__SCAN_IN), .B(keyinput113), .ZN(n15121) );
  XNOR2_X1 U16663 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput77), .ZN(n15120)
         );
  NAND4_X1 U16664 ( .A1(n15123), .A2(n15122), .A3(n15121), .A4(n15120), .ZN(
        n15124) );
  NOR3_X1 U16665 ( .A1(n15126), .A2(n15125), .A3(n15124), .ZN(n15155) );
  AOI22_X1 U16666 ( .A1(n15248), .A2(keyinput75), .B1(n15128), .B2(keyinput66), 
        .ZN(n15127) );
  OAI221_X1 U16667 ( .B1(n15248), .B2(keyinput75), .C1(n15128), .C2(keyinput66), .A(n15127), .ZN(n15138) );
  INV_X1 U16668 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n15257) );
  AOI22_X1 U16669 ( .A1(n15274), .A2(keyinput107), .B1(keyinput86), .B2(n15257), .ZN(n15129) );
  OAI221_X1 U16670 ( .B1(n15274), .B2(keyinput107), .C1(n15257), .C2(
        keyinput86), .A(n15129), .ZN(n15137) );
  AOI22_X1 U16671 ( .A1(n15132), .A2(keyinput94), .B1(n15131), .B2(keyinput68), 
        .ZN(n15130) );
  OAI221_X1 U16672 ( .B1(n15132), .B2(keyinput94), .C1(n15131), .C2(keyinput68), .A(n15130), .ZN(n15136) );
  XNOR2_X1 U16673 ( .A(P3_IR_REG_5__SCAN_IN), .B(keyinput82), .ZN(n15134) );
  XNOR2_X1 U16674 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput118), .ZN(n15133) );
  NAND2_X1 U16675 ( .A1(n15134), .A2(n15133), .ZN(n15135) );
  NOR4_X1 U16676 ( .A1(n15138), .A2(n15137), .A3(n15136), .A4(n15135), .ZN(
        n15154) );
  AOI22_X1 U16677 ( .A1(n15141), .A2(keyinput87), .B1(keyinput96), .B2(n15140), 
        .ZN(n15139) );
  OAI221_X1 U16678 ( .B1(n15141), .B2(keyinput87), .C1(n15140), .C2(keyinput96), .A(n15139), .ZN(n15152) );
  AOI22_X1 U16679 ( .A1(n15143), .A2(keyinput93), .B1(keyinput115), .B2(n9776), 
        .ZN(n15142) );
  OAI221_X1 U16680 ( .B1(n15143), .B2(keyinput93), .C1(n9776), .C2(keyinput115), .A(n15142), .ZN(n15151) );
  AOI22_X1 U16681 ( .A1(n15146), .A2(keyinput91), .B1(n15145), .B2(keyinput110), .ZN(n15144) );
  OAI221_X1 U16682 ( .B1(n15146), .B2(keyinput91), .C1(n15145), .C2(
        keyinput110), .A(n15144), .ZN(n15150) );
  XOR2_X1 U16683 ( .A(n15271), .B(keyinput114), .Z(n15148) );
  XNOR2_X1 U16684 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput125), .ZN(n15147) );
  NAND2_X1 U16685 ( .A1(n15148), .A2(n15147), .ZN(n15149) );
  NOR4_X1 U16686 ( .A1(n15152), .A2(n15151), .A3(n15150), .A4(n15149), .ZN(
        n15153) );
  AND4_X1 U16687 ( .A1(n15156), .A2(n15155), .A3(n15154), .A4(n15153), .ZN(
        n15289) );
  OAI22_X1 U16688 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(keyinput98), .B1(
        P3_DATAO_REG_21__SCAN_IN), .B2(keyinput83), .ZN(n15157) );
  AOI221_X1 U16689 ( .B1(P1_DATAO_REG_19__SCAN_IN), .B2(keyinput98), .C1(
        keyinput83), .C2(P3_DATAO_REG_21__SCAN_IN), .A(n15157), .ZN(n15164) );
  OAI22_X1 U16690 ( .A1(P3_REG2_REG_29__SCAN_IN), .A2(keyinput74), .B1(
        P3_REG0_REG_25__SCAN_IN), .B2(keyinput64), .ZN(n15158) );
  AOI221_X1 U16691 ( .B1(P3_REG2_REG_29__SCAN_IN), .B2(keyinput74), .C1(
        keyinput64), .C2(P3_REG0_REG_25__SCAN_IN), .A(n15158), .ZN(n15163) );
  OAI22_X1 U16692 ( .A1(SI_5_), .A2(keyinput99), .B1(P2_IR_REG_19__SCAN_IN), 
        .B2(keyinput123), .ZN(n15159) );
  AOI221_X1 U16693 ( .B1(SI_5_), .B2(keyinput99), .C1(keyinput123), .C2(
        P2_IR_REG_19__SCAN_IN), .A(n15159), .ZN(n15162) );
  OAI22_X1 U16694 ( .A1(P2_D_REG_0__SCAN_IN), .A2(keyinput105), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput88), .ZN(n15160) );
  AOI221_X1 U16695 ( .B1(P2_D_REG_0__SCAN_IN), .B2(keyinput105), .C1(
        keyinput88), .C2(P2_REG3_REG_17__SCAN_IN), .A(n15160), .ZN(n15161) );
  NAND4_X1 U16696 ( .A1(n15164), .A2(n15163), .A3(n15162), .A4(n15161), .ZN(
        n15192) );
  OAI22_X1 U16697 ( .A1(P3_D_REG_28__SCAN_IN), .A2(keyinput119), .B1(
        keyinput106), .B2(P2_WR_REG_SCAN_IN), .ZN(n15165) );
  AOI221_X1 U16698 ( .B1(P3_D_REG_28__SCAN_IN), .B2(keyinput119), .C1(
        P2_WR_REG_SCAN_IN), .C2(keyinput106), .A(n15165), .ZN(n15172) );
  OAI22_X1 U16699 ( .A1(P2_REG0_REG_22__SCAN_IN), .A2(keyinput80), .B1(
        keyinput78), .B2(P2_ADDR_REG_14__SCAN_IN), .ZN(n15166) );
  AOI221_X1 U16700 ( .B1(P2_REG0_REG_22__SCAN_IN), .B2(keyinput80), .C1(
        P2_ADDR_REG_14__SCAN_IN), .C2(keyinput78), .A(n15166), .ZN(n15171) );
  OAI22_X1 U16701 ( .A1(P2_REG0_REG_9__SCAN_IN), .A2(keyinput97), .B1(
        P1_ADDR_REG_0__SCAN_IN), .B2(keyinput102), .ZN(n15167) );
  AOI221_X1 U16702 ( .B1(P2_REG0_REG_9__SCAN_IN), .B2(keyinput97), .C1(
        keyinput102), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n15167), .ZN(n15170) );
  OAI22_X1 U16703 ( .A1(P2_D_REG_8__SCAN_IN), .A2(keyinput120), .B1(keyinput95), .B2(P2_REG3_REG_27__SCAN_IN), .ZN(n15168) );
  AOI221_X1 U16704 ( .B1(P2_D_REG_8__SCAN_IN), .B2(keyinput120), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput95), .A(n15168), .ZN(n15169) );
  NAND4_X1 U16705 ( .A1(n15172), .A2(n15171), .A3(n15170), .A4(n15169), .ZN(
        n15191) );
  OAI22_X1 U16706 ( .A1(P3_D_REG_18__SCAN_IN), .A2(keyinput101), .B1(
        P1_REG0_REG_24__SCAN_IN), .B2(keyinput92), .ZN(n15173) );
  AOI221_X1 U16707 ( .B1(P3_D_REG_18__SCAN_IN), .B2(keyinput101), .C1(
        keyinput92), .C2(P1_REG0_REG_24__SCAN_IN), .A(n15173), .ZN(n15180) );
  OAI22_X1 U16708 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(keyinput69), .B1(
        P1_REG1_REG_19__SCAN_IN), .B2(keyinput84), .ZN(n15174) );
  AOI221_X1 U16709 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(keyinput69), .C1(
        keyinput84), .C2(P1_REG1_REG_19__SCAN_IN), .A(n15174), .ZN(n15179) );
  OAI22_X1 U16710 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput65), .B1(
        P1_D_REG_31__SCAN_IN), .B2(keyinput117), .ZN(n15175) );
  AOI221_X1 U16711 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput65), .C1(
        keyinput117), .C2(P1_D_REG_31__SCAN_IN), .A(n15175), .ZN(n15178) );
  OAI22_X1 U16712 ( .A1(P3_REG1_REG_19__SCAN_IN), .A2(keyinput70), .B1(
        keyinput103), .B2(P2_D_REG_29__SCAN_IN), .ZN(n15176) );
  AOI221_X1 U16713 ( .B1(P3_REG1_REG_19__SCAN_IN), .B2(keyinput70), .C1(
        P2_D_REG_29__SCAN_IN), .C2(keyinput103), .A(n15176), .ZN(n15177) );
  NAND4_X1 U16714 ( .A1(n15180), .A2(n15179), .A3(n15178), .A4(n15177), .ZN(
        n15190) );
  OAI22_X1 U16715 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(keyinput124), .B1(
        P2_REG2_REG_5__SCAN_IN), .B2(keyinput67), .ZN(n15181) );
  AOI221_X1 U16716 ( .B1(P2_REG2_REG_24__SCAN_IN), .B2(keyinput124), .C1(
        keyinput67), .C2(P2_REG2_REG_5__SCAN_IN), .A(n15181), .ZN(n15188) );
  OAI22_X1 U16717 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(keyinput104), .B1(
        keyinput90), .B2(P3_REG2_REG_31__SCAN_IN), .ZN(n15182) );
  AOI221_X1 U16718 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput104), .C1(
        P3_REG2_REG_31__SCAN_IN), .C2(keyinput90), .A(n15182), .ZN(n15187) );
  OAI22_X1 U16719 ( .A1(P1_D_REG_26__SCAN_IN), .A2(keyinput121), .B1(
        keyinput108), .B2(P1_REG0_REG_25__SCAN_IN), .ZN(n15183) );
  AOI221_X1 U16720 ( .B1(P1_D_REG_26__SCAN_IN), .B2(keyinput121), .C1(
        P1_REG0_REG_25__SCAN_IN), .C2(keyinput108), .A(n15183), .ZN(n15186) );
  OAI22_X1 U16721 ( .A1(P3_REG0_REG_14__SCAN_IN), .A2(keyinput112), .B1(
        P1_REG1_REG_17__SCAN_IN), .B2(keyinput89), .ZN(n15184) );
  AOI221_X1 U16722 ( .B1(P3_REG0_REG_14__SCAN_IN), .B2(keyinput112), .C1(
        keyinput89), .C2(P1_REG1_REG_17__SCAN_IN), .A(n15184), .ZN(n15185) );
  NAND4_X1 U16723 ( .A1(n15188), .A2(n15187), .A3(n15186), .A4(n15185), .ZN(
        n15189) );
  NOR4_X1 U16724 ( .A1(n15192), .A2(n15191), .A3(n15190), .A4(n15189), .ZN(
        n15288) );
  AOI22_X1 U16725 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput8), .B1(
        P3_REG2_REG_31__SCAN_IN), .B2(keyinput26), .ZN(n15193) );
  OAI221_X1 U16726 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput8), .C1(
        P3_REG2_REG_31__SCAN_IN), .C2(keyinput26), .A(n15193), .ZN(n15200) );
  AOI22_X1 U16727 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput30), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(keyinput29), .ZN(n15194) );
  OAI221_X1 U16728 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput30), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput29), .A(n15194), .ZN(n15199) );
  AOI22_X1 U16729 ( .A1(P3_DATAO_REG_1__SCAN_IN), .A2(keyinput27), .B1(
        P1_REG1_REG_17__SCAN_IN), .B2(keyinput25), .ZN(n15195) );
  OAI221_X1 U16730 ( .B1(P3_DATAO_REG_1__SCAN_IN), .B2(keyinput27), .C1(
        P1_REG1_REG_17__SCAN_IN), .C2(keyinput25), .A(n15195), .ZN(n15198) );
  AOI22_X1 U16731 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput23), .B1(
        P3_D_REG_18__SCAN_IN), .B2(keyinput37), .ZN(n15196) );
  OAI221_X1 U16732 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput23), .C1(
        P3_D_REG_18__SCAN_IN), .C2(keyinput37), .A(n15196), .ZN(n15197) );
  NOR4_X1 U16733 ( .A1(n15200), .A2(n15199), .A3(n15198), .A4(n15197), .ZN(
        n15228) );
  AOI22_X1 U16734 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput1), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput12), .ZN(n15201) );
  OAI221_X1 U16735 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput1), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput12), .A(n15201), .ZN(n15208) );
  AOI22_X1 U16736 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(keyinput38), .B1(SI_5_), 
        .B2(keyinput35), .ZN(n15202) );
  OAI221_X1 U16737 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(keyinput38), .C1(SI_5_), 
        .C2(keyinput35), .A(n15202), .ZN(n15207) );
  AOI22_X1 U16738 ( .A1(P2_D_REG_0__SCAN_IN), .A2(keyinput41), .B1(
        P3_REG0_REG_25__SCAN_IN), .B2(keyinput0), .ZN(n15203) );
  OAI221_X1 U16739 ( .B1(P2_D_REG_0__SCAN_IN), .B2(keyinput41), .C1(
        P3_REG0_REG_25__SCAN_IN), .C2(keyinput0), .A(n15203), .ZN(n15206) );
  AOI22_X1 U16740 ( .A1(P3_DATAO_REG_10__SCAN_IN), .A2(keyinput32), .B1(
        P3_REG2_REG_29__SCAN_IN), .B2(keyinput10), .ZN(n15204) );
  OAI221_X1 U16741 ( .B1(P3_DATAO_REG_10__SCAN_IN), .B2(keyinput32), .C1(
        P3_REG2_REG_29__SCAN_IN), .C2(keyinput10), .A(n15204), .ZN(n15205) );
  NOR4_X1 U16742 ( .A1(n15208), .A2(n15207), .A3(n15206), .A4(n15205), .ZN(
        n15227) );
  AOI22_X1 U16743 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(keyinput4), .B1(
        P2_IR_REG_31__SCAN_IN), .B2(keyinput61), .ZN(n15209) );
  OAI221_X1 U16744 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(keyinput4), .C1(
        P2_IR_REG_31__SCAN_IN), .C2(keyinput61), .A(n15209), .ZN(n15216) );
  AOI22_X1 U16745 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(keyinput46), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(keyinput34), .ZN(n15210) );
  OAI221_X1 U16746 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(keyinput46), .C1(
        P1_DATAO_REG_19__SCAN_IN), .C2(keyinput34), .A(n15210), .ZN(n15215) );
  AOI22_X1 U16747 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(keyinput9), .B1(
        P3_REG0_REG_14__SCAN_IN), .B2(keyinput48), .ZN(n15211) );
  OAI221_X1 U16748 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(keyinput9), .C1(
        P3_REG0_REG_14__SCAN_IN), .C2(keyinput48), .A(n15211), .ZN(n15214) );
  AOI22_X1 U16749 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput31), .B1(
        P3_IR_REG_5__SCAN_IN), .B2(keyinput18), .ZN(n15212) );
  OAI221_X1 U16750 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput31), .C1(
        P3_IR_REG_5__SCAN_IN), .C2(keyinput18), .A(n15212), .ZN(n15213) );
  NOR4_X1 U16751 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        n15226) );
  AOI22_X1 U16752 ( .A1(P1_REG1_REG_19__SCAN_IN), .A2(keyinput20), .B1(
        P2_REG0_REG_1__SCAN_IN), .B2(keyinput15), .ZN(n15217) );
  OAI221_X1 U16753 ( .B1(P1_REG1_REG_19__SCAN_IN), .B2(keyinput20), .C1(
        P2_REG0_REG_1__SCAN_IN), .C2(keyinput15), .A(n15217), .ZN(n15224) );
  AOI22_X1 U16754 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput42), .B1(
        P2_IR_REG_26__SCAN_IN), .B2(keyinput58), .ZN(n15218) );
  OAI221_X1 U16755 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput42), .C1(
        P2_IR_REG_26__SCAN_IN), .C2(keyinput58), .A(n15218), .ZN(n15223) );
  AOI22_X1 U16756 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(keyinput60), .B1(
        P3_REG2_REG_25__SCAN_IN), .B2(keyinput47), .ZN(n15219) );
  OAI221_X1 U16757 ( .B1(P2_REG2_REG_24__SCAN_IN), .B2(keyinput60), .C1(
        P3_REG2_REG_25__SCAN_IN), .C2(keyinput47), .A(n15219), .ZN(n15222) );
  AOI22_X1 U16758 ( .A1(P1_D_REG_26__SCAN_IN), .A2(keyinput57), .B1(
        P3_D_REG_28__SCAN_IN), .B2(keyinput55), .ZN(n15220) );
  OAI221_X1 U16759 ( .B1(P1_D_REG_26__SCAN_IN), .B2(keyinput57), .C1(
        P3_D_REG_28__SCAN_IN), .C2(keyinput55), .A(n15220), .ZN(n15221) );
  NOR4_X1 U16760 ( .A1(n15224), .A2(n15223), .A3(n15222), .A4(n15221), .ZN(
        n15225) );
  NAND4_X1 U16761 ( .A1(n15228), .A2(n15227), .A3(n15226), .A4(n15225), .ZN(
        n15287) );
  AOI22_X1 U16762 ( .A1(n15231), .A2(keyinput7), .B1(n15230), .B2(keyinput13), 
        .ZN(n15229) );
  OAI221_X1 U16763 ( .B1(n15231), .B2(keyinput7), .C1(n15230), .C2(keyinput13), 
        .A(n15229), .ZN(n15235) );
  XOR2_X1 U16764 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput59), .Z(n15234) );
  XNOR2_X1 U16765 ( .A(n15232), .B(keyinput19), .ZN(n15233) );
  OR3_X1 U16766 ( .A1(n15235), .A2(n15234), .A3(n15233), .ZN(n15244) );
  AOI22_X1 U16767 ( .A1(n15238), .A2(keyinput21), .B1(keyinput36), .B2(n15237), 
        .ZN(n15236) );
  OAI221_X1 U16768 ( .B1(n15238), .B2(keyinput21), .C1(n15237), .C2(keyinput36), .A(n15236), .ZN(n15243) );
  INV_X1 U16769 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n15240) );
  AOI22_X1 U16770 ( .A1(n15241), .A2(keyinput17), .B1(keyinput28), .B2(n15240), 
        .ZN(n15239) );
  OAI221_X1 U16771 ( .B1(n15241), .B2(keyinput17), .C1(n15240), .C2(keyinput28), .A(n15239), .ZN(n15242) );
  NOR3_X1 U16772 ( .A1(n15244), .A2(n15243), .A3(n15242), .ZN(n15285) );
  AOI22_X1 U16773 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(keyinput14), .B1(
        P2_D_REG_8__SCAN_IN), .B2(keyinput56), .ZN(n15245) );
  OAI221_X1 U16774 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(keyinput14), .C1(
        P2_D_REG_8__SCAN_IN), .C2(keyinput56), .A(n15245), .ZN(n15254) );
  AOI22_X1 U16775 ( .A1(P2_REG2_REG_5__SCAN_IN), .A2(keyinput3), .B1(
        P3_REG0_REG_12__SCAN_IN), .B2(keyinput2), .ZN(n15246) );
  OAI221_X1 U16776 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(keyinput3), .C1(
        P3_REG0_REG_12__SCAN_IN), .C2(keyinput2), .A(n15246), .ZN(n15253) );
  AOI22_X1 U16777 ( .A1(n15249), .A2(keyinput45), .B1(n15248), .B2(keyinput11), 
        .ZN(n15247) );
  OAI221_X1 U16778 ( .B1(n15249), .B2(keyinput45), .C1(n15248), .C2(keyinput11), .A(n15247), .ZN(n15252) );
  AOI22_X1 U16779 ( .A1(P1_REG1_REG_1__SCAN_IN), .A2(keyinput63), .B1(
        P3_REG3_REG_9__SCAN_IN), .B2(keyinput62), .ZN(n15250) );
  OAI221_X1 U16780 ( .B1(P1_REG1_REG_1__SCAN_IN), .B2(keyinput63), .C1(
        P3_REG3_REG_9__SCAN_IN), .C2(keyinput62), .A(n15250), .ZN(n15251) );
  NOR4_X1 U16781 ( .A1(n15254), .A2(n15253), .A3(n15252), .A4(n15251), .ZN(
        n15284) );
  AOI22_X1 U16782 ( .A1(n15257), .A2(keyinput22), .B1(n15256), .B2(keyinput39), 
        .ZN(n15255) );
  OAI221_X1 U16783 ( .B1(n15257), .B2(keyinput22), .C1(n15256), .C2(keyinput39), .A(n15255), .ZN(n15269) );
  AOI22_X1 U16784 ( .A1(n15260), .A2(keyinput16), .B1(n15259), .B2(keyinput5), 
        .ZN(n15258) );
  OAI221_X1 U16785 ( .B1(n15260), .B2(keyinput16), .C1(n15259), .C2(keyinput5), 
        .A(n15258), .ZN(n15268) );
  INV_X1 U16786 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15262) );
  AOI22_X1 U16787 ( .A1(n15263), .A2(keyinput53), .B1(n15262), .B2(keyinput40), 
        .ZN(n15261) );
  OAI221_X1 U16788 ( .B1(n15263), .B2(keyinput53), .C1(n15262), .C2(keyinput40), .A(n15261), .ZN(n15267) );
  AOI22_X1 U16789 ( .A1(n15265), .A2(keyinput24), .B1(keyinput52), .B2(n11996), 
        .ZN(n15264) );
  OAI221_X1 U16790 ( .B1(n15265), .B2(keyinput24), .C1(n11996), .C2(keyinput52), .A(n15264), .ZN(n15266) );
  NOR4_X1 U16791 ( .A1(n15269), .A2(n15268), .A3(n15267), .A4(n15266), .ZN(
        n15283) );
  AOI22_X1 U16792 ( .A1(n15271), .A2(keyinput50), .B1(n9776), .B2(keyinput51), 
        .ZN(n15270) );
  OAI221_X1 U16793 ( .B1(n15271), .B2(keyinput50), .C1(n9776), .C2(keyinput51), 
        .A(n15270), .ZN(n15281) );
  AOI22_X1 U16794 ( .A1(n8702), .A2(keyinput33), .B1(n15273), .B2(keyinput6), 
        .ZN(n15272) );
  OAI221_X1 U16795 ( .B1(n8702), .B2(keyinput33), .C1(n15273), .C2(keyinput6), 
        .A(n15272), .ZN(n15280) );
  XOR2_X1 U16796 ( .A(n15274), .B(keyinput43), .Z(n15278) );
  XNOR2_X1 U16797 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput54), .ZN(n15277) );
  XNOR2_X1 U16798 ( .A(P1_REG0_REG_25__SCAN_IN), .B(keyinput44), .ZN(n15276)
         );
  XNOR2_X1 U16799 ( .A(P3_IR_REG_28__SCAN_IN), .B(keyinput49), .ZN(n15275) );
  NAND4_X1 U16800 ( .A1(n15278), .A2(n15277), .A3(n15276), .A4(n15275), .ZN(
        n15279) );
  NOR3_X1 U16801 ( .A1(n15281), .A2(n15280), .A3(n15279), .ZN(n15282) );
  NAND4_X1 U16802 ( .A1(n15285), .A2(n15284), .A3(n15283), .A4(n15282), .ZN(
        n15286) );
  AOI211_X1 U16803 ( .C1(n15289), .C2(n15288), .A(n15287), .B(n15286), .ZN(
        n15290) );
  XNOR2_X1 U16804 ( .A(n15291), .B(n15290), .ZN(n15296) );
  INV_X1 U16805 ( .A(n15292), .ZN(n15293) );
  NAND2_X1 U16806 ( .A1(n15294), .A2(n15293), .ZN(n15295) );
  XNOR2_X1 U16807 ( .A(n15296), .B(n15295), .ZN(SUB_1596_U69) );
  XOR2_X1 U16808 ( .A(n15297), .B(n15298), .Z(SUB_1596_U59) );
  XNOR2_X1 U16809 ( .A(n15299), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16810 ( .B1(n15301), .B2(n15300), .A(n15310), .ZN(SUB_1596_U53) );
  XOR2_X1 U16811 ( .A(n15303), .B(n15302), .Z(SUB_1596_U56) );
  OAI21_X1 U16812 ( .B1(n15306), .B2(n15305), .A(n15304), .ZN(n15308) );
  XOR2_X1 U16813 ( .A(n15308), .B(n15307), .Z(SUB_1596_U60) );
  XOR2_X1 U16814 ( .A(n15310), .B(n15309), .Z(SUB_1596_U5) );
  XNOR2_X1 U7232 ( .A(n10280), .B(n10254), .ZN(n10245) );
  CLKBUF_X3 U7262 ( .A(n7552), .Z(n8107) );
  NAND2_X2 U7276 ( .A1(n12521), .A2(n13141), .ZN(n7550) );
  CLKBUF_X1 U7305 ( .A(n8589), .Z(n9046) );
  CLKBUF_X1 U7337 ( .A(n8063), .Z(n10521) );
  CLKBUF_X1 U7413 ( .A(n8477), .Z(n6485) );
  INV_X1 U8990 ( .A(n8648), .ZN(n8754) );
  INV_X2 U9022 ( .A(n13595), .ZN(n13642) );
endmodule

