

module b20_C_SARLock_k_64_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112;

  NAND2_X1 U4818 ( .A1(n4846), .A2(n4847), .ZN(n5544) );
  OAI21_X1 U4819 ( .B1(n8275), .B2(n8062), .A(n7903), .ZN(n6441) );
  BUF_X1 U4821 ( .A(n5702), .Z(n4315) );
  INV_X2 U4822 ( .A(n5823), .ZN(n5880) );
  INV_X1 U4823 ( .A(n4985), .ZN(n5086) );
  INV_X1 U4824 ( .A(n5702), .ZN(n5654) );
  NAND2_X1 U4827 ( .A1(n4942), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4941) );
  AND2_X1 U4828 ( .A1(n4606), .A2(n4605), .ZN(n4982) );
  AND2_X1 U4829 ( .A1(n6314), .A2(n6313), .ZN(n6315) );
  OR2_X1 U4830 ( .A1(n6991), .A2(n4769), .ZN(n4768) );
  AOI21_X1 U4831 ( .B1(n4429), .B2(n4428), .A(n4426), .ZN(n6457) );
  INV_X1 U4832 ( .A(n7027), .ZN(n6207) );
  AND2_X1 U4833 ( .A1(n7933), .A2(n8100), .ZN(n8085) );
  INV_X2 U4834 ( .A(n5658), .ZN(n5705) );
  AOI21_X1 U4836 ( .B1(n9370), .B2(n9372), .A(n8987), .ZN(n9362) );
  NAND2_X1 U4837 ( .A1(n4312), .A2(n4320), .ZN(n5452) );
  CLKBUF_X2 U4838 ( .A(n5050), .Z(n5101) );
  NOR2_X1 U4839 ( .A1(n7015), .A2(n9761), .ZN(n7095) );
  NAND2_X1 U4840 ( .A1(n6205), .A2(n6206), .ZN(n5829) );
  XNOR2_X1 U4841 ( .A(n6298), .B(n6705), .ZN(n8151) );
  INV_X1 U4842 ( .A(n6054), .ZN(n7893) );
  BUF_X1 U4843 ( .A(n4948), .Z(n9136) );
  NAND2_X1 U4844 ( .A1(n4964), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4966) );
  XNOR2_X1 U4845 ( .A(n4937), .B(P1_IR_REG_19__SCAN_IN), .ZN(n4948) );
  XNOR2_X1 U4846 ( .A(n4966), .B(n4965), .ZN(n7497) );
  XNOR2_X1 U4847 ( .A(n4941), .B(n4943), .ZN(n7342) );
  INV_X2 U4848 ( .A(n5697), .ZN(n4321) );
  OR2_X1 U4849 ( .A1(n6434), .A2(n5735), .ZN(n4311) );
  AND2_X4 U4850 ( .A1(n4998), .A2(n9572), .ZN(n5072) );
  NAND2_X1 U4851 ( .A1(n6711), .A2(n5740), .ZN(n4312) );
  NOR2_X2 U4852 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4929) );
  NAND4_X2 U4853 ( .A1(n5653), .A2(n5652), .A3(n5651), .A4(n5650), .ZN(n9242)
         );
  NOR2_X2 U4854 ( .A1(n4933), .A2(n4932), .ZN(n4934) );
  NAND2_X2 U4855 ( .A1(n7679), .A2(n5815), .ZN(n5823) );
  XNOR2_X2 U4856 ( .A(n5796), .B(n8576), .ZN(n7679) );
  INV_X1 U4857 ( .A(n8098), .ZN(n4313) );
  INV_X1 U4858 ( .A(n8098), .ZN(n4314) );
  INV_X1 U4859 ( .A(n6206), .ZN(n8098) );
  OAI21_X2 U4860 ( .B1(n4842), .B2(n5246), .A(n4841), .ZN(n8634) );
  NAND3_X1 U4861 ( .A1(n4970), .A2(n7094), .A3(n5019), .ZN(n5702) );
  AND2_X1 U4862 ( .A1(n4998), .A2(n4997), .ZN(n5562) );
  NAND2_X1 U4863 ( .A1(n4972), .A2(n5019), .ZN(n5658) );
  AND2_X4 U4864 ( .A1(n5019), .A2(n5003), .ZN(n5697) );
  AOI21_X2 U4865 ( .B1(n4859), .B2(n4858), .A(n4855), .ZN(n6902) );
  XNOR2_X2 U4867 ( .A(n5876), .B(n5875), .ZN(n6856) );
  NAND2_X1 U4868 ( .A1(n4430), .A2(n6459), .ZN(n4318) );
  NAND2_X2 U4869 ( .A1(n4430), .A2(n6459), .ZN(n4319) );
  XNOR2_X1 U4870 ( .A(n5790), .B(n5789), .ZN(n7231) );
  NAND2_X2 U4871 ( .A1(n4349), .A2(n5850), .ZN(n6588) );
  INV_X2 U4872 ( .A(n4982), .ZN(n4320) );
  NOR2_X1 U4873 ( .A1(n8744), .A2(n4431), .ZN(n6434) );
  OAI21_X1 U4874 ( .B1(n4343), .B2(n8746), .A(n8745), .ZN(n8747) );
  AOI21_X1 U4875 ( .B1(n8320), .B2(n7904), .A(n6088), .ZN(n8310) );
  AOI21_X1 U4876 ( .B1(n8387), .B2(n8393), .A(n6043), .ZN(n8372) );
  XNOR2_X1 U4877 ( .A(n4768), .B(n6593), .ZN(n9822) );
  NAND2_X1 U4878 ( .A1(n5731), .A2(n9010), .ZN(n4970) );
  INV_X1 U4879 ( .A(n9749), .ZN(n7699) );
  INV_X1 U4880 ( .A(n9040), .ZN(n6631) );
  INV_X4 U4881 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OAI21_X1 U4882 ( .B1(n8744), .B2(n6431), .A(n6430), .ZN(n6432) );
  AND2_X1 U4883 ( .A1(n5544), .A2(n5543), .ZN(n8713) );
  AND2_X1 U4884 ( .A1(n4473), .A2(n4472), .ZN(n8945) );
  NOR2_X1 U4885 ( .A1(n9398), .A2(n9397), .ZN(n9399) );
  OAI21_X1 U4886 ( .B1(n6428), .B2(n9906), .A(n6427), .ZN(n6429) );
  NAND2_X1 U4887 ( .A1(n4475), .A2(n8936), .ZN(n8941) );
  NAND2_X1 U4888 ( .A1(n7785), .A2(n7787), .ZN(n7739) );
  OAI21_X1 U4889 ( .B1(n4677), .B2(n4681), .A(n4680), .ZN(n8271) );
  NAND2_X1 U4890 ( .A1(n4671), .A2(n4686), .ZN(n8291) );
  NAND2_X1 U4891 ( .A1(n4433), .A2(n4432), .ZN(n4431) );
  INV_X1 U4892 ( .A(n6430), .ZN(n4433) );
  NAND2_X1 U4893 ( .A1(n4435), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4791) );
  INV_X1 U4894 ( .A(n6431), .ZN(n4432) );
  OAI21_X1 U4895 ( .B1(n4704), .B2(n8369), .A(n4702), .ZN(n8338) );
  AOI21_X1 U4896 ( .B1(n4506), .B2(n4786), .A(n8168), .ZN(n8167) );
  OAI21_X1 U4897 ( .B1(n6192), .B2(n4729), .A(n4727), .ZN(n8394) );
  NAND2_X1 U4898 ( .A1(n7634), .A2(n7996), .ZN(n7602) );
  MUX2_X1 U4899 ( .A(n8883), .B(n8882), .S(n8943), .Z(n8892) );
  OR2_X1 U4900 ( .A1(n7636), .A2(n7637), .ZN(n7634) );
  AOI21_X1 U4901 ( .B1(n7437), .B2(n6499), .A(n4887), .ZN(n4886) );
  NAND2_X1 U4902 ( .A1(n7252), .A2(n7253), .ZN(n7402) );
  INV_X1 U4903 ( .A(n8721), .ZN(n4844) );
  NOR2_X1 U4904 ( .A1(n7607), .A2(n7606), .ZN(n7605) );
  AND2_X1 U4905 ( .A1(n7205), .A2(n8872), .ZN(n7207) );
  NAND2_X1 U4906 ( .A1(n5382), .A2(n5381), .ZN(n9494) );
  OR2_X1 U4907 ( .A1(n9779), .A2(n7265), .ZN(n8870) );
  NAND2_X1 U4908 ( .A1(n5254), .A2(n5253), .ZN(n5278) );
  INV_X2 U4909 ( .A(n9366), .ZN(n4322) );
  NOR2_X1 U4910 ( .A1(n6994), .A2(n6285), .ZN(n6286) );
  NOR2_X1 U4911 ( .A1(n9822), .A2(n5906), .ZN(n9821) );
  NAND2_X1 U4912 ( .A1(n4826), .A2(n4825), .ZN(n5200) );
  NAND2_X1 U4913 ( .A1(n5865), .A2(n6983), .ZN(n7962) );
  NAND2_X1 U4914 ( .A1(n5135), .A2(n5134), .ZN(n5154) );
  NAND4_X1 U4915 ( .A1(n5827), .A2(n5826), .A3(n5825), .A4(n5824), .ZN(n5842)
         );
  AND2_X1 U4916 ( .A1(n6690), .A2(n4971), .ZN(n4972) );
  NAND2_X1 U4917 ( .A1(n5003), .A2(n9136), .ZN(n7094) );
  AND2_X2 U4918 ( .A1(n7703), .A2(n7342), .ZN(n5731) );
  NAND2_X1 U4919 ( .A1(n4969), .A2(n4968), .ZN(n5019) );
  BUF_X2 U4920 ( .A(n6684), .Z(n9041) );
  NAND2_X1 U4921 ( .A1(n5085), .A2(n5084), .ZN(n5108) );
  NAND4_X1 U4922 ( .A1(n5028), .A2(n4739), .A3(n4738), .A4(n4737), .ZN(n9040)
         );
  NAND2_X1 U4923 ( .A1(n5788), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5790) );
  INV_X1 U4924 ( .A(n4971), .ZN(n5003) );
  NAND2_X1 U4925 ( .A1(n5456), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U4926 ( .A1(n4348), .A2(n4741), .ZN(n4742) );
  NAND2_X1 U4927 ( .A1(n5829), .A2(n4586), .ZN(n6054) );
  NAND2_X1 U4928 ( .A1(n6711), .A2(n5740), .ZN(n4985) );
  NAND2_X1 U4929 ( .A1(n5786), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6055) );
  NAND2_X1 U4930 ( .A1(n6223), .A2(n6224), .ZN(n7454) );
  XNOR2_X1 U4931 ( .A(n4991), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4998) );
  NAND2_X1 U4932 ( .A1(n4996), .A2(n4995), .ZN(n9572) );
  INV_X2 U4933 ( .A(n9568), .ZN(n7708) );
  OR2_X1 U4934 ( .A1(n5794), .A2(n6031), .ZN(n5776) );
  NAND2_X1 U4935 ( .A1(n4995), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4991) );
  AND2_X1 U4936 ( .A1(n5989), .A2(n5783), .ZN(n6029) );
  OAI21_X1 U4937 ( .B1(n6175), .B2(n4891), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6251) );
  XNOR2_X1 U4938 ( .A(n5082), .B(SI_3_), .ZN(n5080) );
  XNOR2_X1 U4939 ( .A(n5889), .B(n5888), .ZN(n6585) );
  NAND2_X1 U4940 ( .A1(n5861), .A2(n5860), .ZN(n6649) );
  AND2_X1 U4941 ( .A1(n5780), .A2(n5781), .ZN(n5989) );
  NOR2_X1 U4942 ( .A1(n4892), .A2(n4639), .ZN(n4638) );
  NOR2_X1 U4943 ( .A1(n4958), .A2(n4957), .ZN(n4959) );
  AND2_X1 U4944 ( .A1(n4917), .A2(n4965), .ZN(n4752) );
  NOR2_X1 U4945 ( .A1(n5766), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n4895) );
  XNOR2_X1 U4946 ( .A(n5828), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6364) );
  INV_X1 U4947 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5875) );
  INV_X1 U4948 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4950) );
  INV_X1 U4949 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10038) );
  AND2_X1 U4950 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5102) );
  INV_X1 U4951 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5207) );
  INV_X1 U4952 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5206) );
  NOR2_X1 U4953 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5764) );
  INV_X1 U4954 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4955) );
  INV_X1 U4955 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5330) );
  INV_X1 U4956 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9982) );
  INV_X1 U4957 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5453) );
  INV_X1 U4958 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5729) );
  INV_X1 U4959 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4954) );
  INV_X1 U4960 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5726) );
  INV_X1 U4961 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6225) );
  INV_X1 U4962 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5329) );
  INV_X1 U4963 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6030) );
  INV_X1 U4964 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5782) );
  INV_X1 U4965 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6221) );
  INV_X1 U4966 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5784) );
  INV_X4 U4967 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4968 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5787) );
  INV_X1 U4969 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6252) );
  INV_X1 U4970 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4928) );
  INV_X1 U4971 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5781) );
  NOR2_X1 U4972 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4930) );
  INV_X1 U4973 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4906) );
  INV_X1 U4974 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n10034) );
  INV_X1 U4975 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5999) );
  NOR2_X1 U4976 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5765) );
  XNOR2_X2 U4977 ( .A(n6684), .B(n6693), .ZN(n6685) );
  NAND3_X1 U4978 ( .A1(n4970), .A2(n7094), .A3(n5019), .ZN(n4323) );
  NAND2_X1 U4979 ( .A1(n5829), .A2(n6574), .ZN(n4325) );
  NAND2_X1 U4980 ( .A1(n5829), .A2(n4320), .ZN(n4326) );
  NAND2_X1 U4981 ( .A1(n5829), .A2(n4320), .ZN(n5849) );
  AOI21_X2 U4982 ( .B1(n6281), .B2(n6313), .A(n6282), .ZN(n6641) );
  NOR2_X2 U4983 ( .A1(n6281), .A2(n6313), .ZN(n6282) );
  OAI21_X2 U4984 ( .B1(n7739), .B2(n4901), .A(n4899), .ZN(n7762) );
  NOR2_X4 U4985 ( .A1(n9374), .A2(n9494), .ZN(n9373) );
  OR2_X2 U4986 ( .A1(n7566), .A2(n9502), .ZN(n9374) );
  NAND2_X1 U4987 ( .A1(n8863), .A2(n8862), .ZN(n4446) );
  MUX2_X1 U4988 ( .A(n8019), .B(n8018), .S(n8070), .Z(n8026) );
  INV_X1 U4989 ( .A(n7679), .ZN(n5816) );
  NAND2_X1 U4990 ( .A1(n7804), .A2(n8293), .ZN(n8055) );
  OR2_X1 U4991 ( .A1(n6255), .A2(n7779), .ZN(n7901) );
  INV_X1 U4992 ( .A(n4893), .ZN(n4891) );
  OR2_X1 U4993 ( .A1(n9394), .A2(n9197), .ZN(n8935) );
  XNOR2_X1 U4994 ( .A(n5301), .B(SI_12_), .ZN(n5300) );
  OR2_X1 U4995 ( .A1(n7836), .A2(n8113), .ZN(n6077) );
  OR2_X1 U4996 ( .A1(n9526), .A2(n9531), .ZN(n8880) );
  NAND2_X1 U4997 ( .A1(n8028), .A2(n8027), .ZN(n4496) );
  NAND2_X1 U4998 ( .A1(n4502), .A2(n4500), .ZN(n4499) );
  NOR2_X1 U4999 ( .A1(n8079), .A2(n4501), .ZN(n4500) );
  INV_X1 U5000 ( .A(n8078), .ZN(n4501) );
  AND2_X1 U5001 ( .A1(n5775), .A2(n4894), .ZN(n4893) );
  INV_X1 U5002 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4894) );
  INV_X1 U5003 ( .A(n8627), .ZN(n4848) );
  INV_X1 U5004 ( .A(n6649), .ZN(n6313) );
  NAND2_X1 U5005 ( .A1(n4516), .A2(n4518), .ZN(n4515) );
  AND2_X1 U5006 ( .A1(n4797), .A2(n4796), .ZN(n6288) );
  NAND2_X1 U5007 ( .A1(n6604), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4796) );
  NAND2_X1 U5008 ( .A1(n8528), .A2(n8293), .ZN(n4684) );
  AND2_X1 U5009 ( .A1(n7877), .A2(n8283), .ZN(n8062) );
  OR2_X1 U5010 ( .A1(n7841), .A2(n8322), .ZN(n8040) );
  OR2_X1 U5011 ( .A1(n7836), .A2(n8346), .ZN(n8030) );
  NOR2_X1 U5012 ( .A1(n5922), .A2(n4645), .ZN(n4644) );
  INV_X1 U5013 ( .A(n5905), .ZN(n4645) );
  NOR2_X1 U5014 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6309) );
  XNOR2_X1 U5015 ( .A(n5044), .B(n5705), .ZN(n5045) );
  OR2_X1 U5016 ( .A1(n9401), .A2(n9408), .ZN(n9160) );
  NAND2_X1 U5017 ( .A1(n9209), .A2(n4810), .ZN(n4809) );
  NOR2_X1 U5018 ( .A1(n9182), .A2(n4361), .ZN(n4552) );
  OAI21_X1 U5019 ( .B1(n9154), .B2(n9281), .A(n4824), .ZN(n4813) );
  NAND2_X1 U5020 ( .A1(n4824), .A2(n9154), .ZN(n4821) );
  OR2_X1 U5021 ( .A1(n9494), .A2(n9499), .ZN(n8952) );
  NOR2_X1 U5022 ( .A1(n4464), .A2(n4462), .ZN(n4461) );
  INV_X1 U5023 ( .A(n8841), .ZN(n4462) );
  AND2_X1 U5024 ( .A1(n5610), .A2(n5586), .ZN(n5611) );
  INV_X1 U5025 ( .A(n5378), .ZN(n4632) );
  AOI21_X1 U5026 ( .B1(n4596), .B2(n4598), .A(n4412), .ZN(n4594) );
  NAND2_X1 U5027 ( .A1(n4615), .A2(n4619), .ZN(n4614) );
  NAND2_X1 U5028 ( .A1(n7219), .A2(n4898), .ZN(n7667) );
  AND2_X1 U5029 ( .A1(n6458), .A2(n6930), .ZN(n6459) );
  OR2_X1 U5030 ( .A1(n4898), .A2(n4897), .ZN(n4896) );
  NAND2_X1 U5031 ( .A1(n6463), .A2(n6672), .ZN(n4881) );
  NAND2_X1 U5032 ( .A1(n7627), .A2(n7626), .ZN(n7625) );
  NAND2_X1 U5033 ( .A1(n8095), .A2(n8094), .ZN(n4505) );
  AOI21_X1 U5034 ( .B1(n8092), .B2(n6418), .A(n4338), .ZN(n4504) );
  NAND2_X1 U5035 ( .A1(n6282), .A2(n4519), .ZN(n4516) );
  XNOR2_X1 U5036 ( .A(n6288), .B(n6377), .ZN(n7319) );
  AOI21_X1 U5037 ( .B1(n4378), .B2(n8238), .A(n8237), .ZN(n8259) );
  NAND2_X1 U5038 ( .A1(n4787), .A2(n4789), .ZN(n8237) );
  OR2_X1 U5039 ( .A1(n7754), .A2(n8273), .ZN(n8063) );
  XNOR2_X1 U5040 ( .A(n7782), .B(n8077), .ZN(n7928) );
  AND2_X1 U5041 ( .A1(n4674), .A2(n4672), .ZN(n6443) );
  NOR2_X1 U5042 ( .A1(n4673), .A2(n4678), .ZN(n4672) );
  AND2_X1 U5043 ( .A1(n4679), .A2(n4687), .ZN(n4673) );
  NAND2_X1 U5044 ( .A1(n6202), .A2(n8055), .ZN(n8275) );
  NAND2_X1 U5045 ( .A1(n4721), .A2(n4334), .ZN(n6202) );
  INV_X1 U5046 ( .A(n4655), .ZN(n8333) );
  AOI21_X1 U5047 ( .B1(n4657), .B2(n4663), .A(n4667), .ZN(n4656) );
  AND2_X1 U5048 ( .A1(n8351), .A2(n8114), .ZN(n4667) );
  OAI21_X1 U5049 ( .B1(n4705), .B2(n4703), .A(n4695), .ZN(n4702) );
  INV_X1 U5050 ( .A(n4696), .ZN(n4695) );
  AND4_X1 U5051 ( .A1(n6024), .A2(n6023), .A3(n6022), .A4(n6021), .ZN(n8389)
         );
  AOI21_X1 U5052 ( .B1(n4653), .B2(n4654), .A(n4350), .ZN(n4649) );
  OR2_X1 U5053 ( .A1(n4391), .A2(n5922), .ZN(n4646) );
  NAND2_X1 U5054 ( .A1(n5905), .A2(n5904), .ZN(n4648) );
  NAND2_X1 U5055 ( .A1(n4636), .A2(n4923), .ZN(n5893) );
  INV_X1 U5056 ( .A(n5849), .ZN(n6057) );
  INV_X1 U5057 ( .A(n5829), .ZN(n6056) );
  NAND2_X1 U5058 ( .A1(n6309), .A2(n4906), .ZN(n5850) );
  AND2_X1 U5059 ( .A1(n7706), .A2(n9572), .ZN(n5050) );
  NAND2_X1 U5060 ( .A1(n4532), .A2(n4528), .ZN(n4527) );
  NAND2_X1 U5061 ( .A1(n4533), .A2(n4531), .ZN(n4528) );
  AND4_X1 U5062 ( .A1(n5750), .A2(n5749), .A3(n5748), .A4(n5747), .ZN(n9197)
         );
  NAND2_X1 U5063 ( .A1(n9282), .A2(n4823), .ZN(n4818) );
  AOI21_X1 U5064 ( .B1(n9260), .B2(n9181), .A(n4911), .ZN(n9248) );
  NAND2_X1 U5065 ( .A1(n4558), .A2(n4556), .ZN(n9355) );
  NAND2_X1 U5066 ( .A1(n4557), .A2(n4757), .ZN(n4556) );
  NAND2_X1 U5067 ( .A1(n4759), .A2(n7563), .ZN(n4557) );
  AND2_X1 U5068 ( .A1(n7487), .A2(n8891), .ZN(n4836) );
  NAND2_X1 U5069 ( .A1(n5309), .A2(n5308), .ZN(n9519) );
  NAND2_X1 U5070 ( .A1(n5282), .A2(n5281), .ZN(n9526) );
  NAND2_X1 U5071 ( .A1(n4584), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4973) );
  AND2_X1 U5072 ( .A1(n5577), .A2(n5556), .ZN(n5578) );
  INV_X1 U5073 ( .A(n5523), .ZN(n5609) );
  INV_X1 U5074 ( .A(n8107), .ZN(n8273) );
  OR2_X1 U5075 ( .A1(P2_U3150), .A2(n6409), .ZN(n8255) );
  AND4_X1 U5076 ( .A1(n5680), .A2(n5679), .A3(n5678), .A4(n5677), .ZN(n9198)
         );
  NOR2_X1 U5077 ( .A1(n7942), .A2(n7937), .ZN(n4478) );
  NAND2_X1 U5078 ( .A1(n8070), .A2(n7938), .ZN(n4479) );
  NAND2_X1 U5079 ( .A1(n7982), .A2(n4486), .ZN(n4488) );
  AND2_X1 U5080 ( .A1(n6194), .A2(n8001), .ZN(n4490) );
  OAI21_X1 U5081 ( .B1(n4621), .B2(n4622), .A(n8905), .ZN(n8906) );
  NAND2_X1 U5082 ( .A1(n4460), .A2(n8902), .ZN(n4456) );
  NAND2_X1 U5083 ( .A1(n8029), .A2(n8070), .ZN(n4497) );
  NAND2_X1 U5084 ( .A1(n4496), .A2(n8085), .ZN(n4495) );
  AND2_X1 U5085 ( .A1(n9235), .A2(n8923), .ZN(n4590) );
  AOI21_X1 U5086 ( .B1(n8918), .B2(n8917), .A(n4592), .ZN(n4591) );
  NAND2_X1 U5087 ( .A1(n8920), .A2(n8919), .ZN(n4592) );
  NAND4_X1 U5088 ( .A1(n5765), .A2(n5764), .A3(n5875), .A4(n5763), .ZN(n5766)
         );
  OR2_X1 U5089 ( .A1(n5736), .A2(n7379), .ZN(n4971) );
  INV_X1 U5090 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4931) );
  NOR2_X1 U5091 ( .A1(n4613), .A2(n5249), .ZN(n4612) );
  INV_X1 U5092 ( .A(n5248), .ZN(n5249) );
  INV_X1 U5093 ( .A(n4616), .ZN(n4613) );
  INV_X1 U5094 ( .A(n4920), .ZN(n4620) );
  INV_X1 U5095 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4608) );
  INV_X1 U5096 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4607) );
  NAND3_X1 U5097 ( .A1(n4981), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4605) );
  INV_X1 U5098 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4981) );
  INV_X1 U5099 ( .A(n6486), .ZN(n4897) );
  AND2_X1 U5100 ( .A1(n7668), .A2(n6484), .ZN(n4898) );
  AND2_X1 U5101 ( .A1(n4499), .A2(n8080), .ZN(n4498) );
  AND2_X1 U5102 ( .A1(n9813), .A2(n6312), .ZN(n6314) );
  NOR2_X1 U5103 ( .A1(n7397), .A2(n7374), .ZN(n4445) );
  NAND2_X1 U5104 ( .A1(n4736), .A2(n4735), .ZN(n4734) );
  INV_X1 U5105 ( .A(n7355), .ZN(n4735) );
  OAI21_X1 U5106 ( .B1(n6441), .B2(n4716), .A(n4714), .ZN(n7883) );
  AOI21_X1 U5107 ( .B1(n4717), .B2(n4715), .A(n4367), .ZN(n4714) );
  INV_X1 U5108 ( .A(n4717), .ZN(n4716) );
  INV_X1 U5109 ( .A(n8064), .ZN(n4715) );
  NAND2_X1 U5110 ( .A1(n6139), .A2(n6138), .ZN(n6150) );
  INV_X1 U5111 ( .A(n6140), .ZN(n6139) );
  AND2_X1 U5112 ( .A1(n4685), .A2(n4684), .ZN(n4683) );
  OR2_X1 U5113 ( .A1(n7829), .A2(n8302), .ZN(n8046) );
  NOR2_X1 U5114 ( .A1(n6098), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4436) );
  OR2_X1 U5115 ( .A1(n6071), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6082) );
  OR2_X1 U5116 ( .A1(n6061), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6063) );
  OR2_X1 U5117 ( .A1(n8395), .A2(n8374), .ZN(n8012) );
  INV_X1 U5118 ( .A(n6019), .ZN(n5811) );
  NOR2_X1 U5119 ( .A1(n5967), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n4437) );
  AOI21_X1 U5120 ( .B1(n5976), .B2(n4331), .A(n4373), .ZN(n4653) );
  INV_X1 U5121 ( .A(n7986), .ZN(n4693) );
  OR2_X1 U5122 ( .A1(n7418), .A2(n7424), .ZN(n7420) );
  NAND2_X1 U5123 ( .A1(n4720), .A2(n8422), .ZN(n6187) );
  INV_X1 U5124 ( .A(n8434), .ZN(n4720) );
  NAND2_X1 U5125 ( .A1(n7231), .A2(n8090), .ZN(n6458) );
  NAND2_X1 U5126 ( .A1(n4375), .A2(n4893), .ZN(n4892) );
  AND2_X1 U5127 ( .A1(n5599), .A2(n5598), .ZN(n5601) );
  OR2_X1 U5128 ( .A1(n9249), .A2(n4321), .ZN(n5599) );
  AOI21_X1 U5129 ( .B1(n4327), .B2(n4853), .A(n4380), .ZN(n4847) );
  NOR2_X1 U5130 ( .A1(n4872), .A2(n4871), .ZN(n4870) );
  INV_X1 U5131 ( .A(n4877), .ZN(n4871) );
  INV_X1 U5132 ( .A(n4879), .ZN(n4872) );
  NOR2_X1 U5133 ( .A1(n8745), .A2(n8746), .ZN(n4879) );
  OAI21_X1 U5134 ( .B1(n8939), .B2(n9148), .A(n4370), .ZN(n4473) );
  INV_X1 U5135 ( .A(n8941), .ZN(n8939) );
  NAND2_X1 U5136 ( .A1(n9148), .A2(n8943), .ZN(n4474) );
  NOR2_X1 U5137 ( .A1(n9229), .A2(n9411), .ZN(n4582) );
  OR2_X1 U5138 ( .A1(n9411), .A2(n9198), .ZN(n8948) );
  NAND2_X1 U5139 ( .A1(n5507), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5535) );
  NOR2_X1 U5140 ( .A1(n9487), .A2(n9350), .ZN(n4577) );
  NOR2_X1 U5141 ( .A1(n4756), .A2(n7487), .ZN(n4555) );
  OR2_X1 U5142 ( .A1(n9510), .A2(n9028), .ZN(n7563) );
  OR2_X1 U5143 ( .A1(n9510), .A2(n9516), .ZN(n8886) );
  OR2_X1 U5144 ( .A1(n9535), .A2(n8643), .ZN(n8875) );
  NOR2_X1 U5145 ( .A1(n5213), .A2(n7333), .ZN(n5233) );
  OAI21_X1 U5146 ( .B1(n7044), .B2(n9755), .A(n9038), .ZN(n6880) );
  INV_X1 U5147 ( .A(n6596), .ZN(n5724) );
  OAI21_X1 U5148 ( .B1(n7678), .B2(SI_29_), .A(n7677), .ZN(n7885) );
  NAND2_X1 U5149 ( .A1(n5690), .A2(n5689), .ZN(n6159) );
  NAND2_X1 U5150 ( .A1(n5688), .A2(n5687), .ZN(n5690) );
  NAND2_X1 U5151 ( .A1(n5666), .A2(n5665), .ZN(n5688) );
  NAND2_X1 U5152 ( .A1(n5664), .A2(n5663), .ZN(n5666) );
  NAND2_X1 U5153 ( .A1(n5640), .A2(n5639), .ZN(n5664) );
  NAND2_X1 U5154 ( .A1(n5638), .A2(n5637), .ZN(n5640) );
  AND2_X1 U5155 ( .A1(n5636), .A2(n5635), .ZN(n5637) );
  OAI21_X1 U5156 ( .B1(n5481), .B2(n5480), .A(n5479), .ZN(n5499) );
  NAND2_X1 U5157 ( .A1(n4935), .A2(n4755), .ZN(n4866) );
  AOI21_X1 U5158 ( .B1(n4631), .B2(n5375), .A(n4413), .ZN(n4629) );
  OAI21_X1 U5159 ( .B1(n5355), .B2(n5354), .A(n5353), .ZN(n5376) );
  AOI21_X1 U5160 ( .B1(n4619), .B2(n4618), .A(n4617), .ZN(n4616) );
  INV_X1 U5161 ( .A(n5228), .ZN(n4617) );
  INV_X1 U5162 ( .A(n5198), .ZN(n4618) );
  XNOR2_X1 U5163 ( .A(n5251), .B(SI_10_), .ZN(n5248) );
  AOI21_X1 U5164 ( .B1(n4828), .B2(n4830), .A(n4381), .ZN(n4825) );
  AND2_X1 U5165 ( .A1(n6476), .A2(n6472), .ZN(n4904) );
  OR2_X1 U5166 ( .A1(n5924), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U5167 ( .A1(n6481), .A2(n6480), .ZN(n7219) );
  XNOR2_X1 U5168 ( .A(n5779), .B(n5778), .ZN(n6206) );
  NAND2_X1 U5169 ( .A1(n5777), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5779) );
  OAI22_X1 U5170 ( .A1(n6060), .A2(n6308), .B1(n7027), .B2(n5835), .ZN(n4485)
         );
  NAND2_X1 U5171 ( .A1(n6617), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U5172 ( .A1(n6278), .A2(n6279), .ZN(n6654) );
  NAND2_X1 U5173 ( .A1(n6364), .A2(n4740), .ZN(n6310) );
  NAND2_X1 U5174 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n6276), .ZN(n4740) );
  NAND2_X1 U5175 ( .A1(n9805), .A2(n9806), .ZN(n9804) );
  NAND2_X1 U5176 ( .A1(n6316), .A2(n4745), .ZN(n4743) );
  NAND2_X1 U5177 ( .A1(n4355), .A2(n6641), .ZN(n4512) );
  OR2_X1 U5178 ( .A1(n4513), .A2(n4515), .ZN(n4434) );
  NOR2_X1 U5179 ( .A1(n6565), .A2(n5881), .ZN(n6564) );
  AND2_X1 U5180 ( .A1(n6990), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4769) );
  OR2_X1 U5181 ( .A1(n9823), .A2(n6287), .ZN(n4799) );
  NAND2_X1 U5182 ( .A1(n4799), .A2(n4798), .ZN(n4797) );
  INV_X1 U5183 ( .A(n7392), .ZN(n4798) );
  OR2_X1 U5184 ( .A1(n5918), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5934) );
  OR2_X1 U5185 ( .A1(n7319), .A2(n4416), .ZN(n4522) );
  NAND2_X1 U5186 ( .A1(n6289), .A2(n4523), .ZN(n4521) );
  NOR2_X1 U5187 ( .A1(n7319), .A2(n5939), .ZN(n7318) );
  OR2_X1 U5188 ( .A1(n8138), .A2(n6296), .ZN(n6298) );
  OR2_X1 U5189 ( .A1(n8177), .A2(n6351), .ZN(n4783) );
  NAND2_X1 U5190 ( .A1(n6329), .A2(n4782), .ZN(n4781) );
  INV_X1 U5191 ( .A(n8177), .ZN(n4782) );
  OR2_X1 U5192 ( .A1(n8155), .A2(n6351), .ZN(n4785) );
  AOI21_X1 U5193 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n6824), .A(n8167), .ZN(
        n6301) );
  OR2_X1 U5194 ( .A1(n8185), .A2(n8498), .ZN(n4795) );
  AND3_X1 U5195 ( .A1(n4793), .A2(n4424), .A3(n4792), .ZN(n6302) );
  NAND2_X1 U5196 ( .A1(n6163), .A2(n6162), .ZN(n6255) );
  XNOR2_X1 U5197 ( .A(n7883), .B(n8079), .ZN(n6217) );
  NOR2_X1 U5198 ( .A1(n8077), .A2(n8392), .ZN(n6445) );
  INV_X1 U5199 ( .A(n4683), .ZN(n4681) );
  AOI22_X1 U5200 ( .A1(n4683), .A2(n6115), .B1(n4682), .B2(n4684), .ZN(n4680)
         );
  OR2_X1 U5201 ( .A1(n8061), .A2(n8062), .ZN(n8274) );
  AOI21_X1 U5202 ( .B1(n8041), .B2(n4724), .A(n4723), .ZN(n4722) );
  INV_X1 U5203 ( .A(n8046), .ZN(n4723) );
  NAND2_X1 U5204 ( .A1(n8532), .A2(n8302), .ZN(n4685) );
  AND2_X1 U5205 ( .A1(n6134), .A2(n6133), .ZN(n8283) );
  AND2_X1 U5206 ( .A1(n8049), .A2(n8046), .ZN(n8296) );
  AND2_X1 U5207 ( .A1(n6126), .A2(n6125), .ZN(n8293) );
  INV_X1 U5208 ( .A(n4662), .ZN(n4661) );
  OAI21_X1 U5209 ( .B1(n4663), .B2(n8371), .A(n4668), .ZN(n4662) );
  NAND2_X1 U5210 ( .A1(n8556), .A2(n8375), .ZN(n4668) );
  NAND2_X1 U5211 ( .A1(n8372), .A2(n4664), .ZN(n4660) );
  AND2_X1 U5212 ( .A1(n4660), .A2(n4657), .ZN(n8344) );
  AND2_X1 U5213 ( .A1(n8023), .A2(n8027), .ZN(n8349) );
  AND4_X1 U5214 ( .A1(n5821), .A2(n5820), .A3(n5819), .A4(n5818), .ZN(n8360)
         );
  NAND2_X1 U5215 ( .A1(n4666), .A2(n8371), .ZN(n4665) );
  INV_X1 U5216 ( .A(n8372), .ZN(n4666) );
  OR2_X1 U5217 ( .A1(n6037), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6048) );
  INV_X1 U5218 ( .A(n4728), .ZN(n4727) );
  OAI21_X1 U5219 ( .B1(n4347), .B2(n4729), .A(n8008), .ZN(n4728) );
  OR2_X1 U5220 ( .A1(n6196), .A2(n4730), .ZN(n4729) );
  AND2_X1 U5221 ( .A1(n8008), .A2(n8006), .ZN(n8002) );
  OR2_X1 U5222 ( .A1(n6007), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U5223 ( .A1(n6192), .A2(n4347), .ZN(n8417) );
  NAND2_X1 U5224 ( .A1(n4437), .A2(n7527), .ZN(n5993) );
  AND2_X1 U5225 ( .A1(n7420), .A2(n7974), .ZN(n6191) );
  AND4_X1 U5226 ( .A1(n5972), .A2(n5971), .A3(n5970), .A4(n5969), .ZN(n7578)
         );
  NAND2_X1 U5227 ( .A1(n7233), .A2(n4644), .ZN(n4641) );
  AOI21_X1 U5228 ( .B1(n7233), .B2(n4357), .A(n4642), .ZN(n7370) );
  NOR2_X1 U5229 ( .A1(n4646), .A2(n4643), .ZN(n4642) );
  INV_X1 U5230 ( .A(n7912), .ZN(n4643) );
  OR2_X1 U5231 ( .A1(n8432), .A2(n9876), .ZN(n8422) );
  OR2_X1 U5232 ( .A1(n5894), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U5233 ( .A1(n6895), .A2(n5801), .ZN(n5882) );
  INV_X1 U5234 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U5235 ( .A1(n8125), .A2(n4635), .ZN(n4634) );
  NAND2_X1 U5236 ( .A1(n6977), .A2(n5868), .ZN(n7109) );
  INV_X1 U5237 ( .A(n8430), .ZN(n8392) );
  INV_X1 U5238 ( .A(n8433), .ZN(n8390) );
  AND2_X1 U5239 ( .A1(n6534), .A2(n8085), .ZN(n8433) );
  NAND2_X1 U5240 ( .A1(n7901), .A2(n7882), .ZN(n8079) );
  AOI22_X1 U5241 ( .A1(n6443), .A2(n6147), .B1(n8273), .B2(n8266), .ZN(n6262)
         );
  NAND2_X1 U5242 ( .A1(n6005), .A2(n6004), .ZN(n8500) );
  NAND2_X1 U5243 ( .A1(n6220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6222) );
  NOR2_X1 U5244 ( .A1(n6178), .A2(n6172), .ZN(n7933) );
  INV_X1 U5245 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5915) );
  AND2_X1 U5246 ( .A1(n5712), .A2(n4967), .ZN(n4968) );
  INV_X1 U5247 ( .A(n7482), .ZN(n4969) );
  AND2_X1 U5248 ( .A1(n8681), .A2(n5575), .ZN(n8597) );
  NAND2_X1 U5249 ( .A1(n5197), .A2(n5196), .ZN(n4862) );
  AND2_X1 U5250 ( .A1(n4876), .A2(n4874), .ZN(n4873) );
  INV_X1 U5251 ( .A(n8649), .ZN(n4874) );
  NAND2_X1 U5252 ( .A1(n8680), .A2(n5605), .ZN(n4876) );
  NAND2_X1 U5253 ( .A1(n5195), .A2(n5194), .ZN(n4863) );
  AND2_X1 U5254 ( .A1(n5233), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U5255 ( .A1(n5263), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U5256 ( .A1(n5122), .A2(n4857), .ZN(n4856) );
  INV_X1 U5257 ( .A(n5100), .ZN(n4857) );
  INV_X1 U5258 ( .A(n6860), .ZN(n5095) );
  AND4_X1 U5259 ( .A1(n5152), .A2(n5151), .A3(n5150), .A4(n5149), .ZN(n8848)
         );
  NAND4_X1 U5260 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n4999), .ZN(n6684)
         );
  NAND2_X1 U5261 ( .A1(n5050), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5001) );
  NAND2_X1 U5262 ( .A1(n8769), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5000) );
  NOR2_X1 U5263 ( .A1(n9604), .A2(n4560), .ZN(n9097) );
  AND2_X1 U5264 ( .A1(n9609), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4560) );
  XNOR2_X1 U5265 ( .A(n9229), .B(n9242), .ZN(n9221) );
  INV_X1 U5266 ( .A(n4552), .ZN(n4551) );
  AOI21_X1 U5267 ( .B1(n4552), .B2(n4550), .A(n4376), .ZN(n4549) );
  INV_X1 U5268 ( .A(n9183), .ZN(n4550) );
  AND2_X1 U5269 ( .A1(n8833), .A2(n9157), .ZN(n9235) );
  INV_X1 U5270 ( .A(n4819), .ZN(n4814) );
  OAI22_X1 U5271 ( .A1(n9275), .A2(n9179), .B1(n9299), .B2(n9446), .ZN(n9260)
         );
  NOR2_X1 U5272 ( .A1(n9280), .A2(n9439), .ZN(n9179) );
  AND2_X1 U5273 ( .A1(n8915), .A2(n9153), .ZN(n9281) );
  NAND2_X1 U5274 ( .A1(n4837), .A2(n9307), .ZN(n9297) );
  NAND2_X1 U5275 ( .A1(n4353), .A2(n4909), .ZN(n4543) );
  OR2_X1 U5276 ( .A1(n9460), .A2(n9466), .ZN(n4910) );
  OR2_X1 U5277 ( .A1(n4623), .A2(n9177), .ZN(n4909) );
  NAND2_X1 U5278 ( .A1(n8907), .A2(n9151), .ZN(n9305) );
  AOI21_X1 U5279 ( .B1(n9334), .B2(n9176), .A(n4908), .ZN(n9321) );
  NAND2_X1 U5280 ( .A1(n9350), .A2(n9465), .ZN(n9176) );
  INV_X1 U5281 ( .A(n9172), .ZN(n4760) );
  NAND2_X1 U5282 ( .A1(n9170), .A2(n9507), .ZN(n9172) );
  AND2_X1 U5283 ( .A1(n8952), .A2(n8986), .ZN(n9372) );
  NAND2_X1 U5284 ( .A1(n7490), .A2(n8884), .ZN(n7564) );
  AND2_X1 U5285 ( .A1(n7407), .A2(n4750), .ZN(n4749) );
  NAND2_X1 U5286 ( .A1(n7253), .A2(n7405), .ZN(n4750) );
  INV_X1 U5287 ( .A(n7405), .ZN(n4751) );
  NAND2_X1 U5288 ( .A1(n7402), .A2(n7401), .ZN(n7485) );
  NAND2_X1 U5289 ( .A1(n7242), .A2(n7241), .ZN(n7243) );
  OR2_X1 U5290 ( .A1(n9535), .A2(n9031), .ZN(n7241) );
  NAND2_X1 U5291 ( .A1(n7243), .A2(n8971), .ZN(n7406) );
  NAND2_X1 U5292 ( .A1(n7210), .A2(n7209), .ZN(n7211) );
  OR2_X1 U5293 ( .A1(n7208), .A2(n9032), .ZN(n7209) );
  NAND2_X1 U5294 ( .A1(n7211), .A2(n8970), .ZN(n7242) );
  INV_X1 U5295 ( .A(n8794), .ZN(n5457) );
  OR2_X1 U5296 ( .A1(n9779), .A2(n9033), .ZN(n7147) );
  NAND3_X1 U5297 ( .A1(n6880), .A2(n6879), .A3(n8843), .ZN(n4463) );
  NAND2_X1 U5298 ( .A1(n6880), .A2(n6879), .ZN(n7013) );
  AND4_X1 U5299 ( .A1(n5106), .A2(n5105), .A3(n5104), .A4(n5103), .ZN(n7046)
         );
  AND2_X1 U5300 ( .A1(n9010), .A2(n7379), .ZN(n6688) );
  INV_X1 U5301 ( .A(n9148), .ZN(n9391) );
  INV_X1 U5302 ( .A(n9393), .ZN(n9396) );
  NAND2_X1 U5303 ( .A1(n9394), .A2(n9762), .ZN(n9395) );
  NAND2_X1 U5304 ( .A1(n9401), .A2(n9762), .ZN(n4834) );
  INV_X1 U5305 ( .A(n9249), .ZN(n9433) );
  INV_X1 U5306 ( .A(n9280), .ZN(n9446) );
  AND2_X1 U5307 ( .A1(n9002), .A2(n5740), .ZN(n9475) );
  INV_X1 U5308 ( .A(n9170), .ZN(n9502) );
  INV_X1 U5309 ( .A(n9523), .ZN(n9481) );
  XNOR2_X1 U5310 ( .A(n7885), .B(n7884), .ZN(n8773) );
  NOR2_X1 U5311 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4468), .ZN(n4466) );
  XNOR2_X1 U5312 ( .A(n6159), .B(n6158), .ZN(n7585) );
  XNOR2_X1 U5313 ( .A(n5664), .B(n5663), .ZN(n7500) );
  XNOR2_X1 U5314 ( .A(n5619), .B(n5636), .ZN(n7476) );
  AND2_X1 U5315 ( .A1(n5638), .A2(n5635), .ZN(n5619) );
  XNOR2_X1 U5316 ( .A(n5587), .B(n5611), .ZN(n7452) );
  AND2_X1 U5317 ( .A1(n5582), .A2(n5612), .ZN(n5587) );
  OR2_X1 U5318 ( .A1(n5551), .A2(n5550), .ZN(n5579) );
  AND2_X1 U5319 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  XNOR2_X1 U5320 ( .A(n5532), .B(n5547), .ZN(n7478) );
  NAND2_X1 U5321 ( .A1(n5527), .A2(n5549), .ZN(n5532) );
  INV_X1 U5322 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U5323 ( .A1(n4595), .A2(n4597), .ZN(n5326) );
  NAND2_X1 U5324 ( .A1(n5278), .A2(n4600), .ZN(n4595) );
  NAND2_X1 U5325 ( .A1(n4602), .A2(n5276), .ZN(n5305) );
  NAND2_X1 U5326 ( .A1(n4604), .A2(n4603), .ZN(n4602) );
  INV_X1 U5327 ( .A(n5278), .ZN(n4604) );
  XNOR2_X1 U5328 ( .A(n5173), .B(SI_7_), .ZN(n5172) );
  XNOR2_X1 U5329 ( .A(n5155), .B(SI_6_), .ZN(n5153) );
  INV_X1 U5330 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4864) );
  NOR2_X2 U5331 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4987) );
  AND3_X1 U5332 ( .A1(n6095), .A2(n6094), .A3(n6093), .ZN(n8322) );
  NAND2_X1 U5333 ( .A1(n6097), .A2(n6096), .ZN(n7767) );
  AND4_X1 U5334 ( .A1(n6076), .A2(n6075), .A3(n6074), .A4(n6073), .ZN(n8346)
         );
  NAND2_X1 U5335 ( .A1(n7739), .A2(n7786), .ZN(n7789) );
  NAND2_X1 U5336 ( .A1(n4885), .A2(n6499), .ZN(n7525) );
  NAND2_X1 U5337 ( .A1(n7436), .A2(n6498), .ZN(n4885) );
  INV_X1 U5338 ( .A(n8111), .ZN(n8312) );
  AOI21_X1 U5339 ( .B1(n4886), .B2(n4888), .A(n4884), .ZN(n4883) );
  INV_X1 U5340 ( .A(n7524), .ZN(n4884) );
  INV_X1 U5341 ( .A(n8121), .ZN(n7549) );
  INV_X1 U5342 ( .A(n8524), .ZN(n7877) );
  NAND4_X1 U5343 ( .A1(n5914), .A2(n5913), .A3(n5912), .A4(n5911), .ZN(n8123)
         );
  OR2_X1 U5344 ( .A1(n7027), .A2(n5822), .ZN(n5827) );
  OAI21_X1 U5345 ( .B1(n6588), .B2(n6307), .A(n6306), .ZN(n9815) );
  OR2_X1 U5346 ( .A1(n8185), .A2(n4794), .ZN(n4792) );
  OR2_X1 U5347 ( .A1(n8203), .A2(n8498), .ZN(n4794) );
  OR2_X1 U5348 ( .A1(n4330), .A2(n8203), .ZN(n4793) );
  NAND2_X1 U5349 ( .A1(n4763), .A2(n4762), .ZN(n8211) );
  INV_X1 U5350 ( .A(n8256), .ZN(n4442) );
  OR2_X1 U5351 ( .A1(n8259), .A2(n9825), .ZN(n4443) );
  INV_X1 U5352 ( .A(n8247), .ZN(n8250) );
  XNOR2_X1 U5353 ( .A(n4525), .B(n6305), .ZN(n4524) );
  NOR2_X1 U5354 ( .A1(n8241), .A2(n8240), .ZN(n8239) );
  NOR2_X1 U5355 ( .A1(n9832), .A2(n4773), .ZN(n4771) );
  NOR2_X1 U5356 ( .A1(n4774), .A2(n4779), .ZN(n4773) );
  INV_X1 U5357 ( .A(n4776), .ZN(n4774) );
  INV_X1 U5358 ( .A(n8518), .ZN(n7896) );
  INV_X1 U5359 ( .A(n6255), .ZN(n7724) );
  NAND2_X1 U5360 ( .A1(n4719), .A2(n8063), .ZN(n6265) );
  INV_X1 U5361 ( .A(n8076), .ZN(n7782) );
  NAND2_X1 U5362 ( .A1(n6047), .A2(n6046), .ZN(n8383) );
  INV_X1 U5363 ( .A(n8398), .ZN(n8418) );
  OR2_X1 U5364 ( .A1(n6834), .A2(n8413), .ZN(n8429) );
  NAND2_X1 U5365 ( .A1(n7895), .A2(n7894), .ZN(n8513) );
  AND2_X1 U5366 ( .A1(n4713), .A2(n6219), .ZN(n4711) );
  NAND2_X1 U5367 ( .A1(n6218), .A2(n9901), .ZN(n6219) );
  AND2_X1 U5368 ( .A1(n6235), .A2(n6234), .ZN(n8574) );
  OAI22_X1 U5369 ( .A1(n6575), .A2(n4586), .B1(n4611), .B2(n6574), .ZN(n4585)
         );
  INV_X1 U5370 ( .A(n9295), .ZN(n9451) );
  INV_X1 U5371 ( .A(n9458), .ZN(n9283) );
  NAND2_X1 U5372 ( .A1(n5050), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n4737) );
  NAND2_X1 U5373 ( .A1(n4317), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4738) );
  NOR2_X1 U5374 ( .A1(n9592), .A2(n4561), .ZN(n9606) );
  AND2_X1 U5375 ( .A1(n9597), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4561) );
  OAI21_X1 U5376 ( .B1(n9168), .B2(n9523), .A(n9167), .ZN(n9398) );
  AOI21_X1 U5377 ( .B1(n9166), .B2(n9474), .A(n9165), .ZN(n9167) );
  OAI21_X1 U5378 ( .B1(n9185), .B2(n4532), .A(n4527), .ZN(n4526) );
  NAND2_X1 U5379 ( .A1(n4545), .A2(n4358), .ZN(n4529) );
  OR2_X1 U5380 ( .A1(n4545), .A2(n4399), .ZN(n4530) );
  NAND2_X1 U5381 ( .A1(n4328), .A2(n9195), .ZN(n4807) );
  OAI21_X1 U5382 ( .B1(n4328), .B2(n4806), .A(n4804), .ZN(n4803) );
  NAND2_X1 U5383 ( .A1(n4746), .A2(n9193), .ZN(n9406) );
  NAND2_X1 U5384 ( .A1(n4535), .A2(n4534), .ZN(n9193) );
  NAND2_X1 U5385 ( .A1(n4341), .A2(n9195), .ZN(n4746) );
  NAND2_X1 U5386 ( .A1(n5559), .A2(n5558), .ZN(n9441) );
  OAI21_X1 U5387 ( .B1(n4480), .B2(n4477), .A(n4476), .ZN(n7963) );
  NOR2_X1 U5388 ( .A1(n4479), .A2(n4478), .ZN(n4477) );
  OR2_X1 U5389 ( .A1(n7949), .A2(n7948), .ZN(n4476) );
  AOI22_X1 U5390 ( .A1(n4487), .A2(n4489), .B1(n4490), .B2(n4491), .ZN(n8003)
         );
  NAND2_X1 U5391 ( .A1(n7998), .A2(n7997), .ZN(n4491) );
  AND3_X1 U5392 ( .A1(n4392), .A2(n4488), .A3(n4490), .ZN(n4487) );
  NAND2_X1 U5393 ( .A1(n7487), .A2(n8893), .ZN(n4454) );
  NAND2_X1 U5394 ( .A1(n4459), .A2(n4458), .ZN(n4457) );
  NOR2_X1 U5395 ( .A1(n8903), .A2(n8943), .ZN(n4458) );
  NAND2_X1 U5396 ( .A1(n4460), .A2(n8904), .ZN(n4459) );
  NAND2_X1 U5397 ( .A1(n4493), .A2(n4492), .ZN(n8043) );
  AND2_X1 U5398 ( .A1(n8313), .A2(n8036), .ZN(n4492) );
  NAND2_X1 U5399 ( .A1(n4494), .A2(n8033), .ZN(n4493) );
  NAND2_X1 U5400 ( .A1(n8922), .A2(n4590), .ZN(n4589) );
  MUX2_X1 U5401 ( .A(n8072), .B(n8071), .S(n8085), .Z(n8073) );
  NAND2_X1 U5402 ( .A1(n7896), .A2(n8105), .ZN(n7902) );
  AND2_X1 U5403 ( .A1(n8222), .A2(n6396), .ZN(n6399) );
  NOR2_X1 U5404 ( .A1(n7928), .A2(n4718), .ZN(n4717) );
  INV_X1 U5405 ( .A(n8063), .ZN(n4718) );
  AND2_X1 U5406 ( .A1(n7829), .A2(n8302), .ZN(n8045) );
  INV_X1 U5407 ( .A(n7342), .ZN(n5736) );
  NAND2_X1 U5408 ( .A1(n6161), .A2(n6160), .ZN(n7676) );
  NAND2_X1 U5409 ( .A1(n6159), .A2(n6158), .ZN(n6161) );
  INV_X1 U5410 ( .A(n5402), .ZN(n5404) );
  INV_X1 U5411 ( .A(n5374), .ZN(n5377) );
  AOI21_X1 U5412 ( .B1(n4597), .B2(n4599), .A(n5325), .ZN(n4596) );
  NAND2_X1 U5413 ( .A1(n5203), .A2(n5202), .ZN(n5228) );
  INV_X1 U5414 ( .A(n5157), .ZN(n4830) );
  INV_X1 U5415 ( .A(n4829), .ZN(n4828) );
  OAI21_X1 U5416 ( .B1(n5153), .B2(n4830), .A(n5172), .ZN(n4829) );
  NAND3_X1 U5417 ( .A1(n4742), .A2(n4383), .A3(n4743), .ZN(n6317) );
  OR2_X1 U5418 ( .A1(n7315), .A2(n6322), .ZN(n4736) );
  AND2_X1 U5419 ( .A1(n4734), .A2(n4733), .ZN(n6325) );
  NAND2_X1 U5420 ( .A1(n7361), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4733) );
  AOI21_X1 U5421 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8146), .A(n8137), .ZN(
        n6328) );
  AND3_X1 U5422 ( .A1(n4780), .A2(n4781), .A3(n4422), .ZN(n6331) );
  AND3_X1 U5423 ( .A1(n4763), .A2(n4425), .A3(n4762), .ZN(n6335) );
  OR2_X1 U5424 ( .A1(n6150), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7720) );
  NOR2_X1 U5425 ( .A1(n4681), .A2(n4332), .ZN(n4679) );
  NAND2_X1 U5426 ( .A1(n4679), .A2(n4676), .ZN(n4675) );
  INV_X1 U5427 ( .A(n6105), .ZN(n4676) );
  OAI21_X1 U5428 ( .B1(n4680), .B2(n4332), .A(n4382), .ZN(n4678) );
  OR2_X1 U5429 ( .A1(n7877), .A2(n8283), .ZN(n7903) );
  OR2_X1 U5430 ( .A1(n7738), .A2(n8336), .ZN(n8034) );
  INV_X1 U5431 ( .A(n6082), .ZN(n6081) );
  INV_X1 U5432 ( .A(n8349), .ZN(n4659) );
  NAND2_X1 U5433 ( .A1(n8027), .A2(n6199), .ZN(n4697) );
  OR2_X1 U5434 ( .A1(n4703), .A2(n4707), .ZN(n4698) );
  INV_X1 U5435 ( .A(n6063), .ZN(n5813) );
  INV_X1 U5436 ( .A(n6195), .ZN(n4730) );
  NAND2_X1 U5437 ( .A1(n4331), .A2(n5977), .ZN(n4654) );
  INV_X1 U5438 ( .A(n4437), .ZN(n5982) );
  OR2_X1 U5439 ( .A1(n8123), .A2(n9882), .ZN(n7975) );
  OR2_X1 U5440 ( .A1(n8125), .A2(n9867), .ZN(n7952) );
  NAND2_X1 U5441 ( .A1(n5834), .A2(n9850), .ZN(n6942) );
  CLKBUF_X1 U5442 ( .A(n6457), .Z(n6417) );
  AND2_X1 U5443 ( .A1(n7931), .A2(n6193), .ZN(n8407) );
  NAND2_X1 U5444 ( .A1(n4647), .A2(n5905), .ZN(n8435) );
  OR2_X1 U5445 ( .A1(n7233), .A2(n5904), .ZN(n4647) );
  OR2_X1 U5446 ( .A1(n6233), .A2(n6248), .ZN(n6537) );
  NAND2_X1 U5447 ( .A1(n4640), .A2(n5773), .ZN(n4639) );
  INV_X1 U5448 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4640) );
  INV_X1 U5449 ( .A(n5766), .ZN(n5767) );
  NAND2_X1 U5450 ( .A1(n4323), .A2(n5658), .ZN(n5043) );
  NOR2_X1 U5451 ( .A1(n5606), .A2(n4878), .ZN(n4877) );
  INV_X1 U5452 ( .A(n8681), .ZN(n4878) );
  NAND2_X1 U5453 ( .A1(n8934), .A2(n9185), .ZN(n4475) );
  NOR2_X1 U5454 ( .A1(n9001), .A2(n8998), .ZN(n4472) );
  INV_X1 U5455 ( .A(n4534), .ZN(n4533) );
  NAND2_X1 U5456 ( .A1(n4821), .A2(n4820), .ZN(n4819) );
  NOR2_X1 U5457 ( .A1(n9251), .A2(n4822), .ZN(n4820) );
  INV_X1 U5458 ( .A(n4922), .ZN(n4758) );
  NOR2_X1 U5459 ( .A1(n4579), .A2(n9519), .ZN(n4578) );
  INV_X1 U5460 ( .A(n4580), .ZN(n4579) );
  NOR2_X1 U5461 ( .A1(n9526), .A2(n9535), .ZN(n4580) );
  INV_X1 U5462 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5184) );
  NOR2_X1 U5463 ( .A1(n9433), .A2(n9266), .ZN(n9254) );
  NAND2_X1 U5464 ( .A1(n9265), .A2(n9138), .ZN(n9266) );
  NOR2_X1 U5465 ( .A1(n7039), .A2(n7699), .ZN(n7038) );
  XNOR2_X1 U5466 ( .A(n7676), .B(n7675), .ZN(n7678) );
  AND2_X1 U5467 ( .A1(n5689), .A2(n5670), .ZN(n5687) );
  AND2_X1 U5468 ( .A1(n5665), .A2(n5644), .ZN(n5663) );
  OR2_X1 U5469 ( .A1(n5614), .A2(n5613), .ZN(n5635) );
  AND2_X1 U5470 ( .A1(n5612), .A2(n5611), .ZN(n5613) );
  NAND2_X1 U5471 ( .A1(n5609), .A2(n5608), .ZN(n5638) );
  AND2_X1 U5472 ( .A1(n5607), .A2(n5610), .ZN(n5608) );
  NAND2_X1 U5473 ( .A1(n4953), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5727) );
  INV_X1 U5474 ( .A(n5276), .ZN(n4601) );
  INV_X1 U5475 ( .A(n5300), .ZN(n5304) );
  INV_X1 U5476 ( .A(n5277), .ZN(n4603) );
  NAND2_X1 U5477 ( .A1(n5252), .A2(SI_10_), .ZN(n5253) );
  NAND2_X1 U5478 ( .A1(n4614), .A2(n4612), .ZN(n5254) );
  NAND2_X1 U5479 ( .A1(n5177), .A2(n5176), .ZN(n5198) );
  OAI21_X1 U5480 ( .B1(n4982), .B2(n4611), .A(n4610), .ZN(n5036) );
  XNOR2_X1 U5481 ( .A(n5036), .B(SI_1_), .ZN(n5033) );
  NOR2_X1 U5482 ( .A1(n7817), .A2(n4890), .ZN(n4889) );
  INV_X1 U5483 ( .A(n6513), .ZN(n4890) );
  AOI21_X1 U5484 ( .B1(n4902), .B2(n4900), .A(n4339), .ZN(n4899) );
  INV_X1 U5485 ( .A(n4902), .ZN(n4901) );
  NAND2_X1 U5486 ( .A1(n7667), .A2(n6486), .ZN(n7544) );
  INV_X1 U5487 ( .A(n6528), .ZN(n4438) );
  INV_X1 U5488 ( .A(n6499), .ZN(n4888) );
  NOR2_X1 U5489 ( .A1(n7842), .A2(n4903), .ZN(n4902) );
  INV_X1 U5490 ( .A(n7742), .ZN(n4903) );
  INV_X1 U5491 ( .A(n7774), .ZN(n7749) );
  NAND2_X1 U5492 ( .A1(n6515), .A2(n8391), .ZN(n7851) );
  AND2_X1 U5493 ( .A1(n6828), .A2(n6537), .ZN(n6548) );
  NAND2_X1 U5494 ( .A1(n4520), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6652) );
  INV_X1 U5495 ( .A(n6654), .ZN(n4520) );
  NAND2_X1 U5496 ( .A1(n6641), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6844) );
  INV_X1 U5497 ( .A(n6315), .ZN(n4744) );
  XNOR2_X1 U5498 ( .A(n6317), .B(n6585), .ZN(n6562) );
  NOR2_X1 U5499 ( .A1(n6562), .A2(n7161), .ZN(n6561) );
  AOI21_X1 U5500 ( .B1(n6585), .B2(n6317), .A(n6561), .ZN(n6993) );
  INV_X1 U5501 ( .A(n4515), .ZN(n4510) );
  XNOR2_X1 U5502 ( .A(n6286), .B(n9829), .ZN(n9824) );
  INV_X1 U5503 ( .A(n4734), .ZN(n7354) );
  INV_X1 U5504 ( .A(n4736), .ZN(n7356) );
  NOR2_X1 U5505 ( .A1(n6382), .A2(n7348), .ZN(n7615) );
  NOR2_X1 U5506 ( .A1(n7605), .A2(n6293), .ZN(n8140) );
  NOR2_X1 U5507 ( .A1(n7615), .A2(n7616), .ZN(n7614) );
  OR2_X1 U5508 ( .A1(n8192), .A2(n4765), .ZN(n4762) );
  OR2_X1 U5509 ( .A1(n8212), .A2(n8191), .ZN(n4765) );
  NAND2_X1 U5510 ( .A1(n6332), .A2(n4764), .ZN(n4763) );
  INV_X1 U5511 ( .A(n8212), .ZN(n4764) );
  OR2_X1 U5512 ( .A1(n8192), .A2(n8191), .ZN(n4767) );
  INV_X1 U5513 ( .A(n8220), .ZN(n4435) );
  OR2_X1 U5514 ( .A1(n8220), .A2(n4423), .ZN(n4789) );
  NAND2_X1 U5515 ( .A1(n6303), .A2(n4788), .ZN(n4787) );
  INV_X1 U5516 ( .A(n8238), .ZN(n4788) );
  NAND2_X1 U5517 ( .A1(n4779), .A2(n6338), .ZN(n4776) );
  INV_X1 U5518 ( .A(n6404), .ZN(n4779) );
  NAND2_X1 U5519 ( .A1(n6150), .A2(n6141), .ZN(n8264) );
  INV_X1 U5520 ( .A(n6120), .ZN(n6119) );
  INV_X1 U5521 ( .A(n4436), .ZN(n6108) );
  NAND2_X1 U5522 ( .A1(n4436), .A2(n7825), .ZN(n6120) );
  OR2_X1 U5523 ( .A1(n8041), .A2(n8044), .ZN(n8303) );
  AND2_X1 U5524 ( .A1(n8040), .A2(n8037), .ZN(n8313) );
  NAND2_X1 U5525 ( .A1(n8371), .A2(n8021), .ZN(n4700) );
  INV_X1 U5526 ( .A(n6048), .ZN(n5812) );
  OR2_X1 U5527 ( .A1(n6014), .A2(n6013), .ZN(n7656) );
  AND4_X1 U5528 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n8374)
         );
  INV_X1 U5529 ( .A(n8407), .ZN(n6194) );
  INV_X1 U5530 ( .A(n5993), .ZN(n5809) );
  INV_X1 U5531 ( .A(n8119), .ZN(n7994) );
  NAND2_X1 U5532 ( .A1(n4651), .A2(n4653), .ZN(n8404) );
  OR2_X1 U5533 ( .A1(n7461), .A2(n4654), .ZN(n4651) );
  AOI21_X1 U5534 ( .B1(n7916), .B2(n4693), .A(n4692), .ZN(n4691) );
  INV_X1 U5535 ( .A(n7989), .ZN(n4692) );
  INV_X1 U5536 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5806) );
  INV_X1 U5537 ( .A(n5940), .ZN(n5807) );
  OR2_X1 U5538 ( .A1(n5956), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5967) );
  AND2_X1 U5539 ( .A1(n7985), .A2(n7986), .ZN(n7915) );
  NAND2_X1 U5540 ( .A1(n6190), .A2(n4365), .ZN(n7418) );
  INV_X1 U5541 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5804) );
  INV_X1 U5542 ( .A(n5908), .ZN(n5805) );
  NAND2_X1 U5543 ( .A1(n7975), .A2(n7368), .ZN(n8434) );
  INV_X1 U5544 ( .A(n6187), .ZN(n7367) );
  INV_X1 U5545 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5802) );
  INV_X1 U5546 ( .A(n5882), .ZN(n5803) );
  OR2_X1 U5547 ( .A1(n6833), .A2(n6204), .ZN(n8440) );
  NAND2_X1 U5548 ( .A1(n6137), .A2(n6136), .ZN(n7754) );
  NAND2_X1 U5549 ( .A1(n6090), .A2(n6089), .ZN(n7841) );
  NAND2_X1 U5550 ( .A1(n6070), .A2(n6069), .ZN(n7836) );
  NAND2_X1 U5551 ( .A1(n6018), .A2(n6017), .ZN(n7645) );
  AND2_X1 U5552 ( .A1(n4652), .A2(n5975), .ZN(n7638) );
  OR2_X1 U5553 ( .A1(n7461), .A2(n5973), .ZN(n4652) );
  AND3_X1 U5554 ( .A1(n5864), .A2(n5863), .A3(n5862), .ZN(n9860) );
  AND2_X1 U5555 ( .A1(n6548), .A2(n8573), .ZN(n6533) );
  XNOR2_X1 U5556 ( .A(P2_IR_REG_1__SCAN_IN), .B(keyinput6), .ZN(n10020) );
  NOR2_X1 U5557 ( .A1(n4892), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n4637) );
  AND3_X2 U5558 ( .A1(n4895), .A2(n5768), .A3(n5772), .ZN(n5774) );
  NOR2_X1 U5559 ( .A1(n5771), .A2(n5770), .ZN(n5772) );
  NAND2_X1 U5560 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5828) );
  AOI22_X1 U5561 ( .A1(n9041), .A2(n5654), .B1(n6692), .B2(n5697), .ZN(n5007)
         );
  AOI21_X1 U5562 ( .B1(n4854), .B2(n4852), .A(n4379), .ZN(n4851) );
  INV_X1 U5563 ( .A(n5474), .ZN(n4852) );
  AND2_X1 U5564 ( .A1(n5462), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5484) );
  OR2_X1 U5565 ( .A1(n5311), .A2(n5310), .ZN(n5338) );
  AND2_X1 U5566 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n5536), .ZN(n5560) );
  AND2_X1 U5567 ( .A1(n8720), .A2(n8605), .ZN(n4843) );
  INV_X1 U5568 ( .A(n5046), .ZN(n7694) );
  AND2_X1 U5569 ( .A1(n5460), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5462) );
  CLKBUF_X1 U5570 ( .A(n8614), .Z(n8616) );
  INV_X1 U5571 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U5572 ( .A1(n4867), .A2(n4868), .ZN(n8744) );
  NAND2_X1 U5573 ( .A1(n4869), .A2(n4879), .ZN(n4868) );
  INV_X1 U5574 ( .A(n4873), .ZN(n4869) );
  NOR2_X1 U5575 ( .A1(n5338), .A2(n5337), .ZN(n5362) );
  NAND2_X1 U5576 ( .A1(n9010), .A2(n9136), .ZN(n9016) );
  NAND2_X1 U5577 ( .A1(n6733), .A2(n6734), .ZN(n6792) );
  AND2_X1 U5578 ( .A1(n6792), .A2(n4562), .ZN(n9070) );
  NAND2_X1 U5579 ( .A1(n6804), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4562) );
  NOR2_X1 U5580 ( .A1(n9070), .A2(n9069), .ZN(n9068) );
  INV_X1 U5581 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7333) );
  NAND2_X1 U5582 ( .A1(n9097), .A2(n9098), .ZN(n9096) );
  NOR2_X1 U5583 ( .A1(n9578), .A2(n4407), .ZN(n9621) );
  NOR2_X1 U5584 ( .A1(n9621), .A2(n9622), .ZN(n9620) );
  NOR2_X1 U5585 ( .A1(n9639), .A2(n4564), .ZN(n9649) );
  AND2_X1 U5586 ( .A1(n9644), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4564) );
  NOR2_X1 U5587 ( .A1(n9649), .A2(n9650), .ZN(n9648) );
  NOR2_X1 U5588 ( .A1(n9648), .A2(n4563), .ZN(n9114) );
  AND2_X1 U5589 ( .A1(n9124), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4563) );
  OR2_X1 U5590 ( .A1(n9713), .A2(n9714), .ZN(n9710) );
  AOI21_X1 U5591 ( .B1(n4534), .B2(n9209), .A(n4366), .ZN(n4532) );
  NOR2_X1 U5592 ( .A1(n4583), .A2(n9394), .ZN(n9186) );
  NAND2_X1 U5593 ( .A1(n4805), .A2(n4328), .ZN(n4804) );
  NAND2_X1 U5594 ( .A1(n4812), .A2(n9195), .ZN(n4805) );
  NOR2_X1 U5595 ( .A1(n9195), .A2(n4916), .ZN(n4534) );
  AND2_X1 U5596 ( .A1(n4354), .A2(n4549), .ZN(n4548) );
  NAND2_X1 U5597 ( .A1(n4547), .A2(n9184), .ZN(n4546) );
  NAND2_X1 U5598 ( .A1(n9237), .A2(n4582), .ZN(n9210) );
  NAND2_X1 U5599 ( .A1(n4808), .A2(n4809), .ZN(n9206) );
  AND2_X1 U5600 ( .A1(n9245), .A2(n9254), .ZN(n9237) );
  NAND2_X1 U5601 ( .A1(n9237), .A2(n9419), .ZN(n9223) );
  NAND2_X1 U5602 ( .A1(n9222), .A2(n9221), .ZN(n9205) );
  NAND2_X1 U5603 ( .A1(n4817), .A2(n4815), .ZN(n9236) );
  NAND2_X1 U5604 ( .A1(n4819), .A2(n9156), .ZN(n4817) );
  NAND2_X1 U5605 ( .A1(n9282), .A2(n4816), .ZN(n4815) );
  AND2_X1 U5606 ( .A1(n4823), .A2(n9156), .ZN(n4816) );
  OAI21_X1 U5607 ( .B1(n4539), .B2(n4538), .A(n4537), .ZN(n9275) );
  AOI21_X1 U5608 ( .B1(n4329), .B2(n4335), .A(n4374), .ZN(n4537) );
  NAND2_X1 U5609 ( .A1(n4329), .A2(n4346), .ZN(n4538) );
  AND2_X1 U5610 ( .A1(n9466), .A2(n5482), .ZN(n4624) );
  NAND2_X1 U5611 ( .A1(n9373), .A2(n4574), .ZN(n9315) );
  NOR2_X1 U5612 ( .A1(n4576), .A2(n9460), .ZN(n4574) );
  OR2_X1 U5613 ( .A1(n9451), .A2(n9315), .ZN(n9291) );
  NAND2_X1 U5614 ( .A1(n8991), .A2(n8990), .ZN(n9306) );
  NAND2_X1 U5615 ( .A1(n8991), .A2(n4839), .ZN(n9307) );
  NOR2_X1 U5616 ( .A1(n9305), .A2(n4840), .ZN(n4839) );
  INV_X1 U5617 ( .A(n8990), .ZN(n4840) );
  AND2_X1 U5618 ( .A1(n8950), .A2(n8990), .ZN(n9322) );
  NAND2_X1 U5619 ( .A1(n9373), .A2(n4577), .ZN(n9341) );
  NOR2_X1 U5620 ( .A1(n5412), .A2(n5411), .ZN(n5460) );
  INV_X1 U5621 ( .A(n8975), .ZN(n7559) );
  AOI21_X1 U5622 ( .B1(n4749), .B2(n4751), .A(n4337), .ZN(n4748) );
  NAND2_X1 U5623 ( .A1(n7243), .A2(n4749), .ZN(n4747) );
  NAND2_X1 U5624 ( .A1(n7214), .A2(n8733), .ZN(n7246) );
  NAND2_X1 U5625 ( .A1(n7214), .A2(n4580), .ZN(n7409) );
  NAND2_X1 U5626 ( .A1(n7207), .A2(n7206), .ZN(n7251) );
  NAND2_X1 U5627 ( .A1(n7141), .A2(n7140), .ZN(n8810) );
  AND2_X1 U5628 ( .A1(n7149), .A2(n8606), .ZN(n7214) );
  OR2_X1 U5629 ( .A1(n8858), .A2(n9034), .ZN(n7145) );
  AND4_X1 U5630 ( .A1(n5129), .A2(n5128), .A3(n5127), .A4(n5126), .ZN(n7088)
         );
  AND4_X1 U5631 ( .A1(n5054), .A2(n5053), .A3(n5052), .A4(n5051), .ZN(n6870)
         );
  NAND2_X1 U5632 ( .A1(n6770), .A2(n8804), .ZN(n8956) );
  NAND2_X1 U5633 ( .A1(n6693), .A2(n6703), .ZN(n7039) );
  AOI21_X1 U5634 ( .B1(n5724), .B2(n5713), .A(n6598), .ZN(n6777) );
  NAND2_X1 U5635 ( .A1(n5672), .A2(n5671), .ZN(n9411) );
  AOI21_X1 U5636 ( .B1(n9282), .B2(n9281), .A(n9154), .ZN(n9263) );
  NAND2_X1 U5637 ( .A1(n4835), .A2(n5232), .ZN(n7208) );
  NAND2_X1 U5638 ( .A1(n5212), .A2(n5211), .ZN(n9779) );
  INV_X1 U5639 ( .A(n9452), .ZN(n9771) );
  AND2_X1 U5640 ( .A1(n6688), .A2(n7342), .ZN(n9452) );
  AND2_X1 U5641 ( .A1(n6453), .A2(n5019), .ZN(n9009) );
  XNOR2_X1 U5642 ( .A(n7678), .B(SI_29_), .ZN(n8793) );
  XNOR2_X1 U5643 ( .A(n5688), .B(n5687), .ZN(n7555) );
  NOR2_X1 U5644 ( .A1(n4950), .A2(n4949), .ZN(n4951) );
  INV_X1 U5645 ( .A(n4964), .ZN(n4961) );
  XNOR2_X1 U5646 ( .A(n5727), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5732) );
  NAND2_X1 U5647 ( .A1(n4753), .A2(n4336), .ZN(n4942) );
  INV_X1 U5648 ( .A(n4866), .ZN(n4865) );
  XNOR2_X1 U5649 ( .A(n5499), .B(n5498), .ZN(n7328) );
  NOR2_X1 U5650 ( .A1(n4630), .A2(n4628), .ZN(n4627) );
  OAI21_X1 U5651 ( .B1(n4629), .B2(n4628), .A(n4414), .ZN(n4626) );
  INV_X1 U5652 ( .A(n5429), .ZN(n4628) );
  NAND2_X1 U5653 ( .A1(n4936), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U5654 ( .A1(n4625), .A2(n4629), .ZN(n5430) );
  NAND2_X1 U5655 ( .A1(n5376), .A2(n4631), .ZN(n4625) );
  XNOR2_X1 U5656 ( .A(n5250), .B(n5248), .ZN(n6612) );
  NAND2_X1 U5657 ( .A1(n4614), .A2(n4616), .ZN(n5250) );
  OR2_X1 U5658 ( .A1(n5209), .A2(n5208), .ZN(n5333) );
  XNOR2_X1 U5659 ( .A(n5227), .B(n4920), .ZN(n6608) );
  OAI21_X1 U5660 ( .B1(n5200), .B2(n5199), .A(n5198), .ZN(n5227) );
  XNOR2_X1 U5661 ( .A(n5109), .B(SI_4_), .ZN(n5107) );
  CLKBUF_X1 U5662 ( .A(n4987), .Z(n4988) );
  AND2_X1 U5663 ( .A1(n7219), .A2(n6484), .ZN(n7669) );
  INV_X1 U5664 ( .A(n6894), .ZN(n6469) );
  NAND2_X1 U5665 ( .A1(n5792), .A2(n5791), .ZN(n8351) );
  OR2_X1 U5666 ( .A1(n4319), .A2(n9848), .ZN(n6464) );
  NAND2_X1 U5667 ( .A1(n4880), .A2(n6465), .ZN(n6671) );
  INV_X1 U5668 ( .A(n4881), .ZN(n4880) );
  AND2_X1 U5669 ( .A1(n6465), .A2(n6463), .ZN(n6673) );
  NAND2_X1 U5670 ( .A1(n6117), .A2(n6116), .ZN(n7804) );
  OR2_X1 U5671 ( .A1(n5849), .A2(n10066), .ZN(n6116) );
  NAND2_X1 U5672 ( .A1(n6036), .A2(n6035), .ZN(n8395) );
  NAND2_X1 U5673 ( .A1(n6514), .A2(n6513), .ZN(n7816) );
  INV_X1 U5674 ( .A(n7861), .ZN(n7871) );
  NAND2_X1 U5675 ( .A1(n6891), .A2(n6472), .ZN(n6964) );
  NAND2_X1 U5676 ( .A1(n5992), .A2(n5991), .ZN(n7599) );
  NAND2_X1 U5677 ( .A1(n7789), .A2(n7742), .ZN(n7843) );
  NAND2_X1 U5678 ( .A1(n7789), .A2(n4902), .ZN(n7844) );
  NAND2_X1 U5679 ( .A1(n6497), .A2(n6496), .ZN(n7436) );
  INV_X1 U5680 ( .A(n7879), .ZN(n7856) );
  OR2_X1 U5681 ( .A1(n6552), .A2(n6551), .ZN(n7860) );
  NAND2_X1 U5682 ( .A1(n6531), .A2(n8427), .ZN(n7876) );
  NAND2_X1 U5683 ( .A1(n7625), .A2(n6506), .ZN(n7647) );
  INV_X1 U5684 ( .A(n7874), .ZN(n7864) );
  NAND2_X1 U5685 ( .A1(n4505), .A2(n4504), .ZN(n4503) );
  INV_X1 U5686 ( .A(n7231), .ZN(n8096) );
  XNOR2_X1 U5687 ( .A(n6174), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8100) );
  AND2_X1 U5688 ( .A1(n7030), .A2(n6170), .ZN(n7779) );
  INV_X1 U5689 ( .A(n8283), .ZN(n8108) );
  OR2_X1 U5690 ( .A1(n5823), .A2(n5844), .ZN(n5846) );
  NOR2_X1 U5691 ( .A1(n4485), .A2(n4484), .ZN(n4483) );
  NOR2_X1 U5692 ( .A1(n5910), .A2(n6680), .ZN(n4484) );
  OAI21_X1 U5693 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6617), .A(n6656), .ZN(n6618) );
  NOR2_X1 U5694 ( .A1(n6839), .A2(n6840), .ZN(n6838) );
  NAND2_X1 U5695 ( .A1(n4743), .A2(n4742), .ZN(n6850) );
  AOI21_X1 U5696 ( .B1(n6370), .B2(n6856), .A(n6838), .ZN(n6560) );
  NOR2_X1 U5697 ( .A1(n6560), .A2(n6559), .ZN(n6558) );
  AOI21_X1 U5698 ( .B1(n6585), .B2(n6371), .A(n6558), .ZN(n6988) );
  NAND2_X1 U5699 ( .A1(n6988), .A2(n6987), .ZN(n6986) );
  INV_X1 U5700 ( .A(n4768), .ZN(n6319) );
  INV_X1 U5701 ( .A(n4799), .ZN(n7393) );
  INV_X1 U5702 ( .A(n4797), .ZN(n7391) );
  AOI21_X1 U5703 ( .B1(n6379), .B2(n7313), .A(n7312), .ZN(n7350) );
  NOR2_X1 U5704 ( .A1(n7350), .A2(n7349), .ZN(n7348) );
  NAND2_X1 U5705 ( .A1(n4522), .A2(n4521), .ZN(n7351) );
  NOR2_X1 U5706 ( .A1(n6385), .A2(n7614), .ZN(n8132) );
  NAND2_X1 U5707 ( .A1(n4781), .A2(n4780), .ZN(n8176) );
  NAND2_X1 U5708 ( .A1(n4507), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4506) );
  INV_X1 U5709 ( .A(n6299), .ZN(n4786) );
  INV_X1 U5710 ( .A(n8151), .ZN(n4507) );
  INV_X1 U5711 ( .A(n8249), .ZN(n9838) );
  NAND2_X1 U5712 ( .A1(n4777), .A2(n4776), .ZN(n4775) );
  OR2_X1 U5713 ( .A1(n4779), .A2(n6338), .ZN(n4777) );
  OAI21_X1 U5714 ( .B1(n6447), .B2(n9845), .A(n6446), .ZN(n8263) );
  NOR2_X1 U5715 ( .A1(n6445), .A2(n6444), .ZN(n6446) );
  NOR2_X1 U5716 ( .A1(n8283), .A2(n8390), .ZN(n6444) );
  INV_X1 U5717 ( .A(n8291), .ZN(n4677) );
  NAND2_X1 U5718 ( .A1(n4721), .A2(n4722), .ZN(n8287) );
  OAI21_X1 U5719 ( .B1(n8291), .B2(n6115), .A(n4685), .ZN(n8281) );
  NAND2_X1 U5720 ( .A1(n4725), .A2(n8038), .ZN(n8297) );
  NAND2_X1 U5721 ( .A1(n4726), .A2(n8047), .ZN(n4725) );
  INV_X1 U5722 ( .A(n8304), .ZN(n4726) );
  NAND2_X1 U5723 ( .A1(n4660), .A2(n4661), .ZN(n8345) );
  NAND2_X1 U5724 ( .A1(n4665), .A2(n4669), .ZN(n8358) );
  NAND2_X1 U5725 ( .A1(n4708), .A2(n8021), .ZN(n8361) );
  OR2_X1 U5726 ( .A1(n8369), .A2(n8371), .ZN(n4708) );
  NAND2_X1 U5727 ( .A1(n8417), .A2(n6195), .ZN(n7661) );
  NAND2_X1 U5728 ( .A1(n5980), .A2(n5979), .ZN(n8509) );
  NAND2_X1 U5729 ( .A1(n4694), .A2(n7986), .ZN(n7512) );
  NAND2_X1 U5730 ( .A1(n6191), .A2(n7421), .ZN(n4694) );
  INV_X1 U5731 ( .A(n8386), .ZN(n8419) );
  AND2_X1 U5732 ( .A1(n5932), .A2(n5931), .ZN(n9888) );
  NAND2_X1 U5733 ( .A1(n4641), .A2(n4646), .ZN(n7371) );
  INV_X1 U5734 ( .A(n4633), .ZN(n7158) );
  AOI21_X1 U5735 ( .B1(n7109), .B2(n4634), .A(n4352), .ZN(n4633) );
  INV_X1 U5736 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6895) );
  AND2_X2 U5737 ( .A1(n6254), .A2(n6253), .ZN(n9920) );
  NAND2_X1 U5738 ( .A1(n7717), .A2(n7716), .ZN(n8518) );
  AND2_X1 U5739 ( .A1(n6149), .A2(n6148), .ZN(n8076) );
  INV_X1 U5740 ( .A(n7712), .ZN(n6267) );
  INV_X1 U5741 ( .A(n7754), .ZN(n8266) );
  AOI21_X1 U5742 ( .B1(n7500), .B2(n7893), .A(n6127), .ZN(n8524) );
  INV_X1 U5743 ( .A(n7804), .ZN(n8528) );
  INV_X1 U5744 ( .A(n7767), .ZN(n8536) );
  OR2_X1 U5745 ( .A1(n8491), .A2(n8490), .ZN(n8557) );
  AND2_X1 U5746 ( .A1(n7458), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6601) );
  NAND2_X1 U5747 ( .A1(n8575), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U5748 ( .A1(n6224), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6226) );
  INV_X1 U5749 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6624) );
  INV_X1 U5750 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6614) );
  INV_X1 U5751 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6610) );
  INV_X1 U5752 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6606) );
  INV_X1 U5753 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6595) );
  INV_X1 U5754 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9991) );
  XNOR2_X1 U5755 ( .A(n5901), .B(n5915), .ZN(n6990) );
  INV_X1 U5756 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6587) );
  INV_X1 U5757 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6584) );
  INV_X1 U5758 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6582) );
  XNOR2_X1 U5759 ( .A(P2_IR_REG_2__SCAN_IN), .B(P2_IR_REG_31__SCAN_IN), .ZN(
        n4801) );
  AND4_X1 U5760 ( .A1(n5190), .A2(n5189), .A3(n5188), .A4(n5187), .ZN(n8854)
         );
  AND2_X1 U5761 ( .A1(n5676), .A2(n5746), .ZN(n9212) );
  INV_X1 U5762 ( .A(n9441), .ZN(n9138) );
  AND4_X1 U5763 ( .A1(n5541), .A2(n5540), .A3(n5539), .A4(n5538), .ZN(n9439)
         );
  AND4_X1 U5764 ( .A1(n5218), .A2(n5217), .A3(n5216), .A4(n5215), .ZN(n7265)
         );
  INV_X1 U5765 ( .A(n4861), .ZN(n4860) );
  NAND2_X1 U5766 ( .A1(n5025), .A2(n5024), .ZN(n6630) );
  NAND2_X1 U5767 ( .A1(n4849), .A2(n4851), .ZN(n8628) );
  NAND2_X1 U5768 ( .A1(n4850), .A2(n4854), .ZN(n4849) );
  INV_X1 U5769 ( .A(n8616), .ZN(n4850) );
  AND4_X1 U5770 ( .A1(n5268), .A2(n5267), .A3(n5266), .A4(n5265), .ZN(n8643)
         );
  NAND2_X1 U5771 ( .A1(n4875), .A2(n4876), .ZN(n8650) );
  NAND2_X1 U5772 ( .A1(n5621), .A2(n5620), .ZN(n9427) );
  AOI21_X1 U5773 ( .B1(n8682), .B2(n8681), .A(n8680), .ZN(n8684) );
  AND4_X1 U5774 ( .A1(n5343), .A2(n5342), .A3(n5341), .A4(n5340), .ZN(n9516)
         );
  AND4_X1 U5775 ( .A1(n5238), .A2(n5237), .A3(n5236), .A4(n5235), .ZN(n9533)
         );
  INV_X1 U5776 ( .A(n8759), .ZN(n8726) );
  AND2_X1 U5777 ( .A1(n5122), .A2(n5095), .ZN(n4858) );
  NAND2_X1 U5778 ( .A1(n4385), .A2(n4856), .ZN(n4855) );
  NAND2_X1 U5779 ( .A1(n5753), .A2(n9024), .ZN(n8763) );
  AOI21_X1 U5780 ( .B1(n9006), .B2(n7703), .A(n7342), .ZN(n4450) );
  NAND2_X1 U5781 ( .A1(n4452), .A2(n9007), .ZN(n4451) );
  AOI21_X1 U5782 ( .B1(n9008), .B2(n7342), .A(n9024), .ZN(n4448) );
  NAND4_X1 U5783 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n9038)
         );
  NOR2_X1 U5784 ( .A1(n9606), .A2(n9605), .ZN(n9604) );
  NOR2_X1 U5785 ( .A1(n9620), .A2(n4559), .ZN(n6799) );
  AND2_X1 U5786 ( .A1(n6813), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4559) );
  NAND2_X1 U5787 ( .A1(n6799), .A2(n6800), .ZN(n9112) );
  XNOR2_X1 U5788 ( .A(n9114), .B(n9126), .ZN(n9668) );
  INV_X1 U5789 ( .A(n9700), .ZN(n9718) );
  NAND2_X1 U5790 ( .A1(n4333), .A2(n9696), .ZN(n4570) );
  NAND2_X1 U5791 ( .A1(n4567), .A2(n9110), .ZN(n4566) );
  NAND2_X1 U5792 ( .A1(n9616), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U5793 ( .A1(n8776), .A2(n8775), .ZN(n9148) );
  OAI21_X1 U5794 ( .B1(n9248), .B2(n4551), .A(n4549), .ZN(n9220) );
  INV_X1 U5795 ( .A(n9427), .ZN(n9245) );
  NOR2_X1 U5796 ( .A1(n4356), .A2(n9182), .ZN(n9233) );
  NAND2_X1 U5797 ( .A1(n4386), .A2(n4818), .ZN(n9250) );
  AND2_X1 U5798 ( .A1(n5589), .A2(n5588), .ZN(n9249) );
  AND2_X1 U5799 ( .A1(n5534), .A2(n5533), .ZN(n9280) );
  AND2_X1 U5800 ( .A1(n5506), .A2(n5505), .ZN(n9295) );
  OAI21_X1 U5801 ( .B1(n9321), .B2(n4543), .A(n4329), .ZN(n9289) );
  AND2_X1 U5802 ( .A1(n5515), .A2(n5514), .ZN(n9458) );
  AOI21_X1 U5803 ( .B1(n9321), .B2(n9178), .A(n4541), .ZN(n4540) );
  INV_X1 U5804 ( .A(n4909), .ZN(n4541) );
  NAND2_X1 U5805 ( .A1(n5459), .A2(n5458), .ZN(n9350) );
  OR2_X1 U5806 ( .A1(n7167), .A2(n5452), .ZN(n5459) );
  NAND2_X1 U5807 ( .A1(n4761), .A2(n9172), .ZN(n9371) );
  NAND2_X1 U5808 ( .A1(n9171), .A2(n4922), .ZN(n4761) );
  AND2_X1 U5809 ( .A1(n5361), .A2(n5360), .ZN(n9170) );
  NAND2_X1 U5810 ( .A1(n7485), .A2(n8891), .ZN(n7486) );
  OAI21_X1 U5811 ( .B1(n7243), .B2(n4751), .A(n4749), .ZN(n7489) );
  NAND2_X1 U5812 ( .A1(n7406), .A2(n7405), .ZN(n7408) );
  AND4_X1 U5813 ( .A1(n5290), .A2(n5289), .A3(n5288), .A4(n5287), .ZN(n9531)
         );
  INV_X1 U5814 ( .A(n8849), .ZN(n8857) );
  NAND2_X1 U5815 ( .A1(n4463), .A2(n8841), .ZN(n7089) );
  OR2_X1 U5816 ( .A1(n8794), .A2(n6573), .ZN(n5039) );
  AND2_X1 U5817 ( .A1(n5040), .A2(n4345), .ZN(n4553) );
  OR2_X1 U5818 ( .A1(n4322), .A2(n7017), .ZN(n9738) );
  OR2_X1 U5819 ( .A1(n7016), .A2(n9136), .ZN(n9735) );
  INV_X1 U5820 ( .A(n9369), .ZN(n9742) );
  INV_X1 U5821 ( .A(n9041), .ZN(n7687) );
  INV_X1 U5822 ( .A(n9733), .ZN(n9722) );
  NAND2_X1 U5823 ( .A1(n9396), .A2(n9395), .ZN(n9397) );
  OAI21_X1 U5824 ( .B1(n9406), .B2(n9766), .A(n4377), .ZN(n9545) );
  AND2_X1 U5825 ( .A1(n9405), .A2(n4834), .ZN(n4833) );
  NAND2_X1 U5826 ( .A1(n6596), .A2(n9009), .ZN(n9745) );
  XNOR2_X1 U5827 ( .A(n7892), .B(n7891), .ZN(n9569) );
  NAND2_X1 U5828 ( .A1(n4994), .A2(n4993), .ZN(n4996) );
  NAND2_X1 U5829 ( .A1(n4468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4993) );
  OAI21_X1 U5830 ( .B1(n4466), .B2(n4360), .A(n4465), .ZN(n4994) );
  NAND2_X1 U5831 ( .A1(n4977), .A2(n4976), .ZN(n4980) );
  NAND2_X1 U5832 ( .A1(n4978), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4976) );
  AOI21_X1 U5833 ( .B1(n4973), .B2(n4975), .A(n4949), .ZN(n4554) );
  NAND2_X1 U5834 ( .A1(n4963), .A2(n4962), .ZN(n7482) );
  NOR2_X1 U5835 ( .A1(n4961), .A2(n4960), .ZN(n4962) );
  OAI21_X1 U5836 ( .B1(n4953), .B2(n4952), .A(n4951), .ZN(n4963) );
  NOR2_X1 U5837 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4960) );
  XNOR2_X1 U5838 ( .A(n5557), .B(n5578), .ZN(n7457) );
  AND2_X1 U5839 ( .A1(n5552), .A2(n5579), .ZN(n5557) );
  INV_X1 U5840 ( .A(n5732), .ZN(n9010) );
  XNOR2_X1 U5841 ( .A(n4947), .B(n4955), .ZN(n7379) );
  INV_X1 U5842 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6625) );
  XNOR2_X1 U5843 ( .A(n5181), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9609) );
  XNOR2_X1 U5844 ( .A(n4689), .B(n5172), .ZN(n6594) );
  NAND2_X1 U5845 ( .A1(n4827), .A2(n5157), .ZN(n4689) );
  AND2_X1 U5846 ( .A1(n5180), .A2(n5160), .ZN(n9597) );
  NOR2_X1 U5847 ( .A1(n5140), .A2(n5139), .ZN(n9089) );
  INV_X1 U5848 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6579) );
  INV_X1 U5849 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6577) );
  INV_X1 U5850 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U5851 ( .A1(n9830), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U5852 ( .A1(n4793), .A2(n4792), .ZN(n8202) );
  NAND2_X1 U5853 ( .A1(n8258), .A2(n9816), .ZN(n4444) );
  NOR2_X1 U5854 ( .A1(n4441), .A2(n8257), .ZN(n4440) );
  NAND2_X1 U5855 ( .A1(n9816), .A2(n4775), .ZN(n4772) );
  AOI21_X1 U5856 ( .B1(n4524), .B2(n9808), .A(n4340), .ZN(n4778) );
  AND2_X1 U5857 ( .A1(n4712), .A2(n4713), .ZN(n7727) );
  NOR2_X1 U5858 ( .A1(n9906), .A2(n9845), .ZN(n4709) );
  NAND2_X1 U5859 ( .A1(n4568), .A2(n4565), .ZN(P1_U3262) );
  NAND2_X1 U5860 ( .A1(n4569), .A2(n9136), .ZN(n4568) );
  AOI21_X1 U5861 ( .B1(n9137), .B2(n7703), .A(n4566), .ZN(n4565) );
  NAND2_X1 U5862 ( .A1(n9135), .A2(n4570), .ZN(n4569) );
  NAND2_X1 U5863 ( .A1(n4832), .A2(n4831), .ZN(P1_U3518) );
  NAND2_X1 U5864 ( .A1(n9787), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n4831) );
  NAND2_X1 U5865 ( .A1(n9545), .A2(n9789), .ZN(n4832) );
  AND2_X1 U5866 ( .A1(n4851), .A2(n4848), .ZN(n4327) );
  AND2_X1 U5867 ( .A1(n4809), .A2(n9194), .ZN(n4328) );
  AND2_X1 U5868 ( .A1(n4542), .A2(n4910), .ZN(n4329) );
  NAND4_X1 U5869 ( .A1(n5848), .A2(n5847), .A3(n5846), .A4(n5845), .ZN(n8126)
         );
  INV_X1 U5870 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U5871 ( .A1(n4754), .A2(n4753), .ZN(n4964) );
  OR2_X1 U5872 ( .A1(n8198), .A2(n6301), .ZN(n4330) );
  NAND2_X1 U5873 ( .A1(n6184), .A2(n7944), .ZN(n7907) );
  NAND2_X1 U5874 ( .A1(n8509), .A2(n8119), .ZN(n4331) );
  AND2_X1 U5875 ( .A1(n8524), .A2(n8283), .ZN(n4332) );
  INV_X1 U5876 ( .A(n9195), .ZN(n4806) );
  AOI21_X1 U5877 ( .B1(n9248), .B2(n4548), .A(n4546), .ZN(n4545) );
  AND2_X1 U5878 ( .A1(n8015), .A2(n8021), .ZN(n8370) );
  INV_X1 U5879 ( .A(n4540), .ZN(n9309) );
  XOR2_X1 U5880 ( .A(n9133), .B(n9132), .Z(n4333) );
  AND2_X1 U5881 ( .A1(n5774), .A2(n4387), .ZN(n5794) );
  INV_X1 U5882 ( .A(n7948), .ZN(n4481) );
  XNOR2_X1 U5883 ( .A(n5799), .B(n5798), .ZN(n5815) );
  AND2_X1 U5884 ( .A1(n4722), .A2(n8054), .ZN(n4334) );
  INV_X1 U5885 ( .A(n4598), .ZN(n4597) );
  OAI21_X1 U5886 ( .B1(n4603), .B2(n4599), .A(n5303), .ZN(n4598) );
  AND2_X1 U5887 ( .A1(n8948), .A2(n9194), .ZN(n9209) );
  AND4_X1 U5888 ( .A1(n6067), .A2(n6066), .A3(n6065), .A4(n6064), .ZN(n8375)
         );
  AND2_X1 U5889 ( .A1(n4543), .A2(n4346), .ZN(n4335) );
  INV_X1 U5890 ( .A(n8302), .ZN(n8110) );
  AND2_X1 U5891 ( .A1(n6114), .A2(n6113), .ZN(n8302) );
  INV_X1 U5892 ( .A(n4854), .ZN(n4853) );
  INV_X1 U5893 ( .A(n9460), .ZN(n9316) );
  NAND2_X1 U5894 ( .A1(n5483), .A2(n5482), .ZN(n9460) );
  AND2_X1 U5895 ( .A1(n4939), .A2(n4865), .ZN(n4336) );
  AND2_X1 U5896 ( .A1(n8708), .A2(n9508), .ZN(n4337) );
  AND2_X1 U5897 ( .A1(n8513), .A2(n8093), .ZN(n4338) );
  AND4_X1 U5898 ( .A1(n5874), .A2(n5873), .A3(n5872), .A4(n5871), .ZN(n7160)
         );
  INV_X1 U5899 ( .A(n7160), .ZN(n8125) );
  AND2_X1 U5900 ( .A1(n7744), .A2(n8112), .ZN(n4339) );
  OR2_X1 U5901 ( .A1(n6416), .A2(n6415), .ZN(n4340) );
  NAND2_X1 U5902 ( .A1(n4535), .A2(n4536), .ZN(n4341) );
  AND3_X1 U5903 ( .A1(n5091), .A2(n5090), .A3(n5089), .ZN(n9755) );
  AND2_X1 U5904 ( .A1(n4581), .A2(n4582), .ZN(n4342) );
  NAND2_X1 U5905 ( .A1(n4843), .A2(n5246), .ZN(n8604) );
  INV_X2 U5906 ( .A(n4948), .ZN(n7703) );
  INV_X1 U5907 ( .A(n6574), .ZN(n4586) );
  NAND2_X1 U5908 ( .A1(n5774), .A2(n5773), .ZN(n6175) );
  AND2_X1 U5909 ( .A1(n4875), .A2(n4873), .ZN(n4343) );
  NAND3_X1 U5910 ( .A1(n5858), .A2(n5857), .A3(n5856), .ZN(n5867) );
  OR2_X1 U5911 ( .A1(n9572), .A2(n4998), .ZN(n5074) );
  NAND2_X1 U5912 ( .A1(n4988), .A2(n4928), .ZN(n5031) );
  AND2_X1 U5913 ( .A1(n5042), .A2(n5041), .ZN(n4344) );
  INV_X1 U5914 ( .A(n4813), .ZN(n4823) );
  OR2_X1 U5915 ( .A1(n4312), .A2(n6747), .ZN(n4345) );
  NAND2_X1 U5916 ( .A1(n9295), .A2(n9458), .ZN(n4346) );
  INV_X1 U5917 ( .A(n5072), .ZN(n5512) );
  INV_X1 U5918 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4468) );
  NOR2_X1 U5919 ( .A1(n6068), .A2(n4670), .ZN(n4664) );
  AND2_X1 U5920 ( .A1(n6194), .A2(n8000), .ZN(n4347) );
  NAND2_X1 U5921 ( .A1(n5276), .A2(n5258), .ZN(n5277) );
  INV_X1 U5922 ( .A(n6692), .ZN(n6693) );
  NAND2_X1 U5923 ( .A1(n5198), .A2(n5179), .ZN(n5199) );
  AND2_X1 U5924 ( .A1(n4745), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4348) );
  NAND2_X1 U5925 ( .A1(n4801), .A2(n4800), .ZN(n4349) );
  NAND2_X1 U5926 ( .A1(n8403), .A2(n6193), .ZN(n4350) );
  OR2_X1 U5927 ( .A1(n9433), .A2(n9438), .ZN(n9156) );
  INV_X1 U5928 ( .A(n8884), .ZN(n7487) );
  AND2_X1 U5929 ( .A1(n4519), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4351) );
  AND2_X1 U5930 ( .A1(n7160), .A2(n9867), .ZN(n4352) );
  NAND2_X1 U5931 ( .A1(n9460), .A2(n9466), .ZN(n4353) );
  OR2_X1 U5932 ( .A1(n9229), .A2(n9242), .ZN(n4354) );
  INV_X1 U5933 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4974) );
  INV_X1 U5934 ( .A(n9159), .ZN(n4810) );
  NAND2_X1 U5935 ( .A1(n4992), .A2(n4468), .ZN(n4995) );
  AND2_X1 U5936 ( .A1(n4351), .A2(n6585), .ZN(n4355) );
  AND2_X1 U5937 ( .A1(n9248), .A2(n9183), .ZN(n4356) );
  AND2_X1 U5938 ( .A1(n8935), .A2(n8997), .ZN(n9185) );
  INV_X1 U5939 ( .A(n9185), .ZN(n4531) );
  NAND2_X1 U5940 ( .A1(n5410), .A2(n5409), .ZN(n9487) );
  NAND2_X1 U5941 ( .A1(n5774), .A2(n4638), .ZN(n5777) );
  AND2_X1 U5942 ( .A1(n7912), .A2(n4644), .ZN(n4357) );
  AND2_X1 U5943 ( .A1(n4532), .A2(n4531), .ZN(n4358) );
  AND2_X1 U5944 ( .A1(n5880), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n4359) );
  AND3_X1 U5945 ( .A1(n4959), .A2(n4752), .A3(n4467), .ZN(n4360) );
  AND2_X1 U5946 ( .A1(n9427), .A2(n9415), .ZN(n4361) );
  INV_X1 U5947 ( .A(n4688), .ZN(n9882) );
  OAI211_X1 U5948 ( .C1(n6594), .C2(n6054), .A(n5921), .B(n5920), .ZN(n4688)
         );
  INV_X1 U5949 ( .A(n8021), .ZN(n4707) );
  NAND2_X1 U5950 ( .A1(n5262), .A2(n5261), .ZN(n9535) );
  INV_X1 U5951 ( .A(n9155), .ZN(n4822) );
  NAND2_X1 U5952 ( .A1(n5438), .A2(n5437), .ZN(n9324) );
  INV_X1 U5953 ( .A(n9324), .ZN(n4623) );
  OR2_X1 U5954 ( .A1(n8070), .A2(n7938), .ZN(n4362) );
  INV_X1 U5955 ( .A(n4583), .ZN(n9199) );
  NAND2_X1 U5956 ( .A1(n9237), .A2(n4342), .ZN(n4583) );
  AOI21_X1 U5957 ( .B1(n5199), .B2(n5198), .A(n4620), .ZN(n4619) );
  AND2_X1 U5958 ( .A1(n9307), .A2(n9151), .ZN(n4363) );
  INV_X1 U5959 ( .A(n6283), .ZN(n4518) );
  INV_X1 U5960 ( .A(n4757), .ZN(n4756) );
  AOI21_X1 U5961 ( .B1(n4759), .B2(n4758), .A(n4372), .ZN(n4757) );
  INV_X1 U5962 ( .A(n9229), .ZN(n9419) );
  NAND2_X1 U5963 ( .A1(n5646), .A2(n5645), .ZN(n9229) );
  INV_X1 U5964 ( .A(n4600), .ZN(n4599) );
  NOR2_X1 U5965 ( .A1(n5304), .A2(n4601), .ZN(n4600) );
  NAND2_X1 U5966 ( .A1(n4510), .A2(n4517), .ZN(n4364) );
  INV_X1 U5967 ( .A(n4664), .ZN(n4663) );
  NAND2_X1 U5968 ( .A1(n7908), .A2(n7969), .ZN(n4365) );
  AND2_X1 U5969 ( .A1(n9401), .A2(n9166), .ZN(n4366) );
  AND2_X1 U5970 ( .A1(n7782), .A2(n8077), .ZN(n4367) );
  OR2_X1 U5971 ( .A1(n5008), .A2(n5007), .ZN(n4368) );
  AND2_X1 U5972 ( .A1(n4814), .A2(n4818), .ZN(n4369) );
  NAND2_X1 U5973 ( .A1(n5336), .A2(n5335), .ZN(n9510) );
  AND2_X1 U5974 ( .A1(n7990), .A2(n7989), .ZN(n7916) );
  AND2_X1 U5975 ( .A1(n9015), .A2(n4474), .ZN(n4370) );
  AND4_X1 U5976 ( .A1(n8861), .A2(n8865), .A3(n8870), .A4(n8860), .ZN(n4371)
         );
  AND2_X1 U5977 ( .A1(n9494), .A2(n9363), .ZN(n4372) );
  NAND2_X1 U5978 ( .A1(n8796), .A2(n8795), .ZN(n9394) );
  OR2_X1 U5979 ( .A1(n7804), .A2(n8293), .ZN(n8054) );
  NOR2_X1 U5980 ( .A1(n8509), .A2(n8119), .ZN(n4373) );
  INV_X1 U5981 ( .A(n4670), .ZN(n4669) );
  NOR2_X1 U5982 ( .A1(n8488), .A2(n8391), .ZN(n4670) );
  INV_X1 U5983 ( .A(n4576), .ZN(n4575) );
  NAND2_X1 U5984 ( .A1(n4577), .A2(n4623), .ZN(n4576) );
  NOR2_X1 U5985 ( .A1(n6175), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n6172) );
  AND2_X1 U5986 ( .A1(n9451), .A2(n9283), .ZN(n4374) );
  AND3_X1 U5987 ( .A1(n6221), .A2(n6252), .A3(n6225), .ZN(n4375) );
  AND2_X1 U5988 ( .A1(n9245), .A2(n9227), .ZN(n4376) );
  INV_X1 U5989 ( .A(n8027), .ZN(n4703) );
  INV_X1 U5990 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5773) );
  NOR2_X1 U5991 ( .A1(n9372), .A2(n4760), .ZN(n4759) );
  AND2_X1 U5992 ( .A1(n4833), .A2(n9404), .ZN(n4377) );
  XNOR2_X1 U5993 ( .A(n5327), .B(SI_13_), .ZN(n5325) );
  AND2_X1 U5994 ( .A1(n4791), .A2(n4790), .ZN(n4378) );
  AND2_X1 U5995 ( .A1(n5497), .A2(n8690), .ZN(n4379) );
  AND2_X1 U5996 ( .A1(n5522), .A2(n5521), .ZN(n4380) );
  AND2_X1 U5997 ( .A1(n5174), .A2(SI_7_), .ZN(n4381) );
  INV_X1 U5998 ( .A(n8556), .ZN(n6198) );
  AND2_X1 U5999 ( .A1(n6059), .A2(n6058), .ZN(n8556) );
  AND2_X1 U6000 ( .A1(n8536), .A2(n8111), .ZN(n8041) );
  NAND2_X1 U6001 ( .A1(n8054), .A2(n8055), .ZN(n8286) );
  INV_X1 U6002 ( .A(n8286), .ZN(n4682) );
  INV_X1 U6003 ( .A(n8532), .ZN(n7829) );
  AND2_X1 U6004 ( .A1(n6107), .A2(n6106), .ZN(n8532) );
  NAND2_X1 U6005 ( .A1(n7877), .A2(n8108), .ZN(n4382) );
  NAND2_X1 U6006 ( .A1(n6856), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4383) );
  AND2_X1 U6007 ( .A1(n8691), .A2(n5496), .ZN(n4384) );
  NAND2_X1 U6008 ( .A1(n6914), .A2(n6913), .ZN(n4385) );
  AND2_X1 U6009 ( .A1(n4821), .A2(n9155), .ZN(n4386) );
  INV_X1 U6010 ( .A(n4812), .ZN(n4811) );
  NAND2_X1 U6011 ( .A1(n9209), .A2(n9221), .ZN(n4812) );
  INV_X1 U6012 ( .A(n7993), .ZN(n4486) );
  AND3_X1 U6013 ( .A1(n5853), .A2(n5852), .A3(n5851), .ZN(n9855) );
  INV_X1 U6014 ( .A(n9855), .ZN(n5854) );
  AND2_X1 U6015 ( .A1(n4638), .A2(n5778), .ZN(n4387) );
  AOI21_X1 U6016 ( .B1(n6264), .B2(n8436), .A(n6263), .ZN(n7709) );
  AND2_X1 U6017 ( .A1(n4578), .A2(n8596), .ZN(n4388) );
  NAND2_X1 U6018 ( .A1(n5833), .A2(n5832), .ZN(n9850) );
  AND2_X1 U6019 ( .A1(n8910), .A2(n8992), .ZN(n4389) );
  NOR2_X1 U6020 ( .A1(n8901), .A2(n9016), .ZN(n4390) );
  AND2_X1 U6021 ( .A1(n4648), .A2(n8434), .ZN(n4391) );
  INV_X1 U6022 ( .A(n7738), .ZN(n8544) );
  NAND2_X1 U6023 ( .A1(n6079), .A2(n6078), .ZN(n7738) );
  AND2_X1 U6024 ( .A1(n7991), .A2(n7992), .ZN(n4392) );
  NOR2_X1 U6025 ( .A1(n8045), .A2(n8044), .ZN(n4724) );
  AND2_X1 U6026 ( .A1(n6507), .A2(n6506), .ZN(n4393) );
  OR2_X1 U6027 ( .A1(n8351), .A2(n8360), .ZN(n8023) );
  AND2_X1 U6028 ( .A1(n4785), .A2(n4784), .ZN(n4394) );
  AND2_X1 U6029 ( .A1(n4811), .A2(n4806), .ZN(n4395) );
  AND2_X1 U6030 ( .A1(n6488), .A2(n4896), .ZN(n4396) );
  AND2_X1 U6031 ( .A1(n4795), .A2(n4330), .ZN(n4397) );
  AND2_X1 U6032 ( .A1(n4469), .A2(n4753), .ZN(n4398) );
  OR2_X1 U6033 ( .A1(n4533), .A2(n4531), .ZN(n4399) );
  AND2_X1 U6034 ( .A1(n5039), .A2(n4553), .ZN(n9749) );
  AND2_X1 U6035 ( .A1(n4767), .A2(n4766), .ZN(n4400) );
  NAND2_X1 U6036 ( .A1(n5774), .A2(n4637), .ZN(n4401) );
  INV_X1 U6037 ( .A(n4658), .ZN(n4657) );
  NAND2_X1 U6038 ( .A1(n4661), .A2(n4659), .ZN(n4658) );
  OR2_X1 U6039 ( .A1(n6198), .A2(n8375), .ZN(n8024) );
  INV_X1 U6040 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4755) );
  INV_X1 U6041 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4905) );
  INV_X1 U6042 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U6043 ( .A1(n6146), .A2(n6145), .ZN(n8107) );
  NAND2_X1 U6044 ( .A1(n5696), .A2(n5695), .ZN(n9401) );
  INV_X1 U6045 ( .A(n9401), .ZN(n4581) );
  INV_X1 U6046 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4611) );
  XOR2_X1 U6047 ( .A(n8524), .B(n4319), .Z(n4402) );
  INV_X1 U6048 ( .A(n7786), .ZN(n4900) );
  AND2_X1 U6049 ( .A1(n7214), .A2(n4578), .ZN(n4403) );
  AND2_X1 U6050 ( .A1(n9373), .A2(n9357), .ZN(n4404) );
  AND2_X1 U6051 ( .A1(n9373), .A2(n4575), .ZN(n4405) );
  INV_X1 U6052 ( .A(n7397), .ZN(n6604) );
  INV_X1 U6053 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U6054 ( .A1(n7564), .A2(n7563), .ZN(n9171) );
  OR2_X1 U6055 ( .A1(n8895), .A2(n8817), .ZN(n4406) );
  INV_X1 U6056 ( .A(n9829), .ZN(n6593) );
  AND2_X1 U6057 ( .A1(n5919), .A2(n5934), .ZN(n9829) );
  AND2_X1 U6058 ( .A1(n9583), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4407) );
  INV_X1 U6059 ( .A(n4699), .ZN(n4705) );
  NAND2_X1 U6060 ( .A1(n5483), .A2(n4624), .ZN(n9151) );
  OR2_X1 U6061 ( .A1(n5358), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n4408) );
  INV_X1 U6062 ( .A(n7352), .ZN(n4523) );
  INV_X1 U6063 ( .A(n4753), .ZN(n5358) );
  AND4_X1 U6064 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n9508)
         );
  NOR2_X1 U6065 ( .A1(n8150), .A2(n6299), .ZN(n4409) );
  OR2_X1 U6066 ( .A1(n5974), .A2(n7505), .ZN(n5975) );
  NAND2_X1 U6067 ( .A1(n5768), .A2(n5767), .ZN(n5950) );
  AND2_X1 U6068 ( .A1(n9160), .A2(n8947), .ZN(n9195) );
  INV_X1 U6069 ( .A(n4631), .ZN(n4630) );
  NOR2_X1 U6070 ( .A1(n5405), .A2(n4632), .ZN(n4631) );
  INV_X1 U6071 ( .A(n9178), .ZN(n4544) );
  AND2_X1 U6072 ( .A1(n4761), .A2(n4759), .ZN(n4410) );
  NOR2_X1 U6073 ( .A1(n9291), .A2(n9446), .ZN(n9265) );
  AND2_X1 U6074 ( .A1(n4708), .A2(n4706), .ZN(n4411) );
  AND2_X1 U6075 ( .A1(n5327), .A2(SI_13_), .ZN(n4412) );
  AND2_X1 U6076 ( .A1(n5404), .A2(n5403), .ZN(n4413) );
  OR2_X1 U6077 ( .A1(n5428), .A2(SI_17_), .ZN(n4414) );
  AND2_X1 U6078 ( .A1(n6192), .A2(n8000), .ZN(n4415) );
  OR2_X1 U6079 ( .A1(n7352), .A2(n5939), .ZN(n4416) );
  AND2_X1 U6080 ( .A1(n5246), .A2(n8720), .ZN(n4417) );
  OR2_X1 U6081 ( .A1(n4918), .A2(n6440), .ZN(n4418) );
  INV_X1 U6082 ( .A(n4687), .ZN(n4686) );
  NOR2_X1 U6083 ( .A1(n8536), .A2(n8312), .ZN(n4687) );
  NOR2_X1 U6084 ( .A1(n5377), .A2(SI_15_), .ZN(n5375) );
  INV_X1 U6085 ( .A(n4916), .ZN(n4536) );
  NOR2_X1 U6086 ( .A1(n4322), .A2(n7094), .ZN(n4419) );
  INV_X2 U6087 ( .A(n9906), .ZN(n9905) );
  NAND2_X1 U6088 ( .A1(n4980), .A2(n4979), .ZN(n5740) );
  OR2_X1 U6089 ( .A1(n6616), .A2(n8098), .ZN(n9825) );
  NAND2_X1 U6090 ( .A1(n6861), .A2(n5100), .ZN(n6912) );
  OR2_X1 U6091 ( .A1(n6323), .A2(n6290), .ZN(n4420) );
  NAND2_X1 U6092 ( .A1(n4860), .A2(n4863), .ZN(n7258) );
  NAND2_X1 U6093 ( .A1(n4859), .A2(n5095), .ZN(n6861) );
  NOR2_X1 U6094 ( .A1(n7318), .A2(n6289), .ZN(n4421) );
  NAND2_X1 U6095 ( .A1(n6824), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4422) );
  XNOR2_X1 U6096 ( .A(n5776), .B(n5793), .ZN(n6205) );
  XNOR2_X1 U6097 ( .A(n4554), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6711) );
  NAND2_X1 U6098 ( .A1(n6419), .A2(n7900), .ZN(n8436) );
  AND3_X1 U6099 ( .A1(n5879), .A2(n5878), .A3(n5877), .ZN(n9867) );
  INV_X1 U6100 ( .A(n9867), .ZN(n4635) );
  NAND2_X1 U6101 ( .A1(n5836), .A2(n4483), .ZN(n8127) );
  INV_X1 U6102 ( .A(n8127), .ZN(n4482) );
  NAND2_X1 U6103 ( .A1(n4573), .A2(n4572), .ZN(n7049) );
  INV_X1 U6104 ( .A(n7049), .ZN(n4571) );
  OR2_X1 U6105 ( .A1(n8238), .A2(n8221), .ZN(n4423) );
  OR2_X1 U6106 ( .A1(n8216), .A2(n8494), .ZN(n4424) );
  OR2_X1 U6107 ( .A1(n8216), .A2(n8397), .ZN(n4425) );
  AND2_X1 U6108 ( .A1(n7502), .A2(n7454), .ZN(n4426) );
  AND2_X1 U6109 ( .A1(n4517), .A2(n4516), .ZN(n4427) );
  INV_X1 U6110 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4609) );
  INV_X1 U6111 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n4428) );
  XNOR2_X1 U6112 ( .A(n6331), .B(n8198), .ZN(n8192) );
  XNOR2_X1 U6113 ( .A(n6335), .B(n8233), .ZN(n8227) );
  XNOR2_X1 U6114 ( .A(n6302), .B(n8233), .ZN(n8220) );
  AOI21_X1 U6115 ( .B1(n9569), .B2(n8792), .A(n8768), .ZN(n9388) );
  NAND2_X1 U6116 ( .A1(n6612), .A2(n8792), .ZN(n4835) );
  NAND2_X1 U6117 ( .A1(n7075), .A2(n6479), .ZN(n7221) );
  NAND2_X1 U6118 ( .A1(n6782), .A2(n6468), .ZN(n6893) );
  NAND2_X1 U6119 ( .A1(n4439), .A2(n4438), .ZN(n7737) );
  NOR2_X1 U6120 ( .A1(n7869), .A2(n4912), .ZN(n7756) );
  INV_X1 U6121 ( .A(n5774), .ZN(n6179) );
  INV_X1 U6122 ( .A(n6233), .ZN(n4429) );
  OAI21_X1 U6123 ( .B1(n7219), .B2(n4897), .A(n4396), .ZN(n6494) );
  NAND2_X1 U6124 ( .A1(n6891), .A2(n4904), .ZN(n7073) );
  NAND2_X4 U6125 ( .A1(n4430), .A2(n6459), .ZN(n7774) );
  NAND2_X1 U6126 ( .A1(n6457), .A2(n6456), .ZN(n4430) );
  NAND2_X1 U6127 ( .A1(n6470), .A2(n6469), .ZN(n6891) );
  NAND2_X1 U6128 ( .A1(n6231), .A2(n6230), .ZN(n6233) );
  NAND2_X1 U6129 ( .A1(n6518), .A2(n7852), .ZN(n7855) );
  NAND3_X1 U6130 ( .A1(n4311), .A2(n5761), .A3(n5760), .ZN(P1_U3220) );
  NAND2_X1 U6131 ( .A1(n4443), .A2(n4442), .ZN(n4441) );
  NOR2_X1 U6132 ( .A1(n9824), .A2(n5907), .ZN(n9823) );
  NAND3_X1 U6133 ( .A1(n4511), .A2(n4512), .A3(n4434), .ZN(n6565) );
  NAND2_X1 U6134 ( .A1(n4444), .A2(n4440), .ZN(P2_U3200) );
  NAND2_X1 U6135 ( .A1(n4881), .A2(n6465), .ZN(n6783) );
  NAND2_X1 U6136 ( .A1(n7801), .A2(n7752), .ZN(n7753) );
  NAND2_X1 U6137 ( .A1(n7855), .A2(n6521), .ZN(n6527) );
  NAND2_X1 U6138 ( .A1(n6081), .A2(n6080), .ZN(n6091) );
  NAND2_X1 U6139 ( .A1(n6119), .A2(n6118), .ZN(n6128) );
  NAND2_X1 U6140 ( .A1(n5813), .A2(n10033), .ZN(n6071) );
  MUX2_X2 U6141 ( .A(n8087), .B(n8086), .S(n8085), .Z(n8089) );
  NAND2_X1 U6142 ( .A1(n5811), .A2(n5810), .ZN(n6037) );
  NAND2_X1 U6143 ( .A1(n5809), .A2(n5808), .ZN(n6007) );
  NAND2_X1 U6144 ( .A1(n5803), .A2(n5802), .ZN(n5894) );
  NAND2_X1 U6145 ( .A1(n5807), .A2(n5806), .ZN(n5956) );
  NAND2_X1 U6146 ( .A1(n5805), .A2(n5804), .ZN(n5924) );
  NAND2_X1 U6147 ( .A1(n5812), .A2(n10048), .ZN(n6061) );
  NAND2_X1 U6148 ( .A1(n6783), .A2(n6784), .ZN(n6782) );
  OAI21_X1 U6149 ( .B1(n4924), .B2(n8079), .A(n4498), .ZN(n8084) );
  INV_X1 U6150 ( .A(n6527), .ZN(n4439) );
  NAND2_X1 U6151 ( .A1(n7648), .A2(n6510), .ZN(n7810) );
  NAND2_X1 U6152 ( .A1(n8075), .A2(n8074), .ZN(n4502) );
  AOI21_X1 U6153 ( .B1(n8091), .B2(n8090), .A(n4503), .ZN(n8097) );
  NOR2_X1 U6154 ( .A1(n8227), .A2(n8380), .ZN(n8226) );
  NOR2_X1 U6155 ( .A1(n6993), .A2(n6992), .ZN(n6991) );
  NOR2_X1 U6156 ( .A1(n9821), .A2(n6320), .ZN(n7384) );
  NOR2_X1 U6157 ( .A1(n7382), .A2(n4445), .ZN(n6321) );
  NAND2_X1 U6158 ( .A1(n8244), .A2(n8245), .ZN(n8247) );
  NAND2_X1 U6159 ( .A1(n8160), .A2(n6392), .ZN(n8170) );
  AOI21_X1 U6160 ( .B1(n6367), .B2(n6588), .A(n9800), .ZN(n6639) );
  INV_X1 U6161 ( .A(n6847), .ZN(n4745) );
  AOI21_X1 U6162 ( .B1(n7536), .B2(n6504), .A(n6503), .ZN(n7627) );
  NAND2_X1 U6163 ( .A1(n6327), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n8133) );
  NOR2_X1 U6164 ( .A1(n7316), .A2(n7430), .ZN(n7315) );
  NAND2_X2 U6165 ( .A1(n5027), .A2(n5026), .ZN(n6627) );
  OR2_X1 U6166 ( .A1(n4940), .A2(n4949), .ZN(n5408) );
  NAND2_X1 U6167 ( .A1(n4861), .A2(n4863), .ZN(n7330) );
  MUX2_X1 U6168 ( .A(n8890), .B(n8889), .S(n9016), .Z(n8898) );
  MUX2_X2 U6169 ( .A(n8929), .B(n8943), .S(n9161), .Z(n8930) );
  NAND2_X1 U6170 ( .A1(n8899), .A2(n9361), .ZN(n4460) );
  NAND2_X1 U6171 ( .A1(n4456), .A2(n4390), .ZN(n4455) );
  NAND3_X1 U6172 ( .A1(n8864), .A2(n4446), .A3(n4371), .ZN(n8871) );
  NAND2_X1 U6173 ( .A1(n4451), .A2(n4450), .ZN(n4449) );
  NAND2_X1 U6174 ( .A1(n4449), .A2(n4448), .ZN(n4447) );
  OAI21_X1 U6175 ( .B1(n4591), .B2(n4589), .A(n8924), .ZN(n8925) );
  OAI22_X1 U6176 ( .A1(n9013), .A2(n8946), .B1(n7703), .B2(n8957), .ZN(n4452)
         );
  NAND2_X1 U6177 ( .A1(n8162), .A2(n8161), .ZN(n8160) );
  NAND3_X1 U6178 ( .A1(n9022), .A2(n9023), .A3(n4447), .ZN(P1_U3242) );
  OAI21_X1 U6179 ( .B1(n4453), .B2(n4406), .A(n8952), .ZN(n8894) );
  AOI21_X1 U6180 ( .B1(n8892), .B2(n8891), .A(n4454), .ZN(n4453) );
  AND3_X1 U6181 ( .A1(n4457), .A2(n4455), .A3(n4389), .ZN(n8914) );
  NAND2_X1 U6182 ( .A1(n4463), .A2(n4461), .ZN(n7139) );
  INV_X1 U6183 ( .A(n8845), .ZN(n4464) );
  NAND2_X1 U6184 ( .A1(n4470), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4465) );
  NAND3_X1 U6185 ( .A1(n5137), .A2(n4934), .A3(n4978), .ZN(n4470) );
  NAND3_X1 U6186 ( .A1(n4959), .A2(n4752), .A3(n4755), .ZN(n4471) );
  NOR2_X1 U6187 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(n4468), .ZN(n4467) );
  INV_X1 U6188 ( .A(n4471), .ZN(n4469) );
  AND2_X1 U6189 ( .A1(n4959), .A2(n4755), .ZN(n4754) );
  NOR2_X2 U6190 ( .A1(n4471), .A2(n4470), .ZN(n4992) );
  AND2_X2 U6191 ( .A1(n4934), .A2(n5137), .ZN(n4753) );
  NAND2_X1 U6192 ( .A1(n5795), .A2(n5798), .ZN(n8575) );
  NAND3_X1 U6193 ( .A1(n4362), .A2(n7943), .A3(n4481), .ZN(n4480) );
  NAND2_X1 U6194 ( .A1(n9848), .A2(n4482), .ZN(n7935) );
  NAND2_X2 U6195 ( .A1(n5800), .A2(n5816), .ZN(n5910) );
  NAND2_X2 U6196 ( .A1(n7679), .A2(n5800), .ZN(n7027) );
  NAND2_X2 U6197 ( .A1(n5816), .A2(n5815), .ZN(n6060) );
  NAND3_X1 U6198 ( .A1(n7984), .A2(n7983), .A3(n4486), .ZN(n4489) );
  NAND3_X1 U6199 ( .A1(n4497), .A2(n4495), .A3(n8323), .ZN(n4494) );
  XNOR2_X1 U6200 ( .A(n6301), .B(n8198), .ZN(n8185) );
  NAND2_X1 U6201 ( .A1(n6641), .A2(n4351), .ZN(n4517) );
  OAI21_X1 U6202 ( .B1(n6282), .B2(n6283), .A(n4508), .ZN(n4511) );
  INV_X1 U6203 ( .A(n4509), .ZN(n4508) );
  OAI21_X1 U6204 ( .B1(n6283), .B2(n4519), .A(n6585), .ZN(n4509) );
  NAND2_X1 U6205 ( .A1(n4517), .A2(n4514), .ZN(n4513) );
  INV_X1 U6206 ( .A(n6585), .ZN(n4514) );
  INV_X1 U6207 ( .A(n6843), .ZN(n4519) );
  MUX2_X1 U6208 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n5843), .S(n6588), .Z(n9806)
         );
  NAND2_X1 U6209 ( .A1(n6652), .A2(n6279), .ZN(n9805) );
  NAND3_X1 U6210 ( .A1(n4522), .A2(n4420), .A3(n4521), .ZN(n6292) );
  NAND3_X1 U6211 ( .A1(n4789), .A2(n4787), .A3(n6304), .ZN(n4525) );
  NAND2_X1 U6212 ( .A1(n4545), .A2(n9158), .ZN(n4535) );
  NAND3_X1 U6213 ( .A1(n4530), .A2(n4529), .A3(n4526), .ZN(n9392) );
  INV_X1 U6214 ( .A(n9321), .ZN(n4539) );
  NAND3_X1 U6215 ( .A1(n4353), .A2(n4909), .A3(n4544), .ZN(n4542) );
  INV_X1 U6216 ( .A(n4545), .ZN(n9208) );
  NAND3_X1 U6217 ( .A1(n4354), .A2(n4549), .A3(n4551), .ZN(n4547) );
  NAND2_X1 U6218 ( .A1(n9749), .A2(n9040), .ZN(n8804) );
  NAND2_X1 U6219 ( .A1(n7490), .A2(n4555), .ZN(n4558) );
  NAND2_X1 U6220 ( .A1(n4571), .A2(n9755), .ZN(n7050) );
  AND2_X1 U6221 ( .A1(n9749), .A2(n9739), .ZN(n4572) );
  INV_X1 U6222 ( .A(n7039), .ZN(n4573) );
  NAND2_X1 U6223 ( .A1(n7214), .A2(n4388), .ZN(n7566) );
  NAND3_X1 U6224 ( .A1(n4754), .A2(n4753), .A3(n4965), .ZN(n4584) );
  NAND2_X1 U6225 ( .A1(n4585), .A2(n4312), .ZN(n4587) );
  NAND2_X2 U6226 ( .A1(n4985), .A2(n4586), .ZN(n8794) );
  OAI21_X2 U6227 ( .B1(n4985), .B2(n6726), .A(n4587), .ZN(n6692) );
  NAND2_X1 U6228 ( .A1(n4588), .A2(n5058), .ZN(n5062) );
  XNOR2_X1 U6229 ( .A(n4588), .B(n5058), .ZN(n6589) );
  NAND2_X1 U6230 ( .A1(n5038), .A2(n5037), .ZN(n4588) );
  NAND2_X1 U6231 ( .A1(n5278), .A2(n4596), .ZN(n4593) );
  NAND2_X1 U6232 ( .A1(n4593), .A2(n4594), .ZN(n5355) );
  NAND3_X1 U6233 ( .A1(n4606), .A2(P1_DATAO_REG_1__SCAN_IN), .A3(n4605), .ZN(
        n4610) );
  NAND3_X1 U6234 ( .A1(n4608), .A2(n4609), .A3(n4607), .ZN(n4606) );
  INV_X1 U6235 ( .A(n5200), .ZN(n4615) );
  NAND2_X1 U6236 ( .A1(n4623), .A2(n9151), .ZN(n4622) );
  INV_X1 U6237 ( .A(n8907), .ZN(n4621) );
  OAI21_X1 U6238 ( .B1(n5376), .B2(n5375), .A(n5378), .ZN(n5406) );
  AOI21_X1 U6239 ( .B1(n5376), .B2(n4627), .A(n4626), .ZN(n5447) );
  NAND2_X1 U6240 ( .A1(n6941), .A2(n6978), .ZN(n5866) );
  NAND2_X1 U6241 ( .A1(n5855), .A2(n7907), .ZN(n6941) );
  OAI21_X1 U6242 ( .B1(n7109), .B2(n4352), .A(n4634), .ZN(n4636) );
  NAND2_X1 U6243 ( .A1(n4650), .A2(n4649), .ZN(n7657) );
  NAND2_X1 U6244 ( .A1(n7461), .A2(n4653), .ZN(n4650) );
  OAI21_X1 U6245 ( .B1(n4658), .B2(n8372), .A(n4656), .ZN(n4655) );
  OR2_X1 U6246 ( .A1(n8300), .A2(n6105), .ZN(n4671) );
  OR2_X1 U6247 ( .A1(n8300), .A2(n4675), .ZN(n4674) );
  OAI22_X1 U6248 ( .A1(n8310), .A2(n8313), .B1(n8112), .B2(n7841), .ZN(n8300)
         );
  NAND2_X1 U6249 ( .A1(n5834), .A2(n6460), .ZN(n7938) );
  XNOR2_X1 U6250 ( .A(n6171), .B(n8079), .ZN(n6216) );
  NAND2_X1 U6251 ( .A1(n5949), .A2(n5948), .ZN(n7461) );
  NAND2_X1 U6252 ( .A1(n5866), .A2(n7906), .ZN(n6977) );
  AOI22_X1 U6253 ( .A1(n6262), .A2(n6157), .B1(n7782), .B2(n8106), .ZN(n6171)
         );
  NAND2_X1 U6254 ( .A1(n8333), .A2(n8337), .ZN(n8332) );
  NAND2_X1 U6255 ( .A1(n7370), .A2(n5933), .ZN(n7425) );
  NAND2_X1 U6256 ( .A1(n5503), .A2(n5502), .ZN(n5523) );
  NAND2_X1 U6257 ( .A1(n5451), .A2(n5436), .ZN(n5481) );
  NAND2_X1 U6258 ( .A1(n5447), .A2(n5435), .ZN(n5451) );
  NAND3_X1 U6259 ( .A1(n6191), .A2(n7421), .A3(n7916), .ZN(n4690) );
  NAND2_X1 U6260 ( .A1(n4690), .A2(n4691), .ZN(n7636) );
  OAI21_X1 U6261 ( .B1(n8362), .B2(n4700), .A(n8024), .ZN(n4699) );
  NOR2_X1 U6262 ( .A1(n8362), .A2(n4707), .ZN(n4706) );
  OAI21_X1 U6263 ( .B1(n8362), .B2(n4698), .A(n4697), .ZN(n4696) );
  NAND2_X1 U6264 ( .A1(n4701), .A2(n4705), .ZN(n8350) );
  NAND2_X1 U6265 ( .A1(n8369), .A2(n4706), .ZN(n4701) );
  NAND2_X1 U6266 ( .A1(n4705), .A2(n8023), .ZN(n4704) );
  AOI21_X1 U6267 ( .B1(n6216), .B2(n4709), .A(n4418), .ZN(n4710) );
  NAND2_X1 U6268 ( .A1(n6216), .A2(n8436), .ZN(n4712) );
  NAND2_X1 U6269 ( .A1(n4711), .A2(n4712), .ZN(n6439) );
  OAI21_X1 U6270 ( .B1(n4711), .B2(n9906), .A(n4710), .ZN(P2_U3456) );
  INV_X1 U6271 ( .A(n6215), .ZN(n4713) );
  NAND2_X1 U6272 ( .A1(n6441), .A2(n8064), .ZN(n4719) );
  NAND2_X1 U6273 ( .A1(n8304), .A2(n4724), .ZN(n4721) );
  NAND2_X1 U6274 ( .A1(n4982), .A2(n4732), .ZN(n4731) );
  INV_X4 U6275 ( .A(n4982), .ZN(n6574) );
  OAI21_X1 U6276 ( .B1(n4982), .B2(P2_DATAO_REG_2__SCAN_IN), .A(n4731), .ZN(
        n5059) );
  NAND2_X1 U6277 ( .A1(n8769), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4739) );
  MUX2_X1 U6278 ( .A(n8583), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  MUX2_X1 U6279 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8583), .S(n5829), .Z(n9848) );
  NOR2_X1 U6280 ( .A1(n6315), .A2(n6316), .ZN(n4741) );
  NAND3_X1 U6281 ( .A1(n6846), .A2(n4744), .A3(P2_REG2_REG_3__SCAN_IN), .ZN(
        n6848) );
  NOR2_X1 U6282 ( .A1(n6316), .A2(n6315), .ZN(n6643) );
  NAND2_X1 U6283 ( .A1(n4747), .A2(n4748), .ZN(n7490) );
  INV_X1 U6284 ( .A(n4767), .ZN(n8190) );
  INV_X1 U6285 ( .A(n6332), .ZN(n4766) );
  NAND2_X1 U6286 ( .A1(n8239), .A2(n4771), .ZN(n4770) );
  OAI211_X1 U6287 ( .C1(n8239), .C2(n4772), .A(n4770), .B(n4778), .ZN(P2_U3201) );
  OR2_X2 U6288 ( .A1(n8155), .A2(n4783), .ZN(n4780) );
  INV_X1 U6289 ( .A(n4785), .ZN(n8154) );
  INV_X1 U6290 ( .A(n6329), .ZN(n4784) );
  NOR2_X1 U6291 ( .A1(n8151), .A2(n8506), .ZN(n8150) );
  INV_X1 U6292 ( .A(n4791), .ZN(n8219) );
  INV_X1 U6293 ( .A(n6303), .ZN(n4790) );
  INV_X1 U6294 ( .A(n4795), .ZN(n8184) );
  NAND3_X1 U6295 ( .A1(n6276), .A2(n4905), .A3(P2_IR_REG_2__SCAN_IN), .ZN(
        n4800) );
  NAND2_X1 U6296 ( .A1(n9222), .A2(n4395), .ZN(n4802) );
  NAND2_X1 U6297 ( .A1(n9222), .A2(n4811), .ZN(n4808) );
  OAI211_X1 U6298 ( .C1(n9222), .C2(n4807), .A(n4803), .B(n4802), .ZN(n9196)
         );
  INV_X1 U6299 ( .A(n9262), .ZN(n4824) );
  NAND2_X1 U6300 ( .A1(n5154), .A2(n4828), .ZN(n4826) );
  NAND2_X1 U6301 ( .A1(n5154), .A2(n5153), .ZN(n4827) );
  NAND2_X1 U6302 ( .A1(n4836), .A2(n7485), .ZN(n7558) );
  NOR2_X1 U6303 ( .A1(n9296), .A2(n4838), .ZN(n4837) );
  INV_X1 U6304 ( .A(n9151), .ZN(n4838) );
  NAND3_X1 U6305 ( .A1(n8810), .A2(n7142), .A3(n8808), .ZN(n7205) );
  INV_X1 U6306 ( .A(n8720), .ZN(n4842) );
  AOI21_X2 U6307 ( .B1(n8720), .B2(n4845), .A(n4844), .ZN(n4841) );
  INV_X1 U6308 ( .A(n8605), .ZN(n4845) );
  NAND2_X1 U6309 ( .A1(n8614), .A2(n4327), .ZN(n4846) );
  OAI21_X1 U6310 ( .B1(n8616), .B2(n5475), .A(n5474), .ZN(n8689) );
  AOI21_X1 U6311 ( .B1(n5474), .B2(n5475), .A(n4384), .ZN(n4854) );
  NAND2_X1 U6312 ( .A1(n4862), .A2(n7260), .ZN(n4861) );
  AND2_X1 U6313 ( .A1(n4862), .A2(n4863), .ZN(n7259) );
  AND4_X2 U6314 ( .A1(n4987), .A2(n4929), .A3(n4864), .A4(n4928), .ZN(n5137)
         );
  NAND3_X1 U6315 ( .A1(n4987), .A2(n4929), .A3(n4928), .ZN(n5113) );
  INV_X1 U6316 ( .A(n4942), .ZN(n4944) );
  NOR2_X1 U6317 ( .A1(n5358), .A2(n4866), .ZN(n4940) );
  NAND2_X1 U6318 ( .A1(n8682), .A2(n4870), .ZN(n4867) );
  NAND2_X1 U6319 ( .A1(n8682), .A2(n4877), .ZN(n4875) );
  NAND2_X1 U6320 ( .A1(n7935), .A2(n6464), .ZN(n6672) );
  NAND2_X1 U6321 ( .A1(n7436), .A2(n4886), .ZN(n4882) );
  NAND2_X1 U6322 ( .A1(n4882), .A2(n4883), .ZN(n7536) );
  INV_X1 U6323 ( .A(n7523), .ZN(n4887) );
  NAND2_X1 U6324 ( .A1(n6514), .A2(n4889), .ZN(n7815) );
  NAND2_X1 U6325 ( .A1(n7815), .A2(n7851), .ZN(n6518) );
  NAND2_X1 U6326 ( .A1(n7625), .A2(n4393), .ZN(n7648) );
  AND2_X1 U6327 ( .A1(n4895), .A2(n5768), .ZN(n5780) );
  NAND4_X1 U6328 ( .A1(n5762), .A2(n4906), .A3(n6276), .A4(n4905), .ZN(n5860)
         );
  AND2_X1 U6329 ( .A1(n7421), .A2(n7420), .ZN(n7464) );
  OAI21_X1 U6330 ( .B1(n4398), .B2(n4949), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n4977) );
  NAND2_X1 U6331 ( .A1(n7899), .A2(n7898), .ZN(n8095) );
  INV_X1 U6332 ( .A(n7139), .ZN(n7141) );
  INV_X1 U6333 ( .A(n9275), .ZN(n9276) );
  NAND2_X1 U6334 ( .A1(n5732), .A2(n7703), .ZN(n6690) );
  NAND2_X1 U6335 ( .A1(n9815), .A2(n9814), .ZN(n9813) );
  INV_X1 U6336 ( .A(n6685), .ZN(n8960) );
  AOI21_X1 U6337 ( .B1(n7883), .B2(n7901), .A(n8072), .ZN(n7897) );
  OAI21_X1 U6338 ( .B1(n9206), .B2(n9161), .A(n9160), .ZN(n9162) );
  XNOR2_X2 U6339 ( .A(n6226), .B(n6225), .ZN(n7477) );
  OAI21_X2 U6340 ( .B1(n8709), .B2(n8713), .A(n8597), .ZN(n8682) );
  OAI21_X1 U6341 ( .B1(n8954), .B2(n7136), .A(n8865), .ZN(n8953) );
  INV_X1 U6342 ( .A(n8953), .ZN(n7140) );
  NOR2_X1 U6343 ( .A1(n7027), .A2(n6359), .ZN(n4907) );
  INV_X1 U6344 ( .A(n5596), .ZN(n5622) );
  INV_X1 U6345 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4949) );
  INV_X1 U6346 ( .A(n5867), .ZN(n5865) );
  AND2_X1 U6347 ( .A1(n9479), .A2(n9175), .ZN(n4908) );
  AND2_X1 U6348 ( .A1(n9138), .A2(n9180), .ZN(n4911) );
  AND2_X1 U6349 ( .A1(n7753), .A2(n4402), .ZN(n4912) );
  OR2_X1 U6350 ( .A1(n8266), .A2(n8508), .ZN(n4913) );
  OR2_X1 U6351 ( .A1(n8266), .A2(n8570), .ZN(n4914) );
  OR2_X1 U6352 ( .A1(n9216), .A2(n8760), .ZN(n4915) );
  XNOR2_X1 U6353 ( .A(n7753), .B(n4402), .ZN(n7868) );
  AND2_X1 U6354 ( .A1(n9216), .A2(n9198), .ZN(n4916) );
  AND2_X1 U6355 ( .A1(n4975), .A2(n4974), .ZN(n4917) );
  AND2_X1 U6356 ( .A1(n9906), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4918) );
  AND4_X1 U6357 ( .A1(n5701), .A2(n5700), .A3(n5699), .A4(n5698), .ZN(n9408)
         );
  INV_X1 U6358 ( .A(n9408), .ZN(n9166) );
  AND2_X1 U6359 ( .A1(n6688), .A2(n6689), .ZN(n9762) );
  INV_X1 U6360 ( .A(n9762), .ZN(n9781) );
  OR2_X1 U6361 ( .A1(n6687), .A2(n5740), .ZN(n9532) );
  NOR2_X1 U6362 ( .A1(n5263), .A2(n5234), .ZN(n4919) );
  NOR2_X1 U6363 ( .A1(n7724), .A2(n8570), .ZN(n6440) );
  AND2_X1 U6364 ( .A1(n5228), .A2(n5205), .ZN(n4920) );
  OR2_X1 U6365 ( .A1(n5829), .A2(n6364), .ZN(n4921) );
  NOR2_X1 U6366 ( .A1(n7724), .A2(n8508), .ZN(n6256) );
  AND3_X1 U6367 ( .A1(n6086), .A2(n6085), .A3(n6084), .ZN(n8336) );
  INV_X1 U6368 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6307) );
  NAND2_X1 U6369 ( .A1(n7016), .A2(n9733), .ZN(n9366) );
  INV_X1 U6370 ( .A(n9789), .ZN(n9787) );
  AND2_X1 U6371 ( .A1(n8440), .A2(n9893), .ZN(n9877) );
  INV_X1 U6372 ( .A(n9877), .ZN(n6266) );
  OR2_X1 U6373 ( .A1(n6421), .A2(n8100), .ZN(n9893) );
  AND4_X1 U6374 ( .A1(n5367), .A2(n5366), .A3(n5365), .A4(n5364), .ZN(n9507)
         );
  INV_X1 U6375 ( .A(n6217), .ZN(n6218) );
  OR2_X1 U6376 ( .A1(n9170), .A2(n9507), .ZN(n4922) );
  OR2_X1 U6377 ( .A1(n8124), .A2(n7078), .ZN(n4923) );
  OR2_X1 U6378 ( .A1(n8075), .A2(n8074), .ZN(n4924) );
  OR2_X1 U6379 ( .A1(n8076), .A2(n8570), .ZN(n4925) );
  OR2_X1 U6380 ( .A1(n8076), .A2(n8508), .ZN(n4926) );
  AND2_X1 U6381 ( .A1(n8657), .A2(n5395), .ZN(n4927) );
  MUX2_X1 U6382 ( .A(n7935), .B(n7934), .S(n7933), .Z(n7942) );
  INV_X1 U6383 ( .A(n8056), .ZN(n8057) );
  NOR2_X1 U6384 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  NAND2_X1 U6385 ( .A1(n8060), .A2(n8059), .ZN(n8069) );
  INV_X1 U6386 ( .A(n8073), .ZN(n8080) );
  INV_X1 U6387 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5763) );
  AND2_X1 U6388 ( .A1(n6990), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6285) );
  INV_X1 U6389 ( .A(n8336), .ZN(n6087) );
  INV_X1 U6390 ( .A(n9476), .ZN(n9177) );
  NOR2_X1 U6391 ( .A1(n7738), .A2(n6087), .ZN(n6088) );
  INV_X1 U6392 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5775) );
  OAI22_X1 U6393 ( .A1(n5079), .A2(n9749), .B1(n6631), .B2(n4321), .ZN(n5044)
         );
  OR2_X1 U6394 ( .A1(n7751), .A2(n8109), .ZN(n7752) );
  AND2_X1 U6395 ( .A1(n6856), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6283) );
  AND2_X1 U6396 ( .A1(n7231), .A2(n8100), .ZN(n6232) );
  INV_X1 U6397 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5762) );
  INV_X1 U6398 ( .A(n5196), .ZN(n5194) );
  INV_X1 U6399 ( .A(n6630), .ZN(n5026) );
  OR2_X1 U6400 ( .A1(n5185), .A2(n5184), .ZN(n5213) );
  AND2_X1 U6401 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  INV_X1 U6402 ( .A(n5350), .ZN(n5352) );
  INV_X1 U6403 ( .A(n7437), .ZN(n6498) );
  INV_X1 U6404 ( .A(n6963), .ZN(n6476) );
  INV_X1 U6405 ( .A(n7222), .ZN(n6480) );
  NAND2_X1 U6406 ( .A1(n6588), .A2(n6307), .ZN(n6306) );
  INV_X1 U6407 ( .A(n6298), .ZN(n6297) );
  INV_X1 U6408 ( .A(n8296), .ZN(n8290) );
  INV_X1 U6409 ( .A(n5535), .ZN(n5536) );
  NOR2_X1 U6410 ( .A1(n9164), .A2(n9163), .ZN(n9165) );
  INV_X1 U6411 ( .A(n9415), .ZN(n9227) );
  OR2_X1 U6412 ( .A1(n9526), .A2(n9030), .ZN(n7405) );
  OR2_X1 U6413 ( .A1(n7129), .A2(n8858), .ZN(n7178) );
  OR2_X1 U6414 ( .A1(n5581), .A2(n5580), .ZN(n5612) );
  NOR2_X1 U6415 ( .A1(n5352), .A2(n5351), .ZN(n5354) );
  NAND2_X1 U6416 ( .A1(n5256), .A2(n5255), .ZN(n5276) );
  INV_X1 U6417 ( .A(n5910), .ZN(n6164) );
  INV_X1 U6418 ( .A(n8239), .ZN(n8243) );
  XNOR2_X1 U6419 ( .A(n6443), .B(n6442), .ZN(n6447) );
  INV_X1 U6420 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6257) );
  AND3_X1 U6421 ( .A1(n6537), .A2(n8573), .A3(n6541), .ZN(n6831) );
  NAND2_X1 U6422 ( .A1(n6267), .A2(n6266), .ZN(n6268) );
  AND2_X1 U6423 ( .A1(n6551), .A2(n8085), .ZN(n8430) );
  INV_X1 U6424 ( .A(n8436), .ZN(n9845) );
  AND2_X1 U6425 ( .A1(n5560), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5590) );
  AND2_X1 U6426 ( .A1(n5662), .A2(n5661), .ZN(n6431) );
  OR2_X1 U6427 ( .A1(n5285), .A2(n5284), .ZN(n5311) );
  OR2_X1 U6428 ( .A1(n5384), .A2(n5383), .ZN(n5412) );
  AND2_X1 U6429 ( .A1(n5590), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5623) );
  OR2_X1 U6430 ( .A1(n5751), .A2(n6632), .ZN(n5742) );
  AND2_X1 U6431 ( .A1(n5484), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5507) );
  AND2_X1 U6432 ( .A1(n9600), .A2(n9601), .ZN(n9602) );
  OR2_X1 U6433 ( .A1(n9618), .A2(n9614), .ZN(n9706) );
  INV_X1 U6434 ( .A(n9487), .ZN(n9357) );
  OR2_X1 U6435 ( .A1(n8953), .A2(n7138), .ZN(n8808) );
  INV_X1 U6436 ( .A(n9761), .ZN(n7084) );
  INV_X1 U6437 ( .A(n6766), .ZN(n9739) );
  INV_X1 U6438 ( .A(n5452), .ZN(n8792) );
  AND2_X1 U6439 ( .A1(n5639), .A2(n5618), .ZN(n5636) );
  OR2_X1 U6440 ( .A1(n6552), .A2(n6534), .ZN(n7874) );
  INV_X1 U6441 ( .A(n7860), .ZN(n7870) );
  AND2_X1 U6442 ( .A1(n6550), .A2(n6549), .ZN(n7861) );
  AND2_X1 U6443 ( .A1(n6156), .A2(n6155), .ZN(n8077) );
  AND4_X1 U6444 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n8391)
         );
  INV_X1 U6445 ( .A(n8255), .ZN(n9840) );
  INV_X1 U6446 ( .A(n8246), .ZN(n9830) );
  NAND2_X1 U6447 ( .A1(n8573), .A2(n6530), .ZN(n8427) );
  AND2_X1 U6448 ( .A1(n8422), .A2(n7964), .ZN(n7908) );
  INV_X1 U6449 ( .A(n8429), .ZN(n8382) );
  NOR2_X1 U6450 ( .A1(n9920), .A2(n6257), .ZN(n6258) );
  AND2_X1 U6451 ( .A1(n6540), .A2(n6831), .ZN(n6253) );
  NAND2_X1 U6452 ( .A1(n7932), .A2(n7347), .ZN(n9894) );
  INV_X1 U6453 ( .A(n9894), .ZN(n9900) );
  NAND2_X1 U6454 ( .A1(n5102), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5124) );
  INV_X1 U6455 ( .A(n8760), .ZN(n8741) );
  NAND2_X1 U6456 ( .A1(n5738), .A2(n9009), .ZN(n9733) );
  AND4_X1 U6457 ( .A1(n5595), .A2(n5594), .A3(n5593), .A4(n5592), .ZN(n9438)
         );
  AND4_X1 U6458 ( .A1(n5389), .A2(n5388), .A3(n5387), .A4(n5386), .ZN(n9499)
         );
  INV_X1 U6459 ( .A(n9711), .ZN(n9692) );
  INV_X1 U6460 ( .A(n9706), .ZN(n9696) );
  NAND2_X1 U6461 ( .A1(n9156), .A2(n8921), .ZN(n9251) );
  INV_X1 U6462 ( .A(n9289), .ZN(n9290) );
  INV_X1 U6463 ( .A(n9735), .ZN(n9724) );
  INV_X1 U6464 ( .A(n9532), .ZN(n9474) );
  INV_X1 U6465 ( .A(n9738), .ZN(n9349) );
  INV_X1 U6466 ( .A(n9475), .ZN(n9530) );
  AND2_X1 U6467 ( .A1(n8946), .A2(n9017), .ZN(n9523) );
  INV_X1 U6468 ( .A(n9786), .ZN(n9766) );
  AND3_X1 U6469 ( .A1(n6683), .A2(n6682), .A3(n7008), .ZN(n6778) );
  NAND2_X1 U6470 ( .A1(n7083), .A2(n9769), .ZN(n9786) );
  AND2_X1 U6471 ( .A1(n5259), .A2(n5231), .ZN(n9583) );
  XNOR2_X1 U6472 ( .A(n5132), .B(SI_5_), .ZN(n5130) );
  INV_X1 U6473 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9993) );
  AND2_X1 U6474 ( .A1(n6526), .A2(n6525), .ZN(n7879) );
  AND2_X1 U6475 ( .A1(n7030), .A2(n7029), .ZN(n8093) );
  OR2_X1 U6476 ( .A1(n6542), .A2(n6273), .ZN(n8248) );
  INV_X1 U6477 ( .A(n9816), .ZN(n9832) );
  AND2_X1 U6478 ( .A1(n6834), .A2(n8427), .ZN(n8441) );
  OR2_X1 U6479 ( .A1(n8441), .A2(n6976), .ZN(n8386) );
  NOR2_X1 U6480 ( .A1(n6256), .A2(n6258), .ZN(n6259) );
  NAND2_X1 U6481 ( .A1(n9920), .A2(n9900), .ZN(n8508) );
  INV_X1 U6482 ( .A(n9920), .ZN(n9918) );
  OR2_X1 U6483 ( .A1(n9906), .A2(n9894), .ZN(n8570) );
  AND2_X1 U6484 ( .A1(n6425), .A2(n6424), .ZN(n9906) );
  AND2_X1 U6485 ( .A1(n6542), .A2(n6601), .ZN(n8573) );
  INV_X1 U6486 ( .A(n6418), .ZN(n8090) );
  INV_X1 U6487 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6651) );
  AND2_X1 U6488 ( .A1(n6602), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6453) );
  AND2_X1 U6489 ( .A1(n5739), .A2(n9733), .ZN(n8760) );
  INV_X1 U6490 ( .A(n8748), .ZN(n8766) );
  OR2_X1 U6491 ( .A1(n9618), .A2(n6732), .ZN(n9711) );
  INV_X1 U6492 ( .A(n9616), .ZN(n9721) );
  AND3_X1 U6493 ( .A1(n7128), .A2(n7127), .A3(n7126), .ZN(n9777) );
  OR2_X1 U6494 ( .A1(n4322), .A2(n7012), .ZN(n9369) );
  AND2_X1 U6495 ( .A1(n9777), .A2(n9776), .ZN(n9795) );
  INV_X1 U6496 ( .A(n9745), .ZN(n9746) );
  INV_X1 U6497 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6667) );
  INV_X1 U6498 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6573) );
  INV_X1 U6499 ( .A(n8248), .ZN(P2_U3893) );
  NAND2_X1 U6500 ( .A1(n6272), .A2(n6271), .ZN(P2_U3487) );
  NAND4_X1 U6501 ( .A1(n4930), .A2(n5329), .A3(n9982), .A4(n5207), .ZN(n4933)
         );
  NAND4_X1 U6502 ( .A1(n10038), .A2(n5330), .A3(n5206), .A4(n4931), .ZN(n4932)
         );
  INV_X1 U6503 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U6504 ( .A1(n5408), .A2(n4954), .ZN(n4936) );
  NAND2_X1 U6505 ( .A1(n5454), .A2(n5453), .ZN(n5456) );
  INV_X1 U6506 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4938) );
  AND3_X1 U6507 ( .A1(n4954), .A2(n5453), .A3(n4938), .ZN(n4939) );
  NAND2_X1 U6508 ( .A1(n4944), .A2(n4943), .ZN(n4946) );
  INV_X1 U6509 ( .A(n4946), .ZN(n4945) );
  NAND2_X1 U6510 ( .A1(n4945), .A2(n4955), .ZN(n4953) );
  NAND2_X1 U6511 ( .A1(n4946), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4947) );
  NAND2_X1 U6512 ( .A1(n5726), .A2(n5729), .ZN(n4952) );
  NOR2_X1 U6513 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n4956) );
  NAND4_X1 U6514 ( .A1(n4956), .A2(n4955), .A3(n4935), .A4(n4954), .ZN(n4958)
         );
  NAND4_X1 U6515 ( .A1(n5729), .A2(n5726), .A3(n5453), .A4(n4950), .ZN(n4957)
         );
  XNOR2_X1 U6516 ( .A(n4973), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5712) );
  INV_X1 U6517 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4965) );
  INV_X1 U6518 ( .A(n7497), .ZN(n4967) );
  INV_X1 U6519 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4975) );
  INV_X1 U6520 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4978) );
  INV_X1 U6521 ( .A(n4992), .ZN(n4979) );
  AND2_X1 U6522 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4983) );
  NAND2_X1 U6523 ( .A1(n4320), .A2(n4983), .ZN(n5015) );
  AND2_X1 U6524 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6525 ( .A1(n4982), .A2(n4984), .ZN(n5839) );
  NAND2_X1 U6526 ( .A1(n5015), .A2(n5839), .ZN(n5034) );
  XNOR2_X1 U6527 ( .A(n5033), .B(n5034), .ZN(n5831) );
  INV_X1 U6528 ( .A(n5831), .ZN(n6575) );
  NAND2_X1 U6529 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4986) );
  MUX2_X1 U6530 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4986), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n4990) );
  INV_X1 U6531 ( .A(n4988), .ZN(n4989) );
  NAND2_X1 U6532 ( .A1(n4990), .A2(n4989), .ZN(n6726) );
  INV_X1 U6533 ( .A(n6726), .ZN(n9049) );
  NAND2_X1 U6534 ( .A1(n5043), .A2(n6692), .ZN(n5005) );
  INV_X1 U6535 ( .A(n9572), .ZN(n4997) );
  NAND2_X1 U6536 ( .A1(n5562), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5002) );
  INV_X1 U6537 ( .A(n4998), .ZN(n7706) );
  NAND2_X1 U6538 ( .A1(n5072), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4999) );
  NAND2_X1 U6539 ( .A1(n6684), .A2(n5697), .ZN(n5004) );
  NAND2_X1 U6540 ( .A1(n5005), .A2(n5004), .ZN(n5006) );
  XNOR2_X1 U6541 ( .A(n5006), .B(n5705), .ZN(n5008) );
  NAND2_X1 U6542 ( .A1(n5008), .A2(n5007), .ZN(n7692) );
  NAND2_X1 U6543 ( .A1(n4368), .A2(n7692), .ZN(n6629) );
  INV_X1 U6544 ( .A(n6629), .ZN(n5027) );
  NAND2_X1 U6545 ( .A1(n4316), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5012) );
  NAND2_X1 U6546 ( .A1(n5072), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5011) );
  NAND2_X1 U6547 ( .A1(n8769), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5010) );
  NAND2_X1 U6548 ( .A1(n5050), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5009) );
  NAND4_X2 U6549 ( .A1(n5012), .A2(n5011), .A3(n5010), .A4(n5009), .ZN(n9042)
         );
  NAND2_X1 U6550 ( .A1(n9042), .A2(n5697), .ZN(n5018) );
  INV_X1 U6551 ( .A(SI_0_), .ZN(n5014) );
  INV_X1 U6552 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5013) );
  OAI21_X1 U6553 ( .B1(n4586), .B2(n5014), .A(n5013), .ZN(n5016) );
  AND2_X1 U6554 ( .A1(n5016), .A2(n5015), .ZN(n9574) );
  MUX2_X1 U6555 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9574), .S(n4985), .Z(n7688) );
  NAND2_X1 U6556 ( .A1(n5043), .A2(n7688), .ZN(n5017) );
  AND2_X1 U6557 ( .A1(n5018), .A2(n5017), .ZN(n5023) );
  INV_X1 U6558 ( .A(n5019), .ZN(n6454) );
  NAND2_X1 U6559 ( .A1(n6454), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U6560 ( .A1(n5023), .A2(n5020), .ZN(n6708) );
  NAND2_X1 U6561 ( .A1(n9042), .A2(n5654), .ZN(n5022) );
  AOI22_X1 U6562 ( .A1(n5697), .A2(n7688), .B1(n6454), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U6563 ( .A1(n5022), .A2(n5021), .ZN(n6709) );
  NAND2_X1 U6564 ( .A1(n6708), .A2(n6709), .ZN(n5025) );
  NAND2_X1 U6565 ( .A1(n5023), .A2(n5705), .ZN(n5024) );
  NAND2_X1 U6566 ( .A1(n6627), .A2(n7692), .ZN(n5047) );
  NAND2_X1 U6567 ( .A1(n5072), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5028) );
  OR2_X1 U6568 ( .A1(n6631), .A2(n4315), .ZN(n5042) );
  NOR2_X1 U6569 ( .A1(n4988), .A2(n4949), .ZN(n5029) );
  MUX2_X1 U6570 ( .A(n4949), .B(n5029), .S(P1_IR_REG_2__SCAN_IN), .Z(n5030) );
  INV_X1 U6571 ( .A(n5030), .ZN(n5032) );
  NAND2_X1 U6572 ( .A1(n5032), .A2(n5031), .ZN(n6747) );
  XNOR2_X1 U6573 ( .A(n5059), .B(SI_2_), .ZN(n5058) );
  INV_X1 U6574 ( .A(n5033), .ZN(n5035) );
  NAND2_X1 U6575 ( .A1(n5035), .A2(n5034), .ZN(n5038) );
  NAND2_X1 U6576 ( .A1(n5036), .A2(SI_1_), .ZN(n5037) );
  OR2_X1 U6577 ( .A1(n5452), .A2(n6589), .ZN(n5040) );
  NAND2_X1 U6578 ( .A1(n5697), .A2(n7699), .ZN(n5041) );
  INV_X1 U6579 ( .A(n5043), .ZN(n5079) );
  NAND2_X1 U6580 ( .A1(n5045), .A2(n4344), .ZN(n5048) );
  OAI21_X1 U6581 ( .B1(n4344), .B2(n5045), .A(n5048), .ZN(n5046) );
  NAND2_X1 U6582 ( .A1(n5047), .A2(n7694), .ZN(n7695) );
  NAND2_X1 U6583 ( .A1(n7695), .A2(n5048), .ZN(n6758) );
  INV_X1 U6584 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U6585 ( .A1(n4316), .A2(n5049), .ZN(n5054) );
  NAND2_X1 U6586 ( .A1(n5072), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U6587 ( .A1(n8769), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U6588 ( .A1(n5050), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U6589 ( .A1(n5031), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5056) );
  INV_X1 U6590 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5055) );
  NAND2_X1 U6591 ( .A1(n5056), .A2(n5055), .ZN(n5087) );
  OR2_X1 U6592 ( .A1(n5056), .A2(n5055), .ZN(n5057) );
  NAND2_X1 U6593 ( .A1(n5087), .A2(n5057), .ZN(n9054) );
  INV_X1 U6594 ( .A(n5059), .ZN(n5060) );
  NAND2_X1 U6595 ( .A1(n5060), .A2(SI_2_), .ZN(n5061) );
  NAND2_X1 U6596 ( .A1(n5062), .A2(n5061), .ZN(n5081) );
  MUX2_X1 U6597 ( .A(n6582), .B(n6572), .S(n6574), .Z(n5082) );
  XNOR2_X1 U6598 ( .A(n5081), .B(n5080), .ZN(n6581) );
  OR2_X1 U6599 ( .A1(n5452), .A2(n6581), .ZN(n5064) );
  OR2_X1 U6600 ( .A1(n8794), .A2(n6572), .ZN(n5063) );
  OAI211_X1 U6601 ( .C1(n4312), .C2(n9054), .A(n5064), .B(n5063), .ZN(n6766)
         );
  OAI22_X1 U6602 ( .A1(n6870), .A2(n4321), .B1(n9739), .B2(n5079), .ZN(n5065)
         );
  XNOR2_X1 U6603 ( .A(n5065), .B(n5705), .ZN(n5070) );
  OR2_X1 U6604 ( .A1(n6870), .A2(n4315), .ZN(n5067) );
  NAND2_X1 U6605 ( .A1(n5697), .A2(n6766), .ZN(n5066) );
  NAND2_X1 U6606 ( .A1(n5067), .A2(n5066), .ZN(n5068) );
  XNOR2_X1 U6607 ( .A(n5070), .B(n5068), .ZN(n6759) );
  NAND2_X1 U6608 ( .A1(n6758), .A2(n6759), .ZN(n6757) );
  INV_X1 U6609 ( .A(n5068), .ZN(n5069) );
  NAND2_X1 U6610 ( .A1(n5070), .A2(n5069), .ZN(n5071) );
  NAND2_X1 U6611 ( .A1(n6757), .A2(n5071), .ZN(n6859) );
  NAND2_X1 U6612 ( .A1(n5072), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6613 ( .A1(n5101), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5077) );
  NOR2_X1 U6614 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5073) );
  NOR2_X1 U6615 ( .A1(n5102), .A2(n5073), .ZN(n7052) );
  NAND2_X1 U6616 ( .A1(n4317), .A2(n7052), .ZN(n5076) );
  INV_X4 U6617 ( .A(n5074), .ZN(n8769) );
  NAND2_X1 U6618 ( .A1(n8769), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6619 ( .A1(n9038), .A2(n5697), .ZN(n5093) );
  INV_X1 U6620 ( .A(n5079), .ZN(n5283) );
  NAND2_X1 U6621 ( .A1(n5081), .A2(n5080), .ZN(n5085) );
  INV_X1 U6622 ( .A(n5082), .ZN(n5083) );
  NAND2_X1 U6623 ( .A1(n5083), .A2(SI_3_), .ZN(n5084) );
  MUX2_X1 U6624 ( .A(n6584), .B(n6577), .S(n6574), .Z(n5109) );
  XNOR2_X1 U6625 ( .A(n5108), .B(n5107), .ZN(n6583) );
  OR2_X1 U6626 ( .A1(n5452), .A2(n6583), .ZN(n5091) );
  OR2_X1 U6627 ( .A1(n8794), .A2(n6577), .ZN(n5090) );
  NAND2_X1 U6628 ( .A1(n5087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5088) );
  XNOR2_X1 U6629 ( .A(n5088), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U6630 ( .A1(n5086), .A2(n6804), .ZN(n5089) );
  INV_X1 U6631 ( .A(n9755), .ZN(n7051) );
  NAND2_X1 U6632 ( .A1(n5283), .A2(n7051), .ZN(n5092) );
  NAND2_X1 U6633 ( .A1(n5093), .A2(n5092), .ZN(n5094) );
  XNOR2_X1 U6634 ( .A(n5094), .B(n5705), .ZN(n5096) );
  AOI22_X1 U6635 ( .A1(n9038), .A2(n5654), .B1(n7051), .B2(n5697), .ZN(n5097)
         );
  XNOR2_X1 U6636 ( .A(n5096), .B(n5097), .ZN(n6860) );
  INV_X1 U6637 ( .A(n5096), .ZN(n5099) );
  INV_X1 U6638 ( .A(n5097), .ZN(n5098) );
  NAND2_X1 U6639 ( .A1(n5099), .A2(n5098), .ZN(n5100) );
  NAND2_X1 U6640 ( .A1(n5101), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U6641 ( .A1(n5072), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5105) );
  OAI21_X1 U6642 ( .B1(n5102), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5124), .ZN(
        n6921) );
  INV_X1 U6643 ( .A(n6921), .ZN(n9723) );
  NAND2_X1 U6644 ( .A1(n4316), .A2(n9723), .ZN(n5104) );
  NAND2_X1 U6645 ( .A1(n8769), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U6646 ( .A1(n5108), .A2(n5107), .ZN(n5112) );
  INV_X1 U6647 ( .A(n5109), .ZN(n5110) );
  NAND2_X1 U6648 ( .A1(n5110), .A2(SI_4_), .ZN(n5111) );
  NAND2_X1 U6649 ( .A1(n5112), .A2(n5111), .ZN(n5131) );
  MUX2_X1 U6650 ( .A(n6587), .B(n6579), .S(n6574), .Z(n5132) );
  XNOR2_X1 U6651 ( .A(n5131), .B(n5130), .ZN(n6586) );
  OR2_X1 U6652 ( .A1(n6586), .A2(n5452), .ZN(n5116) );
  NAND2_X1 U6653 ( .A1(n5113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5114) );
  XNOR2_X1 U6654 ( .A(n5114), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U6655 ( .A1(n5086), .A2(n9075), .ZN(n5115) );
  OAI211_X1 U6656 ( .C1(n8794), .C2(n6579), .A(n5116), .B(n5115), .ZN(n6883)
         );
  INV_X1 U6657 ( .A(n6883), .ZN(n9728) );
  INV_X1 U6658 ( .A(n5283), .ZN(n5596) );
  OAI22_X1 U6659 ( .A1(n7046), .A2(n4321), .B1(n9728), .B2(n5596), .ZN(n5117)
         );
  XNOR2_X1 U6660 ( .A(n5117), .B(n4324), .ZN(n6914) );
  INV_X1 U6661 ( .A(n6914), .ZN(n5121) );
  OR2_X1 U6662 ( .A1(n7046), .A2(n4315), .ZN(n5119) );
  NAND2_X1 U6663 ( .A1(n5697), .A2(n6883), .ZN(n5118) );
  NAND2_X1 U6664 ( .A1(n5119), .A2(n5118), .ZN(n6913) );
  INV_X1 U6665 ( .A(n6913), .ZN(n5120) );
  NAND2_X1 U6666 ( .A1(n5121), .A2(n5120), .ZN(n5122) );
  NAND2_X1 U6667 ( .A1(n5101), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6668 ( .A1(n5072), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5128) );
  NOR2_X2 U6669 ( .A1(n5124), .A2(n5123), .ZN(n5147) );
  AND2_X1 U6670 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  NOR2_X1 U6671 ( .A1(n5147), .A2(n5125), .ZN(n7018) );
  NAND2_X1 U6672 ( .A1(n4316), .A2(n7018), .ZN(n5127) );
  NAND2_X1 U6673 ( .A1(n8769), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U6674 ( .A1(n5131), .A2(n5130), .ZN(n5135) );
  INV_X1 U6675 ( .A(n5132), .ZN(n5133) );
  NAND2_X1 U6676 ( .A1(n5133), .A2(SI_5_), .ZN(n5134) );
  INV_X1 U6677 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5136) );
  MUX2_X1 U6678 ( .A(n9991), .B(n5136), .S(n6574), .Z(n5155) );
  XNOR2_X1 U6679 ( .A(n5154), .B(n5153), .ZN(n6591) );
  OR2_X1 U6680 ( .A1(n6591), .A2(n5452), .ZN(n5142) );
  NOR2_X1 U6681 ( .A1(n5137), .A2(n4949), .ZN(n5138) );
  MUX2_X1 U6682 ( .A(n4949), .B(n5138), .S(P1_IR_REG_6__SCAN_IN), .Z(n5140) );
  INV_X1 U6683 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U6684 ( .A1(n5137), .A2(n10069), .ZN(n5209) );
  INV_X1 U6685 ( .A(n5209), .ZN(n5139) );
  AOI22_X1 U6686 ( .A1(n5457), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5086), .B2(
        n9089), .ZN(n5141) );
  NAND2_X1 U6687 ( .A1(n5142), .A2(n5141), .ZN(n9761) );
  OAI22_X1 U6688 ( .A1(n7088), .A2(n4321), .B1(n7084), .B2(n5596), .ZN(n5143)
         );
  XNOR2_X1 U6689 ( .A(n5143), .B(n4324), .ZN(n5145) );
  OAI22_X1 U6690 ( .A1(n7088), .A2(n4315), .B1(n7084), .B2(n4321), .ZN(n5144)
         );
  NAND2_X1 U6691 ( .A1(n5145), .A2(n5144), .ZN(n6903) );
  NAND2_X1 U6692 ( .A1(n6902), .A2(n6903), .ZN(n5146) );
  OR2_X1 U6693 ( .A1(n5145), .A2(n5144), .ZN(n6904) );
  NAND2_X1 U6694 ( .A1(n5146), .A2(n6904), .ZN(n6952) );
  NAND2_X1 U6695 ( .A1(n5072), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5152) );
  NAND2_X1 U6696 ( .A1(n5101), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5151) );
  NAND2_X1 U6697 ( .A1(n5147), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5185) );
  OR2_X1 U6698 ( .A1(n5147), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5148) );
  AND2_X1 U6699 ( .A1(n5185), .A2(n5148), .ZN(n7098) );
  NAND2_X1 U6700 ( .A1(n4317), .A2(n7098), .ZN(n5150) );
  NAND2_X1 U6701 ( .A1(n8769), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5149) );
  OR2_X1 U6702 ( .A1(n8848), .A2(n4323), .ZN(n5164) );
  INV_X1 U6703 ( .A(n5155), .ZN(n5156) );
  NAND2_X1 U6704 ( .A1(n5156), .A2(SI_6_), .ZN(n5157) );
  INV_X1 U6705 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5158) );
  MUX2_X1 U6706 ( .A(n6595), .B(n5158), .S(n6574), .Z(n5173) );
  OR2_X1 U6707 ( .A1(n6594), .A2(n5452), .ZN(n5162) );
  NAND2_X1 U6708 ( .A1(n5209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U6709 ( .A1(n5159), .A2(n5207), .ZN(n5180) );
  OR2_X1 U6710 ( .A1(n5159), .A2(n5207), .ZN(n5160) );
  AOI22_X1 U6711 ( .A1(n5457), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5086), .B2(
        n9597), .ZN(n5161) );
  NAND2_X1 U6712 ( .A1(n5162), .A2(n5161), .ZN(n8849) );
  NAND2_X1 U6713 ( .A1(n8849), .A2(n5697), .ZN(n5163) );
  AND2_X1 U6714 ( .A1(n5164), .A2(n5163), .ZN(n6954) );
  NAND2_X1 U6715 ( .A1(n6952), .A2(n6954), .ZN(n5167) );
  NAND2_X1 U6716 ( .A1(n8849), .A2(n5283), .ZN(n5165) );
  OAI21_X1 U6717 ( .B1(n8848), .B2(n4321), .A(n5165), .ZN(n5166) );
  XNOR2_X1 U6718 ( .A(n5166), .B(n4324), .ZN(n6953) );
  NAND2_X1 U6719 ( .A1(n5167), .A2(n6953), .ZN(n5171) );
  INV_X1 U6720 ( .A(n6952), .ZN(n5169) );
  INV_X1 U6721 ( .A(n6954), .ZN(n5168) );
  NAND2_X1 U6722 ( .A1(n5169), .A2(n5168), .ZN(n5170) );
  NAND2_X1 U6723 ( .A1(n5171), .A2(n5170), .ZN(n5197) );
  INV_X1 U6724 ( .A(n5197), .ZN(n5195) );
  INV_X1 U6725 ( .A(n5173), .ZN(n5174) );
  INV_X1 U6726 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5175) );
  MUX2_X1 U6727 ( .A(n6606), .B(n5175), .S(n4320), .Z(n5177) );
  INV_X1 U6728 ( .A(SI_8_), .ZN(n5176) );
  INV_X1 U6729 ( .A(n5177), .ZN(n5178) );
  NAND2_X1 U6730 ( .A1(n5178), .A2(SI_8_), .ZN(n5179) );
  XNOR2_X1 U6731 ( .A(n5200), .B(n5199), .ZN(n6599) );
  NAND2_X1 U6732 ( .A1(n6599), .A2(n8792), .ZN(n5183) );
  NAND2_X1 U6733 ( .A1(n5180), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5181) );
  AOI22_X1 U6734 ( .A1(n5457), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5086), .B2(
        n9609), .ZN(n5182) );
  NAND2_X1 U6735 ( .A1(n5183), .A2(n5182), .ZN(n8858) );
  NAND2_X1 U6736 ( .A1(n8858), .A2(n5283), .ZN(n5192) );
  NAND2_X1 U6737 ( .A1(n5072), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6738 ( .A1(n8769), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5189) );
  NAND2_X1 U6739 ( .A1(n5185), .A2(n5184), .ZN(n5186) );
  AND2_X1 U6740 ( .A1(n5213), .A2(n5186), .ZN(n7261) );
  NAND2_X1 U6741 ( .A1(n4317), .A2(n7261), .ZN(n5188) );
  NAND2_X1 U6742 ( .A1(n5101), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5187) );
  OR2_X1 U6743 ( .A1(n8854), .A2(n4321), .ZN(n5191) );
  NAND2_X1 U6744 ( .A1(n5192), .A2(n5191), .ZN(n5193) );
  XNOR2_X1 U6745 ( .A(n5193), .B(n4324), .ZN(n5196) );
  INV_X1 U6746 ( .A(n8854), .ZN(n9034) );
  AOI22_X1 U6747 ( .A1(n8858), .A2(n5697), .B1(n9034), .B2(n5654), .ZN(n7260)
         );
  INV_X1 U6748 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5201) );
  MUX2_X1 U6749 ( .A(n6610), .B(n5201), .S(n4320), .Z(n5203) );
  INV_X1 U6750 ( .A(SI_9_), .ZN(n5202) );
  INV_X1 U6751 ( .A(n5203), .ZN(n5204) );
  NAND2_X1 U6752 ( .A1(n5204), .A2(SI_9_), .ZN(n5205) );
  NAND2_X1 U6753 ( .A1(n6608), .A2(n8792), .ZN(n5212) );
  NAND2_X1 U6754 ( .A1(n5207), .A2(n5206), .ZN(n5208) );
  NAND2_X1 U6755 ( .A1(n5333), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5210) );
  XNOR2_X1 U6756 ( .A(n5210), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9105) );
  AOI22_X1 U6757 ( .A1(n5457), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5086), .B2(
        n9105), .ZN(n5211) );
  NAND2_X1 U6758 ( .A1(n9779), .A2(n5622), .ZN(n5220) );
  NAND2_X1 U6759 ( .A1(n5072), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5218) );
  NAND2_X1 U6760 ( .A1(n8769), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5217) );
  AND2_X1 U6761 ( .A1(n5213), .A2(n7333), .ZN(n5214) );
  NOR2_X1 U6762 ( .A1(n5233), .A2(n5214), .ZN(n7334) );
  NAND2_X1 U6763 ( .A1(n4316), .A2(n7334), .ZN(n5216) );
  NAND2_X1 U6764 ( .A1(n5101), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5215) );
  OR2_X1 U6765 ( .A1(n7265), .A2(n4321), .ZN(n5219) );
  NAND2_X1 U6766 ( .A1(n5220), .A2(n5219), .ZN(n5221) );
  XNOR2_X1 U6767 ( .A(n5221), .B(n4324), .ZN(n5223) );
  NOR2_X1 U6768 ( .A1(n7265), .A2(n4315), .ZN(n5222) );
  AOI21_X1 U6769 ( .B1(n9779), .B2(n5697), .A(n5222), .ZN(n5224) );
  XNOR2_X1 U6770 ( .A(n5223), .B(n5224), .ZN(n7332) );
  NAND2_X1 U6771 ( .A1(n7330), .A2(n7332), .ZN(n7331) );
  INV_X1 U6772 ( .A(n5223), .ZN(n5225) );
  NAND2_X1 U6773 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  NAND2_X1 U6774 ( .A1(n7331), .A2(n5226), .ZN(n5245) );
  INV_X1 U6775 ( .A(n5245), .ZN(n5243) );
  INV_X1 U6776 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5229) );
  MUX2_X1 U6777 ( .A(n6614), .B(n5229), .S(n6574), .Z(n5251) );
  OAI21_X1 U6778 ( .B1(n5333), .B2(P1_IR_REG_9__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5280) );
  INV_X1 U6779 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6780 ( .A1(n5280), .A2(n5230), .ZN(n5259) );
  OR2_X1 U6781 ( .A1(n5280), .A2(n5230), .ZN(n5231) );
  AOI22_X1 U6782 ( .A1(n5457), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5086), .B2(
        n9583), .ZN(n5232) );
  NAND2_X1 U6783 ( .A1(n7208), .A2(n5283), .ZN(n5240) );
  NAND2_X1 U6784 ( .A1(n5072), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6785 ( .A1(n5101), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5237) );
  NOR2_X1 U6786 ( .A1(n5233), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U6787 ( .A1(n4316), .A2(n4919), .ZN(n5236) );
  NAND2_X1 U6788 ( .A1(n8769), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5235) );
  OR2_X1 U6789 ( .A1(n9533), .A2(n4321), .ZN(n5239) );
  NAND2_X1 U6790 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  XNOR2_X1 U6791 ( .A(n5241), .B(n5705), .ZN(n5244) );
  INV_X1 U6792 ( .A(n5244), .ZN(n5242) );
  NAND2_X1 U6793 ( .A1(n5243), .A2(n5242), .ZN(n5246) );
  NAND2_X2 U6794 ( .A1(n5245), .A2(n5244), .ZN(n8720) );
  NOR2_X1 U6795 ( .A1(n9533), .A2(n4315), .ZN(n5247) );
  AOI21_X1 U6796 ( .B1(n7208), .B2(n5697), .A(n5247), .ZN(n8605) );
  INV_X1 U6797 ( .A(n5251), .ZN(n5252) );
  MUX2_X1 U6798 ( .A(n6624), .B(n6625), .S(n4320), .Z(n5256) );
  INV_X1 U6799 ( .A(SI_11_), .ZN(n5255) );
  INV_X1 U6800 ( .A(n5256), .ZN(n5257) );
  NAND2_X1 U6801 ( .A1(n5257), .A2(SI_11_), .ZN(n5258) );
  XNOR2_X1 U6802 ( .A(n5278), .B(n5277), .ZN(n6623) );
  NAND2_X1 U6803 ( .A1(n6623), .A2(n8792), .ZN(n5262) );
  NAND2_X1 U6804 ( .A1(n5259), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5260) );
  XNOR2_X1 U6805 ( .A(n5260), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6813) );
  AOI22_X1 U6806 ( .A1(n5457), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5086), .B2(
        n6813), .ZN(n5261) );
  NAND2_X1 U6807 ( .A1(n9535), .A2(n5283), .ZN(n5270) );
  NAND2_X1 U6808 ( .A1(n5101), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6809 ( .A1(n5072), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5267) );
  OR2_X1 U6810 ( .A1(n5263), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5264) );
  AND2_X1 U6811 ( .A1(n5285), .A2(n5264), .ZN(n8730) );
  NAND2_X1 U6812 ( .A1(n4317), .A2(n8730), .ZN(n5266) );
  NAND2_X1 U6813 ( .A1(n8769), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5265) );
  OR2_X1 U6814 ( .A1(n8643), .A2(n4321), .ZN(n5269) );
  NAND2_X1 U6815 ( .A1(n5270), .A2(n5269), .ZN(n5271) );
  XNOR2_X1 U6816 ( .A(n5271), .B(n5705), .ZN(n5274) );
  NOR2_X1 U6817 ( .A1(n8643), .A2(n4315), .ZN(n5272) );
  AOI21_X1 U6818 ( .B1(n9535), .B2(n5697), .A(n5272), .ZN(n5273) );
  NAND2_X1 U6819 ( .A1(n5274), .A2(n5273), .ZN(n8635) );
  OR2_X1 U6820 ( .A1(n5274), .A2(n5273), .ZN(n5275) );
  AND2_X1 U6821 ( .A1(n8635), .A2(n5275), .ZN(n8721) );
  NAND2_X1 U6822 ( .A1(n8634), .A2(n8635), .ZN(n5298) );
  MUX2_X1 U6823 ( .A(n6651), .B(n6667), .S(n6574), .Z(n5301) );
  XNOR2_X1 U6824 ( .A(n5305), .B(n5300), .ZN(n6650) );
  NAND2_X1 U6825 ( .A1(n6650), .A2(n8792), .ZN(n5282) );
  OAI21_X1 U6826 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6827 ( .A1(n5280), .A2(n5279), .ZN(n5306) );
  XNOR2_X1 U6828 ( .A(n5306), .B(n5329), .ZN(n9123) );
  AOI22_X1 U6829 ( .A1(n5457), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5086), .B2(
        n9123), .ZN(n5281) );
  NAND2_X1 U6830 ( .A1(n9526), .A2(n5283), .ZN(n5292) );
  NAND2_X1 U6831 ( .A1(n5101), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6832 ( .A1(n5072), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5289) );
  INV_X1 U6833 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U6834 ( .A1(n5285), .A2(n5284), .ZN(n5286) );
  AND2_X1 U6835 ( .A1(n5311), .A2(n5286), .ZN(n8645) );
  NAND2_X1 U6836 ( .A1(n4317), .A2(n8645), .ZN(n5288) );
  NAND2_X1 U6837 ( .A1(n8769), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5287) );
  OR2_X1 U6838 ( .A1(n9531), .A2(n4321), .ZN(n5291) );
  NAND2_X1 U6839 ( .A1(n5292), .A2(n5291), .ZN(n5293) );
  XNOR2_X1 U6840 ( .A(n5293), .B(n5705), .ZN(n5296) );
  NOR2_X1 U6841 ( .A1(n9531), .A2(n4315), .ZN(n5294) );
  AOI21_X1 U6842 ( .B1(n9526), .B2(n5697), .A(n5294), .ZN(n5295) );
  NAND2_X1 U6843 ( .A1(n5296), .A2(n5295), .ZN(n5299) );
  OR2_X1 U6844 ( .A1(n5296), .A2(n5295), .ZN(n5297) );
  AND2_X1 U6845 ( .A1(n5299), .A2(n5297), .ZN(n8636) );
  NAND2_X1 U6846 ( .A1(n5298), .A2(n8636), .ZN(n8638) );
  NAND2_X1 U6847 ( .A1(n8638), .A2(n5299), .ZN(n8699) );
  INV_X1 U6848 ( .A(n5301), .ZN(n5302) );
  NAND2_X1 U6849 ( .A1(n5302), .A2(SI_12_), .ZN(n5303) );
  MUX2_X1 U6850 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6574), .Z(n5327) );
  XNOR2_X1 U6851 ( .A(n5326), .B(n5325), .ZN(n6668) );
  NAND2_X1 U6852 ( .A1(n6668), .A2(n8792), .ZN(n5309) );
  OAI21_X1 U6853 ( .B1(n5306), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5307) );
  XNOR2_X1 U6854 ( .A(n5307), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9644) );
  AOI22_X1 U6855 ( .A1(n5457), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5086), .B2(
        n9644), .ZN(n5308) );
  NAND2_X1 U6856 ( .A1(n9519), .A2(n5622), .ZN(n5318) );
  NAND2_X1 U6857 ( .A1(n5101), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6858 ( .A1(n5072), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5315) );
  INV_X1 U6859 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6860 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  AND2_X1 U6861 ( .A1(n5338), .A2(n5312), .ZN(n8705) );
  NAND2_X1 U6862 ( .A1(n4317), .A2(n8705), .ZN(n5314) );
  NAND2_X1 U6863 ( .A1(n8769), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5313) );
  OR2_X1 U6864 ( .A1(n9508), .A2(n4321), .ZN(n5317) );
  NAND2_X1 U6865 ( .A1(n5318), .A2(n5317), .ZN(n5319) );
  XNOR2_X1 U6866 ( .A(n5319), .B(n4324), .ZN(n5321) );
  NOR2_X1 U6867 ( .A1(n9508), .A2(n4315), .ZN(n5320) );
  AOI21_X1 U6868 ( .B1(n9519), .B2(n5697), .A(n5320), .ZN(n5322) );
  XNOR2_X1 U6869 ( .A(n5321), .B(n5322), .ZN(n8700) );
  NAND2_X1 U6870 ( .A1(n8699), .A2(n8700), .ZN(n8698) );
  INV_X1 U6871 ( .A(n5321), .ZN(n5323) );
  NAND2_X1 U6872 ( .A1(n5323), .A2(n5322), .ZN(n5324) );
  NAND2_X1 U6873 ( .A1(n8698), .A2(n5324), .ZN(n8585) );
  MUX2_X1 U6874 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4320), .Z(n5350) );
  XNOR2_X1 U6875 ( .A(n5350), .B(SI_14_), .ZN(n5328) );
  XNOR2_X1 U6876 ( .A(n5355), .B(n5328), .ZN(n6823) );
  NAND2_X1 U6877 ( .A1(n6823), .A2(n8792), .ZN(n5336) );
  NOR2_X1 U6878 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5331) );
  NAND4_X1 U6879 ( .A1(n5331), .A2(n5330), .A3(n5329), .A4(n9982), .ZN(n5332)
         );
  OAI21_X1 U6880 ( .B1(n5333), .B2(n5332), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5334) );
  XNOR2_X1 U6881 ( .A(n5334), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9124) );
  AOI22_X1 U6882 ( .A1(n5457), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5086), .B2(
        n9124), .ZN(n5335) );
  NAND2_X1 U6883 ( .A1(n9510), .A2(n5622), .ZN(n5345) );
  NAND2_X1 U6884 ( .A1(n5101), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6885 ( .A1(n5072), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5342) );
  INV_X1 U6886 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5337) );
  AND2_X1 U6887 ( .A1(n5338), .A2(n5337), .ZN(n5339) );
  NOR2_X1 U6888 ( .A1(n5362), .A2(n5339), .ZN(n8593) );
  NAND2_X1 U6889 ( .A1(n4316), .A2(n8593), .ZN(n5341) );
  NAND2_X1 U6890 ( .A1(n8769), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5340) );
  OR2_X1 U6891 ( .A1(n9516), .A2(n4321), .ZN(n5344) );
  NAND2_X1 U6892 ( .A1(n5345), .A2(n5344), .ZN(n5346) );
  XNOR2_X1 U6893 ( .A(n5346), .B(n4324), .ZN(n8586) );
  NAND2_X1 U6894 ( .A1(n9510), .A2(n5697), .ZN(n5348) );
  OR2_X1 U6895 ( .A1(n9516), .A2(n4315), .ZN(n5347) );
  NAND2_X1 U6896 ( .A1(n5348), .A2(n5347), .ZN(n8584) );
  NAND2_X1 U6897 ( .A1(n8586), .A2(n8584), .ZN(n5349) );
  NAND2_X1 U6898 ( .A1(n8585), .A2(n5349), .ZN(n5373) );
  INV_X1 U6899 ( .A(SI_14_), .ZN(n5351) );
  NAND2_X1 U6900 ( .A1(n5352), .A2(n5351), .ZN(n5353) );
  INV_X1 U6901 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5356) );
  INV_X1 U6902 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6868) );
  MUX2_X1 U6903 ( .A(n5356), .B(n6868), .S(n6574), .Z(n5374) );
  XNOR2_X1 U6904 ( .A(n5374), .B(SI_15_), .ZN(n5357) );
  XNOR2_X1 U6905 ( .A(n5376), .B(n5357), .ZN(n6866) );
  NAND2_X1 U6906 ( .A1(n6866), .A2(n8792), .ZN(n5361) );
  NAND2_X1 U6907 ( .A1(n5358), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5359) );
  XNOR2_X1 U6908 ( .A(n5359), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9671) );
  AOI22_X1 U6909 ( .A1(n5457), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5086), .B2(
        n9671), .ZN(n5360) );
  NAND2_X1 U6910 ( .A1(n5101), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U6911 ( .A1(n5072), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5366) );
  OR2_X1 U6912 ( .A1(n5362), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6913 ( .A1(n5362), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5384) );
  AND2_X1 U6914 ( .A1(n5363), .A2(n5384), .ZN(n8764) );
  NAND2_X1 U6915 ( .A1(n4316), .A2(n8764), .ZN(n5365) );
  NAND2_X1 U6916 ( .A1(n8769), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5364) );
  OAI22_X1 U6917 ( .A1(n9170), .A2(n5596), .B1(n9507), .B2(n4321), .ZN(n5368)
         );
  XNOR2_X1 U6918 ( .A(n5368), .B(n4324), .ZN(n8661) );
  OR2_X1 U6919 ( .A1(n9170), .A2(n4321), .ZN(n5370) );
  OR2_X1 U6920 ( .A1(n9507), .A2(n5702), .ZN(n5369) );
  NAND2_X1 U6921 ( .A1(n5370), .A2(n5369), .ZN(n8756) );
  OAI22_X1 U6922 ( .A1(n8661), .A2(n8756), .B1(n8584), .B2(n8586), .ZN(n5371)
         );
  INV_X1 U6923 ( .A(n5371), .ZN(n5372) );
  NAND2_X1 U6924 ( .A1(n5373), .A2(n5372), .ZN(n5396) );
  NAND2_X1 U6925 ( .A1(n5377), .A2(SI_15_), .ZN(n5378) );
  MUX2_X1 U6926 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6574), .Z(n5402) );
  XNOR2_X1 U6927 ( .A(n5402), .B(SI_16_), .ZN(n5379) );
  XNOR2_X1 U6928 ( .A(n5406), .B(n5379), .ZN(n6935) );
  NAND2_X1 U6929 ( .A1(n6935), .A2(n8792), .ZN(n5382) );
  NAND2_X1 U6930 ( .A1(n4408), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5380) );
  XNOR2_X1 U6931 ( .A(n5380), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9128) );
  AOI22_X1 U6932 ( .A1(n5457), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5086), .B2(
        n9128), .ZN(n5381) );
  NAND2_X1 U6933 ( .A1(n9494), .A2(n5622), .ZN(n5391) );
  NAND2_X1 U6934 ( .A1(n5072), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6935 ( .A1(n8769), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5388) );
  INV_X1 U6936 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U6937 ( .A1(n5384), .A2(n5383), .ZN(n5385) );
  AND2_X1 U6938 ( .A1(n5412), .A2(n5385), .ZN(n9375) );
  NAND2_X1 U6939 ( .A1(n4316), .A2(n9375), .ZN(n5387) );
  NAND2_X1 U6940 ( .A1(n5101), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5386) );
  OR2_X1 U6941 ( .A1(n9499), .A2(n4321), .ZN(n5390) );
  NAND2_X1 U6942 ( .A1(n5391), .A2(n5390), .ZN(n5392) );
  XNOR2_X1 U6943 ( .A(n5392), .B(n4324), .ZN(n5397) );
  NAND2_X1 U6944 ( .A1(n9494), .A2(n5697), .ZN(n5394) );
  OR2_X1 U6945 ( .A1(n9499), .A2(n4323), .ZN(n5393) );
  NAND2_X1 U6946 ( .A1(n5394), .A2(n5393), .ZN(n5398) );
  NAND2_X1 U6947 ( .A1(n5397), .A2(n5398), .ZN(n8657) );
  NAND2_X1 U6948 ( .A1(n8661), .A2(n8756), .ZN(n5395) );
  NAND2_X1 U6949 ( .A1(n5396), .A2(n4927), .ZN(n5401) );
  INV_X1 U6950 ( .A(n5397), .ZN(n5400) );
  INV_X1 U6951 ( .A(n5398), .ZN(n5399) );
  NAND2_X1 U6952 ( .A1(n5400), .A2(n5399), .ZN(n8656) );
  NAND2_X1 U6953 ( .A1(n5401), .A2(n8656), .ZN(n8674) );
  INV_X1 U6954 ( .A(SI_16_), .ZN(n5403) );
  NOR2_X1 U6955 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  INV_X1 U6956 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7103) );
  INV_X1 U6957 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5407) );
  MUX2_X1 U6958 ( .A(n7103), .B(n5407), .S(n6574), .Z(n5427) );
  XNOR2_X1 U6959 ( .A(n5427), .B(SI_17_), .ZN(n5429) );
  XNOR2_X1 U6960 ( .A(n5430), .B(n5429), .ZN(n7058) );
  NAND2_X1 U6961 ( .A1(n7058), .A2(n8792), .ZN(n5410) );
  XNOR2_X1 U6962 ( .A(n5408), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9688) );
  AOI22_X1 U6963 ( .A1(n5457), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5086), .B2(
        n9688), .ZN(n5409) );
  NAND2_X1 U6964 ( .A1(n9487), .A2(n5622), .ZN(n5419) );
  INV_X1 U6965 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5411) );
  AND2_X1 U6966 ( .A1(n5412), .A2(n5411), .ZN(n5413) );
  OR2_X1 U6967 ( .A1(n5413), .A2(n5460), .ZN(n9358) );
  INV_X1 U6968 ( .A(n4317), .ZN(n5491) );
  NAND2_X1 U6969 ( .A1(n5072), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6970 ( .A1(n8769), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5414) );
  AND2_X1 U6971 ( .A1(n5415), .A2(n5414), .ZN(n5417) );
  NAND2_X1 U6972 ( .A1(n5101), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5416) );
  OAI211_X1 U6973 ( .C1(n9358), .C2(n5491), .A(n5417), .B(n5416), .ZN(n9473)
         );
  NAND2_X1 U6974 ( .A1(n9473), .A2(n5697), .ZN(n5418) );
  NAND2_X1 U6975 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  XNOR2_X1 U6976 ( .A(n5420), .B(n4324), .ZN(n5422) );
  AND2_X1 U6977 ( .A1(n9473), .A2(n5654), .ZN(n5421) );
  AOI21_X1 U6978 ( .B1(n9487), .B2(n5697), .A(n5421), .ZN(n5423) );
  XNOR2_X1 U6979 ( .A(n5422), .B(n5423), .ZN(n8673) );
  NAND2_X1 U6980 ( .A1(n8674), .A2(n8673), .ZN(n5426) );
  INV_X1 U6981 ( .A(n5422), .ZN(n5424) );
  NAND2_X1 U6982 ( .A1(n5424), .A2(n5423), .ZN(n5425) );
  NAND2_X1 U6983 ( .A1(n5426), .A2(n5425), .ZN(n8614) );
  INV_X1 U6984 ( .A(n5427), .ZN(n5428) );
  MUX2_X1 U6985 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6574), .Z(n5431) );
  NAND2_X1 U6986 ( .A1(n5431), .A2(SI_18_), .ZN(n5436) );
  INV_X1 U6987 ( .A(n5431), .ZN(n5433) );
  INV_X1 U6988 ( .A(SI_18_), .ZN(n5432) );
  NAND2_X1 U6989 ( .A1(n5433), .A2(n5432), .ZN(n5434) );
  NAND2_X1 U6990 ( .A1(n5436), .A2(n5434), .ZN(n5448) );
  INV_X1 U6991 ( .A(n5448), .ZN(n5435) );
  MUX2_X1 U6992 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n4320), .Z(n5476) );
  XNOR2_X1 U6993 ( .A(n5476), .B(SI_19_), .ZN(n5480) );
  XNOR2_X1 U6994 ( .A(n5481), .B(n5480), .ZN(n7230) );
  NAND2_X1 U6995 ( .A1(n7230), .A2(n8792), .ZN(n5438) );
  AOI22_X1 U6996 ( .A1(n5457), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9136), .B2(
        n5086), .ZN(n5437) );
  NAND2_X1 U6997 ( .A1(n9324), .A2(n5622), .ZN(n5443) );
  NOR2_X1 U6998 ( .A1(n5462), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5439) );
  OR2_X1 U6999 ( .A1(n5484), .A2(n5439), .ZN(n9325) );
  AOI22_X1 U7000 ( .A1(n5072), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n5101), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U7001 ( .A1(n8769), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5440) );
  OAI211_X1 U7002 ( .C1(n9325), .C2(n5491), .A(n5441), .B(n5440), .ZN(n9476)
         );
  NAND2_X1 U7003 ( .A1(n9476), .A2(n5697), .ZN(n5442) );
  NAND2_X1 U7004 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  XNOR2_X1 U7005 ( .A(n5444), .B(n4324), .ZN(n8619) );
  NAND2_X1 U7006 ( .A1(n9324), .A2(n5697), .ZN(n5446) );
  NAND2_X1 U7007 ( .A1(n9476), .A2(n5654), .ZN(n5445) );
  NAND2_X1 U7008 ( .A1(n5446), .A2(n5445), .ZN(n5471) );
  INV_X1 U7009 ( .A(n5447), .ZN(n5449) );
  NAND2_X1 U7010 ( .A1(n5449), .A2(n5448), .ZN(n5450) );
  NAND2_X1 U7011 ( .A1(n5451), .A2(n5450), .ZN(n7167) );
  OR2_X1 U7012 ( .A1(n5454), .A2(n5453), .ZN(n5455) );
  AND2_X1 U7013 ( .A1(n5456), .A2(n5455), .ZN(n9717) );
  AOI22_X1 U7014 ( .A1(n5457), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5086), .B2(
        n9717), .ZN(n5458) );
  NAND2_X1 U7015 ( .A1(n9350), .A2(n5697), .ZN(n5466) );
  NOR2_X1 U7016 ( .A1(n5460), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5461) );
  OR2_X1 U7017 ( .A1(n5462), .A2(n5461), .ZN(n9342) );
  AOI22_X1 U7018 ( .A1(n8769), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n5072), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U7019 ( .A1(n5101), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5463) );
  OAI211_X1 U7020 ( .C1(n9342), .C2(n5491), .A(n5464), .B(n5463), .ZN(n9465)
         );
  NAND2_X1 U7021 ( .A1(n9465), .A2(n5654), .ZN(n5465) );
  NAND2_X1 U7022 ( .A1(n5466), .A2(n5465), .ZN(n8735) );
  NAND2_X1 U7023 ( .A1(n9350), .A2(n5622), .ZN(n5468) );
  NAND2_X1 U7024 ( .A1(n9465), .A2(n5697), .ZN(n5467) );
  NAND2_X1 U7025 ( .A1(n5468), .A2(n5467), .ZN(n5469) );
  XNOR2_X1 U7026 ( .A(n5469), .B(n4324), .ZN(n8615) );
  OAI22_X1 U7027 ( .A1(n8619), .A2(n5471), .B1(n8735), .B2(n8615), .ZN(n5475)
         );
  NAND2_X1 U7028 ( .A1(n8615), .A2(n8735), .ZN(n5470) );
  INV_X1 U7029 ( .A(n5471), .ZN(n8618) );
  NAND2_X1 U7030 ( .A1(n5470), .A2(n8618), .ZN(n5473) );
  INV_X1 U7031 ( .A(n5470), .ZN(n5472) );
  AOI22_X1 U7032 ( .A1(n8619), .A2(n5473), .B1(n5472), .B2(n5471), .ZN(n5474)
         );
  INV_X1 U7033 ( .A(n5476), .ZN(n5478) );
  INV_X1 U7034 ( .A(SI_19_), .ZN(n5477) );
  NAND2_X1 U7035 ( .A1(n5478), .A2(n5477), .ZN(n5479) );
  INV_X1 U7036 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7329) );
  INV_X1 U7037 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7344) );
  MUX2_X1 U7038 ( .A(n7329), .B(n7344), .S(n4320), .Z(n5501) );
  XNOR2_X1 U7039 ( .A(n5501), .B(SI_20_), .ZN(n5498) );
  NAND2_X1 U7040 ( .A1(n7328), .A2(n8792), .ZN(n5483) );
  OR2_X1 U7041 ( .A1(n8794), .A2(n7344), .ZN(n5482) );
  NAND2_X1 U7042 ( .A1(n9460), .A2(n5622), .ZN(n5493) );
  NOR2_X1 U7043 ( .A1(n5484), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5485) );
  OR2_X1 U7044 ( .A1(n5507), .A2(n5485), .ZN(n9311) );
  INV_X1 U7045 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U7046 ( .A1(n5072), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U7047 ( .A1(n5101), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5486) );
  OAI211_X1 U7048 ( .C1(n5488), .C2(n5074), .A(n5487), .B(n5486), .ZN(n5489)
         );
  INV_X1 U7049 ( .A(n5489), .ZN(n5490) );
  OAI21_X1 U7050 ( .B1(n9311), .B2(n5491), .A(n5490), .ZN(n9466) );
  NAND2_X1 U7051 ( .A1(n9466), .A2(n5697), .ZN(n5492) );
  NAND2_X1 U7052 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  XNOR2_X1 U7053 ( .A(n5494), .B(n5705), .ZN(n8691) );
  AND2_X1 U7054 ( .A1(n9466), .A2(n5654), .ZN(n5495) );
  AOI21_X1 U7055 ( .B1(n9460), .B2(n5697), .A(n5495), .ZN(n5496) );
  INV_X1 U7056 ( .A(n8691), .ZN(n5497) );
  INV_X1 U7057 ( .A(n5496), .ZN(n8690) );
  NAND2_X1 U7058 ( .A1(n5499), .A2(n5498), .ZN(n5503) );
  INV_X1 U7059 ( .A(SI_20_), .ZN(n5500) );
  NAND2_X1 U7060 ( .A1(n5501), .A2(n5500), .ZN(n5502) );
  INV_X1 U7061 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7346) );
  INV_X1 U7062 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7381) );
  MUX2_X1 U7063 ( .A(n7346), .B(n7381), .S(n4320), .Z(n5525) );
  XNOR2_X1 U7064 ( .A(n5525), .B(SI_21_), .ZN(n5504) );
  XNOR2_X1 U7065 ( .A(n5523), .B(n5504), .ZN(n7345) );
  NAND2_X1 U7066 ( .A1(n7345), .A2(n8792), .ZN(n5506) );
  OR2_X1 U7067 ( .A1(n8794), .A2(n7381), .ZN(n5505) );
  OR2_X1 U7068 ( .A1(n5507), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5508) );
  AND2_X1 U7069 ( .A1(n5508), .A2(n5535), .ZN(n9293) );
  NAND2_X1 U7070 ( .A1(n9293), .A2(n4316), .ZN(n5515) );
  INV_X1 U7071 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7072 ( .A1(n5101), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7073 ( .A1(n8769), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5509) );
  OAI211_X1 U7074 ( .C1(n5512), .C2(n5511), .A(n5510), .B(n5509), .ZN(n5513)
         );
  INV_X1 U7075 ( .A(n5513), .ZN(n5514) );
  OAI22_X1 U7076 ( .A1(n9295), .A2(n5596), .B1(n9458), .B2(n4321), .ZN(n5516)
         );
  XNOR2_X1 U7077 ( .A(n5516), .B(n4324), .ZN(n5519) );
  OR2_X1 U7078 ( .A1(n9295), .A2(n4321), .ZN(n5518) );
  NAND2_X1 U7079 ( .A1(n9283), .A2(n5654), .ZN(n5517) );
  NAND2_X1 U7080 ( .A1(n5518), .A2(n5517), .ZN(n5520) );
  XNOR2_X1 U7081 ( .A(n5519), .B(n5520), .ZN(n8627) );
  INV_X1 U7082 ( .A(n5519), .ZN(n5522) );
  INV_X1 U7083 ( .A(n5520), .ZN(n5521) );
  INV_X1 U7084 ( .A(SI_21_), .ZN(n5524) );
  NAND2_X1 U7085 ( .A1(n5525), .A2(n5524), .ZN(n5545) );
  NAND2_X1 U7086 ( .A1(n5609), .A2(n5545), .ZN(n5527) );
  INV_X1 U7087 ( .A(n5525), .ZN(n5526) );
  NAND2_X1 U7088 ( .A1(n5526), .A2(SI_21_), .ZN(n5549) );
  INV_X1 U7089 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7479) );
  INV_X1 U7090 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7481) );
  MUX2_X1 U7091 ( .A(n7479), .B(n7481), .S(n4320), .Z(n5529) );
  INV_X1 U7092 ( .A(SI_22_), .ZN(n5528) );
  NAND2_X1 U7093 ( .A1(n5529), .A2(n5528), .ZN(n5546) );
  INV_X1 U7094 ( .A(n5529), .ZN(n5530) );
  NAND2_X1 U7095 ( .A1(n5530), .A2(SI_22_), .ZN(n5531) );
  NAND2_X1 U7096 ( .A1(n5546), .A2(n5531), .ZN(n5547) );
  NAND2_X1 U7097 ( .A1(n7478), .A2(n8792), .ZN(n5534) );
  OR2_X1 U7098 ( .A1(n8794), .A2(n7481), .ZN(n5533) );
  NAND2_X1 U7099 ( .A1(n5101), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7100 ( .A1(n5072), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5540) );
  NOR2_X1 U7101 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n5536), .ZN(n5537) );
  NOR2_X1 U7102 ( .A1(n5560), .A2(n5537), .ZN(n9278) );
  NAND2_X1 U7103 ( .A1(n4316), .A2(n9278), .ZN(n5539) );
  NAND2_X1 U7104 ( .A1(n8769), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5538) );
  OAI22_X1 U7105 ( .A1(n9280), .A2(n5596), .B1(n9439), .B2(n4321), .ZN(n5542)
         );
  XNOR2_X1 U7106 ( .A(n5542), .B(n5705), .ZN(n5543) );
  NOR2_X2 U7107 ( .A1(n5544), .A2(n5543), .ZN(n8711) );
  OAI22_X1 U7108 ( .A1(n9280), .A2(n4321), .B1(n9439), .B2(n4315), .ZN(n8710)
         );
  NOR2_X2 U7109 ( .A1(n8711), .A2(n8710), .ZN(n8709) );
  AND2_X1 U7110 ( .A1(n5545), .A2(n5546), .ZN(n5576) );
  NAND2_X1 U7111 ( .A1(n5609), .A2(n5576), .ZN(n5552) );
  INV_X1 U7112 ( .A(n5546), .ZN(n5551) );
  INV_X1 U7113 ( .A(n5547), .ZN(n5548) );
  INV_X1 U7114 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7460) );
  INV_X1 U7115 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7456) );
  MUX2_X1 U7116 ( .A(n7460), .B(n7456), .S(n4320), .Z(n5554) );
  INV_X1 U7117 ( .A(SI_23_), .ZN(n5553) );
  NAND2_X1 U7118 ( .A1(n5554), .A2(n5553), .ZN(n5577) );
  INV_X1 U7119 ( .A(n5554), .ZN(n5555) );
  NAND2_X1 U7120 ( .A1(n5555), .A2(SI_23_), .ZN(n5556) );
  NAND2_X1 U7121 ( .A1(n7457), .A2(n8792), .ZN(n5559) );
  OR2_X1 U7122 ( .A1(n8794), .A2(n7456), .ZN(n5558) );
  NAND2_X1 U7123 ( .A1(n9441), .A2(n5622), .ZN(n5568) );
  NAND2_X1 U7124 ( .A1(n5101), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7125 ( .A1(n5072), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5565) );
  NOR2_X1 U7126 ( .A1(n5560), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5561) );
  NOR2_X1 U7127 ( .A1(n5590), .A2(n5561), .ZN(n9268) );
  NAND2_X1 U7128 ( .A1(n4316), .A2(n9268), .ZN(n5564) );
  NAND2_X1 U7129 ( .A1(n8769), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5563) );
  NAND4_X1 U7130 ( .A1(n5566), .A2(n5565), .A3(n5564), .A4(n5563), .ZN(n9284)
         );
  NAND2_X1 U7131 ( .A1(n9284), .A2(n5697), .ZN(n5567) );
  NAND2_X1 U7132 ( .A1(n5568), .A2(n5567), .ZN(n5569) );
  XNOR2_X1 U7133 ( .A(n5569), .B(n5705), .ZN(n5571) );
  AND2_X1 U7134 ( .A1(n9284), .A2(n5654), .ZN(n5570) );
  AOI21_X1 U7135 ( .B1(n9441), .B2(n5697), .A(n5570), .ZN(n5572) );
  NAND2_X1 U7136 ( .A1(n5571), .A2(n5572), .ZN(n8681) );
  INV_X1 U7137 ( .A(n5571), .ZN(n5574) );
  INV_X1 U7138 ( .A(n5572), .ZN(n5573) );
  NAND2_X1 U7139 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  AND2_X1 U7140 ( .A1(n5576), .A2(n5577), .ZN(n5607) );
  NAND2_X1 U7141 ( .A1(n5609), .A2(n5607), .ZN(n5582) );
  INV_X1 U7142 ( .A(n5577), .ZN(n5581) );
  INV_X1 U7143 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7453) );
  INV_X1 U7144 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7484) );
  MUX2_X1 U7145 ( .A(n7453), .B(n7484), .S(n6574), .Z(n5584) );
  INV_X1 U7146 ( .A(SI_24_), .ZN(n5583) );
  NAND2_X1 U7147 ( .A1(n5584), .A2(n5583), .ZN(n5610) );
  INV_X1 U7148 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U7149 ( .A1(n5585), .A2(SI_24_), .ZN(n5586) );
  NAND2_X1 U7150 ( .A1(n7452), .A2(n8792), .ZN(n5589) );
  OR2_X1 U7151 ( .A1(n8794), .A2(n7484), .ZN(n5588) );
  NAND2_X1 U7152 ( .A1(n5072), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7153 ( .A1(n8769), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5594) );
  NOR2_X1 U7154 ( .A1(n5590), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5591) );
  NOR2_X1 U7155 ( .A1(n5623), .A2(n5591), .ZN(n9255) );
  NAND2_X1 U7156 ( .A1(n4317), .A2(n9255), .ZN(n5593) );
  NAND2_X1 U7157 ( .A1(n5101), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5592) );
  OAI22_X1 U7158 ( .A1(n9249), .A2(n5596), .B1(n9438), .B2(n4321), .ZN(n5597)
         );
  XNOR2_X1 U7159 ( .A(n5597), .B(n5705), .ZN(n5600) );
  OR2_X1 U7160 ( .A1(n9438), .A2(n4315), .ZN(n5598) );
  NAND2_X1 U7161 ( .A1(n5600), .A2(n5601), .ZN(n5605) );
  INV_X1 U7162 ( .A(n5600), .ZN(n5603) );
  INV_X1 U7163 ( .A(n5601), .ZN(n5602) );
  NAND2_X1 U7164 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  NAND2_X1 U7165 ( .A1(n5605), .A2(n5604), .ZN(n8680) );
  INV_X1 U7166 ( .A(n5605), .ZN(n5606) );
  INV_X1 U7167 ( .A(n5610), .ZN(n5614) );
  INV_X1 U7168 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n10066) );
  INV_X1 U7169 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7499) );
  MUX2_X1 U7170 ( .A(n10066), .B(n7499), .S(n6574), .Z(n5616) );
  INV_X1 U7171 ( .A(SI_25_), .ZN(n5615) );
  NAND2_X1 U7172 ( .A1(n5616), .A2(n5615), .ZN(n5639) );
  INV_X1 U7173 ( .A(n5616), .ZN(n5617) );
  NAND2_X1 U7174 ( .A1(n5617), .A2(SI_25_), .ZN(n5618) );
  NAND2_X1 U7175 ( .A1(n7476), .A2(n8792), .ZN(n5621) );
  OR2_X1 U7176 ( .A1(n8794), .A2(n7499), .ZN(n5620) );
  NAND2_X1 U7177 ( .A1(n9427), .A2(n5622), .ZN(n5631) );
  NAND2_X1 U7178 ( .A1(n5072), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7179 ( .A1(n5101), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5628) );
  INV_X1 U7180 ( .A(n5623), .ZN(n5625) );
  INV_X1 U7181 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U7182 ( .A1(n5623), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5648) );
  INV_X1 U7183 ( .A(n5648), .ZN(n5647) );
  AOI21_X1 U7184 ( .B1(n5625), .B2(n5624), .A(n5647), .ZN(n9239) );
  NAND2_X1 U7185 ( .A1(n4317), .A2(n9239), .ZN(n5627) );
  NAND2_X1 U7186 ( .A1(n8769), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5626) );
  NAND4_X1 U7187 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n5626), .ZN(n9415)
         );
  NAND2_X1 U7188 ( .A1(n9415), .A2(n5697), .ZN(n5630) );
  NAND2_X1 U7189 ( .A1(n5631), .A2(n5630), .ZN(n5632) );
  XNOR2_X1 U7190 ( .A(n5632), .B(n4324), .ZN(n5634) );
  OAI22_X1 U7191 ( .A1(n9245), .A2(n4321), .B1(n9227), .B2(n5702), .ZN(n5633)
         );
  XNOR2_X1 U7192 ( .A(n5634), .B(n5633), .ZN(n8649) );
  NOR2_X1 U7193 ( .A1(n5634), .A2(n5633), .ZN(n8746) );
  INV_X1 U7194 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7501) );
  INV_X1 U7195 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7521) );
  MUX2_X1 U7196 ( .A(n7501), .B(n7521), .S(n4320), .Z(n5642) );
  INV_X1 U7197 ( .A(SI_26_), .ZN(n5641) );
  NAND2_X1 U7198 ( .A1(n5642), .A2(n5641), .ZN(n5665) );
  INV_X1 U7199 ( .A(n5642), .ZN(n5643) );
  NAND2_X1 U7200 ( .A1(n5643), .A2(SI_26_), .ZN(n5644) );
  NAND2_X1 U7201 ( .A1(n7500), .A2(n8792), .ZN(n5646) );
  OR2_X1 U7202 ( .A1(n8794), .A2(n7521), .ZN(n5645) );
  NAND2_X1 U7203 ( .A1(n5101), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7204 ( .A1(n5072), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5652) );
  INV_X1 U7205 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7206 ( .A1(n5647), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5673) );
  INV_X1 U7207 ( .A(n5673), .ZN(n5675) );
  AOI21_X1 U7208 ( .B1(n5649), .B2(n5648), .A(n5675), .ZN(n9224) );
  NAND2_X1 U7209 ( .A1(n4317), .A2(n9224), .ZN(n5651) );
  NAND2_X1 U7210 ( .A1(n8769), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5650) );
  AND2_X1 U7211 ( .A1(n9242), .A2(n5654), .ZN(n5655) );
  AOI21_X1 U7212 ( .B1(n9229), .B2(n5697), .A(n5655), .ZN(n5660) );
  NAND2_X1 U7213 ( .A1(n9229), .A2(n5622), .ZN(n5657) );
  NAND2_X1 U7214 ( .A1(n9242), .A2(n5697), .ZN(n5656) );
  NAND2_X1 U7215 ( .A1(n5657), .A2(n5656), .ZN(n5659) );
  XNOR2_X1 U7216 ( .A(n5659), .B(n4324), .ZN(n5662) );
  XOR2_X1 U7217 ( .A(n5660), .B(n5662), .Z(n8745) );
  INV_X1 U7218 ( .A(n5660), .ZN(n5661) );
  INV_X1 U7219 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6135) );
  INV_X1 U7220 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7596) );
  MUX2_X1 U7221 ( .A(n6135), .B(n7596), .S(n6574), .Z(n5668) );
  INV_X1 U7222 ( .A(SI_27_), .ZN(n5667) );
  NAND2_X1 U7223 ( .A1(n5668), .A2(n5667), .ZN(n5689) );
  INV_X1 U7224 ( .A(n5668), .ZN(n5669) );
  NAND2_X1 U7225 ( .A1(n5669), .A2(SI_27_), .ZN(n5670) );
  NAND2_X1 U7226 ( .A1(n7555), .A2(n8792), .ZN(n5672) );
  OR2_X1 U7227 ( .A1(n8794), .A2(n7596), .ZN(n5671) );
  NAND2_X1 U7228 ( .A1(n9411), .A2(n5622), .ZN(n5682) );
  NAND2_X1 U7229 ( .A1(n5072), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7230 ( .A1(n8769), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5679) );
  INV_X1 U7231 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7232 ( .A1(n5674), .A2(n5673), .ZN(n5676) );
  NAND2_X1 U7233 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n5675), .ZN(n5746) );
  NAND2_X1 U7234 ( .A1(n4316), .A2(n9212), .ZN(n5678) );
  NAND2_X1 U7235 ( .A1(n5101), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5677) );
  OR2_X1 U7236 ( .A1(n9198), .A2(n4321), .ZN(n5681) );
  NAND2_X1 U7237 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  XNOR2_X1 U7238 ( .A(n5683), .B(n5705), .ZN(n5686) );
  NOR2_X1 U7239 ( .A1(n9198), .A2(n4323), .ZN(n5684) );
  AOI21_X1 U7240 ( .B1(n9411), .B2(n5697), .A(n5684), .ZN(n5685) );
  NAND2_X1 U7241 ( .A1(n5686), .A2(n5685), .ZN(n5756) );
  OAI21_X1 U7242 ( .B1(n5686), .B2(n5685), .A(n5756), .ZN(n6430) );
  INV_X1 U7243 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10080) );
  INV_X1 U7244 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7654) );
  MUX2_X1 U7245 ( .A(n10080), .B(n7654), .S(n4320), .Z(n5692) );
  INV_X1 U7246 ( .A(SI_28_), .ZN(n5691) );
  NAND2_X1 U7247 ( .A1(n5692), .A2(n5691), .ZN(n6160) );
  INV_X1 U7248 ( .A(n5692), .ZN(n5693) );
  NAND2_X1 U7249 ( .A1(n5693), .A2(SI_28_), .ZN(n5694) );
  AND2_X1 U7250 ( .A1(n6160), .A2(n5694), .ZN(n6158) );
  NAND2_X1 U7251 ( .A1(n7585), .A2(n8792), .ZN(n5696) );
  OR2_X1 U7252 ( .A1(n8794), .A2(n7654), .ZN(n5695) );
  NAND2_X1 U7253 ( .A1(n9401), .A2(n5697), .ZN(n5704) );
  NAND2_X1 U7254 ( .A1(n5072), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U7255 ( .A1(n5101), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5700) );
  XNOR2_X1 U7256 ( .A(n5746), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9200) );
  NAND2_X1 U7257 ( .A1(n4317), .A2(n9200), .ZN(n5699) );
  NAND2_X1 U7258 ( .A1(n8769), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5698) );
  OR2_X1 U7259 ( .A1(n9408), .A2(n4315), .ZN(n5703) );
  NAND2_X1 U7260 ( .A1(n5704), .A2(n5703), .ZN(n5706) );
  XNOR2_X1 U7261 ( .A(n5706), .B(n5705), .ZN(n5709) );
  NAND2_X1 U7262 ( .A1(n9401), .A2(n5622), .ZN(n5707) );
  OAI21_X1 U7263 ( .B1(n9408), .B2(n4321), .A(n5707), .ZN(n5708) );
  XNOR2_X1 U7264 ( .A(n5709), .B(n5708), .ZN(n5734) );
  NAND2_X1 U7265 ( .A1(n7497), .A2(P1_B_REG_SCAN_IN), .ZN(n5710) );
  MUX2_X1 U7266 ( .A(P1_B_REG_SCAN_IN), .B(n5710), .S(n7482), .Z(n5711) );
  NAND2_X1 U7267 ( .A1(n5711), .A2(n5712), .ZN(n6596) );
  INV_X1 U7268 ( .A(n5712), .ZN(n7519) );
  NAND2_X1 U7269 ( .A1(n7519), .A2(n7497), .ZN(n9563) );
  OAI21_X1 U7270 ( .B1(n6596), .B2(P1_D_REG_1__SCAN_IN), .A(n9563), .ZN(n6683)
         );
  INV_X1 U7271 ( .A(n6683), .ZN(n5725) );
  INV_X1 U7272 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5713) );
  AND2_X1 U7273 ( .A1(n7482), .A2(n7519), .ZN(n6598) );
  NOR4_X1 U7274 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5722) );
  NOR4_X1 U7275 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5721) );
  INV_X1 U7276 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9976) );
  INV_X1 U7277 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9975) );
  INV_X1 U7278 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9979) );
  INV_X1 U7279 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10019) );
  NAND4_X1 U7280 ( .A1(n9976), .A2(n9975), .A3(n9979), .A4(n10019), .ZN(n5719)
         );
  NOR4_X1 U7281 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5717) );
  NOR4_X1 U7282 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5716) );
  NOR4_X1 U7283 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5715) );
  NOR4_X1 U7284 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5714) );
  NAND4_X1 U7285 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n5718)
         );
  NOR4_X1 U7286 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5719), .A4(n5718), .ZN(n5720) );
  NAND3_X1 U7287 ( .A1(n5722), .A2(n5721), .A3(n5720), .ZN(n5723) );
  NAND2_X1 U7288 ( .A1(n5724), .A2(n5723), .ZN(n7008) );
  NAND3_X1 U7289 ( .A1(n5725), .A2(n6777), .A3(n7008), .ZN(n5751) );
  NAND2_X1 U7290 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  NAND2_X1 U7291 ( .A1(n5728), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5730) );
  XNOR2_X1 U7292 ( .A(n5730), .B(n5729), .ZN(n6602) );
  INV_X1 U7293 ( .A(n9009), .ZN(n6632) );
  INV_X1 U7294 ( .A(n5731), .ZN(n6689) );
  INV_X1 U7295 ( .A(n7379), .ZN(n8957) );
  NAND2_X1 U7296 ( .A1(n5732), .A2(n8957), .ZN(n6687) );
  INV_X1 U7297 ( .A(n6687), .ZN(n9002) );
  OR2_X1 U7298 ( .A1(n9762), .A2(n9002), .ZN(n5733) );
  NOR2_X2 U7299 ( .A1(n5742), .A2(n5733), .ZN(n8748) );
  NAND3_X1 U7300 ( .A1(n6434), .A2(n5734), .A3(n8748), .ZN(n5761) );
  INV_X1 U7301 ( .A(n5734), .ZN(n5757) );
  NAND3_X1 U7302 ( .A1(n5757), .A2(n8748), .A3(n5756), .ZN(n5735) );
  INV_X1 U7303 ( .A(n5742), .ZN(n5744) );
  NAND2_X1 U7304 ( .A1(n6688), .A2(n5736), .ZN(n7017) );
  INV_X1 U7305 ( .A(n7017), .ZN(n5737) );
  NAND2_X1 U7306 ( .A1(n5744), .A2(n5737), .ZN(n5739) );
  NAND2_X1 U7307 ( .A1(n9452), .A2(n9136), .ZN(n6681) );
  INV_X1 U7308 ( .A(n6681), .ZN(n5738) );
  NAND2_X1 U7309 ( .A1(n9474), .A2(n5731), .ZN(n5741) );
  NOR2_X2 U7310 ( .A1(n5742), .A2(n5741), .ZN(n8757) );
  INV_X1 U7311 ( .A(n8757), .ZN(n8728) );
  AND2_X1 U7312 ( .A1(n9475), .A2(n5731), .ZN(n5743) );
  NAND2_X1 U7313 ( .A1(n5744), .A2(n5743), .ZN(n8759) );
  NAND2_X1 U7314 ( .A1(n5072), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7315 ( .A1(n8769), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5749) );
  INV_X1 U7316 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5745) );
  NOR2_X1 U7317 ( .A1(n5746), .A2(n5745), .ZN(n9169) );
  NAND2_X1 U7318 ( .A1(n4316), .A2(n9169), .ZN(n5748) );
  NAND2_X1 U7319 ( .A1(n5101), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5747) );
  INV_X1 U7320 ( .A(n9197), .ZN(n9026) );
  AOI22_X1 U7321 ( .A1(n8726), .A2(n9026), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5755) );
  NAND2_X1 U7322 ( .A1(n5751), .A2(n6681), .ZN(n5752) );
  OR2_X1 U7323 ( .A1(n6687), .A2(n5731), .ZN(n7007) );
  NAND2_X1 U7324 ( .A1(n5752), .A2(n7007), .ZN(n6633) );
  OAI21_X1 U7325 ( .B1(n6633), .B2(n6454), .A(P1_STATE_REG_SCAN_IN), .ZN(n5753) );
  OR2_X1 U7326 ( .A1(n6602), .A2(P1_U3086), .ZN(n9024) );
  NAND2_X1 U7327 ( .A1(n8763), .A2(n9200), .ZN(n5754) );
  OAI211_X1 U7328 ( .C1(n9198), .C2(n8728), .A(n5755), .B(n5754), .ZN(n5759)
         );
  NOR3_X1 U7329 ( .A1(n5757), .A2(n5756), .A3(n8766), .ZN(n5758) );
  AOI211_X1 U7330 ( .C1(n9401), .C2(n8741), .A(n5759), .B(n5758), .ZN(n5760)
         );
  INV_X1 U7331 ( .A(n5860), .ZN(n5768) );
  NOR2_X1 U7332 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5769) );
  NAND4_X1 U7333 ( .A1(n5769), .A2(n5784), .A3(n5999), .A4(n10034), .ZN(n5771)
         );
  NAND4_X1 U7334 ( .A1(n5787), .A2(n6030), .A3(n5781), .A4(n5782), .ZN(n5770)
         );
  INV_X1 U7335 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5793) );
  INV_X1 U7336 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7337 ( .A1(n7230), .A2(n7893), .ZN(n5792) );
  INV_X1 U7338 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5988) );
  AND4_X1 U7339 ( .A1(n5988), .A2(n5999), .A3(n10034), .A4(n5782), .ZN(n5783)
         );
  NAND2_X1 U7340 ( .A1(n6029), .A2(n6030), .ZN(n6044) );
  INV_X1 U7341 ( .A(n6044), .ZN(n5785) );
  NAND2_X1 U7342 ( .A1(n5785), .A2(n5784), .ZN(n5786) );
  NAND2_X1 U7343 ( .A1(n6055), .A2(n5787), .ZN(n5788) );
  INV_X1 U7344 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5789) );
  AOI22_X1 U7345 ( .A1(n6057), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8096), .B2(
        n6056), .ZN(n5791) );
  NAND2_X1 U7346 ( .A1(n5794), .A2(n5793), .ZN(n5797) );
  INV_X1 U7347 ( .A(n5797), .ZN(n5795) );
  INV_X1 U7348 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5798) );
  INV_X1 U7349 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U7350 ( .A1(n5797), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5799) );
  INV_X1 U7351 ( .A(n5815), .ZN(n5800) );
  INV_X1 U7352 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7527) );
  INV_X1 U7353 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5808) );
  INV_X1 U7354 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5810) );
  INV_X1 U7355 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10048) );
  INV_X1 U7356 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10033) );
  NAND2_X1 U7357 ( .A1(n6063), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7358 ( .A1(n6071), .A2(n5814), .ZN(n8352) );
  NAND2_X1 U7359 ( .A1(n6164), .A2(n8352), .ZN(n5821) );
  INV_X1 U7360 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8482) );
  OR2_X1 U7361 ( .A1(n7027), .A2(n8482), .ZN(n5820) );
  INV_X1 U7362 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5817) );
  OR2_X1 U7363 ( .A1(n6060), .A2(n5817), .ZN(n5819) );
  INV_X1 U7364 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8550) );
  OR2_X1 U7365 ( .A1(n5823), .A2(n8550), .ZN(n5818) );
  INV_X1 U7366 ( .A(n8360), .ZN(n8114) );
  INV_X1 U7367 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5822) );
  OR2_X1 U7368 ( .A1(n6060), .A2(n9990), .ZN(n5826) );
  NAND2_X1 U7369 ( .A1(n5880), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5825) );
  INV_X1 U7370 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6677) );
  OR2_X1 U7371 ( .A1(n5910), .A2(n6677), .ZN(n5824) );
  INV_X1 U7372 ( .A(n5842), .ZN(n5834) );
  OR2_X1 U7373 ( .A1(n4325), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5830) );
  AND2_X1 U7374 ( .A1(n5830), .A2(n4921), .ZN(n5833) );
  OR2_X1 U7375 ( .A1(n6054), .A2(n5831), .ZN(n5832) );
  INV_X1 U7376 ( .A(n9850), .ZN(n6460) );
  NAND2_X1 U7377 ( .A1(n5842), .A2(n9850), .ZN(n7936) );
  NAND2_X1 U7378 ( .A1(n7938), .A2(n7936), .ZN(n6181) );
  NAND2_X1 U7379 ( .A1(n5880), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5836) );
  INV_X1 U7380 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6308) );
  INV_X1 U7381 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5835) );
  INV_X1 U7382 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6680) );
  NAND2_X1 U7383 ( .A1(n4586), .A2(SI_0_), .ZN(n5838) );
  INV_X1 U7384 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U7385 ( .A1(n5838), .A2(n5837), .ZN(n5840) );
  AND2_X1 U7386 ( .A1(n5840), .A2(n5839), .ZN(n8583) );
  NAND2_X1 U7387 ( .A1(n8127), .A2(n9848), .ZN(n5841) );
  NAND2_X1 U7388 ( .A1(n6181), .A2(n5841), .ZN(n6924) );
  NAND2_X1 U7389 ( .A1(n6924), .A2(n6942), .ZN(n5855) );
  NAND2_X1 U7390 ( .A1(n5938), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5848) );
  INV_X1 U7391 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5843) );
  OR2_X1 U7392 ( .A1(n7027), .A2(n5843), .ZN(n5847) );
  INV_X1 U7393 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5844) );
  INV_X1 U7394 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6788) );
  OR2_X1 U7395 ( .A1(n5910), .A2(n6788), .ZN(n5845) );
  OR2_X1 U7396 ( .A1(n6054), .A2(n6589), .ZN(n5853) );
  OR2_X1 U7397 ( .A1(n4326), .A2(n4732), .ZN(n5852) );
  OR2_X1 U7398 ( .A1(n5829), .A2(n6588), .ZN(n5851) );
  NAND2_X1 U7399 ( .A1(n6466), .A2(n5854), .ZN(n6184) );
  NAND2_X1 U7400 ( .A1(n8126), .A2(n9855), .ZN(n7944) );
  OR2_X1 U7401 ( .A1(n8126), .A2(n5854), .ZN(n6978) );
  INV_X1 U7402 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6359) );
  NOR2_X1 U7403 ( .A1(n4907), .A2(n4359), .ZN(n5858) );
  INV_X1 U7404 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6982) );
  OR2_X1 U7405 ( .A1(n6060), .A2(n6982), .ZN(n5857) );
  OR2_X1 U7406 ( .A1(n5910), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5856) );
  OR2_X1 U7407 ( .A1(n6054), .A2(n6581), .ZN(n5864) );
  OR2_X1 U7408 ( .A1(n5849), .A2(n6582), .ZN(n5863) );
  NAND2_X1 U7409 ( .A1(n5850), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5859) );
  MUX2_X1 U7410 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5859), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5861) );
  OR2_X1 U7411 ( .A1(n5829), .A2(n6649), .ZN(n5862) );
  NAND2_X1 U7412 ( .A1(n5867), .A2(n9860), .ZN(n7950) );
  NAND2_X1 U7413 ( .A1(n7962), .A2(n7950), .ZN(n7906) );
  INV_X1 U7414 ( .A(n9860), .ZN(n6983) );
  OR2_X1 U7415 ( .A1(n5867), .A2(n6983), .ZN(n5868) );
  NAND2_X1 U7416 ( .A1(n6207), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5874) );
  INV_X1 U7417 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7111) );
  OR2_X1 U7418 ( .A1(n6060), .A2(n7111), .ZN(n5873) );
  NAND2_X1 U7419 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5869) );
  AND2_X1 U7420 ( .A1(n5882), .A2(n5869), .ZN(n6968) );
  OR2_X1 U7421 ( .A1(n5910), .A2(n6968), .ZN(n5872) );
  INV_X1 U7422 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5870) );
  OR2_X1 U7423 ( .A1(n5823), .A2(n5870), .ZN(n5871) );
  OR2_X1 U7424 ( .A1(n6054), .A2(n6583), .ZN(n5879) );
  OR2_X1 U7425 ( .A1(n5849), .A2(n6584), .ZN(n5878) );
  NAND2_X1 U7426 ( .A1(n5860), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5876) );
  OR2_X1 U7427 ( .A1(n5829), .A2(n6856), .ZN(n5877) );
  NAND2_X1 U7428 ( .A1(n5880), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5887) );
  INV_X1 U7429 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5881) );
  OR2_X1 U7430 ( .A1(n7027), .A2(n5881), .ZN(n5886) );
  NAND2_X1 U7431 ( .A1(n5882), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5883) );
  AND2_X1 U7432 ( .A1(n5894), .A2(n5883), .ZN(n7162) );
  OR2_X1 U7433 ( .A1(n5910), .A2(n7162), .ZN(n5885) );
  OR2_X1 U7434 ( .A1(n6060), .A2(n7161), .ZN(n5884) );
  NAND4_X1 U7435 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n8124)
         );
  OR2_X1 U7436 ( .A1(n5860), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7437 ( .A1(n5900), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5889) );
  INV_X1 U7438 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5888) );
  OR2_X1 U7439 ( .A1(n6054), .A2(n6586), .ZN(n5891) );
  OR2_X1 U7440 ( .A1(n5849), .A2(n6587), .ZN(n5890) );
  OAI211_X1 U7441 ( .C1(n5829), .C2(n6585), .A(n5891), .B(n5890), .ZN(n7078)
         );
  NAND2_X1 U7442 ( .A1(n8124), .A2(n7078), .ZN(n5892) );
  NAND2_X1 U7443 ( .A1(n5893), .A2(n5892), .ZN(n7233) );
  NAND2_X1 U7444 ( .A1(n5880), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5899) );
  INV_X1 U7445 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7235) );
  OR2_X1 U7446 ( .A1(n6060), .A2(n7235), .ZN(n5898) );
  INV_X1 U7447 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6357) );
  OR2_X1 U7448 ( .A1(n7027), .A2(n6357), .ZN(n5897) );
  NAND2_X1 U7449 ( .A1(n5894), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5895) );
  AND2_X1 U7450 ( .A1(n5908), .A2(n5895), .ZN(n7236) );
  OR2_X1 U7451 ( .A1(n5910), .A2(n7236), .ZN(n5896) );
  NAND4_X1 U7452 ( .A1(n5899), .A2(n5898), .A3(n5897), .A4(n5896), .ZN(n8432)
         );
  NOR2_X1 U7453 ( .A1(n5900), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5916) );
  OR2_X1 U7454 ( .A1(n5916), .A2(n6031), .ZN(n5901) );
  OR2_X1 U7455 ( .A1(n6054), .A2(n6591), .ZN(n5903) );
  OR2_X1 U7456 ( .A1(n5849), .A2(n9991), .ZN(n5902) );
  OAI211_X1 U7457 ( .C1(n5829), .C2(n6990), .A(n5903), .B(n5902), .ZN(n7238)
         );
  AND2_X1 U7458 ( .A1(n8432), .A2(n7238), .ZN(n5904) );
  OR2_X1 U7459 ( .A1(n8432), .A2(n7238), .ZN(n5905) );
  NAND2_X1 U7460 ( .A1(n5880), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5914) );
  INV_X1 U7461 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5906) );
  OR2_X1 U7462 ( .A1(n6060), .A2(n5906), .ZN(n5913) );
  INV_X1 U7463 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5907) );
  OR2_X1 U7464 ( .A1(n7027), .A2(n5907), .ZN(n5912) );
  NAND2_X1 U7465 ( .A1(n5908), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5909) );
  AND2_X1 U7466 ( .A1(n5924), .A2(n5909), .ZN(n8428) );
  OR2_X1 U7467 ( .A1(n5910), .A2(n8428), .ZN(n5911) );
  OR2_X1 U7468 ( .A1(n5849), .A2(n6595), .ZN(n5921) );
  NAND2_X1 U7469 ( .A1(n5916), .A2(n5915), .ZN(n5918) );
  NAND2_X1 U7470 ( .A1(n5918), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5917) );
  MUX2_X1 U7471 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5917), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5919) );
  OR2_X1 U7472 ( .A1(n5829), .A2(n6593), .ZN(n5920) );
  NAND2_X1 U7473 ( .A1(n8123), .A2(n9882), .ZN(n7368) );
  NOR2_X1 U7474 ( .A1(n8123), .A2(n4688), .ZN(n5922) );
  NAND2_X1 U7475 ( .A1(n5880), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5929) );
  INV_X1 U7476 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7374) );
  OR2_X1 U7477 ( .A1(n6060), .A2(n7374), .ZN(n5928) );
  INV_X1 U7478 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5923) );
  OR2_X1 U7479 ( .A1(n7027), .A2(n5923), .ZN(n5927) );
  NAND2_X1 U7480 ( .A1(n5924), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5925) );
  AND2_X1 U7481 ( .A1(n5940), .A2(n5925), .ZN(n7445) );
  OR2_X1 U7482 ( .A1(n5910), .A2(n7445), .ZN(n5926) );
  NAND4_X1 U7483 ( .A1(n5929), .A2(n5928), .A3(n5927), .A4(n5926), .ZN(n8431)
         );
  NAND2_X1 U7484 ( .A1(n6599), .A2(n7893), .ZN(n5932) );
  NAND2_X1 U7485 ( .A1(n5934), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5930) );
  XNOR2_X1 U7486 ( .A(n5930), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7397) );
  AOI22_X1 U7487 ( .A1(n6057), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6056), .B2(
        n7397), .ZN(n5931) );
  OR2_X1 U7488 ( .A1(n8431), .A2(n9888), .ZN(n7976) );
  NAND2_X1 U7489 ( .A1(n8431), .A2(n9888), .ZN(n7971) );
  NAND2_X1 U7490 ( .A1(n7976), .A2(n7971), .ZN(n7912) );
  INV_X1 U7491 ( .A(n9888), .ZN(n7448) );
  NAND2_X1 U7492 ( .A1(n8431), .A2(n7448), .ZN(n5933) );
  NAND2_X1 U7493 ( .A1(n6608), .A2(n7893), .ZN(n5937) );
  OAI21_X1 U7494 ( .B1(n5934), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5935) );
  XNOR2_X1 U7495 ( .A(n5935), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6377) );
  AOI22_X1 U7496 ( .A1(n6057), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6056), .B2(
        n6377), .ZN(n5936) );
  NAND2_X1 U7497 ( .A1(n5937), .A2(n5936), .ZN(n7541) );
  NAND2_X1 U7498 ( .A1(n5938), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5946) );
  INV_X1 U7499 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5939) );
  OR2_X1 U7500 ( .A1(n7027), .A2(n5939), .ZN(n5945) );
  NAND2_X1 U7501 ( .A1(n5940), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5941) );
  AND2_X1 U7502 ( .A1(n5956), .A2(n5941), .ZN(n7550) );
  OR2_X1 U7503 ( .A1(n5910), .A2(n7550), .ZN(n5944) );
  INV_X1 U7504 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5942) );
  OR2_X1 U7505 ( .A1(n5823), .A2(n5942), .ZN(n5943) );
  NAND4_X1 U7506 ( .A1(n5946), .A2(n5945), .A3(n5944), .A4(n5943), .ZN(n8122)
         );
  OR2_X1 U7507 ( .A1(n7541), .A2(n8122), .ZN(n5947) );
  NAND2_X1 U7508 ( .A1(n7425), .A2(n5947), .ZN(n5949) );
  NAND2_X1 U7509 ( .A1(n7541), .A2(n8122), .ZN(n5948) );
  NAND2_X1 U7510 ( .A1(n6612), .A2(n7893), .ZN(n5955) );
  NAND2_X1 U7511 ( .A1(n5950), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5951) );
  MUX2_X1 U7512 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5951), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n5952) );
  INV_X1 U7513 ( .A(n5952), .ZN(n5953) );
  NOR2_X1 U7514 ( .A1(n5953), .A2(n5780), .ZN(n6323) );
  AOI22_X1 U7515 ( .A1(n6057), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6056), .B2(
        n6323), .ZN(n5954) );
  NAND2_X1 U7516 ( .A1(n5955), .A2(n5954), .ZN(n9899) );
  NAND2_X1 U7517 ( .A1(n5938), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5962) );
  INV_X1 U7518 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6290) );
  OR2_X1 U7519 ( .A1(n7027), .A2(n6290), .ZN(n5961) );
  NAND2_X1 U7520 ( .A1(n5956), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5957) );
  AND2_X1 U7521 ( .A1(n5967), .A2(n5957), .ZN(n7579) );
  OR2_X1 U7522 ( .A1(n5910), .A2(n7579), .ZN(n5960) );
  INV_X1 U7523 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5958) );
  OR2_X1 U7524 ( .A1(n5823), .A2(n5958), .ZN(n5959) );
  NAND4_X1 U7525 ( .A1(n5962), .A2(n5961), .A3(n5960), .A4(n5959), .ZN(n8121)
         );
  AND2_X1 U7526 ( .A1(n9899), .A2(n8121), .ZN(n7503) );
  NAND2_X1 U7527 ( .A1(n6623), .A2(n7893), .ZN(n5966) );
  NOR2_X1 U7528 ( .A1(n5780), .A2(n6031), .ZN(n5963) );
  MUX2_X1 U7529 ( .A(n6031), .B(n5963), .S(P2_IR_REG_11__SCAN_IN), .Z(n5964)
         );
  NOR2_X1 U7530 ( .A1(n5964), .A2(n5989), .ZN(n6324) );
  AOI22_X1 U7531 ( .A1(n6057), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6056), .B2(
        n6324), .ZN(n5965) );
  NAND2_X1 U7532 ( .A1(n5966), .A2(n5965), .ZN(n7513) );
  NAND2_X1 U7533 ( .A1(n5880), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5972) );
  INV_X1 U7534 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7606) );
  OR2_X1 U7535 ( .A1(n7027), .A2(n7606), .ZN(n5971) );
  INV_X1 U7536 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7609) );
  OR2_X1 U7537 ( .A1(n6060), .A2(n7609), .ZN(n5970) );
  NAND2_X1 U7538 ( .A1(n5967), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5968) );
  AND2_X1 U7539 ( .A1(n5982), .A2(n5968), .ZN(n7514) );
  OR2_X1 U7540 ( .A1(n5910), .A2(n7514), .ZN(n5969) );
  INV_X1 U7541 ( .A(n7578), .ZN(n8120) );
  AND2_X1 U7542 ( .A1(n7513), .A2(n8120), .ZN(n5974) );
  OR2_X1 U7543 ( .A1(n7503), .A2(n5974), .ZN(n5973) );
  INV_X1 U7544 ( .A(n5973), .ZN(n5977) );
  OR2_X1 U7545 ( .A1(n7513), .A2(n7578), .ZN(n7990) );
  NAND2_X1 U7546 ( .A1(n7513), .A2(n7578), .ZN(n7989) );
  INV_X1 U7547 ( .A(n7916), .ZN(n7508) );
  OR2_X1 U7548 ( .A1(n9899), .A2(n8121), .ZN(n7504) );
  AND2_X1 U7549 ( .A1(n7508), .A2(n7504), .ZN(n7505) );
  INV_X1 U7550 ( .A(n5975), .ZN(n5976) );
  NAND2_X1 U7551 ( .A1(n6650), .A2(n7893), .ZN(n5980) );
  OR2_X1 U7552 ( .A1(n5989), .A2(n6031), .ZN(n5978) );
  XNOR2_X1 U7553 ( .A(n5978), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6387) );
  AOI22_X1 U7554 ( .A1(n6057), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6056), .B2(
        n6387), .ZN(n5979) );
  NAND2_X1 U7555 ( .A1(n5880), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5987) );
  INV_X1 U7556 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6388) );
  OR2_X1 U7557 ( .A1(n7027), .A2(n6388), .ZN(n5986) );
  INV_X1 U7558 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5981) );
  OR2_X1 U7559 ( .A1(n6060), .A2(n5981), .ZN(n5985) );
  NAND2_X1 U7560 ( .A1(n5982), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5983) );
  AND2_X1 U7561 ( .A1(n5993), .A2(n5983), .ZN(n7640) );
  OR2_X1 U7562 ( .A1(n5910), .A2(n7640), .ZN(n5984) );
  NAND4_X1 U7563 ( .A1(n5987), .A2(n5986), .A3(n5985), .A4(n5984), .ZN(n8119)
         );
  NAND2_X1 U7564 ( .A1(n6668), .A2(n7893), .ZN(n5992) );
  NAND2_X1 U7565 ( .A1(n5989), .A2(n5988), .ZN(n5990) );
  NAND2_X1 U7566 ( .A1(n5990), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6000) );
  XNOR2_X1 U7567 ( .A(n6000), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8159) );
  AOI22_X1 U7568 ( .A1(n6057), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6056), .B2(
        n8159), .ZN(n5991) );
  NAND2_X1 U7569 ( .A1(n5880), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5998) );
  INV_X1 U7570 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6351) );
  OR2_X1 U7571 ( .A1(n6060), .A2(n6351), .ZN(n5997) );
  INV_X1 U7572 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8506) );
  OR2_X1 U7573 ( .A1(n7027), .A2(n8506), .ZN(n5996) );
  NAND2_X1 U7574 ( .A1(n5993), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5994) );
  AND2_X1 U7575 ( .A1(n6007), .A2(n5994), .ZN(n7600) );
  OR2_X1 U7576 ( .A1(n5910), .A2(n7600), .ZN(n5995) );
  NAND4_X1 U7577 ( .A1(n5998), .A2(n5997), .A3(n5996), .A4(n5995), .ZN(n8409)
         );
  NAND2_X1 U7578 ( .A1(n7599), .A2(n8409), .ZN(n8403) );
  NAND2_X1 U7579 ( .A1(n6823), .A2(n7893), .ZN(n6005) );
  NAND2_X1 U7580 ( .A1(n6000), .A2(n5999), .ZN(n6001) );
  NAND2_X1 U7581 ( .A1(n6001), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7582 ( .A1(n6002), .A2(n10034), .ZN(n6015) );
  OR2_X1 U7583 ( .A1(n6002), .A2(n10034), .ZN(n6003) );
  NAND2_X1 U7584 ( .A1(n6015), .A2(n6003), .ZN(n6824) );
  INV_X1 U7585 ( .A(n6824), .ZN(n8181) );
  AOI22_X1 U7586 ( .A1(n6057), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6056), .B2(
        n8181), .ZN(n6004) );
  NAND2_X1 U7587 ( .A1(n5880), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6012) );
  INV_X1 U7588 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7589 ( .A1(n7027), .A2(n6006), .ZN(n6011) );
  INV_X1 U7590 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6348) );
  OR2_X1 U7591 ( .A1(n6060), .A2(n6348), .ZN(n6010) );
  NAND2_X1 U7592 ( .A1(n6007), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6008) );
  AND2_X1 U7593 ( .A1(n6019), .A2(n6008), .ZN(n8412) );
  OR2_X1 U7594 ( .A1(n5910), .A2(n8412), .ZN(n6009) );
  NAND4_X1 U7595 ( .A1(n6012), .A2(n6011), .A3(n6010), .A4(n6009), .ZN(n8118)
         );
  NAND2_X1 U7596 ( .A1(n8500), .A2(n8118), .ZN(n6193) );
  INV_X1 U7597 ( .A(n6193), .ZN(n6014) );
  OR2_X1 U7598 ( .A1(n7599), .A2(n8409), .ZN(n8405) );
  OR2_X1 U7599 ( .A1(n8500), .A2(n8118), .ZN(n7931) );
  AND2_X1 U7600 ( .A1(n8405), .A2(n7931), .ZN(n6013) );
  NAND2_X1 U7601 ( .A1(n6866), .A2(n7893), .ZN(n6018) );
  NAND2_X1 U7602 ( .A1(n6015), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6016) );
  XNOR2_X1 U7603 ( .A(n6016), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8198) );
  AOI22_X1 U7604 ( .A1(n6057), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6056), .B2(
        n8198), .ZN(n6017) );
  NAND2_X1 U7605 ( .A1(n5880), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6024) );
  INV_X1 U7606 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8498) );
  OR2_X1 U7607 ( .A1(n7027), .A2(n8498), .ZN(n6023) );
  INV_X1 U7608 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8191) );
  OR2_X1 U7609 ( .A1(n6060), .A2(n8191), .ZN(n6022) );
  NAND2_X1 U7610 ( .A1(n6019), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6020) );
  AND2_X1 U7611 ( .A1(n6037), .A2(n6020), .ZN(n7662) );
  OR2_X1 U7612 ( .A1(n5910), .A2(n7662), .ZN(n6021) );
  OR2_X1 U7613 ( .A1(n7645), .A2(n8389), .ZN(n8008) );
  NAND2_X1 U7614 ( .A1(n7645), .A2(n8389), .ZN(n8006) );
  INV_X1 U7615 ( .A(n8002), .ZN(n6025) );
  AND2_X1 U7616 ( .A1(n7656), .A2(n6025), .ZN(n6026) );
  NAND2_X1 U7617 ( .A1(n7657), .A2(n6026), .ZN(n6028) );
  INV_X1 U7618 ( .A(n8389), .ZN(n8410) );
  NAND2_X1 U7619 ( .A1(n7645), .A2(n8410), .ZN(n6027) );
  NAND2_X1 U7620 ( .A1(n6028), .A2(n6027), .ZN(n8387) );
  NAND2_X1 U7621 ( .A1(n6935), .A2(n7893), .ZN(n6036) );
  NOR2_X1 U7622 ( .A1(n6029), .A2(n6031), .ZN(n6032) );
  MUX2_X1 U7623 ( .A(n6032), .B(n6031), .S(n6030), .Z(n6033) );
  INV_X1 U7624 ( .A(n6033), .ZN(n6034) );
  AND2_X1 U7625 ( .A1(n6044), .A2(n6034), .ZN(n8216) );
  AOI22_X1 U7626 ( .A1(n6057), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6056), .B2(
        n8216), .ZN(n6035) );
  NAND2_X1 U7627 ( .A1(n5880), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6042) );
  INV_X1 U7628 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8397) );
  OR2_X1 U7629 ( .A1(n6060), .A2(n8397), .ZN(n6041) );
  INV_X1 U7630 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8494) );
  OR2_X1 U7631 ( .A1(n7027), .A2(n8494), .ZN(n6040) );
  NAND2_X1 U7632 ( .A1(n6037), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6038) );
  AND2_X1 U7633 ( .A1(n6048), .A2(n6038), .ZN(n8396) );
  OR2_X1 U7634 ( .A1(n5910), .A2(n8396), .ZN(n6039) );
  NAND2_X1 U7635 ( .A1(n8395), .A2(n8374), .ZN(n8014) );
  NAND2_X1 U7636 ( .A1(n8012), .A2(n8014), .ZN(n8393) );
  INV_X1 U7637 ( .A(n8374), .ZN(n8117) );
  AND2_X1 U7638 ( .A1(n8395), .A2(n8117), .ZN(n6043) );
  NAND2_X1 U7639 ( .A1(n7058), .A2(n7893), .ZN(n6047) );
  NAND2_X1 U7640 ( .A1(n6044), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6045) );
  XNOR2_X1 U7641 ( .A(n6045), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8233) );
  AOI22_X1 U7642 ( .A1(n6057), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6056), .B2(
        n8233), .ZN(n6046) );
  NAND2_X1 U7643 ( .A1(n5880), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6053) );
  INV_X1 U7644 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8380) );
  OR2_X1 U7645 ( .A1(n6060), .A2(n8380), .ZN(n6052) );
  INV_X1 U7646 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8221) );
  OR2_X1 U7647 ( .A1(n7027), .A2(n8221), .ZN(n6051) );
  NAND2_X1 U7648 ( .A1(n6048), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6049) );
  AND2_X1 U7649 ( .A1(n6061), .A2(n6049), .ZN(n8379) );
  OR2_X1 U7650 ( .A1(n5910), .A2(n8379), .ZN(n6050) );
  OR2_X1 U7651 ( .A1(n8383), .A2(n8391), .ZN(n8015) );
  NAND2_X1 U7652 ( .A1(n8383), .A2(n8391), .ZN(n8021) );
  INV_X1 U7653 ( .A(n8383), .ZN(n8488) );
  OR2_X1 U7654 ( .A1(n7167), .A2(n6054), .ZN(n6059) );
  XNOR2_X1 U7655 ( .A(n6055), .B(P2_IR_REG_18__SCAN_IN), .ZN(n6398) );
  AOI22_X1 U7656 ( .A1(n6057), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6056), .B2(
        n6398), .ZN(n6058) );
  NAND2_X1 U7657 ( .A1(n6207), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6067) );
  INV_X1 U7658 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8364) );
  OR2_X1 U7659 ( .A1(n6060), .A2(n8364), .ZN(n6066) );
  NAND2_X1 U7660 ( .A1(n6061), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6062) );
  AND2_X1 U7661 ( .A1(n6063), .A2(n6062), .ZN(n8363) );
  OR2_X1 U7662 ( .A1(n5910), .A2(n8363), .ZN(n6065) );
  INV_X1 U7663 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8554) );
  OR2_X1 U7664 ( .A1(n5823), .A2(n8554), .ZN(n6064) );
  NOR2_X1 U7665 ( .A1(n8556), .A2(n8375), .ZN(n6068) );
  INV_X1 U7666 ( .A(n8375), .ZN(n8115) );
  NAND2_X1 U7667 ( .A1(n8351), .A2(n8360), .ZN(n8027) );
  NAND2_X1 U7668 ( .A1(n7328), .A2(n7893), .ZN(n6070) );
  OR2_X1 U7669 ( .A1(n5849), .A2(n7329), .ZN(n6069) );
  NAND2_X1 U7670 ( .A1(n6071), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7671 ( .A1(n6082), .A2(n6072), .ZN(n8339) );
  NAND2_X1 U7672 ( .A1(n8339), .A2(n6164), .ZN(n6076) );
  NAND2_X1 U7673 ( .A1(n5938), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7674 ( .A1(n6207), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7675 ( .A1(n5880), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6073) );
  NAND2_X1 U7676 ( .A1(n7836), .A2(n8346), .ZN(n8323) );
  NAND2_X1 U7677 ( .A1(n8030), .A2(n8323), .ZN(n8337) );
  INV_X1 U7678 ( .A(n8346), .ZN(n8113) );
  NAND2_X1 U7679 ( .A1(n8332), .A2(n6077), .ZN(n8320) );
  NAND2_X1 U7680 ( .A1(n7345), .A2(n7893), .ZN(n6079) );
  OR2_X1 U7681 ( .A1(n5849), .A2(n7346), .ZN(n6078) );
  INV_X1 U7682 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7683 ( .A1(n6082), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7684 ( .A1(n6091), .A2(n6083), .ZN(n8327) );
  NAND2_X1 U7685 ( .A1(n8327), .A2(n6164), .ZN(n6086) );
  AOI22_X1 U7686 ( .A1(n6207), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5938), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U7687 ( .A1(n5880), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7688 ( .A1(n7738), .A2(n8336), .ZN(n8035) );
  NAND2_X1 U7689 ( .A1(n8034), .A2(n8035), .ZN(n7904) );
  NAND2_X1 U7690 ( .A1(n7478), .A2(n7893), .ZN(n6090) );
  OR2_X1 U7691 ( .A1(n5849), .A2(n7479), .ZN(n6089) );
  OR2_X2 U7692 ( .A1(n6091), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7693 ( .A1(n6091), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7694 ( .A1(n6098), .A2(n6092), .ZN(n8315) );
  NAND2_X1 U7695 ( .A1(n8315), .A2(n6164), .ZN(n6095) );
  AOI22_X1 U7696 ( .A1(n6207), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n5938), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7697 ( .A1(n5880), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7698 ( .A1(n7841), .A2(n8322), .ZN(n8037) );
  INV_X1 U7699 ( .A(n8322), .ZN(n8112) );
  NAND2_X1 U7700 ( .A1(n7457), .A2(n7893), .ZN(n6097) );
  OR2_X1 U7701 ( .A1(n5849), .A2(n7460), .ZN(n6096) );
  NAND2_X1 U7702 ( .A1(n6098), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7703 ( .A1(n6108), .A2(n6099), .ZN(n8305) );
  NAND2_X1 U7704 ( .A1(n8305), .A2(n6164), .ZN(n6104) );
  INV_X1 U7705 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8534) );
  NAND2_X1 U7706 ( .A1(n5938), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7707 ( .A1(n6207), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6100) );
  OAI211_X1 U7708 ( .C1(n8534), .C2(n5823), .A(n6101), .B(n6100), .ZN(n6102)
         );
  INV_X1 U7709 ( .A(n6102), .ZN(n6103) );
  NAND2_X1 U7710 ( .A1(n6104), .A2(n6103), .ZN(n8111) );
  NOR2_X1 U7711 ( .A1(n7767), .A2(n8111), .ZN(n6105) );
  NAND2_X1 U7712 ( .A1(n7452), .A2(n7893), .ZN(n6107) );
  OR2_X1 U7713 ( .A1(n5849), .A2(n7453), .ZN(n6106) );
  INV_X1 U7714 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U7715 ( .A1(n6108), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7716 ( .A1(n6120), .A2(n6109), .ZN(n8295) );
  NAND2_X1 U7717 ( .A1(n8295), .A2(n6164), .ZN(n6114) );
  INV_X1 U7718 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n10078) );
  NAND2_X1 U7719 ( .A1(n5880), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7720 ( .A1(n6207), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6110) );
  OAI211_X1 U7721 ( .C1(n6060), .C2(n10078), .A(n6111), .B(n6110), .ZN(n6112)
         );
  INV_X1 U7722 ( .A(n6112), .ZN(n6113) );
  NOR2_X1 U7723 ( .A1(n8532), .A2(n8302), .ZN(n6115) );
  NAND2_X1 U7724 ( .A1(n7476), .A2(n7893), .ZN(n6117) );
  INV_X1 U7725 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7726 ( .A1(n6120), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7727 ( .A1(n6128), .A2(n6121), .ZN(n8285) );
  NAND2_X1 U7728 ( .A1(n8285), .A2(n6164), .ZN(n6126) );
  INV_X1 U7729 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8526) );
  NAND2_X1 U7730 ( .A1(n5938), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7731 ( .A1(n6207), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6122) );
  OAI211_X1 U7732 ( .C1(n8526), .C2(n5823), .A(n6123), .B(n6122), .ZN(n6124)
         );
  INV_X1 U7733 ( .A(n6124), .ZN(n6125) );
  NOR2_X1 U7734 ( .A1(n5849), .A2(n7501), .ZN(n6127) );
  OR2_X2 U7735 ( .A1(n6128), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7736 ( .A1(n6128), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7737 ( .A1(n6140), .A2(n6129), .ZN(n8276) );
  NAND2_X1 U7738 ( .A1(n8276), .A2(n6164), .ZN(n6134) );
  INV_X1 U7739 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8522) );
  NAND2_X1 U7740 ( .A1(n6207), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7741 ( .A1(n5938), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6130) );
  OAI211_X1 U7742 ( .C1(n8522), .C2(n5823), .A(n6131), .B(n6130), .ZN(n6132)
         );
  INV_X1 U7743 ( .A(n6132), .ZN(n6133) );
  NAND2_X1 U7744 ( .A1(n7555), .A2(n7893), .ZN(n6137) );
  OR2_X1 U7745 ( .A1(n5849), .A2(n6135), .ZN(n6136) );
  INV_X1 U7746 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7747 ( .A1(n6140), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7748 ( .A1(n8264), .A2(n6164), .ZN(n6146) );
  INV_X1 U7749 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U7750 ( .A1(n5938), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7751 ( .A1(n6207), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6142) );
  OAI211_X1 U7752 ( .C1(n6448), .C2(n5823), .A(n6143), .B(n6142), .ZN(n6144)
         );
  INV_X1 U7753 ( .A(n6144), .ZN(n6145) );
  NAND2_X1 U7754 ( .A1(n7754), .A2(n8107), .ZN(n6147) );
  NAND2_X1 U7755 ( .A1(n7585), .A2(n7893), .ZN(n6149) );
  OR2_X1 U7756 ( .A1(n4326), .A2(n10080), .ZN(n6148) );
  NAND2_X1 U7757 ( .A1(n6150), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7758 ( .A1(n7720), .A2(n6151), .ZN(n7710) );
  NAND2_X1 U7759 ( .A1(n7710), .A2(n6164), .ZN(n6156) );
  INV_X1 U7760 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n7711) );
  NAND2_X1 U7761 ( .A1(n6207), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7762 ( .A1(n5880), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6152) );
  OAI211_X1 U7763 ( .C1(n6060), .C2(n7711), .A(n6153), .B(n6152), .ZN(n6154)
         );
  INV_X1 U7764 ( .A(n6154), .ZN(n6155) );
  NAND2_X1 U7765 ( .A1(n8076), .A2(n8077), .ZN(n6157) );
  INV_X1 U7766 ( .A(n8077), .ZN(n8106) );
  INV_X1 U7767 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7729) );
  INV_X1 U7768 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10018) );
  MUX2_X1 U7769 ( .A(n7729), .B(n10018), .S(n6574), .Z(n7675) );
  NAND2_X1 U7770 ( .A1(n8793), .A2(n7893), .ZN(n6163) );
  OR2_X1 U7771 ( .A1(n4326), .A2(n7729), .ZN(n6162) );
  INV_X1 U7772 ( .A(n7720), .ZN(n6165) );
  NAND2_X1 U7773 ( .A1(n6165), .A2(n6164), .ZN(n7030) );
  INV_X1 U7774 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7775 ( .A1(n6207), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7776 ( .A1(n5938), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6166) );
  OAI211_X1 U7777 ( .C1(n5823), .C2(n6168), .A(n6167), .B(n6166), .ZN(n6169)
         );
  INV_X1 U7778 ( .A(n6169), .ZN(n6170) );
  NAND2_X1 U7779 ( .A1(n6255), .A2(n7779), .ZN(n7882) );
  INV_X1 U7780 ( .A(n6172), .ZN(n6173) );
  NAND2_X1 U7781 ( .A1(n6173), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7782 ( .A1(n8096), .A2(n8100), .ZN(n6419) );
  NAND2_X1 U7783 ( .A1(n6175), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6176) );
  MUX2_X1 U7784 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6176), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n6177) );
  INV_X1 U7785 ( .A(n6177), .ZN(n6178) );
  NAND2_X1 U7786 ( .A1(n6179), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6180) );
  XNOR2_X1 U7787 ( .A(n6180), .B(P2_IR_REG_20__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U7788 ( .A1(n7933), .A2(n6418), .ZN(n7900) );
  INV_X1 U7789 ( .A(n6181), .ZN(n6183) );
  INV_X1 U7790 ( .A(n9848), .ZN(n6926) );
  INV_X1 U7791 ( .A(n7935), .ZN(n6182) );
  NAND2_X1 U7792 ( .A1(n6183), .A2(n6182), .ZN(n6922) );
  NAND2_X1 U7793 ( .A1(n6922), .A2(n7938), .ZN(n6940) );
  INV_X1 U7794 ( .A(n7907), .ZN(n6943) );
  NAND2_X1 U7795 ( .A1(n6940), .A2(n6943), .ZN(n6972) );
  NAND2_X1 U7796 ( .A1(n6972), .A2(n6184), .ZN(n6185) );
  INV_X1 U7797 ( .A(n7906), .ZN(n6979) );
  NAND2_X1 U7798 ( .A1(n6185), .A2(n6979), .ZN(n6974) );
  NAND2_X1 U7799 ( .A1(n6974), .A2(n7962), .ZN(n7108) );
  NAND2_X1 U7800 ( .A1(n8125), .A2(n9867), .ZN(n7960) );
  NAND2_X1 U7801 ( .A1(n7108), .A2(n7960), .ZN(n6186) );
  NAND2_X1 U7802 ( .A1(n6186), .A2(n7952), .ZN(n7157) );
  XNOR2_X1 U7803 ( .A(n8124), .B(n7078), .ZN(n7911) );
  NAND2_X1 U7804 ( .A1(n7157), .A2(n7911), .ZN(n7417) );
  INV_X1 U7805 ( .A(n7078), .ZN(n9870) );
  OR2_X1 U7806 ( .A1(n8124), .A2(n9870), .ZN(n7951) );
  AND2_X1 U7807 ( .A1(n7971), .A2(n7368), .ZN(n7969) );
  INV_X1 U7808 ( .A(n7238), .ZN(n9876) );
  NAND2_X1 U7809 ( .A1(n7969), .A2(n6187), .ZN(n6188) );
  AND2_X1 U7810 ( .A1(n7976), .A2(n6188), .ZN(n6190) );
  AND2_X1 U7811 ( .A1(n7951), .A2(n6190), .ZN(n7416) );
  INV_X1 U7812 ( .A(n8122), .ZN(n7545) );
  OR2_X1 U7813 ( .A1(n7545), .A2(n7541), .ZN(n7463) );
  NAND2_X1 U7814 ( .A1(n7545), .A2(n7541), .ZN(n7977) );
  NAND2_X1 U7815 ( .A1(n7463), .A2(n7977), .ZN(n7424) );
  INV_X1 U7816 ( .A(n7424), .ZN(n7972) );
  AND2_X1 U7817 ( .A1(n7416), .A2(n7972), .ZN(n6189) );
  NAND2_X1 U7818 ( .A1(n7417), .A2(n6189), .ZN(n7421) );
  NAND2_X1 U7819 ( .A1(n8432), .A2(n9876), .ZN(n7964) );
  OR2_X1 U7820 ( .A1(n9899), .A2(n7549), .ZN(n7985) );
  AND2_X1 U7821 ( .A1(n7985), .A2(n7463), .ZN(n7974) );
  NAND2_X1 U7822 ( .A1(n9899), .A2(n7549), .ZN(n7986) );
  XNOR2_X1 U7823 ( .A(n8509), .B(n7994), .ZN(n7637) );
  OR2_X1 U7824 ( .A1(n8509), .A2(n7994), .ZN(n7996) );
  INV_X1 U7825 ( .A(n8409), .ZN(n7629) );
  NAND2_X1 U7826 ( .A1(n7599), .A2(n7629), .ZN(n7999) );
  NAND2_X1 U7827 ( .A1(n7602), .A2(n7999), .ZN(n6192) );
  OR2_X1 U7828 ( .A1(n7599), .A2(n7629), .ZN(n8000) );
  INV_X1 U7829 ( .A(n8118), .ZN(n7660) );
  NAND2_X1 U7830 ( .A1(n8500), .A2(n7660), .ZN(n6195) );
  INV_X1 U7831 ( .A(n8006), .ZN(n6196) );
  NAND2_X1 U7832 ( .A1(n8394), .A2(n8014), .ZN(n6197) );
  NAND2_X1 U7833 ( .A1(n6197), .A2(n8012), .ZN(n8369) );
  INV_X1 U7834 ( .A(n8370), .ZN(n8371) );
  NAND2_X1 U7835 ( .A1(n6198), .A2(n8375), .ZN(n8022) );
  NAND2_X1 U7836 ( .A1(n8024), .A2(n8022), .ZN(n8362) );
  INV_X1 U7837 ( .A(n8023), .ZN(n6199) );
  NAND2_X1 U7838 ( .A1(n8338), .A2(n8030), .ZN(n8324) );
  AND2_X1 U7839 ( .A1(n8035), .A2(n8323), .ZN(n8031) );
  NAND2_X1 U7840 ( .A1(n8324), .A2(n8031), .ZN(n6200) );
  NAND2_X1 U7841 ( .A1(n6200), .A2(n8034), .ZN(n8314) );
  NAND2_X1 U7842 ( .A1(n8314), .A2(n8037), .ZN(n6201) );
  NAND2_X1 U7843 ( .A1(n6201), .A2(n8040), .ZN(n8304) );
  NAND2_X1 U7844 ( .A1(n7767), .A2(n8312), .ZN(n8038) );
  NAND2_X1 U7845 ( .A1(n7754), .A2(n8273), .ZN(n8064) );
  INV_X1 U7846 ( .A(n6232), .ZN(n6203) );
  NAND2_X1 U7847 ( .A1(n7933), .A2(n8090), .ZN(n6930) );
  OR2_X1 U7848 ( .A1(n6203), .A2(n6930), .ZN(n6532) );
  INV_X1 U7849 ( .A(n8100), .ZN(n7932) );
  INV_X1 U7850 ( .A(n7933), .ZN(n7347) );
  NAND2_X1 U7851 ( .A1(n6532), .A2(n9894), .ZN(n6833) );
  AND2_X1 U7852 ( .A1(n6203), .A2(n6458), .ZN(n6204) );
  INV_X1 U7853 ( .A(n6205), .ZN(n6413) );
  XNOR2_X1 U7854 ( .A(n6413), .B(n8098), .ZN(n6551) );
  INV_X1 U7855 ( .A(n6551), .ZN(n6534) );
  INV_X1 U7856 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7857 ( .A1(n5938), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7858 ( .A1(n6207), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6208) );
  OAI211_X1 U7859 ( .C1(n6210), .C2(n5823), .A(n6209), .B(n6208), .ZN(n6211)
         );
  INV_X1 U7860 ( .A(n6211), .ZN(n6212) );
  NAND2_X1 U7861 ( .A1(n7030), .A2(n6212), .ZN(n8105) );
  NAND2_X1 U7862 ( .A1(n5829), .A2(P2_B_REG_SCAN_IN), .ZN(n6213) );
  AND2_X1 U7863 ( .A1(n8430), .A2(n6213), .ZN(n7718) );
  AOI22_X1 U7864 ( .A1(n8433), .A2(n8106), .B1(n8105), .B2(n7718), .ZN(n6214)
         );
  OAI21_X1 U7865 ( .B1(n6217), .B2(n8440), .A(n6214), .ZN(n6215) );
  NAND2_X1 U7866 ( .A1(n8096), .A2(n8090), .ZN(n6421) );
  NAND2_X1 U7867 ( .A1(n6251), .A2(n6252), .ZN(n6220) );
  NAND2_X1 U7868 ( .A1(n6222), .A2(n6221), .ZN(n6224) );
  OR2_X1 U7869 ( .A1(n6222), .A2(n6221), .ZN(n6223) );
  XNOR2_X1 U7870 ( .A(n7454), .B(P2_B_REG_SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7871 ( .A1(n6227), .A2(n7477), .ZN(n6231) );
  NAND2_X1 U7872 ( .A1(n4401), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6228) );
  MUX2_X1 U7873 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6228), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6229) );
  NAND2_X1 U7874 ( .A1(n6229), .A2(n5777), .ZN(n7502) );
  INV_X1 U7875 ( .A(n7502), .ZN(n6230) );
  AOI21_X1 U7876 ( .B1(n6232), .B2(n6418), .A(n8085), .ZN(n6236) );
  NAND2_X1 U7877 ( .A1(n6417), .A2(n6236), .ZN(n6830) );
  NOR2_X1 U7878 ( .A1(n9893), .A2(n7933), .ZN(n6530) );
  OR2_X1 U7879 ( .A1(n6233), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U7880 ( .A1(n7477), .A2(n7502), .ZN(n6234) );
  INV_X1 U7881 ( .A(n6236), .ZN(n6237) );
  NAND2_X1 U7882 ( .A1(n8574), .A2(n6237), .ZN(n6829) );
  OAI21_X1 U7883 ( .B1(n6830), .B2(n6530), .A(n6829), .ZN(n6254) );
  NAND2_X1 U7884 ( .A1(n6417), .A2(n8574), .ZN(n6540) );
  NOR2_X1 U7885 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .ZN(
        n6241) );
  NOR4_X1 U7886 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6240) );
  NOR4_X1 U7887 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6239) );
  NOR4_X1 U7888 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6238) );
  NAND4_X1 U7889 ( .A1(n6241), .A2(n6240), .A3(n6239), .A4(n6238), .ZN(n6247)
         );
  NOR4_X1 U7890 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6245) );
  NOR4_X1 U7891 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6244) );
  NOR4_X1 U7892 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6243) );
  NOR4_X1 U7893 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n6242) );
  NAND4_X1 U7894 ( .A1(n6245), .A2(n6244), .A3(n6243), .A4(n6242), .ZN(n6246)
         );
  NOR2_X1 U7895 ( .A1(n6247), .A2(n6246), .ZN(n6248) );
  INV_X1 U7896 ( .A(n7477), .ZN(n6250) );
  NOR2_X1 U7897 ( .A1(n7454), .A2(n7502), .ZN(n6249) );
  NAND2_X1 U7898 ( .A1(n6250), .A2(n6249), .ZN(n6542) );
  XNOR2_X1 U7899 ( .A(n6251), .B(n6252), .ZN(n7458) );
  NAND2_X1 U7900 ( .A1(n6458), .A2(n8085), .ZN(n6541) );
  NAND2_X1 U7901 ( .A1(n6439), .A2(n9920), .ZN(n6260) );
  NAND2_X1 U7902 ( .A1(n6260), .A2(n6259), .ZN(P2_U3488) );
  INV_X1 U7903 ( .A(n7928), .ZN(n6261) );
  XNOR2_X1 U7904 ( .A(n6262), .B(n6261), .ZN(n6264) );
  OAI22_X1 U7905 ( .A1(n7779), .A2(n8392), .B1(n8273), .B2(n8390), .ZN(n6263)
         );
  XOR2_X1 U7906 ( .A(n7928), .B(n6265), .Z(n7712) );
  NAND2_X1 U7907 ( .A1(n7709), .A2(n6268), .ZN(n6428) );
  NAND2_X1 U7908 ( .A1(n6428), .A2(n9920), .ZN(n6272) );
  INV_X1 U7909 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6269) );
  OR2_X1 U7910 ( .A1(n9920), .A2(n6269), .ZN(n6270) );
  AND2_X1 U7911 ( .A1(n4926), .A2(n6270), .ZN(n6271) );
  INV_X1 U7912 ( .A(n6601), .ZN(n6273) );
  INV_X1 U7913 ( .A(n8085), .ZN(n8070) );
  NAND2_X1 U7914 ( .A1(n6542), .A2(n8070), .ZN(n6274) );
  NAND2_X1 U7915 ( .A1(n6274), .A2(n7458), .ZN(n6412) );
  NAND2_X1 U7916 ( .A1(n6412), .A2(n5829), .ZN(n6275) );
  NAND2_X1 U7917 ( .A1(n6275), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7918 ( .A(n8216), .ZN(n6936) );
  INV_X1 U7919 ( .A(n6377), .ZN(n7323) );
  NAND2_X1 U7920 ( .A1(n6276), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7921 ( .A1(n6364), .A2(n6277), .ZN(n6278) );
  NAND2_X1 U7922 ( .A1(n6309), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7923 ( .A1(n6588), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6280) );
  AND2_X2 U7924 ( .A1(n9804), .A2(n6280), .ZN(n6281) );
  INV_X1 U7925 ( .A(n6282), .ZN(n6842) );
  XNOR2_X1 U7926 ( .A(n6856), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6843) );
  AOI21_X1 U7927 ( .B1(n6585), .B2(n4364), .A(n6564), .ZN(n6996) );
  NAND2_X1 U7928 ( .A1(P2_REG1_REG_6__SCAN_IN), .A2(n6990), .ZN(n6284) );
  OAI21_X1 U7929 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n6990), .A(n6284), .ZN(
        n6995) );
  NOR2_X1 U7930 ( .A1(n6996), .A2(n6995), .ZN(n6994) );
  NOR2_X1 U7931 ( .A1(n9829), .A2(n6286), .ZN(n6287) );
  AOI22_X1 U7932 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n7397), .B1(n6604), .B2(
        n5923), .ZN(n7392) );
  NOR2_X1 U7933 ( .A1(n6377), .A2(n6288), .ZN(n6289) );
  INV_X1 U7934 ( .A(n6323), .ZN(n7361) );
  AOI22_X1 U7935 ( .A1(n6323), .A2(P2_REG1_REG_10__SCAN_IN), .B1(n6290), .B2(
        n7361), .ZN(n7352) );
  INV_X1 U7936 ( .A(n6324), .ZN(n7612) );
  NAND2_X1 U7937 ( .A1(n6292), .A2(n7612), .ZN(n6291) );
  INV_X1 U7938 ( .A(n6291), .ZN(n6293) );
  OAI21_X1 U7939 ( .B1(n6292), .B2(n7612), .A(n6291), .ZN(n7607) );
  INV_X1 U7940 ( .A(n6387), .ZN(n8146) );
  NAND2_X1 U7941 ( .A1(n8146), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7942 ( .A1(n6387), .A2(n6388), .ZN(n6294) );
  NAND2_X1 U7943 ( .A1(n6295), .A2(n6294), .ZN(n8139) );
  NOR2_X1 U7944 ( .A1(n8140), .A2(n8139), .ZN(n8138) );
  INV_X1 U7945 ( .A(n6295), .ZN(n6296) );
  NOR2_X1 U7946 ( .A1(n8159), .A2(n6297), .ZN(n6299) );
  INV_X1 U7947 ( .A(n8159), .ZN(n6705) );
  NAND2_X1 U7948 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6824), .ZN(n6300) );
  OAI21_X1 U7949 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n6824), .A(n6300), .ZN(
        n8168) );
  AOI22_X1 U7950 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8216), .B1(n6936), .B2(
        n8494), .ZN(n8203) );
  NOR2_X1 U7951 ( .A1(n8233), .A2(n6302), .ZN(n6303) );
  INV_X1 U7952 ( .A(n6398), .ZN(n8251) );
  NAND2_X1 U7953 ( .A1(n8251), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6304) );
  OAI21_X1 U7954 ( .B1(n8251), .B2(P2_REG1_REG_18__SCAN_IN), .A(n6304), .ZN(
        n8238) );
  XNOR2_X1 U7955 ( .A(n7231), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6405) );
  INV_X1 U7956 ( .A(n6405), .ZN(n6305) );
  NOR2_X1 U7957 ( .A1(n6205), .A2(P2_U3151), .ZN(n7586) );
  AND2_X1 U7958 ( .A1(n6412), .A2(n7586), .ZN(n6339) );
  INV_X1 U7959 ( .A(n6339), .ZN(n6616) );
  NAND2_X1 U7960 ( .A1(n6309), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U7961 ( .A1(n6310), .A2(n6311), .ZN(n6660) );
  INV_X1 U7962 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9990) );
  OAI21_X1 U7963 ( .B1(n6660), .B2(n9990), .A(n6311), .ZN(n9814) );
  NAND2_X1 U7964 ( .A1(n6588), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6312) );
  NOR2_X2 U7965 ( .A1(n6314), .A2(n6313), .ZN(n6316) );
  INV_X1 U7966 ( .A(n6316), .ZN(n6846) );
  XNOR2_X1 U7967 ( .A(n6856), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6847) );
  INV_X1 U7968 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7161) );
  NAND2_X1 U7969 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n6990), .ZN(n6318) );
  OAI21_X1 U7970 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6990), .A(n6318), .ZN(
        n6992) );
  NOR2_X1 U7971 ( .A1(n9829), .A2(n6319), .ZN(n6320) );
  AOI22_X1 U7972 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n7397), .B1(n6604), .B2(
        n7374), .ZN(n7383) );
  NOR2_X1 U7973 ( .A1(n7384), .A2(n7383), .ZN(n7382) );
  NOR2_X1 U7974 ( .A1(n6377), .A2(n6321), .ZN(n6322) );
  INV_X1 U7975 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7430) );
  XNOR2_X1 U7976 ( .A(n6321), .B(n6377), .ZN(n7316) );
  INV_X1 U7977 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7472) );
  AOI22_X1 U7978 ( .A1(n6323), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7472), .B2(
        n7361), .ZN(n7355) );
  INV_X1 U7979 ( .A(n6325), .ZN(n6326) );
  OR2_X2 U7980 ( .A1(n6325), .A2(n6324), .ZN(n8135) );
  OAI21_X1 U7981 ( .B1(n6326), .B2(n7612), .A(n8135), .ZN(n7610) );
  INV_X1 U7982 ( .A(n7610), .ZN(n6327) );
  XOR2_X1 U7983 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6387), .Z(n8134) );
  AOI21_X1 U7984 ( .B1(n8133), .B2(n8135), .A(n8134), .ZN(n8137) );
  NOR2_X1 U7985 ( .A1(n8159), .A2(n6328), .ZN(n6329) );
  XNOR2_X1 U7986 ( .A(n6328), .B(n8159), .ZN(n8155) );
  NAND2_X1 U7987 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6824), .ZN(n6330) );
  OAI21_X1 U7988 ( .B1(n6824), .B2(P2_REG2_REG_14__SCAN_IN), .A(n6330), .ZN(
        n8177) );
  NOR2_X1 U7989 ( .A1(n8198), .A2(n6331), .ZN(n6332) );
  NAND2_X1 U7990 ( .A1(n6936), .A2(n8397), .ZN(n6334) );
  NAND2_X1 U7991 ( .A1(n8216), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6333) );
  AND2_X1 U7992 ( .A1(n6334), .A2(n6333), .ZN(n8212) );
  NOR2_X1 U7993 ( .A1(n8233), .A2(n6335), .ZN(n6336) );
  NOR2_X1 U7994 ( .A1(n8226), .A2(n6336), .ZN(n8241) );
  NAND2_X1 U7995 ( .A1(n8251), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6337) );
  OAI21_X1 U7996 ( .B1(n8251), .B2(P2_REG2_REG_18__SCAN_IN), .A(n6337), .ZN(
        n8240) );
  INV_X1 U7997 ( .A(n6337), .ZN(n6338) );
  MUX2_X1 U7998 ( .A(n5817), .B(P2_REG2_REG_19__SCAN_IN), .S(n7231), .Z(n6404)
         );
  AND2_X1 U7999 ( .A1(n6339), .A2(n8098), .ZN(n9816) );
  NAND2_X1 U8000 ( .A1(n4314), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6340) );
  OAI21_X1 U8001 ( .B1(n4314), .B2(n8380), .A(n6340), .ZN(n6341) );
  INV_X1 U8002 ( .A(n8233), .ZN(n7104) );
  OR2_X1 U8003 ( .A1(n6341), .A2(n7104), .ZN(n6396) );
  XNOR2_X1 U8004 ( .A(n6341), .B(n8233), .ZN(n8224) );
  NAND2_X1 U8005 ( .A1(n4314), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6342) );
  OAI21_X1 U8006 ( .B1(n4313), .B2(n8397), .A(n6342), .ZN(n6343) );
  OR2_X1 U8007 ( .A1(n6936), .A2(n6343), .ZN(n6395) );
  XNOR2_X1 U8008 ( .A(n6343), .B(n8216), .ZN(n8206) );
  NAND2_X1 U8009 ( .A1(n4314), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6344) );
  OAI21_X1 U8010 ( .B1(n4314), .B2(n8191), .A(n6344), .ZN(n6346) );
  INV_X1 U8011 ( .A(n6346), .ZN(n6345) );
  NAND2_X1 U8012 ( .A1(n8198), .A2(n6345), .ZN(n6394) );
  XNOR2_X1 U8013 ( .A(n6346), .B(n8198), .ZN(n8188) );
  NAND2_X1 U8014 ( .A1(n4314), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6347) );
  OAI21_X1 U8015 ( .B1(n4313), .B2(n6348), .A(n6347), .ZN(n6349) );
  OR2_X1 U8016 ( .A1(n6824), .A2(n6349), .ZN(n6393) );
  XNOR2_X1 U8017 ( .A(n6349), .B(n8181), .ZN(n8171) );
  NAND2_X1 U8018 ( .A1(n4314), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6350) );
  OAI21_X1 U8019 ( .B1(n4313), .B2(n6351), .A(n6350), .ZN(n6391) );
  OR2_X1 U8020 ( .A1(n6705), .A2(n6391), .ZN(n6392) );
  OR2_X1 U8021 ( .A1(n4314), .A2(n7609), .ZN(n6353) );
  NAND2_X1 U8022 ( .A1(n4314), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U8023 ( .A1(n6353), .A2(n6352), .ZN(n6383) );
  NOR2_X1 U8024 ( .A1(n6383), .A2(n7612), .ZN(n6385) );
  MUX2_X1 U8025 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n4313), .Z(n6380) );
  NOR2_X1 U8026 ( .A1(n6380), .A2(n7361), .ZN(n6382) );
  OR2_X1 U8027 ( .A1(n4314), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8028 ( .A1(n4313), .A2(n5939), .ZN(n6354) );
  NAND2_X1 U8029 ( .A1(n6355), .A2(n6354), .ZN(n6378) );
  NOR2_X1 U8030 ( .A1(n6378), .A2(n6377), .ZN(n7311) );
  INV_X1 U8031 ( .A(n7311), .ZN(n6379) );
  NAND2_X1 U8032 ( .A1(n4314), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6356) );
  OAI21_X1 U8033 ( .B1(n4314), .B2(n7374), .A(n6356), .ZN(n6375) );
  OR2_X1 U8034 ( .A1(n6375), .A2(n6604), .ZN(n6376) );
  MUX2_X1 U8035 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n4314), .Z(n6374) );
  XNOR2_X1 U8036 ( .A(n6374), .B(n9829), .ZN(n9837) );
  INV_X1 U8037 ( .A(n6990), .ZN(n6358) );
  MUX2_X1 U8038 ( .A(n7235), .B(n6357), .S(n4314), .Z(n6372) );
  NAND2_X1 U8039 ( .A1(n6358), .A2(n6372), .ZN(n6373) );
  MUX2_X1 U8040 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n4314), .Z(n6371) );
  MUX2_X1 U8041 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n4314), .Z(n6370) );
  MUX2_X1 U8042 ( .A(n6982), .B(n6359), .S(n4313), .Z(n6368) );
  INV_X1 U8043 ( .A(n6368), .ZN(n6369) );
  MUX2_X1 U8044 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6206), .Z(n6367) );
  OR2_X1 U8045 ( .A1(n6206), .A2(n9990), .ZN(n6361) );
  NAND2_X1 U8046 ( .A1(n6206), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U8047 ( .A1(n6361), .A2(n6360), .ZN(n6365) );
  XNOR2_X1 U8048 ( .A(n6365), .B(n6364), .ZN(n6657) );
  OR2_X1 U8049 ( .A1(n6206), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8050 ( .A1(n6206), .A2(n5835), .ZN(n6362) );
  NAND2_X1 U8051 ( .A1(n6363), .A2(n6362), .ZN(n6617) );
  NAND2_X1 U8052 ( .A1(n6657), .A2(n6656), .ZN(n6655) );
  INV_X1 U8053 ( .A(n6364), .ZN(n6665) );
  NAND2_X1 U8054 ( .A1(n6365), .A2(n6665), .ZN(n6366) );
  NAND2_X1 U8055 ( .A1(n6655), .A2(n6366), .ZN(n9802) );
  INV_X1 U8056 ( .A(n6588), .ZN(n9809) );
  XNOR2_X1 U8057 ( .A(n6367), .B(n9809), .ZN(n9803) );
  AND2_X1 U8058 ( .A1(n9802), .A2(n9803), .ZN(n9800) );
  XNOR2_X1 U8059 ( .A(n6368), .B(n6649), .ZN(n6638) );
  NAND2_X1 U8060 ( .A1(n6639), .A2(n6638), .ZN(n6637) );
  OAI21_X1 U8061 ( .B1(n6369), .B2(n6649), .A(n6637), .ZN(n6839) );
  XNOR2_X1 U8062 ( .A(n6370), .B(n6856), .ZN(n6840) );
  XNOR2_X1 U8063 ( .A(n6371), .B(n6585), .ZN(n6559) );
  XNOR2_X1 U8064 ( .A(n6372), .B(n6990), .ZN(n6987) );
  NAND2_X1 U8065 ( .A1(n6373), .A2(n6986), .ZN(n9836) );
  NAND2_X1 U8066 ( .A1(n9837), .A2(n9836), .ZN(n9835) );
  OAI21_X1 U8067 ( .B1(n6374), .B2(n6593), .A(n9835), .ZN(n7386) );
  XNOR2_X1 U8068 ( .A(n6375), .B(n7397), .ZN(n7387) );
  NAND2_X1 U8069 ( .A1(n7386), .A2(n7387), .ZN(n7385) );
  NAND2_X1 U8070 ( .A1(n6376), .A2(n7385), .ZN(n7313) );
  AND2_X1 U8071 ( .A1(n6378), .A2(n6377), .ZN(n7312) );
  AOI21_X1 U8072 ( .B1(n7361), .B2(n6380), .A(n6382), .ZN(n6381) );
  INV_X1 U8073 ( .A(n6381), .ZN(n7349) );
  AND2_X1 U8074 ( .A1(n6383), .A2(n7612), .ZN(n6384) );
  OR2_X1 U8075 ( .A1(n6385), .A2(n6384), .ZN(n7616) );
  NAND2_X1 U8076 ( .A1(n8098), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6386) );
  OAI211_X1 U8077 ( .C1(n8098), .C2(n6388), .A(n6387), .B(n6386), .ZN(n8129)
         );
  OR2_X1 U8078 ( .A1(n4313), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6390) );
  AOI21_X1 U8079 ( .B1(n4313), .B2(n6388), .A(n6387), .ZN(n6389) );
  AND2_X1 U8080 ( .A1(n6390), .A2(n6389), .ZN(n8128) );
  AOI21_X1 U8081 ( .B1(n8132), .B2(n8129), .A(n8128), .ZN(n8162) );
  XNOR2_X1 U8082 ( .A(n6391), .B(n8159), .ZN(n8161) );
  NAND2_X1 U8083 ( .A1(n8171), .A2(n8170), .ZN(n8169) );
  NAND2_X1 U8084 ( .A1(n6393), .A2(n8169), .ZN(n8187) );
  NAND2_X1 U8085 ( .A1(n8188), .A2(n8187), .ZN(n8186) );
  NAND2_X1 U8086 ( .A1(n6394), .A2(n8186), .ZN(n8205) );
  NAND2_X1 U8087 ( .A1(n8206), .A2(n8205), .ZN(n8204) );
  NAND2_X1 U8088 ( .A1(n6395), .A2(n8204), .ZN(n8223) );
  NAND2_X1 U8089 ( .A1(n8224), .A2(n8223), .ZN(n8222) );
  NAND2_X1 U8090 ( .A1(n4314), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6397) );
  OAI21_X1 U8091 ( .B1(n6206), .B2(n8364), .A(n6397), .ZN(n6400) );
  NAND2_X1 U8092 ( .A1(n6399), .A2(n6400), .ZN(n8245) );
  NAND2_X1 U8093 ( .A1(n8245), .A2(n6398), .ZN(n6403) );
  INV_X1 U8094 ( .A(n6399), .ZN(n6402) );
  INV_X1 U8095 ( .A(n6400), .ZN(n6401) );
  NAND2_X1 U8096 ( .A1(n6402), .A2(n6401), .ZN(n8244) );
  NAND2_X1 U8097 ( .A1(n6403), .A2(n8244), .ZN(n6407) );
  MUX2_X1 U8098 ( .A(n6405), .B(n6404), .S(n8098), .Z(n6406) );
  XNOR2_X1 U8099 ( .A(n6407), .B(n6406), .ZN(n6411) );
  NAND2_X1 U8100 ( .A1(P2_U3893), .A2(n6205), .ZN(n8249) );
  INV_X1 U8101 ( .A(n7458), .ZN(n6408) );
  NOR2_X1 U8102 ( .A1(n6542), .A2(n6408), .ZN(n6409) );
  AND2_X1 U8103 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6535) );
  AOI21_X1 U8104 ( .B1(n9840), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n6535), .ZN(
        n6410) );
  OAI21_X1 U8105 ( .B1(n6411), .B2(n8249), .A(n6410), .ZN(n6416) );
  NOR2_X1 U8106 ( .A1(n6206), .A2(P2_U3151), .ZN(n7556) );
  NAND2_X1 U8107 ( .A1(n6412), .A2(n7556), .ZN(n6414) );
  MUX2_X1 U8108 ( .A(n6414), .B(n8248), .S(n6413), .Z(n8246) );
  NOR2_X1 U8109 ( .A1(n8246), .A2(n7231), .ZN(n6415) );
  NOR2_X1 U8110 ( .A1(n6417), .A2(n8574), .ZN(n6828) );
  NAND2_X1 U8111 ( .A1(n7347), .A2(n6418), .ZN(n6455) );
  OR2_X1 U8112 ( .A1(n6419), .A2(n6455), .ZN(n6545) );
  NOR2_X1 U8113 ( .A1(n9900), .A2(n8085), .ZN(n6420) );
  NAND2_X1 U8114 ( .A1(n6545), .A2(n6420), .ZN(n6523) );
  NAND2_X1 U8115 ( .A1(n6421), .A2(n9900), .ZN(n8413) );
  NAND2_X1 U8116 ( .A1(n6523), .A2(n8413), .ZN(n6538) );
  NAND2_X1 U8117 ( .A1(n6533), .A2(n6538), .ZN(n6425) );
  NAND2_X1 U8118 ( .A1(n6537), .A2(n8573), .ZN(n6422) );
  NOR2_X1 U8119 ( .A1(n6540), .A2(n6422), .ZN(n6529) );
  NAND2_X1 U8120 ( .A1(n6532), .A2(n6545), .ZN(n6423) );
  NAND2_X1 U8121 ( .A1(n6529), .A2(n6423), .ZN(n6424) );
  INV_X1 U8122 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U8123 ( .A1(n9906), .A2(n6426), .ZN(n6427) );
  NAND2_X1 U8124 ( .A1(n6429), .A2(n4925), .ZN(P2_U3455) );
  INV_X1 U8125 ( .A(n6432), .ZN(n6433) );
  OAI21_X1 U8126 ( .B1(n6434), .B2(n6433), .A(n8748), .ZN(n6438) );
  AOI22_X1 U8127 ( .A1(n8757), .A2(n9242), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6435) );
  OAI21_X1 U8128 ( .B1(n9408), .B2(n8759), .A(n6435), .ZN(n6436) );
  AOI21_X1 U8129 ( .B1(n9212), .B2(n8763), .A(n6436), .ZN(n6437) );
  INV_X1 U8130 ( .A(n9411), .ZN(n9216) );
  NAND3_X1 U8131 ( .A1(n6438), .A2(n6437), .A3(n4915), .ZN(P1_U3214) );
  NAND2_X1 U8132 ( .A1(n8063), .A2(n8064), .ZN(n8067) );
  XNOR2_X1 U8133 ( .A(n6441), .B(n8067), .ZN(n8268) );
  INV_X1 U8134 ( .A(n8067), .ZN(n6442) );
  AOI21_X1 U8135 ( .B1(n6266), .B2(n8268), .A(n8263), .ZN(n6450) );
  MUX2_X1 U8136 ( .A(n6448), .B(n6450), .S(n9905), .Z(n6449) );
  NAND2_X1 U8137 ( .A1(n6449), .A2(n4914), .ZN(P2_U3454) );
  INV_X1 U8138 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6451) );
  MUX2_X1 U8139 ( .A(n6451), .B(n6450), .S(n9920), .Z(n6452) );
  NAND2_X1 U8140 ( .A1(n6452), .A2(n4913), .ZN(P2_U3486) );
  AND2_X2 U8141 ( .A1(n6454), .A2(n6453), .ZN(P1_U3973) );
  INV_X1 U8142 ( .A(n6455), .ZN(n6456) );
  XNOR2_X1 U8143 ( .A(n8351), .B(n7774), .ZN(n7734) );
  XNOR2_X1 U8144 ( .A(n7734), .B(n8360), .ZN(n6528) );
  XNOR2_X1 U8145 ( .A(n6460), .B(n4318), .ZN(n6461) );
  NAND2_X1 U8146 ( .A1(n6461), .A2(n5834), .ZN(n6465) );
  INV_X1 U8147 ( .A(n6461), .ZN(n6462) );
  NAND2_X1 U8148 ( .A1(n6462), .A2(n5842), .ZN(n6463) );
  XNOR2_X1 U8149 ( .A(n7774), .B(n9855), .ZN(n6467) );
  INV_X1 U8150 ( .A(n8126), .ZN(n6466) );
  XNOR2_X1 U8151 ( .A(n6467), .B(n6466), .ZN(n6784) );
  OR2_X1 U8152 ( .A1(n6467), .A2(n8126), .ZN(n6468) );
  INV_X1 U8153 ( .A(n6893), .ZN(n6470) );
  XNOR2_X1 U8154 ( .A(n7774), .B(n9860), .ZN(n6471) );
  XNOR2_X1 U8155 ( .A(n6471), .B(n5867), .ZN(n6894) );
  NAND2_X1 U8156 ( .A1(n6471), .A2(n5867), .ZN(n6472) );
  XNOR2_X1 U8157 ( .A(n7749), .B(n9867), .ZN(n6473) );
  NAND2_X1 U8158 ( .A1(n6473), .A2(n7160), .ZN(n7071) );
  INV_X1 U8159 ( .A(n6473), .ZN(n6474) );
  NAND2_X1 U8160 ( .A1(n8125), .A2(n6474), .ZN(n6475) );
  NAND2_X1 U8161 ( .A1(n7071), .A2(n6475), .ZN(n6963) );
  NAND2_X1 U8162 ( .A1(n7073), .A2(n7071), .ZN(n6477) );
  XNOR2_X1 U8163 ( .A(n4319), .B(n7078), .ZN(n6478) );
  XNOR2_X1 U8164 ( .A(n6478), .B(n8124), .ZN(n7070) );
  NAND2_X1 U8165 ( .A1(n6477), .A2(n7070), .ZN(n7075) );
  INV_X1 U8166 ( .A(n8124), .ZN(n7223) );
  NAND2_X1 U8167 ( .A1(n6478), .A2(n7223), .ZN(n6479) );
  INV_X1 U8168 ( .A(n7221), .ZN(n6481) );
  XNOR2_X1 U8169 ( .A(n7238), .B(n7774), .ZN(n6482) );
  INV_X1 U8170 ( .A(n8432), .ZN(n7671) );
  XNOR2_X1 U8171 ( .A(n6482), .B(n7671), .ZN(n7222) );
  INV_X1 U8172 ( .A(n6482), .ZN(n6483) );
  NAND2_X1 U8173 ( .A1(n6483), .A2(n8432), .ZN(n6484) );
  XNOR2_X1 U8174 ( .A(n4319), .B(n9882), .ZN(n6485) );
  INV_X1 U8175 ( .A(n8123), .ZN(n7444) );
  XNOR2_X1 U8176 ( .A(n6485), .B(n7444), .ZN(n7668) );
  OR2_X1 U8177 ( .A1(n6485), .A2(n8123), .ZN(n6486) );
  XNOR2_X1 U8178 ( .A(n7541), .B(n7749), .ZN(n7546) );
  NAND2_X1 U8179 ( .A1(n7546), .A2(n8122), .ZN(n7573) );
  XNOR2_X1 U8180 ( .A(n9888), .B(n7774), .ZN(n6489) );
  NAND2_X1 U8181 ( .A1(n6489), .A2(n8431), .ZN(n6487) );
  AND2_X1 U8182 ( .A1(n7573), .A2(n6487), .ZN(n6488) );
  XNOR2_X1 U8183 ( .A(n9899), .B(n4319), .ZN(n7575) );
  NAND2_X1 U8184 ( .A1(n7575), .A2(n7549), .ZN(n6491) );
  INV_X1 U8185 ( .A(n8431), .ZN(n7426) );
  INV_X1 U8186 ( .A(n6489), .ZN(n7543) );
  NAND3_X1 U8187 ( .A1(n7573), .A2(n7426), .A3(n7543), .ZN(n6490) );
  OAI211_X1 U8188 ( .C1(n7546), .C2(n8122), .A(n6491), .B(n6490), .ZN(n6492)
         );
  INV_X1 U8189 ( .A(n6492), .ZN(n6493) );
  NAND2_X1 U8190 ( .A1(n6494), .A2(n6493), .ZN(n6497) );
  INV_X1 U8191 ( .A(n7575), .ZN(n6495) );
  NAND2_X1 U8192 ( .A1(n6495), .A2(n8121), .ZN(n6496) );
  XNOR2_X1 U8193 ( .A(n7916), .B(n7749), .ZN(n7437) );
  NAND2_X1 U8194 ( .A1(n7437), .A2(n8120), .ZN(n6499) );
  XNOR2_X1 U8195 ( .A(n8509), .B(n7774), .ZN(n6500) );
  NAND2_X1 U8196 ( .A1(n6500), .A2(n7994), .ZN(n7523) );
  INV_X1 U8197 ( .A(n6500), .ZN(n6501) );
  NAND2_X1 U8198 ( .A1(n6501), .A2(n8119), .ZN(n7524) );
  XNOR2_X1 U8199 ( .A(n7599), .B(n7749), .ZN(n7534) );
  INV_X1 U8200 ( .A(n7534), .ZN(n6502) );
  NAND2_X1 U8201 ( .A1(n6502), .A2(n7629), .ZN(n6504) );
  AND2_X1 U8202 ( .A1(n7534), .A2(n8409), .ZN(n6503) );
  XNOR2_X1 U8203 ( .A(n8500), .B(n7774), .ZN(n6505) );
  XNOR2_X1 U8204 ( .A(n6505), .B(n8118), .ZN(n7626) );
  NAND2_X1 U8205 ( .A1(n6505), .A2(n7660), .ZN(n6506) );
  XNOR2_X1 U8206 ( .A(n7645), .B(n4319), .ZN(n6508) );
  XNOR2_X1 U8207 ( .A(n6508), .B(n8389), .ZN(n7646) );
  INV_X1 U8208 ( .A(n7646), .ZN(n6507) );
  INV_X1 U8209 ( .A(n6508), .ZN(n6509) );
  NAND2_X1 U8210 ( .A1(n6509), .A2(n8410), .ZN(n6510) );
  XNOR2_X1 U8211 ( .A(n8395), .B(n4319), .ZN(n6511) );
  XNOR2_X1 U8212 ( .A(n6511), .B(n8117), .ZN(n7809) );
  NAND2_X1 U8213 ( .A1(n7810), .A2(n7809), .ZN(n6514) );
  INV_X1 U8214 ( .A(n6511), .ZN(n6512) );
  NAND2_X1 U8215 ( .A1(n6512), .A2(n8117), .ZN(n6513) );
  XNOR2_X1 U8216 ( .A(n8383), .B(n7774), .ZN(n6515) );
  INV_X1 U8217 ( .A(n6515), .ZN(n6516) );
  INV_X1 U8218 ( .A(n8391), .ZN(n8116) );
  NAND2_X1 U8219 ( .A1(n6516), .A2(n8116), .ZN(n6517) );
  NAND2_X1 U8220 ( .A1(n7851), .A2(n6517), .ZN(n7817) );
  XNOR2_X1 U8221 ( .A(n8556), .B(n4319), .ZN(n6519) );
  XNOR2_X1 U8222 ( .A(n6519), .B(n8375), .ZN(n7852) );
  INV_X1 U8223 ( .A(n6519), .ZN(n6520) );
  NAND2_X1 U8224 ( .A1(n6520), .A2(n8375), .ZN(n6521) );
  INV_X1 U8225 ( .A(n6545), .ZN(n6522) );
  NAND2_X1 U8226 ( .A1(n6533), .A2(n6522), .ZN(n6526) );
  INV_X1 U8227 ( .A(n6523), .ZN(n6524) );
  NAND2_X1 U8228 ( .A1(n6529), .A2(n6524), .ZN(n6525) );
  INV_X1 U8229 ( .A(n7737), .ZN(n7834) );
  AOI211_X1 U8230 ( .C1(n6528), .C2(n6527), .A(n7879), .B(n7834), .ZN(n6557)
         );
  NAND2_X1 U8231 ( .A1(n6529), .A2(n9900), .ZN(n6531) );
  AND2_X1 U8232 ( .A1(n8351), .A2(n7876), .ZN(n6556) );
  INV_X1 U8233 ( .A(n6532), .ZN(n6547) );
  NAND2_X1 U8234 ( .A1(n6533), .A2(n6547), .ZN(n6552) );
  INV_X1 U8235 ( .A(n6535), .ZN(n6536) );
  OAI21_X1 U8236 ( .B1(n7874), .B2(n8346), .A(n6536), .ZN(n6555) );
  INV_X1 U8237 ( .A(n8352), .ZN(n6553) );
  INV_X1 U8238 ( .A(n6537), .ZN(n6539) );
  OAI21_X1 U8239 ( .B1(n6540), .B2(n6539), .A(n6538), .ZN(n6543) );
  AND4_X1 U8240 ( .A1(n6543), .A2(n6542), .A3(n7458), .A4(n6541), .ZN(n6544)
         );
  OAI21_X1 U8241 ( .B1(n6548), .B2(n6545), .A(n6544), .ZN(n6546) );
  NAND2_X1 U8242 ( .A1(n6546), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6550) );
  NAND2_X1 U8243 ( .A1(n8573), .A2(n6547), .ZN(n8099) );
  OR2_X1 U8244 ( .A1(n6548), .A2(n8099), .ZN(n6549) );
  OAI22_X1 U8245 ( .A1(n6553), .A2(n7861), .B1(n7860), .B2(n8375), .ZN(n6554)
         );
  OR4_X1 U8246 ( .A1(n6557), .A2(n6556), .A3(n6555), .A4(n6554), .ZN(P2_U3159)
         );
  AOI211_X1 U8247 ( .C1(n6560), .C2(n6559), .A(n8249), .B(n6558), .ZN(n6571)
         );
  NOR2_X1 U8248 ( .A1(n8246), .A2(n6585), .ZN(n6570) );
  AOI21_X1 U8249 ( .B1(n7161), .B2(n6562), .A(n6561), .ZN(n6563) );
  NAND2_X1 U8250 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7076) );
  OAI21_X1 U8251 ( .B1(n6563), .B2(n9832), .A(n7076), .ZN(n6569) );
  AOI21_X1 U8252 ( .B1(n5881), .B2(n6565), .A(n6564), .ZN(n6567) );
  INV_X1 U8253 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6566) );
  OAI22_X1 U8254 ( .A1(n6567), .A2(n9825), .B1(n8255), .B2(n6566), .ZN(n6568)
         );
  OR4_X1 U8255 ( .A1(n6571), .A2(n6570), .A3(n6569), .A4(n6568), .ZN(P2_U3187)
         );
  AND2_X1 U8256 ( .A1(n4586), .A2(P1_U3086), .ZN(n7106) );
  INV_X1 U8257 ( .A(n7106), .ZN(n7522) );
  NOR2_X1 U8258 ( .A1(n4586), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9568) );
  OAI222_X1 U8259 ( .A1(n7522), .A2(n4611), .B1(n7708), .B2(n6575), .C1(n6726), 
        .C2(P1_U3086), .ZN(P1_U3354) );
  OAI222_X1 U8260 ( .A1(n9054), .A2(P1_U3086), .B1(n7708), .B2(n6581), .C1(
        n6572), .C2(n7522), .ZN(P1_U3352) );
  OAI222_X1 U8261 ( .A1(n6747), .A2(P1_U3086), .B1(n7708), .B2(n6589), .C1(
        n6573), .C2(n7522), .ZN(P1_U3353) );
  NAND2_X1 U8262 ( .A1(n6574), .A2(P2_U3151), .ZN(n7728) );
  INV_X1 U8263 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6576) );
  AND2_X1 U8264 ( .A1(n4586), .A2(P2_U3151), .ZN(n8581) );
  INV_X2 U8265 ( .A(n8581), .ZN(n7730) );
  OAI222_X1 U8266 ( .A1(n7728), .A2(n6576), .B1(n7730), .B2(n6575), .C1(
        P2_U3151), .C2(n6665), .ZN(P2_U3294) );
  INV_X1 U8267 ( .A(n6804), .ZN(n6578) );
  OAI222_X1 U8268 ( .A1(n6578), .A2(P1_U3086), .B1(n7708), .B2(n6583), .C1(
        n6577), .C2(n7522), .ZN(P1_U3351) );
  INV_X1 U8269 ( .A(n9075), .ZN(n6580) );
  OAI222_X1 U8270 ( .A1(n6580), .A2(P1_U3086), .B1(n7708), .B2(n6586), .C1(
        n6579), .C2(n7522), .ZN(P1_U3350) );
  INV_X1 U8271 ( .A(n7728), .ZN(n7587) );
  INV_X1 U8272 ( .A(n7587), .ZN(n8577) );
  OAI222_X1 U8273 ( .A1(n8577), .A2(n6582), .B1(n7730), .B2(n6581), .C1(
        P2_U3151), .C2(n6649), .ZN(P2_U3292) );
  OAI222_X1 U8274 ( .A1(n8577), .A2(n6584), .B1(n7730), .B2(n6583), .C1(
        P2_U3151), .C2(n6856), .ZN(P2_U3291) );
  OAI222_X1 U8275 ( .A1(n8577), .A2(n6587), .B1(n7730), .B2(n6586), .C1(
        P2_U3151), .C2(n6585), .ZN(P2_U3290) );
  OAI222_X1 U8276 ( .A1(n8577), .A2(n4732), .B1(n7730), .B2(n6589), .C1(
        P2_U3151), .C2(n6588), .ZN(P2_U3293) );
  AOI22_X1 U8277 ( .A1(n9089), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n7106), .ZN(n6590) );
  OAI21_X1 U8278 ( .B1(n6591), .B2(n7708), .A(n6590), .ZN(P1_U3349) );
  OAI222_X1 U8279 ( .A1(n8577), .A2(n9991), .B1(n7730), .B2(n6591), .C1(
        P2_U3151), .C2(n6990), .ZN(P2_U3289) );
  AOI22_X1 U8280 ( .A1(n9597), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n7106), .ZN(n6592) );
  OAI21_X1 U8281 ( .B1(n6594), .B2(n7708), .A(n6592), .ZN(P1_U3348) );
  OAI222_X1 U8282 ( .A1(n8577), .A2(n6595), .B1(n7730), .B2(n6594), .C1(
        P2_U3151), .C2(n6593), .ZN(P2_U3288) );
  NAND2_X1 U8283 ( .A1(n9745), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6597) );
  OAI21_X1 U8284 ( .B1(n9745), .B2(n6598), .A(n6597), .ZN(P1_U3439) );
  INV_X1 U8285 ( .A(n6599), .ZN(n6605) );
  AOI22_X1 U8286 ( .A1(n9609), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7106), .ZN(n6600) );
  OAI21_X1 U8287 ( .B1(n6605), .B2(n7708), .A(n6600), .ZN(P1_U3347) );
  NAND2_X1 U8288 ( .A1(n8573), .A2(n6233), .ZN(n9946) );
  AOI22_X1 U8289 ( .A1(n9946), .A2(n4428), .B1(n6601), .B2(n4426), .ZN(
        P2_U3376) );
  AND2_X1 U8290 ( .A1(n9946), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8291 ( .A1(n9946), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8292 ( .A1(n9946), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8293 ( .A1(n9946), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8294 ( .A1(n9946), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8295 ( .A1(n9946), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8296 ( .A1(n9946), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8297 ( .A1(n9946), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8298 ( .A1(n9946), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8299 ( .A1(n9946), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8300 ( .A1(n9946), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8301 ( .A1(n9946), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8302 ( .A1(n9946), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8303 ( .A1(n9946), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8304 ( .A1(n9946), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8305 ( .A1(n9946), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8306 ( .A1(n9946), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8307 ( .A1(n9946), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8308 ( .A1(n9946), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8309 ( .A1(n9946), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8310 ( .A1(n9946), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8311 ( .A1(n9946), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8312 ( .A1(n9946), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  NAND2_X1 U8313 ( .A1(n6632), .A2(n9024), .ZN(n6722) );
  AOI21_X1 U8314 ( .B1(n9002), .B2(n6602), .A(n5086), .ZN(n6721) );
  INV_X1 U8315 ( .A(n6721), .ZN(n6603) );
  AND2_X1 U8316 ( .A1(n6722), .A2(n6603), .ZN(n9616) );
  NOR2_X1 U8317 ( .A1(n9616), .A2(P1_U3973), .ZN(P1_U3085) );
  OAI222_X1 U8318 ( .A1(n8577), .A2(n6606), .B1(n7730), .B2(n6605), .C1(
        P2_U3151), .C2(n6604), .ZN(P2_U3287) );
  INV_X1 U8319 ( .A(n9946), .ZN(n6607) );
  INV_X1 U8320 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10008) );
  NOR2_X1 U8321 ( .A1(n6607), .A2(n10008), .ZN(P2_U3234) );
  INV_X1 U8322 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10071) );
  NOR2_X1 U8323 ( .A1(n6607), .A2(n10071), .ZN(P2_U3255) );
  INV_X1 U8324 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10007) );
  NOR2_X1 U8325 ( .A1(n6607), .A2(n10007), .ZN(P2_U3235) );
  INV_X1 U8326 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10068) );
  NOR2_X1 U8327 ( .A1(n6607), .A2(n10068), .ZN(P2_U3248) );
  INV_X1 U8328 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9997) );
  NOR2_X1 U8329 ( .A1(n6607), .A2(n9997), .ZN(P2_U3245) );
  INV_X1 U8330 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10081) );
  NOR2_X1 U8331 ( .A1(n6607), .A2(n10081), .ZN(P2_U3256) );
  INV_X1 U8332 ( .A(n6608), .ZN(n6611) );
  AOI22_X1 U8333 ( .A1(n9105), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n7106), .ZN(n6609) );
  OAI21_X1 U8334 ( .B1(n6611), .B2(n7708), .A(n6609), .ZN(P1_U3346) );
  OAI222_X1 U8335 ( .A1(n7730), .A2(n6611), .B1(n7323), .B2(P2_U3151), .C1(
        n6610), .C2(n8577), .ZN(P2_U3286) );
  INV_X1 U8336 ( .A(n6612), .ZN(n6615) );
  AOI22_X1 U8337 ( .A1(n9583), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7106), .ZN(n6613) );
  OAI21_X1 U8338 ( .B1(n6615), .B2(n7708), .A(n6613), .ZN(P1_U3345) );
  OAI222_X1 U8339 ( .A1(n7730), .A2(n6615), .B1(n7361), .B2(P2_U3151), .C1(
        n6614), .C2(n8577), .ZN(P2_U3285) );
  INV_X1 U8340 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6622) );
  NAND2_X1 U8341 ( .A1(n6616), .A2(n8249), .ZN(n6619) );
  AOI22_X1 U8342 ( .A1(n6619), .A2(n6618), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6621) );
  OAI211_X1 U8343 ( .C1(n8255), .C2(n6622), .A(n6621), .B(n6620), .ZN(P2_U3182) );
  INV_X1 U8344 ( .A(n6623), .ZN(n6626) );
  OAI222_X1 U8345 ( .A1(n7728), .A2(n6624), .B1(n7730), .B2(n6626), .C1(
        P2_U3151), .C2(n7612), .ZN(P2_U3284) );
  INV_X1 U8346 ( .A(n6813), .ZN(n9630) );
  OAI222_X1 U8347 ( .A1(n9630), .A2(P1_U3086), .B1(n7708), .B2(n6626), .C1(
        n6625), .C2(n7522), .ZN(P1_U3344) );
  INV_X1 U8348 ( .A(n6627), .ZN(n6628) );
  AOI21_X1 U8349 ( .B1(n6630), .B2(n6629), .A(n6628), .ZN(n6636) );
  AOI22_X1 U8350 ( .A1(n8726), .A2(n9040), .B1(n8757), .B2(n9042), .ZN(n6635)
         );
  OR2_X1 U8351 ( .A1(n6633), .A2(n6632), .ZN(n7698) );
  AOI22_X1 U8352 ( .A1(n8741), .A2(n6692), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n7698), .ZN(n6634) );
  OAI211_X1 U8353 ( .C1(n6636), .C2(n8766), .A(n6635), .B(n6634), .ZN(P1_U3222) );
  OAI21_X1 U8354 ( .B1(n6639), .B2(n6638), .A(n6637), .ZN(n6640) );
  NAND2_X1 U8355 ( .A1(n6640), .A2(n9838), .ZN(n6648) );
  INV_X1 U8356 ( .A(n9825), .ZN(n9808) );
  OAI21_X1 U8357 ( .B1(n6641), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6844), .ZN(
        n6642) );
  AOI22_X1 U8358 ( .A1(n9840), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(n9808), .B2(
        n6642), .ZN(n6646) );
  NAND2_X1 U8359 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6896) );
  OAI21_X1 U8360 ( .B1(n6643), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6848), .ZN(
        n6644) );
  NAND2_X1 U8361 ( .A1(n9816), .A2(n6644), .ZN(n6645) );
  AND3_X1 U8362 ( .A1(n6646), .A2(n6896), .A3(n6645), .ZN(n6647) );
  OAI211_X1 U8363 ( .C1(n8246), .C2(n6649), .A(n6648), .B(n6647), .ZN(P2_U3185) );
  INV_X1 U8364 ( .A(n6650), .ZN(n6666) );
  OAI222_X1 U8365 ( .A1(n7730), .A2(n6666), .B1(n8146), .B2(P2_U3151), .C1(
        n6651), .C2(n8577), .ZN(P2_U3283) );
  INV_X1 U8366 ( .A(n6652), .ZN(n6653) );
  AOI21_X1 U8367 ( .B1(n5822), .B2(n6654), .A(n6653), .ZN(n6659) );
  OAI211_X1 U8368 ( .C1(n6657), .C2(n6656), .A(n9838), .B(n6655), .ZN(n6658)
         );
  OAI21_X1 U8369 ( .B1(n6659), .B2(n9825), .A(n6658), .ZN(n6663) );
  XOR2_X1 U8370 ( .A(n9990), .B(n6660), .Z(n6661) );
  OAI22_X1 U8371 ( .A1(n9832), .A2(n6661), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6677), .ZN(n6662) );
  AOI211_X1 U8372 ( .C1(n9840), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6663), .B(
        n6662), .ZN(n6664) );
  OAI21_X1 U8373 ( .B1(n6665), .B2(n8246), .A(n6664), .ZN(P2_U3183) );
  INV_X1 U8374 ( .A(n9123), .ZN(n6818) );
  OAI222_X1 U8375 ( .A1(n7522), .A2(n6667), .B1(P1_U3086), .B2(n6818), .C1(
        n6666), .C2(n7708), .ZN(P1_U3343) );
  INV_X1 U8376 ( .A(n6668), .ZN(n6706) );
  AOI22_X1 U8377 ( .A1(n9644), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7106), .ZN(n6669) );
  OAI21_X1 U8378 ( .B1(n6706), .B2(n7708), .A(n6669), .ZN(P1_U3342) );
  NOR2_X1 U8379 ( .A1(n7871), .A2(P2_U3151), .ZN(n6789) );
  INV_X1 U8380 ( .A(n7876), .ZN(n7867) );
  OAI22_X1 U8381 ( .A1(n7860), .A2(n4482), .B1(n7867), .B2(n9850), .ZN(n6670)
         );
  AOI21_X1 U8382 ( .B1(n7864), .B2(n8126), .A(n6670), .ZN(n6676) );
  OAI21_X1 U8383 ( .B1(n6673), .B2(n6672), .A(n6671), .ZN(n6674) );
  NAND2_X1 U8384 ( .A1(n6674), .A2(n7856), .ZN(n6675) );
  OAI211_X1 U8385 ( .C1(n6789), .C2(n6677), .A(n6676), .B(n6675), .ZN(P2_U3162) );
  NAND2_X1 U8386 ( .A1(n8127), .A2(n6926), .ZN(n7939) );
  NAND2_X1 U8387 ( .A1(n7935), .A2(n7939), .ZN(n7905) );
  AOI22_X1 U8388 ( .A1(n7856), .A2(n7905), .B1(n9848), .B2(n7876), .ZN(n6679)
         );
  NAND2_X1 U8389 ( .A1(n7864), .A2(n5842), .ZN(n6678) );
  OAI211_X1 U8390 ( .C1(n6789), .C2(n6680), .A(n6679), .B(n6678), .ZN(P2_U3172) );
  INV_X1 U8391 ( .A(n6777), .ZN(n7010) );
  AND3_X1 U8392 ( .A1(n9009), .A2(n6681), .A3(n7007), .ZN(n6682) );
  AND2_X2 U8393 ( .A1(n7010), .A2(n6778), .ZN(n9789) );
  INV_X1 U8394 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U8395 ( .A1(n9042), .A2(n7688), .ZN(n6686) );
  NAND2_X1 U8396 ( .A1(n6685), .A2(n6686), .ZN(n6769) );
  OAI21_X1 U8397 ( .B1(n6685), .B2(n6686), .A(n6769), .ZN(n7066) );
  OR2_X1 U8398 ( .A1(n6687), .A2(n6689), .ZN(n7682) );
  INV_X1 U8399 ( .A(n6688), .ZN(n7681) );
  NAND2_X1 U8400 ( .A1(n6690), .A2(n6689), .ZN(n6691) );
  NAND3_X1 U8401 ( .A1(n7682), .A2(n7681), .A3(n6691), .ZN(n7083) );
  OR2_X1 U8402 ( .A1(n9016), .A2(n5736), .ZN(n9769) );
  AOI22_X1 U8403 ( .A1(n9042), .A2(n9474), .B1(n6692), .B2(n9762), .ZN(n6694)
         );
  INV_X1 U8404 ( .A(n7688), .ZN(n6703) );
  OAI211_X1 U8405 ( .C1(n6703), .C2(n6693), .A(n9452), .B(n7039), .ZN(n7061)
         );
  OAI211_X1 U8406 ( .C1(n6631), .C2(n9530), .A(n6694), .B(n7061), .ZN(n6695)
         );
  AOI21_X1 U8407 ( .B1(n7066), .B2(n9786), .A(n6695), .ZN(n6697) );
  NOR2_X1 U8408 ( .A1(n9042), .A2(n6703), .ZN(n6764) );
  INV_X1 U8409 ( .A(n6764), .ZN(n6700) );
  XNOR2_X1 U8410 ( .A(n6700), .B(n6685), .ZN(n6696) );
  NAND2_X1 U8411 ( .A1(n5732), .A2(n9136), .ZN(n8946) );
  NAND2_X1 U8412 ( .A1(n8957), .A2(n5736), .ZN(n9017) );
  NAND2_X1 U8413 ( .A1(n6696), .A2(n9481), .ZN(n7069) );
  NAND2_X1 U8414 ( .A1(n6697), .A2(n7069), .ZN(n9540) );
  NAND2_X1 U8415 ( .A1(n9540), .A2(n9789), .ZN(n6698) );
  OAI21_X1 U8416 ( .B1(n9789), .B2(n6699), .A(n6698), .ZN(P1_U3456) );
  INV_X1 U8417 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U8418 ( .A1(n9042), .A2(n6703), .ZN(n8803) );
  NAND2_X1 U8419 ( .A1(n6700), .A2(n8803), .ZN(n8955) );
  INV_X1 U8420 ( .A(n8955), .ZN(n6702) );
  NOR2_X1 U8421 ( .A1(n9786), .A2(n9481), .ZN(n6701) );
  OAI222_X1 U8422 ( .A1(n6703), .A2(n7681), .B1(n6702), .B2(n6701), .C1(n9530), 
        .C2(n7687), .ZN(n9541) );
  NAND2_X1 U8423 ( .A1(n9541), .A2(n9789), .ZN(n6704) );
  OAI21_X1 U8424 ( .B1(n9789), .B2(n10041), .A(n6704), .ZN(P1_U3453) );
  INV_X1 U8425 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6707) );
  OAI222_X1 U8426 ( .A1(n7728), .A2(n6707), .B1(n7730), .B2(n6706), .C1(
        P2_U3151), .C2(n6705), .ZN(P2_U3282) );
  XOR2_X1 U8427 ( .A(n6709), .B(n6708), .Z(n7689) );
  INV_X1 U8428 ( .A(n7689), .ZN(n6712) );
  INV_X1 U8429 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6710) );
  INV_X1 U8430 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7680) );
  NOR2_X1 U8431 ( .A1(n6710), .A2(n7680), .ZN(n9047) );
  INV_X1 U8432 ( .A(n6711), .ZN(n9614) );
  MUX2_X1 U8433 ( .A(n6712), .B(n9047), .S(n9614), .Z(n6714) );
  INV_X1 U8434 ( .A(n5740), .ZN(n6735) );
  AOI21_X1 U8435 ( .B1(n9614), .B2(n7680), .A(n5740), .ZN(n9613) );
  OAI21_X1 U8436 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n9613), .A(P1_U3973), .ZN(
        n6713) );
  AOI21_X1 U8437 ( .B1(n6714), .B2(n6735), .A(n6713), .ZN(n6754) );
  INV_X1 U8438 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6715) );
  XNOR2_X1 U8439 ( .A(n6804), .B(n6715), .ZN(n6724) );
  XNOR2_X1 U8440 ( .A(n6747), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6746) );
  XNOR2_X1 U8441 ( .A(n6726), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9045) );
  AND2_X1 U8442 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9044) );
  NAND2_X1 U8443 ( .A1(n9045), .A2(n9044), .ZN(n9043) );
  NAND2_X1 U8444 ( .A1(n9049), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6716) );
  NAND2_X1 U8445 ( .A1(n9043), .A2(n6716), .ZN(n6745) );
  NAND2_X1 U8446 ( .A1(n6746), .A2(n6745), .ZN(n6744) );
  INV_X1 U8447 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6717) );
  OR2_X1 U8448 ( .A1(n6747), .A2(n6717), .ZN(n6718) );
  NAND2_X1 U8449 ( .A1(n6744), .A2(n6718), .ZN(n9063) );
  XNOR2_X1 U8450 ( .A(n9054), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U8451 ( .A1(n9063), .A2(n9064), .ZN(n9062) );
  INV_X1 U8452 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6719) );
  OR2_X1 U8453 ( .A1(n9054), .A2(n6719), .ZN(n6720) );
  NAND2_X1 U8454 ( .A1(n9062), .A2(n6720), .ZN(n6723) );
  NAND2_X1 U8455 ( .A1(n6722), .A2(n6721), .ZN(n9618) );
  NAND2_X1 U8456 ( .A1(n6723), .A2(n6724), .ZN(n6806) );
  OAI211_X1 U8457 ( .C1(n6724), .C2(n6723), .A(n9696), .B(n6806), .ZN(n6739)
         );
  INV_X1 U8458 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6725) );
  XNOR2_X1 U8459 ( .A(n6804), .B(n6725), .ZN(n6734) );
  XNOR2_X1 U8460 ( .A(n6747), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6743) );
  XNOR2_X1 U8461 ( .A(n6726), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U8462 ( .A1(n9048), .A2(n9047), .ZN(n9046) );
  NAND2_X1 U8463 ( .A1(n9049), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6727) );
  NAND2_X1 U8464 ( .A1(n9046), .A2(n6727), .ZN(n6742) );
  NAND2_X1 U8465 ( .A1(n6743), .A2(n6742), .ZN(n6741) );
  INV_X1 U8466 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6728) );
  OR2_X1 U8467 ( .A1(n6747), .A2(n6728), .ZN(n6729) );
  NAND2_X1 U8468 ( .A1(n6741), .A2(n6729), .ZN(n9060) );
  XNOR2_X1 U8469 ( .A(n9054), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9061) );
  NAND2_X1 U8470 ( .A1(n9060), .A2(n9061), .ZN(n9059) );
  INV_X1 U8471 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6730) );
  OR2_X1 U8472 ( .A1(n9054), .A2(n6730), .ZN(n6731) );
  NAND2_X1 U8473 ( .A1(n9059), .A2(n6731), .ZN(n6733) );
  NAND2_X1 U8474 ( .A1(n6735), .A2(n9614), .ZN(n6732) );
  OAI211_X1 U8475 ( .C1(n6734), .C2(n6733), .A(n9692), .B(n6792), .ZN(n6738)
         );
  AND2_X1 U8476 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6858) );
  AOI21_X1 U8477 ( .B1(n9616), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6858), .ZN(
        n6737) );
  OR2_X1 U8478 ( .A1(n9618), .A2(n6735), .ZN(n9700) );
  NAND2_X1 U8479 ( .A1(n9718), .A2(n6804), .ZN(n6736) );
  NAND4_X1 U8480 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6740)
         );
  OR2_X1 U8481 ( .A1(n6754), .A2(n6740), .ZN(P1_U3247) );
  OAI211_X1 U8482 ( .C1(n6743), .C2(n6742), .A(n9692), .B(n6741), .ZN(n6752)
         );
  OAI211_X1 U8483 ( .C1(n6746), .C2(n6745), .A(n9696), .B(n6744), .ZN(n6751)
         );
  AOI22_X1 U8484 ( .A1(n9616), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6750) );
  INV_X1 U8485 ( .A(n6747), .ZN(n6748) );
  NAND2_X1 U8486 ( .A1(n9718), .A2(n6748), .ZN(n6749) );
  NAND4_X1 U8487 ( .A1(n6752), .A2(n6751), .A3(n6750), .A4(n6749), .ZN(n6753)
         );
  OR2_X1 U8488 ( .A1(n6754), .A2(n6753), .ZN(P1_U3245) );
  INV_X1 U8489 ( .A(n8763), .ZN(n8739) );
  NAND2_X1 U8490 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9055) );
  INV_X1 U8491 ( .A(n9055), .ZN(n6756) );
  INV_X1 U8492 ( .A(n9038), .ZN(n6873) );
  OAI22_X1 U8493 ( .A1(n8760), .A2(n9739), .B1(n6873), .B2(n8759), .ZN(n6755)
         );
  AOI211_X1 U8494 ( .C1(n8757), .C2(n9040), .A(n6756), .B(n6755), .ZN(n6762)
         );
  OAI21_X1 U8495 ( .B1(n6759), .B2(n6758), .A(n6757), .ZN(n6760) );
  NAND2_X1 U8496 ( .A1(n6760), .A2(n8748), .ZN(n6761) );
  OAI211_X1 U8497 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n8739), .A(n6762), .B(
        n6761), .ZN(P1_U3218) );
  INV_X1 U8498 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6776) );
  NOR2_X1 U8499 ( .A1(n9041), .A2(n6693), .ZN(n6763) );
  AOI21_X2 U8500 ( .B1(n8960), .B2(n6764), .A(n6763), .ZN(n7032) );
  NAND2_X1 U8501 ( .A1(n6631), .A2(n7699), .ZN(n6770) );
  NAND2_X1 U8502 ( .A1(n7032), .A2(n6770), .ZN(n6765) );
  NAND2_X1 U8503 ( .A1(n6765), .A2(n8804), .ZN(n6877) );
  NAND2_X1 U8504 ( .A1(n6870), .A2(n6766), .ZN(n6876) );
  INV_X1 U8505 ( .A(n6870), .ZN(n9039) );
  NAND2_X1 U8506 ( .A1(n9039), .A2(n9739), .ZN(n8806) );
  NAND2_X1 U8507 ( .A1(n6876), .A2(n8806), .ZN(n8958) );
  XNOR2_X1 U8508 ( .A(n6877), .B(n8958), .ZN(n6767) );
  AOI222_X1 U8509 ( .A1(n9481), .A2(n6767), .B1(n9038), .B2(n9475), .C1(n9040), 
        .C2(n9474), .ZN(n9744) );
  NAND2_X1 U8510 ( .A1(n7687), .A2(n6693), .ZN(n6768) );
  NAND2_X1 U8511 ( .A1(n6769), .A2(n6768), .ZN(n7037) );
  NAND2_X1 U8512 ( .A1(n7037), .A2(n8956), .ZN(n7036) );
  NAND2_X1 U8513 ( .A1(n6631), .A2(n9749), .ZN(n6771) );
  NAND2_X1 U8514 ( .A1(n7036), .A2(n6771), .ZN(n6772) );
  NAND2_X1 U8515 ( .A1(n6772), .A2(n8958), .ZN(n6872) );
  OAI21_X1 U8516 ( .B1(n6772), .B2(n8958), .A(n6872), .ZN(n9741) );
  OAI211_X1 U8517 ( .C1(n7038), .C2(n9739), .A(n9452), .B(n7049), .ZN(n9734)
         );
  OAI21_X1 U8518 ( .B1(n9739), .B2(n9781), .A(n9734), .ZN(n6773) );
  AOI21_X1 U8519 ( .B1(n9741), .B2(n9786), .A(n6773), .ZN(n6774) );
  NAND2_X1 U8520 ( .A1(n9744), .A2(n6774), .ZN(n6779) );
  NAND2_X1 U8521 ( .A1(n6779), .A2(n9789), .ZN(n6775) );
  OAI21_X1 U8522 ( .B1(n9789), .B2(n6776), .A(n6775), .ZN(P1_U3462) );
  NAND2_X1 U8523 ( .A1(n6778), .A2(n6777), .ZN(n9796) );
  INV_X2 U8524 ( .A(n9796), .ZN(n9799) );
  NAND2_X1 U8525 ( .A1(n6779), .A2(n9799), .ZN(n6780) );
  OAI21_X1 U8526 ( .B1(n9799), .B2(n6719), .A(n6780), .ZN(P1_U3525) );
  OAI22_X1 U8527 ( .A1(n7860), .A2(n5834), .B1(n9855), .B2(n7867), .ZN(n6781)
         );
  AOI21_X1 U8528 ( .B1(n7864), .B2(n5867), .A(n6781), .ZN(n6787) );
  OAI21_X1 U8529 ( .B1(n6784), .B2(n6783), .A(n6782), .ZN(n6785) );
  NAND2_X1 U8530 ( .A1(n6785), .A2(n7856), .ZN(n6786) );
  OAI211_X1 U8531 ( .C1(n6789), .C2(n6788), .A(n6787), .B(n6786), .ZN(P2_U3177) );
  INV_X1 U8532 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7248) );
  AOI22_X1 U8533 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9123), .B1(n6818), .B2(
        n7248), .ZN(n6800) );
  NAND2_X1 U8534 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n9583), .ZN(n6790) );
  OAI21_X1 U8535 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9583), .A(n6790), .ZN(
        n9579) );
  NOR2_X1 U8536 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n9105), .ZN(n6791) );
  AOI21_X1 U8537 ( .B1(n9105), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6791), .ZN(
        n9098) );
  INV_X1 U8538 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6793) );
  MUX2_X1 U8539 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6793), .S(n9075), .Z(n6794)
         );
  INV_X1 U8540 ( .A(n6794), .ZN(n9069) );
  AOI21_X1 U8541 ( .B1(n9075), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9068), .ZN(
        n9084) );
  INV_X1 U8542 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6795) );
  MUX2_X1 U8543 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6795), .S(n9089), .Z(n6796)
         );
  INV_X1 U8544 ( .A(n6796), .ZN(n9083) );
  NOR2_X1 U8545 ( .A1(n9084), .A2(n9083), .ZN(n9082) );
  AOI21_X1 U8546 ( .B1(n9089), .B2(P1_REG2_REG_6__SCAN_IN), .A(n9082), .ZN(
        n9594) );
  XNOR2_X1 U8547 ( .A(n9597), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n9593) );
  NOR2_X1 U8548 ( .A1(n9594), .A2(n9593), .ZN(n9592) );
  NAND2_X1 U8549 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n9609), .ZN(n6797) );
  OAI21_X1 U8550 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9609), .A(n6797), .ZN(
        n9605) );
  OAI21_X1 U8551 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9105), .A(n9096), .ZN(
        n9580) );
  NOR2_X1 U8552 ( .A1(n9579), .A2(n9580), .ZN(n9578) );
  INV_X1 U8553 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6798) );
  AOI22_X1 U8554 ( .A1(n6813), .A2(n6798), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n9630), .ZN(n9622) );
  OAI21_X1 U8555 ( .B1(n6800), .B2(n6799), .A(n9112), .ZN(n6801) );
  INV_X1 U8556 ( .A(n6801), .ZN(n6822) );
  NAND2_X1 U8557 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n9583), .ZN(n6802) );
  OAI21_X1 U8558 ( .B1(n9583), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6802), .ZN(
        n9576) );
  NOR2_X1 U8559 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9105), .ZN(n6803) );
  AOI21_X1 U8560 ( .B1(n9105), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6803), .ZN(
        n9102) );
  NAND2_X1 U8561 ( .A1(n6804), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6805) );
  NAND2_X1 U8562 ( .A1(n6806), .A2(n6805), .ZN(n9077) );
  INV_X1 U8563 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6890) );
  MUX2_X1 U8564 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6890), .S(n9075), .Z(n9078)
         );
  NAND2_X1 U8565 ( .A1(n9077), .A2(n9078), .ZN(n9076) );
  NAND2_X1 U8566 ( .A1(n9075), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6807) );
  NAND2_X1 U8567 ( .A1(n9076), .A2(n6807), .ZN(n9091) );
  INV_X1 U8568 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9792) );
  MUX2_X1 U8569 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n9792), .S(n9089), .Z(n9092)
         );
  NAND2_X1 U8570 ( .A1(n9091), .A2(n9092), .ZN(n9090) );
  NAND2_X1 U8571 ( .A1(n9089), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6808) );
  NAND2_X1 U8572 ( .A1(n9090), .A2(n6808), .ZN(n9587) );
  INV_X1 U8573 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6809) );
  XNOR2_X1 U8574 ( .A(n9597), .B(n6809), .ZN(n9588) );
  AND2_X1 U8575 ( .A1(n9587), .A2(n9588), .ZN(n9589) );
  AND2_X1 U8576 ( .A1(n9597), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6810) );
  OR2_X1 U8577 ( .A1(n9589), .A2(n6810), .ZN(n9600) );
  OR2_X1 U8578 ( .A1(n9609), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6812) );
  NAND2_X1 U8579 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n9609), .ZN(n6811) );
  AND2_X1 U8580 ( .A1(n6812), .A2(n6811), .ZN(n9601) );
  AOI21_X1 U8581 ( .B1(n9609), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9602), .ZN(
        n9101) );
  NAND2_X1 U8582 ( .A1(n9102), .A2(n9101), .ZN(n9100) );
  OAI21_X1 U8583 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9105), .A(n9100), .ZN(
        n9577) );
  NOR2_X1 U8584 ( .A1(n9576), .A2(n9577), .ZN(n9575) );
  AOI21_X1 U8585 ( .B1(n9583), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9575), .ZN(
        n9625) );
  XNOR2_X1 U8586 ( .A(n6813), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n9626) );
  NOR2_X1 U8587 ( .A1(n9625), .A2(n9626), .ZN(n9624) );
  AOI21_X1 U8588 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6813), .A(n9624), .ZN(
        n6816) );
  INV_X1 U8589 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6814) );
  AOI22_X1 U8590 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n9123), .B1(n6818), .B2(
        n6814), .ZN(n6815) );
  NAND2_X1 U8591 ( .A1(n6816), .A2(n6815), .ZN(n9122) );
  OAI21_X1 U8592 ( .B1(n6816), .B2(n6815), .A(n9122), .ZN(n6820) );
  AND2_X1 U8593 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8641) );
  AOI21_X1 U8594 ( .B1(n9616), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n8641), .ZN(
        n6817) );
  OAI21_X1 U8595 ( .B1(n9700), .B2(n6818), .A(n6817), .ZN(n6819) );
  AOI21_X1 U8596 ( .B1(n6820), .B2(n9696), .A(n6819), .ZN(n6821) );
  OAI21_X1 U8597 ( .B1(n6822), .B2(n9711), .A(n6821), .ZN(P1_U3255) );
  INV_X1 U8598 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6825) );
  INV_X1 U8599 ( .A(n6823), .ZN(n6827) );
  OAI222_X1 U8600 ( .A1(n7728), .A2(n6825), .B1(n7730), .B2(n6827), .C1(
        P2_U3151), .C2(n6824), .ZN(P2_U3281) );
  INV_X1 U8601 ( .A(n9124), .ZN(n9658) );
  INV_X1 U8602 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6826) );
  OAI222_X1 U8603 ( .A1(n9658), .A2(P1_U3086), .B1(n7708), .B2(n6827), .C1(
        n6826), .C2(n7522), .ZN(P1_U3341) );
  INV_X1 U8604 ( .A(n6828), .ZN(n6832) );
  NAND4_X1 U8605 ( .A1(n6832), .A2(n6831), .A3(n6830), .A4(n6829), .ZN(n6834)
         );
  INV_X1 U8606 ( .A(n7905), .ZN(n9844) );
  NAND2_X1 U8607 ( .A1(n5842), .A2(n8430), .ZN(n9843) );
  OAI21_X1 U8608 ( .B1(n9844), .B2(n6833), .A(n9843), .ZN(n6835) );
  INV_X2 U8609 ( .A(n8441), .ZN(n8398) );
  NAND2_X1 U8610 ( .A1(n6835), .A2(n8398), .ZN(n6837) );
  INV_X1 U8611 ( .A(n8427), .ZN(n8353) );
  AOI22_X1 U8612 ( .A1(n8441), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n8353), .ZN(n6836) );
  OAI211_X1 U8613 ( .C1(n8429), .C2(n6926), .A(n6837), .B(n6836), .ZN(P2_U3233) );
  AOI211_X1 U8614 ( .C1(n6840), .C2(n6839), .A(n8249), .B(n6838), .ZN(n6841)
         );
  INV_X1 U8615 ( .A(n6841), .ZN(n6855) );
  NAND3_X1 U8616 ( .A1(n6844), .A2(n6843), .A3(n6842), .ZN(n6845) );
  AOI21_X1 U8617 ( .B1(n4427), .B2(n6845), .A(n9825), .ZN(n6853) );
  AND3_X1 U8618 ( .A1(n6848), .A2(n6847), .A3(n6846), .ZN(n6849) );
  OAI21_X1 U8619 ( .B1(n6850), .B2(n6849), .A(n9816), .ZN(n6851) );
  NAND2_X1 U8620 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6965) );
  NAND2_X1 U8621 ( .A1(n6851), .A2(n6965), .ZN(n6852) );
  AOI211_X1 U8622 ( .C1(n9840), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6853), .B(
        n6852), .ZN(n6854) );
  OAI211_X1 U8623 ( .C1(n8246), .C2(n6856), .A(n6855), .B(n6854), .ZN(P2_U3186) );
  INV_X1 U8624 ( .A(n7052), .ZN(n6865) );
  INV_X1 U8625 ( .A(n7046), .ZN(n9037) );
  OAI22_X1 U8626 ( .A1(n9755), .A2(n8760), .B1(n8728), .B2(n6870), .ZN(n6857)
         );
  AOI211_X1 U8627 ( .C1(n8726), .C2(n9037), .A(n6858), .B(n6857), .ZN(n6864)
         );
  AOI21_X1 U8628 ( .B1(n6859), .B2(n6860), .A(n8766), .ZN(n6862) );
  NAND2_X1 U8629 ( .A1(n6862), .A2(n6861), .ZN(n6863) );
  OAI211_X1 U8630 ( .C1(n8739), .C2(n6865), .A(n6864), .B(n6863), .ZN(P1_U3230) );
  INV_X1 U8631 ( .A(n6866), .ZN(n6869) );
  AOI22_X1 U8632 ( .A1(n8198), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n7587), .ZN(n6867) );
  OAI21_X1 U8633 ( .B1(n6869), .B2(n7730), .A(n6867), .ZN(P2_U3280) );
  INV_X1 U8634 ( .A(n9671), .ZN(n9126) );
  OAI222_X1 U8635 ( .A1(P1_U3086), .A2(n9126), .B1(n7708), .B2(n6869), .C1(
        n6868), .C2(n7522), .ZN(P1_U3340) );
  INV_X1 U8636 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U8637 ( .A1(n6870), .A2(n9739), .ZN(n6871) );
  NAND2_X1 U8638 ( .A1(n6872), .A2(n6871), .ZN(n7048) );
  XNOR2_X1 U8639 ( .A(n9038), .B(n9755), .ZN(n8963) );
  NAND2_X1 U8640 ( .A1(n7048), .A2(n8963), .ZN(n7047) );
  NAND2_X1 U8641 ( .A1(n6873), .A2(n9755), .ZN(n6874) );
  NAND2_X1 U8642 ( .A1(n7047), .A2(n6874), .ZN(n6875) );
  NAND2_X1 U8643 ( .A1(n7046), .A2(n6883), .ZN(n8841) );
  NAND2_X1 U8644 ( .A1(n9037), .A2(n9728), .ZN(n8843) );
  NAND2_X1 U8645 ( .A1(n8841), .A2(n8843), .ZN(n8961) );
  NAND2_X1 U8646 ( .A1(n6875), .A2(n8961), .ZN(n7004) );
  OAI21_X1 U8647 ( .B1(n6875), .B2(n8961), .A(n7004), .ZN(n9730) );
  INV_X1 U8648 ( .A(n9730), .ZN(n6885) );
  NAND2_X1 U8649 ( .A1(n6877), .A2(n6876), .ZN(n6878) );
  NAND2_X2 U8650 ( .A1(n6878), .A2(n8806), .ZN(n7044) );
  NAND2_X1 U8651 ( .A1(n7044), .A2(n9755), .ZN(n6879) );
  XNOR2_X1 U8652 ( .A(n7013), .B(n8961), .ZN(n6881) );
  INV_X1 U8653 ( .A(n7088), .ZN(n9036) );
  AOI222_X1 U8654 ( .A1(n9481), .A2(n6881), .B1(n9036), .B2(n9475), .C1(n9038), 
        .C2(n9474), .ZN(n9732) );
  OR2_X1 U8655 ( .A1(n7050), .A2(n6883), .ZN(n7015) );
  AOI21_X1 U8656 ( .B1(n7050), .B2(n6883), .A(n9771), .ZN(n6882) );
  AND2_X1 U8657 ( .A1(n7015), .A2(n6882), .ZN(n9725) );
  AOI21_X1 U8658 ( .B1(n9762), .B2(n6883), .A(n9725), .ZN(n6884) );
  OAI211_X1 U8659 ( .C1(n9766), .C2(n6885), .A(n9732), .B(n6884), .ZN(n6888)
         );
  NAND2_X1 U8660 ( .A1(n6888), .A2(n9789), .ZN(n6886) );
  OAI21_X1 U8661 ( .B1(n9789), .B2(n6887), .A(n6886), .ZN(P1_U3468) );
  NAND2_X1 U8662 ( .A1(n6888), .A2(n9799), .ZN(n6889) );
  OAI21_X1 U8663 ( .B1(n9799), .B2(n6890), .A(n6889), .ZN(P1_U3527) );
  INV_X1 U8664 ( .A(n6891), .ZN(n6892) );
  AOI211_X1 U8665 ( .C1(n6894), .C2(n6893), .A(n7879), .B(n6892), .ZN(n6901)
         );
  AOI22_X1 U8666 ( .A1(n6895), .A2(n7871), .B1(n7870), .B2(n8126), .ZN(n6899)
         );
  INV_X1 U8667 ( .A(n6896), .ZN(n6897) );
  AOI21_X1 U8668 ( .B1(n7876), .B2(n6983), .A(n6897), .ZN(n6898) );
  OAI211_X1 U8669 ( .C1(n7160), .C2(n7874), .A(n6899), .B(n6898), .ZN(n6900)
         );
  OR2_X1 U8670 ( .A1(n6901), .A2(n6900), .ZN(P2_U3158) );
  NAND2_X1 U8671 ( .A1(n6904), .A2(n6903), .ZN(n6905) );
  XNOR2_X1 U8672 ( .A(n6902), .B(n6905), .ZN(n6911) );
  NAND2_X1 U8673 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9086) );
  INV_X1 U8674 ( .A(n9086), .ZN(n6906) );
  AOI21_X1 U8675 ( .B1(n8757), .B2(n9037), .A(n6906), .ZN(n6908) );
  INV_X1 U8676 ( .A(n8848), .ZN(n9035) );
  NAND2_X1 U8677 ( .A1(n8726), .A2(n9035), .ZN(n6907) );
  OAI211_X1 U8678 ( .C1(n8760), .C2(n7084), .A(n6908), .B(n6907), .ZN(n6909)
         );
  AOI21_X1 U8679 ( .B1(n7018), .B2(n8763), .A(n6909), .ZN(n6910) );
  OAI21_X1 U8680 ( .B1(n6911), .B2(n8766), .A(n6910), .ZN(P1_U3239) );
  XNOR2_X1 U8681 ( .A(n6914), .B(n6913), .ZN(n6915) );
  XNOR2_X1 U8682 ( .A(n6912), .B(n6915), .ZN(n6916) );
  NAND2_X1 U8683 ( .A1(n6916), .A2(n8748), .ZN(n6920) );
  NAND2_X1 U8684 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9072) );
  INV_X1 U8685 ( .A(n9072), .ZN(n6918) );
  OAI22_X1 U8686 ( .A1(n8760), .A2(n9728), .B1(n7088), .B2(n8759), .ZN(n6917)
         );
  AOI211_X1 U8687 ( .C1(n8757), .C2(n9038), .A(n6918), .B(n6917), .ZN(n6919)
         );
  OAI211_X1 U8688 ( .C1(n8739), .C2(n6921), .A(n6920), .B(n6919), .ZN(P1_U3227) );
  INV_X1 U8689 ( .A(n6922), .ZN(n6923) );
  AOI21_X1 U8690 ( .B1(n7935), .B2(n6181), .A(n6923), .ZN(n9851) );
  INV_X1 U8691 ( .A(n6924), .ZN(n6925) );
  AOI22_X1 U8692 ( .A1(n6925), .A2(n8436), .B1(n8430), .B2(n8126), .ZN(n6929)
         );
  NOR3_X1 U8693 ( .A1(n6181), .A2(n9845), .A3(n6926), .ZN(n6927) );
  OAI21_X1 U8694 ( .B1(n6927), .B2(n8433), .A(n8127), .ZN(n6928) );
  OAI211_X1 U8695 ( .C1(n9851), .C2(n8440), .A(n6929), .B(n6928), .ZN(n9853)
         );
  AOI21_X1 U8696 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n8353), .A(n9853), .ZN(
        n6934) );
  OR2_X1 U8697 ( .A1(n7231), .A2(n6930), .ZN(n6975) );
  NOR2_X1 U8698 ( .A1(n8441), .A2(n6975), .ZN(n8444) );
  INV_X1 U8699 ( .A(n9851), .ZN(n6932) );
  OAI22_X1 U8700 ( .A1(n8398), .A2(n9990), .B1(n9850), .B2(n8429), .ZN(n6931)
         );
  AOI21_X1 U8701 ( .B1(n8444), .B2(n6932), .A(n6931), .ZN(n6933) );
  OAI21_X1 U8702 ( .B1(n6934), .B2(n8418), .A(n6933), .ZN(P2_U3232) );
  INV_X1 U8703 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6937) );
  INV_X1 U8704 ( .A(n6935), .ZN(n6939) );
  OAI222_X1 U8705 ( .A1(n7728), .A2(n6937), .B1(n7730), .B2(n6939), .C1(
        P2_U3151), .C2(n6936), .ZN(P2_U3279) );
  INV_X1 U8706 ( .A(n9128), .ZN(n9678) );
  INV_X1 U8707 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6938) );
  OAI222_X1 U8708 ( .A1(n9678), .A2(P1_U3086), .B1(n7708), .B2(n6939), .C1(
        n6938), .C2(n7522), .ZN(P1_U3339) );
  OAI21_X1 U8709 ( .B1(n6940), .B2(n6943), .A(n6972), .ZN(n6947) );
  INV_X1 U8710 ( .A(n6947), .ZN(n9856) );
  INV_X1 U8711 ( .A(n8444), .ZN(n7434) );
  INV_X1 U8712 ( .A(n8440), .ZN(n7469) );
  OAI22_X1 U8713 ( .A1(n5834), .A2(n8390), .B1(n5865), .B2(n8392), .ZN(n6946)
         );
  NAND3_X1 U8714 ( .A1(n6924), .A2(n6943), .A3(n6942), .ZN(n6944) );
  AOI21_X1 U8715 ( .B1(n6941), .B2(n6944), .A(n9845), .ZN(n6945) );
  AOI211_X1 U8716 ( .C1(n7469), .C2(n6947), .A(n6946), .B(n6945), .ZN(n6948)
         );
  INV_X1 U8717 ( .A(n6948), .ZN(n9858) );
  OAI22_X1 U8718 ( .A1(n9855), .A2(n8413), .B1(n6788), .B2(n8427), .ZN(n6949)
         );
  NOR2_X1 U8719 ( .A1(n9858), .A2(n6949), .ZN(n6950) );
  MUX2_X1 U8720 ( .A(n6307), .B(n6950), .S(n8398), .Z(n6951) );
  OAI21_X1 U8721 ( .B1(n9856), .B2(n7434), .A(n6951), .ZN(P2_U3231) );
  XOR2_X1 U8722 ( .A(n6954), .B(n6953), .Z(n6955) );
  XNOR2_X1 U8723 ( .A(n6952), .B(n6955), .ZN(n6961) );
  NAND2_X1 U8724 ( .A1(n8763), .A2(n7098), .ZN(n6958) );
  NAND2_X1 U8725 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9598) );
  INV_X1 U8726 ( .A(n9598), .ZN(n6956) );
  AOI21_X1 U8727 ( .B1(n8757), .B2(n9036), .A(n6956), .ZN(n6957) );
  OAI211_X1 U8728 ( .C1(n8854), .C2(n8759), .A(n6958), .B(n6957), .ZN(n6959)
         );
  AOI21_X1 U8729 ( .B1(n8849), .B2(n8741), .A(n6959), .ZN(n6960) );
  OAI21_X1 U8730 ( .B1(n6961), .B2(n8766), .A(n6960), .ZN(P1_U3213) );
  INV_X1 U8731 ( .A(n7073), .ZN(n6962) );
  AOI21_X1 U8732 ( .B1(n6964), .B2(n6963), .A(n6962), .ZN(n6971) );
  INV_X1 U8733 ( .A(n6965), .ZN(n6967) );
  NOR2_X1 U8734 ( .A1(n7867), .A2(n9867), .ZN(n6966) );
  AOI211_X1 U8735 ( .C1(n7864), .C2(n8124), .A(n6967), .B(n6966), .ZN(n6970)
         );
  INV_X1 U8736 ( .A(n6968), .ZN(n7112) );
  AOI22_X1 U8737 ( .A1(n7112), .A2(n7871), .B1(n7870), .B2(n5867), .ZN(n6969)
         );
  OAI211_X1 U8738 ( .C1(n6971), .C2(n7879), .A(n6970), .B(n6969), .ZN(P2_U3170) );
  NAND3_X1 U8739 ( .A1(n6972), .A2(n6184), .A3(n7906), .ZN(n6973) );
  AND2_X1 U8740 ( .A1(n6974), .A2(n6973), .ZN(n9861) );
  AND2_X1 U8741 ( .A1(n8440), .A2(n6975), .ZN(n6976) );
  NAND3_X1 U8742 ( .A1(n6941), .A2(n6979), .A3(n6978), .ZN(n6980) );
  NAND2_X1 U8743 ( .A1(n6977), .A2(n6980), .ZN(n6981) );
  AOI222_X1 U8744 ( .A1(n8436), .A2(n6981), .B1(n8126), .B2(n8433), .C1(n8125), 
        .C2(n8430), .ZN(n9859) );
  MUX2_X1 U8745 ( .A(n6982), .B(n9859), .S(n8398), .Z(n6985) );
  AOI22_X1 U8746 ( .A1(n8382), .A2(n6983), .B1(n6895), .B2(n8353), .ZN(n6984)
         );
  OAI211_X1 U8747 ( .C1(n9861), .C2(n8386), .A(n6985), .B(n6984), .ZN(P2_U3230) );
  OAI21_X1 U8748 ( .B1(n6988), .B2(n6987), .A(n6986), .ZN(n7001) );
  NAND2_X1 U8749 ( .A1(n9840), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n6989) );
  NAND2_X1 U8750 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7224) );
  OAI211_X1 U8751 ( .C1(n8246), .C2(n6990), .A(n6989), .B(n7224), .ZN(n7000)
         );
  AOI21_X1 U8752 ( .B1(n6993), .B2(n6992), .A(n6991), .ZN(n6998) );
  AOI21_X1 U8753 ( .B1(n6996), .B2(n6995), .A(n6994), .ZN(n6997) );
  OAI22_X1 U8754 ( .A1(n6998), .A2(n9832), .B1(n6997), .B2(n9825), .ZN(n6999)
         );
  AOI211_X1 U8755 ( .C1(n7001), .C2(n9838), .A(n7000), .B(n6999), .ZN(n7002)
         );
  INV_X1 U8756 ( .A(n7002), .ZN(P2_U3188) );
  NAND2_X1 U8757 ( .A1(n7046), .A2(n9728), .ZN(n7003) );
  NAND2_X1 U8758 ( .A1(n7004), .A2(n7003), .ZN(n7005) );
  NAND2_X1 U8759 ( .A1(n7088), .A2(n9761), .ZN(n8845) );
  NAND2_X1 U8760 ( .A1(n9036), .A2(n7084), .ZN(n8842) );
  NAND2_X1 U8761 ( .A1(n8845), .A2(n8842), .ZN(n8962) );
  NAND2_X1 U8762 ( .A1(n7005), .A2(n8962), .ZN(n7086) );
  OAI21_X1 U8763 ( .B1(n7005), .B2(n8962), .A(n7086), .ZN(n7006) );
  INV_X1 U8764 ( .A(n7006), .ZN(n9765) );
  AND2_X1 U8765 ( .A1(n9009), .A2(P1_D_REG_1__SCAN_IN), .ZN(n7011) );
  AND3_X1 U8766 ( .A1(n7008), .A2(n9563), .A3(n7007), .ZN(n7009) );
  OAI211_X1 U8767 ( .C1(n9746), .C2(n7011), .A(n7010), .B(n7009), .ZN(n7016)
         );
  AND2_X1 U8768 ( .A1(n7083), .A2(n7094), .ZN(n7012) );
  XOR2_X1 U8769 ( .A(n7089), .B(n8962), .Z(n7014) );
  AOI222_X1 U8770 ( .A1(n9481), .A2(n7014), .B1(n9035), .B2(n9475), .C1(n9037), 
        .C2(n9474), .ZN(n9764) );
  MUX2_X1 U8771 ( .A(n6795), .B(n9764), .S(n9366), .Z(n7022) );
  AOI211_X1 U8772 ( .C1(n9761), .C2(n7015), .A(n9771), .B(n7095), .ZN(n9760)
         );
  INV_X1 U8773 ( .A(n7018), .ZN(n7019) );
  OAI22_X1 U8774 ( .A1(n9738), .A2(n7084), .B1(n7019), .B2(n9733), .ZN(n7020)
         );
  AOI21_X1 U8775 ( .B1(n9760), .B2(n9724), .A(n7020), .ZN(n7021) );
  OAI211_X1 U8776 ( .C1(n9765), .C2(n9369), .A(n7022), .B(n7021), .ZN(P1_U3287) );
  NAND2_X1 U8777 ( .A1(n8248), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7023) );
  OAI21_X1 U8778 ( .B1(n7779), .B2(n8248), .A(n7023), .ZN(P2_U3520) );
  INV_X1 U8779 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7026) );
  NAND2_X1 U8780 ( .A1(n5880), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7025) );
  INV_X1 U8781 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8262) );
  OR2_X1 U8782 ( .A1(n6060), .A2(n8262), .ZN(n7024) );
  OAI211_X1 U8783 ( .C1(n7027), .C2(n7026), .A(n7025), .B(n7024), .ZN(n7028)
         );
  INV_X1 U8784 ( .A(n7028), .ZN(n7029) );
  NAND2_X1 U8785 ( .A1(n8248), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7031) );
  OAI21_X1 U8786 ( .B1(n8093), .B2(n8248), .A(n7031), .ZN(P2_U3522) );
  XNOR2_X1 U8787 ( .A(n7032), .B(n8956), .ZN(n7033) );
  NAND2_X1 U8788 ( .A1(n7033), .A2(n9481), .ZN(n7035) );
  AOI22_X1 U8789 ( .A1(n9039), .A2(n9475), .B1(n9474), .B2(n9041), .ZN(n7034)
         );
  NAND2_X1 U8790 ( .A1(n7035), .A2(n7034), .ZN(n9751) );
  AOI21_X1 U8791 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n9722), .A(n9751), .ZN(
        n7043) );
  OAI21_X1 U8792 ( .B1(n7037), .B2(n8956), .A(n7036), .ZN(n9752) );
  AOI211_X1 U8793 ( .C1(n7699), .C2(n7039), .A(n9771), .B(n7038), .ZN(n9747)
         );
  AOI22_X1 U8794 ( .A1(n9747), .A2(n9724), .B1(P1_REG2_REG_2__SCAN_IN), .B2(
        n4322), .ZN(n7040) );
  OAI21_X1 U8795 ( .B1(n9749), .B2(n9738), .A(n7040), .ZN(n7041) );
  AOI21_X1 U8796 ( .B1(n9742), .B2(n9752), .A(n7041), .ZN(n7042) );
  OAI21_X1 U8797 ( .B1(n4322), .B2(n7043), .A(n7042), .ZN(P1_U3291) );
  XOR2_X1 U8798 ( .A(n8963), .B(n7044), .Z(n7045) );
  OAI222_X1 U8799 ( .A1(n9530), .A2(n7046), .B1(n9532), .B2(n6870), .C1(n7045), 
        .C2(n9523), .ZN(n9756) );
  INV_X1 U8800 ( .A(n9756), .ZN(n7057) );
  OAI21_X1 U8801 ( .B1(n7048), .B2(n8963), .A(n7047), .ZN(n9758) );
  OAI211_X1 U8802 ( .C1(n4571), .C2(n9755), .A(n9452), .B(n7050), .ZN(n9754)
         );
  NAND2_X1 U8803 ( .A1(n9349), .A2(n7051), .ZN(n7054) );
  AOI22_X1 U8804 ( .A1(n4322), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7052), .B2(
        n9722), .ZN(n7053) );
  OAI211_X1 U8805 ( .C1(n9735), .C2(n9754), .A(n7054), .B(n7053), .ZN(n7055)
         );
  AOI21_X1 U8806 ( .B1(n9758), .B2(n9742), .A(n7055), .ZN(n7056) );
  OAI21_X1 U8807 ( .B1(n7057), .B2(n4322), .A(n7056), .ZN(P1_U3289) );
  INV_X1 U8808 ( .A(n7058), .ZN(n7105) );
  AOI22_X1 U8809 ( .A1(n9688), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7106), .ZN(n7059) );
  OAI21_X1 U8810 ( .B1(n7105), .B2(n7708), .A(n7059), .ZN(P1_U3338) );
  INV_X1 U8811 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7060) );
  OAI22_X1 U8812 ( .A1(n9735), .A2(n7061), .B1(n7060), .B2(n9733), .ZN(n7064)
         );
  OR2_X1 U8813 ( .A1(n4322), .A2(n9532), .ZN(n9347) );
  INV_X1 U8814 ( .A(n9042), .ZN(n7062) );
  NOR2_X1 U8815 ( .A1(n9347), .A2(n7062), .ZN(n7063) );
  AOI211_X1 U8816 ( .C1(n4322), .C2(P1_REG2_REG_1__SCAN_IN), .A(n7064), .B(
        n7063), .ZN(n7068) );
  OR2_X1 U8817 ( .A1(n4322), .A2(n9530), .ZN(n9377) );
  OAI22_X1 U8818 ( .A1(n6693), .A2(n9738), .B1(n9377), .B2(n6631), .ZN(n7065)
         );
  AOI21_X1 U8819 ( .B1(n9742), .B2(n7066), .A(n7065), .ZN(n7067) );
  OAI211_X1 U8820 ( .C1(n4322), .C2(n7069), .A(n7068), .B(n7067), .ZN(P1_U3292) );
  INV_X1 U8821 ( .A(n7070), .ZN(n7072) );
  NAND3_X1 U8822 ( .A1(n7073), .A2(n7072), .A3(n7071), .ZN(n7074) );
  AOI21_X1 U8823 ( .B1(n7075), .B2(n7074), .A(n7879), .ZN(n7082) );
  INV_X1 U8824 ( .A(n7076), .ZN(n7077) );
  AOI21_X1 U8825 ( .B1(n7876), .B2(n7078), .A(n7077), .ZN(n7079) );
  OAI21_X1 U8826 ( .B1(n7874), .B2(n7671), .A(n7079), .ZN(n7081) );
  OAI22_X1 U8827 ( .A1(n7162), .A2(n7861), .B1(n7860), .B2(n7160), .ZN(n7080)
         );
  OR3_X1 U8828 ( .A1(n7082), .A2(n7081), .A3(n7080), .ZN(P2_U3167) );
  INV_X1 U8829 ( .A(n7083), .ZN(n7125) );
  NAND2_X1 U8830 ( .A1(n7088), .A2(n7084), .ZN(n7085) );
  NAND2_X1 U8831 ( .A1(n7086), .A2(n7085), .ZN(n7087) );
  OR2_X1 U8832 ( .A1(n8848), .A2(n8849), .ZN(n8965) );
  NAND2_X1 U8833 ( .A1(n8849), .A2(n8848), .ZN(n8838) );
  NAND2_X1 U8834 ( .A1(n8965), .A2(n8838), .ZN(n7090) );
  NAND2_X1 U8835 ( .A1(n7087), .A2(n7090), .ZN(n7121) );
  OAI21_X1 U8836 ( .B1(n7087), .B2(n7090), .A(n7121), .ZN(n7185) );
  OAI22_X1 U8837 ( .A1(n7088), .A2(n9532), .B1(n8854), .B2(n9530), .ZN(n7093)
         );
  NAND2_X1 U8838 ( .A1(n7139), .A2(n8842), .ZN(n8840) );
  OR2_X1 U8839 ( .A1(n8840), .A2(n7090), .ZN(n7115) );
  NAND2_X1 U8840 ( .A1(n8840), .A2(n7090), .ZN(n7091) );
  AOI21_X1 U8841 ( .B1(n7115), .B2(n7091), .A(n9523), .ZN(n7092) );
  AOI211_X1 U8842 ( .C1(n7125), .C2(n7185), .A(n7093), .B(n7092), .ZN(n7188)
         );
  INV_X1 U8843 ( .A(n7095), .ZN(n7097) );
  NAND2_X1 U8844 ( .A1(n7095), .A2(n8857), .ZN(n7129) );
  INV_X1 U8845 ( .A(n7129), .ZN(n7096) );
  AOI21_X1 U8846 ( .B1(n8849), .B2(n7097), .A(n7096), .ZN(n7186) );
  NOR2_X1 U8847 ( .A1(n9735), .A2(n9771), .ZN(n9303) );
  NAND2_X1 U8848 ( .A1(n7186), .A2(n9303), .ZN(n7100) );
  AOI22_X1 U8849 ( .A1(n4322), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7098), .B2(
        n9722), .ZN(n7099) );
  OAI211_X1 U8850 ( .C1(n8857), .C2(n9738), .A(n7100), .B(n7099), .ZN(n7101)
         );
  AOI21_X1 U8851 ( .B1(n7185), .B2(n4419), .A(n7101), .ZN(n7102) );
  OAI21_X1 U8852 ( .B1(n7188), .B2(n4322), .A(n7102), .ZN(P1_U3286) );
  OAI222_X1 U8853 ( .A1(n7730), .A2(n7105), .B1(n7104), .B2(P2_U3151), .C1(
        n7103), .C2(n8577), .ZN(P2_U3278) );
  AOI22_X1 U8854 ( .A1(n9717), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7106), .ZN(n7107) );
  OAI21_X1 U8855 ( .B1(n7167), .B2(n7708), .A(n7107), .ZN(P1_U3337) );
  NAND2_X1 U8856 ( .A1(n7952), .A2(n7960), .ZN(n7948) );
  XNOR2_X1 U8857 ( .A(n7108), .B(n7948), .ZN(n9865) );
  XNOR2_X1 U8858 ( .A(n7109), .B(n7948), .ZN(n7110) );
  AOI222_X1 U8859 ( .A1(n8436), .A2(n7110), .B1(n5867), .B2(n8433), .C1(n8124), 
        .C2(n8430), .ZN(n9866) );
  MUX2_X1 U8860 ( .A(n7111), .B(n9866), .S(n8398), .Z(n7114) );
  AOI22_X1 U8861 ( .A1(n8382), .A2(n4635), .B1(n8353), .B2(n7112), .ZN(n7113)
         );
  OAI211_X1 U8862 ( .C1(n8386), .C2(n9865), .A(n7114), .B(n7113), .ZN(P2_U3229) );
  OR2_X1 U8863 ( .A1(n8858), .A2(n8854), .ZN(n8847) );
  NAND2_X1 U8864 ( .A1(n8858), .A2(n8854), .ZN(n8839) );
  NAND2_X1 U8865 ( .A1(n8847), .A2(n8839), .ZN(n7122) );
  INV_X1 U8866 ( .A(n7122), .ZN(n7117) );
  NAND2_X1 U8867 ( .A1(n7115), .A2(n8838), .ZN(n7116) );
  NAND2_X1 U8868 ( .A1(n7116), .A2(n7117), .ZN(n7169) );
  OAI21_X1 U8869 ( .B1(n7117), .B2(n7116), .A(n7169), .ZN(n7118) );
  NAND2_X1 U8870 ( .A1(n7118), .A2(n9481), .ZN(n7128) );
  OAI22_X1 U8871 ( .A1(n8848), .A2(n9532), .B1(n7265), .B2(n9530), .ZN(n7119)
         );
  INV_X1 U8872 ( .A(n7119), .ZN(n7127) );
  NAND2_X1 U8873 ( .A1(n8857), .A2(n8848), .ZN(n7120) );
  NAND2_X1 U8874 ( .A1(n7121), .A2(n7120), .ZN(n7123) );
  NAND2_X1 U8875 ( .A1(n7123), .A2(n7122), .ZN(n7146) );
  OR2_X1 U8876 ( .A1(n7123), .A2(n7122), .ZN(n7124) );
  NAND2_X1 U8877 ( .A1(n7146), .A2(n7124), .ZN(n9775) );
  NAND2_X1 U8878 ( .A1(n9775), .A2(n7125), .ZN(n7126) );
  NAND2_X1 U8879 ( .A1(n7129), .A2(n8858), .ZN(n7130) );
  NAND2_X1 U8880 ( .A1(n7178), .A2(n7130), .ZN(n9772) );
  INV_X1 U8881 ( .A(n9303), .ZN(n7133) );
  AOI22_X1 U8882 ( .A1(n4322), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7261), .B2(
        n9722), .ZN(n7132) );
  NAND2_X1 U8883 ( .A1(n9349), .A2(n8858), .ZN(n7131) );
  OAI211_X1 U8884 ( .C1(n9772), .C2(n7133), .A(n7132), .B(n7131), .ZN(n7134)
         );
  AOI21_X1 U8885 ( .B1(n9775), .B2(n4419), .A(n7134), .ZN(n7135) );
  OAI21_X1 U8886 ( .B1(n9777), .B2(n4322), .A(n7135), .ZN(P1_U3285) );
  NAND2_X1 U8887 ( .A1(n8870), .A2(n8847), .ZN(n8954) );
  AND2_X1 U8888 ( .A1(n8839), .A2(n8838), .ZN(n7136) );
  NAND2_X1 U8889 ( .A1(n9779), .A2(n7265), .ZN(n8865) );
  NAND2_X1 U8890 ( .A1(n8965), .A2(n8842), .ZN(n7137) );
  NOR2_X1 U8891 ( .A1(n8954), .A2(n7137), .ZN(n7138) );
  OR2_X1 U8892 ( .A1(n7208), .A2(n9533), .ZN(n8874) );
  NAND2_X1 U8893 ( .A1(n7208), .A2(n9533), .ZN(n8872) );
  NAND2_X1 U8894 ( .A1(n8874), .A2(n8872), .ZN(n8969) );
  INV_X1 U8895 ( .A(n8969), .ZN(n7142) );
  INV_X1 U8896 ( .A(n7205), .ZN(n7144) );
  AOI21_X1 U8897 ( .B1(n8810), .B2(n8808), .A(n7142), .ZN(n7143) );
  NOR2_X1 U8898 ( .A1(n7144), .A2(n7143), .ZN(n7199) );
  OR2_X1 U8899 ( .A1(n4322), .A2(n9523), .ZN(n9386) );
  NAND2_X1 U8900 ( .A1(n7146), .A2(n7145), .ZN(n7177) );
  NAND2_X1 U8901 ( .A1(n8870), .A2(n8865), .ZN(n7176) );
  NAND2_X1 U8902 ( .A1(n7177), .A2(n7176), .ZN(n7175) );
  INV_X1 U8903 ( .A(n7265), .ZN(n9033) );
  NAND2_X1 U8904 ( .A1(n7175), .A2(n7147), .ZN(n7148) );
  NAND2_X1 U8905 ( .A1(n7148), .A2(n8969), .ZN(n7210) );
  OAI21_X1 U8906 ( .B1(n7148), .B2(n8969), .A(n7210), .ZN(n7194) );
  NAND2_X1 U8907 ( .A1(n7194), .A2(n9742), .ZN(n7156) );
  NOR2_X2 U8908 ( .A1(n7178), .A2(n9779), .ZN(n7149) );
  INV_X1 U8909 ( .A(n7149), .ZN(n7150) );
  INV_X1 U8910 ( .A(n7208), .ZN(n8606) );
  AOI211_X1 U8911 ( .C1(n7208), .C2(n7150), .A(n9771), .B(n7214), .ZN(n7195)
         );
  INV_X1 U8912 ( .A(n9347), .ZN(n9380) );
  AOI22_X1 U8913 ( .A1(n4322), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n4919), .B2(
        n9722), .ZN(n7151) );
  OAI21_X1 U8914 ( .B1(n9377), .B2(n8643), .A(n7151), .ZN(n7152) );
  AOI21_X1 U8915 ( .B1(n9380), .B2(n9033), .A(n7152), .ZN(n7153) );
  OAI21_X1 U8916 ( .B1(n8606), .B2(n9738), .A(n7153), .ZN(n7154) );
  AOI21_X1 U8917 ( .B1(n7195), .B2(n9724), .A(n7154), .ZN(n7155) );
  OAI211_X1 U8918 ( .C1(n7199), .C2(n9386), .A(n7156), .B(n7155), .ZN(P1_U3283) );
  XNOR2_X1 U8919 ( .A(n7157), .B(n7911), .ZN(n9873) );
  XNOR2_X1 U8920 ( .A(n7158), .B(n7911), .ZN(n7159) );
  OAI222_X1 U8921 ( .A1(n8390), .A2(n7160), .B1(n8392), .B2(n7671), .C1(n7159), 
        .C2(n9845), .ZN(n9871) );
  AOI21_X1 U8922 ( .B1(n7469), .B2(n9873), .A(n9871), .ZN(n7166) );
  NOR2_X1 U8923 ( .A1(n8398), .A2(n7161), .ZN(n7164) );
  OAI22_X1 U8924 ( .A1(n8429), .A2(n9870), .B1(n7162), .B2(n8427), .ZN(n7163)
         );
  AOI211_X1 U8925 ( .C1(n9873), .C2(n8444), .A(n7164), .B(n7163), .ZN(n7165)
         );
  OAI21_X1 U8926 ( .B1(n7166), .B2(n8418), .A(n7165), .ZN(P2_U3228) );
  INV_X1 U8927 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7168) );
  OAI222_X1 U8928 ( .A1(n7728), .A2(n7168), .B1(n8251), .B2(P2_U3151), .C1(
        n7730), .C2(n7167), .ZN(P2_U3277) );
  NAND2_X1 U8929 ( .A1(n7169), .A2(n8839), .ZN(n7171) );
  INV_X1 U8930 ( .A(n7176), .ZN(n7170) );
  XNOR2_X1 U8931 ( .A(n7171), .B(n7170), .ZN(n7172) );
  NAND2_X1 U8932 ( .A1(n7172), .A2(n9481), .ZN(n7174) );
  OR2_X1 U8933 ( .A1(n8854), .A2(n9532), .ZN(n7173) );
  NAND2_X1 U8934 ( .A1(n7174), .A2(n7173), .ZN(n9783) );
  INV_X1 U8935 ( .A(n9783), .ZN(n7184) );
  OAI21_X1 U8936 ( .B1(n7177), .B2(n7176), .A(n7175), .ZN(n9785) );
  XOR2_X1 U8937 ( .A(n9779), .B(n7178), .Z(n7179) );
  INV_X1 U8938 ( .A(n9533), .ZN(n9032) );
  AOI22_X1 U8939 ( .A1(n7179), .A2(n9452), .B1(n9475), .B2(n9032), .ZN(n9780)
         );
  AOI22_X1 U8940 ( .A1(n4322), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7334), .B2(
        n9722), .ZN(n7181) );
  NAND2_X1 U8941 ( .A1(n9349), .A2(n9779), .ZN(n7180) );
  OAI211_X1 U8942 ( .C1(n9780), .C2(n9735), .A(n7181), .B(n7180), .ZN(n7182)
         );
  AOI21_X1 U8943 ( .B1(n9785), .B2(n9742), .A(n7182), .ZN(n7183) );
  OAI21_X1 U8944 ( .B1(n7184), .B2(n4322), .A(n7183), .ZN(P1_U3284) );
  INV_X1 U8945 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7191) );
  INV_X1 U8946 ( .A(n7185), .ZN(n7189) );
  AOI22_X1 U8947 ( .A1(n7186), .A2(n9452), .B1(n9762), .B2(n8849), .ZN(n7187)
         );
  OAI211_X1 U8948 ( .C1(n7189), .C2(n9769), .A(n7188), .B(n7187), .ZN(n7192)
         );
  NAND2_X1 U8949 ( .A1(n7192), .A2(n9789), .ZN(n7190) );
  OAI21_X1 U8950 ( .B1(n9789), .B2(n7191), .A(n7190), .ZN(P1_U3474) );
  NAND2_X1 U8951 ( .A1(n7192), .A2(n9799), .ZN(n7193) );
  OAI21_X1 U8952 ( .B1(n9799), .B2(n6809), .A(n7193), .ZN(P1_U3529) );
  INV_X1 U8953 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7201) );
  NAND2_X1 U8954 ( .A1(n7194), .A2(n9786), .ZN(n7198) );
  OAI22_X1 U8955 ( .A1(n7265), .A2(n9532), .B1(n8643), .B2(n9530), .ZN(n7196)
         );
  AOI211_X1 U8956 ( .C1(n9762), .C2(n7208), .A(n7196), .B(n7195), .ZN(n7197)
         );
  OAI211_X1 U8957 ( .C1(n9523), .C2(n7199), .A(n7198), .B(n7197), .ZN(n7202)
         );
  NAND2_X1 U8958 ( .A1(n7202), .A2(n9789), .ZN(n7200) );
  OAI21_X1 U8959 ( .B1(n9789), .B2(n7201), .A(n7200), .ZN(P1_U3483) );
  INV_X1 U8960 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7204) );
  NAND2_X1 U8961 ( .A1(n7202), .A2(n9799), .ZN(n7203) );
  OAI21_X1 U8962 ( .B1(n9799), .B2(n7204), .A(n7203), .ZN(P1_U3532) );
  NAND2_X1 U8963 ( .A1(n9535), .A2(n8643), .ZN(n8878) );
  NAND2_X1 U8964 ( .A1(n8875), .A2(n8878), .ZN(n8970) );
  INV_X1 U8965 ( .A(n8970), .ZN(n7206) );
  OAI211_X1 U8966 ( .C1(n7207), .C2(n7206), .A(n9481), .B(n7251), .ZN(n9537)
         );
  OAI21_X1 U8967 ( .B1(n7211), .B2(n8970), .A(n7242), .ZN(n9529) );
  NAND2_X1 U8968 ( .A1(n9529), .A2(n9742), .ZN(n7218) );
  NAND2_X1 U8969 ( .A1(n9380), .A2(n9032), .ZN(n7213) );
  AOI22_X1 U8970 ( .A1(n4322), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n8730), .B2(
        n9722), .ZN(n7212) );
  OAI211_X1 U8971 ( .C1(n9531), .C2(n9377), .A(n7213), .B(n7212), .ZN(n7216)
         );
  INV_X1 U8972 ( .A(n9535), .ZN(n8733) );
  OAI211_X1 U8973 ( .C1(n7214), .C2(n8733), .A(n9452), .B(n7246), .ZN(n9536)
         );
  NOR2_X1 U8974 ( .A1(n9536), .A2(n9735), .ZN(n7215) );
  AOI211_X1 U8975 ( .C1(n9349), .C2(n9535), .A(n7216), .B(n7215), .ZN(n7217)
         );
  OAI211_X1 U8976 ( .C1(n4322), .C2(n9537), .A(n7218), .B(n7217), .ZN(P1_U3282) );
  INV_X1 U8977 ( .A(n7219), .ZN(n7220) );
  AOI211_X1 U8978 ( .C1(n7222), .C2(n7221), .A(n7879), .B(n7220), .ZN(n7229)
         );
  OAI22_X1 U8979 ( .A1(n7860), .A2(n7223), .B1(n9876), .B2(n7867), .ZN(n7228)
         );
  INV_X1 U8980 ( .A(n7224), .ZN(n7225) );
  AOI21_X1 U8981 ( .B1(n7864), .B2(n8123), .A(n7225), .ZN(n7226) );
  OAI21_X1 U8982 ( .B1(n7236), .B2(n7861), .A(n7226), .ZN(n7227) );
  OR3_X1 U8983 ( .A1(n7229), .A2(n7228), .A3(n7227), .ZN(P2_U3179) );
  INV_X1 U8984 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7232) );
  INV_X1 U8985 ( .A(n7230), .ZN(n7705) );
  OAI222_X1 U8986 ( .A1(n7728), .A2(n7232), .B1(n7730), .B2(n7705), .C1(n7231), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  NAND2_X1 U8987 ( .A1(n7417), .A2(n7951), .ZN(n7366) );
  XOR2_X1 U8988 ( .A(n7908), .B(n7366), .Z(n9878) );
  XNOR2_X1 U8989 ( .A(n7233), .B(n7908), .ZN(n7234) );
  AOI222_X1 U8990 ( .A1(n8436), .A2(n7234), .B1(n8123), .B2(n8430), .C1(n8124), 
        .C2(n8433), .ZN(n9875) );
  MUX2_X1 U8991 ( .A(n7235), .B(n9875), .S(n8398), .Z(n7240) );
  INV_X1 U8992 ( .A(n7236), .ZN(n7237) );
  AOI22_X1 U8993 ( .A1(n8382), .A2(n7238), .B1(n8353), .B2(n7237), .ZN(n7239)
         );
  OAI211_X1 U8994 ( .C1(n8386), .C2(n9878), .A(n7240), .B(n7239), .ZN(P2_U3227) );
  INV_X1 U8995 ( .A(n8643), .ZN(n9031) );
  NAND2_X1 U8996 ( .A1(n9526), .A2(n9531), .ZN(n8877) );
  NAND2_X1 U8997 ( .A1(n8880), .A2(n8877), .ZN(n8971) );
  OAI21_X1 U8998 ( .B1(n7243), .B2(n8971), .A(n7406), .ZN(n7244) );
  INV_X1 U8999 ( .A(n7244), .ZN(n9528) );
  INV_X1 U9000 ( .A(n7409), .ZN(n7245) );
  AOI211_X1 U9001 ( .C1(n9526), .C2(n7246), .A(n9771), .B(n7245), .ZN(n9525)
         );
  INV_X1 U9002 ( .A(n9526), .ZN(n8648) );
  NOR2_X1 U9003 ( .A1(n8648), .A2(n9738), .ZN(n7250) );
  INV_X1 U9004 ( .A(n8645), .ZN(n7247) );
  OAI22_X1 U9005 ( .A1(n9366), .A2(n7248), .B1(n7247), .B2(n9733), .ZN(n7249)
         );
  AOI211_X1 U9006 ( .C1(n9525), .C2(n9724), .A(n7250), .B(n7249), .ZN(n7257)
         );
  INV_X1 U9007 ( .A(n8971), .ZN(n7253) );
  NAND2_X1 U9008 ( .A1(n7251), .A2(n8875), .ZN(n7252) );
  OAI211_X1 U9009 ( .C1(n7253), .C2(n7252), .A(n7402), .B(n9481), .ZN(n7255)
         );
  OR2_X1 U9010 ( .A1(n8643), .A2(n9532), .ZN(n7254) );
  OAI211_X1 U9011 ( .C1(n9508), .C2(n9530), .A(n7255), .B(n7254), .ZN(n9524)
         );
  NAND2_X1 U9012 ( .A1(n9524), .A2(n9366), .ZN(n7256) );
  OAI211_X1 U9013 ( .C1(n9528), .C2(n9369), .A(n7257), .B(n7256), .ZN(P1_U3281) );
  OAI21_X1 U9014 ( .B1(n7260), .B2(n7259), .A(n7258), .ZN(n7268) );
  INV_X1 U9015 ( .A(n8858), .ZN(n9770) );
  NOR2_X1 U9016 ( .A1(n8760), .A2(n9770), .ZN(n7267) );
  NAND2_X1 U9017 ( .A1(n8763), .A2(n7261), .ZN(n7264) );
  NAND2_X1 U9018 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9610) );
  INV_X1 U9019 ( .A(n9610), .ZN(n7262) );
  AOI21_X1 U9020 ( .B1(n8757), .B2(n9035), .A(n7262), .ZN(n7263) );
  OAI211_X1 U9021 ( .C1(n7265), .C2(n8759), .A(n7264), .B(n7263), .ZN(n7266)
         );
  AOI211_X1 U9022 ( .C1(n7268), .C2(n8748), .A(n7267), .B(n7266), .ZN(n7269)
         );
  INV_X1 U9023 ( .A(n7269), .ZN(P1_U3221) );
  INV_X1 U9024 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9928) );
  NOR2_X1 U9025 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7307) );
  NOR2_X1 U9026 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7305) );
  NOR2_X1 U9027 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7303) );
  NOR2_X1 U9028 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7301) );
  NOR2_X1 U9029 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7299) );
  NOR2_X1 U9030 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7297) );
  INV_X1 U9031 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7271) );
  INV_X1 U9032 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7270) );
  AOI22_X1 U9033 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7271), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n7270), .ZN(n9941) );
  NAND2_X1 U9034 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7295) );
  XOR2_X1 U9035 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(P2_ADDR_REG_11__SCAN_IN), 
        .Z(n9943) );
  NAND2_X1 U9036 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7293) );
  INV_X1 U9037 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9586) );
  XNOR2_X1 U9038 ( .A(n9586), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(n9945) );
  NOR2_X1 U9039 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7277) );
  XNOR2_X1 U9040 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10112) );
  NAND2_X1 U9041 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7275) );
  XNOR2_X1 U9042 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n9993), .ZN(n10110) );
  NAND2_X1 U9043 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7273) );
  XOR2_X1 U9044 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10108) );
  AOI21_X1 U9045 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9921) );
  INV_X1 U9046 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9925) );
  NAND3_X1 U9047 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9923) );
  OAI21_X1 U9048 ( .B1(n9921), .B2(n9925), .A(n9923), .ZN(n10107) );
  NAND2_X1 U9049 ( .A1(n10108), .A2(n10107), .ZN(n7272) );
  NAND2_X1 U9050 ( .A1(n7273), .A2(n7272), .ZN(n10109) );
  NAND2_X1 U9051 ( .A1(n10110), .A2(n10109), .ZN(n7274) );
  NAND2_X1 U9052 ( .A1(n7275), .A2(n7274), .ZN(n10111) );
  NOR2_X1 U9053 ( .A1(n10112), .A2(n10111), .ZN(n7276) );
  NOR2_X1 U9054 ( .A1(n7277), .A2(n7276), .ZN(n7278) );
  NOR2_X1 U9055 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7278), .ZN(n10101) );
  AND2_X1 U9056 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7278), .ZN(n10100) );
  NOR2_X1 U9057 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10100), .ZN(n7279) );
  NOR2_X1 U9058 ( .A1(n10101), .A2(n7279), .ZN(n7280) );
  NAND2_X1 U9059 ( .A1(n7280), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7282) );
  INV_X1 U9060 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9087) );
  XNOR2_X1 U9061 ( .A(n7280), .B(n9087), .ZN(n10099) );
  NAND2_X1 U9062 ( .A1(n10099), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7281) );
  NAND2_X1 U9063 ( .A1(n7282), .A2(n7281), .ZN(n7283) );
  NAND2_X1 U9064 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7283), .ZN(n7285) );
  INV_X1 U9065 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10006) );
  XNOR2_X1 U9066 ( .A(n10006), .B(n7283), .ZN(n10105) );
  NAND2_X1 U9067 ( .A1(n10105), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7284) );
  NAND2_X1 U9068 ( .A1(n7285), .A2(n7284), .ZN(n7286) );
  NAND2_X1 U9069 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7286), .ZN(n7288) );
  INV_X1 U9070 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9612) );
  XNOR2_X1 U9071 ( .A(n9612), .B(n7286), .ZN(n10106) );
  NAND2_X1 U9072 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10106), .ZN(n7287) );
  NAND2_X1 U9073 ( .A1(n7288), .A2(n7287), .ZN(n7289) );
  NAND2_X1 U9074 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7289), .ZN(n7291) );
  XOR2_X1 U9075 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7289), .Z(n10104) );
  NAND2_X1 U9076 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10104), .ZN(n7290) );
  NAND2_X1 U9077 ( .A1(n7291), .A2(n7290), .ZN(n9944) );
  NAND2_X1 U9078 ( .A1(n9945), .A2(n9944), .ZN(n7292) );
  NAND2_X1 U9079 ( .A1(n7293), .A2(n7292), .ZN(n9942) );
  NAND2_X1 U9080 ( .A1(n9943), .A2(n9942), .ZN(n7294) );
  NAND2_X1 U9081 ( .A1(n7295), .A2(n7294), .ZN(n9940) );
  NOR2_X1 U9082 ( .A1(n9941), .A2(n9940), .ZN(n7296) );
  NOR2_X1 U9083 ( .A1(n7297), .A2(n7296), .ZN(n9939) );
  INV_X1 U9084 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9647) );
  INV_X1 U9085 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8153) );
  AOI22_X1 U9086 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n9647), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n8153), .ZN(n9938) );
  NOR2_X1 U9087 ( .A1(n9939), .A2(n9938), .ZN(n7298) );
  NOR2_X1 U9088 ( .A1(n7299), .A2(n7298), .ZN(n9937) );
  INV_X1 U9089 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9662) );
  INV_X1 U9090 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8175) );
  AOI22_X1 U9091 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n9662), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n8175), .ZN(n9936) );
  NOR2_X1 U9092 ( .A1(n9937), .A2(n9936), .ZN(n7300) );
  NOR2_X1 U9093 ( .A1(n7301), .A2(n7300), .ZN(n9935) );
  INV_X1 U9094 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9674) );
  INV_X1 U9095 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8189) );
  AOI22_X1 U9096 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9674), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8189), .ZN(n9934) );
  NOR2_X1 U9097 ( .A1(n9935), .A2(n9934), .ZN(n7302) );
  NOR2_X1 U9098 ( .A1(n7303), .A2(n7302), .ZN(n9933) );
  INV_X1 U9099 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9687) );
  INV_X1 U9100 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8210) );
  AOI22_X1 U9101 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9687), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n8210), .ZN(n9932) );
  NOR2_X1 U9102 ( .A1(n9933), .A2(n9932), .ZN(n7304) );
  NOR2_X1 U9103 ( .A1(n7305), .A2(n7304), .ZN(n9931) );
  INV_X1 U9104 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9704) );
  INV_X1 U9105 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8225) );
  AOI22_X1 U9106 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9704), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n8225), .ZN(n9930) );
  NOR2_X1 U9107 ( .A1(n9931), .A2(n9930), .ZN(n7306) );
  NOR2_X1 U9108 ( .A1(n7307), .A2(n7306), .ZN(n9927) );
  NOR2_X1 U9109 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9927), .ZN(n7308) );
  NAND2_X1 U9110 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9927), .ZN(n9926) );
  OAI21_X1 U9111 ( .B1(n9928), .B2(n7308), .A(n9926), .ZN(n7310) );
  XNOR2_X1 U9112 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7309) );
  XNOR2_X1 U9113 ( .A(n7310), .B(n7309), .ZN(ADD_1068_U4) );
  NOR2_X1 U9114 ( .A1(n7312), .A2(n7311), .ZN(n7314) );
  XNOR2_X1 U9115 ( .A(n7314), .B(n7313), .ZN(n7326) );
  AOI21_X1 U9116 ( .B1(n7316), .B2(n7430), .A(n7315), .ZN(n7317) );
  NOR2_X1 U9117 ( .A1(n7317), .A2(n9832), .ZN(n7325) );
  AOI21_X1 U9118 ( .B1(n5939), .B2(n7319), .A(n7318), .ZN(n7320) );
  OR2_X1 U9119 ( .A1(n7320), .A2(n9825), .ZN(n7322) );
  AND2_X1 U9120 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7552) );
  AOI21_X1 U9121 ( .B1(n9840), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7552), .ZN(
        n7321) );
  OAI211_X1 U9122 ( .C1(n8246), .C2(n7323), .A(n7322), .B(n7321), .ZN(n7324)
         );
  AOI211_X1 U9123 ( .C1(n7326), .C2(n9838), .A(n7325), .B(n7324), .ZN(n7327)
         );
  INV_X1 U9124 ( .A(n7327), .ZN(P2_U3191) );
  INV_X1 U9125 ( .A(n7328), .ZN(n7343) );
  OAI222_X1 U9126 ( .A1(n7730), .A2(n7343), .B1(P2_U3151), .B2(n8090), .C1(
        n7329), .C2(n8577), .ZN(P2_U3275) );
  OAI21_X1 U9127 ( .B1(n7332), .B2(n7330), .A(n7331), .ZN(n7340) );
  NAND2_X1 U9128 ( .A1(n8741), .A2(n9779), .ZN(n7338) );
  NOR2_X1 U9129 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7333), .ZN(n9104) );
  AOI21_X1 U9130 ( .B1(n8726), .B2(n9032), .A(n9104), .ZN(n7337) );
  NAND2_X1 U9131 ( .A1(n8763), .A2(n7334), .ZN(n7336) );
  NAND2_X1 U9132 ( .A1(n8757), .A2(n9034), .ZN(n7335) );
  NAND4_X1 U9133 ( .A1(n7338), .A2(n7337), .A3(n7336), .A4(n7335), .ZN(n7339)
         );
  AOI21_X1 U9134 ( .B1(n7340), .B2(n8748), .A(n7339), .ZN(n7341) );
  INV_X1 U9135 ( .A(n7341), .ZN(P1_U3231) );
  OAI222_X1 U9136 ( .A1(n7522), .A2(n7344), .B1(n7708), .B2(n7343), .C1(
        P1_U3086), .C2(n7342), .ZN(P1_U3335) );
  INV_X1 U9137 ( .A(n7345), .ZN(n7380) );
  OAI222_X1 U9138 ( .A1(n7730), .A2(n7380), .B1(P2_U3151), .B2(n7347), .C1(
        n7346), .C2(n8577), .ZN(P2_U3274) );
  AOI21_X1 U9139 ( .B1(n7350), .B2(n7349), .A(n7348), .ZN(n7365) );
  AOI21_X1 U9140 ( .B1(n4421), .B2(n7352), .A(n7351), .ZN(n7353) );
  NOR2_X1 U9141 ( .A1(n7353), .A2(n9825), .ZN(n7363) );
  AOI21_X1 U9142 ( .B1(n7356), .B2(n7355), .A(n7354), .ZN(n7357) );
  OR2_X1 U9143 ( .A1(n7357), .A2(n9832), .ZN(n7360) );
  INV_X1 U9144 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7358) );
  NOR2_X1 U9145 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7358), .ZN(n7581) );
  AOI21_X1 U9146 ( .B1(n9840), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7581), .ZN(
        n7359) );
  OAI211_X1 U9147 ( .C1(n8246), .C2(n7361), .A(n7360), .B(n7359), .ZN(n7362)
         );
  NOR2_X1 U9148 ( .A1(n7363), .A2(n7362), .ZN(n7364) );
  OAI21_X1 U9149 ( .B1(n7365), .B2(n8249), .A(n7364), .ZN(P2_U3192) );
  NAND2_X1 U9150 ( .A1(n7366), .A2(n7908), .ZN(n8423) );
  NAND2_X1 U9151 ( .A1(n8423), .A2(n7367), .ZN(n8426) );
  NAND2_X1 U9152 ( .A1(n8426), .A2(n7368), .ZN(n7369) );
  XNOR2_X1 U9153 ( .A(n7369), .B(n7912), .ZN(n9887) );
  INV_X1 U9154 ( .A(n9887), .ZN(n7378) );
  OAI211_X1 U9155 ( .C1(n7371), .C2(n7912), .A(n7370), .B(n8436), .ZN(n7373)
         );
  AOI22_X1 U9156 ( .A1(n8433), .A2(n8123), .B1(n8122), .B2(n8430), .ZN(n7372)
         );
  NAND2_X1 U9157 ( .A1(n7373), .A2(n7372), .ZN(n9890) );
  NOR2_X1 U9158 ( .A1(n8429), .A2(n9888), .ZN(n7376) );
  OAI22_X1 U9159 ( .A1(n8398), .A2(n7374), .B1(n7445), .B2(n8427), .ZN(n7375)
         );
  AOI211_X1 U9160 ( .C1(n9890), .C2(n8398), .A(n7376), .B(n7375), .ZN(n7377)
         );
  OAI21_X1 U9161 ( .B1(n7378), .B2(n8386), .A(n7377), .ZN(P2_U3225) );
  OAI222_X1 U9162 ( .A1(n7522), .A2(n7381), .B1(n7708), .B2(n7380), .C1(
        P1_U3086), .C2(n7379), .ZN(P1_U3334) );
  AOI21_X1 U9163 ( .B1(n7384), .B2(n7383), .A(n7382), .ZN(n7399) );
  INV_X1 U9164 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7390) );
  OAI21_X1 U9165 ( .B1(n7387), .B2(n7386), .A(n7385), .ZN(n7388) );
  NAND2_X1 U9166 ( .A1(n7388), .A2(n9838), .ZN(n7389) );
  NAND2_X1 U9167 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7443) );
  OAI211_X1 U9168 ( .C1(n8255), .C2(n7390), .A(n7389), .B(n7443), .ZN(n7396)
         );
  AOI21_X1 U9169 ( .B1(n7393), .B2(n7392), .A(n7391), .ZN(n7394) );
  NOR2_X1 U9170 ( .A1(n7394), .A2(n9825), .ZN(n7395) );
  AOI211_X1 U9171 ( .C1(n9830), .C2(n7397), .A(n7396), .B(n7395), .ZN(n7398)
         );
  OAI21_X1 U9172 ( .B1(n7399), .B2(n9832), .A(n7398), .ZN(P2_U3190) );
  OR2_X1 U9173 ( .A1(n9519), .A2(n9508), .ZN(n8893) );
  NAND2_X1 U9174 ( .A1(n9519), .A2(n9508), .ZN(n8891) );
  NAND2_X1 U9175 ( .A1(n8893), .A2(n8891), .ZN(n7407) );
  INV_X1 U9176 ( .A(n8880), .ZN(n7400) );
  NOR2_X1 U9177 ( .A1(n7407), .A2(n7400), .ZN(n7401) );
  INV_X1 U9178 ( .A(n7485), .ZN(n7404) );
  INV_X1 U9179 ( .A(n7407), .ZN(n8973) );
  AOI21_X1 U9180 ( .B1(n7402), .B2(n8880), .A(n8973), .ZN(n7403) );
  NOR2_X1 U9181 ( .A1(n7404), .A2(n7403), .ZN(n9522) );
  INV_X1 U9182 ( .A(n9531), .ZN(n9030) );
  OAI21_X1 U9183 ( .B1(n7408), .B2(n7407), .A(n7489), .ZN(n9515) );
  NAND2_X1 U9184 ( .A1(n9515), .A2(n9742), .ZN(n7415) );
  AOI211_X1 U9185 ( .C1(n9519), .C2(n7409), .A(n9771), .B(n4403), .ZN(n9517)
         );
  INV_X1 U9186 ( .A(n9519), .ZN(n8708) );
  AOI22_X1 U9187 ( .A1(n4322), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8705), .B2(
        n9722), .ZN(n7410) );
  OAI21_X1 U9188 ( .B1(n9377), .B2(n9516), .A(n7410), .ZN(n7411) );
  AOI21_X1 U9189 ( .B1(n9380), .B2(n9030), .A(n7411), .ZN(n7412) );
  OAI21_X1 U9190 ( .B1(n8708), .B2(n9738), .A(n7412), .ZN(n7413) );
  AOI21_X1 U9191 ( .B1(n9517), .B2(n9724), .A(n7413), .ZN(n7414) );
  OAI211_X1 U9192 ( .C1(n9522), .C2(n9386), .A(n7415), .B(n7414), .ZN(P1_U3280) );
  NAND2_X1 U9193 ( .A1(n7417), .A2(n7416), .ZN(n7419) );
  AND2_X1 U9194 ( .A1(n7419), .A2(n7418), .ZN(n7423) );
  INV_X1 U9195 ( .A(n7464), .ZN(n7422) );
  AOI21_X1 U9196 ( .B1(n7424), .B2(n7423), .A(n7422), .ZN(n9898) );
  INV_X1 U9197 ( .A(n9898), .ZN(n7435) );
  XNOR2_X1 U9198 ( .A(n7425), .B(n7424), .ZN(n7429) );
  OAI22_X1 U9199 ( .A1(n7426), .A2(n8390), .B1(n7549), .B2(n8392), .ZN(n7427)
         );
  AOI21_X1 U9200 ( .B1(n9898), .B2(n7469), .A(n7427), .ZN(n7428) );
  OAI21_X1 U9201 ( .B1(n9845), .B2(n7429), .A(n7428), .ZN(n9896) );
  NAND2_X1 U9202 ( .A1(n9896), .A2(n8398), .ZN(n7433) );
  OAI22_X1 U9203 ( .A1(n8398), .A2(n7430), .B1(n7550), .B2(n8427), .ZN(n7431)
         );
  AOI21_X1 U9204 ( .B1(n8382), .B2(n7541), .A(n7431), .ZN(n7432) );
  OAI211_X1 U9205 ( .C1(n7435), .C2(n7434), .A(n7433), .B(n7432), .ZN(P2_U3224) );
  XOR2_X1 U9206 ( .A(n7436), .B(n7437), .Z(n7441) );
  NAND2_X1 U9207 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7617) );
  OAI21_X1 U9208 ( .B1(n7860), .B2(n7549), .A(n7617), .ZN(n7439) );
  OAI22_X1 U9209 ( .A1(n7514), .A2(n7861), .B1(n7874), .B2(n7994), .ZN(n7438)
         );
  AOI211_X1 U9210 ( .C1(n7513), .C2(n7876), .A(n7439), .B(n7438), .ZN(n7440)
         );
  OAI21_X1 U9211 ( .B1(n7441), .B2(n7879), .A(n7440), .ZN(P2_U3176) );
  XNOR2_X1 U9212 ( .A(n7544), .B(n7543), .ZN(n7442) );
  NOR2_X1 U9213 ( .A1(n7442), .A2(n8431), .ZN(n7542) );
  AOI21_X1 U9214 ( .B1(n8431), .B2(n7442), .A(n7542), .ZN(n7451) );
  INV_X1 U9215 ( .A(n7443), .ZN(n7447) );
  OAI22_X1 U9216 ( .A1(n7445), .A2(n7861), .B1(n7860), .B2(n7444), .ZN(n7446)
         );
  AOI211_X1 U9217 ( .C1(n7864), .C2(n8122), .A(n7447), .B(n7446), .ZN(n7450)
         );
  NAND2_X1 U9218 ( .A1(n7876), .A2(n7448), .ZN(n7449) );
  OAI211_X1 U9219 ( .C1(n7451), .C2(n7879), .A(n7450), .B(n7449), .ZN(P2_U3161) );
  INV_X1 U9220 ( .A(n7452), .ZN(n7483) );
  OAI222_X1 U9221 ( .A1(n7730), .A2(n7483), .B1(P2_U3151), .B2(n7454), .C1(
        n7453), .C2(n8577), .ZN(P2_U3271) );
  NAND2_X1 U9222 ( .A1(n7457), .A2(n9568), .ZN(n7455) );
  OAI211_X1 U9223 ( .C1(n7456), .C2(n7522), .A(n7455), .B(n9024), .ZN(P1_U3332) );
  NAND2_X1 U9224 ( .A1(n7457), .A2(n8581), .ZN(n7459) );
  OR2_X1 U9225 ( .A1(n7458), .A2(P2_U3151), .ZN(n8103) );
  OAI211_X1 U9226 ( .C1(n7460), .C2(n8577), .A(n7459), .B(n8103), .ZN(P2_U3272) );
  XNOR2_X1 U9227 ( .A(n7461), .B(n7915), .ZN(n7462) );
  NAND2_X1 U9228 ( .A1(n7462), .A2(n8436), .ZN(n7471) );
  NAND2_X1 U9229 ( .A1(n7464), .A2(n7463), .ZN(n7466) );
  INV_X1 U9230 ( .A(n7915), .ZN(n7465) );
  XNOR2_X1 U9231 ( .A(n7466), .B(n7465), .ZN(n9902) );
  NAND2_X1 U9232 ( .A1(n8122), .A2(n8433), .ZN(n7467) );
  OAI21_X1 U9233 ( .B1(n7578), .B2(n8392), .A(n7467), .ZN(n7468) );
  AOI21_X1 U9234 ( .B1(n9902), .B2(n7469), .A(n7468), .ZN(n7470) );
  AND2_X1 U9235 ( .A1(n7471), .A2(n7470), .ZN(n9904) );
  OAI22_X1 U9236 ( .A1(n8398), .A2(n7472), .B1(n7579), .B2(n8427), .ZN(n7473)
         );
  AOI21_X1 U9237 ( .B1(n8382), .B2(n9899), .A(n7473), .ZN(n7475) );
  NAND2_X1 U9238 ( .A1(n9902), .A2(n8444), .ZN(n7474) );
  OAI211_X1 U9239 ( .C1(n9904), .C2(n8441), .A(n7475), .B(n7474), .ZN(P2_U3223) );
  INV_X1 U9240 ( .A(n7476), .ZN(n7498) );
  OAI222_X1 U9241 ( .A1(n7730), .A2(n7498), .B1(P2_U3151), .B2(n7477), .C1(
        n10066), .C2(n8577), .ZN(P2_U3270) );
  INV_X1 U9242 ( .A(n7478), .ZN(n7480) );
  OAI222_X1 U9243 ( .A1(n7728), .A2(n7479), .B1(n7730), .B2(n7480), .C1(n7932), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9244 ( .A1(n7522), .A2(n7481), .B1(n7708), .B2(n7480), .C1(n9010), 
        .C2(P1_U3086), .ZN(P1_U3333) );
  OAI222_X1 U9245 ( .A1(n7522), .A2(n7484), .B1(n7708), .B2(n7483), .C1(
        P1_U3086), .C2(n7482), .ZN(P1_U3331) );
  NAND2_X1 U9246 ( .A1(n9510), .A2(n9516), .ZN(n8816) );
  NAND2_X1 U9247 ( .A1(n8886), .A2(n8816), .ZN(n8884) );
  AOI21_X1 U9248 ( .B1(n7486), .B2(n8884), .A(n9523), .ZN(n7488) );
  NAND2_X1 U9249 ( .A1(n7488), .A2(n7558), .ZN(n9512) );
  INV_X1 U9250 ( .A(n9508), .ZN(n9029) );
  OAI21_X1 U9251 ( .B1(n7490), .B2(n8884), .A(n7564), .ZN(n9506) );
  NAND2_X1 U9252 ( .A1(n9506), .A2(n9742), .ZN(n7496) );
  NAND2_X1 U9253 ( .A1(n9380), .A2(n9029), .ZN(n7492) );
  AOI22_X1 U9254 ( .A1(n4322), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8593), .B2(
        n9722), .ZN(n7491) );
  OAI211_X1 U9255 ( .C1(n9507), .C2(n9377), .A(n7492), .B(n7491), .ZN(n7494)
         );
  INV_X1 U9256 ( .A(n9510), .ZN(n8596) );
  OAI211_X1 U9257 ( .C1(n4403), .C2(n8596), .A(n9452), .B(n7566), .ZN(n9511)
         );
  NOR2_X1 U9258 ( .A1(n9511), .A2(n9735), .ZN(n7493) );
  AOI211_X1 U9259 ( .C1(n9349), .C2(n9510), .A(n7494), .B(n7493), .ZN(n7495)
         );
  OAI211_X1 U9260 ( .C1(n4322), .C2(n9512), .A(n7496), .B(n7495), .ZN(P1_U3279) );
  OAI222_X1 U9261 ( .A1(n7522), .A2(n7499), .B1(n7708), .B2(n7498), .C1(
        P1_U3086), .C2(n7497), .ZN(P1_U3330) );
  INV_X1 U9262 ( .A(n7500), .ZN(n7520) );
  OAI222_X1 U9263 ( .A1(n7730), .A2(n7520), .B1(P2_U3151), .B2(n7502), .C1(
        n7501), .C2(n8577), .ZN(P2_U3269) );
  OR2_X1 U9264 ( .A1(n7461), .A2(n7503), .ZN(n7506) );
  AND2_X1 U9265 ( .A1(n7506), .A2(n7504), .ZN(n7509) );
  NAND2_X1 U9266 ( .A1(n7506), .A2(n7505), .ZN(n7507) );
  OAI211_X1 U9267 ( .C1(n7509), .C2(n7508), .A(n8436), .B(n7507), .ZN(n7511)
         );
  AOI22_X1 U9268 ( .A1(n8430), .A2(n8119), .B1(n8121), .B2(n8433), .ZN(n7510)
         );
  NAND2_X1 U9269 ( .A1(n7511), .A2(n7510), .ZN(n7589) );
  INV_X1 U9270 ( .A(n7589), .ZN(n7518) );
  XNOR2_X1 U9271 ( .A(n7512), .B(n7916), .ZN(n7590) );
  INV_X1 U9272 ( .A(n7513), .ZN(n7595) );
  NOR2_X1 U9273 ( .A1(n7595), .A2(n8429), .ZN(n7516) );
  OAI22_X1 U9274 ( .A1(n8398), .A2(n7609), .B1(n7514), .B2(n8427), .ZN(n7515)
         );
  AOI211_X1 U9275 ( .C1(n7590), .C2(n8419), .A(n7516), .B(n7515), .ZN(n7517)
         );
  OAI21_X1 U9276 ( .B1(n7518), .B2(n8418), .A(n7517), .ZN(P2_U3222) );
  OAI222_X1 U9277 ( .A1(n7522), .A2(n7521), .B1(n7708), .B2(n7520), .C1(
        P1_U3086), .C2(n7519), .ZN(P1_U3329) );
  NAND2_X1 U9278 ( .A1(n7524), .A2(n7523), .ZN(n7526) );
  XOR2_X1 U9279 ( .A(n7526), .B(n7525), .Z(n7533) );
  OAI22_X1 U9280 ( .A1(n7640), .A2(n7861), .B1(n7874), .B2(n7629), .ZN(n7530)
         );
  NOR2_X1 U9281 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7527), .ZN(n8143) );
  INV_X1 U9282 ( .A(n8143), .ZN(n7528) );
  OAI21_X1 U9283 ( .B1(n7860), .B2(n7578), .A(n7528), .ZN(n7529) );
  NOR2_X1 U9284 ( .A1(n7530), .A2(n7529), .ZN(n7532) );
  NAND2_X1 U9285 ( .A1(n8509), .A2(n7876), .ZN(n7531) );
  OAI211_X1 U9286 ( .C1(n7533), .C2(n7879), .A(n7532), .B(n7531), .ZN(P2_U3164) );
  XNOR2_X1 U9287 ( .A(n7534), .B(n7629), .ZN(n7535) );
  XNOR2_X1 U9288 ( .A(n7536), .B(n7535), .ZN(n7540) );
  NAND2_X1 U9289 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8152) );
  OAI21_X1 U9290 ( .B1(n7874), .B2(n7660), .A(n8152), .ZN(n7538) );
  OAI22_X1 U9291 ( .A1(n7600), .A2(n7861), .B1(n7860), .B2(n7994), .ZN(n7537)
         );
  AOI211_X1 U9292 ( .C1(n7599), .C2(n7876), .A(n7538), .B(n7537), .ZN(n7539)
         );
  OAI21_X1 U9293 ( .B1(n7540), .B2(n7879), .A(n7539), .ZN(P2_U3174) );
  INV_X1 U9294 ( .A(n7541), .ZN(n9895) );
  AOI21_X1 U9295 ( .B1(n7544), .B2(n7543), .A(n7542), .ZN(n7548) );
  XNOR2_X1 U9296 ( .A(n7546), .B(n7545), .ZN(n7547) );
  NAND2_X1 U9297 ( .A1(n7548), .A2(n7547), .ZN(n7574) );
  OAI211_X1 U9298 ( .C1(n7548), .C2(n7547), .A(n7574), .B(n7856), .ZN(n7554)
         );
  OAI22_X1 U9299 ( .A1(n7550), .A2(n7861), .B1(n7874), .B2(n7549), .ZN(n7551)
         );
  AOI211_X1 U9300 ( .C1(n7870), .C2(n8431), .A(n7552), .B(n7551), .ZN(n7553)
         );
  OAI211_X1 U9301 ( .C1(n9895), .C2(n7867), .A(n7554), .B(n7553), .ZN(P2_U3171) );
  INV_X1 U9302 ( .A(n7555), .ZN(n7597) );
  AOI21_X1 U9303 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n7587), .A(n7556), .ZN(
        n7557) );
  OAI21_X1 U9304 ( .B1(n7597), .B2(n7730), .A(n7557), .ZN(P2_U3268) );
  XNOR2_X1 U9305 ( .A(n9502), .B(n9507), .ZN(n8975) );
  NAND2_X1 U9306 ( .A1(n7558), .A2(n8886), .ZN(n7562) );
  INV_X1 U9307 ( .A(n7562), .ZN(n7560) );
  NAND2_X1 U9308 ( .A1(n7560), .A2(n7559), .ZN(n8985) );
  INV_X1 U9309 ( .A(n8985), .ZN(n7561) );
  AOI21_X1 U9310 ( .B1(n8975), .B2(n7562), .A(n7561), .ZN(n9505) );
  INV_X1 U9311 ( .A(n9516), .ZN(n9028) );
  XNOR2_X1 U9312 ( .A(n9171), .B(n8975), .ZN(n9498) );
  NAND2_X1 U9313 ( .A1(n9498), .A2(n9742), .ZN(n7572) );
  INV_X1 U9314 ( .A(n9374), .ZN(n7565) );
  AOI211_X1 U9315 ( .C1(n9502), .C2(n7566), .A(n9771), .B(n7565), .ZN(n9500)
         );
  AOI22_X1 U9316 ( .A1(n4322), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8764), .B2(
        n9722), .ZN(n7567) );
  OAI21_X1 U9317 ( .B1(n9377), .B2(n9499), .A(n7567), .ZN(n7568) );
  AOI21_X1 U9318 ( .B1(n9380), .B2(n9028), .A(n7568), .ZN(n7569) );
  OAI21_X1 U9319 ( .B1(n9170), .B2(n9738), .A(n7569), .ZN(n7570) );
  AOI21_X1 U9320 ( .B1(n9500), .B2(n9724), .A(n7570), .ZN(n7571) );
  OAI211_X1 U9321 ( .C1(n9505), .C2(n9386), .A(n7572), .B(n7571), .ZN(P1_U3278) );
  NAND2_X1 U9322 ( .A1(n7574), .A2(n7573), .ZN(n7577) );
  XNOR2_X1 U9323 ( .A(n7575), .B(n8121), .ZN(n7576) );
  XNOR2_X1 U9324 ( .A(n7577), .B(n7576), .ZN(n7584) );
  OAI22_X1 U9325 ( .A1(n7579), .A2(n7861), .B1(n7874), .B2(n7578), .ZN(n7580)
         );
  AOI211_X1 U9326 ( .C1(n7870), .C2(n8122), .A(n7581), .B(n7580), .ZN(n7583)
         );
  NAND2_X1 U9327 ( .A1(n9899), .A2(n7876), .ZN(n7582) );
  OAI211_X1 U9328 ( .C1(n7584), .C2(n7879), .A(n7583), .B(n7582), .ZN(P2_U3157) );
  INV_X1 U9329 ( .A(n7585), .ZN(n7655) );
  AOI21_X1 U9330 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n7587), .A(n7586), .ZN(
        n7588) );
  OAI21_X1 U9331 ( .B1(n7655), .B2(n7730), .A(n7588), .ZN(P2_U3267) );
  AOI21_X1 U9332 ( .B1(n7590), .B2(n6266), .A(n7589), .ZN(n7592) );
  MUX2_X1 U9333 ( .A(n7606), .B(n7592), .S(n9920), .Z(n7591) );
  OAI21_X1 U9334 ( .B1(n7595), .B2(n8508), .A(n7591), .ZN(P2_U3470) );
  INV_X1 U9335 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7593) );
  MUX2_X1 U9336 ( .A(n7593), .B(n7592), .S(n9905), .Z(n7594) );
  OAI21_X1 U9337 ( .B1(n7595), .B2(n8570), .A(n7594), .ZN(P2_U3423) );
  OAI222_X1 U9338 ( .A1(P1_U3086), .A2(n6711), .B1(n7708), .B2(n7597), .C1(
        n7596), .C2(n7522), .ZN(P1_U3328) );
  NAND2_X1 U9339 ( .A1(n8405), .A2(n8403), .ZN(n7997) );
  XNOR2_X1 U9340 ( .A(n8404), .B(n7997), .ZN(n7598) );
  OAI222_X1 U9341 ( .A1(n8390), .A2(n7994), .B1(n8392), .B2(n7660), .C1(n7598), 
        .C2(n9845), .ZN(n8504) );
  INV_X1 U9342 ( .A(n7599), .ZN(n8571) );
  OAI22_X1 U9343 ( .A1(n8571), .A2(n8413), .B1(n7600), .B2(n8427), .ZN(n7601)
         );
  OAI21_X1 U9344 ( .B1(n8504), .B2(n7601), .A(n8398), .ZN(n7604) );
  XOR2_X1 U9345 ( .A(n7997), .B(n7602), .Z(n8505) );
  AOI22_X1 U9346 ( .A1(n8505), .A2(n8419), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8418), .ZN(n7603) );
  NAND2_X1 U9347 ( .A1(n7604), .A2(n7603), .ZN(P2_U3220) );
  AOI21_X1 U9348 ( .B1(n7607), .B2(n7606), .A(n7605), .ZN(n7624) );
  INV_X1 U9349 ( .A(n8133), .ZN(n7608) );
  AOI21_X1 U9350 ( .B1(n7610), .B2(n7609), .A(n7608), .ZN(n7611) );
  NOR2_X1 U9351 ( .A1(n7611), .A2(n9832), .ZN(n7622) );
  NOR2_X1 U9352 ( .A1(n8246), .A2(n7612), .ZN(n7621) );
  INV_X1 U9353 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7613) );
  NOR2_X1 U9354 ( .A1(n8255), .A2(n7613), .ZN(n7620) );
  AOI21_X1 U9355 ( .B1(n7616), .B2(n7615), .A(n7614), .ZN(n7618) );
  OAI21_X1 U9356 ( .B1(n7618), .B2(n8249), .A(n7617), .ZN(n7619) );
  NOR4_X1 U9357 ( .A1(n7622), .A2(n7621), .A3(n7620), .A4(n7619), .ZN(n7623)
         );
  OAI21_X1 U9358 ( .B1(n7624), .B2(n9825), .A(n7623), .ZN(P2_U3193) );
  INV_X1 U9359 ( .A(n8500), .ZN(n8414) );
  OAI21_X1 U9360 ( .B1(n7627), .B2(n7626), .A(n7625), .ZN(n7628) );
  NAND2_X1 U9361 ( .A1(n7628), .A2(n7856), .ZN(n7633) );
  NAND2_X1 U9362 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8173) );
  INV_X1 U9363 ( .A(n8173), .ZN(n7631) );
  OAI22_X1 U9364 ( .A1(n8412), .A2(n7861), .B1(n7860), .B2(n7629), .ZN(n7630)
         );
  AOI211_X1 U9365 ( .C1(n7864), .C2(n8410), .A(n7631), .B(n7630), .ZN(n7632)
         );
  OAI211_X1 U9366 ( .C1(n8414), .C2(n7867), .A(n7633), .B(n7632), .ZN(P2_U3155) );
  INV_X1 U9367 ( .A(n7634), .ZN(n7635) );
  AOI21_X1 U9368 ( .B1(n7637), .B2(n7636), .A(n7635), .ZN(n8510) );
  INV_X1 U9369 ( .A(n8510), .ZN(n7644) );
  INV_X1 U9370 ( .A(n7637), .ZN(n7991) );
  XNOR2_X1 U9371 ( .A(n7638), .B(n7991), .ZN(n7639) );
  AOI222_X1 U9372 ( .A1(n8436), .A2(n7639), .B1(n8120), .B2(n8433), .C1(n8409), 
        .C2(n8430), .ZN(n8512) );
  OAI21_X1 U9373 ( .B1(n7640), .B2(n8427), .A(n8512), .ZN(n7641) );
  NAND2_X1 U9374 ( .A1(n7641), .A2(n8398), .ZN(n7643) );
  AOI22_X1 U9375 ( .A1(n8509), .A2(n8382), .B1(P2_REG2_REG_12__SCAN_IN), .B2(
        n8418), .ZN(n7642) );
  OAI211_X1 U9376 ( .C1(n7644), .C2(n8386), .A(n7643), .B(n7642), .ZN(P2_U3221) );
  INV_X1 U9377 ( .A(n7645), .ZN(n8565) );
  AOI21_X1 U9378 ( .B1(n7647), .B2(n7646), .A(n7879), .ZN(n7649) );
  NAND2_X1 U9379 ( .A1(n7649), .A2(n7648), .ZN(n7653) );
  NAND2_X1 U9380 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8193) );
  INV_X1 U9381 ( .A(n8193), .ZN(n7651) );
  OAI22_X1 U9382 ( .A1(n7662), .A2(n7861), .B1(n7860), .B2(n7660), .ZN(n7650)
         );
  AOI211_X1 U9383 ( .C1(n7864), .C2(n8117), .A(n7651), .B(n7650), .ZN(n7652)
         );
  OAI211_X1 U9384 ( .C1(n8565), .C2(n7867), .A(n7653), .B(n7652), .ZN(P2_U3181) );
  OAI222_X1 U9385 ( .A1(P1_U3086), .A2(n5740), .B1(n7708), .B2(n7655), .C1(
        n7654), .C2(n7522), .ZN(P1_U3327) );
  NAND2_X1 U9386 ( .A1(n7657), .A2(n7656), .ZN(n7658) );
  XNOR2_X1 U9387 ( .A(n7658), .B(n8002), .ZN(n7659) );
  OAI222_X1 U9388 ( .A1(n8392), .A2(n8374), .B1(n8390), .B2(n7660), .C1(n9845), 
        .C2(n7659), .ZN(n8496) );
  INV_X1 U9389 ( .A(n8496), .ZN(n7666) );
  XNOR2_X1 U9390 ( .A(n7661), .B(n8002), .ZN(n8497) );
  NOR2_X1 U9391 ( .A1(n8565), .A2(n8429), .ZN(n7664) );
  OAI22_X1 U9392 ( .A1(n8398), .A2(n8191), .B1(n7662), .B2(n8427), .ZN(n7663)
         );
  AOI211_X1 U9393 ( .C1(n8497), .C2(n8419), .A(n7664), .B(n7663), .ZN(n7665)
         );
  OAI21_X1 U9394 ( .B1(n7666), .B2(n8418), .A(n7665), .ZN(P2_U3218) );
  OAI21_X1 U9395 ( .B1(n7669), .B2(n7668), .A(n7667), .ZN(n7670) );
  NAND2_X1 U9396 ( .A1(n7670), .A2(n7856), .ZN(n7674) );
  AND2_X1 U9397 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9828) );
  OAI22_X1 U9398 ( .A1(n8428), .A2(n7861), .B1(n7860), .B2(n7671), .ZN(n7672)
         );
  AOI211_X1 U9399 ( .C1(n7864), .C2(n8431), .A(n9828), .B(n7672), .ZN(n7673)
         );
  OAI211_X1 U9400 ( .C1(n9882), .C2(n7867), .A(n7674), .B(n7673), .ZN(P2_U3153) );
  NAND2_X1 U9401 ( .A1(n7676), .A2(n7675), .ZN(n7677) );
  INV_X1 U9402 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8774) );
  INV_X1 U9403 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n10039) );
  MUX2_X1 U9404 ( .A(n8774), .B(n10039), .S(n4586), .Z(n7887) );
  XNOR2_X1 U9405 ( .A(n7887), .B(SI_30_), .ZN(n7884) );
  INV_X1 U9406 ( .A(n8773), .ZN(n7707) );
  OAI222_X1 U9407 ( .A1(n7730), .A2(n7707), .B1(n7679), .B2(P2_U3151), .C1(
        n10039), .C2(n7728), .ZN(P2_U3265) );
  NOR2_X1 U9408 ( .A1(n9366), .A2(n7680), .ZN(n7684) );
  AND4_X1 U9409 ( .A1(n9366), .A2(n8955), .A3(n7682), .A4(n7681), .ZN(n7683)
         );
  AOI211_X1 U9410 ( .C1(n9722), .C2(P1_REG3_REG_0__SCAN_IN), .A(n7684), .B(
        n7683), .ZN(n7686) );
  OAI21_X1 U9411 ( .B1(n9349), .B2(n9303), .A(n7688), .ZN(n7685) );
  OAI211_X1 U9412 ( .C1(n7687), .C2(n9377), .A(n7686), .B(n7685), .ZN(P1_U3293) );
  AOI22_X1 U9413 ( .A1(n8741), .A2(n7688), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n7698), .ZN(n7691) );
  AOI22_X1 U9414 ( .A1(n8726), .A2(n9041), .B1(n7689), .B2(n8748), .ZN(n7690)
         );
  NAND2_X1 U9415 ( .A1(n7691), .A2(n7690), .ZN(P1_U3232) );
  INV_X1 U9416 ( .A(n7692), .ZN(n7693) );
  NOR2_X1 U9417 ( .A1(n7694), .A2(n7693), .ZN(n7697) );
  INV_X1 U9418 ( .A(n7695), .ZN(n7696) );
  AOI21_X1 U9419 ( .B1(n7697), .B2(n6627), .A(n7696), .ZN(n7702) );
  AOI22_X1 U9420 ( .A1(n8726), .A2(n9039), .B1(n8757), .B2(n9041), .ZN(n7701)
         );
  AOI22_X1 U9421 ( .A1(n8741), .A2(n7699), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n7698), .ZN(n7700) );
  OAI211_X1 U9422 ( .C1(n7702), .C2(n8766), .A(n7701), .B(n7700), .ZN(P1_U3237) );
  INV_X1 U9423 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7704) );
  OAI222_X1 U9424 ( .A1(n7703), .A2(P1_U3086), .B1(n7708), .B2(n7705), .C1(
        n7704), .C2(n7522), .ZN(P1_U3336) );
  OAI222_X1 U9425 ( .A1(P1_U3086), .A2(n7706), .B1(n7708), .B2(n7707), .C1(
        n8774), .C2(n7522), .ZN(P1_U3325) );
  INV_X1 U9426 ( .A(n7710), .ZN(n7778) );
  OAI22_X1 U9427 ( .A1(n7778), .A2(n8427), .B1(n8398), .B2(n7711), .ZN(n7714)
         );
  NOR2_X1 U9428 ( .A1(n7712), .A2(n8386), .ZN(n7713) );
  AOI211_X1 U9429 ( .C1(n8382), .C2(n7782), .A(n7714), .B(n7713), .ZN(n7715)
         );
  OAI21_X1 U9430 ( .B1(n7709), .B2(n8418), .A(n7715), .ZN(P2_U3205) );
  NAND2_X1 U9431 ( .A1(n8773), .A2(n7893), .ZN(n7717) );
  OR2_X1 U9432 ( .A1(n5849), .A2(n10039), .ZN(n7716) );
  INV_X1 U9433 ( .A(n7718), .ZN(n7719) );
  NOR2_X1 U9434 ( .A1(n8093), .A2(n7719), .ZN(n8514) );
  NOR2_X1 U9435 ( .A1(n7720), .A2(n8427), .ZN(n7722) );
  AOI21_X1 U9436 ( .B1(n8514), .B2(n8398), .A(n7722), .ZN(n8260) );
  NAND2_X1 U9437 ( .A1(n8441), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7721) );
  OAI211_X1 U9438 ( .C1(n7896), .C2(n8429), .A(n8260), .B(n7721), .ZN(P2_U3203) );
  AOI21_X1 U9439 ( .B1(n8441), .B2(P2_REG2_REG_29__SCAN_IN), .A(n7722), .ZN(
        n7723) );
  OAI21_X1 U9440 ( .B1(n7724), .B2(n8429), .A(n7723), .ZN(n7725) );
  AOI21_X1 U9441 ( .B1(n6218), .B2(n8444), .A(n7725), .ZN(n7726) );
  OAI21_X1 U9442 ( .B1(n7727), .B2(n8418), .A(n7726), .ZN(P2_U3204) );
  INV_X1 U9443 ( .A(n8793), .ZN(n9571) );
  OAI222_X1 U9444 ( .A1(n7730), .A2(n9571), .B1(n5815), .B2(P2_U3151), .C1(
        n7729), .C2(n7728), .ZN(P2_U3266) );
  XNOR2_X1 U9445 ( .A(n7836), .B(n4319), .ZN(n7731) );
  NAND2_X1 U9446 ( .A1(n7731), .A2(n8346), .ZN(n7787) );
  INV_X1 U9447 ( .A(n7731), .ZN(n7732) );
  NAND2_X1 U9448 ( .A1(n7732), .A2(n8113), .ZN(n7733) );
  NAND2_X1 U9449 ( .A1(n7787), .A2(n7733), .ZN(n7832) );
  INV_X1 U9450 ( .A(n7734), .ZN(n7735) );
  AND2_X1 U9451 ( .A1(n7735), .A2(n8114), .ZN(n7833) );
  NOR2_X1 U9452 ( .A1(n7832), .A2(n7833), .ZN(n7736) );
  NAND2_X1 U9453 ( .A1(n7737), .A2(n7736), .ZN(n7785) );
  XNOR2_X1 U9454 ( .A(n7738), .B(n7749), .ZN(n7740) );
  XNOR2_X1 U9455 ( .A(n7740), .B(n8336), .ZN(n7786) );
  INV_X1 U9456 ( .A(n7740), .ZN(n7741) );
  NAND2_X1 U9457 ( .A1(n7741), .A2(n8336), .ZN(n7742) );
  XNOR2_X1 U9458 ( .A(n7841), .B(n7774), .ZN(n7743) );
  XNOR2_X1 U9459 ( .A(n7743), .B(n8322), .ZN(n7842) );
  INV_X1 U9460 ( .A(n7743), .ZN(n7744) );
  XNOR2_X1 U9461 ( .A(n7767), .B(n7774), .ZN(n7794) );
  XNOR2_X1 U9462 ( .A(n8532), .B(n4319), .ZN(n7745) );
  NAND2_X1 U9463 ( .A1(n7745), .A2(n8110), .ZN(n7797) );
  OAI21_X1 U9464 ( .B1(n8312), .B2(n7794), .A(n7797), .ZN(n7748) );
  INV_X1 U9465 ( .A(n7745), .ZN(n7746) );
  NAND2_X1 U9466 ( .A1(n7746), .A2(n8302), .ZN(n7798) );
  NAND3_X1 U9467 ( .A1(n7797), .A2(n8312), .A3(n7794), .ZN(n7747) );
  OAI211_X1 U9468 ( .C1(n7762), .C2(n7748), .A(n7798), .B(n7747), .ZN(n7750)
         );
  XNOR2_X1 U9469 ( .A(n7804), .B(n7749), .ZN(n7751) );
  XNOR2_X1 U9470 ( .A(n7751), .B(n8293), .ZN(n7799) );
  NAND2_X1 U9471 ( .A1(n7750), .A2(n7799), .ZN(n7801) );
  INV_X1 U9472 ( .A(n8293), .ZN(n8109) );
  NOR2_X1 U9473 ( .A1(n7868), .A2(n8108), .ZN(n7869) );
  XNOR2_X1 U9474 ( .A(n7754), .B(n4318), .ZN(n7770) );
  XNOR2_X1 U9475 ( .A(n7770), .B(n8107), .ZN(n7755) );
  NAND2_X1 U9476 ( .A1(n7756), .A2(n7755), .ZN(n7773) );
  OAI211_X1 U9477 ( .C1(n7756), .C2(n7755), .A(n7773), .B(n7856), .ZN(n7761)
         );
  INV_X1 U9478 ( .A(n8264), .ZN(n7758) );
  AOI22_X1 U9479 ( .A1(n8108), .A2(n7870), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7757) );
  OAI21_X1 U9480 ( .B1(n7758), .B2(n7861), .A(n7757), .ZN(n7759) );
  AOI21_X1 U9481 ( .B1(n7864), .B2(n8106), .A(n7759), .ZN(n7760) );
  OAI211_X1 U9482 ( .C1(n8266), .C2(n7867), .A(n7761), .B(n7760), .ZN(P2_U3154) );
  XOR2_X1 U9483 ( .A(n7794), .B(n7762), .Z(n7796) );
  XNOR2_X1 U9484 ( .A(n7796), .B(n8312), .ZN(n7769) );
  INV_X1 U9485 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n7763) );
  OAI22_X1 U9486 ( .A1(n8302), .A2(n7874), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7763), .ZN(n7766) );
  INV_X1 U9487 ( .A(n8305), .ZN(n7764) );
  OAI22_X1 U9488 ( .A1(n7764), .A2(n7861), .B1(n7860), .B2(n8322), .ZN(n7765)
         );
  AOI211_X1 U9489 ( .C1(n7767), .C2(n7876), .A(n7766), .B(n7765), .ZN(n7768)
         );
  OAI21_X1 U9490 ( .B1(n7769), .B2(n7879), .A(n7768), .ZN(P2_U3156) );
  INV_X1 U9491 ( .A(n7770), .ZN(n7771) );
  NAND2_X1 U9492 ( .A1(n7771), .A2(n8107), .ZN(n7772) );
  NAND2_X1 U9493 ( .A1(n7773), .A2(n7772), .ZN(n7776) );
  XOR2_X1 U9494 ( .A(n7774), .B(n7928), .Z(n7775) );
  XNOR2_X1 U9495 ( .A(n7776), .B(n7775), .ZN(n7784) );
  INV_X1 U9496 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7777) );
  OAI22_X1 U9497 ( .A1(n7778), .A2(n7861), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7777), .ZN(n7781) );
  OAI22_X1 U9498 ( .A1(n7779), .A2(n7874), .B1(n8273), .B2(n7860), .ZN(n7780)
         );
  AOI211_X1 U9499 ( .C1(n7782), .C2(n7876), .A(n7781), .B(n7780), .ZN(n7783)
         );
  OAI21_X1 U9500 ( .B1(n7784), .B2(n7879), .A(n7783), .ZN(P2_U3160) );
  NAND3_X1 U9501 ( .A1(n7785), .A2(n4900), .A3(n7787), .ZN(n7788) );
  AOI21_X1 U9502 ( .B1(n7789), .B2(n7788), .A(n7879), .ZN(n7793) );
  AOI22_X1 U9503 ( .A1(n7864), .A2(n8112), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7791) );
  AOI22_X1 U9504 ( .A1(n8327), .A2(n7871), .B1(n7870), .B2(n8113), .ZN(n7790)
         );
  OAI211_X1 U9505 ( .C1(n8544), .C2(n7867), .A(n7791), .B(n7790), .ZN(n7792)
         );
  OR2_X1 U9506 ( .A1(n7793), .A2(n7792), .ZN(P2_U3163) );
  INV_X1 U9507 ( .A(n7762), .ZN(n7795) );
  OAI22_X1 U9508 ( .A1(n7796), .A2(n8312), .B1(n7795), .B2(n7794), .ZN(n7823)
         );
  NAND2_X1 U9509 ( .A1(n7797), .A2(n7798), .ZN(n7824) );
  NOR2_X1 U9510 ( .A1(n7823), .A2(n7824), .ZN(n7822) );
  INV_X1 U9511 ( .A(n7798), .ZN(n7800) );
  NOR3_X1 U9512 ( .A1(n7822), .A2(n7800), .A3(n7799), .ZN(n7803) );
  INV_X1 U9513 ( .A(n7801), .ZN(n7802) );
  OAI21_X1 U9514 ( .B1(n7803), .B2(n7802), .A(n7856), .ZN(n7808) );
  AOI22_X1 U9515 ( .A1(n8108), .A2(n7864), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7807) );
  AOI22_X1 U9516 ( .A1(n8110), .A2(n7870), .B1(n8285), .B2(n7871), .ZN(n7806)
         );
  NAND2_X1 U9517 ( .A1(n7804), .A2(n7876), .ZN(n7805) );
  NAND4_X1 U9518 ( .A1(n7808), .A2(n7807), .A3(n7806), .A4(n7805), .ZN(
        P2_U3165) );
  XNOR2_X1 U9519 ( .A(n7810), .B(n7809), .ZN(n7814) );
  NAND2_X1 U9520 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8208) );
  OAI21_X1 U9521 ( .B1(n7874), .B2(n8391), .A(n8208), .ZN(n7812) );
  OAI22_X1 U9522 ( .A1(n8396), .A2(n7861), .B1(n7860), .B2(n8389), .ZN(n7811)
         );
  AOI211_X1 U9523 ( .C1(n8395), .C2(n7876), .A(n7812), .B(n7811), .ZN(n7813)
         );
  OAI21_X1 U9524 ( .B1(n7814), .B2(n7879), .A(n7813), .ZN(P2_U3166) );
  INV_X1 U9525 ( .A(n7815), .ZN(n7854) );
  AOI21_X1 U9526 ( .B1(n7817), .B2(n7816), .A(n7854), .ZN(n7821) );
  NAND2_X1 U9527 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8228) );
  OAI21_X1 U9528 ( .B1(n7874), .B2(n8375), .A(n8228), .ZN(n7819) );
  OAI22_X1 U9529 ( .A1(n8379), .A2(n7861), .B1(n7860), .B2(n8374), .ZN(n7818)
         );
  AOI211_X1 U9530 ( .C1(n8383), .C2(n7876), .A(n7819), .B(n7818), .ZN(n7820)
         );
  OAI21_X1 U9531 ( .B1(n7821), .B2(n7879), .A(n7820), .ZN(P2_U3168) );
  AOI21_X1 U9532 ( .B1(n7824), .B2(n7823), .A(n7822), .ZN(n7831) );
  OAI22_X1 U9533 ( .A1(n8293), .A2(n7874), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7825), .ZN(n7828) );
  INV_X1 U9534 ( .A(n8295), .ZN(n7826) );
  OAI22_X1 U9535 ( .A1(n7826), .A2(n7861), .B1(n8312), .B2(n7860), .ZN(n7827)
         );
  AOI211_X1 U9536 ( .C1(n7829), .C2(n7876), .A(n7828), .B(n7827), .ZN(n7830)
         );
  OAI21_X1 U9537 ( .B1(n7831), .B2(n7879), .A(n7830), .ZN(P2_U3169) );
  OAI21_X1 U9538 ( .B1(n7834), .B2(n7833), .A(n7832), .ZN(n7835) );
  AOI21_X1 U9539 ( .B1(n7835), .B2(n7785), .A(n7879), .ZN(n7840) );
  INV_X1 U9540 ( .A(n7836), .ZN(n8548) );
  AOI22_X1 U9541 ( .A1(n7864), .A2(n6087), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7838) );
  AOI22_X1 U9542 ( .A1(n8339), .A2(n7871), .B1(n7870), .B2(n8114), .ZN(n7837)
         );
  OAI211_X1 U9543 ( .C1(n8548), .C2(n7867), .A(n7838), .B(n7837), .ZN(n7839)
         );
  OR2_X1 U9544 ( .A1(n7840), .A2(n7839), .ZN(P2_U3173) );
  INV_X1 U9545 ( .A(n7841), .ZN(n8540) );
  AOI21_X1 U9546 ( .B1(n7843), .B2(n7842), .A(n7879), .ZN(n7845) );
  NAND2_X1 U9547 ( .A1(n7845), .A2(n7844), .ZN(n7850) );
  NOR2_X1 U9548 ( .A1(n7860), .A2(n8336), .ZN(n7848) );
  INV_X1 U9549 ( .A(n8315), .ZN(n7846) );
  OAI22_X1 U9550 ( .A1(n8312), .A2(n7874), .B1(n7861), .B2(n7846), .ZN(n7847)
         );
  AOI211_X1 U9551 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3151), .A(n7848), 
        .B(n7847), .ZN(n7849) );
  OAI211_X1 U9552 ( .C1(n8540), .C2(n7867), .A(n7850), .B(n7849), .ZN(P2_U3175) );
  INV_X1 U9553 ( .A(n7851), .ZN(n7853) );
  NOR3_X1 U9554 ( .A1(n7854), .A2(n7853), .A3(n7852), .ZN(n7858) );
  INV_X1 U9555 ( .A(n7855), .ZN(n7857) );
  OAI21_X1 U9556 ( .B1(n7858), .B2(n7857), .A(n7856), .ZN(n7866) );
  NAND2_X1 U9557 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8254) );
  INV_X1 U9558 ( .A(n8254), .ZN(n7863) );
  OAI22_X1 U9559 ( .A1(n8363), .A2(n7861), .B1(n7860), .B2(n8391), .ZN(n7862)
         );
  AOI211_X1 U9560 ( .C1(n7864), .C2(n8114), .A(n7863), .B(n7862), .ZN(n7865)
         );
  OAI211_X1 U9561 ( .C1(n8556), .C2(n7867), .A(n7866), .B(n7865), .ZN(P2_U3178) );
  AOI21_X1 U9562 ( .B1(n8108), .B2(n7868), .A(n7869), .ZN(n7880) );
  AOI22_X1 U9563 ( .A1(n8109), .A2(n7870), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n7873) );
  NAND2_X1 U9564 ( .A1(n8276), .A2(n7871), .ZN(n7872) );
  OAI211_X1 U9565 ( .C1(n8273), .C2(n7874), .A(n7873), .B(n7872), .ZN(n7875)
         );
  AOI21_X1 U9566 ( .B1(n7877), .B2(n7876), .A(n7875), .ZN(n7878) );
  OAI21_X1 U9567 ( .B1(n7880), .B2(n7879), .A(n7878), .ZN(P2_U3180) );
  INV_X1 U9568 ( .A(n8105), .ZN(n7881) );
  NAND2_X1 U9569 ( .A1(n8518), .A2(n7881), .ZN(n8083) );
  NAND2_X1 U9570 ( .A1(n8083), .A2(n7882), .ZN(n8072) );
  INV_X1 U9571 ( .A(n7902), .ZN(n8081) );
  NAND2_X1 U9572 ( .A1(n7885), .A2(n7884), .ZN(n7889) );
  INV_X1 U9573 ( .A(SI_30_), .ZN(n7886) );
  NAND2_X1 U9574 ( .A1(n7887), .A2(n7886), .ZN(n7888) );
  NAND2_X1 U9575 ( .A1(n7889), .A2(n7888), .ZN(n7892) );
  INV_X1 U9576 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9565) );
  INV_X1 U9577 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8578) );
  MUX2_X1 U9578 ( .A(n9565), .B(n8578), .S(n4586), .Z(n7890) );
  XNOR2_X1 U9579 ( .A(n7890), .B(SI_31_), .ZN(n7891) );
  NAND2_X1 U9580 ( .A1(n9569), .A2(n7893), .ZN(n7895) );
  OR2_X1 U9581 ( .A1(n5849), .A2(n8578), .ZN(n7894) );
  OAI21_X1 U9582 ( .B1(n7897), .B2(n8081), .A(n8513), .ZN(n7899) );
  NAND3_X1 U9583 ( .A1(n7897), .A2(n8093), .A3(n7896), .ZN(n7898) );
  INV_X1 U9584 ( .A(n7900), .ZN(n8094) );
  NOR2_X1 U9585 ( .A1(n8513), .A2(n8093), .ZN(n8088) );
  NAND2_X1 U9586 ( .A1(n7902), .A2(n7901), .ZN(n8071) );
  NOR2_X1 U9587 ( .A1(n8088), .A2(n8071), .ZN(n7930) );
  INV_X1 U9588 ( .A(n7903), .ZN(n8061) );
  OR2_X1 U9589 ( .A1(n8067), .A2(n8274), .ZN(n8058) );
  INV_X1 U9590 ( .A(n8045), .ZN(n8049) );
  INV_X1 U9591 ( .A(n8038), .ZN(n8044) );
  INV_X1 U9592 ( .A(n7904), .ZN(n8325) );
  INV_X1 U9593 ( .A(n8362), .ZN(n7923) );
  NOR2_X1 U9594 ( .A1(n7906), .A2(n7905), .ZN(n7910) );
  NOR2_X1 U9595 ( .A1(n7907), .A2(n6181), .ZN(n7909) );
  NAND4_X1 U9596 ( .A1(n7910), .A2(n7909), .A3(n4481), .A4(n7908), .ZN(n7914)
         );
  INV_X1 U9597 ( .A(n7911), .ZN(n7913) );
  NOR4_X1 U9598 ( .A1(n7914), .A2(n7913), .A3(n7912), .A4(n8434), .ZN(n7917)
         );
  AND4_X1 U9599 ( .A1(n7917), .A2(n7972), .A3(n7916), .A4(n7915), .ZN(n7918)
         );
  NAND3_X1 U9600 ( .A1(n7997), .A2(n7918), .A3(n7991), .ZN(n7919) );
  NOR2_X1 U9601 ( .A1(n8407), .A2(n7919), .ZN(n7920) );
  NAND2_X1 U9602 ( .A1(n8002), .A2(n7920), .ZN(n7921) );
  NOR2_X1 U9603 ( .A1(n8393), .A2(n7921), .ZN(n7922) );
  NAND4_X1 U9604 ( .A1(n8349), .A2(n8370), .A3(n7923), .A4(n7922), .ZN(n7924)
         );
  NOR2_X1 U9605 ( .A1(n8337), .A2(n7924), .ZN(n7925) );
  NAND3_X1 U9606 ( .A1(n8313), .A2(n8325), .A3(n7925), .ZN(n7926) );
  OR4_X1 U9607 ( .A1(n8290), .A2(n8286), .A3(n8303), .A4(n7926), .ZN(n7927) );
  NOR4_X1 U9608 ( .A1(n8072), .A2(n7928), .A3(n8058), .A4(n7927), .ZN(n7929)
         );
  AOI21_X1 U9609 ( .B1(n7930), .B2(n7929), .A(n7933), .ZN(n8092) );
  INV_X1 U9610 ( .A(n7931), .ZN(n8005) );
  MUX2_X1 U9611 ( .A(n8118), .B(n8500), .S(n8085), .Z(n8004) );
  NAND2_X1 U9612 ( .A1(n7939), .A2(n7932), .ZN(n7934) );
  INV_X1 U9613 ( .A(n7936), .ZN(n7937) );
  INV_X1 U9614 ( .A(n7939), .ZN(n7940) );
  NOR2_X1 U9615 ( .A1(n6181), .A2(n7940), .ZN(n7941) );
  AOI21_X1 U9616 ( .B1(n7942), .B2(n7941), .A(n7907), .ZN(n7943) );
  NAND2_X1 U9617 ( .A1(n7962), .A2(n6184), .ZN(n7946) );
  NAND2_X1 U9618 ( .A1(n7950), .A2(n7944), .ZN(n7945) );
  MUX2_X1 U9619 ( .A(n7946), .B(n7945), .S(n8085), .Z(n7947) );
  INV_X1 U9620 ( .A(n7947), .ZN(n7949) );
  NAND2_X1 U9621 ( .A1(n7963), .A2(n7950), .ZN(n7958) );
  NAND2_X1 U9622 ( .A1(n8422), .A2(n7951), .ZN(n7965) );
  INV_X1 U9623 ( .A(n7952), .ZN(n7953) );
  NOR2_X1 U9624 ( .A1(n7965), .A2(n7953), .ZN(n7957) );
  NAND2_X1 U9625 ( .A1(n8124), .A2(n9870), .ZN(n7959) );
  INV_X1 U9626 ( .A(n7959), .ZN(n7954) );
  NAND2_X1 U9627 ( .A1(n7954), .A2(n8422), .ZN(n7955) );
  NAND2_X1 U9628 ( .A1(n7955), .A2(n7964), .ZN(n7956) );
  AOI21_X1 U9629 ( .B1(n7958), .B2(n7957), .A(n7956), .ZN(n7968) );
  NAND2_X1 U9630 ( .A1(n7960), .A2(n7959), .ZN(n7961) );
  AOI21_X1 U9631 ( .B1(n7963), .B2(n7962), .A(n7961), .ZN(n7966) );
  OAI21_X1 U9632 ( .B1(n7966), .B2(n7965), .A(n7964), .ZN(n7967) );
  MUX2_X1 U9633 ( .A(n7968), .B(n7967), .S(n8085), .Z(n7970) );
  OAI22_X1 U9634 ( .A1(n7970), .A2(n8434), .B1(n8085), .B2(n7969), .ZN(n7984)
         );
  MUX2_X1 U9635 ( .A(n7976), .B(n7971), .S(n8085), .Z(n7973) );
  NAND2_X1 U9636 ( .A1(n7973), .A2(n7972), .ZN(n7979) );
  INV_X1 U9637 ( .A(n7979), .ZN(n7983) );
  INV_X1 U9638 ( .A(n7974), .ZN(n7981) );
  AND2_X1 U9639 ( .A1(n7976), .A2(n7975), .ZN(n7978) );
  OAI211_X1 U9640 ( .C1(n7979), .C2(n7978), .A(n7986), .B(n7977), .ZN(n7980)
         );
  MUX2_X1 U9641 ( .A(n7981), .B(n7980), .S(n8085), .Z(n7982) );
  NAND2_X1 U9642 ( .A1(n7990), .A2(n7985), .ZN(n7988) );
  NAND2_X1 U9643 ( .A1(n7989), .A2(n7986), .ZN(n7987) );
  MUX2_X1 U9644 ( .A(n7988), .B(n7987), .S(n8070), .Z(n7993) );
  MUX2_X1 U9645 ( .A(n7990), .B(n7989), .S(n8085), .Z(n7992) );
  NAND2_X1 U9646 ( .A1(n8509), .A2(n7994), .ZN(n7995) );
  MUX2_X1 U9647 ( .A(n7996), .B(n7995), .S(n8070), .Z(n7998) );
  MUX2_X1 U9648 ( .A(n8000), .B(n7999), .S(n8085), .Z(n8001) );
  OAI211_X1 U9649 ( .C1(n8005), .C2(n8004), .A(n8003), .B(n8002), .ZN(n8010)
         );
  AND2_X1 U9650 ( .A1(n8014), .A2(n8006), .ZN(n8007) );
  MUX2_X1 U9651 ( .A(n8008), .B(n8007), .S(n8085), .Z(n8009) );
  NAND3_X1 U9652 ( .A1(n8010), .A2(n8009), .A3(n8012), .ZN(n8011) );
  NAND2_X1 U9653 ( .A1(n8011), .A2(n8370), .ZN(n8017) );
  INV_X1 U9654 ( .A(n8012), .ZN(n8013) );
  NOR2_X1 U9655 ( .A1(n8017), .A2(n8013), .ZN(n8019) );
  INV_X1 U9656 ( .A(n8014), .ZN(n8016) );
  OAI211_X1 U9657 ( .C1(n8017), .C2(n8016), .A(n8024), .B(n8015), .ZN(n8018)
         );
  NAND3_X1 U9658 ( .A1(n8026), .A2(n8027), .A3(n8022), .ZN(n8020) );
  NAND3_X1 U9659 ( .A1(n8020), .A2(n8030), .A3(n8023), .ZN(n8029) );
  NAND2_X1 U9660 ( .A1(n8022), .A2(n8021), .ZN(n8025) );
  OAI211_X1 U9661 ( .C1(n8026), .C2(n8025), .A(n8024), .B(n8023), .ZN(n8028)
         );
  AND2_X1 U9662 ( .A1(n8034), .A2(n8030), .ZN(n8032) );
  MUX2_X1 U9663 ( .A(n8032), .B(n8031), .S(n8070), .Z(n8033) );
  MUX2_X1 U9664 ( .A(n8035), .B(n8034), .S(n8070), .Z(n8036) );
  AND2_X1 U9665 ( .A1(n8038), .A2(n8037), .ZN(n8039) );
  MUX2_X1 U9666 ( .A(n8040), .B(n8039), .S(n8070), .Z(n8042) );
  INV_X1 U9667 ( .A(n8041), .ZN(n8047) );
  NAND4_X1 U9668 ( .A1(n8043), .A2(n8296), .A3(n8042), .A4(n8047), .ZN(n8053)
         );
  OAI21_X1 U9669 ( .B1(n8045), .B2(n8044), .A(n8046), .ZN(n8051) );
  NAND2_X1 U9670 ( .A1(n8047), .A2(n8046), .ZN(n8048) );
  NAND2_X1 U9671 ( .A1(n8049), .A2(n8048), .ZN(n8050) );
  MUX2_X1 U9672 ( .A(n8051), .B(n8050), .S(n8070), .Z(n8052) );
  NAND3_X1 U9673 ( .A1(n8053), .A2(n4682), .A3(n8052), .ZN(n8060) );
  MUX2_X1 U9674 ( .A(n8055), .B(n8054), .S(n8085), .Z(n8056) );
  MUX2_X1 U9675 ( .A(n8062), .B(n8061), .S(n8070), .Z(n8066) );
  MUX2_X1 U9676 ( .A(n8064), .B(n8063), .S(n8085), .Z(n8065) );
  OAI21_X1 U9677 ( .B1(n8067), .B2(n8066), .A(n8065), .ZN(n8068) );
  NAND2_X1 U9678 ( .A1(n8069), .A2(n8068), .ZN(n8075) );
  MUX2_X1 U9679 ( .A(n8077), .B(n8076), .S(n8070), .Z(n8074) );
  MUX2_X1 U9680 ( .A(n8077), .B(n8076), .S(n8085), .Z(n8078) );
  INV_X1 U9681 ( .A(n8084), .ZN(n8082) );
  NOR2_X1 U9682 ( .A1(n8082), .A2(n8081), .ZN(n8087) );
  NAND2_X1 U9683 ( .A1(n8084), .A2(n8083), .ZN(n8086) );
  NOR2_X1 U9684 ( .A1(n8089), .A2(n8088), .ZN(n8091) );
  XNOR2_X1 U9685 ( .A(n8097), .B(n8096), .ZN(n8104) );
  NOR3_X1 U9686 ( .A1(n8099), .A2(n8098), .A3(n6205), .ZN(n8102) );
  OAI21_X1 U9687 ( .B1(n8103), .B2(n8100), .A(P2_B_REG_SCAN_IN), .ZN(n8101) );
  OAI22_X1 U9688 ( .A1(n8104), .A2(n8103), .B1(n8102), .B2(n8101), .ZN(
        P2_U3296) );
  MUX2_X1 U9689 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8105), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9690 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8106), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9691 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8107), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9692 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8108), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9693 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8109), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9694 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8110), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9695 ( .A(n8111), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8248), .Z(
        P2_U3514) );
  MUX2_X1 U9696 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8112), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9697 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n6087), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9698 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8113), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9699 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8114), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9700 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8115), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9701 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8116), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9702 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8117), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9703 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8410), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9704 ( .A(n8118), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8248), .Z(
        P2_U3505) );
  MUX2_X1 U9705 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8409), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U9706 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8119), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9707 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8120), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9708 ( .A(n8121), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8248), .Z(
        P2_U3501) );
  MUX2_X1 U9709 ( .A(n8122), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8248), .Z(
        P2_U3500) );
  MUX2_X1 U9710 ( .A(n8431), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8248), .Z(
        P2_U3499) );
  MUX2_X1 U9711 ( .A(n8123), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8248), .Z(
        P2_U3498) );
  MUX2_X1 U9712 ( .A(n8432), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8248), .Z(
        P2_U3497) );
  MUX2_X1 U9713 ( .A(n8124), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8248), .Z(
        P2_U3496) );
  MUX2_X1 U9714 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8125), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U9715 ( .A(n5867), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8248), .Z(
        P2_U3494) );
  MUX2_X1 U9716 ( .A(n8126), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8248), .Z(
        P2_U3493) );
  MUX2_X1 U9717 ( .A(n5842), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8248), .Z(
        P2_U3492) );
  MUX2_X1 U9718 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8127), .S(P2_U3893), .Z(
        P2_U3491) );
  INV_X1 U9719 ( .A(n8128), .ZN(n8130) );
  NAND2_X1 U9720 ( .A1(n8130), .A2(n8129), .ZN(n8131) );
  XNOR2_X1 U9721 ( .A(n8132), .B(n8131), .ZN(n8148) );
  AND3_X1 U9722 ( .A1(n8135), .A2(n8134), .A3(n8133), .ZN(n8136) );
  OAI21_X1 U9723 ( .B1(n8137), .B2(n8136), .A(n9816), .ZN(n8145) );
  AOI21_X1 U9724 ( .B1(n8140), .B2(n8139), .A(n8138), .ZN(n8141) );
  NOR2_X1 U9725 ( .A1(n9825), .A2(n8141), .ZN(n8142) );
  AOI211_X1 U9726 ( .C1(n9840), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n8143), .B(
        n8142), .ZN(n8144) );
  OAI211_X1 U9727 ( .C1(n8246), .C2(n8146), .A(n8145), .B(n8144), .ZN(n8147)
         );
  AOI21_X1 U9728 ( .B1(n8148), .B2(n9838), .A(n8147), .ZN(n8149) );
  INV_X1 U9729 ( .A(n8149), .ZN(P2_U3194) );
  AOI21_X1 U9730 ( .B1(n8506), .B2(n8151), .A(n8150), .ZN(n8166) );
  OAI21_X1 U9731 ( .B1(n8255), .B2(n8153), .A(n8152), .ZN(n8158) );
  AOI21_X1 U9732 ( .B1(n8155), .B2(n6351), .A(n8154), .ZN(n8156) );
  NOR2_X1 U9733 ( .A1(n8156), .A2(n9832), .ZN(n8157) );
  AOI211_X1 U9734 ( .C1(n9830), .C2(n8159), .A(n8158), .B(n8157), .ZN(n8165)
         );
  OAI21_X1 U9735 ( .B1(n8162), .B2(n8161), .A(n8160), .ZN(n8163) );
  NAND2_X1 U9736 ( .A1(n8163), .A2(n9838), .ZN(n8164) );
  OAI211_X1 U9737 ( .C1(n8166), .C2(n9825), .A(n8165), .B(n8164), .ZN(P2_U3195) );
  AOI21_X1 U9738 ( .B1(n4409), .B2(n8168), .A(n8167), .ZN(n8183) );
  OAI21_X1 U9739 ( .B1(n8171), .B2(n8170), .A(n8169), .ZN(n8172) );
  NAND2_X1 U9740 ( .A1(n8172), .A2(n9838), .ZN(n8174) );
  OAI211_X1 U9741 ( .C1(n8255), .C2(n8175), .A(n8174), .B(n8173), .ZN(n8180)
         );
  AOI21_X1 U9742 ( .B1(n4394), .B2(n8177), .A(n8176), .ZN(n8178) );
  NOR2_X1 U9743 ( .A1(n8178), .A2(n9832), .ZN(n8179) );
  AOI211_X1 U9744 ( .C1(n9830), .C2(n8181), .A(n8180), .B(n8179), .ZN(n8182)
         );
  OAI21_X1 U9745 ( .B1(n8183), .B2(n9825), .A(n8182), .ZN(P2_U3196) );
  AOI21_X1 U9746 ( .B1(n8498), .B2(n8185), .A(n8184), .ZN(n8201) );
  OAI21_X1 U9747 ( .B1(n8188), .B2(n8187), .A(n8186), .ZN(n8197) );
  NOR2_X1 U9748 ( .A1(n8255), .A2(n8189), .ZN(n8196) );
  AOI21_X1 U9749 ( .B1(n8192), .B2(n8191), .A(n8190), .ZN(n8194) );
  OAI21_X1 U9750 ( .B1(n9832), .B2(n8194), .A(n8193), .ZN(n8195) );
  AOI211_X1 U9751 ( .C1(n9838), .C2(n8197), .A(n8196), .B(n8195), .ZN(n8200)
         );
  NAND2_X1 U9752 ( .A1(n9830), .A2(n8198), .ZN(n8199) );
  OAI211_X1 U9753 ( .C1(n8201), .C2(n9825), .A(n8200), .B(n8199), .ZN(P2_U3197) );
  AOI21_X1 U9754 ( .B1(n4397), .B2(n8203), .A(n8202), .ZN(n8218) );
  OAI21_X1 U9755 ( .B1(n8206), .B2(n8205), .A(n8204), .ZN(n8207) );
  NAND2_X1 U9756 ( .A1(n8207), .A2(n9838), .ZN(n8209) );
  OAI211_X1 U9757 ( .C1(n8255), .C2(n8210), .A(n8209), .B(n8208), .ZN(n8215)
         );
  AOI21_X1 U9758 ( .B1(n4400), .B2(n8212), .A(n8211), .ZN(n8213) );
  NOR2_X1 U9759 ( .A1(n8213), .A2(n9832), .ZN(n8214) );
  AOI211_X1 U9760 ( .C1(n9830), .C2(n8216), .A(n8215), .B(n8214), .ZN(n8217)
         );
  OAI21_X1 U9761 ( .B1(n8218), .B2(n9825), .A(n8217), .ZN(P2_U3198) );
  AOI21_X1 U9762 ( .B1(n8221), .B2(n8220), .A(n8219), .ZN(n8236) );
  OAI21_X1 U9763 ( .B1(n8224), .B2(n8223), .A(n8222), .ZN(n8232) );
  NOR2_X1 U9764 ( .A1(n8255), .A2(n8225), .ZN(n8231) );
  AOI21_X1 U9765 ( .B1(n8227), .B2(n8380), .A(n8226), .ZN(n8229) );
  OAI21_X1 U9766 ( .B1(n9832), .B2(n8229), .A(n8228), .ZN(n8230) );
  AOI211_X1 U9767 ( .C1(n9838), .C2(n8232), .A(n8231), .B(n8230), .ZN(n8235)
         );
  NAND2_X1 U9768 ( .A1(n9830), .A2(n8233), .ZN(n8234) );
  OAI211_X1 U9769 ( .C1(n8236), .C2(n9825), .A(n8235), .B(n8234), .ZN(P2_U3199) );
  NAND2_X1 U9770 ( .A1(n8241), .A2(n8240), .ZN(n8242) );
  NAND2_X1 U9771 ( .A1(n8243), .A2(n8242), .ZN(n8258) );
  OAI21_X1 U9772 ( .B1(n8248), .B2(n8247), .A(n8246), .ZN(n8253) );
  NOR2_X1 U9773 ( .A1(n8250), .A2(n8249), .ZN(n8252) );
  MUX2_X1 U9774 ( .A(n8253), .B(n8252), .S(n8251), .Z(n8257) );
  OAI21_X1 U9775 ( .B1(n8255), .B2(n9928), .A(n8254), .ZN(n8256) );
  NAND2_X1 U9776 ( .A1(n8513), .A2(n8382), .ZN(n8261) );
  OAI211_X1 U9777 ( .C1(n8398), .C2(n8262), .A(n8261), .B(n8260), .ZN(P2_U3202) );
  INV_X1 U9778 ( .A(n8263), .ZN(n8270) );
  AOI22_X1 U9779 ( .A1(n8264), .A2(n8353), .B1(n8441), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8265) );
  OAI21_X1 U9780 ( .B1(n8266), .B2(n8429), .A(n8265), .ZN(n8267) );
  AOI21_X1 U9781 ( .B1(n8268), .B2(n8419), .A(n8267), .ZN(n8269) );
  OAI21_X1 U9782 ( .B1(n8270), .B2(n8418), .A(n8269), .ZN(P2_U3206) );
  XNOR2_X1 U9783 ( .A(n8271), .B(n8274), .ZN(n8272) );
  OAI222_X1 U9784 ( .A1(n8392), .A2(n8273), .B1(n8390), .B2(n8293), .C1(n9845), 
        .C2(n8272), .ZN(n8452) );
  INV_X1 U9785 ( .A(n8452), .ZN(n8280) );
  XOR2_X1 U9786 ( .A(n8275), .B(n8274), .Z(n8453) );
  AOI22_X1 U9787 ( .A1(n8276), .A2(n8353), .B1(n8441), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8277) );
  OAI21_X1 U9788 ( .B1(n8524), .B2(n8429), .A(n8277), .ZN(n8278) );
  AOI21_X1 U9789 ( .B1(n8453), .B2(n8419), .A(n8278), .ZN(n8279) );
  OAI21_X1 U9790 ( .B1(n8280), .B2(n8418), .A(n8279), .ZN(P2_U3207) );
  NOR2_X1 U9791 ( .A1(n8528), .A2(n8413), .ZN(n8284) );
  XNOR2_X1 U9792 ( .A(n8281), .B(n4682), .ZN(n8282) );
  OAI222_X1 U9793 ( .A1(n8392), .A2(n8283), .B1(n8390), .B2(n8302), .C1(n9845), 
        .C2(n8282), .ZN(n8456) );
  AOI211_X1 U9794 ( .C1(n8353), .C2(n8285), .A(n8284), .B(n8456), .ZN(n8289)
         );
  XNOR2_X1 U9795 ( .A(n8287), .B(n8286), .ZN(n8457) );
  AOI22_X1 U9796 ( .A1(n8457), .A2(n8419), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8418), .ZN(n8288) );
  OAI21_X1 U9797 ( .B1(n8289), .B2(n8418), .A(n8288), .ZN(P2_U3208) );
  NOR2_X1 U9798 ( .A1(n8532), .A2(n8413), .ZN(n8294) );
  XNOR2_X1 U9799 ( .A(n8291), .B(n8290), .ZN(n8292) );
  OAI222_X1 U9800 ( .A1(n8390), .A2(n8312), .B1(n8392), .B2(n8293), .C1(n8292), 
        .C2(n9845), .ZN(n8460) );
  AOI211_X1 U9801 ( .C1(n8353), .C2(n8295), .A(n8294), .B(n8460), .ZN(n8299)
         );
  XNOR2_X1 U9802 ( .A(n8297), .B(n8296), .ZN(n8461) );
  AOI22_X1 U9803 ( .A1(n8461), .A2(n8419), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8418), .ZN(n8298) );
  OAI21_X1 U9804 ( .B1(n8299), .B2(n8418), .A(n8298), .ZN(P2_U3209) );
  XOR2_X1 U9805 ( .A(n8303), .B(n8300), .Z(n8301) );
  OAI222_X1 U9806 ( .A1(n8390), .A2(n8322), .B1(n8392), .B2(n8302), .C1(n9845), 
        .C2(n8301), .ZN(n8464) );
  INV_X1 U9807 ( .A(n8464), .ZN(n8309) );
  XNOR2_X1 U9808 ( .A(n8304), .B(n8303), .ZN(n8465) );
  AOI22_X1 U9809 ( .A1(n8441), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8353), .B2(
        n8305), .ZN(n8306) );
  OAI21_X1 U9810 ( .B1(n8536), .B2(n8429), .A(n8306), .ZN(n8307) );
  AOI21_X1 U9811 ( .B1(n8465), .B2(n8419), .A(n8307), .ZN(n8308) );
  OAI21_X1 U9812 ( .B1(n8309), .B2(n8418), .A(n8308), .ZN(P2_U3210) );
  XOR2_X1 U9813 ( .A(n8310), .B(n8313), .Z(n8311) );
  OAI222_X1 U9814 ( .A1(n8390), .A2(n8336), .B1(n8392), .B2(n8312), .C1(n9845), 
        .C2(n8311), .ZN(n8468) );
  INV_X1 U9815 ( .A(n8468), .ZN(n8319) );
  XOR2_X1 U9816 ( .A(n8314), .B(n8313), .Z(n8469) );
  AOI22_X1 U9817 ( .A1(n8441), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8353), .B2(
        n8315), .ZN(n8316) );
  OAI21_X1 U9818 ( .B1(n8540), .B2(n8429), .A(n8316), .ZN(n8317) );
  AOI21_X1 U9819 ( .B1(n8469), .B2(n8419), .A(n8317), .ZN(n8318) );
  OAI21_X1 U9820 ( .B1(n8319), .B2(n8441), .A(n8318), .ZN(P2_U3211) );
  XNOR2_X1 U9821 ( .A(n8320), .B(n8325), .ZN(n8321) );
  OAI222_X1 U9822 ( .A1(n8390), .A2(n8346), .B1(n8392), .B2(n8322), .C1(n9845), 
        .C2(n8321), .ZN(n8472) );
  INV_X1 U9823 ( .A(n8472), .ZN(n8331) );
  NAND2_X1 U9824 ( .A1(n8324), .A2(n8323), .ZN(n8326) );
  XNOR2_X1 U9825 ( .A(n8326), .B(n8325), .ZN(n8473) );
  AOI22_X1 U9826 ( .A1(n8441), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8353), .B2(
        n8327), .ZN(n8328) );
  OAI21_X1 U9827 ( .B1(n8544), .B2(n8429), .A(n8328), .ZN(n8329) );
  AOI21_X1 U9828 ( .B1(n8473), .B2(n8419), .A(n8329), .ZN(n8330) );
  OAI21_X1 U9829 ( .B1(n8331), .B2(n8441), .A(n8330), .ZN(P2_U3212) );
  OAI21_X1 U9830 ( .B1(n8333), .B2(n8337), .A(n8332), .ZN(n8334) );
  INV_X1 U9831 ( .A(n8334), .ZN(n8335) );
  OAI222_X1 U9832 ( .A1(n8392), .A2(n8336), .B1(n8390), .B2(n8360), .C1(n9845), 
        .C2(n8335), .ZN(n8476) );
  INV_X1 U9833 ( .A(n8476), .ZN(n8343) );
  XOR2_X1 U9834 ( .A(n8338), .B(n8337), .Z(n8477) );
  AOI22_X1 U9835 ( .A1(n8441), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8353), .B2(
        n8339), .ZN(n8340) );
  OAI21_X1 U9836 ( .B1(n8548), .B2(n8429), .A(n8340), .ZN(n8341) );
  AOI21_X1 U9837 ( .B1(n8477), .B2(n8419), .A(n8341), .ZN(n8342) );
  OAI21_X1 U9838 ( .B1(n8343), .B2(n8441), .A(n8342), .ZN(P2_U3213) );
  AOI211_X1 U9839 ( .C1(n8349), .C2(n8345), .A(n9845), .B(n8344), .ZN(n8348)
         );
  OAI22_X1 U9840 ( .A1(n8346), .A2(n8392), .B1(n8375), .B2(n8390), .ZN(n8347)
         );
  OR2_X1 U9841 ( .A1(n8348), .A2(n8347), .ZN(n8480) );
  INV_X1 U9842 ( .A(n8480), .ZN(n8357) );
  XOR2_X1 U9843 ( .A(n8350), .B(n8349), .Z(n8481) );
  INV_X1 U9844 ( .A(n8351), .ZN(n8552) );
  AOI22_X1 U9845 ( .A1(n8441), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8353), .B2(
        n8352), .ZN(n8354) );
  OAI21_X1 U9846 ( .B1(n8552), .B2(n8429), .A(n8354), .ZN(n8355) );
  AOI21_X1 U9847 ( .B1(n8481), .B2(n8419), .A(n8355), .ZN(n8356) );
  OAI21_X1 U9848 ( .B1(n8357), .B2(n8441), .A(n8356), .ZN(P2_U3214) );
  XNOR2_X1 U9849 ( .A(n8358), .B(n8362), .ZN(n8359) );
  OAI222_X1 U9850 ( .A1(n8390), .A2(n8391), .B1(n8392), .B2(n8360), .C1(n8359), 
        .C2(n9845), .ZN(n8484) );
  INV_X1 U9851 ( .A(n8484), .ZN(n8368) );
  AOI21_X1 U9852 ( .B1(n8362), .B2(n8361), .A(n4411), .ZN(n8485) );
  NOR2_X1 U9853 ( .A1(n8556), .A2(n8429), .ZN(n8366) );
  OAI22_X1 U9854 ( .A1(n8398), .A2(n8364), .B1(n8363), .B2(n8427), .ZN(n8365)
         );
  AOI211_X1 U9855 ( .C1(n8485), .C2(n8419), .A(n8366), .B(n8365), .ZN(n8367)
         );
  OAI21_X1 U9856 ( .B1(n8368), .B2(n8441), .A(n8367), .ZN(P2_U3215) );
  XNOR2_X1 U9857 ( .A(n8369), .B(n8370), .ZN(n8489) );
  XNOR2_X1 U9858 ( .A(n8372), .B(n8371), .ZN(n8373) );
  NAND2_X1 U9859 ( .A1(n8373), .A2(n8436), .ZN(n8378) );
  OAI22_X1 U9860 ( .A1(n8375), .A2(n8392), .B1(n8374), .B2(n8390), .ZN(n8376)
         );
  INV_X1 U9861 ( .A(n8376), .ZN(n8377) );
  NAND2_X1 U9862 ( .A1(n8378), .A2(n8377), .ZN(n8491) );
  NAND2_X1 U9863 ( .A1(n8491), .A2(n8398), .ZN(n8385) );
  OAI22_X1 U9864 ( .A1(n8398), .A2(n8380), .B1(n8379), .B2(n8427), .ZN(n8381)
         );
  AOI21_X1 U9865 ( .B1(n8383), .B2(n8382), .A(n8381), .ZN(n8384) );
  OAI211_X1 U9866 ( .C1(n8489), .C2(n8386), .A(n8385), .B(n8384), .ZN(P2_U3216) );
  XNOR2_X1 U9867 ( .A(n8387), .B(n8393), .ZN(n8388) );
  OAI222_X1 U9868 ( .A1(n8392), .A2(n8391), .B1(n8390), .B2(n8389), .C1(n8388), 
        .C2(n9845), .ZN(n8492) );
  INV_X1 U9869 ( .A(n8492), .ZN(n8402) );
  XNOR2_X1 U9870 ( .A(n8394), .B(n8393), .ZN(n8493) );
  INV_X1 U9871 ( .A(n8395), .ZN(n8561) );
  NOR2_X1 U9872 ( .A1(n8561), .A2(n8429), .ZN(n8400) );
  OAI22_X1 U9873 ( .A1(n8398), .A2(n8397), .B1(n8396), .B2(n8427), .ZN(n8399)
         );
  AOI211_X1 U9874 ( .C1(n8493), .C2(n8419), .A(n8400), .B(n8399), .ZN(n8401)
         );
  OAI21_X1 U9875 ( .B1(n8402), .B2(n8441), .A(n8401), .ZN(P2_U3217) );
  NAND2_X1 U9876 ( .A1(n8404), .A2(n8403), .ZN(n8406) );
  NAND2_X1 U9877 ( .A1(n8406), .A2(n8405), .ZN(n8408) );
  XNOR2_X1 U9878 ( .A(n8408), .B(n8407), .ZN(n8411) );
  AOI222_X1 U9879 ( .A1(n8436), .A2(n8411), .B1(n8410), .B2(n8430), .C1(n8409), 
        .C2(n8433), .ZN(n8503) );
  INV_X1 U9880 ( .A(n8503), .ZN(n8416) );
  OAI22_X1 U9881 ( .A1(n8414), .A2(n8413), .B1(n8412), .B2(n8427), .ZN(n8415)
         );
  OAI21_X1 U9882 ( .B1(n8416), .B2(n8415), .A(n8398), .ZN(n8421) );
  OAI21_X1 U9883 ( .B1(n4415), .B2(n6194), .A(n8417), .ZN(n8501) );
  AOI22_X1 U9884 ( .A1(n8501), .A2(n8419), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8418), .ZN(n8420) );
  NAND2_X1 U9885 ( .A1(n8421), .A2(n8420), .ZN(P2_U3219) );
  NAND2_X1 U9886 ( .A1(n8423), .A2(n8422), .ZN(n8424) );
  NAND2_X1 U9887 ( .A1(n8424), .A2(n8434), .ZN(n8425) );
  NAND2_X1 U9888 ( .A1(n8426), .A2(n8425), .ZN(n9883) );
  INV_X1 U9889 ( .A(n9883), .ZN(n8445) );
  OAI22_X1 U9890 ( .A1(n8429), .A2(n9882), .B1(n8428), .B2(n8427), .ZN(n8443)
         );
  AOI22_X1 U9891 ( .A1(n8433), .A2(n8432), .B1(n8431), .B2(n8430), .ZN(n8439)
         );
  XNOR2_X1 U9892 ( .A(n8435), .B(n8434), .ZN(n8437) );
  NAND2_X1 U9893 ( .A1(n8437), .A2(n8436), .ZN(n8438) );
  OAI211_X1 U9894 ( .C1(n9883), .C2(n8440), .A(n8439), .B(n8438), .ZN(n9885)
         );
  MUX2_X1 U9895 ( .A(n9885), .B(P2_REG2_REG_7__SCAN_IN), .S(n8441), .Z(n8442)
         );
  AOI211_X1 U9896 ( .C1(n8445), .C2(n8444), .A(n8443), .B(n8442), .ZN(n8446)
         );
  INV_X1 U9897 ( .A(n8446), .ZN(P2_U3226) );
  INV_X1 U9898 ( .A(n8508), .ZN(n8448) );
  NAND2_X1 U9899 ( .A1(n8513), .A2(n8448), .ZN(n8447) );
  NAND2_X1 U9900 ( .A1(n8514), .A2(n9920), .ZN(n8449) );
  OAI211_X1 U9901 ( .C1(n9920), .C2(n7026), .A(n8447), .B(n8449), .ZN(P2_U3490) );
  INV_X1 U9902 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U9903 ( .A1(n8518), .A2(n8448), .ZN(n8450) );
  OAI211_X1 U9904 ( .C1(n9920), .C2(n8451), .A(n8450), .B(n8449), .ZN(P2_U3489) );
  INV_X1 U9905 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8454) );
  AOI21_X1 U9906 ( .B1(n8453), .B2(n6266), .A(n8452), .ZN(n8521) );
  MUX2_X1 U9907 ( .A(n8454), .B(n8521), .S(n9920), .Z(n8455) );
  OAI21_X1 U9908 ( .B1(n8524), .B2(n8508), .A(n8455), .ZN(P2_U3485) );
  INV_X1 U9909 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8458) );
  AOI21_X1 U9910 ( .B1(n6266), .B2(n8457), .A(n8456), .ZN(n8525) );
  MUX2_X1 U9911 ( .A(n8458), .B(n8525), .S(n9920), .Z(n8459) );
  OAI21_X1 U9912 ( .B1(n8528), .B2(n8508), .A(n8459), .ZN(P2_U3484) );
  INV_X1 U9913 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8462) );
  AOI21_X1 U9914 ( .B1(n8461), .B2(n6266), .A(n8460), .ZN(n8529) );
  MUX2_X1 U9915 ( .A(n8462), .B(n8529), .S(n9920), .Z(n8463) );
  OAI21_X1 U9916 ( .B1(n8532), .B2(n8508), .A(n8463), .ZN(P2_U3483) );
  INV_X1 U9917 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8466) );
  AOI21_X1 U9918 ( .B1(n6266), .B2(n8465), .A(n8464), .ZN(n8533) );
  MUX2_X1 U9919 ( .A(n8466), .B(n8533), .S(n9920), .Z(n8467) );
  OAI21_X1 U9920 ( .B1(n8536), .B2(n8508), .A(n8467), .ZN(P2_U3482) );
  INV_X1 U9921 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8470) );
  AOI21_X1 U9922 ( .B1(n6266), .B2(n8469), .A(n8468), .ZN(n8537) );
  MUX2_X1 U9923 ( .A(n8470), .B(n8537), .S(n9920), .Z(n8471) );
  OAI21_X1 U9924 ( .B1(n8540), .B2(n8508), .A(n8471), .ZN(P2_U3481) );
  INV_X1 U9925 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8474) );
  AOI21_X1 U9926 ( .B1(n8473), .B2(n6266), .A(n8472), .ZN(n8541) );
  MUX2_X1 U9927 ( .A(n8474), .B(n8541), .S(n9920), .Z(n8475) );
  OAI21_X1 U9928 ( .B1(n8544), .B2(n8508), .A(n8475), .ZN(P2_U3480) );
  INV_X1 U9929 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8478) );
  AOI21_X1 U9930 ( .B1(n8477), .B2(n6266), .A(n8476), .ZN(n8545) );
  MUX2_X1 U9931 ( .A(n8478), .B(n8545), .S(n9920), .Z(n8479) );
  OAI21_X1 U9932 ( .B1(n8548), .B2(n8508), .A(n8479), .ZN(P2_U3479) );
  AOI21_X1 U9933 ( .B1(n6266), .B2(n8481), .A(n8480), .ZN(n8549) );
  MUX2_X1 U9934 ( .A(n8482), .B(n8549), .S(n9920), .Z(n8483) );
  OAI21_X1 U9935 ( .B1(n8552), .B2(n8508), .A(n8483), .ZN(P2_U3478) );
  INV_X1 U9936 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8486) );
  AOI21_X1 U9937 ( .B1(n8485), .B2(n6266), .A(n8484), .ZN(n8553) );
  MUX2_X1 U9938 ( .A(n8486), .B(n8553), .S(n9920), .Z(n8487) );
  OAI21_X1 U9939 ( .B1(n8556), .B2(n8508), .A(n8487), .ZN(P2_U3477) );
  OAI22_X1 U9940 ( .A1(n8489), .A2(n9877), .B1(n8488), .B2(n9894), .ZN(n8490)
         );
  MUX2_X1 U9941 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8557), .S(n9920), .Z(
        P2_U3476) );
  AOI21_X1 U9942 ( .B1(n6266), .B2(n8493), .A(n8492), .ZN(n8558) );
  MUX2_X1 U9943 ( .A(n8494), .B(n8558), .S(n9920), .Z(n8495) );
  OAI21_X1 U9944 ( .B1(n8561), .B2(n8508), .A(n8495), .ZN(P2_U3475) );
  AOI21_X1 U9945 ( .B1(n8497), .B2(n6266), .A(n8496), .ZN(n8562) );
  MUX2_X1 U9946 ( .A(n8498), .B(n8562), .S(n9920), .Z(n8499) );
  OAI21_X1 U9947 ( .B1(n8565), .B2(n8508), .A(n8499), .ZN(P2_U3474) );
  AOI22_X1 U9948 ( .A1(n8501), .A2(n6266), .B1(n9900), .B2(n8500), .ZN(n8502)
         );
  NAND2_X1 U9949 ( .A1(n8503), .A2(n8502), .ZN(n8566) );
  MUX2_X1 U9950 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8566), .S(n9920), .Z(
        P2_U3473) );
  AOI21_X1 U9951 ( .B1(n8505), .B2(n6266), .A(n8504), .ZN(n8567) );
  MUX2_X1 U9952 ( .A(n8506), .B(n8567), .S(n9920), .Z(n8507) );
  OAI21_X1 U9953 ( .B1(n8571), .B2(n8508), .A(n8507), .ZN(P2_U3472) );
  AOI22_X1 U9954 ( .A1(n8510), .A2(n6266), .B1(n9900), .B2(n8509), .ZN(n8511)
         );
  NAND2_X1 U9955 ( .A1(n8512), .A2(n8511), .ZN(n8572) );
  MUX2_X1 U9956 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8572), .S(n9920), .Z(
        P2_U3471) );
  INV_X1 U9957 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8516) );
  INV_X1 U9958 ( .A(n8570), .ZN(n8517) );
  NAND2_X1 U9959 ( .A1(n8513), .A2(n8517), .ZN(n8515) );
  NAND2_X1 U9960 ( .A1(n8514), .A2(n9905), .ZN(n8519) );
  OAI211_X1 U9961 ( .C1(n8516), .C2(n9905), .A(n8515), .B(n8519), .ZN(P2_U3458) );
  NAND2_X1 U9962 ( .A1(n8518), .A2(n8517), .ZN(n8520) );
  OAI211_X1 U9963 ( .C1(n6210), .C2(n9905), .A(n8520), .B(n8519), .ZN(P2_U3457) );
  MUX2_X1 U9964 ( .A(n8522), .B(n8521), .S(n9905), .Z(n8523) );
  OAI21_X1 U9965 ( .B1(n8524), .B2(n8570), .A(n8523), .ZN(P2_U3453) );
  MUX2_X1 U9966 ( .A(n8526), .B(n8525), .S(n9905), .Z(n8527) );
  OAI21_X1 U9967 ( .B1(n8528), .B2(n8570), .A(n8527), .ZN(P2_U3452) );
  INV_X1 U9968 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8530) );
  MUX2_X1 U9969 ( .A(n8530), .B(n8529), .S(n9905), .Z(n8531) );
  OAI21_X1 U9970 ( .B1(n8532), .B2(n8570), .A(n8531), .ZN(P2_U3451) );
  MUX2_X1 U9971 ( .A(n8534), .B(n8533), .S(n9905), .Z(n8535) );
  OAI21_X1 U9972 ( .B1(n8536), .B2(n8570), .A(n8535), .ZN(P2_U3450) );
  INV_X1 U9973 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8538) );
  MUX2_X1 U9974 ( .A(n8538), .B(n8537), .S(n9905), .Z(n8539) );
  OAI21_X1 U9975 ( .B1(n8540), .B2(n8570), .A(n8539), .ZN(P2_U3449) );
  INV_X1 U9976 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8542) );
  MUX2_X1 U9977 ( .A(n8542), .B(n8541), .S(n9905), .Z(n8543) );
  OAI21_X1 U9978 ( .B1(n8544), .B2(n8570), .A(n8543), .ZN(P2_U3448) );
  INV_X1 U9979 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8546) );
  MUX2_X1 U9980 ( .A(n8546), .B(n8545), .S(n9905), .Z(n8547) );
  OAI21_X1 U9981 ( .B1(n8548), .B2(n8570), .A(n8547), .ZN(P2_U3447) );
  MUX2_X1 U9982 ( .A(n8550), .B(n8549), .S(n9905), .Z(n8551) );
  OAI21_X1 U9983 ( .B1(n8552), .B2(n8570), .A(n8551), .ZN(P2_U3446) );
  MUX2_X1 U9984 ( .A(n8554), .B(n8553), .S(n9905), .Z(n8555) );
  OAI21_X1 U9985 ( .B1(n8556), .B2(n8570), .A(n8555), .ZN(P2_U3444) );
  MUX2_X1 U9986 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8557), .S(n9905), .Z(
        P2_U3441) );
  INV_X1 U9987 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8559) );
  MUX2_X1 U9988 ( .A(n8559), .B(n8558), .S(n9905), .Z(n8560) );
  OAI21_X1 U9989 ( .B1(n8561), .B2(n8570), .A(n8560), .ZN(P2_U3438) );
  INV_X1 U9990 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8563) );
  MUX2_X1 U9991 ( .A(n8563), .B(n8562), .S(n9905), .Z(n8564) );
  OAI21_X1 U9992 ( .B1(n8565), .B2(n8570), .A(n8564), .ZN(P2_U3435) );
  MUX2_X1 U9993 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8566), .S(n9905), .Z(
        P2_U3432) );
  INV_X1 U9994 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8568) );
  MUX2_X1 U9995 ( .A(n8568), .B(n8567), .S(n9905), .Z(n8569) );
  OAI21_X1 U9996 ( .B1(n8571), .B2(n8570), .A(n8569), .ZN(P2_U3429) );
  MUX2_X1 U9997 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n8572), .S(n9905), .Z(
        P2_U3426) );
  MUX2_X1 U9998 ( .A(P2_D_REG_1__SCAN_IN), .B(n8574), .S(n8573), .Z(P2_U3377)
         );
  NAND3_X1 U9999 ( .A1(n8576), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8579) );
  OAI22_X1 U10000 ( .A1(n8575), .A2(n8579), .B1(n8578), .B2(n8577), .ZN(n8580)
         );
  AOI21_X1 U10001 ( .B1(n9569), .B2(n8581), .A(n8580), .ZN(n8582) );
  INV_X1 U10002 ( .A(n8582), .ZN(P2_U3264) );
  INV_X1 U10003 ( .A(n8584), .ZN(n8589) );
  INV_X1 U10004 ( .A(n8585), .ZN(n8587) );
  NOR2_X1 U10005 ( .A1(n8587), .A2(n8586), .ZN(n8658) );
  AOI21_X1 U10006 ( .B1(n8587), .B2(n8586), .A(n8658), .ZN(n8588) );
  NAND2_X1 U10007 ( .A1(n8588), .A2(n8589), .ZN(n8660) );
  OAI21_X1 U10008 ( .B1(n8589), .B2(n8588), .A(n8660), .ZN(n8590) );
  NAND2_X1 U10009 ( .A1(n8590), .A2(n8748), .ZN(n8595) );
  NAND2_X1 U10010 ( .A1(n8757), .A2(n9029), .ZN(n8591) );
  NAND2_X1 U10011 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9660) );
  OAI211_X1 U10012 ( .C1(n8759), .C2(n9507), .A(n8591), .B(n9660), .ZN(n8592)
         );
  AOI21_X1 U10013 ( .B1(n8593), .B2(n8763), .A(n8592), .ZN(n8594) );
  OAI211_X1 U10014 ( .C1(n8596), .C2(n8760), .A(n8595), .B(n8594), .ZN(
        P1_U3215) );
  INV_X1 U10015 ( .A(n8682), .ZN(n8599) );
  NOR3_X1 U10016 ( .A1(n8709), .A2(n8713), .A3(n8597), .ZN(n8598) );
  OAI21_X1 U10017 ( .B1(n8599), .B2(n8598), .A(n8748), .ZN(n8603) );
  INV_X1 U10018 ( .A(n9438), .ZN(n9027) );
  AOI22_X1 U10019 ( .A1(n8726), .A2(n9027), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n8600) );
  OAI21_X1 U10020 ( .B1(n9439), .B2(n8728), .A(n8600), .ZN(n8601) );
  AOI21_X1 U10021 ( .B1(n9268), .B2(n8763), .A(n8601), .ZN(n8602) );
  OAI211_X1 U10022 ( .C1(n9138), .C2(n8760), .A(n8603), .B(n8602), .ZN(
        P1_U3216) );
  OAI21_X1 U10023 ( .B1(n8605), .B2(n4417), .A(n8604), .ZN(n8612) );
  NOR2_X1 U10024 ( .A1(n8760), .A2(n8606), .ZN(n8611) );
  NAND2_X1 U10025 ( .A1(n8763), .A2(n4919), .ZN(n8609) );
  NAND2_X1 U10026 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9584) );
  INV_X1 U10027 ( .A(n9584), .ZN(n8607) );
  AOI21_X1 U10028 ( .B1(n8757), .B2(n9033), .A(n8607), .ZN(n8608) );
  OAI211_X1 U10029 ( .C1(n8643), .C2(n8759), .A(n8609), .B(n8608), .ZN(n8610)
         );
  AOI211_X1 U10030 ( .C1(n8612), .C2(n8748), .A(n8611), .B(n8610), .ZN(n8613)
         );
  INV_X1 U10031 ( .A(n8613), .ZN(P1_U3217) );
  INV_X1 U10032 ( .A(n8615), .ZN(n8617) );
  XOR2_X1 U10033 ( .A(n8616), .B(n8615), .Z(n8736) );
  NOR2_X1 U10034 ( .A1(n8736), .A2(n8735), .ZN(n8734) );
  AOI21_X1 U10035 ( .B1(n8617), .B2(n8616), .A(n8734), .ZN(n8621) );
  XNOR2_X1 U10036 ( .A(n8619), .B(n8618), .ZN(n8620) );
  XNOR2_X1 U10037 ( .A(n8621), .B(n8620), .ZN(n8626) );
  INV_X1 U10038 ( .A(n9466), .ZN(n9328) );
  NAND2_X1 U10039 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9110) );
  OAI21_X1 U10040 ( .B1(n8759), .B2(n9328), .A(n9110), .ZN(n8622) );
  AOI21_X1 U10041 ( .B1(n8757), .B2(n9465), .A(n8622), .ZN(n8623) );
  OAI21_X1 U10042 ( .B1(n8739), .B2(n9325), .A(n8623), .ZN(n8624) );
  AOI21_X1 U10043 ( .B1(n9324), .B2(n8741), .A(n8624), .ZN(n8625) );
  OAI21_X1 U10044 ( .B1(n8626), .B2(n8766), .A(n8625), .ZN(P1_U3219) );
  XOR2_X1 U10045 ( .A(n8628), .B(n8627), .Z(n8633) );
  INV_X1 U10046 ( .A(n9439), .ZN(n9299) );
  AOI22_X1 U10047 ( .A1(n8726), .A2(n9299), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8630) );
  NAND2_X1 U10048 ( .A1(n8763), .A2(n9293), .ZN(n8629) );
  OAI211_X1 U10049 ( .C1(n9328), .C2(n8728), .A(n8630), .B(n8629), .ZN(n8631)
         );
  AOI21_X1 U10050 ( .B1(n9451), .B2(n8741), .A(n8631), .ZN(n8632) );
  OAI21_X1 U10051 ( .B1(n8633), .B2(n8766), .A(n8632), .ZN(P1_U3223) );
  INV_X1 U10052 ( .A(n8634), .ZN(n8723) );
  INV_X1 U10053 ( .A(n8635), .ZN(n8637) );
  NOR3_X1 U10054 ( .A1(n8723), .A2(n8637), .A3(n8636), .ZN(n8640) );
  INV_X1 U10055 ( .A(n8638), .ZN(n8639) );
  OAI21_X1 U10056 ( .B1(n8640), .B2(n8639), .A(n8748), .ZN(n8647) );
  AOI21_X1 U10057 ( .B1(n8726), .B2(n9029), .A(n8641), .ZN(n8642) );
  OAI21_X1 U10058 ( .B1(n8643), .B2(n8728), .A(n8642), .ZN(n8644) );
  AOI21_X1 U10059 ( .B1(n8645), .B2(n8763), .A(n8644), .ZN(n8646) );
  OAI211_X1 U10060 ( .C1(n8648), .C2(n8760), .A(n8647), .B(n8646), .ZN(
        P1_U3224) );
  AOI21_X1 U10061 ( .B1(n8650), .B2(n8649), .A(n4343), .ZN(n8655) );
  AOI22_X1 U10062 ( .A1(n8726), .A2(n9242), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8652) );
  NAND2_X1 U10063 ( .A1(n8763), .A2(n9239), .ZN(n8651) );
  OAI211_X1 U10064 ( .C1(n9438), .C2(n8728), .A(n8652), .B(n8651), .ZN(n8653)
         );
  AOI21_X1 U10065 ( .B1(n9427), .B2(n8741), .A(n8653), .ZN(n8654) );
  OAI21_X1 U10066 ( .B1(n8655), .B2(n8766), .A(n8654), .ZN(P1_U3225) );
  NAND2_X1 U10067 ( .A1(n8657), .A2(n8656), .ZN(n8667) );
  INV_X1 U10068 ( .A(n8658), .ZN(n8659) );
  NAND2_X1 U10069 ( .A1(n8660), .A2(n8659), .ZN(n8663) );
  INV_X1 U10070 ( .A(n8661), .ZN(n8662) );
  NAND2_X1 U10071 ( .A1(n8663), .A2(n8662), .ZN(n8664) );
  OAI21_X1 U10072 ( .B1(n8663), .B2(n8662), .A(n8664), .ZN(n8755) );
  NOR2_X1 U10073 ( .A1(n8755), .A2(n8756), .ZN(n8754) );
  INV_X1 U10074 ( .A(n8664), .ZN(n8665) );
  NOR2_X1 U10075 ( .A1(n8754), .A2(n8665), .ZN(n8666) );
  XOR2_X1 U10076 ( .A(n8667), .B(n8666), .Z(n8672) );
  INV_X1 U10077 ( .A(n9473), .ZN(n9491) );
  INV_X1 U10078 ( .A(n9507), .ZN(n9379) );
  NAND2_X1 U10079 ( .A1(n8757), .A2(n9379), .ZN(n8668) );
  NAND2_X1 U10080 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9685) );
  OAI211_X1 U10081 ( .C1(n8759), .C2(n9491), .A(n8668), .B(n9685), .ZN(n8669)
         );
  AOI21_X1 U10082 ( .B1(n9375), .B2(n8763), .A(n8669), .ZN(n8671) );
  NAND2_X1 U10083 ( .A1(n9494), .A2(n8741), .ZN(n8670) );
  OAI211_X1 U10084 ( .C1(n8672), .C2(n8766), .A(n8671), .B(n8670), .ZN(
        P1_U3226) );
  XOR2_X1 U10085 ( .A(n8674), .B(n8673), .Z(n8679) );
  INV_X1 U10086 ( .A(n9499), .ZN(n9363) );
  INV_X1 U10087 ( .A(n9465), .ZN(n9175) );
  NAND2_X1 U10088 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9702) );
  OAI21_X1 U10089 ( .B1(n8759), .B2(n9175), .A(n9702), .ZN(n8675) );
  AOI21_X1 U10090 ( .B1(n8757), .B2(n9363), .A(n8675), .ZN(n8676) );
  OAI21_X1 U10091 ( .B1(n8739), .B2(n9358), .A(n8676), .ZN(n8677) );
  AOI21_X1 U10092 ( .B1(n9487), .B2(n8741), .A(n8677), .ZN(n8678) );
  OAI21_X1 U10093 ( .B1(n8679), .B2(n8766), .A(n8678), .ZN(P1_U3228) );
  AND3_X1 U10094 ( .A1(n8682), .A2(n8681), .A3(n8680), .ZN(n8683) );
  OAI21_X1 U10095 ( .B1(n8684), .B2(n8683), .A(n8748), .ZN(n8688) );
  INV_X1 U10096 ( .A(n9284), .ZN(n9180) );
  AOI22_X1 U10097 ( .A1(n8726), .A2(n9415), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8685) );
  OAI21_X1 U10098 ( .B1(n9180), .B2(n8728), .A(n8685), .ZN(n8686) );
  AOI21_X1 U10099 ( .B1(n9255), .B2(n8763), .A(n8686), .ZN(n8687) );
  OAI211_X1 U10100 ( .C1(n9249), .C2(n8760), .A(n8688), .B(n8687), .ZN(
        P1_U3229) );
  XNOR2_X1 U10101 ( .A(n8691), .B(n8690), .ZN(n8692) );
  XNOR2_X1 U10102 ( .A(n8689), .B(n8692), .ZN(n8697) );
  AOI22_X1 U10103 ( .A1(n8726), .A2(n9283), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n8694) );
  NAND2_X1 U10104 ( .A1(n8757), .A2(n9476), .ZN(n8693) );
  OAI211_X1 U10105 ( .C1(n8739), .C2(n9311), .A(n8694), .B(n8693), .ZN(n8695)
         );
  AOI21_X1 U10106 ( .B1(n9460), .B2(n8741), .A(n8695), .ZN(n8696) );
  OAI21_X1 U10107 ( .B1(n8697), .B2(n8766), .A(n8696), .ZN(P1_U3233) );
  OAI21_X1 U10108 ( .B1(n8700), .B2(n8699), .A(n8698), .ZN(n8701) );
  NAND2_X1 U10109 ( .A1(n8701), .A2(n8748), .ZN(n8707) );
  NAND2_X1 U10110 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9645) );
  INV_X1 U10111 ( .A(n9645), .ZN(n8702) );
  AOI21_X1 U10112 ( .B1(n8757), .B2(n9030), .A(n8702), .ZN(n8703) );
  OAI21_X1 U10113 ( .B1(n9516), .B2(n8759), .A(n8703), .ZN(n8704) );
  AOI21_X1 U10114 ( .B1(n8705), .B2(n8763), .A(n8704), .ZN(n8706) );
  OAI211_X1 U10115 ( .C1(n8708), .C2(n8760), .A(n8707), .B(n8706), .ZN(
        P1_U3234) );
  INV_X1 U10116 ( .A(n8709), .ZN(n8714) );
  OAI21_X1 U10117 ( .B1(n8711), .B2(n8713), .A(n8710), .ZN(n8712) );
  OAI21_X1 U10118 ( .B1(n8714), .B2(n8713), .A(n8712), .ZN(n8715) );
  NAND2_X1 U10119 ( .A1(n8715), .A2(n8748), .ZN(n8719) );
  AOI22_X1 U10120 ( .A1(n8726), .A2(n9284), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8716) );
  OAI21_X1 U10121 ( .B1(n9458), .B2(n8728), .A(n8716), .ZN(n8717) );
  AOI21_X1 U10122 ( .B1(n9278), .B2(n8763), .A(n8717), .ZN(n8718) );
  OAI211_X1 U10123 ( .C1(n9280), .C2(n8760), .A(n8719), .B(n8718), .ZN(
        P1_U3235) );
  INV_X1 U10124 ( .A(n8604), .ZN(n8722) );
  NOR3_X1 U10125 ( .A1(n8722), .A2(n4842), .A3(n8721), .ZN(n8724) );
  OAI21_X1 U10126 ( .B1(n8724), .B2(n8723), .A(n8748), .ZN(n8732) );
  INV_X1 U10127 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8725) );
  NOR2_X1 U10128 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8725), .ZN(n9632) );
  AOI21_X1 U10129 ( .B1(n8726), .B2(n9030), .A(n9632), .ZN(n8727) );
  OAI21_X1 U10130 ( .B1(n9533), .B2(n8728), .A(n8727), .ZN(n8729) );
  AOI21_X1 U10131 ( .B1(n8730), .B2(n8763), .A(n8729), .ZN(n8731) );
  OAI211_X1 U10132 ( .C1(n8733), .C2(n8760), .A(n8732), .B(n8731), .ZN(
        P1_U3236) );
  AOI21_X1 U10133 ( .B1(n8736), .B2(n8735), .A(n8734), .ZN(n8743) );
  NAND2_X1 U10134 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9719) );
  OAI21_X1 U10135 ( .B1(n8759), .B2(n9177), .A(n9719), .ZN(n8737) );
  AOI21_X1 U10136 ( .B1(n8757), .B2(n9473), .A(n8737), .ZN(n8738) );
  OAI21_X1 U10137 ( .B1(n8739), .B2(n9342), .A(n8738), .ZN(n8740) );
  AOI21_X1 U10138 ( .B1(n9350), .B2(n8741), .A(n8740), .ZN(n8742) );
  OAI21_X1 U10139 ( .B1(n8743), .B2(n8766), .A(n8742), .ZN(P1_U3238) );
  INV_X1 U10140 ( .A(n8744), .ZN(n8749) );
  NAND3_X1 U10141 ( .A1(n8749), .A2(n8748), .A3(n8747), .ZN(n8753) );
  AOI22_X1 U10142 ( .A1(n8757), .A2(n9415), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8750) );
  OAI21_X1 U10143 ( .B1(n9198), .B2(n8759), .A(n8750), .ZN(n8751) );
  AOI21_X1 U10144 ( .B1(n9224), .B2(n8763), .A(n8751), .ZN(n8752) );
  OAI211_X1 U10145 ( .C1(n9419), .C2(n8760), .A(n8753), .B(n8752), .ZN(
        P1_U3240) );
  AOI21_X1 U10146 ( .B1(n8756), .B2(n8755), .A(n8754), .ZN(n8767) );
  NAND2_X1 U10147 ( .A1(n8757), .A2(n9028), .ZN(n8758) );
  NAND2_X1 U10148 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9672) );
  OAI211_X1 U10149 ( .C1(n8759), .C2(n9499), .A(n8758), .B(n9672), .ZN(n8762)
         );
  NOR2_X1 U10150 ( .A1(n9170), .A2(n8760), .ZN(n8761) );
  AOI211_X1 U10151 ( .C1(n8764), .C2(n8763), .A(n8762), .B(n8761), .ZN(n8765)
         );
  OAI21_X1 U10152 ( .B1(n8767), .B2(n8766), .A(n8765), .ZN(P1_U3241) );
  NOR2_X1 U10153 ( .A1(n8794), .A2(n9565), .ZN(n8768) );
  INV_X1 U10154 ( .A(n9388), .ZN(n8940) );
  NAND2_X1 U10155 ( .A1(n8769), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U10156 ( .A1(n5072), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U10157 ( .A1(n5101), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8770) );
  NAND3_X1 U10158 ( .A1(n8772), .A2(n8771), .A3(n8770), .ZN(n9142) );
  INV_X1 U10159 ( .A(n9142), .ZN(n8937) );
  NAND2_X1 U10160 ( .A1(n8940), .A2(n8937), .ZN(n9015) );
  INV_X1 U10161 ( .A(n9015), .ZN(n8780) );
  NAND2_X1 U10162 ( .A1(n8773), .A2(n8792), .ZN(n8776) );
  OR2_X1 U10163 ( .A1(n8794), .A2(n8774), .ZN(n8775) );
  NAND2_X1 U10164 ( .A1(n8769), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8779) );
  NAND2_X1 U10165 ( .A1(n5072), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U10166 ( .A1(n5101), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8777) );
  AND3_X1 U10167 ( .A1(n8779), .A2(n8778), .A3(n8777), .ZN(n9164) );
  NOR2_X1 U10168 ( .A1(n9148), .A2(n9164), .ZN(n8938) );
  NOR2_X1 U10169 ( .A1(n8780), .A2(n8938), .ZN(n8983) );
  INV_X1 U10170 ( .A(n9242), .ZN(n9424) );
  OR2_X1 U10171 ( .A1(n9229), .A2(n9424), .ZN(n8923) );
  NAND2_X1 U10172 ( .A1(n8948), .A2(n8923), .ZN(n8790) );
  INV_X1 U10173 ( .A(n8790), .ZN(n8797) );
  NAND2_X1 U10174 ( .A1(n9401), .A2(n9408), .ZN(n8947) );
  NAND2_X1 U10175 ( .A1(n9411), .A2(n9198), .ZN(n9194) );
  NAND2_X1 U10176 ( .A1(n8947), .A2(n9194), .ZN(n9161) );
  OR2_X1 U10177 ( .A1(n9427), .A2(n9227), .ZN(n8833) );
  OR2_X1 U10178 ( .A1(n9441), .A2(n9180), .ZN(n8949) );
  OR2_X1 U10179 ( .A1(n9446), .A2(n9439), .ZN(n8915) );
  AND2_X1 U10180 ( .A1(n8949), .A2(n8915), .ZN(n8834) );
  INV_X1 U10181 ( .A(n8834), .ZN(n8781) );
  NAND2_X1 U10182 ( .A1(n9441), .A2(n9180), .ZN(n9155) );
  NAND2_X1 U10183 ( .A1(n8781), .A2(n9155), .ZN(n8782) );
  NAND2_X1 U10184 ( .A1(n9156), .A2(n8782), .ZN(n8783) );
  NAND2_X1 U10185 ( .A1(n9433), .A2(n9438), .ZN(n8921) );
  NAND2_X1 U10186 ( .A1(n8783), .A2(n8921), .ZN(n8784) );
  AND2_X1 U10187 ( .A1(n8833), .A2(n8784), .ZN(n8799) );
  NAND2_X1 U10188 ( .A1(n9446), .A2(n9439), .ZN(n9153) );
  AND2_X1 U10189 ( .A1(n9155), .A2(n9153), .ZN(n8835) );
  NAND2_X1 U10190 ( .A1(n9295), .A2(n9283), .ZN(n8992) );
  NAND2_X1 U10191 ( .A1(n9460), .A2(n9328), .ZN(n8907) );
  NAND2_X1 U10192 ( .A1(n8992), .A2(n4621), .ZN(n8785) );
  NAND2_X1 U10193 ( .A1(n9451), .A2(n9458), .ZN(n9152) );
  NAND2_X1 U10194 ( .A1(n8785), .A2(n9152), .ZN(n8911) );
  INV_X1 U10195 ( .A(n8911), .ZN(n8786) );
  NAND3_X1 U10196 ( .A1(n8921), .A2(n8835), .A3(n8786), .ZN(n8788) );
  NAND2_X1 U10197 ( .A1(n9427), .A2(n9227), .ZN(n9157) );
  INV_X1 U10198 ( .A(n9157), .ZN(n8787) );
  AOI21_X1 U10199 ( .B1(n8799), .B2(n8788), .A(n8787), .ZN(n8789) );
  NOR2_X1 U10200 ( .A1(n8790), .A2(n8789), .ZN(n8791) );
  OR2_X1 U10201 ( .A1(n9161), .A2(n8791), .ZN(n8798) );
  NAND2_X1 U10202 ( .A1(n8793), .A2(n8792), .ZN(n8796) );
  OR2_X1 U10203 ( .A1(n8794), .A2(n10018), .ZN(n8795) );
  OAI211_X1 U10204 ( .C1(n8797), .C2(n8798), .A(n8935), .B(n9160), .ZN(n8994)
         );
  NAND2_X1 U10205 ( .A1(n9229), .A2(n9424), .ZN(n9159) );
  NOR2_X1 U10206 ( .A1(n8798), .A2(n4810), .ZN(n8996) );
  INV_X1 U10207 ( .A(n8996), .ZN(n8827) );
  INV_X1 U10208 ( .A(n8799), .ZN(n8800) );
  NOR2_X1 U10209 ( .A1(n8800), .A2(n4838), .ZN(n8993) );
  INV_X1 U10210 ( .A(n8993), .ZN(n8825) );
  OR2_X1 U10211 ( .A1(n9324), .A2(n9177), .ZN(n8950) );
  OR2_X1 U10212 ( .A1(n9350), .A2(n9175), .ZN(n8951) );
  NAND2_X1 U10213 ( .A1(n8950), .A2(n8951), .ZN(n8903) );
  NAND2_X1 U10214 ( .A1(n9350), .A2(n9175), .ZN(n8989) );
  NAND2_X1 U10215 ( .A1(n9487), .A2(n9491), .ZN(n8801) );
  AND2_X1 U10216 ( .A1(n8989), .A2(n8801), .ZN(n8904) );
  NAND2_X1 U10217 ( .A1(n9041), .A2(n6693), .ZN(n8802) );
  AND4_X1 U10218 ( .A1(n8804), .A2(n8803), .A3(n8957), .A4(n8802), .ZN(n8807)
         );
  NAND2_X1 U10219 ( .A1(n9038), .A2(n9755), .ZN(n8805) );
  AND4_X1 U10220 ( .A1(n8807), .A2(n8843), .A3(n8806), .A4(n8805), .ZN(n8809)
         );
  OAI211_X1 U10221 ( .C1(n8810), .C2(n8809), .A(n8874), .B(n8808), .ZN(n8812)
         );
  NAND2_X1 U10222 ( .A1(n8878), .A2(n8872), .ZN(n8866) );
  INV_X1 U10223 ( .A(n8866), .ZN(n8811) );
  NAND2_X1 U10224 ( .A1(n8880), .A2(n8875), .ZN(n8868) );
  AOI21_X1 U10225 ( .B1(n8812), .B2(n8811), .A(n8868), .ZN(n8814) );
  NAND2_X1 U10226 ( .A1(n8891), .A2(n8877), .ZN(n8813) );
  OAI211_X1 U10227 ( .C1(n8814), .C2(n8813), .A(n8886), .B(n8893), .ZN(n8815)
         );
  INV_X1 U10228 ( .A(n8815), .ZN(n8820) );
  NAND2_X1 U10229 ( .A1(n9494), .A2(n9499), .ZN(n8986) );
  NAND2_X1 U10230 ( .A1(n9502), .A2(n9507), .ZN(n8984) );
  NAND2_X1 U10231 ( .A1(n8986), .A2(n8984), .ZN(n8895) );
  INV_X1 U10232 ( .A(n8816), .ZN(n8817) );
  AND2_X1 U10233 ( .A1(n9357), .A2(n9473), .ZN(n9337) );
  INV_X1 U10234 ( .A(n9337), .ZN(n8900) );
  NAND2_X1 U10235 ( .A1(n9170), .A2(n9379), .ZN(n8836) );
  AND2_X1 U10236 ( .A1(n8952), .A2(n8836), .ZN(n8887) );
  INV_X1 U10237 ( .A(n8887), .ZN(n8818) );
  NAND2_X1 U10238 ( .A1(n8818), .A2(n8986), .ZN(n8819) );
  OAI211_X1 U10239 ( .C1(n8820), .C2(n4406), .A(n8900), .B(n8819), .ZN(n8821)
         );
  AND2_X1 U10240 ( .A1(n8904), .A2(n8821), .ZN(n8822) );
  NAND2_X1 U10241 ( .A1(n9324), .A2(n9177), .ZN(n8990) );
  OAI21_X1 U10242 ( .B1(n8903), .B2(n8822), .A(n8990), .ZN(n8823) );
  NAND2_X1 U10243 ( .A1(n8992), .A2(n8823), .ZN(n8824) );
  NOR2_X1 U10244 ( .A1(n8825), .A2(n8824), .ZN(n8826) );
  NOR2_X1 U10245 ( .A1(n8827), .A2(n8826), .ZN(n8828) );
  NAND2_X1 U10246 ( .A1(n9148), .A2(n9164), .ZN(n8981) );
  NAND2_X1 U10247 ( .A1(n9394), .A2(n9197), .ZN(n8997) );
  OAI211_X1 U10248 ( .C1(n8994), .C2(n8828), .A(n8981), .B(n8997), .ZN(n8829)
         );
  AND2_X1 U10249 ( .A1(n9388), .A2(n9142), .ZN(n9001) );
  AOI21_X1 U10250 ( .B1(n8983), .B2(n8829), .A(n9001), .ZN(n8830) );
  XNOR2_X1 U10251 ( .A(n8830), .B(n7703), .ZN(n9008) );
  NAND2_X1 U10252 ( .A1(n9159), .A2(n9157), .ZN(n8831) );
  INV_X1 U10253 ( .A(n9016), .ZN(n8943) );
  NAND3_X1 U10254 ( .A1(n8831), .A2(n8943), .A3(n8923), .ZN(n8928) );
  NAND2_X1 U10255 ( .A1(n8923), .A2(n8833), .ZN(n8832) );
  NAND2_X1 U10256 ( .A1(n8832), .A2(n9016), .ZN(n8924) );
  MUX2_X1 U10257 ( .A(n8835), .B(n8834), .S(n8943), .Z(n8918) );
  INV_X1 U10258 ( .A(n8836), .ZN(n8837) );
  NAND2_X1 U10259 ( .A1(n8986), .A2(n8837), .ZN(n8890) );
  NAND4_X1 U10260 ( .A1(n8840), .A2(n8839), .A3(n8838), .A4(n9016), .ZN(n8864)
         );
  NAND2_X1 U10261 ( .A1(n7013), .A2(n8841), .ZN(n8844) );
  NAND3_X1 U10262 ( .A1(n8844), .A2(n8843), .A3(n8842), .ZN(n8846) );
  NAND2_X1 U10263 ( .A1(n8846), .A2(n8845), .ZN(n8863) );
  AND3_X1 U10264 ( .A1(n8847), .A2(n8943), .A3(n8965), .ZN(n8862) );
  NAND2_X1 U10265 ( .A1(n8848), .A2(n8943), .ZN(n8856) );
  OAI21_X1 U10266 ( .B1(n8856), .B2(n9034), .A(n8849), .ZN(n8853) );
  OR2_X1 U10267 ( .A1(n8848), .A2(n8943), .ZN(n8850) );
  OAI21_X1 U10268 ( .B1(n8850), .B2(n8854), .A(n8857), .ZN(n8852) );
  OAI22_X1 U10269 ( .A1(n8850), .A2(n8849), .B1(n8854), .B2(n8943), .ZN(n8851)
         );
  AOI22_X1 U10270 ( .A1(n8853), .A2(n8852), .B1(n8851), .B2(n9770), .ZN(n8861)
         );
  NAND2_X1 U10271 ( .A1(n8854), .A2(n8943), .ZN(n8855) );
  OAI21_X1 U10272 ( .B1(n8857), .B2(n8856), .A(n8855), .ZN(n8859) );
  NAND2_X1 U10273 ( .A1(n8859), .A2(n8858), .ZN(n8860) );
  NAND2_X1 U10274 ( .A1(n8871), .A2(n8865), .ZN(n8867) );
  AOI21_X1 U10275 ( .B1(n8867), .B2(n8874), .A(n8866), .ZN(n8869) );
  OAI21_X1 U10276 ( .B1(n8869), .B2(n8868), .A(n8877), .ZN(n8883) );
  NAND2_X1 U10277 ( .A1(n8871), .A2(n8870), .ZN(n8873) );
  NAND2_X1 U10278 ( .A1(n8873), .A2(n8872), .ZN(n8876) );
  NAND3_X1 U10279 ( .A1(n8876), .A2(n8875), .A3(n8874), .ZN(n8879) );
  NAND3_X1 U10280 ( .A1(n8879), .A2(n8878), .A3(n8877), .ZN(n8881) );
  NAND2_X1 U10281 ( .A1(n8881), .A2(n8880), .ZN(n8882) );
  NAND2_X1 U10282 ( .A1(n8892), .A2(n8893), .ZN(n8885) );
  NAND3_X1 U10283 ( .A1(n8885), .A2(n7487), .A3(n8891), .ZN(n8888) );
  NAND3_X1 U10284 ( .A1(n8888), .A2(n8887), .A3(n8886), .ZN(n8889) );
  NAND2_X1 U10285 ( .A1(n8894), .A2(n8943), .ZN(n8897) );
  NAND3_X1 U10286 ( .A1(n8895), .A2(n8952), .A3(n9016), .ZN(n8896) );
  NAND3_X1 U10287 ( .A1(n8898), .A2(n8897), .A3(n8896), .ZN(n8899) );
  XNOR2_X1 U10288 ( .A(n9487), .B(n9473), .ZN(n9361) );
  AND2_X1 U10289 ( .A1(n8951), .A2(n8900), .ZN(n8902) );
  NAND2_X1 U10290 ( .A1(n8990), .A2(n8989), .ZN(n8901) );
  NAND2_X1 U10291 ( .A1(n9151), .A2(n8943), .ZN(n8905) );
  NAND2_X1 U10292 ( .A1(n8906), .A2(n8950), .ZN(n8909) );
  NAND3_X1 U10293 ( .A1(n8907), .A2(n9476), .A3(n9016), .ZN(n8908) );
  NAND2_X1 U10294 ( .A1(n8909), .A2(n8908), .ZN(n8910) );
  NAND2_X1 U10295 ( .A1(n8992), .A2(n9151), .ZN(n8912) );
  MUX2_X1 U10296 ( .A(n8912), .B(n8911), .S(n8943), .Z(n8913) );
  OAI22_X1 U10297 ( .A1(n8914), .A2(n8913), .B1(n8943), .B2(n9152), .ZN(n8916)
         );
  NAND2_X1 U10298 ( .A1(n8916), .A2(n9281), .ZN(n8917) );
  INV_X1 U10299 ( .A(n9251), .ZN(n8920) );
  MUX2_X1 U10300 ( .A(n9155), .B(n8949), .S(n9016), .Z(n8919) );
  MUX2_X1 U10301 ( .A(n8921), .B(n9156), .S(n8943), .Z(n8922) );
  NAND2_X1 U10302 ( .A1(n8925), .A2(n9159), .ZN(n8927) );
  INV_X1 U10303 ( .A(n8948), .ZN(n8926) );
  AOI21_X1 U10304 ( .B1(n8928), .B2(n8927), .A(n8926), .ZN(n8929) );
  NAND2_X1 U10305 ( .A1(n8930), .A2(n9160), .ZN(n8933) );
  OAI21_X1 U10306 ( .B1(n9161), .B2(n8948), .A(n9160), .ZN(n8931) );
  NAND2_X1 U10307 ( .A1(n8931), .A2(n9016), .ZN(n8932) );
  NAND2_X1 U10308 ( .A1(n8933), .A2(n8932), .ZN(n8934) );
  MUX2_X1 U10309 ( .A(n8997), .B(n8935), .S(n9016), .Z(n8936) );
  NOR2_X1 U10310 ( .A1(n8937), .A2(n9164), .ZN(n8998) );
  NAND2_X1 U10311 ( .A1(n8938), .A2(n8940), .ZN(n9003) );
  INV_X1 U10312 ( .A(n9164), .ZN(n9025) );
  NAND4_X1 U10313 ( .A1(n8941), .A2(n8940), .A3(n9025), .A4(n9148), .ZN(n8942)
         );
  OAI21_X1 U10314 ( .B1(n9003), .B2(n8943), .A(n8942), .ZN(n8944) );
  NOR2_X1 U10315 ( .A1(n8945), .A2(n8944), .ZN(n9013) );
  XNOR2_X1 U10316 ( .A(n9451), .B(n9458), .ZN(n9296) );
  NAND2_X1 U10317 ( .A1(n8949), .A2(n9155), .ZN(n9262) );
  INV_X1 U10318 ( .A(n9305), .ZN(n9310) );
  NAND2_X1 U10319 ( .A1(n8951), .A2(n8989), .ZN(n9336) );
  INV_X1 U10320 ( .A(n9361), .ZN(n8976) );
  INV_X1 U10321 ( .A(n8954), .ZN(n8967) );
  NOR4_X1 U10322 ( .A1(n8958), .A2(n8957), .A3(n8956), .A4(n8955), .ZN(n8959)
         );
  NAND2_X1 U10323 ( .A1(n8960), .A2(n8959), .ZN(n8964) );
  NOR4_X1 U10324 ( .A1(n8964), .A2(n8963), .A3(n8962), .A4(n8961), .ZN(n8966)
         );
  NAND4_X1 U10325 ( .A1(n7140), .A2(n8967), .A3(n8966), .A4(n8965), .ZN(n8968)
         );
  NOR4_X1 U10326 ( .A1(n8971), .A2(n8970), .A3(n8969), .A4(n8968), .ZN(n8972)
         );
  NAND4_X1 U10327 ( .A1(n9372), .A2(n7487), .A3(n8973), .A4(n8972), .ZN(n8974)
         );
  NOR4_X1 U10328 ( .A1(n9336), .A2(n8976), .A3(n8975), .A4(n8974), .ZN(n8977)
         );
  NAND4_X1 U10329 ( .A1(n9281), .A2(n9322), .A3(n9310), .A4(n8977), .ZN(n8978)
         );
  NOR4_X1 U10330 ( .A1(n9251), .A2(n9296), .A3(n9262), .A4(n8978), .ZN(n8979)
         );
  NAND4_X1 U10331 ( .A1(n9209), .A2(n9235), .A3(n8979), .A4(n9221), .ZN(n8980)
         );
  NOR3_X1 U10332 ( .A1(n4531), .A2(n4806), .A3(n8980), .ZN(n8982) );
  INV_X1 U10333 ( .A(n9001), .ZN(n9021) );
  NAND4_X1 U10334 ( .A1(n8983), .A2(n8982), .A3(n9021), .A4(n8981), .ZN(n9007)
         );
  NAND2_X1 U10335 ( .A1(n8985), .A2(n8984), .ZN(n9370) );
  INV_X1 U10336 ( .A(n8986), .ZN(n8987) );
  NAND2_X1 U10337 ( .A1(n9362), .A2(n9361), .ZN(n9335) );
  NOR2_X1 U10338 ( .A1(n9336), .A2(n9337), .ZN(n8988) );
  NAND2_X1 U10339 ( .A1(n9335), .A2(n8988), .ZN(n9339) );
  NAND2_X1 U10340 ( .A1(n9339), .A2(n8989), .ZN(n9323) );
  NAND2_X1 U10341 ( .A1(n9323), .A2(n9322), .ZN(n8991) );
  NAND3_X1 U10342 ( .A1(n8993), .A2(n8992), .A3(n9306), .ZN(n8995) );
  AOI21_X1 U10343 ( .B1(n8996), .B2(n8995), .A(n8994), .ZN(n9000) );
  OAI21_X1 U10344 ( .B1(n9391), .B2(n8998), .A(n8997), .ZN(n8999) );
  NOR3_X1 U10345 ( .A1(n9001), .A2(n9000), .A3(n8999), .ZN(n9005) );
  NAND3_X1 U10346 ( .A1(n9003), .A2(n9002), .A3(n9015), .ZN(n9004) );
  OAI21_X1 U10347 ( .B1(n9005), .B2(n9004), .A(n9007), .ZN(n9006) );
  NAND4_X1 U10348 ( .A1(n9009), .A2(n9614), .A3(n9474), .A4(n5731), .ZN(n9012)
         );
  INV_X1 U10349 ( .A(n9024), .ZN(n9011) );
  NAND2_X1 U10350 ( .A1(n9011), .A2(n9010), .ZN(n9018) );
  NAND3_X1 U10351 ( .A1(n9012), .A2(P1_B_REG_SCAN_IN), .A3(n9018), .ZN(n9023)
         );
  INV_X1 U10352 ( .A(n9013), .ZN(n9014) );
  OAI21_X1 U10353 ( .B1(n9016), .B2(n9015), .A(n9014), .ZN(n9020) );
  NOR2_X1 U10354 ( .A1(n9018), .A2(n9017), .ZN(n9019) );
  OAI211_X1 U10355 ( .C1(n9021), .C2(n7703), .A(n9020), .B(n9019), .ZN(n9022)
         );
  MUX2_X1 U10356 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9142), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10357 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9025), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10358 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9026), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10359 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9166), .S(P1_U3973), .Z(
        P1_U3582) );
  INV_X1 U10360 ( .A(n9198), .ZN(n9416) );
  MUX2_X1 U10361 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9416), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10362 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9242), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9415), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10364 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9027), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10365 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9284), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10366 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9299), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9283), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10368 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9466), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10369 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9476), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10370 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9465), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10371 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9473), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10372 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9363), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10373 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9379), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10374 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9028), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10375 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9029), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10376 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9030), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9031), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10378 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9032), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10379 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9033), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10380 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9034), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9035), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10382 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9036), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9037), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10384 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9038), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9039), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9040), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9041), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10388 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9042), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10389 ( .C1(n9045), .C2(n9044), .A(n9696), .B(n9043), .ZN(n9053)
         );
  OAI211_X1 U10390 ( .C1(n9048), .C2(n9047), .A(n9692), .B(n9046), .ZN(n9052)
         );
  AOI22_X1 U10391 ( .A1(n9616), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9051) );
  NAND2_X1 U10392 ( .A1(n9718), .A2(n9049), .ZN(n9050) );
  NAND4_X1 U10393 ( .A1(n9053), .A2(n9052), .A3(n9051), .A4(n9050), .ZN(
        P1_U3244) );
  INV_X1 U10394 ( .A(n9054), .ZN(n9058) );
  INV_X1 U10395 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9056) );
  OAI21_X1 U10396 ( .B1(n9721), .B2(n9056), .A(n9055), .ZN(n9057) );
  AOI21_X1 U10397 ( .B1(n9058), .B2(n9718), .A(n9057), .ZN(n9067) );
  OAI211_X1 U10398 ( .C1(n9061), .C2(n9060), .A(n9692), .B(n9059), .ZN(n9066)
         );
  OAI211_X1 U10399 ( .C1(n9064), .C2(n9063), .A(n9696), .B(n9062), .ZN(n9065)
         );
  NAND3_X1 U10400 ( .A1(n9067), .A2(n9066), .A3(n9065), .ZN(P1_U3246) );
  AOI211_X1 U10401 ( .C1(n9070), .C2(n9069), .A(n9068), .B(n9711), .ZN(n9071)
         );
  INV_X1 U10402 ( .A(n9071), .ZN(n9081) );
  INV_X1 U10403 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9073) );
  OAI21_X1 U10404 ( .B1(n9721), .B2(n9073), .A(n9072), .ZN(n9074) );
  AOI21_X1 U10405 ( .B1(n9075), .B2(n9718), .A(n9074), .ZN(n9080) );
  OAI211_X1 U10406 ( .C1(n9078), .C2(n9077), .A(n9696), .B(n9076), .ZN(n9079)
         );
  NAND3_X1 U10407 ( .A1(n9081), .A2(n9080), .A3(n9079), .ZN(P1_U3248) );
  AOI211_X1 U10408 ( .C1(n9084), .C2(n9083), .A(n9082), .B(n9711), .ZN(n9085)
         );
  INV_X1 U10409 ( .A(n9085), .ZN(n9095) );
  OAI21_X1 U10410 ( .B1(n9721), .B2(n9087), .A(n9086), .ZN(n9088) );
  AOI21_X1 U10411 ( .B1(n9089), .B2(n9718), .A(n9088), .ZN(n9094) );
  OAI211_X1 U10412 ( .C1(n9092), .C2(n9091), .A(n9696), .B(n9090), .ZN(n9093)
         );
  NAND3_X1 U10413 ( .A1(n9095), .A2(n9094), .A3(n9093), .ZN(P1_U3249) );
  OAI21_X1 U10414 ( .B1(n9098), .B2(n9097), .A(n9096), .ZN(n9099) );
  NAND2_X1 U10415 ( .A1(n9099), .A2(n9692), .ZN(n9109) );
  OAI21_X1 U10416 ( .B1(n9102), .B2(n9101), .A(n9100), .ZN(n9103) );
  NAND2_X1 U10417 ( .A1(n9103), .A2(n9696), .ZN(n9108) );
  AOI21_X1 U10418 ( .B1(n9616), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9104), .ZN(
        n9107) );
  NAND2_X1 U10419 ( .A1(n9718), .A2(n9105), .ZN(n9106) );
  NAND4_X1 U10420 ( .A1(n9109), .A2(n9108), .A3(n9107), .A4(n9106), .ZN(
        P1_U3252) );
  INV_X1 U10421 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9981) );
  XNOR2_X1 U10422 ( .A(n9688), .B(n9981), .ZN(n9690) );
  NAND2_X1 U10423 ( .A1(n9644), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9111) );
  OAI21_X1 U10424 ( .B1(n9644), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9111), .ZN(
        n9640) );
  OAI21_X1 U10425 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9123), .A(n9112), .ZN(
        n9641) );
  NOR2_X1 U10426 ( .A1(n9640), .A2(n9641), .ZN(n9639) );
  INV_X1 U10427 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9113) );
  AOI22_X1 U10428 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9658), .B1(n9124), .B2(
        n9113), .ZN(n9650) );
  NOR2_X1 U10429 ( .A1(n9114), .A2(n9126), .ZN(n9115) );
  INV_X1 U10430 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9667) );
  NOR2_X1 U10431 ( .A1(n9667), .A2(n9668), .ZN(n9666) );
  NOR2_X1 U10432 ( .A1(n9115), .A2(n9666), .ZN(n9681) );
  NAND2_X1 U10433 ( .A1(n9128), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9116) );
  OAI21_X1 U10434 ( .B1(n9128), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9116), .ZN(
        n9680) );
  NOR2_X1 U10435 ( .A1(n9681), .A2(n9680), .ZN(n9679) );
  AOI21_X1 U10436 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9128), .A(n9679), .ZN(
        n9689) );
  NAND2_X1 U10437 ( .A1(n9690), .A2(n9689), .ZN(n9118) );
  OR2_X1 U10438 ( .A1(n9688), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9117) );
  NAND2_X1 U10439 ( .A1(n9118), .A2(n9117), .ZN(n9713) );
  NAND2_X1 U10440 ( .A1(n9717), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9119) );
  OAI21_X1 U10441 ( .B1(n9717), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9119), .ZN(
        n9714) );
  NAND2_X1 U10442 ( .A1(n9710), .A2(n9119), .ZN(n9120) );
  XNOR2_X1 U10443 ( .A(n9120), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9134) );
  INV_X1 U10444 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9121) );
  XNOR2_X1 U10445 ( .A(n9688), .B(n9121), .ZN(n9694) );
  XOR2_X1 U10446 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9128), .Z(n9676) );
  XNOR2_X1 U10447 ( .A(n9644), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9637) );
  OAI21_X1 U10448 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n9123), .A(n9122), .ZN(
        n9638) );
  NOR2_X1 U10449 ( .A1(n9637), .A2(n9638), .ZN(n9636) );
  AOI21_X1 U10450 ( .B1(n9644), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9636), .ZN(
        n9654) );
  XNOR2_X1 U10451 ( .A(n9124), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9653) );
  NOR2_X1 U10452 ( .A1(n9654), .A2(n9653), .ZN(n9652) );
  AOI21_X1 U10453 ( .B1(n9124), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9652), .ZN(
        n9125) );
  NOR2_X1 U10454 ( .A1(n9125), .A2(n9126), .ZN(n9127) );
  INV_X1 U10455 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9664) );
  XNOR2_X1 U10456 ( .A(n9126), .B(n9125), .ZN(n9665) );
  NOR2_X1 U10457 ( .A1(n9664), .A2(n9665), .ZN(n9663) );
  NOR2_X1 U10458 ( .A1(n9127), .A2(n9663), .ZN(n9677) );
  NAND2_X1 U10459 ( .A1(n9676), .A2(n9677), .ZN(n9675) );
  OAI21_X1 U10460 ( .B1(n9128), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9675), .ZN(
        n9693) );
  NAND2_X1 U10461 ( .A1(n9694), .A2(n9693), .ZN(n9130) );
  OR2_X1 U10462 ( .A1(n9688), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U10463 ( .A1(n9130), .A2(n9129), .ZN(n9709) );
  NAND2_X1 U10464 ( .A1(n9717), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9131) );
  OAI21_X1 U10465 ( .B1(n9717), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9131), .ZN(
        n9708) );
  OR2_X1 U10466 ( .A1(n9709), .A2(n9708), .ZN(n9705) );
  NAND2_X1 U10467 ( .A1(n9705), .A2(n9131), .ZN(n9133) );
  INV_X1 U10468 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9132) );
  OAI22_X1 U10469 ( .A1(n9134), .A2(n9711), .B1(n9706), .B2(n4333), .ZN(n9137)
         );
  AOI21_X1 U10470 ( .B1(n9692), .B2(n9134), .A(n9718), .ZN(n9135) );
  INV_X1 U10471 ( .A(n9394), .ZN(n9188) );
  NAND2_X1 U10472 ( .A1(n9391), .A2(n9186), .ZN(n9145) );
  XNOR2_X1 U10473 ( .A(n9388), .B(n9145), .ZN(n9139) );
  NAND2_X1 U10474 ( .A1(n9139), .A2(n9452), .ZN(n9387) );
  NAND2_X1 U10475 ( .A1(n9614), .A2(P1_B_REG_SCAN_IN), .ZN(n9140) );
  NAND2_X1 U10476 ( .A1(n9475), .A2(n9140), .ZN(n9163) );
  INV_X1 U10477 ( .A(n9163), .ZN(n9141) );
  NAND2_X1 U10478 ( .A1(n9142), .A2(n9141), .ZN(n9389) );
  NOR2_X1 U10479 ( .A1(n4322), .A2(n9389), .ZN(n9147) );
  NOR2_X1 U10480 ( .A1(n9388), .A2(n9738), .ZN(n9143) );
  AOI211_X1 U10481 ( .C1(n4322), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9147), .B(
        n9143), .ZN(n9144) );
  OAI21_X1 U10482 ( .B1(n9387), .B2(n9735), .A(n9144), .ZN(P1_U3263) );
  OAI211_X1 U10483 ( .C1(n9391), .C2(n9186), .A(n9452), .B(n9145), .ZN(n9390)
         );
  AND2_X1 U10484 ( .A1(n4322), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9146) );
  NOR2_X1 U10485 ( .A1(n9147), .A2(n9146), .ZN(n9150) );
  NAND2_X1 U10486 ( .A1(n9148), .A2(n9349), .ZN(n9149) );
  OAI211_X1 U10487 ( .C1(n9390), .C2(n9735), .A(n9150), .B(n9149), .ZN(
        P1_U3264) );
  NAND2_X2 U10488 ( .A1(n9297), .A2(n9152), .ZN(n9282) );
  INV_X1 U10489 ( .A(n9153), .ZN(n9154) );
  NAND2_X1 U10490 ( .A1(n9236), .A2(n9235), .ZN(n9234) );
  NAND2_X1 U10491 ( .A1(n9234), .A2(n9157), .ZN(n9222) );
  INV_X1 U10492 ( .A(n9209), .ZN(n9158) );
  XNOR2_X1 U10493 ( .A(n9162), .B(n9185), .ZN(n9168) );
  AOI21_X1 U10494 ( .B1(n9169), .B2(n9722), .A(n9398), .ZN(n9192) );
  NOR2_X1 U10495 ( .A1(n9487), .A2(n9473), .ZN(n9173) );
  OAI22_X1 U10496 ( .A1(n9355), .A2(n9173), .B1(n9491), .B2(n9357), .ZN(n9174)
         );
  INV_X1 U10497 ( .A(n9174), .ZN(n9334) );
  INV_X1 U10498 ( .A(n9350), .ZN(n9479) );
  NAND2_X1 U10499 ( .A1(n4623), .A2(n9177), .ZN(n9178) );
  NAND2_X1 U10500 ( .A1(n9441), .A2(n9284), .ZN(n9181) );
  NAND2_X1 U10501 ( .A1(n9249), .A2(n9438), .ZN(n9183) );
  NOR2_X1 U10502 ( .A1(n9249), .A2(n9438), .ZN(n9182) );
  NAND2_X1 U10503 ( .A1(n9229), .A2(n9242), .ZN(n9184) );
  NAND2_X1 U10504 ( .A1(n9392), .A2(n9742), .ZN(n9191) );
  AOI211_X1 U10505 ( .C1(n9394), .C2(n4583), .A(n9771), .B(n9186), .ZN(n9393)
         );
  INV_X1 U10506 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9187) );
  OAI22_X1 U10507 ( .A1(n9188), .A2(n9738), .B1(n9187), .B2(n9366), .ZN(n9189)
         );
  AOI21_X1 U10508 ( .B1(n9393), .B2(n9724), .A(n9189), .ZN(n9190) );
  OAI211_X1 U10509 ( .C1(n4322), .C2(n9192), .A(n9191), .B(n9190), .ZN(
        P1_U3356) );
  OAI222_X1 U10510 ( .A1(n9532), .A2(n9198), .B1(n9530), .B2(n9197), .C1(n9196), .C2(n9523), .ZN(n9403) );
  AOI211_X1 U10511 ( .C1(n9401), .C2(n9210), .A(n9771), .B(n9199), .ZN(n9402)
         );
  NAND2_X1 U10512 ( .A1(n9402), .A2(n9724), .ZN(n9202) );
  AOI22_X1 U10513 ( .A1(n4322), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9200), .B2(
        n9722), .ZN(n9201) );
  OAI211_X1 U10514 ( .C1(n4581), .C2(n9738), .A(n9202), .B(n9201), .ZN(n9203)
         );
  AOI21_X1 U10515 ( .B1(n9403), .B2(n9366), .A(n9203), .ZN(n9204) );
  OAI21_X1 U10516 ( .B1(n9406), .B2(n9369), .A(n9204), .ZN(P1_U3265) );
  NOR2_X1 U10517 ( .A1(n9209), .A2(n4810), .ZN(n9207) );
  AOI21_X1 U10518 ( .B1(n9207), .B2(n9205), .A(n9206), .ZN(n9414) );
  XNOR2_X1 U10519 ( .A(n9208), .B(n9209), .ZN(n9407) );
  NAND2_X1 U10520 ( .A1(n9407), .A2(n9742), .ZN(n9219) );
  INV_X1 U10521 ( .A(n9210), .ZN(n9211) );
  AOI211_X1 U10522 ( .C1(n9411), .C2(n9223), .A(n9771), .B(n9211), .ZN(n9409)
         );
  INV_X1 U10523 ( .A(n9377), .ZN(n9345) );
  AOI22_X1 U10524 ( .A1(n4322), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9212), .B2(
        n9722), .ZN(n9213) );
  OAI21_X1 U10525 ( .B1(n9347), .B2(n9424), .A(n9213), .ZN(n9214) );
  AOI21_X1 U10526 ( .B1(n9345), .B2(n9166), .A(n9214), .ZN(n9215) );
  OAI21_X1 U10527 ( .B1(n9216), .B2(n9738), .A(n9215), .ZN(n9217) );
  AOI21_X1 U10528 ( .B1(n9409), .B2(n9724), .A(n9217), .ZN(n9218) );
  OAI211_X1 U10529 ( .C1(n9414), .C2(n9386), .A(n9219), .B(n9218), .ZN(
        P1_U3266) );
  XNOR2_X1 U10530 ( .A(n9220), .B(n9221), .ZN(n9423) );
  OAI21_X1 U10531 ( .B1(n9222), .B2(n9221), .A(n9205), .ZN(n9421) );
  INV_X1 U10532 ( .A(n9386), .ZN(n9353) );
  OAI211_X1 U10533 ( .C1(n9419), .C2(n9237), .A(n9452), .B(n9223), .ZN(n9418)
         );
  NAND2_X1 U10534 ( .A1(n9345), .A2(n9416), .ZN(n9226) );
  AOI22_X1 U10535 ( .A1(n4322), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9224), .B2(
        n9722), .ZN(n9225) );
  OAI211_X1 U10536 ( .C1(n9227), .C2(n9347), .A(n9226), .B(n9225), .ZN(n9228)
         );
  AOI21_X1 U10537 ( .B1(n9229), .B2(n9349), .A(n9228), .ZN(n9230) );
  OAI21_X1 U10538 ( .B1(n9418), .B2(n9735), .A(n9230), .ZN(n9231) );
  AOI21_X1 U10539 ( .B1(n9421), .B2(n9353), .A(n9231), .ZN(n9232) );
  OAI21_X1 U10540 ( .B1(n9423), .B2(n9369), .A(n9232), .ZN(P1_U3267) );
  XNOR2_X1 U10541 ( .A(n9233), .B(n9235), .ZN(n9431) );
  OAI21_X1 U10542 ( .B1(n9236), .B2(n9235), .A(n9234), .ZN(n9428) );
  INV_X1 U10543 ( .A(n9254), .ZN(n9238) );
  AOI211_X1 U10544 ( .C1(n9427), .C2(n9238), .A(n9771), .B(n9237), .ZN(n9425)
         );
  NAND2_X1 U10545 ( .A1(n9425), .A2(n9724), .ZN(n9244) );
  AOI22_X1 U10546 ( .A1(n4322), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9239), .B2(
        n9722), .ZN(n9240) );
  OAI21_X1 U10547 ( .B1(n9347), .B2(n9438), .A(n9240), .ZN(n9241) );
  AOI21_X1 U10548 ( .B1(n9345), .B2(n9242), .A(n9241), .ZN(n9243) );
  OAI211_X1 U10549 ( .C1(n9245), .C2(n9738), .A(n9244), .B(n9243), .ZN(n9246)
         );
  AOI21_X1 U10550 ( .B1(n9428), .B2(n9353), .A(n9246), .ZN(n9247) );
  OAI21_X1 U10551 ( .B1(n9431), .B2(n9369), .A(n9247), .ZN(P1_U3268) );
  XNOR2_X1 U10552 ( .A(n9248), .B(n9251), .ZN(n9436) );
  NOR2_X1 U10553 ( .A1(n9249), .A2(n9738), .ZN(n9258) );
  AND2_X1 U10554 ( .A1(n9284), .A2(n9474), .ZN(n9253) );
  AOI211_X1 U10555 ( .C1(n9251), .C2(n9250), .A(n9523), .B(n4369), .ZN(n9252)
         );
  AOI211_X1 U10556 ( .C1(n9475), .C2(n9415), .A(n9253), .B(n9252), .ZN(n9435)
         );
  AOI211_X1 U10557 ( .C1(n9433), .C2(n9266), .A(n9771), .B(n9254), .ZN(n9432)
         );
  AOI22_X1 U10558 ( .A1(n9432), .A2(n7703), .B1(n9722), .B2(n9255), .ZN(n9256)
         );
  AOI21_X1 U10559 ( .B1(n9435), .B2(n9256), .A(n4322), .ZN(n9257) );
  AOI211_X1 U10560 ( .C1(n4322), .C2(P1_REG2_REG_24__SCAN_IN), .A(n9258), .B(
        n9257), .ZN(n9259) );
  OAI21_X1 U10561 ( .B1(n9436), .B2(n9369), .A(n9259), .ZN(P1_U3269) );
  XNOR2_X1 U10562 ( .A(n9260), .B(n9262), .ZN(n9437) );
  INV_X1 U10563 ( .A(n9437), .ZN(n9274) );
  AOI22_X1 U10564 ( .A1(n9380), .A2(n9299), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n4322), .ZN(n9261) );
  OAI21_X1 U10565 ( .B1(n9438), .B2(n9377), .A(n9261), .ZN(n9272) );
  XNOR2_X1 U10566 ( .A(n9263), .B(n9262), .ZN(n9264) );
  NAND2_X1 U10567 ( .A1(n9264), .A2(n9481), .ZN(n9443) );
  INV_X1 U10568 ( .A(n9265), .ZN(n9277) );
  AOI21_X1 U10569 ( .B1(n9441), .B2(n9277), .A(n9771), .ZN(n9267) );
  NAND2_X1 U10570 ( .A1(n9267), .A2(n9266), .ZN(n9442) );
  INV_X1 U10571 ( .A(n9442), .ZN(n9269) );
  AOI22_X1 U10572 ( .A1(n9269), .A2(n7703), .B1(n9722), .B2(n9268), .ZN(n9270)
         );
  AOI21_X1 U10573 ( .B1(n9443), .B2(n9270), .A(n4322), .ZN(n9271) );
  AOI211_X1 U10574 ( .C1(n9349), .C2(n9441), .A(n9272), .B(n9271), .ZN(n9273)
         );
  OAI21_X1 U10575 ( .B1(n9274), .B2(n9369), .A(n9273), .ZN(P1_U3270) );
  XNOR2_X1 U10576 ( .A(n9276), .B(n9281), .ZN(n9450) );
  AOI21_X1 U10577 ( .B1(n9446), .B2(n9291), .A(n9265), .ZN(n9447) );
  AOI22_X1 U10578 ( .A1(n4322), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9278), .B2(
        n9722), .ZN(n9279) );
  OAI21_X1 U10579 ( .B1(n9280), .B2(n9738), .A(n9279), .ZN(n9287) );
  XNOR2_X1 U10580 ( .A(n9282), .B(n9281), .ZN(n9285) );
  AOI222_X1 U10581 ( .A1(n9481), .A2(n9285), .B1(n9284), .B2(n9475), .C1(n9283), .C2(n9474), .ZN(n9449) );
  NOR2_X1 U10582 ( .A1(n9449), .A2(n4322), .ZN(n9286) );
  AOI211_X1 U10583 ( .C1(n9447), .C2(n9303), .A(n9287), .B(n9286), .ZN(n9288)
         );
  OAI21_X1 U10584 ( .B1(n9450), .B2(n9369), .A(n9288), .ZN(P1_U3271) );
  XNOR2_X1 U10585 ( .A(n9290), .B(n9296), .ZN(n9456) );
  INV_X1 U10586 ( .A(n9291), .ZN(n9292) );
  AOI21_X1 U10587 ( .B1(n9451), .B2(n9315), .A(n9292), .ZN(n9453) );
  AOI22_X1 U10588 ( .A1(n4322), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9293), .B2(
        n9722), .ZN(n9294) );
  OAI21_X1 U10589 ( .B1(n9295), .B2(n9738), .A(n9294), .ZN(n9302) );
  INV_X1 U10590 ( .A(n9296), .ZN(n9298) );
  OAI21_X1 U10591 ( .B1(n4363), .B2(n9298), .A(n9297), .ZN(n9300) );
  AOI222_X1 U10592 ( .A1(n9481), .A2(n9300), .B1(n9466), .B2(n9474), .C1(n9299), .C2(n9475), .ZN(n9455) );
  NOR2_X1 U10593 ( .A1(n9455), .A2(n4322), .ZN(n9301) );
  AOI211_X1 U10594 ( .C1(n9303), .C2(n9453), .A(n9302), .B(n9301), .ZN(n9304)
         );
  OAI21_X1 U10595 ( .B1(n9456), .B2(n9369), .A(n9304), .ZN(P1_U3272) );
  AOI21_X1 U10596 ( .B1(n9306), .B2(n9305), .A(n9523), .ZN(n9308) );
  NAND2_X1 U10597 ( .A1(n9308), .A2(n9307), .ZN(n9462) );
  XNOR2_X1 U10598 ( .A(n9309), .B(n9310), .ZN(n9457) );
  NAND2_X1 U10599 ( .A1(n9457), .A2(n9742), .ZN(n9320) );
  NAND2_X1 U10600 ( .A1(n9380), .A2(n9476), .ZN(n9314) );
  INV_X1 U10601 ( .A(n9311), .ZN(n9312) );
  AOI22_X1 U10602 ( .A1(n4322), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9312), .B2(
        n9722), .ZN(n9313) );
  OAI211_X1 U10603 ( .C1(n9458), .C2(n9377), .A(n9314), .B(n9313), .ZN(n9318)
         );
  OAI211_X1 U10604 ( .C1(n9316), .C2(n4405), .A(n9452), .B(n9315), .ZN(n9461)
         );
  NOR2_X1 U10605 ( .A1(n9461), .A2(n9735), .ZN(n9317) );
  AOI211_X1 U10606 ( .C1(n9349), .C2(n9460), .A(n9318), .B(n9317), .ZN(n9319)
         );
  OAI211_X1 U10607 ( .C1(n4322), .C2(n9462), .A(n9320), .B(n9319), .ZN(
        P1_U3273) );
  XOR2_X1 U10608 ( .A(n9321), .B(n9322), .Z(n9472) );
  XNOR2_X1 U10609 ( .A(n9323), .B(n9322), .ZN(n9470) );
  AOI211_X1 U10610 ( .C1(n9324), .C2(n9341), .A(n9771), .B(n4405), .ZN(n9469)
         );
  NAND2_X1 U10611 ( .A1(n9469), .A2(n9724), .ZN(n9331) );
  INV_X1 U10612 ( .A(n9325), .ZN(n9326) );
  AOI22_X1 U10613 ( .A1(n4322), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9326), .B2(
        n9722), .ZN(n9327) );
  OAI21_X1 U10614 ( .B1(n9377), .B2(n9328), .A(n9327), .ZN(n9329) );
  AOI21_X1 U10615 ( .B1(n9380), .B2(n9465), .A(n9329), .ZN(n9330) );
  OAI211_X1 U10616 ( .C1(n4623), .C2(n9738), .A(n9331), .B(n9330), .ZN(n9332)
         );
  AOI21_X1 U10617 ( .B1(n9470), .B2(n9353), .A(n9332), .ZN(n9333) );
  OAI21_X1 U10618 ( .B1(n9472), .B2(n9369), .A(n9333), .ZN(P1_U3274) );
  XNOR2_X1 U10619 ( .A(n9174), .B(n9336), .ZN(n9484) );
  INV_X1 U10620 ( .A(n9335), .ZN(n9338) );
  OAI21_X1 U10621 ( .B1(n9338), .B2(n9337), .A(n9336), .ZN(n9340) );
  NAND2_X1 U10622 ( .A1(n9340), .A2(n9339), .ZN(n9482) );
  OAI211_X1 U10623 ( .C1(n4404), .C2(n9479), .A(n9452), .B(n9341), .ZN(n9478)
         );
  INV_X1 U10624 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9343) );
  OAI22_X1 U10625 ( .A1(n9366), .A2(n9343), .B1(n9342), .B2(n9733), .ZN(n9344)
         );
  AOI21_X1 U10626 ( .B1(n9345), .B2(n9476), .A(n9344), .ZN(n9346) );
  OAI21_X1 U10627 ( .B1(n9491), .B2(n9347), .A(n9346), .ZN(n9348) );
  AOI21_X1 U10628 ( .B1(n9350), .B2(n9349), .A(n9348), .ZN(n9351) );
  OAI21_X1 U10629 ( .B1(n9478), .B2(n9735), .A(n9351), .ZN(n9352) );
  AOI21_X1 U10630 ( .B1(n9482), .B2(n9353), .A(n9352), .ZN(n9354) );
  OAI21_X1 U10631 ( .B1(n9484), .B2(n9369), .A(n9354), .ZN(P1_U3275) );
  XNOR2_X1 U10632 ( .A(n9355), .B(n9361), .ZN(n9489) );
  INV_X1 U10633 ( .A(n9373), .ZN(n9356) );
  AOI211_X1 U10634 ( .C1(n9487), .C2(n9356), .A(n9771), .B(n4404), .ZN(n9486)
         );
  NOR2_X1 U10635 ( .A1(n9357), .A2(n9738), .ZN(n9360) );
  OAI22_X1 U10636 ( .A1(n9366), .A2(n9981), .B1(n9358), .B2(n9733), .ZN(n9359)
         );
  AOI211_X1 U10637 ( .C1(n9486), .C2(n9724), .A(n9360), .B(n9359), .ZN(n9368)
         );
  OAI211_X1 U10638 ( .C1(n9362), .C2(n9361), .A(n9335), .B(n9481), .ZN(n9365)
         );
  AOI22_X1 U10639 ( .A1(n9475), .A2(n9465), .B1(n9363), .B2(n9474), .ZN(n9364)
         );
  NAND2_X1 U10640 ( .A1(n9365), .A2(n9364), .ZN(n9485) );
  NAND2_X1 U10641 ( .A1(n9485), .A2(n9366), .ZN(n9367) );
  OAI211_X1 U10642 ( .C1(n9489), .C2(n9369), .A(n9368), .B(n9367), .ZN(
        P1_U3276) );
  XOR2_X1 U10643 ( .A(n9372), .B(n9370), .Z(n9497) );
  AOI21_X1 U10644 ( .B1(n9372), .B2(n9371), .A(n4410), .ZN(n9490) );
  NAND2_X1 U10645 ( .A1(n9490), .A2(n9742), .ZN(n9385) );
  AOI211_X1 U10646 ( .C1(n9494), .C2(n9374), .A(n9771), .B(n9373), .ZN(n9492)
         );
  INV_X1 U10647 ( .A(n9494), .ZN(n9382) );
  AOI22_X1 U10648 ( .A1(n4322), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9375), .B2(
        n9722), .ZN(n9376) );
  OAI21_X1 U10649 ( .B1(n9377), .B2(n9491), .A(n9376), .ZN(n9378) );
  AOI21_X1 U10650 ( .B1(n9380), .B2(n9379), .A(n9378), .ZN(n9381) );
  OAI21_X1 U10651 ( .B1(n9382), .B2(n9738), .A(n9381), .ZN(n9383) );
  AOI21_X1 U10652 ( .B1(n9492), .B2(n9724), .A(n9383), .ZN(n9384) );
  OAI211_X1 U10653 ( .C1(n9497), .C2(n9386), .A(n9385), .B(n9384), .ZN(
        P1_U3277) );
  OAI211_X1 U10654 ( .C1(n9388), .C2(n9781), .A(n9387), .B(n9389), .ZN(n9542)
         );
  MUX2_X1 U10655 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9542), .S(n9799), .Z(
        P1_U3553) );
  OAI211_X1 U10656 ( .C1(n9391), .C2(n9781), .A(n9390), .B(n9389), .ZN(n9543)
         );
  MUX2_X1 U10657 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9543), .S(n9799), .Z(
        P1_U3552) );
  NAND2_X1 U10658 ( .A1(n9392), .A2(n9786), .ZN(n9400) );
  NAND2_X1 U10659 ( .A1(n9400), .A2(n9399), .ZN(n9544) );
  MUX2_X1 U10660 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9544), .S(n9799), .Z(
        P1_U3551) );
  INV_X1 U10661 ( .A(n9402), .ZN(n9405) );
  INV_X1 U10662 ( .A(n9403), .ZN(n9404) );
  MUX2_X1 U10663 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9545), .S(n9799), .Z(
        P1_U3550) );
  NAND2_X1 U10664 ( .A1(n9407), .A2(n9786), .ZN(n9413) );
  OAI22_X1 U10665 ( .A1(n9424), .A2(n9532), .B1(n9408), .B2(n9530), .ZN(n9410)
         );
  AOI211_X1 U10666 ( .C1(n9762), .C2(n9411), .A(n9410), .B(n9409), .ZN(n9412)
         );
  OAI211_X1 U10667 ( .C1(n9523), .C2(n9414), .A(n9413), .B(n9412), .ZN(n9546)
         );
  MUX2_X1 U10668 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9546), .S(n9799), .Z(
        P1_U3549) );
  AOI22_X1 U10669 ( .A1(n9416), .A2(n9475), .B1(n9474), .B2(n9415), .ZN(n9417)
         );
  OAI211_X1 U10670 ( .C1(n9419), .C2(n9781), .A(n9418), .B(n9417), .ZN(n9420)
         );
  AOI21_X1 U10671 ( .B1(n9421), .B2(n9481), .A(n9420), .ZN(n9422) );
  OAI21_X1 U10672 ( .B1(n9423), .B2(n9766), .A(n9422), .ZN(n9547) );
  MUX2_X1 U10673 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9547), .S(n9799), .Z(
        P1_U3548) );
  OAI22_X1 U10674 ( .A1(n9424), .A2(n9530), .B1(n9438), .B2(n9532), .ZN(n9426)
         );
  AOI211_X1 U10675 ( .C1(n9762), .C2(n9427), .A(n9426), .B(n9425), .ZN(n9430)
         );
  NAND2_X1 U10676 ( .A1(n9428), .A2(n9481), .ZN(n9429) );
  OAI211_X1 U10677 ( .C1(n9431), .C2(n9766), .A(n9430), .B(n9429), .ZN(n9548)
         );
  MUX2_X1 U10678 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9548), .S(n9799), .Z(
        P1_U3547) );
  AOI21_X1 U10679 ( .B1(n9762), .B2(n9433), .A(n9432), .ZN(n9434) );
  OAI211_X1 U10680 ( .C1(n9436), .C2(n9766), .A(n9435), .B(n9434), .ZN(n9549)
         );
  MUX2_X1 U10681 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9549), .S(n9799), .Z(
        P1_U3546) );
  NAND2_X1 U10682 ( .A1(n9437), .A2(n9786), .ZN(n9445) );
  OAI22_X1 U10683 ( .A1(n9439), .A2(n9532), .B1(n9438), .B2(n9530), .ZN(n9440)
         );
  AOI21_X1 U10684 ( .B1(n9441), .B2(n9762), .A(n9440), .ZN(n9444) );
  NAND4_X1 U10685 ( .A1(n9445), .A2(n9444), .A3(n9443), .A4(n9442), .ZN(n9550)
         );
  MUX2_X1 U10686 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9550), .S(n9799), .Z(
        P1_U3545) );
  AOI22_X1 U10687 ( .A1(n9447), .A2(n9452), .B1(n9762), .B2(n9446), .ZN(n9448)
         );
  OAI211_X1 U10688 ( .C1(n9450), .C2(n9766), .A(n9449), .B(n9448), .ZN(n9551)
         );
  MUX2_X1 U10689 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9551), .S(n9799), .Z(
        P1_U3544) );
  AOI22_X1 U10690 ( .A1(n9453), .A2(n9452), .B1(n9762), .B2(n9451), .ZN(n9454)
         );
  OAI211_X1 U10691 ( .C1(n9456), .C2(n9766), .A(n9455), .B(n9454), .ZN(n9552)
         );
  MUX2_X1 U10692 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9552), .S(n9799), .Z(
        P1_U3543) );
  NAND2_X1 U10693 ( .A1(n9457), .A2(n9786), .ZN(n9464) );
  OAI22_X1 U10694 ( .A1(n9458), .A2(n9530), .B1(n9177), .B2(n9532), .ZN(n9459)
         );
  AOI21_X1 U10695 ( .B1(n9460), .B2(n9762), .A(n9459), .ZN(n9463) );
  NAND4_X1 U10696 ( .A1(n9464), .A2(n9463), .A3(n9462), .A4(n9461), .ZN(n9553)
         );
  MUX2_X1 U10697 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9553), .S(n9799), .Z(
        P1_U3542) );
  AOI22_X1 U10698 ( .A1(n9466), .A2(n9475), .B1(n9474), .B2(n9465), .ZN(n9467)
         );
  OAI21_X1 U10699 ( .B1(n4623), .B2(n9781), .A(n9467), .ZN(n9468) );
  AOI211_X1 U10700 ( .C1(n9470), .C2(n9481), .A(n9469), .B(n9468), .ZN(n9471)
         );
  OAI21_X1 U10701 ( .B1(n9472), .B2(n9766), .A(n9471), .ZN(n9554) );
  MUX2_X1 U10702 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9554), .S(n9799), .Z(
        P1_U3541) );
  AOI22_X1 U10703 ( .A1(n9476), .A2(n9475), .B1(n9474), .B2(n9473), .ZN(n9477)
         );
  OAI211_X1 U10704 ( .C1(n9479), .C2(n9781), .A(n9478), .B(n9477), .ZN(n9480)
         );
  AOI21_X1 U10705 ( .B1(n9482), .B2(n9481), .A(n9480), .ZN(n9483) );
  OAI21_X1 U10706 ( .B1(n9484), .B2(n9766), .A(n9483), .ZN(n9555) );
  MUX2_X1 U10707 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9555), .S(n9799), .Z(
        P1_U3540) );
  AOI211_X1 U10708 ( .C1(n9762), .C2(n9487), .A(n9486), .B(n9485), .ZN(n9488)
         );
  OAI21_X1 U10709 ( .B1(n9489), .B2(n9766), .A(n9488), .ZN(n9556) );
  MUX2_X1 U10710 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9556), .S(n9799), .Z(
        P1_U3539) );
  NAND2_X1 U10711 ( .A1(n9490), .A2(n9786), .ZN(n9496) );
  OAI22_X1 U10712 ( .A1(n9491), .A2(n9530), .B1(n9507), .B2(n9532), .ZN(n9493)
         );
  AOI211_X1 U10713 ( .C1(n9762), .C2(n9494), .A(n9493), .B(n9492), .ZN(n9495)
         );
  OAI211_X1 U10714 ( .C1(n9523), .C2(n9497), .A(n9496), .B(n9495), .ZN(n9557)
         );
  MUX2_X1 U10715 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9557), .S(n9799), .Z(
        P1_U3538) );
  NAND2_X1 U10716 ( .A1(n9498), .A2(n9786), .ZN(n9504) );
  OAI22_X1 U10717 ( .A1(n9499), .A2(n9530), .B1(n9516), .B2(n9532), .ZN(n9501)
         );
  AOI211_X1 U10718 ( .C1(n9762), .C2(n9502), .A(n9501), .B(n9500), .ZN(n9503)
         );
  OAI211_X1 U10719 ( .C1(n9523), .C2(n9505), .A(n9504), .B(n9503), .ZN(n9558)
         );
  MUX2_X1 U10720 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9558), .S(n9799), .Z(
        P1_U3537) );
  NAND2_X1 U10721 ( .A1(n9506), .A2(n9786), .ZN(n9514) );
  OAI22_X1 U10722 ( .A1(n9508), .A2(n9532), .B1(n9507), .B2(n9530), .ZN(n9509)
         );
  AOI21_X1 U10723 ( .B1(n9510), .B2(n9762), .A(n9509), .ZN(n9513) );
  NAND4_X1 U10724 ( .A1(n9514), .A2(n9513), .A3(n9512), .A4(n9511), .ZN(n9559)
         );
  MUX2_X1 U10725 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9559), .S(n9799), .Z(
        P1_U3536) );
  NAND2_X1 U10726 ( .A1(n9515), .A2(n9786), .ZN(n9521) );
  OAI22_X1 U10727 ( .A1(n9531), .A2(n9532), .B1(n9516), .B2(n9530), .ZN(n9518)
         );
  AOI211_X1 U10728 ( .C1(n9762), .C2(n9519), .A(n9518), .B(n9517), .ZN(n9520)
         );
  OAI211_X1 U10729 ( .C1(n9523), .C2(n9522), .A(n9521), .B(n9520), .ZN(n9560)
         );
  MUX2_X1 U10730 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9560), .S(n9799), .Z(
        P1_U3535) );
  AOI211_X1 U10731 ( .C1(n9762), .C2(n9526), .A(n9525), .B(n9524), .ZN(n9527)
         );
  OAI21_X1 U10732 ( .B1(n9528), .B2(n9766), .A(n9527), .ZN(n9561) );
  MUX2_X1 U10733 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9561), .S(n9799), .Z(
        P1_U3534) );
  NAND2_X1 U10734 ( .A1(n9529), .A2(n9786), .ZN(n9539) );
  OAI22_X1 U10735 ( .A1(n9533), .A2(n9532), .B1(n9531), .B2(n9530), .ZN(n9534)
         );
  AOI21_X1 U10736 ( .B1(n9535), .B2(n9762), .A(n9534), .ZN(n9538) );
  NAND4_X1 U10737 ( .A1(n9539), .A2(n9538), .A3(n9537), .A4(n9536), .ZN(n9562)
         );
  MUX2_X1 U10738 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9562), .S(n9799), .Z(
        P1_U3533) );
  MUX2_X1 U10739 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9540), .S(n9799), .Z(
        P1_U3523) );
  MUX2_X1 U10740 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9541), .S(n9799), .Z(
        P1_U3522) );
  MUX2_X1 U10741 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9542), .S(n9789), .Z(
        P1_U3521) );
  MUX2_X1 U10742 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9543), .S(n9789), .Z(
        P1_U3520) );
  MUX2_X1 U10743 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9544), .S(n9789), .Z(
        P1_U3519) );
  MUX2_X1 U10744 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9546), .S(n9789), .Z(
        P1_U3517) );
  MUX2_X1 U10745 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9547), .S(n9789), .Z(
        P1_U3516) );
  MUX2_X1 U10746 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9548), .S(n9789), .Z(
        P1_U3515) );
  MUX2_X1 U10747 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9549), .S(n9789), .Z(
        P1_U3514) );
  MUX2_X1 U10748 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9550), .S(n9789), .Z(
        P1_U3513) );
  MUX2_X1 U10749 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9551), .S(n9789), .Z(
        P1_U3512) );
  MUX2_X1 U10750 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9552), .S(n9789), .Z(
        P1_U3511) );
  MUX2_X1 U10751 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9553), .S(n9789), .Z(
        P1_U3510) );
  MUX2_X1 U10752 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9554), .S(n9789), .Z(
        P1_U3509) );
  MUX2_X1 U10753 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9555), .S(n9789), .Z(
        P1_U3507) );
  MUX2_X1 U10754 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9556), .S(n9789), .Z(
        P1_U3504) );
  MUX2_X1 U10755 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9557), .S(n9789), .Z(
        P1_U3501) );
  MUX2_X1 U10756 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9558), .S(n9789), .Z(
        P1_U3498) );
  MUX2_X1 U10757 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9559), .S(n9789), .Z(
        P1_U3495) );
  MUX2_X1 U10758 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9560), .S(n9789), .Z(
        P1_U3492) );
  MUX2_X1 U10759 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9561), .S(n9789), .Z(
        P1_U3489) );
  MUX2_X1 U10760 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9562), .S(n9789), .Z(
        P1_U3486) );
  MUX2_X1 U10761 ( .A(n9563), .B(P1_D_REG_1__SCAN_IN), .S(n9745), .Z(P1_U3440)
         );
  INV_X1 U10762 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9564) );
  NAND3_X1 U10763 ( .A1(n9564), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9566) );
  OAI22_X1 U10764 ( .A1(n4995), .A2(n9566), .B1(n9565), .B2(n7522), .ZN(n9567)
         );
  AOI21_X1 U10765 ( .B1(n9569), .B2(n9568), .A(n9567), .ZN(n9570) );
  INV_X1 U10766 ( .A(n9570), .ZN(P1_U3324) );
  OAI222_X1 U10767 ( .A1(P1_U3086), .A2(n9572), .B1(n7708), .B2(n9571), .C1(
        n10018), .C2(n7522), .ZN(P1_U3326) );
  MUX2_X1 U10768 ( .A(n9574), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI211_X1 U10769 ( .C1(n9577), .C2(n9576), .A(n9575), .B(n9706), .ZN(n9582)
         );
  AOI211_X1 U10770 ( .C1(n9580), .C2(n9579), .A(n9578), .B(n9711), .ZN(n9581)
         );
  AOI211_X1 U10771 ( .C1(n9718), .C2(n9583), .A(n9582), .B(n9581), .ZN(n9585)
         );
  OAI211_X1 U10772 ( .C1(n9586), .C2(n9721), .A(n9585), .B(n9584), .ZN(
        P1_U3253) );
  INV_X1 U10773 ( .A(n9587), .ZN(n9591) );
  INV_X1 U10774 ( .A(n9588), .ZN(n9590) );
  AOI211_X1 U10775 ( .C1(n9591), .C2(n9590), .A(n9589), .B(n9706), .ZN(n9596)
         );
  AOI211_X1 U10776 ( .C1(n9594), .C2(n9593), .A(n9711), .B(n9592), .ZN(n9595)
         );
  AOI211_X1 U10777 ( .C1(n9718), .C2(n9597), .A(n9596), .B(n9595), .ZN(n9599)
         );
  OAI211_X1 U10778 ( .C1(n9721), .C2(n10006), .A(n9599), .B(n9598), .ZN(
        P1_U3250) );
  OAI21_X1 U10779 ( .B1(n9601), .B2(n9600), .A(n9696), .ZN(n9603) );
  NOR2_X1 U10780 ( .A1(n9603), .A2(n9602), .ZN(n9608) );
  AOI211_X1 U10781 ( .C1(n9606), .C2(n9605), .A(n9604), .B(n9711), .ZN(n9607)
         );
  AOI211_X1 U10782 ( .C1(n9718), .C2(n9609), .A(n9608), .B(n9607), .ZN(n9611)
         );
  OAI211_X1 U10783 ( .C1(n9721), .C2(n9612), .A(n9611), .B(n9610), .ZN(
        P1_U3251) );
  XNOR2_X1 U10784 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10785 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U10786 ( .B1(n9614), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9613), .ZN(
        n9615) );
  XOR2_X1 U10787 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9615), .Z(n9619) );
  AOI22_X1 U10788 ( .A1(n9616), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9617) );
  OAI21_X1 U10789 ( .B1(n9619), .B2(n9618), .A(n9617), .ZN(P1_U3243) );
  INV_X1 U10790 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9635) );
  AOI21_X1 U10791 ( .B1(n9622), .B2(n9621), .A(n9620), .ZN(n9623) );
  NAND2_X1 U10792 ( .A1(n9692), .A2(n9623), .ZN(n9629) );
  AOI21_X1 U10793 ( .B1(n9626), .B2(n9625), .A(n9624), .ZN(n9627) );
  NAND2_X1 U10794 ( .A1(n9696), .A2(n9627), .ZN(n9628) );
  OAI211_X1 U10795 ( .C1(n9700), .C2(n9630), .A(n9629), .B(n9628), .ZN(n9631)
         );
  INV_X1 U10796 ( .A(n9631), .ZN(n9634) );
  INV_X1 U10797 ( .A(n9632), .ZN(n9633) );
  OAI211_X1 U10798 ( .C1(n9635), .C2(n9721), .A(n9634), .B(n9633), .ZN(
        P1_U3254) );
  AOI211_X1 U10799 ( .C1(n9638), .C2(n9637), .A(n9636), .B(n9706), .ZN(n9643)
         );
  AOI211_X1 U10800 ( .C1(n9641), .C2(n9640), .A(n9639), .B(n9711), .ZN(n9642)
         );
  AOI211_X1 U10801 ( .C1(n9718), .C2(n9644), .A(n9643), .B(n9642), .ZN(n9646)
         );
  OAI211_X1 U10802 ( .C1(n9647), .C2(n9721), .A(n9646), .B(n9645), .ZN(
        P1_U3256) );
  AOI21_X1 U10803 ( .B1(n9650), .B2(n9649), .A(n9648), .ZN(n9651) );
  NAND2_X1 U10804 ( .A1(n9692), .A2(n9651), .ZN(n9657) );
  AOI21_X1 U10805 ( .B1(n9654), .B2(n9653), .A(n9652), .ZN(n9655) );
  NAND2_X1 U10806 ( .A1(n9696), .A2(n9655), .ZN(n9656) );
  OAI211_X1 U10807 ( .C1(n9700), .C2(n9658), .A(n9657), .B(n9656), .ZN(n9659)
         );
  INV_X1 U10808 ( .A(n9659), .ZN(n9661) );
  OAI211_X1 U10809 ( .C1(n9662), .C2(n9721), .A(n9661), .B(n9660), .ZN(
        P1_U3257) );
  AOI211_X1 U10810 ( .C1(n9665), .C2(n9664), .A(n9663), .B(n9706), .ZN(n9670)
         );
  AOI211_X1 U10811 ( .C1(n9668), .C2(n9667), .A(n9666), .B(n9711), .ZN(n9669)
         );
  AOI211_X1 U10812 ( .C1(n9718), .C2(n9671), .A(n9670), .B(n9669), .ZN(n9673)
         );
  OAI211_X1 U10813 ( .C1(n9674), .C2(n9721), .A(n9673), .B(n9672), .ZN(
        P1_U3258) );
  OAI21_X1 U10814 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9684) );
  NOR2_X1 U10815 ( .A1(n9700), .A2(n9678), .ZN(n9683) );
  AOI211_X1 U10816 ( .C1(n9681), .C2(n9680), .A(n9679), .B(n9711), .ZN(n9682)
         );
  AOI211_X1 U10817 ( .C1(n9696), .C2(n9684), .A(n9683), .B(n9682), .ZN(n9686)
         );
  OAI211_X1 U10818 ( .C1(n9687), .C2(n9721), .A(n9686), .B(n9685), .ZN(
        P1_U3259) );
  INV_X1 U10819 ( .A(n9688), .ZN(n9699) );
  XNOR2_X1 U10820 ( .A(n9690), .B(n9689), .ZN(n9691) );
  NAND2_X1 U10821 ( .A1(n9692), .A2(n9691), .ZN(n9698) );
  XNOR2_X1 U10822 ( .A(n9694), .B(n9693), .ZN(n9695) );
  NAND2_X1 U10823 ( .A1(n9696), .A2(n9695), .ZN(n9697) );
  OAI211_X1 U10824 ( .C1(n9700), .C2(n9699), .A(n9698), .B(n9697), .ZN(n9701)
         );
  INV_X1 U10825 ( .A(n9701), .ZN(n9703) );
  OAI211_X1 U10826 ( .C1(n9704), .C2(n9721), .A(n9703), .B(n9702), .ZN(
        P1_U3260) );
  INV_X1 U10827 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10077) );
  INV_X1 U10828 ( .A(n9705), .ZN(n9707) );
  AOI211_X1 U10829 ( .C1(n9709), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9716)
         );
  INV_X1 U10830 ( .A(n9710), .ZN(n9712) );
  AOI211_X1 U10831 ( .C1(n9714), .C2(n9713), .A(n9712), .B(n9711), .ZN(n9715)
         );
  AOI211_X1 U10832 ( .C1(n9718), .C2(n9717), .A(n9716), .B(n9715), .ZN(n9720)
         );
  OAI211_X1 U10833 ( .C1(n10077), .C2(n9721), .A(n9720), .B(n9719), .ZN(
        P1_U3261) );
  AOI22_X1 U10834 ( .A1(n4322), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n9723), .B2(
        n9722), .ZN(n9727) );
  NAND2_X1 U10835 ( .A1(n9725), .A2(n9724), .ZN(n9726) );
  OAI211_X1 U10836 ( .C1(n9738), .C2(n9728), .A(n9727), .B(n9726), .ZN(n9729)
         );
  AOI21_X1 U10837 ( .B1(n9730), .B2(n9742), .A(n9729), .ZN(n9731) );
  OAI21_X1 U10838 ( .B1(n4322), .B2(n9732), .A(n9731), .ZN(P1_U3288) );
  OAI22_X1 U10839 ( .A1(n9735), .A2(n9734), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9733), .ZN(n9736) );
  AOI21_X1 U10840 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n4322), .A(n9736), .ZN(
        n9737) );
  OAI21_X1 U10841 ( .B1(n9739), .B2(n9738), .A(n9737), .ZN(n9740) );
  AOI21_X1 U10842 ( .B1(n9742), .B2(n9741), .A(n9740), .ZN(n9743) );
  OAI21_X1 U10843 ( .B1(n4322), .B2(n9744), .A(n9743), .ZN(P1_U3290) );
  AND2_X1 U10844 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9745), .ZN(P1_U3294) );
  AND2_X1 U10845 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9745), .ZN(P1_U3295) );
  AND2_X1 U10846 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9745), .ZN(P1_U3296) );
  NOR2_X1 U10847 ( .A1(n9746), .A2(n9976), .ZN(P1_U3297) );
  AND2_X1 U10848 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9745), .ZN(P1_U3298) );
  AND2_X1 U10849 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9745), .ZN(P1_U3299) );
  AND2_X1 U10850 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9745), .ZN(P1_U3300) );
  AND2_X1 U10851 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9745), .ZN(P1_U3301) );
  AND2_X1 U10852 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9745), .ZN(P1_U3302) );
  AND2_X1 U10853 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9745), .ZN(P1_U3303) );
  INV_X1 U10854 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U10855 ( .A1(n9746), .A2(n10062), .ZN(P1_U3304) );
  AND2_X1 U10856 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9745), .ZN(P1_U3305) );
  AND2_X1 U10857 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9745), .ZN(P1_U3306) );
  AND2_X1 U10858 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9745), .ZN(P1_U3307) );
  AND2_X1 U10859 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9745), .ZN(P1_U3308) );
  NOR2_X1 U10860 ( .A1(n9746), .A2(n9975), .ZN(P1_U3309) );
  AND2_X1 U10861 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9745), .ZN(P1_U3310) );
  AND2_X1 U10862 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9745), .ZN(P1_U3311) );
  AND2_X1 U10863 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9745), .ZN(P1_U3312) );
  AND2_X1 U10864 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9745), .ZN(P1_U3313) );
  AND2_X1 U10865 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9745), .ZN(P1_U3314) );
  INV_X1 U10866 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10051) );
  NOR2_X1 U10867 ( .A1(n9746), .A2(n10051), .ZN(P1_U3315) );
  AND2_X1 U10868 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9745), .ZN(P1_U3316) );
  AND2_X1 U10869 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9745), .ZN(P1_U3317) );
  INV_X1 U10870 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U10871 ( .A1(n9746), .A2(n10049), .ZN(P1_U3318) );
  AND2_X1 U10872 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9745), .ZN(P1_U3319) );
  AND2_X1 U10873 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9745), .ZN(P1_U3320) );
  AND2_X1 U10874 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9745), .ZN(P1_U3321) );
  NOR2_X1 U10875 ( .A1(n9746), .A2(n9979), .ZN(P1_U3322) );
  NOR2_X1 U10876 ( .A1(n9746), .A2(n10019), .ZN(P1_U3323) );
  INV_X1 U10877 ( .A(n9747), .ZN(n9748) );
  OAI21_X1 U10878 ( .B1(n9749), .B2(n9781), .A(n9748), .ZN(n9750) );
  AOI211_X1 U10879 ( .C1(n9786), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9790)
         );
  INV_X1 U10880 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9753) );
  AOI22_X1 U10881 ( .A1(n9789), .A2(n9790), .B1(n9753), .B2(n9787), .ZN(
        P1_U3459) );
  OAI21_X1 U10882 ( .B1(n9755), .B2(n9781), .A(n9754), .ZN(n9757) );
  AOI211_X1 U10883 ( .C1(n9786), .C2(n9758), .A(n9757), .B(n9756), .ZN(n9791)
         );
  INV_X1 U10884 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9759) );
  AOI22_X1 U10885 ( .A1(n9789), .A2(n9791), .B1(n9759), .B2(n9787), .ZN(
        P1_U3465) );
  AOI21_X1 U10886 ( .B1(n9762), .B2(n9761), .A(n9760), .ZN(n9763) );
  OAI211_X1 U10887 ( .C1(n9766), .C2(n9765), .A(n9764), .B(n9763), .ZN(n9767)
         );
  INV_X1 U10888 ( .A(n9767), .ZN(n9793) );
  INV_X1 U10889 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9768) );
  AOI22_X1 U10890 ( .A1(n9789), .A2(n9793), .B1(n9768), .B2(n9787), .ZN(
        P1_U3471) );
  INV_X1 U10891 ( .A(n9769), .ZN(n9774) );
  OAI22_X1 U10892 ( .A1(n9772), .A2(n9771), .B1(n9770), .B2(n9781), .ZN(n9773)
         );
  AOI21_X1 U10893 ( .B1(n9775), .B2(n9774), .A(n9773), .ZN(n9776) );
  INV_X1 U10894 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U10895 ( .A1(n9789), .A2(n9795), .B1(n9778), .B2(n9787), .ZN(
        P1_U3477) );
  INV_X1 U10896 ( .A(n9779), .ZN(n9782) );
  OAI21_X1 U10897 ( .B1(n9782), .B2(n9781), .A(n9780), .ZN(n9784) );
  AOI211_X1 U10898 ( .C1(n9786), .C2(n9785), .A(n9784), .B(n9783), .ZN(n9798)
         );
  INV_X1 U10899 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9788) );
  AOI22_X1 U10900 ( .A1(n9789), .A2(n9798), .B1(n9788), .B2(n9787), .ZN(
        P1_U3480) );
  AOI22_X1 U10901 ( .A1(n9799), .A2(n9790), .B1(n6717), .B2(n9796), .ZN(
        P1_U3524) );
  AOI22_X1 U10902 ( .A1(n9799), .A2(n9791), .B1(n6715), .B2(n9796), .ZN(
        P1_U3526) );
  AOI22_X1 U10903 ( .A1(n9799), .A2(n9793), .B1(n9792), .B2(n9796), .ZN(
        P1_U3528) );
  INV_X1 U10904 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9794) );
  AOI22_X1 U10905 ( .A1(n9799), .A2(n9795), .B1(n9794), .B2(n9796), .ZN(
        P1_U3530) );
  INV_X1 U10906 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9797) );
  AOI22_X1 U10907 ( .A1(n9799), .A2(n9798), .B1(n9797), .B2(n9796), .ZN(
        P1_U3531) );
  INV_X1 U10908 ( .A(n9800), .ZN(n9801) );
  OAI211_X1 U10909 ( .C1(n9803), .C2(n9802), .A(n9801), .B(n9838), .ZN(n9812)
         );
  OAI21_X1 U10910 ( .B1(n9806), .B2(n9805), .A(n9804), .ZN(n9807) );
  AOI22_X1 U10911 ( .A1(n9840), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n9808), .B2(
        n9807), .ZN(n9811) );
  NAND2_X1 U10912 ( .A1(n9830), .A2(n9809), .ZN(n9810) );
  AND3_X1 U10913 ( .A1(n9812), .A2(n9811), .A3(n9810), .ZN(n9820) );
  INV_X1 U10914 ( .A(n9813), .ZN(n9818) );
  NOR2_X1 U10915 ( .A1(n9815), .A2(n9814), .ZN(n9817) );
  OAI21_X1 U10916 ( .B1(n9818), .B2(n9817), .A(n9816), .ZN(n9819) );
  OAI211_X1 U10917 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6788), .A(n9820), .B(
        n9819), .ZN(P2_U3184) );
  AOI21_X1 U10918 ( .B1(n5906), .B2(n9822), .A(n9821), .ZN(n9833) );
  AOI21_X1 U10919 ( .B1(n5907), .B2(n9824), .A(n9823), .ZN(n9826) );
  NOR2_X1 U10920 ( .A1(n9826), .A2(n9825), .ZN(n9827) );
  AOI211_X1 U10921 ( .C1(n9830), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9831)
         );
  OAI21_X1 U10922 ( .B1(n9833), .B2(n9832), .A(n9831), .ZN(n9834) );
  INV_X1 U10923 ( .A(n9834), .ZN(n9842) );
  OAI21_X1 U10924 ( .B1(n9837), .B2(n9836), .A(n9835), .ZN(n9839) );
  AOI22_X1 U10925 ( .A1(n9840), .A2(P2_ADDR_REG_7__SCAN_IN), .B1(n9839), .B2(
        n9838), .ZN(n9841) );
  NAND2_X1 U10926 ( .A1(n9842), .A2(n9841), .ZN(P2_U3189) );
  INV_X1 U10927 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9849) );
  INV_X1 U10928 ( .A(n9843), .ZN(n9847) );
  AOI21_X1 U10929 ( .B1(n9845), .B2(n9877), .A(n9844), .ZN(n9846) );
  AOI211_X1 U10930 ( .C1(n9900), .C2(n9848), .A(n9847), .B(n9846), .ZN(n9907)
         );
  AOI22_X1 U10931 ( .A1(n9906), .A2(n9849), .B1(n9907), .B2(n9905), .ZN(
        P2_U3390) );
  INV_X1 U10932 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9854) );
  OAI22_X1 U10933 ( .A1(n9851), .A2(n9893), .B1(n9850), .B2(n9894), .ZN(n9852)
         );
  NOR2_X1 U10934 ( .A1(n9853), .A2(n9852), .ZN(n9908) );
  AOI22_X1 U10935 ( .A1(n9906), .A2(n9854), .B1(n9908), .B2(n9905), .ZN(
        P2_U3393) );
  OAI22_X1 U10936 ( .A1(n9856), .A2(n9893), .B1(n9855), .B2(n9894), .ZN(n9857)
         );
  NOR2_X1 U10937 ( .A1(n9858), .A2(n9857), .ZN(n9909) );
  AOI22_X1 U10938 ( .A1(n9906), .A2(n5844), .B1(n9909), .B2(n9905), .ZN(
        P2_U3396) );
  INV_X1 U10939 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9864) );
  INV_X1 U10940 ( .A(n9859), .ZN(n9863) );
  OAI22_X1 U10941 ( .A1(n9861), .A2(n9877), .B1(n9860), .B2(n9894), .ZN(n9862)
         );
  NOR2_X1 U10942 ( .A1(n9863), .A2(n9862), .ZN(n9910) );
  AOI22_X1 U10943 ( .A1(n9906), .A2(n9864), .B1(n9910), .B2(n9905), .ZN(
        P2_U3399) );
  INV_X1 U10944 ( .A(n9865), .ZN(n9869) );
  OAI21_X1 U10945 ( .B1(n9867), .B2(n9894), .A(n9866), .ZN(n9868) );
  AOI21_X1 U10946 ( .B1(n9869), .B2(n6266), .A(n9868), .ZN(n9912) );
  AOI22_X1 U10947 ( .A1(n9906), .A2(n5870), .B1(n9912), .B2(n9905), .ZN(
        P2_U3402) );
  INV_X1 U10948 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9874) );
  NOR2_X1 U10949 ( .A1(n9870), .A2(n9894), .ZN(n9872) );
  AOI211_X1 U10950 ( .C1(n6266), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9913)
         );
  AOI22_X1 U10951 ( .A1(n9906), .A2(n9874), .B1(n9913), .B2(n9905), .ZN(
        P2_U3405) );
  INV_X1 U10952 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9881) );
  INV_X1 U10953 ( .A(n9875), .ZN(n9880) );
  OAI22_X1 U10954 ( .A1(n9878), .A2(n9877), .B1(n9876), .B2(n9894), .ZN(n9879)
         );
  NOR2_X1 U10955 ( .A1(n9880), .A2(n9879), .ZN(n9914) );
  AOI22_X1 U10956 ( .A1(n9906), .A2(n9881), .B1(n9914), .B2(n9905), .ZN(
        P2_U3408) );
  INV_X1 U10957 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9886) );
  OAI22_X1 U10958 ( .A1(n9883), .A2(n9893), .B1(n9882), .B2(n9894), .ZN(n9884)
         );
  NOR2_X1 U10959 ( .A1(n9885), .A2(n9884), .ZN(n9915) );
  AOI22_X1 U10960 ( .A1(n9906), .A2(n9886), .B1(n9915), .B2(n9905), .ZN(
        P2_U3411) );
  INV_X1 U10961 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9892) );
  AND2_X1 U10962 ( .A1(n9887), .A2(n6266), .ZN(n9891) );
  NOR2_X1 U10963 ( .A1(n9888), .A2(n9894), .ZN(n9889) );
  NOR3_X1 U10964 ( .A1(n9891), .A2(n9890), .A3(n9889), .ZN(n9916) );
  AOI22_X1 U10965 ( .A1(n9906), .A2(n9892), .B1(n9916), .B2(n9905), .ZN(
        P2_U3414) );
  INV_X1 U10966 ( .A(n9893), .ZN(n9901) );
  NOR2_X1 U10967 ( .A1(n9895), .A2(n9894), .ZN(n9897) );
  AOI211_X1 U10968 ( .C1(n9898), .C2(n9901), .A(n9897), .B(n9896), .ZN(n9917)
         );
  AOI22_X1 U10969 ( .A1(n9906), .A2(n5942), .B1(n9917), .B2(n9905), .ZN(
        P2_U3417) );
  AOI22_X1 U10970 ( .A1(n9902), .A2(n9901), .B1(n9900), .B2(n9899), .ZN(n9903)
         );
  AND2_X1 U10971 ( .A1(n9904), .A2(n9903), .ZN(n9919) );
  AOI22_X1 U10972 ( .A1(n9906), .A2(n5958), .B1(n9919), .B2(n9905), .ZN(
        P2_U3420) );
  AOI22_X1 U10973 ( .A1(n9920), .A2(n9907), .B1(n5835), .B2(n9918), .ZN(
        P2_U3459) );
  AOI22_X1 U10974 ( .A1(n9920), .A2(n9908), .B1(n5822), .B2(n9918), .ZN(
        P2_U3460) );
  AOI22_X1 U10975 ( .A1(n9920), .A2(n9909), .B1(n5843), .B2(n9918), .ZN(
        P2_U3461) );
  AOI22_X1 U10976 ( .A1(n9920), .A2(n9910), .B1(n6359), .B2(n9918), .ZN(
        P2_U3462) );
  INV_X1 U10977 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9911) );
  AOI22_X1 U10978 ( .A1(n9920), .A2(n9912), .B1(n9911), .B2(n9918), .ZN(
        P2_U3463) );
  AOI22_X1 U10979 ( .A1(n9920), .A2(n9913), .B1(n5881), .B2(n9918), .ZN(
        P2_U3464) );
  AOI22_X1 U10980 ( .A1(n9920), .A2(n9914), .B1(n6357), .B2(n9918), .ZN(
        P2_U3465) );
  AOI22_X1 U10981 ( .A1(n9920), .A2(n9915), .B1(n5907), .B2(n9918), .ZN(
        P2_U3466) );
  AOI22_X1 U10982 ( .A1(n9920), .A2(n9916), .B1(n5923), .B2(n9918), .ZN(
        P2_U3467) );
  AOI22_X1 U10983 ( .A1(n9920), .A2(n9917), .B1(n5939), .B2(n9918), .ZN(
        P2_U3468) );
  AOI22_X1 U10984 ( .A1(n9920), .A2(n9919), .B1(n6290), .B2(n9918), .ZN(
        P2_U3469) );
  INV_X1 U10985 ( .A(n9921), .ZN(n9922) );
  NAND2_X1 U10986 ( .A1(n9923), .A2(n9922), .ZN(n9924) );
  XOR2_X1 U10987 ( .A(n9925), .B(n9924), .Z(ADD_1068_U5) );
  XOR2_X1 U10988 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U10989 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9927), .A(n9926), .ZN(
        n9929) );
  XOR2_X1 U10990 ( .A(n9929), .B(n9928), .Z(ADD_1068_U55) );
  XNOR2_X1 U10991 ( .A(n9931), .B(n9930), .ZN(ADD_1068_U56) );
  XNOR2_X1 U10992 ( .A(n9933), .B(n9932), .ZN(ADD_1068_U57) );
  XNOR2_X1 U10993 ( .A(n9935), .B(n9934), .ZN(ADD_1068_U58) );
  XNOR2_X1 U10994 ( .A(n9937), .B(n9936), .ZN(ADD_1068_U59) );
  XNOR2_X1 U10995 ( .A(n9939), .B(n9938), .ZN(ADD_1068_U60) );
  XNOR2_X1 U10996 ( .A(n9941), .B(n9940), .ZN(ADD_1068_U61) );
  XOR2_X1 U10997 ( .A(n9943), .B(n9942), .Z(ADD_1068_U62) );
  XOR2_X1 U10998 ( .A(n9945), .B(n9944), .Z(ADD_1068_U63) );
  NAND2_X1 U10999 ( .A1(n9946), .A2(P2_D_REG_4__SCAN_IN), .ZN(n10098) );
  NAND2_X1 U11000 ( .A1(keyinput54), .A2(keyinput8), .ZN(n9953) );
  NOR2_X1 U11001 ( .A1(keyinput61), .A2(keyinput27), .ZN(n9951) );
  NAND3_X1 U11002 ( .A1(keyinput46), .A2(keyinput53), .A3(keyinput0), .ZN(
        n9949) );
  INV_X1 U11003 ( .A(keyinput47), .ZN(n9947) );
  NAND3_X1 U11004 ( .A1(keyinput2), .A2(keyinput10), .A3(n9947), .ZN(n9948) );
  NOR4_X1 U11005 ( .A1(keyinput23), .A2(keyinput45), .A3(n9949), .A4(n9948), 
        .ZN(n9950) );
  NAND4_X1 U11006 ( .A1(keyinput35), .A2(keyinput22), .A3(n9951), .A4(n9950), 
        .ZN(n9952) );
  NOR4_X1 U11007 ( .A1(keyinput59), .A2(keyinput21), .A3(n9953), .A4(n9952), 
        .ZN(n10096) );
  NAND3_X1 U11008 ( .A1(keyinput19), .A2(keyinput48), .A3(keyinput26), .ZN(
        n9973) );
  NOR2_X1 U11009 ( .A1(keyinput57), .A2(keyinput60), .ZN(n9957) );
  NAND4_X1 U11010 ( .A1(keyinput29), .A2(keyinput4), .A3(keyinput52), .A4(
        keyinput14), .ZN(n9955) );
  NAND2_X1 U11011 ( .A1(keyinput43), .A2(keyinput28), .ZN(n9954) );
  NOR4_X1 U11012 ( .A1(keyinput34), .A2(keyinput1), .A3(n9955), .A4(n9954), 
        .ZN(n9956) );
  NAND4_X1 U11013 ( .A1(keyinput63), .A2(keyinput40), .A3(n9957), .A4(n9956), 
        .ZN(n9972) );
  NOR3_X1 U11014 ( .A1(keyinput33), .A2(keyinput38), .A3(keyinput37), .ZN(
        n9970) );
  NAND3_X1 U11015 ( .A1(keyinput20), .A2(keyinput3), .A3(keyinput15), .ZN(
        n9961) );
  NOR4_X1 U11016 ( .A1(keyinput16), .A2(keyinput55), .A3(keyinput42), .A4(
        keyinput30), .ZN(n9959) );
  NOR2_X1 U11017 ( .A1(keyinput17), .A2(keyinput44), .ZN(n9958) );
  NAND4_X1 U11018 ( .A1(n9959), .A2(keyinput6), .A3(keyinput5), .A4(n9958), 
        .ZN(n9960) );
  NOR3_X1 U11019 ( .A1(keyinput39), .A2(n9961), .A3(n9960), .ZN(n9969) );
  NOR2_X1 U11020 ( .A1(keyinput13), .A2(keyinput51), .ZN(n9962) );
  NAND3_X1 U11021 ( .A1(keyinput32), .A2(keyinput7), .A3(n9962), .ZN(n9967) );
  NAND3_X1 U11022 ( .A1(keyinput41), .A2(keyinput12), .A3(keyinput9), .ZN(
        n9966) );
  NOR4_X1 U11023 ( .A1(keyinput49), .A2(keyinput56), .A3(keyinput25), .A4(
        keyinput24), .ZN(n9964) );
  NOR2_X1 U11024 ( .A1(keyinput36), .A2(keyinput50), .ZN(n9963) );
  NAND4_X1 U11025 ( .A1(n9964), .A2(keyinput62), .A3(keyinput31), .A4(n9963), 
        .ZN(n9965) );
  NOR4_X1 U11026 ( .A1(keyinput58), .A2(n9967), .A3(n9966), .A4(n9965), .ZN(
        n9968) );
  NAND4_X1 U11027 ( .A1(keyinput11), .A2(n9970), .A3(n9969), .A4(n9968), .ZN(
        n9971) );
  NOR4_X1 U11028 ( .A1(keyinput18), .A2(n9973), .A3(n9972), .A4(n9971), .ZN(
        n10095) );
  AOI22_X1 U11029 ( .A1(n9976), .A2(keyinput46), .B1(keyinput23), .B2(n9975), 
        .ZN(n9974) );
  OAI221_X1 U11030 ( .B1(n9976), .B2(keyinput46), .C1(n9975), .C2(keyinput23), 
        .A(n9974), .ZN(n9988) );
  INV_X1 U11031 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U11032 ( .A1(n9979), .A2(keyinput21), .B1(keyinput8), .B2(n9978), 
        .ZN(n9977) );
  OAI221_X1 U11033 ( .B1(n9979), .B2(keyinput21), .C1(n9978), .C2(keyinput8), 
        .A(n9977), .ZN(n9987) );
  AOI22_X1 U11034 ( .A1(n9982), .A2(keyinput54), .B1(keyinput59), .B2(n9981), 
        .ZN(n9980) );
  OAI221_X1 U11035 ( .B1(n9982), .B2(keyinput54), .C1(n9981), .C2(keyinput59), 
        .A(n9980), .ZN(n9986) );
  XNOR2_X1 U11036 ( .A(P1_REG0_REG_22__SCAN_IN), .B(keyinput0), .ZN(n9984) );
  XNOR2_X1 U11037 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput53), .ZN(n9983) );
  NAND2_X1 U11038 ( .A1(n9984), .A2(n9983), .ZN(n9985) );
  NOR4_X1 U11039 ( .A1(n9988), .A2(n9987), .A3(n9986), .A4(n9985), .ZN(n10031)
         );
  AOI22_X1 U11040 ( .A1(n9991), .A2(keyinput2), .B1(keyinput45), .B2(n9990), 
        .ZN(n9989) );
  OAI221_X1 U11041 ( .B1(n9991), .B2(keyinput2), .C1(n9990), .C2(keyinput45), 
        .A(n9989), .ZN(n10003) );
  INV_X1 U11042 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U11043 ( .A1(n9994), .A2(keyinput35), .B1(keyinput61), .B2(n9993), 
        .ZN(n9992) );
  OAI221_X1 U11044 ( .B1(n9994), .B2(keyinput35), .C1(n9993), .C2(keyinput61), 
        .A(n9992), .ZN(n10002) );
  INV_X1 U11045 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9996) );
  AOI22_X1 U11046 ( .A1(n9997), .A2(keyinput47), .B1(keyinput10), .B2(n9996), 
        .ZN(n9995) );
  OAI221_X1 U11047 ( .B1(n9997), .B2(keyinput47), .C1(n9996), .C2(keyinput10), 
        .A(n9995), .ZN(n10001) );
  XNOR2_X1 U11048 ( .A(P2_REG0_REG_20__SCAN_IN), .B(keyinput22), .ZN(n9999) );
  XNOR2_X1 U11049 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput27), .ZN(n9998) );
  NAND2_X1 U11050 ( .A1(n9999), .A2(n9998), .ZN(n10000) );
  NOR4_X1 U11051 ( .A1(n10003), .A2(n10002), .A3(n10001), .A4(n10000), .ZN(
        n10030) );
  INV_X1 U11052 ( .A(SI_29_), .ZN(n10005) );
  AOI22_X1 U11053 ( .A1(n10006), .A2(keyinput3), .B1(n10005), .B2(keyinput15), 
        .ZN(n10004) );
  OAI221_X1 U11054 ( .B1(n10006), .B2(keyinput3), .C1(n10005), .C2(keyinput15), 
        .A(n10004), .ZN(n10016) );
  XNOR2_X1 U11055 ( .A(n10007), .B(keyinput33), .ZN(n10015) );
  XNOR2_X1 U11056 ( .A(n10008), .B(keyinput37), .ZN(n10014) );
  XNOR2_X1 U11057 ( .A(P2_IR_REG_30__SCAN_IN), .B(keyinput38), .ZN(n10012) );
  XNOR2_X1 U11058 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput11), .ZN(n10011) );
  XNOR2_X1 U11059 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput20), .ZN(n10010) );
  XNOR2_X1 U11060 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput39), .ZN(n10009) );
  NAND4_X1 U11061 ( .A1(n10012), .A2(n10011), .A3(n10010), .A4(n10009), .ZN(
        n10013) );
  NOR4_X1 U11062 ( .A1(n10016), .A2(n10015), .A3(n10014), .A4(n10013), .ZN(
        n10029) );
  AOI22_X1 U11063 ( .A1(n10019), .A2(keyinput16), .B1(n10018), .B2(keyinput55), 
        .ZN(n10017) );
  OAI221_X1 U11064 ( .B1(n10019), .B2(keyinput16), .C1(n10018), .C2(keyinput55), .A(n10017), .ZN(n10027) );
  XOR2_X1 U11065 ( .A(P1_REG0_REG_14__SCAN_IN), .B(keyinput5), .Z(n10026) );
  XNOR2_X1 U11066 ( .A(n4609), .B(keyinput44), .ZN(n10025) );
  XNOR2_X1 U11067 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput42), .ZN(n10023) );
  XNOR2_X1 U11068 ( .A(P1_REG0_REG_31__SCAN_IN), .B(keyinput30), .ZN(n10022)
         );
  XNOR2_X1 U11069 ( .A(P2_REG1_REG_16__SCAN_IN), .B(keyinput17), .ZN(n10021)
         );
  NAND4_X1 U11070 ( .A1(n10023), .A2(n10022), .A3(n10021), .A4(n10020), .ZN(
        n10024) );
  NOR4_X1 U11071 ( .A1(n10027), .A2(n10026), .A3(n10025), .A4(n10024), .ZN(
        n10028) );
  NAND4_X1 U11072 ( .A1(n10031), .A2(n10030), .A3(n10029), .A4(n10028), .ZN(
        n10094) );
  AOI22_X1 U11073 ( .A1(n10034), .A2(keyinput34), .B1(keyinput28), .B2(n10033), 
        .ZN(n10032) );
  OAI221_X1 U11074 ( .B1(n10034), .B2(keyinput34), .C1(n10033), .C2(keyinput28), .A(n10032), .ZN(n10046) );
  INV_X1 U11075 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10036) );
  AOI22_X1 U11076 ( .A1(n6359), .A2(keyinput1), .B1(keyinput43), .B2(n10036), 
        .ZN(n10035) );
  OAI221_X1 U11077 ( .B1(n6359), .B2(keyinput1), .C1(n10036), .C2(keyinput43), 
        .A(n10035), .ZN(n10045) );
  AOI22_X1 U11078 ( .A1(n10039), .A2(keyinput48), .B1(n10038), .B2(keyinput26), 
        .ZN(n10037) );
  OAI221_X1 U11079 ( .B1(n10039), .B2(keyinput48), .C1(n10038), .C2(keyinput26), .A(n10037), .ZN(n10044) );
  INV_X1 U11080 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10042) );
  AOI22_X1 U11081 ( .A1(n10042), .A2(keyinput19), .B1(keyinput18), .B2(n10041), 
        .ZN(n10040) );
  OAI221_X1 U11082 ( .B1(n10042), .B2(keyinput19), .C1(n10041), .C2(keyinput18), .A(n10040), .ZN(n10043) );
  NOR4_X1 U11083 ( .A1(n10046), .A2(n10045), .A3(n10044), .A4(n10043), .ZN(
        n10092) );
  AOI22_X1 U11084 ( .A1(n10049), .A2(keyinput52), .B1(n10048), .B2(keyinput14), 
        .ZN(n10047) );
  OAI221_X1 U11085 ( .B1(n10049), .B2(keyinput52), .C1(n10048), .C2(keyinput14), .A(n10047), .ZN(n10060) );
  AOI22_X1 U11086 ( .A1(n10051), .A2(keyinput40), .B1(keyinput60), .B2(n5511), 
        .ZN(n10050) );
  OAI221_X1 U11087 ( .B1(n10051), .B2(keyinput40), .C1(n5511), .C2(keyinput60), 
        .A(n10050), .ZN(n10059) );
  INV_X1 U11088 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10054) );
  INV_X1 U11089 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10053) );
  AOI22_X1 U11090 ( .A1(n10054), .A2(keyinput29), .B1(n10053), .B2(keyinput4), 
        .ZN(n10052) );
  OAI221_X1 U11091 ( .B1(n10054), .B2(keyinput29), .C1(n10053), .C2(keyinput4), 
        .A(n10052), .ZN(n10058) );
  XOR2_X1 U11092 ( .A(n7711), .B(keyinput63), .Z(n10056) );
  XNOR2_X1 U11093 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput57), .ZN(n10055) );
  NAND2_X1 U11094 ( .A1(n10056), .A2(n10055), .ZN(n10057) );
  NOR4_X1 U11095 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n10091) );
  INV_X1 U11096 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10063) );
  AOI22_X1 U11097 ( .A1(n10063), .A2(keyinput25), .B1(n10062), .B2(keyinput24), 
        .ZN(n10061) );
  OAI221_X1 U11098 ( .B1(n10063), .B2(keyinput25), .C1(n10062), .C2(keyinput24), .A(n10061), .ZN(n10075) );
  INV_X1 U11099 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n10065) );
  AOI22_X1 U11100 ( .A1(n10066), .A2(keyinput49), .B1(keyinput56), .B2(n10065), 
        .ZN(n10064) );
  OAI221_X1 U11101 ( .B1(n10066), .B2(keyinput49), .C1(n10065), .C2(keyinput56), .A(n10064), .ZN(n10074) );
  AOI22_X1 U11102 ( .A1(n10069), .A2(keyinput36), .B1(n10068), .B2(keyinput50), 
        .ZN(n10067) );
  OAI221_X1 U11103 ( .B1(n10069), .B2(keyinput36), .C1(n10068), .C2(keyinput50), .A(n10067), .ZN(n10073) );
  AOI22_X1 U11104 ( .A1(n10071), .A2(keyinput62), .B1(keyinput31), .B2(n6290), 
        .ZN(n10070) );
  OAI221_X1 U11105 ( .B1(n10071), .B2(keyinput62), .C1(n6290), .C2(keyinput31), 
        .A(n10070), .ZN(n10072) );
  NOR4_X1 U11106 ( .A1(n10075), .A2(n10074), .A3(n10073), .A4(n10072), .ZN(
        n10090) );
  AOI22_X1 U11107 ( .A1(n10078), .A2(keyinput58), .B1(keyinput41), .B2(n10077), 
        .ZN(n10076) );
  OAI221_X1 U11108 ( .B1(n10078), .B2(keyinput58), .C1(n10077), .C2(keyinput41), .A(n10076), .ZN(n10088) );
  AOI22_X1 U11109 ( .A1(n10081), .A2(keyinput7), .B1(keyinput32), .B2(n10080), 
        .ZN(n10079) );
  OAI221_X1 U11110 ( .B1(n10081), .B2(keyinput7), .C1(n10080), .C2(keyinput32), 
        .A(n10079), .ZN(n10087) );
  XNOR2_X1 U11111 ( .A(SI_0_), .B(keyinput13), .ZN(n10085) );
  XNOR2_X1 U11112 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput51), .ZN(n10084) );
  XNOR2_X1 U11113 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput9), .ZN(n10083) );
  XNOR2_X1 U11114 ( .A(SI_13_), .B(keyinput12), .ZN(n10082) );
  NAND4_X1 U11115 ( .A1(n10085), .A2(n10084), .A3(n10083), .A4(n10082), .ZN(
        n10086) );
  NOR3_X1 U11116 ( .A1(n10088), .A2(n10087), .A3(n10086), .ZN(n10089) );
  NAND4_X1 U11117 ( .A1(n10092), .A2(n10091), .A3(n10090), .A4(n10089), .ZN(
        n10093) );
  AOI211_X1 U11118 ( .C1(n10096), .C2(n10095), .A(n10094), .B(n10093), .ZN(
        n10097) );
  XNOR2_X1 U11119 ( .A(n10098), .B(n10097), .ZN(P2_U3261) );
  XOR2_X1 U11120 ( .A(n10099), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1068_U50) );
  NOR2_X1 U11121 ( .A1(n10101), .A2(n10100), .ZN(n10102) );
  XOR2_X1 U11122 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10102), .Z(ADD_1068_U51) );
  INV_X1 U11123 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10103) );
  XNOR2_X1 U11124 ( .A(n10104), .B(n10103), .ZN(ADD_1068_U47) );
  XOR2_X1 U11125 ( .A(n10105), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1068_U49) );
  XOR2_X1 U11126 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10106), .Z(ADD_1068_U48) );
  XOR2_X1 U11127 ( .A(n10108), .B(n10107), .Z(ADD_1068_U54) );
  XOR2_X1 U11128 ( .A(n10110), .B(n10109), .Z(ADD_1068_U53) );
  XNOR2_X1 U11129 ( .A(n10112), .B(n10111), .ZN(ADD_1068_U52) );
  BUF_X1 U4826 ( .A(n5562), .Z(n4316) );
  CLKBUF_X1 U4825 ( .A(n5562), .Z(n4317) );
  INV_X1 U4820 ( .A(n6060), .ZN(n5938) );
  CLKBUF_X1 U4835 ( .A(n5658), .Z(n4324) );
  INV_X1 U4866 ( .A(n6859), .ZN(n4859) );
endmodule

