

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, 
        READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, 
        M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, 
        STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, 
        W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N,
         BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
         CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
         REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
         FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276;

  CLKBUF_X2 U3457 ( .A(n3866), .Z(n3833) );
  BUF_X2 U3458 ( .A(n3860), .Z(n3825) );
  CLKBUF_X2 U34590 ( .A(n3834), .Z(n3835) );
  NOR2_X1 U34600 ( .A1(n3439), .A2(n3798), .ZN(n4713) );
  AND2_X1 U34610 ( .A1(n3716), .A2(n3752), .ZN(n3809) );
  CLKBUF_X2 U34620 ( .A(n3785), .Z(n4354) );
  NAND3_X2 U34630 ( .A1(n3778), .A2(n3777), .A3(n3776), .ZN(n5169) );
  AND4_X1 U34640 ( .A1(n3738), .A2(n3737), .A3(n3736), .A4(n3735), .ZN(n3745)
         );
  NAND4_X1 U34650 ( .A1(n3667), .A2(n3666), .A3(n3665), .A4(n3664), .ZN(n3848)
         );
  AND4_X2 U3466 ( .A1(n3714), .A2(n3713), .A3(n3712), .A4(n3711), .ZN(n3750)
         );
  AND4_X1 U3467 ( .A1(n3702), .A2(n3701), .A3(n3700), .A4(n3699), .ZN(n3713)
         );
  AND4_X1 U34680 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3711)
         );
  AND2_X1 U34690 ( .A1(n6555), .A2(n4917), .ZN(n3866) );
  AND2_X2 U34700 ( .A1(n3549), .A2(n4949), .ZN(n3442) );
  AND2_X2 U34710 ( .A1(n4934), .A2(n4949), .ZN(n3761) );
  INV_X2 U34720 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4927) );
  OR2_X1 U34730 ( .A1(n4418), .A2(n7067), .ZN(n3448) );
  CLKBUF_X2 U34740 ( .A(n3442), .Z(n4273) );
  NOR3_X1 U3475 ( .A1(n4531), .A2(n5169), .A3(n3795), .ZN(n3814) );
  AND2_X1 U3476 ( .A1(n4680), .A2(n3854), .ZN(n3435) );
  AOI21_X1 U3477 ( .B1(n3797), .B2(n3448), .A(n3435), .ZN(n3800) );
  AND2_X1 U3478 ( .A1(n3796), .A2(n3814), .ZN(n4680) );
  INV_X1 U3479 ( .A(n4490), .ZN(n4705) );
  CLKBUF_X2 U3480 ( .A(n4405), .Z(n4490) );
  OAI21_X1 U3481 ( .B1(n3890), .B2(n3489), .A(n3432), .ZN(n3920) );
  AND4_X1 U3482 ( .A1(n3706), .A2(n3705), .A3(n3704), .A4(n3703), .ZN(n3712)
         );
  NOR2_X1 U3483 ( .A1(n4822), .A2(n4823), .ZN(n3918) );
  AND4_X1 U3484 ( .A1(n3743), .A2(n3742), .A3(n3741), .A4(n3740), .ZN(n3744)
         );
  NAND2_X1 U3485 ( .A1(n3785), .A2(n4871), .ZN(n4627) );
  INV_X2 U3486 ( .A(n5843), .ZN(n4833) );
  XNOR2_X1 U3488 ( .A(n6137), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5611)
         );
  OAI21_X1 U3489 ( .B1(n5379), .B2(n5380), .A(n4560), .ZN(n4902) );
  INV_X1 U3490 ( .A(n5169), .ZN(n4855) );
  NOR2_X4 U3492 ( .A1(n5776), .A2(n3523), .ZN(n5971) );
  OAI21_X2 U3493 ( .B1(n6087), .B2(n4690), .A(n4689), .ZN(n5783) );
  AOI211_X2 U3494 ( .C1(n6146), .C2(n6147), .A(n6117), .B(n6145), .ZN(n6139)
         );
  NOR2_X2 U3495 ( .A1(n6161), .A2(n6115), .ZN(n6146) );
  AND2_X1 U3496 ( .A1(n5714), .A2(n3466), .ZN(n5774) );
  CLKBUF_X1 U3497 ( .A(n5562), .Z(n5619) );
  INV_X1 U3499 ( .A(n4614), .ZN(n6089) );
  OR2_X1 U3500 ( .A1(n4593), .A2(n4592), .ZN(n4614) );
  BUF_X1 U3501 ( .A(n4883), .Z(n3445) );
  NAND2_X1 U3502 ( .A1(n3939), .A2(n3938), .ZN(n4849) );
  BUF_X1 U3503 ( .A(n4842), .Z(n3444) );
  XNOR2_X1 U3504 ( .A(n4921), .B(n4919), .ZN(n4842) );
  OR2_X1 U3507 ( .A1(n4406), .A2(n4863), .ZN(n3813) );
  AND3_X1 U3508 ( .A1(n3848), .A2(n5169), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n4389) );
  AND4_X1 U3509 ( .A1(n3733), .A2(n3732), .A3(n3731), .A4(n3730), .ZN(n3746)
         );
  BUF_X2 U3510 ( .A(n3762), .Z(n4648) );
  CLKBUF_X2 U3511 ( .A(n3865), .Z(n3832) );
  CLKBUF_X2 U3512 ( .A(n3739), .Z(n4649) );
  BUF_X2 U3513 ( .A(n3767), .Z(n4177) );
  CLKBUF_X2 U3514 ( .A(n3768), .Z(n3557) );
  INV_X1 U3515 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3921) );
  AND2_X1 U3516 ( .A1(n3495), .A2(n3493), .ZN(n6104) );
  AND2_X1 U3517 ( .A1(n3423), .A2(n3424), .ZN(n6097) );
  OAI21_X1 U3518 ( .B1(n5842), .B2(n6961), .A(n3485), .ZN(n3484) );
  AOI21_X1 U3519 ( .B1(n4345), .B2(n4344), .A(n4703), .ZN(n4636) );
  XNOR2_X1 U3520 ( .A(n4671), .B(n4670), .ZN(n5850) );
  CLKBUF_X1 U3521 ( .A(n5897), .Z(n5898) );
  NAND2_X1 U3522 ( .A1(n5910), .A2(n5911), .ZN(n5897) );
  NAND2_X1 U3523 ( .A1(n3525), .A2(n4212), .ZN(n5983) );
  NAND2_X1 U3524 ( .A1(n6700), .A2(n4591), .ZN(n5479) );
  OAI21_X1 U3525 ( .B1(n5562), .B2(n5618), .A(n4121), .ZN(n4122) );
  AND2_X1 U3526 ( .A1(n3506), .A2(n4602), .ZN(n3505) );
  NAND2_X1 U3527 ( .A1(n4589), .A2(n4588), .ZN(n4590) );
  OR2_X1 U3528 ( .A1(n4579), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6694)
         );
  OR2_X1 U3529 ( .A1(n4583), .A2(n4582), .ZN(n4589) );
  NAND2_X1 U3530 ( .A1(n4543), .A2(n4542), .ZN(n4809) );
  NAND2_X1 U3531 ( .A1(n4012), .A2(n4011), .ZN(n4573) );
  NOR2_X1 U3532 ( .A1(n5523), .A2(n6726), .ZN(n6954) );
  NAND2_X2 U3533 ( .A1(n5839), .A2(n5029), .ZN(n7086) );
  OAI21_X1 U3534 ( .B1(n5055), .B2(INSTADDRPOINTER_REG_1__SCAN_IN), .A(n5053), 
        .ZN(n4537) );
  NAND2_X1 U3535 ( .A1(n3948), .A2(n4849), .ZN(n3971) );
  NAND2_X1 U3536 ( .A1(n4530), .A2(n4529), .ZN(n5055) );
  AND2_X2 U3537 ( .A1(n4881), .A2(n3947), .ZN(n4960) );
  OR2_X1 U3538 ( .A1(n3915), .A2(n3914), .ZN(n4881) );
  NAND2_X1 U3539 ( .A1(n3915), .A2(n3914), .ZN(n3947) );
  NOR2_X1 U3540 ( .A1(n5717), .A2(n5718), .ZN(n5734) );
  OR2_X1 U3541 ( .A1(n5564), .A2(n4473), .ZN(n5717) );
  NAND2_X1 U3542 ( .A1(n3911), .A2(n3910), .ZN(n3915) );
  NAND2_X1 U3543 ( .A1(n4842), .A2(n7046), .ZN(n3939) );
  CLKBUF_X1 U3544 ( .A(n4783), .Z(n3447) );
  NAND2_X1 U3545 ( .A1(n3878), .A2(n3877), .ZN(n7057) );
  NAND2_X1 U3546 ( .A1(n3889), .A2(n3807), .ZN(n3891) );
  NAND2_X1 U3547 ( .A1(n3896), .A2(n3895), .ZN(n3919) );
  CLKBUF_X1 U3548 ( .A(n4404), .Z(n3431) );
  AND2_X1 U3549 ( .A1(n3823), .A2(n3822), .ZN(n4404) );
  AND3_X1 U3550 ( .A1(n3819), .A2(n3429), .A3(n3455), .ZN(n3824) );
  NAND2_X1 U3551 ( .A1(n4410), .A2(n3434), .ZN(n4672) );
  NOR2_X1 U3552 ( .A1(n3792), .A2(n4406), .ZN(n4410) );
  NAND2_X1 U3553 ( .A1(n4705), .A2(n4833), .ZN(n4431) );
  AND2_X1 U3554 ( .A1(n3794), .A2(n5169), .ZN(n3434) );
  OR2_X1 U3555 ( .A1(n4627), .A2(n4405), .ZN(n4785) );
  CLKBUF_X1 U3556 ( .A(n3881), .Z(n4668) );
  INV_X4 U3557 ( .A(n4418), .ZN(n5184) );
  AND2_X1 U3558 ( .A1(n4867), .A2(n4531), .ZN(n4626) );
  INV_X2 U3559 ( .A(n3848), .ZN(n4871) );
  AND2_X1 U3560 ( .A1(n3775), .A2(n3774), .ZN(n3776) );
  NAND2_X1 U3561 ( .A1(n3647), .A2(n3646), .ZN(n3781) );
  NAND2_X1 U3562 ( .A1(n3454), .A2(n3449), .ZN(n4531) );
  AND4_X1 U3563 ( .A1(n3671), .A2(n3670), .A3(n3669), .A4(n3668), .ZN(n3687)
         );
  AND4_X1 U3564 ( .A1(n3679), .A2(n3678), .A3(n3677), .A4(n3676), .ZN(n3685)
         );
  AND4_X1 U3565 ( .A1(n3675), .A2(n3674), .A3(n3673), .A4(n3672), .ZN(n3686)
         );
  AND4_X1 U3566 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3775)
         );
  AND4_X1 U3567 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3778)
         );
  AND4_X1 U3568 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3774)
         );
  AND4_X1 U3569 ( .A1(n3645), .A2(n3644), .A3(n3643), .A4(n3642), .ZN(n3646)
         );
  AND4_X1 U3570 ( .A1(n3729), .A2(n3728), .A3(n3727), .A4(n3726), .ZN(n3747)
         );
  AND4_X1 U3571 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3647)
         );
  AND4_X1 U3572 ( .A1(n3760), .A2(n3759), .A3(n3758), .A4(n3757), .ZN(n3777)
         );
  AND4_X1 U3573 ( .A1(n3655), .A2(n3654), .A3(n3653), .A4(n3652), .ZN(n3666)
         );
  AND4_X1 U3574 ( .A1(n3698), .A2(n3697), .A3(n3696), .A4(n3695), .ZN(n3714)
         );
  AND4_X1 U3575 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(n3667)
         );
  AND4_X1 U3576 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3660), .ZN(n3664)
         );
  AND4_X1 U3577 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(n3665)
         );
  BUF_X2 U3578 ( .A(n3725), .Z(n4643) );
  BUF_X2 U3579 ( .A(n3761), .Z(n4642) );
  AND2_X2 U3580 ( .A1(n3550), .A2(n6554), .ZN(n3860) );
  AND2_X2 U3581 ( .A1(n6555), .A2(n3549), .ZN(n3739) );
  AND2_X2 U3582 ( .A1(n4927), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4934)
         );
  INV_X1 U3583 ( .A(STATE_REG_2__SCAN_IN), .ZN(n7074) );
  INV_X2 U3584 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7046) );
  NAND2_X1 U3585 ( .A1(n6112), .A2(n3426), .ZN(n3423) );
  OR2_X1 U3586 ( .A1(n3425), .A2(n3493), .ZN(n3424) );
  INV_X1 U3587 ( .A(n4616), .ZN(n3425) );
  AND2_X1 U3588 ( .A1(n3497), .A2(n4616), .ZN(n3426) );
  INV_X1 U3589 ( .A(n6189), .ZN(n3427) );
  INV_X1 U3590 ( .A(n3793), .ZN(n3428) );
  NOR2_X2 U3591 ( .A1(n5887), .A2(n5869), .ZN(n5870) );
  OR2_X1 U3592 ( .A1(n3453), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U3593 ( .A1(n5169), .A2(n4418), .ZN(n5843) );
  AND2_X2 U3594 ( .A1(n5882), .A2(n3463), .ZN(n4703) );
  NOR2_X2 U3595 ( .A1(n5045), .A2(n5122), .ZN(n5123) );
  AND2_X1 U3596 ( .A1(n3779), .A2(n4785), .ZN(n3429) );
  NAND2_X1 U3597 ( .A1(n3784), .A2(n3783), .ZN(n3430) );
  NAND2_X1 U3598 ( .A1(n3784), .A2(n3783), .ZN(n3786) );
  INV_X1 U3599 ( .A(n6089), .ZN(n6187) );
  XNOR2_X1 U3600 ( .A(n4573), .B(n4025), .ZN(n4581) );
  NAND2_X1 U3601 ( .A1(n3802), .A2(n3801), .ZN(n3432) );
  OAI21_X1 U3602 ( .B1(n3799), .B2(n4418), .A(n4855), .ZN(n3433) );
  NAND2_X1 U3603 ( .A1(n3802), .A2(n3801), .ZN(n3889) );
  OAI21_X1 U3604 ( .B1(n3799), .B2(n4418), .A(n4855), .ZN(n3820) );
  INV_X1 U3605 ( .A(n3435), .ZN(n4733) );
  CLKBUF_X1 U3606 ( .A(n5691), .Z(n3436) );
  NAND2_X1 U3607 ( .A1(n4604), .A2(n5679), .ZN(n5691) );
  AND2_X1 U3608 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4809), .ZN(n3437)
         );
  NAND3_X1 U3609 ( .A1(n3430), .A2(n3813), .A3(n3456), .ZN(n3439) );
  NAND3_X1 U3610 ( .A1(n3786), .A2(n3813), .A3(n3456), .ZN(n3799) );
  NOR2_X2 U3611 ( .A1(n5951), .A2(n3518), .ZN(n5910) );
  NAND2_X2 U3612 ( .A1(n5971), .A2(n5972), .ZN(n5951) );
  NAND2_X1 U3613 ( .A1(n3878), .A2(n3852), .ZN(n3912) );
  AND2_X1 U3614 ( .A1(n5837), .A2(n3781), .ZN(n3854) );
  AND2_X1 U3615 ( .A1(n3913), .A2(n3912), .ZN(n3914) );
  NAND2_X1 U3616 ( .A1(n3824), .A2(n4404), .ZN(n3846) );
  AND2_X1 U3617 ( .A1(n3550), .A2(n6554), .ZN(n3440) );
  AND2_X4 U3618 ( .A1(n3468), .A2(n3467), .ZN(n4949) );
  AND2_X1 U3619 ( .A1(n6555), .A2(n4917), .ZN(n3441) );
  AND2_X4 U3620 ( .A1(n6555), .A2(n4934), .ZN(n3734) );
  AND2_X4 U3621 ( .A1(n4934), .A2(n4790), .ZN(n3903) );
  AND2_X2 U3622 ( .A1(n4934), .A2(n6554), .ZN(n3859) );
  NAND2_X2 U3623 ( .A1(n6126), .A2(n4613), .ZN(n6112) );
  OR2_X1 U3624 ( .A1(n3816), .A2(n3815), .ZN(n4742) );
  AND2_X2 U3625 ( .A1(n3785), .A2(n3793), .ZN(n4406) );
  INV_X2 U3626 ( .A(n3781), .ZN(n3793) );
  NAND2_X2 U3627 ( .A1(n5774), .A2(n5777), .ZN(n5776) );
  AND2_X2 U3628 ( .A1(n4835), .A2(n4836), .ZN(n4767) );
  NOR2_X2 U3629 ( .A1(n4821), .A2(n4910), .ZN(n4835) );
  XNOR2_X2 U3630 ( .A(n4703), .B(n4702), .ZN(n5821) );
  XNOR2_X1 U3631 ( .A(n3847), .B(n3846), .ZN(n3880) );
  AND2_X2 U3632 ( .A1(n5882), .A2(n5881), .ZN(n5872) );
  NOR2_X4 U3633 ( .A1(n5897), .A2(n5899), .ZN(n5882) );
  XNOR2_X2 U3634 ( .A(n3891), .B(n3890), .ZN(n4843) );
  XNOR2_X1 U3635 ( .A(n4849), .B(n3947), .ZN(n4883) );
  BUF_X1 U3636 ( .A(n4525), .Z(n3446) );
  INV_X1 U3637 ( .A(n3947), .ZN(n3948) );
  NOR2_X2 U3638 ( .A1(n3428), .A2(n7128), .ZN(n4154) );
  NOR2_X1 U3639 ( .A1(n3970), .A2(n3450), .ZN(n3514) );
  INV_X1 U3640 ( .A(n3971), .ZN(n3513) );
  AND2_X2 U3641 ( .A1(n3921), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3550)
         );
  INV_X1 U3642 ( .A(n6186), .ZN(n3492) );
  NOR2_X1 U3643 ( .A1(n5307), .A2(n3473), .ZN(n3472) );
  INV_X1 U3644 ( .A(n5535), .ZN(n3473) );
  OR2_X1 U3645 ( .A1(n3848), .A2(n7046), .ZN(n3898) );
  NAND2_X1 U3646 ( .A1(n3898), .A2(n3897), .ZN(n4397) );
  AND2_X1 U3647 ( .A1(n6732), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4417) );
  AND2_X1 U3648 ( .A1(n4626), .A2(n3793), .ZN(n3794) );
  AND2_X1 U3649 ( .A1(n6875), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5852) );
  OR2_X1 U3650 ( .A1(n4729), .A2(n4784), .ZN(n4774) );
  AOI21_X1 U3651 ( .B1(n4581), .B2(n4154), .A(n4032), .ZN(n5046) );
  NAND2_X1 U3652 ( .A1(n6112), .A2(n3497), .ZN(n3495) );
  NAND2_X1 U3653 ( .A1(n6171), .A2(n3498), .ZN(n3497) );
  INV_X1 U3654 ( .A(n5809), .ZN(n3498) );
  AND2_X1 U3655 ( .A1(n4002), .A2(n4001), .ZN(n4010) );
  OR2_X1 U3656 ( .A1(n3981), .A2(n3980), .ZN(n4564) );
  INV_X1 U3657 ( .A(n3512), .ZN(n3511) );
  AOI21_X1 U3658 ( .B1(n3970), .B2(n3450), .A(n4582), .ZN(n3512) );
  NOR2_X1 U3659 ( .A1(n3532), .A2(n4345), .ZN(n3531) );
  INV_X1 U3660 ( .A(n5873), .ZN(n3532) );
  NAND2_X1 U3661 ( .A1(n3527), .A2(n4212), .ZN(n3526) );
  INV_X1 U3662 ( .A(n5984), .ZN(n3527) );
  INV_X1 U3663 ( .A(n3517), .ZN(n3516) );
  INV_X1 U3664 ( .A(n3881), .ZN(n4662) );
  OR2_X1 U3665 ( .A1(n3909), .A2(n3908), .ZN(n4545) );
  INV_X1 U3666 ( .A(n4960), .ZN(n5208) );
  NAND2_X1 U3667 ( .A1(n4509), .A2(n3477), .ZN(n3476) );
  INV_X1 U3668 ( .A(n5954), .ZN(n3477) );
  INV_X1 U3669 ( .A(n6041), .ZN(n3479) );
  INV_X1 U3670 ( .A(n5748), .ZN(n3503) );
  NOR2_X1 U3671 ( .A1(n3504), .A2(n3501), .ZN(n3500) );
  INV_X1 U3672 ( .A(n4608), .ZN(n3504) );
  INV_X1 U3673 ( .A(n5722), .ZN(n3501) );
  AND2_X1 U3674 ( .A1(n3470), .A2(n3472), .ZN(n3469) );
  INV_X1 U3675 ( .A(n5566), .ZN(n3470) );
  INV_X1 U3676 ( .A(n4770), .ZN(n3482) );
  NAND2_X1 U3677 ( .A1(n4833), .A2(n4490), .ZN(n4513) );
  AND2_X1 U3678 ( .A1(n4844), .A2(n3894), .ZN(n4877) );
  INV_X1 U3679 ( .A(n3446), .ZN(n5207) );
  OR2_X1 U3680 ( .A1(n4431), .A2(EBX_REG_1__SCAN_IN), .ZN(n4425) );
  NAND2_X1 U3681 ( .A1(n5160), .A2(n5159), .ZN(n6875) );
  AND2_X1 U3682 ( .A1(n4248), .A2(n4247), .ZN(n6019) );
  OAI21_X1 U3683 ( .B1(n6099), .B2(n3690), .A(n4325), .ZN(n5899) );
  NAND2_X1 U3684 ( .A1(n3519), .A2(n5924), .ZN(n3518) );
  INV_X1 U3685 ( .A(n3521), .ZN(n3519) );
  NAND2_X1 U3686 ( .A1(n4265), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4287)
         );
  NAND2_X1 U3687 ( .A1(n3520), .A2(n4286), .ZN(n5936) );
  INV_X1 U3688 ( .A(n5951), .ZN(n3520) );
  OR2_X1 U3689 ( .A1(n6966), .A2(n3690), .ZN(n4211) );
  INV_X1 U3690 ( .A(n5046), .ZN(n4033) );
  OR2_X1 U3691 ( .A1(n6988), .A2(n7051), .ZN(n5110) );
  AND2_X1 U3692 ( .A1(n6077), .A2(n4620), .ZN(n4689) );
  NOR2_X1 U3693 ( .A1(n6105), .A2(n3494), .ZN(n3493) );
  INV_X1 U3694 ( .A(n3496), .ZN(n3494) );
  AND2_X1 U3695 ( .A1(n3460), .A2(n3533), .ZN(n3491) );
  AND2_X1 U3696 ( .A1(n6034), .A2(n5987), .ZN(n6022) );
  NAND2_X1 U3697 ( .A1(n4732), .A2(n6992), .ZN(n4756) );
  OR2_X1 U3698 ( .A1(n4731), .A2(n4730), .ZN(n4732) );
  OR2_X1 U3699 ( .A1(n7057), .A2(n4582), .ZN(n4535) );
  NAND2_X1 U3700 ( .A1(n3880), .A2(n7046), .ZN(n3878) );
  INV_X1 U3701 ( .A(n7057), .ZN(n5629) );
  NOR2_X1 U3702 ( .A1(n3487), .A2(n5855), .ZN(n3486) );
  INV_X1 U3703 ( .A(n5858), .ZN(n3487) );
  OR2_X1 U3704 ( .A1(n4681), .A2(n4419), .ZN(n4420) );
  NAND2_X1 U3705 ( .A1(n6047), .A2(n5028), .ZN(n6045) );
  NAND2_X1 U3706 ( .A1(n5277), .A2(n4683), .ZN(n5839) );
  XNOR2_X1 U3707 ( .A(n4697), .B(n5854), .ZN(n5179) );
  OR2_X1 U3708 ( .A1(n4696), .A2(n5817), .ZN(n4697) );
  INV_X1 U3709 ( .A(n4701), .ZN(n4702) );
  XNOR2_X1 U3710 ( .A(n4708), .B(n3488), .ZN(n5834) );
  INV_X1 U3711 ( .A(n5846), .ZN(n3488) );
  OAI21_X1 U3712 ( .B1(n4707), .B2(n4706), .A(n5845), .ZN(n4708) );
  OR2_X1 U3713 ( .A1(n4299), .A2(n4297), .ZN(n4310) );
  CLKBUF_X2 U3714 ( .A(n3859), .Z(n4650) );
  INV_X1 U3715 ( .A(n4009), .ZN(n4012) );
  OR2_X1 U3716 ( .A1(n4022), .A2(n4021), .ZN(n4595) );
  OR2_X1 U3717 ( .A1(n4000), .A2(n3999), .ZN(n4585) );
  NAND2_X1 U3718 ( .A1(n4573), .A2(n4572), .ZN(n4593) );
  OR2_X1 U3719 ( .A1(n3958), .A2(n3957), .ZN(n4561) );
  OR2_X1 U3720 ( .A1(n4406), .A2(n4871), .ZN(n3810) );
  INV_X1 U3721 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4393) );
  NAND2_X1 U3722 ( .A1(n4406), .A2(n4871), .ZN(n3716) );
  OAI21_X1 U3723 ( .B1(n3971), .B2(n3970), .A(n3450), .ZN(n3515) );
  NAND2_X1 U3724 ( .A1(n3522), .A2(n4286), .ZN(n3521) );
  INV_X1 U3725 ( .A(n5937), .ZN(n3522) );
  AND2_X1 U3726 ( .A1(n4161), .A2(n5716), .ZN(n3517) );
  NAND2_X1 U3727 ( .A1(n3529), .A2(n3465), .ZN(n4126) );
  NAND2_X1 U3728 ( .A1(n5304), .A2(n3528), .ZN(n5562) );
  AND2_X1 U3729 ( .A1(n5532), .A2(n5563), .ZN(n3528) );
  AND2_X1 U3730 ( .A1(n5611), .A2(n5478), .ZN(n3508) );
  INV_X1 U3731 ( .A(n4600), .ZN(n3509) );
  AOI21_X1 U3732 ( .B1(n3971), .B2(n3450), .A(n3511), .ZN(n3510) );
  OR2_X1 U3733 ( .A1(n5169), .A2(n7046), .ZN(n3897) );
  INV_X1 U3734 ( .A(n4848), .ZN(n4853) );
  AOI21_X1 U3735 ( .B1(n7048), .B2(n7040), .A(n4847), .ZN(n4848) );
  OR2_X1 U3736 ( .A1(n3892), .A2(n3921), .ZN(n3926) );
  NOR2_X1 U3737 ( .A1(n5309), .A2(n5307), .ZN(n5536) );
  AND2_X1 U3738 ( .A1(n4430), .A2(n4429), .ZN(n4813) );
  AND4_X1 U3739 ( .A1(n4049), .A2(n4048), .A3(n4047), .A4(n4046), .ZN(n5122)
         );
  OR2_X1 U3740 ( .A1(n5275), .A2(n5111), .ZN(n5112) );
  INV_X1 U3741 ( .A(n5277), .ZN(n5255) );
  AND2_X1 U3742 ( .A1(n5156), .A2(n7028), .ZN(n4991) );
  INV_X1 U3743 ( .A(n4300), .ZN(n4667) );
  AND2_X1 U3744 ( .A1(n3531), .A2(n3462), .ZN(n3530) );
  AND2_X1 U3745 ( .A1(n3542), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4334)
         );
  NAND2_X1 U3746 ( .A1(n4334), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4638)
         );
  OR2_X1 U3747 ( .A1(n4287), .A2(n6133), .ZN(n4296) );
  AND2_X1 U3748 ( .A1(n3541), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4265)
         );
  INV_X1 U3749 ( .A(n4249), .ZN(n3541) );
  OR2_X1 U3750 ( .A1(n6141), .A2(n3690), .ZN(n4285) );
  NAND2_X1 U3751 ( .A1(n6019), .A2(n3524), .ZN(n3523) );
  INV_X1 U3752 ( .A(n3526), .ZN(n3524) );
  AND2_X1 U3753 ( .A1(n3540), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4229)
         );
  NAND2_X1 U3754 ( .A1(n4229), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4249)
         );
  INV_X1 U3755 ( .A(n5776), .ZN(n3525) );
  NAND2_X1 U3756 ( .A1(n4162), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4176)
         );
  CLKBUF_X1 U3757 ( .A(n5774), .Z(n5775) );
  NOR2_X1 U3758 ( .A1(n4127), .A2(n4128), .ZN(n4145) );
  NOR2_X1 U3759 ( .A1(n4092), .A2(n5624), .ZN(n4123) );
  NAND2_X1 U3760 ( .A1(n4123), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4127)
         );
  NOR2_X1 U3761 ( .A1(n4063), .A2(n5541), .ZN(n4079) );
  NAND2_X1 U3762 ( .A1(n4050), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4063)
         );
  INV_X1 U3763 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5541) );
  OR2_X1 U3764 ( .A1(n4026), .A2(n4028), .ZN(n4045) );
  INV_X1 U3765 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4028) );
  AOI21_X1 U3766 ( .B1(n4574), .B2(n4154), .A(n4007), .ZN(n5022) );
  NOR2_X1 U3767 ( .A1(n3984), .A2(n3987), .ZN(n4003) );
  INV_X1 U3768 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3987) );
  NAND2_X1 U3769 ( .A1(n3964), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3984)
         );
  AND3_X1 U3770 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A3(PHYADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n3964) );
  AOI21_X1 U3771 ( .B1(n4960), .B2(n4572), .A(n4540), .ZN(n4811) );
  NAND2_X1 U3772 ( .A1(n4617), .A2(n3461), .ZN(n6087) );
  OR3_X1 U3773 ( .A1(n5938), .A2(n3476), .A3(n3475), .ZN(n3474) );
  INV_X1 U3774 ( .A(n5901), .ZN(n3475) );
  NAND2_X1 U3775 ( .A1(n6089), .A2(n4615), .ZN(n3496) );
  NOR3_X1 U3776 ( .A1(n5975), .A2(n5938), .A3(n5954), .ZN(n5939) );
  OR2_X1 U3777 ( .A1(n6024), .A2(n5973), .ZN(n5975) );
  NAND2_X1 U3778 ( .A1(n6022), .A2(n6021), .ZN(n6024) );
  OR2_X1 U3779 ( .A1(n6171), .A2(n4612), .ZN(n4613) );
  AND2_X1 U3780 ( .A1(n6042), .A2(n3464), .ZN(n6034) );
  INV_X1 U3781 ( .A(n6031), .ZN(n3478) );
  NAND2_X1 U3782 ( .A1(n6042), .A2(n3458), .ZN(n6032) );
  NAND2_X1 U3783 ( .A1(n6042), .A2(n6041), .ZN(n6044) );
  AND2_X1 U3784 ( .A1(n5734), .A2(n5735), .ZN(n6042) );
  AOI21_X1 U3785 ( .B1(n3503), .B2(n4608), .A(n3457), .ZN(n3502) );
  OR2_X1 U3786 ( .A1(n6171), .A2(n6832), .ZN(n6195) );
  AND2_X1 U3787 ( .A1(n4477), .A2(n4476), .ZN(n5718) );
  NAND2_X1 U3788 ( .A1(n4607), .A2(n5722), .ZN(n5749) );
  NAND2_X1 U3789 ( .A1(n5749), .A2(n5748), .ZN(n5747) );
  NAND2_X1 U3790 ( .A1(n3471), .A2(n3472), .ZN(n5565) );
  OR2_X1 U3791 ( .A1(n6187), .A2(n5701), .ZN(n5690) );
  AND2_X1 U3792 ( .A1(n4459), .A2(n4458), .ZN(n5126) );
  NOR2_X1 U3793 ( .A1(n4915), .A2(n3480), .ZN(n5049) );
  NAND2_X1 U3794 ( .A1(n3482), .A2(n3451), .ZN(n3480) );
  AND2_X1 U3795 ( .A1(n4454), .A2(n4453), .ZN(n5048) );
  NAND2_X1 U3796 ( .A1(n5049), .A2(n5048), .ZN(n5125) );
  NOR2_X1 U3797 ( .A1(n4915), .A2(n3481), .ZN(n5024) );
  NAND2_X1 U3798 ( .A1(n3482), .A2(n4445), .ZN(n3481) );
  OR2_X1 U3799 ( .A1(n4915), .A2(n4840), .ZN(n4838) );
  AND2_X1 U3800 ( .A1(n4813), .A2(n4812), .ZN(n4913) );
  NAND2_X1 U3801 ( .A1(n4913), .A2(n4912), .ZN(n4915) );
  NAND2_X1 U3802 ( .A1(n4751), .A2(n6982), .ZN(n6744) );
  NAND2_X1 U3803 ( .A1(n4439), .A2(n4490), .ZN(n5844) );
  INV_X1 U3804 ( .A(n4756), .ZN(n4751) );
  OR2_X1 U3805 ( .A1(n3892), .A2(n4927), .ZN(n3896) );
  INV_X1 U3806 ( .A(n3807), .ZN(n3489) );
  NAND2_X1 U3807 ( .A1(n7046), .A2(n4853), .ZN(n4953) );
  OR2_X1 U3808 ( .A1(n4401), .A2(n4400), .ZN(n4402) );
  AND2_X2 U3809 ( .A1(n3467), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6554)
         );
  NAND2_X1 U3810 ( .A1(n4713), .A2(n5184), .ZN(n4923) );
  NOR2_X1 U3811 ( .A1(n3445), .A2(n5415), .ZN(n5214) );
  OR2_X1 U3812 ( .A1(n4955), .A2(n3446), .ZN(n4971) );
  AND2_X1 U3813 ( .A1(n5286), .A2(n5285), .ZN(n5641) );
  AND2_X1 U3814 ( .A1(n5416), .A2(n3445), .ZN(n7125) );
  NOR2_X1 U3815 ( .A1(n3444), .A2(n7139), .ZN(n5569) );
  NOR2_X1 U3816 ( .A1(n5282), .A2(n7139), .ZN(n5571) );
  INV_X1 U3817 ( .A(n4531), .ZN(n4863) );
  NOR2_X1 U3818 ( .A1(n5089), .A2(n4880), .ZN(n4856) );
  NAND2_X1 U3819 ( .A1(n4854), .A2(n4853), .ZN(n5193) );
  AND2_X1 U3820 ( .A1(n4417), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6992) );
  NOR2_X1 U3821 ( .A1(n5110), .A2(n4672), .ZN(n5156) );
  INV_X2 U3822 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n7128) );
  OR2_X1 U3823 ( .A1(n5156), .A2(n5155), .ZN(n6739) );
  INV_X1 U3824 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U3825 ( .A1(n5852), .A2(n5166), .ZN(n6905) );
  INV_X1 U3826 ( .A(n6973), .ZN(n6950) );
  AND2_X1 U3827 ( .A1(n6875), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6955) );
  INV_X1 U3828 ( .A(n6045), .ZN(n6037) );
  OAI21_X1 U3829 ( .B1(n5872), .B2(n5873), .A(n4344), .ZN(n6054) );
  INV_X1 U3830 ( .A(n5839), .ZN(n7096) );
  INV_X1 U3831 ( .A(n5836), .ZN(n7093) );
  NAND2_X1 U3832 ( .A1(n5839), .A2(n5030), .ZN(n5745) );
  CLKBUF_X2 U3833 ( .A(n5269), .Z(n5275) );
  AOI21_X1 U3834 ( .B1(n5884), .B2(n5883), .A(n5872), .ZN(n6094) );
  INV_X1 U3835 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6180) );
  NAND2_X2 U3836 ( .A1(n4628), .A2(n7021), .ZN(n6993) );
  INV_X1 U3837 ( .A(n5110), .ZN(n4628) );
  XNOR2_X1 U3838 ( .A(n4624), .B(n4623), .ZN(n6230) );
  OR2_X1 U3839 ( .A1(n4756), .A2(n4755), .ZN(n6836) );
  NAND2_X1 U3840 ( .A1(n5612), .A2(n5611), .ZN(n5610) );
  NAND2_X1 U3841 ( .A1(n5477), .A2(n4600), .ZN(n5612) );
  INV_X1 U3843 ( .A(n6836), .ZN(n6846) );
  INV_X1 U3844 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7123) );
  INV_X1 U3845 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7008) );
  INV_X1 U3846 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5128) );
  INV_X1 U3847 ( .A(n3444), .ZN(n5282) );
  INV_X1 U3848 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6732) );
  NOR2_X1 U3849 ( .A1(n4629), .A2(n6988), .ZN(n4847) );
  NOR2_X1 U3850 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6560) );
  NAND2_X1 U3851 ( .A1(n5214), .A2(n5629), .ZN(n5458) );
  INV_X1 U3852 ( .A(n5197), .ZN(n5361) );
  NOR2_X1 U3853 ( .A1(n4971), .A2(n7057), .ZN(n5198) );
  INV_X1 U3854 ( .A(n5198), .ZN(n5334) );
  AND2_X1 U3855 ( .A1(n5417), .A2(n5629), .ZN(n7270) );
  INV_X1 U3856 ( .A(n7259), .ZN(n5451) );
  INV_X1 U3857 ( .A(n7270), .ZN(n5450) );
  AOI22_X1 U3858 ( .A1(n5637), .A2(n7114), .B1(n5635), .B2(n5634), .ZN(n5676)
         );
  INV_X1 U3859 ( .A(n5392), .ZN(n7243) );
  OR2_X1 U3860 ( .A1(n5132), .A2(n7057), .ZN(n5392) );
  NAND2_X1 U3861 ( .A1(DATAI_1_), .A2(n5285), .ZN(n7170) );
  NAND2_X1 U3862 ( .A1(DATAI_2_), .A2(n5285), .ZN(n7185) );
  NAND2_X1 U3863 ( .A1(DATAI_3_), .A2(n5285), .ZN(n7199) );
  NAND2_X1 U3864 ( .A1(DATAI_5_), .A2(n5285), .ZN(n7226) );
  NAND2_X1 U3865 ( .A1(DATAI_6_), .A2(n5285), .ZN(n7242) );
  NAND2_X1 U3866 ( .A1(n4856), .A2(n5629), .ZN(n5603) );
  NAND2_X1 U3867 ( .A1(n4856), .A2(n7057), .ZN(n5393) );
  NAND2_X1 U3868 ( .A1(DATAI_7_), .A2(n5285), .ZN(n7275) );
  OAI21_X1 U3869 ( .B1(n5834), .B2(n6975), .A(n3483), .ZN(U2797) );
  INV_X1 U3870 ( .A(n3484), .ZN(n3483) );
  NOR2_X1 U3871 ( .A1(n5835), .A2(n3486), .ZN(n3485) );
  NAND2_X1 U3872 ( .A1(n5821), .A2(n4704), .ZN(n4712) );
  OAI21_X1 U3873 ( .B1(n6051), .B2(n6039), .A(n4524), .ZN(U2830) );
  OR2_X1 U3874 ( .A1(n5861), .A2(n6045), .ZN(n4523) );
  AND2_X2 U3875 ( .A1(n3550), .A2(n4949), .ZN(n3834) );
  AND2_X2 U3876 ( .A1(n3550), .A2(n6555), .ZN(n3865) );
  AND2_X2 U3877 ( .A1(n4949), .A2(n4917), .ZN(n3725) );
  AND4_X1 U3878 ( .A1(n3724), .A2(n3723), .A3(n3722), .A4(n3721), .ZN(n3449)
         );
  AND2_X1 U3879 ( .A1(n3983), .A2(n3982), .ZN(n3450) );
  AND2_X1 U3880 ( .A1(n4445), .A2(n5023), .ZN(n3451) );
  AND2_X1 U3881 ( .A1(n3515), .A2(n4009), .ZN(n3452) );
  NOR3_X1 U3882 ( .A1(n5975), .A2(n5938), .A3(n3476), .ZN(n5900) );
  NAND2_X1 U3883 ( .A1(n3427), .A2(n3533), .ZN(n6170) );
  NOR2_X1 U3884 ( .A1(n5951), .A2(n3521), .ZN(n5923) );
  OR2_X1 U3885 ( .A1(n5975), .A2(n3474), .ZN(n3453) );
  INV_X1 U3886 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3467) );
  NOR2_X1 U3887 ( .A1(n5776), .A2(n3526), .ZN(n5985) );
  AND4_X1 U3888 ( .A1(n3720), .A2(n3719), .A3(n3718), .A4(n3717), .ZN(n3454)
         );
  NAND2_X1 U3889 ( .A1(n5872), .A2(n5873), .ZN(n4344) );
  NAND2_X1 U3890 ( .A1(n3495), .A2(n3496), .ZN(n6103) );
  AND3_X1 U3891 ( .A1(n3818), .A2(n3817), .A3(n4742), .ZN(n3455) );
  NAND2_X1 U3892 ( .A1(n4425), .A2(n4424), .ZN(n4429) );
  OR2_X1 U3893 ( .A1(n4354), .A2(n4867), .ZN(n3456) );
  NOR2_X1 U3894 ( .A1(n6171), .A2(n5769), .ZN(n3457) );
  NAND2_X1 U3895 ( .A1(n3513), .A2(n3514), .ZN(n4009) );
  AND2_X1 U3896 ( .A1(n3715), .A2(n5837), .ZN(n3752) );
  INV_X1 U3897 ( .A(n3445), .ZN(n5063) );
  AND2_X2 U3898 ( .A1(n3550), .A2(n4790), .ZN(n3768) );
  NAND2_X1 U3899 ( .A1(n5714), .A2(n3517), .ZN(n5731) );
  NAND2_X1 U3900 ( .A1(n5714), .A2(n5716), .ZN(n5715) );
  AND2_X2 U3901 ( .A1(n4917), .A2(n4790), .ZN(n3827) );
  NOR2_X1 U3902 ( .A1(n5778), .A2(n3479), .ZN(n3458) );
  AND2_X1 U3903 ( .A1(n5123), .A2(n5305), .ZN(n5304) );
  AND2_X1 U3904 ( .A1(n5304), .A2(n5532), .ZN(n5531) );
  AND4_X2 U3905 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n4867)
         );
  OR2_X1 U3906 ( .A1(n5975), .A2(n5954), .ZN(n3459) );
  NAND2_X1 U3907 ( .A1(n3507), .A2(n3505), .ZN(n5677) );
  NAND2_X1 U3908 ( .A1(n5747), .A2(n4608), .ZN(n5762) );
  AND2_X1 U3909 ( .A1(n4126), .A2(n4122), .ZN(n5705) );
  NAND2_X1 U3910 ( .A1(n6171), .A2(n5791), .ZN(n3460) );
  NAND2_X1 U3911 ( .A1(n6171), .A2(n6252), .ZN(n3461) );
  AND2_X1 U3912 ( .A1(n4418), .A2(n4354), .ZN(n4572) );
  AND2_X1 U3913 ( .A1(n4701), .A2(n5881), .ZN(n3462) );
  AND2_X1 U3914 ( .A1(n3531), .A2(n5881), .ZN(n3463) );
  AND2_X1 U3915 ( .A1(n3458), .A2(n3478), .ZN(n3464) );
  OR2_X1 U3916 ( .A1(n5125), .A2(n5126), .ZN(n5309) );
  INV_X1 U3917 ( .A(n5309), .ZN(n3471) );
  AND2_X1 U3918 ( .A1(n4120), .A2(n4119), .ZN(n3465) );
  NOR2_X1 U3919 ( .A1(n3516), .A2(n6040), .ZN(n3466) );
  INV_X1 U3920 ( .A(n4840), .ZN(n4445) );
  AND2_X1 U3921 ( .A1(n4444), .A2(n4443), .ZN(n4840) );
  NAND2_X2 U3922 ( .A1(n6047), .A2(n5837), .ZN(n6039) );
  AND2_X2 U3923 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4917) );
  INV_X2 U3924 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3468) );
  NAND2_X1 U3925 ( .A1(n3471), .A2(n3469), .ZN(n5564) );
  INV_X1 U3926 ( .A(n3919), .ZN(n3490) );
  AND2_X2 U3927 ( .A1(n3846), .A2(n3845), .ZN(n3890) );
  OR2_X2 U3928 ( .A1(n3920), .A2(n3490), .ZN(n4921) );
  NAND2_X1 U3929 ( .A1(n3492), .A2(n3491), .ZN(n6126) );
  NAND2_X1 U3930 ( .A1(n3499), .A2(n3502), .ZN(n4610) );
  NAND2_X1 U3931 ( .A1(n4607), .A2(n3500), .ZN(n3499) );
  NAND2_X1 U3932 ( .A1(n5479), .A2(n5478), .ZN(n5477) );
  NAND2_X1 U3933 ( .A1(n5611), .A2(n3509), .ZN(n3506) );
  NAND2_X1 U3934 ( .A1(n5479), .A2(n3508), .ZN(n3507) );
  NAND2_X1 U3935 ( .A1(n4009), .A2(n3510), .ZN(n4567) );
  INV_X1 U3936 ( .A(n5562), .ZN(n3529) );
  NAND2_X1 U3937 ( .A1(n5882), .A2(n3530), .ZN(n4671) );
  NAND3_X1 U3938 ( .A1(n4767), .A2(n4008), .A3(n4769), .ZN(n5021) );
  INV_X1 U3939 ( .A(n5021), .ZN(n4034) );
  NAND2_X1 U3940 ( .A1(n4767), .A2(n4769), .ZN(n4768) );
  NAND2_X1 U3941 ( .A1(n5783), .A2(n4622), .ZN(n4693) );
  INV_X1 U3942 ( .A(n5821), .ZN(n5842) );
  OR2_X1 U3943 ( .A1(n4786), .A2(n4753), .ZN(n7030) );
  AND2_X2 U3944 ( .A1(n6554), .A2(n4917), .ZN(n3762) );
  OR2_X1 U3945 ( .A1(n4627), .A2(n5169), .ZN(n3798) );
  AND2_X2 U3946 ( .A1(n5169), .A2(n5184), .ZN(n4407) );
  INV_X1 U3947 ( .A(n4541), .ZN(n4543) );
  NAND2_X1 U3948 ( .A1(n3781), .A2(n3750), .ZN(n3715) );
  AOI21_X1 U3949 ( .B1(n5850), .B2(n6710), .A(n4699), .ZN(n4700) );
  NAND2_X1 U3950 ( .A1(n5850), .A2(n4684), .ZN(n4687) );
  AOI22_X1 U3951 ( .A1(n6078), .A2(n4689), .B1(n6171), .B2(n4621), .ZN(n4624)
         );
  INV_X2 U3952 ( .A(n6685), .ZN(n6710) );
  INV_X1 U3953 ( .A(n3690), .ZN(n4343) );
  NAND2_X1 U3954 ( .A1(n6171), .A2(n6841), .ZN(n3533) );
  OR2_X1 U3955 ( .A1(n4627), .A2(n5184), .ZN(n3534) );
  NAND2_X1 U3956 ( .A1(n6171), .A2(n6233), .ZN(n3535) );
  NOR2_X1 U3957 ( .A1(n7046), .A2(n3805), .ZN(n3536) );
  NOR2_X1 U3958 ( .A1(n3447), .A2(n5174), .ZN(n3537) );
  NOR2_X1 U3959 ( .A1(n3447), .A2(n4843), .ZN(n3538) );
  OR2_X1 U3960 ( .A1(n5836), .A2(n6424), .ZN(n3539) );
  OAI21_X2 U3961 ( .B1(n4774), .B2(n7051), .A(n4420), .ZN(n6047) );
  INV_X1 U3962 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4128) );
  NOR2_X1 U3963 ( .A1(n5837), .A2(n7128), .ZN(n3881) );
  NAND2_X1 U3964 ( .A1(n4751), .A2(n4737), .ZN(n6756) );
  INV_X1 U3965 ( .A(n5730), .ZN(n4161) );
  NAND2_X1 U3966 ( .A1(n5706), .A2(n4126), .ZN(n5714) );
  AND2_X1 U3967 ( .A1(n4397), .A2(n4369), .ZN(n4374) );
  AND2_X1 U3968 ( .A1(n3790), .A2(n3789), .ZN(n3803) );
  NAND2_X1 U3969 ( .A1(n7123), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4359) );
  INV_X1 U3970 ( .A(n5022), .ZN(n4008) );
  INV_X1 U3971 ( .A(n3969), .ZN(n3970) );
  INV_X1 U3972 ( .A(n4010), .ZN(n4011) );
  OR2_X1 U3973 ( .A1(n3937), .A2(n3936), .ZN(n4554) );
  NAND2_X1 U3974 ( .A1(n3769), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U3975 ( .A1(n3734), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3762), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3643) );
  INV_X1 U3976 ( .A(n4359), .ZN(n4355) );
  INV_X1 U3977 ( .A(n4417), .ZN(n3923) );
  NAND2_X1 U3978 ( .A1(n3821), .A2(n3534), .ZN(n3823) );
  INV_X1 U3979 ( .A(n6030), .ZN(n4212) );
  INV_X1 U3980 ( .A(n5953), .ZN(n4286) );
  OR2_X1 U3981 ( .A1(n3841), .A2(n3840), .ZN(n4526) );
  INV_X1 U3982 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4542) );
  OR2_X1 U3983 ( .A1(n4394), .A2(n4393), .ZN(n4392) );
  NOR2_X1 U3984 ( .A1(n4307), .A2(n4308), .ZN(n4315) );
  INV_X1 U3985 ( .A(n4213), .ZN(n3540) );
  NAND2_X1 U3986 ( .A1(n6553), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4323) );
  NOR2_X1 U3987 ( .A1(n4045), .A2(n5505), .ZN(n4050) );
  INV_X1 U3988 ( .A(n4595), .ZN(n4592) );
  INV_X1 U3989 ( .A(n4392), .ZN(n4353) );
  NAND2_X1 U3990 ( .A1(n4389), .A2(n4572), .ZN(n4401) );
  NAND2_X1 U3991 ( .A1(n3926), .A2(n3925), .ZN(n4919) );
  INV_X1 U3992 ( .A(n6739), .ZN(n5160) );
  OR2_X1 U3993 ( .A1(n6974), .A2(n3690), .ZN(n4248) );
  AOI22_X1 U3994 ( .A1(n3734), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3552) );
  OR2_X1 U3995 ( .A1(n4296), .A2(n4301), .ZN(n4307) );
  INV_X1 U3996 ( .A(n4680), .ZN(n4746) );
  NAND2_X1 U3997 ( .A1(n4315), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4326)
         );
  INV_X1 U3998 ( .A(n4323), .ZN(n4664) );
  NAND2_X1 U3999 ( .A1(n4079), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4092)
         );
  INV_X1 U4000 ( .A(n4614), .ZN(n4603) );
  AND2_X1 U4001 ( .A1(n4488), .A2(n4487), .ZN(n6031) );
  OR2_X1 U4002 ( .A1(n4782), .A2(n4781), .ZN(n4944) );
  AND2_X1 U4003 ( .A1(n4999), .A2(n5063), .ZN(n5319) );
  NAND2_X1 U4004 ( .A1(n4353), .A2(n4352), .ZN(n4678) );
  OR3_X1 U4005 ( .A1(n5891), .A2(n6649), .A3(n6651), .ZN(n5862) );
  NOR2_X1 U4006 ( .A1(n4176), .A2(n6180), .ZN(n4193) );
  AND2_X1 U4007 ( .A1(n4145), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4162)
         );
  INV_X1 U4008 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U4009 ( .A1(n3452), .A2(n4154), .ZN(n3990) );
  NAND2_X1 U4010 ( .A1(n4603), .A2(n4622), .ZN(n5782) );
  NAND2_X1 U4011 ( .A1(n4567), .A2(n4566), .ZN(n4569) );
  OR2_X1 U4012 ( .A1(n6726), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6801) );
  NAND2_X1 U4013 ( .A1(n5214), .A2(n7057), .ZN(n5604) );
  NAND2_X1 U4014 ( .A1(n5630), .A2(n5063), .ZN(n5443) );
  INV_X1 U4015 ( .A(n5319), .ZN(n5360) );
  INV_X1 U4016 ( .A(n7266), .ZN(n5333) );
  NAND2_X1 U4017 ( .A1(n7125), .A2(n5629), .ZN(n7233) );
  OR2_X1 U4018 ( .A1(n5132), .A2(n5629), .ZN(n7108) );
  AND2_X1 U4019 ( .A1(n4403), .A2(n4402), .ZN(n6988) );
  AND2_X1 U4020 ( .A1(n4638), .A2(n4336), .ZN(n6081) );
  NAND2_X1 U4021 ( .A1(n4193), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4213)
         );
  INV_X1 U4022 ( .A(n6961), .ZN(n6978) );
  AND2_X1 U4023 ( .A1(n5852), .A2(n5163), .ZN(n6930) );
  INV_X1 U4024 ( .A(n6039), .ZN(n4704) );
  AND2_X1 U4025 ( .A1(n4479), .A2(n4478), .ZN(n5735) );
  INV_X1 U4026 ( .A(n6047), .ZN(n6012) );
  AND2_X1 U4027 ( .A1(n5839), .A2(n5838), .ZN(n7097) );
  NAND2_X1 U4028 ( .A1(n3990), .A2(n3989), .ZN(n4769) );
  AND2_X1 U4029 ( .A1(n5112), .A2(n6736), .ZN(n6577) );
  NOR2_X1 U4030 ( .A1(n4991), .A2(n5275), .ZN(n5230) );
  NOR2_X1 U4031 ( .A1(n5110), .A2(n7030), .ZN(n5269) );
  INV_X1 U4032 ( .A(n6157), .ZN(n7095) );
  NAND2_X1 U4034 ( .A1(n7128), .A2(n4629), .ZN(n7139) );
  NAND2_X1 U4035 ( .A1(n4003), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4026)
         );
  INV_X1 U4036 ( .A(n6707), .ZN(n6709) );
  INV_X1 U4037 ( .A(n4688), .ZN(n4623) );
  OR2_X1 U4038 ( .A1(n6281), .A2(n5802), .ZN(n6266) );
  INV_X1 U4039 ( .A(n6756), .ZN(n6847) );
  INV_X1 U4040 ( .A(n6744), .ZN(n6768) );
  OR2_X1 U4041 ( .A1(n6525), .A2(n6768), .ZN(n6825) );
  AND2_X1 U4042 ( .A1(n4738), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5053)
         );
  OAI211_X1 U4043 ( .C1(n5288), .C2(n5445), .A(n5641), .B(n5287), .ZN(n5442)
         );
  NOR2_X1 U4044 ( .A1(n4971), .A2(n5629), .ZN(n5197) );
  OR2_X1 U4045 ( .A1(n5140), .A2(n5094), .ZN(n5337) );
  AND2_X1 U4046 ( .A1(n5417), .A2(n7057), .ZN(n7266) );
  AND2_X1 U4047 ( .A1(n7125), .A2(n7057), .ZN(n7259) );
  AND2_X1 U4048 ( .A1(n3537), .A2(n3444), .ZN(n7114) );
  AND2_X1 U4049 ( .A1(n5630), .A2(n3445), .ZN(n7254) );
  OAI21_X1 U4050 ( .B1(n5004), .B2(n5003), .A(n5002), .ZN(n5373) );
  INV_X1 U4051 ( .A(n7108), .ZN(n7245) );
  OR2_X1 U4052 ( .A1(n5140), .A2(n5139), .ZN(n5396) );
  INV_X1 U4053 ( .A(n4953), .ZN(n5285) );
  INV_X1 U4054 ( .A(STATE_REG_0__SCAN_IN), .ZN(n7075) );
  OR2_X1 U4055 ( .A1(n7139), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6726) );
  INV_X1 U4056 ( .A(n6955), .ZN(n6981) );
  INV_X1 U4057 ( .A(n6930), .ZN(n6975) );
  OR2_X1 U4058 ( .A1(n5179), .A2(n5178), .ZN(n6961) );
  NAND2_X1 U4059 ( .A1(n5179), .A2(n5161), .ZN(n6973) );
  AND2_X1 U4060 ( .A1(n4523), .A2(n4522), .ZN(n4524) );
  AND2_X1 U4061 ( .A1(n4685), .A2(n3539), .ZN(n4686) );
  OR2_X1 U4062 ( .A1(n5910), .A2(n5925), .ZN(n6120) );
  INV_X1 U4063 ( .A(n6577), .ZN(n6608) );
  NAND2_X1 U4064 ( .A1(n4991), .A2(n4418), .ZN(n5277) );
  OR2_X1 U4065 ( .A1(n7139), .A2(n6733), .ZN(n6685) );
  OR2_X1 U4066 ( .A1(n6691), .A2(n4760), .ZN(n6707) );
  AND2_X1 U4067 ( .A1(n6778), .A2(n4905), .ZN(n6781) );
  INV_X1 U4068 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n7012) );
  NOR2_X1 U4069 ( .A1(n5206), .A2(n5205), .ZN(n5463) );
  INV_X1 U4070 ( .A(n5061), .ZN(n5326) );
  INV_X1 U4071 ( .A(n7129), .ZN(n7265) );
  NAND2_X1 U4072 ( .A1(DATAI_0_), .A2(n5285), .ZN(n7156) );
  NAND2_X1 U4073 ( .A1(DATAI_4_), .A2(n5285), .ZN(n7214) );
  INV_X1 U4074 ( .A(n6992), .ZN(n7051) );
  INV_X1 U4075 ( .A(n6656), .ZN(n6654) );
  NAND2_X1 U4076 ( .A1(n4712), .A2(n4711), .ZN(U2829) );
  NAND2_X1 U4077 ( .A1(n4687), .A2(n4686), .ZN(U2860) );
  OAI21_X1 U4078 ( .B1(n6230), .B2(n6993), .A(n4637), .ZN(U2957) );
  INV_X1 U4079 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6133) );
  INV_X1 U4080 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4301) );
  INV_X1 U4081 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4308) );
  INV_X1 U4082 ( .A(n4326), .ZN(n3542) );
  INV_X1 U4083 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3543) );
  XNOR2_X1 U4084 ( .A(n4638), .B(n3543), .ZN(n5863) );
  NOR2_X1 U4085 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3544) );
  INV_X1 U4086 ( .A(n3544), .ZN(n3690) );
  AOI22_X1 U4087 ( .A1(n3761), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3762), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3548) );
  AND2_X4 U4088 ( .A1(n3468), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n6555)
         );
  NOR2_X4 U4089 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4090 ( .A1(n3859), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3739), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3547) );
  AND2_X2 U4091 ( .A1(n6554), .A2(n3549), .ZN(n3767) );
  AND2_X4 U4092 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4790) );
  AOI22_X1 U4093 ( .A1(n3767), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4094 ( .A1(n3865), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3545) );
  NAND4_X1 U4095 ( .A1(n3548), .A2(n3547), .A3(n3546), .A4(n3545), .ZN(n3556)
         );
  AND2_X2 U4096 ( .A1(n3549), .A2(n4790), .ZN(n3769) );
  AOI22_X1 U4097 ( .A1(n3903), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4098 ( .A1(n3860), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4099 ( .A1(n3441), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3551) );
  NAND4_X1 U4100 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n3555)
         );
  OR2_X2 U4101 ( .A1(n3556), .A2(n3555), .ZN(n5837) );
  INV_X1 U4102 ( .A(EAX_REG_29__SCAN_IN), .ZN(n3693) );
  AOI22_X1 U4103 ( .A1(n4648), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4104 ( .A1(n4177), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4105 ( .A1(n4650), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4106 ( .A1(n3557), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3558) );
  NAND4_X1 U4107 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3567)
         );
  AOI22_X1 U4108 ( .A1(n3832), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4642), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4109 ( .A1(n3903), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4110 ( .A1(n3833), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4111 ( .A1(n3734), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3562) );
  NAND4_X1 U4112 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n3566)
         );
  NOR2_X1 U4113 ( .A1(n3567), .A2(n3566), .ZN(n4641) );
  AOI22_X1 U4114 ( .A1(n3832), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3571) );
  AOI22_X1 U4115 ( .A1(n3826), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3570) );
  AOI22_X1 U4116 ( .A1(n3833), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4117 ( .A1(n4650), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3568) );
  NAND4_X1 U4118 ( .A1(n3571), .A2(n3570), .A3(n3569), .A4(n3568), .ZN(n3577)
         );
  AOI22_X1 U4119 ( .A1(n4642), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4120 ( .A1(n4649), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4121 ( .A1(n3557), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3573) );
  AOI22_X1 U4122 ( .A1(n3734), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3572) );
  NAND4_X1 U4123 ( .A1(n3575), .A2(n3574), .A3(n3573), .A4(n3572), .ZN(n3576)
         );
  NOR2_X1 U4124 ( .A1(n3577), .A2(n3576), .ZN(n4328) );
  AOI22_X1 U4126 ( .A1(n4650), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3931), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4127 ( .A1(n4642), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4128 ( .A1(n3903), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4129 ( .A1(n4273), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3578) );
  NAND4_X1 U4130 ( .A1(n3581), .A2(n3580), .A3(n3579), .A4(n3578), .ZN(n3587)
         );
  AOI22_X1 U4131 ( .A1(n3832), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4132 ( .A1(n3833), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4133 ( .A1(n3835), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3583) );
  BUF_X1 U4134 ( .A(n3769), .Z(n4651) );
  AOI22_X1 U4135 ( .A1(n4177), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3582) );
  NAND4_X1 U4136 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3586)
         );
  NOR2_X1 U4137 ( .A1(n3587), .A2(n3586), .ZN(n4311) );
  AOI22_X1 U4138 ( .A1(n4642), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4139 ( .A1(n3826), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3590) );
  AOI22_X1 U4140 ( .A1(n3833), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3589) );
  AOI22_X1 U4141 ( .A1(n3557), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3588) );
  NAND4_X1 U4142 ( .A1(n3591), .A2(n3590), .A3(n3589), .A4(n3588), .ZN(n3597)
         );
  AOI22_X1 U4143 ( .A1(n3832), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4144 ( .A1(n4650), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4145 ( .A1(n3931), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4146 ( .A1(n4273), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3592) );
  NAND4_X1 U4147 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3596)
         );
  NOR2_X1 U4148 ( .A1(n3597), .A2(n3596), .ZN(n4288) );
  AOI22_X1 U4149 ( .A1(n3832), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4150 ( .A1(n3931), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4151 ( .A1(n4650), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4152 ( .A1(n3557), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3598) );
  NAND4_X1 U4153 ( .A1(n3601), .A2(n3600), .A3(n3599), .A4(n3598), .ZN(n3607)
         );
  AOI22_X1 U4154 ( .A1(n4642), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3605) );
  AOI22_X1 U4155 ( .A1(n3826), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3604) );
  AOI22_X1 U4156 ( .A1(n3833), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4157 ( .A1(n4649), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3602) );
  NAND4_X1 U4158 ( .A1(n3605), .A2(n3604), .A3(n3603), .A4(n3602), .ZN(n3606)
         );
  NOR2_X1 U4159 ( .A1(n3607), .A2(n3606), .ZN(n4289) );
  OR2_X1 U4160 ( .A1(n4288), .A2(n4289), .ZN(n4299) );
  AOI22_X1 U4161 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n3826), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4162 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n4642), .B1(n3832), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4163 ( .A1(n4648), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4164 ( .A1(n3833), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3608) );
  NAND4_X1 U4165 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3617)
         );
  AOI22_X1 U4166 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n3825), .B1(n3835), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4167 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n4649), .B1(n4651), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4168 ( .A1(n4650), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4169 ( .A1(n3931), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3612) );
  NAND4_X1 U4170 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3616)
         );
  NOR2_X1 U4171 ( .A1(n3617), .A2(n3616), .ZN(n4297) );
  NOR2_X1 U4172 ( .A1(n4311), .A2(n4310), .ZN(n4320) );
  AOI22_X1 U4173 ( .A1(n4642), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4174 ( .A1(n3832), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4175 ( .A1(n4650), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4176 ( .A1(n4273), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3618) );
  NAND4_X1 U4177 ( .A1(n3621), .A2(n3620), .A3(n3619), .A4(n3618), .ZN(n3627)
         );
  AOI22_X1 U4178 ( .A1(n3903), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4179 ( .A1(n3734), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4180 ( .A1(n4649), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4181 ( .A1(n3557), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3622) );
  NAND4_X1 U4182 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(n3626)
         );
  OR2_X1 U4183 ( .A1(n3627), .A2(n3626), .ZN(n4319) );
  NAND2_X1 U4184 ( .A1(n4320), .A2(n4319), .ZN(n4327) );
  NOR2_X1 U4185 ( .A1(n4328), .A2(n4327), .ZN(n4338) );
  AOI22_X1 U4186 ( .A1(n4642), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4187 ( .A1(n3832), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4188 ( .A1(n4650), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4189 ( .A1(n4273), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3628) );
  NAND4_X1 U4190 ( .A1(n3631), .A2(n3630), .A3(n3629), .A4(n3628), .ZN(n3637)
         );
  AOI22_X1 U4191 ( .A1(n3903), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4192 ( .A1(n3931), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4193 ( .A1(n4649), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4194 ( .A1(n3557), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3632) );
  NAND4_X1 U4195 ( .A1(n3635), .A2(n3634), .A3(n3633), .A4(n3632), .ZN(n3636)
         );
  OR2_X1 U4196 ( .A1(n3637), .A2(n3636), .ZN(n4339) );
  NAND2_X1 U4197 ( .A1(n4338), .A2(n4339), .ZN(n4640) );
  XOR2_X1 U4198 ( .A(n4641), .B(n4640), .Z(n3689) );
  AOI22_X1 U4199 ( .A1(n3865), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3440), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4200 ( .A1(n3739), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4201 ( .A1(n3903), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3761), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4202 ( .A1(n3859), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4203 ( .A1(n3441), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4204 ( .A1(n3767), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4205 ( .A1(n3834), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3642) );
  NAND2_X1 U4206 ( .A1(n3734), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3651)
         );
  NAND2_X1 U4207 ( .A1(n3739), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3650) );
  NAND2_X1 U4208 ( .A1(n3834), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3649) );
  NAND2_X1 U4209 ( .A1(n3827), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3648)
         );
  NAND2_X1 U4210 ( .A1(n3761), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3655) );
  NAND2_X1 U4211 ( .A1(n3762), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3654)
         );
  NAND2_X1 U4212 ( .A1(n3860), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3653) );
  NAND2_X1 U4213 ( .A1(n3865), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3652) );
  NAND2_X1 U4214 ( .A1(n3767), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3659) );
  NAND2_X1 U4215 ( .A1(n3903), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3658)
         );
  NAND2_X1 U4216 ( .A1(n3768), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3657) );
  NAND2_X1 U4217 ( .A1(n3769), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3656) );
  NAND2_X1 U4218 ( .A1(n3859), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3663) );
  NAND2_X1 U4219 ( .A1(n3441), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3662)
         );
  NAND2_X1 U4220 ( .A1(n3725), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3661)
         );
  NAND2_X1 U4221 ( .A1(n3442), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3660) );
  NAND3_X1 U4222 ( .A1(n3793), .A2(n5837), .A3(n3848), .ZN(n3815) );
  INV_X1 U4223 ( .A(n3815), .ZN(n3688) );
  NAND2_X1 U4224 ( .A1(n3761), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3671) );
  NAND2_X1 U4225 ( .A1(n3762), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3670)
         );
  NAND2_X1 U4226 ( .A1(n3860), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4227 ( .A1(n3865), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3668) );
  NAND2_X1 U4228 ( .A1(n3734), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3675)
         );
  NAND2_X1 U4229 ( .A1(n3739), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3674) );
  NAND2_X1 U4230 ( .A1(n3834), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3673) );
  NAND2_X1 U4231 ( .A1(n3827), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3672)
         );
  NAND2_X1 U4232 ( .A1(n3767), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3679) );
  NAND2_X1 U4233 ( .A1(n3903), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3678)
         );
  NAND2_X1 U4234 ( .A1(n3768), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3677) );
  NAND2_X1 U4235 ( .A1(n3769), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3676) );
  NAND2_X1 U4236 ( .A1(n3859), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3683) );
  NAND2_X1 U4237 ( .A1(n3866), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3682)
         );
  NAND2_X1 U4238 ( .A1(n3725), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3681)
         );
  NAND2_X1 U4239 ( .A1(n3442), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3680) );
  AND4_X1 U4240 ( .A1(n3683), .A2(n3682), .A3(n3681), .A4(n3680), .ZN(n3684)
         );
  NAND2_X1 U4241 ( .A1(n3688), .A2(n4867), .ZN(n3784) );
  INV_X1 U4242 ( .A(n3784), .ZN(n6553) );
  NAND2_X1 U4243 ( .A1(n3689), .A2(n4664), .ZN(n3692) );
  AOI21_X1 U4244 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n7128), .A(n4343), 
        .ZN(n3691) );
  OAI211_X1 U4245 ( .C1(n4662), .C2(n3693), .A(n3692), .B(n3691), .ZN(n3694)
         );
  OAI21_X1 U4246 ( .B1(n5863), .B2(n3690), .A(n3694), .ZN(n4345) );
  NAND2_X1 U4247 ( .A1(n3767), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3698) );
  NAND2_X1 U4248 ( .A1(n3903), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3697)
         );
  NAND2_X1 U4249 ( .A1(n3768), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3696) );
  NAND2_X1 U4250 ( .A1(n3865), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3702) );
  NAND2_X1 U4251 ( .A1(n3860), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3701) );
  NAND2_X1 U4252 ( .A1(n3866), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3700)
         );
  NAND2_X1 U4253 ( .A1(n3725), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3699)
         );
  NAND2_X1 U4254 ( .A1(n3859), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3706) );
  NAND2_X1 U4255 ( .A1(n3761), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3705) );
  NAND2_X1 U4256 ( .A1(n3762), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3704)
         );
  NAND2_X1 U4257 ( .A1(n3442), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3703) );
  NAND2_X1 U4258 ( .A1(n3734), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3710)
         );
  NAND2_X1 U4259 ( .A1(n3739), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3709) );
  NAND2_X1 U4260 ( .A1(n3834), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3708) );
  NAND2_X1 U4261 ( .A1(n3827), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3707)
         );
  INV_X2 U4262 ( .A(n3750), .ZN(n3785) );
  AOI22_X1 U4263 ( .A1(n3734), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3860), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4264 ( .A1(n3762), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4265 ( .A1(n3859), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4266 ( .A1(n3739), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4267 ( .A1(n3865), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3767), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3724) );
  AOI22_X1 U4268 ( .A1(n3903), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3834), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3723) );
  AOI22_X1 U4269 ( .A1(n3866), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3722) );
  AOI22_X1 U4270 ( .A1(n3761), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3721) );
  NAND2_X1 U4271 ( .A1(n3865), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3729) );
  NAND2_X1 U4272 ( .A1(n3859), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3728) );
  NAND2_X1 U4273 ( .A1(n3866), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3727)
         );
  NAND2_X1 U4274 ( .A1(n3725), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3726)
         );
  NAND2_X1 U4275 ( .A1(n3761), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3733) );
  NAND2_X1 U4276 ( .A1(n3762), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3732)
         );
  NAND2_X1 U4277 ( .A1(n3860), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3731) );
  NAND2_X1 U4278 ( .A1(n3442), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3730) );
  NAND2_X1 U4279 ( .A1(n3734), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3738)
         );
  NAND2_X1 U4280 ( .A1(n3903), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3737)
         );
  NAND2_X1 U4281 ( .A1(n3834), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3736) );
  NAND2_X1 U4282 ( .A1(n3827), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3735)
         );
  NAND2_X1 U4283 ( .A1(n3767), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3743) );
  NAND2_X1 U4284 ( .A1(n3739), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3742) );
  NAND2_X1 U4285 ( .A1(n3768), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3741) );
  NAND2_X1 U4286 ( .A1(n3769), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3740) );
  NAND4_X4 U4287 ( .A1(n3747), .A2(n3746), .A3(n3745), .A4(n3744), .ZN(n4418)
         );
  NAND2_X1 U4288 ( .A1(n7074), .A2(STATE_REG_1__SCAN_IN), .ZN(n7071) );
  INV_X1 U4289 ( .A(STATE_REG_1__SCAN_IN), .ZN(n3748) );
  NAND2_X1 U4290 ( .A1(n3748), .A2(STATE_REG_2__SCAN_IN), .ZN(n3749) );
  NAND2_X1 U4291 ( .A1(n7071), .A2(n3749), .ZN(n7067) );
  NAND2_X1 U4292 ( .A1(n3448), .A2(n3750), .ZN(n3751) );
  NAND4_X1 U4293 ( .A1(n3809), .A2(n3810), .A3(n4626), .A4(n3751), .ZN(n3780)
         );
  NAND2_X1 U4294 ( .A1(n3752), .A2(n4871), .ZN(n3792) );
  NAND2_X1 U4295 ( .A1(n3734), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3756)
         );
  NAND2_X1 U4296 ( .A1(n3739), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U4297 ( .A1(n3834), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3754) );
  NAND2_X1 U4298 ( .A1(n3827), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3753)
         );
  NAND2_X1 U4299 ( .A1(n3859), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3760) );
  NAND2_X1 U4300 ( .A1(n3441), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3759)
         );
  NAND2_X1 U4301 ( .A1(n3725), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3758)
         );
  NAND2_X1 U4302 ( .A1(n3442), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3757) );
  NAND2_X1 U4303 ( .A1(n3761), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3766) );
  NAND2_X1 U4304 ( .A1(n3762), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3765)
         );
  NAND2_X1 U4305 ( .A1(n3860), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3764) );
  NAND2_X1 U4306 ( .A1(n3865), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3763) );
  NAND2_X1 U4307 ( .A1(n3767), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3773) );
  NAND2_X1 U4308 ( .A1(n3903), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3772)
         );
  NAND2_X1 U4309 ( .A1(n3768), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3771) );
  NAND2_X1 U4310 ( .A1(n3769), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3770) );
  NAND2_X1 U4311 ( .A1(n3792), .A2(n4407), .ZN(n3779) );
  NAND2_X1 U4312 ( .A1(n4418), .A2(n4531), .ZN(n4405) );
  NAND2_X1 U4313 ( .A1(n3779), .A2(n4785), .ZN(n3812) );
  NOR2_X1 U4314 ( .A1(n3780), .A2(n3812), .ZN(n3787) );
  OAI21_X1 U4315 ( .B1(n4867), .B2(n3848), .A(n3785), .ZN(n3782) );
  NAND2_X1 U4316 ( .A1(n3782), .A2(n3854), .ZN(n3783) );
  NAND2_X1 U4317 ( .A1(n3787), .A2(n3820), .ZN(n3788) );
  NAND2_X1 U4318 ( .A1(n3788), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3892) );
  INV_X1 U4319 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U4320 ( .A1(n6560), .A2(n7046), .ZN(n4630) );
  NAND2_X1 U4321 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5060) );
  OAI21_X1 U4322 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n5060), .ZN(n5129) );
  OR2_X1 U4323 ( .A1(n4630), .A2(n5129), .ZN(n3790) );
  NAND2_X1 U4324 ( .A1(n3923), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3789) );
  OAI21_X1 U4325 ( .B1(n3892), .B2(n6552), .A(n3803), .ZN(n3791) );
  INV_X1 U4326 ( .A(n3791), .ZN(n3802) );
  NAND2_X1 U4327 ( .A1(n4410), .A2(n3794), .ZN(n4786) );
  INV_X1 U4328 ( .A(n4672), .ZN(n3797) );
  NOR2_X1 U4329 ( .A1(n4418), .A2(n4354), .ZN(n3796) );
  INV_X1 U4330 ( .A(n4867), .ZN(n3795) );
  INV_X1 U4331 ( .A(n3854), .ZN(n4412) );
  NAND2_X1 U4332 ( .A1(n3800), .A2(n4923), .ZN(n3806) );
  NAND2_X1 U4333 ( .A1(n3806), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3801) );
  INV_X1 U4334 ( .A(n3803), .ZN(n3804) );
  NOR2_X1 U4335 ( .A1(n3804), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3805)
         );
  NAND2_X1 U4336 ( .A1(n3806), .A2(n3536), .ZN(n3807) );
  MUX2_X1 U4337 ( .A(n4630), .B(n4417), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3808) );
  OAI21_X1 U4338 ( .B1(n3892), .B2(n3468), .A(n3808), .ZN(n3845) );
  NAND3_X1 U4339 ( .A1(n3809), .A2(n4531), .A3(n3810), .ZN(n3811) );
  NAND2_X1 U4340 ( .A1(n3811), .A2(n4418), .ZN(n3819) );
  NAND2_X1 U4341 ( .A1(n3813), .A2(n4407), .ZN(n3818) );
  NAND2_X1 U4342 ( .A1(n6560), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7034) );
  INV_X1 U4343 ( .A(n7034), .ZN(n3817) );
  INV_X1 U4344 ( .A(n3814), .ZN(n3816) );
  INV_X1 U4345 ( .A(n3433), .ZN(n3821) );
  OR2_X1 U4346 ( .A1(n4855), .A2(n4867), .ZN(n3822) );
  NAND2_X1 U4347 ( .A1(n4843), .A2(n7046), .ZN(n3844) );
  INV_X1 U4348 ( .A(n3898), .ZN(n3842) );
  AOI22_X1 U4349 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n3825), .B1(n4648), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3831) );
  BUF_X1 U4350 ( .A(n3903), .Z(n3826) );
  AOI22_X1 U4351 ( .A1(n3734), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3826), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4352 ( .A1(n4177), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4354 ( .A1(n4649), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3828) );
  NAND4_X1 U4355 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(n3841)
         );
  AOI22_X1 U4356 ( .A1(n3832), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3761), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4357 ( .A1(n4650), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3866), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4358 ( .A1(n3442), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4359 ( .A1(n3835), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3836) );
  NAND4_X1 U4360 ( .A1(n3839), .A2(n3838), .A3(n3837), .A4(n3836), .ZN(n3840)
         );
  NAND2_X1 U4361 ( .A1(n3842), .A2(n4526), .ZN(n3843) );
  NAND2_X1 U4362 ( .A1(n3844), .A2(n3843), .ZN(n3913) );
  INV_X1 U4363 ( .A(n3845), .ZN(n3847) );
  INV_X1 U4364 ( .A(n4526), .ZN(n3850) );
  NAND2_X1 U4365 ( .A1(n4389), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3849) );
  OAI211_X1 U4366 ( .C1(n3850), .C2(n3897), .A(n3849), .B(n3898), .ZN(n3851)
         );
  INV_X1 U4367 ( .A(n3851), .ZN(n3852) );
  INV_X1 U4368 ( .A(n3912), .ZN(n3853) );
  XNOR2_X1 U4369 ( .A(n3913), .B(n3853), .ZN(n4525) );
  NAND2_X1 U4370 ( .A1(n4525), .A2(n4154), .ZN(n3858) );
  AOI22_X1 U4371 ( .A1(n4668), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n7128), .ZN(n3856) );
  AND2_X1 U4372 ( .A1(n3854), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3884) );
  NAND2_X1 U4373 ( .A1(n3884), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3855) );
  AND2_X1 U4374 ( .A1(n3856), .A2(n3855), .ZN(n3857) );
  NAND2_X1 U4375 ( .A1(n3858), .A2(n3857), .ZN(n4831) );
  NAND2_X1 U4376 ( .A1(n4389), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3876) );
  NAND2_X1 U4377 ( .A1(n3898), .A2(n5169), .ZN(n3874) );
  AOI22_X1 U4378 ( .A1(n3859), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3734), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4379 ( .A1(n4648), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4380 ( .A1(n3826), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4381 ( .A1(n4273), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3725), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4382 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3873)
         );
  AOI22_X1 U4383 ( .A1(n3832), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3761), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4384 ( .A1(n3833), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4385 ( .A1(n3835), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4386 ( .A1(n4177), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3868) );
  NAND4_X1 U4387 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3872)
         );
  OR2_X1 U4388 ( .A1(n3873), .A2(n3872), .ZN(n4532) );
  NAND2_X1 U4389 ( .A1(n3874), .A2(n4532), .ZN(n3875) );
  NAND3_X1 U4390 ( .A1(n3876), .A2(n3875), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3877) );
  AND2_X1 U4391 ( .A1(n5837), .A2(n3793), .ZN(n3879) );
  AOI21_X1 U4392 ( .B1(n7057), .B2(n3879), .A(n7128), .ZN(n4718) );
  INV_X1 U4393 ( .A(n3884), .ZN(n3963) );
  NAND2_X1 U4394 ( .A1(n3443), .A2(n4154), .ZN(n3883) );
  AOI22_X1 U4395 ( .A1(n3881), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n7128), .ZN(n3882) );
  OAI211_X1 U4396 ( .C1(n3963), .C2(n3468), .A(n3883), .B(n3882), .ZN(n4717)
         );
  MUX2_X1 U4397 ( .A(n3544), .B(n4718), .S(n4717), .Z(n4830) );
  NAND2_X1 U4398 ( .A1(n4831), .A2(n4830), .ZN(n4822) );
  NAND2_X1 U4399 ( .A1(n3884), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3888) );
  INV_X1 U4400 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U4401 ( .A1(n7128), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4300) );
  NAND2_X1 U4402 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3940) );
  OAI21_X1 U4403 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3940), .ZN(n6690) );
  NAND2_X1 U4404 ( .A1(n3544), .A2(n6690), .ZN(n3885) );
  OAI21_X1 U4405 ( .B1(n5526), .B2(n4300), .A(n3885), .ZN(n3886) );
  AOI21_X1 U4406 ( .B1(n4668), .B2(EAX_REG_2__SCAN_IN), .A(n3886), .ZN(n3887)
         );
  AND2_X1 U4407 ( .A1(n3888), .A2(n3887), .ZN(n4823) );
  INV_X1 U4408 ( .A(n5060), .ZN(n3893) );
  NAND2_X1 U4409 ( .A1(n3893), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4844) );
  NAND2_X1 U4410 ( .A1(n5060), .A2(n7012), .ZN(n3894) );
  INV_X1 U4411 ( .A(n4630), .ZN(n3924) );
  AOI22_X1 U4412 ( .A1(n4877), .A2(n3924), .B1(n3923), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3895) );
  XNOR2_X1 U4413 ( .A(n3920), .B(n3919), .ZN(n4783) );
  NAND2_X1 U4414 ( .A1(n4783), .A2(n7046), .ZN(n3911) );
  AOI22_X1 U4415 ( .A1(n3832), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4416 ( .A1(n3734), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3739), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4417 ( .A1(n4177), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3768), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4418 ( .A1(n3833), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3899) );
  NAND4_X1 U4419 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n3909)
         );
  AOI22_X1 U4420 ( .A1(n4642), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4421 ( .A1(n4650), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4422 ( .A1(n3826), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4423 ( .A1(n3835), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3904) );
  NAND4_X1 U4424 ( .A1(n3907), .A2(n3906), .A3(n3905), .A4(n3904), .ZN(n3908)
         );
  AOI22_X1 U4425 ( .A1(n4397), .A2(n4545), .B1(n4389), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3910) );
  INV_X1 U4426 ( .A(n4154), .ZN(n3916) );
  OAI21_X2 U4427 ( .B1(n5208), .B2(n3916), .A(n4300), .ZN(n4826) );
  NAND2_X1 U4428 ( .A1(n4822), .A2(n4823), .ZN(n3917) );
  OAI21_X1 U4429 ( .B1(n3918), .B2(n4826), .A(n3917), .ZN(n4821) );
  NAND2_X1 U4430 ( .A1(n4844), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3922) );
  NAND3_X1 U4431 ( .A1(n5128), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5088) );
  INV_X1 U4432 ( .A(n5088), .ZN(n7151) );
  NAND2_X1 U4433 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7151), .ZN(n7141) );
  NAND2_X1 U4434 ( .A1(n3922), .A2(n7141), .ZN(n4998) );
  AOI22_X1 U4435 ( .A1(n4998), .A2(n3924), .B1(n3923), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4436 ( .A1(n4642), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4437 ( .A1(n3832), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4438 ( .A1(n4650), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4439 ( .A1(n4273), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3927) );
  NAND4_X1 U4440 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3937)
         );
  AOI22_X1 U4441 ( .A1(n3826), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4442 ( .A1(n3931), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4443 ( .A1(n4649), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4444 ( .A1(n3557), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4445 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3936)
         );
  AOI22_X1 U4446 ( .A1(n4397), .A2(n4554), .B1(n4389), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3938) );
  INV_X1 U4447 ( .A(n3964), .ZN(n3943) );
  INV_X1 U4448 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3941) );
  NAND2_X1 U4449 ( .A1(n3941), .A2(n3940), .ZN(n3942) );
  NAND2_X1 U4450 ( .A1(n3943), .A2(n3942), .ZN(n5518) );
  AOI22_X1 U4451 ( .A1(n5518), .A2(n3544), .B1(n4667), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3945) );
  NAND2_X1 U4452 ( .A1(n4668), .A2(EAX_REG_3__SCAN_IN), .ZN(n3944) );
  OAI211_X1 U4453 ( .C1(n3963), .C2(n3921), .A(n3945), .B(n3944), .ZN(n3946)
         );
  AOI21_X1 U4454 ( .B1(n4883), .B2(n4154), .A(n3946), .ZN(n4910) );
  AOI22_X1 U4455 ( .A1(n4642), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4456 ( .A1(n3832), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4457 ( .A1(n4650), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4458 ( .A1(n4273), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3949) );
  NAND4_X1 U4459 ( .A1(n3952), .A2(n3951), .A3(n3950), .A4(n3949), .ZN(n3958)
         );
  AOI22_X1 U4460 ( .A1(n3826), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4461 ( .A1(n3931), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4462 ( .A1(n4649), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4463 ( .A1(n3557), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3953) );
  NAND4_X1 U4464 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3957)
         );
  NAND2_X1 U4465 ( .A1(n4397), .A2(n4561), .ZN(n3960) );
  NAND2_X1 U4466 ( .A1(n4389), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3959) );
  NAND2_X1 U4467 ( .A1(n3960), .A2(n3959), .ZN(n3969) );
  XNOR2_X1 U4468 ( .A(n3971), .B(n3969), .ZN(n4553) );
  NAND2_X1 U4469 ( .A1(n4553), .A2(n4154), .ZN(n3968) );
  INV_X1 U4470 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4352) );
  NAND2_X1 U4471 ( .A1(n7128), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3962)
         );
  NAND2_X1 U4472 ( .A1(n4668), .A2(EAX_REG_4__SCAN_IN), .ZN(n3961) );
  OAI211_X1 U4473 ( .C1(n3963), .C2(n4352), .A(n3962), .B(n3961), .ZN(n3966)
         );
  OAI21_X1 U4474 ( .B1(n3964), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3984), 
        .ZN(n6857) );
  AND2_X1 U4475 ( .A1(n6857), .A2(n4343), .ZN(n3965) );
  AOI21_X1 U4476 ( .B1(n3966), .B2(n3690), .A(n3965), .ZN(n3967) );
  NAND2_X1 U4477 ( .A1(n3968), .A2(n3967), .ZN(n4836) );
  AOI22_X1 U4478 ( .A1(n3832), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4479 ( .A1(n3931), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4480 ( .A1(n4650), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3973) );
  AOI22_X1 U4481 ( .A1(n4649), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U4482 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3981)
         );
  AOI22_X1 U4483 ( .A1(n3826), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3979) );
  AOI22_X1 U4484 ( .A1(n4648), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4485 ( .A1(n4642), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4486 ( .A1(n3825), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3976) );
  NAND4_X1 U4487 ( .A1(n3979), .A2(n3978), .A3(n3977), .A4(n3976), .ZN(n3980)
         );
  NAND2_X1 U4488 ( .A1(n4397), .A2(n4564), .ZN(n3983) );
  NAND2_X1 U4489 ( .A1(n4389), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3982) );
  AND2_X1 U4490 ( .A1(n3984), .A2(n3987), .ZN(n3985) );
  OR2_X1 U4491 ( .A1(n3985), .A2(n4003), .ZN(n6868) );
  NAND2_X1 U4492 ( .A1(n6868), .A2(n4343), .ZN(n3986) );
  OAI21_X1 U4493 ( .B1(n3987), .B2(n4300), .A(n3986), .ZN(n3988) );
  AOI21_X1 U4494 ( .B1(n4668), .B2(EAX_REG_5__SCAN_IN), .A(n3988), .ZN(n3989)
         );
  AOI22_X1 U4495 ( .A1(n4642), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4496 ( .A1(n3832), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4497 ( .A1(n4650), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4498 ( .A1(n4273), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3991) );
  NAND4_X1 U4499 ( .A1(n3994), .A2(n3993), .A3(n3992), .A4(n3991), .ZN(n4000)
         );
  AOI22_X1 U4500 ( .A1(n3826), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4501 ( .A1(n3931), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4502 ( .A1(n4649), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4503 ( .A1(n3557), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3995) );
  NAND4_X1 U4504 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n3999)
         );
  NAND2_X1 U4505 ( .A1(n4397), .A2(n4585), .ZN(n4002) );
  NAND2_X1 U4506 ( .A1(n4389), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4001) );
  NAND2_X1 U4507 ( .A1(n4009), .A2(n4010), .ZN(n4574) );
  OR2_X1 U4508 ( .A1(n4003), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4004) );
  NAND2_X1 U4509 ( .A1(n4026), .A2(n4004), .ZN(n6885) );
  INV_X1 U4510 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6592) );
  INV_X1 U4511 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4005) );
  OAI22_X1 U4512 ( .A1(n4662), .A2(n6592), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4005), .ZN(n4006) );
  MUX2_X1 U4513 ( .A(n6885), .B(n4006), .S(n3690), .Z(n4007) );
  AOI22_X1 U4514 ( .A1(n4648), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4515 ( .A1(n3931), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4516 ( .A1(n3833), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4517 ( .A1(n3557), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4013) );
  NAND4_X1 U4518 ( .A1(n4016), .A2(n4015), .A3(n4014), .A4(n4013), .ZN(n4022)
         );
  AOI22_X1 U4519 ( .A1(n3832), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4642), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4520 ( .A1(n3826), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4521 ( .A1(n4650), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4522 ( .A1(n4649), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4017) );
  NAND4_X1 U4523 ( .A1(n4020), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(n4021)
         );
  NAND2_X1 U4524 ( .A1(n4397), .A2(n4595), .ZN(n4024) );
  NAND2_X1 U4525 ( .A1(n4389), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4023) );
  NAND2_X1 U4526 ( .A1(n4024), .A2(n4023), .ZN(n4025) );
  INV_X1 U4527 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4031) );
  NAND2_X1 U4528 ( .A1(n4026), .A2(n4028), .ZN(n4027) );
  NAND2_X1 U4529 ( .A1(n4045), .A2(n4027), .ZN(n6902) );
  NOR2_X1 U4530 ( .A1(n4300), .A2(n4028), .ZN(n4029) );
  AOI21_X1 U4531 ( .B1(n6902), .B2(n4343), .A(n4029), .ZN(n4030) );
  OAI21_X1 U4532 ( .B1(n4662), .B2(n4031), .A(n4030), .ZN(n4032) );
  NAND2_X1 U4533 ( .A1(n4034), .A2(n4033), .ZN(n5045) );
  AOI22_X1 U4534 ( .A1(n3832), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4535 ( .A1(n4650), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3826), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4536 ( .A1(n4273), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4537 ( .A1(n3557), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4035) );
  NAND4_X1 U4538 ( .A1(n4038), .A2(n4037), .A3(n4036), .A4(n4035), .ZN(n4044)
         );
  AOI22_X1 U4539 ( .A1(n4642), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4540 ( .A1(n3833), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4541 ( .A1(n4177), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4542 ( .A1(n3931), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4039) );
  NAND4_X1 U4543 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4043)
         );
  OAI21_X1 U4544 ( .B1(n4044), .B2(n4043), .A(n4154), .ZN(n4049) );
  NAND2_X1 U4545 ( .A1(n4668), .A2(EAX_REG_8__SCAN_IN), .ZN(n4048) );
  XNOR2_X1 U4546 ( .A(n4045), .B(n5505), .ZN(n5502) );
  NAND2_X1 U4547 ( .A1(n5502), .A2(n4343), .ZN(n4047) );
  NAND2_X1 U4548 ( .A1(n4667), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4046)
         );
  XOR2_X1 U4549 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n4050), .Z(n5551) );
  AOI22_X1 U4550 ( .A1(n4668), .A2(EAX_REG_9__SCAN_IN), .B1(n4667), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U4551 ( .A1(n3832), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U4552 ( .A1(n4650), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U4553 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n3835), .B1(n3557), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U4554 ( .A1(n3825), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4051) );
  NAND4_X1 U4555 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4060)
         );
  AOI22_X1 U4556 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n3931), .B1(n3826), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U4557 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n4642), .B1(n4643), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U4558 ( .A1(n4177), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U4559 ( .A1(n4649), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4055) );
  NAND4_X1 U4560 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(n4059)
         );
  OAI21_X1 U4561 ( .B1(n4060), .B2(n4059), .A(n4154), .ZN(n4061) );
  OAI211_X1 U4562 ( .C1(n5551), .C2(n3690), .A(n4062), .B(n4061), .ZN(n5305)
         );
  XNOR2_X1 U4563 ( .A(n4063), .B(n5541), .ZN(n5683) );
  NAND2_X1 U4564 ( .A1(n5683), .A2(n4343), .ZN(n4078) );
  AOI22_X1 U4565 ( .A1(n3832), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U4566 ( .A1(n3833), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U4567 ( .A1(n4650), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4568 ( .A1(n3557), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4064) );
  NAND4_X1 U4569 ( .A1(n4067), .A2(n4066), .A3(n4065), .A4(n4064), .ZN(n4073)
         );
  AOI22_X1 U4570 ( .A1(n4642), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U4571 ( .A1(n3826), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U4572 ( .A1(n4649), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4573 ( .A1(n3931), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4068) );
  NAND4_X1 U4574 ( .A1(n4071), .A2(n4070), .A3(n4069), .A4(n4068), .ZN(n4072)
         );
  OAI21_X1 U4575 ( .B1(n4073), .B2(n4072), .A(n4154), .ZN(n4076) );
  NAND2_X1 U4576 ( .A1(n3881), .A2(EAX_REG_10__SCAN_IN), .ZN(n4075) );
  NAND2_X1 U4577 ( .A1(n4667), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4074)
         );
  AND3_X1 U4578 ( .A1(n4076), .A2(n4075), .A3(n4074), .ZN(n4077) );
  NAND2_X1 U4579 ( .A1(n4078), .A2(n4077), .ZN(n5532) );
  XOR2_X1 U4580 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n4079), .Z(n6910) );
  AOI22_X1 U4581 ( .A1(n3881), .A2(EAX_REG_11__SCAN_IN), .B1(n4667), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U4582 ( .A1(n3931), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U4583 ( .A1(n3832), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U4584 ( .A1(n4650), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U4585 ( .A1(n3826), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4080) );
  NAND4_X1 U4586 ( .A1(n4083), .A2(n4082), .A3(n4081), .A4(n4080), .ZN(n4089)
         );
  AOI22_X1 U4587 ( .A1(n4642), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U4588 ( .A1(n3833), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U4589 ( .A1(n4177), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U4590 ( .A1(n3835), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4084) );
  NAND4_X1 U4591 ( .A1(n4087), .A2(n4086), .A3(n4085), .A4(n4084), .ZN(n4088)
         );
  OAI21_X1 U4592 ( .B1(n4089), .B2(n4088), .A(n4154), .ZN(n4090) );
  OAI211_X1 U4593 ( .C1(n6910), .C2(n3690), .A(n4091), .B(n4090), .ZN(n5563)
         );
  XNOR2_X1 U4594 ( .A(n4092), .B(n5624), .ZN(n5725) );
  INV_X1 U4595 ( .A(EAX_REG_12__SCAN_IN), .ZN(n4093) );
  OAI22_X1 U4596 ( .A1(n4662), .A2(n4093), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5624), .ZN(n4094) );
  NAND2_X1 U4597 ( .A1(n4094), .A2(n3690), .ZN(n4106) );
  AOI22_X1 U4598 ( .A1(n3832), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4642), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U4599 ( .A1(n4273), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U4600 ( .A1(n3931), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U4601 ( .A1(n3833), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4095) );
  NAND4_X1 U4602 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(n4104)
         );
  AOI22_X1 U4603 ( .A1(n4648), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U4604 ( .A1(n4650), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U4605 ( .A1(n3826), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U4606 ( .A1(n4177), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4099) );
  NAND4_X1 U4607 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4103)
         );
  OAI21_X1 U4608 ( .B1(n4104), .B2(n4103), .A(n4154), .ZN(n4105) );
  NAND2_X1 U4609 ( .A1(n4106), .A2(n4105), .ZN(n4107) );
  AOI21_X1 U4610 ( .B1(n5725), .B2(n3544), .A(n4107), .ZN(n5618) );
  INV_X1 U4611 ( .A(n5618), .ZN(n4120) );
  AOI22_X1 U4612 ( .A1(n3832), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U4613 ( .A1(n3833), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3826), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U4614 ( .A1(n3825), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U4615 ( .A1(n3557), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4108) );
  NAND4_X1 U4616 ( .A1(n4111), .A2(n4110), .A3(n4109), .A4(n4108), .ZN(n4117)
         );
  AOI22_X1 U4617 ( .A1(n4650), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U4618 ( .A1(n4177), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U4619 ( .A1(n4642), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U4620 ( .A1(n3931), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4112) );
  NAND4_X1 U4621 ( .A1(n4115), .A2(n4114), .A3(n4113), .A4(n4112), .ZN(n4116)
         );
  OR2_X1 U4622 ( .A1(n4117), .A2(n4116), .ZN(n4118) );
  NAND2_X1 U4623 ( .A1(n4154), .A2(n4118), .ZN(n4121) );
  INV_X1 U4624 ( .A(n4121), .ZN(n4119) );
  NAND2_X1 U4625 ( .A1(n4668), .A2(EAX_REG_13__SCAN_IN), .ZN(n4125) );
  OAI21_X1 U4626 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4123), .A(n4127), 
        .ZN(n6920) );
  AOI22_X1 U4627 ( .A1(n4343), .A2(n6920), .B1(n4667), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4124) );
  NAND2_X1 U4628 ( .A1(n4125), .A2(n4124), .ZN(n5707) );
  NAND2_X1 U4629 ( .A1(n5705), .A2(n5707), .ZN(n5706) );
  XOR2_X1 U4630 ( .A(n4128), .B(n4127), .Z(n6938) );
  NAND2_X1 U4631 ( .A1(n6938), .A2(n4343), .ZN(n4132) );
  INV_X1 U4632 ( .A(EAX_REG_14__SCAN_IN), .ZN(n4130) );
  INV_X1 U4633 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7126) );
  OAI21_X1 U4634 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n7126), .A(n7128), 
        .ZN(n4129) );
  OAI21_X1 U4635 ( .B1(n4662), .B2(n4130), .A(n4129), .ZN(n4131) );
  NAND2_X1 U4636 ( .A1(n4132), .A2(n4131), .ZN(n4144) );
  AOI22_X1 U4637 ( .A1(n3832), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U4638 ( .A1(n3833), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U4639 ( .A1(n4177), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4134) );
  AOI22_X1 U4640 ( .A1(n3826), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4133) );
  NAND4_X1 U4641 ( .A1(n4136), .A2(n4135), .A3(n4134), .A4(n4133), .ZN(n4142)
         );
  AOI22_X1 U4642 ( .A1(n4642), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U4643 ( .A1(n3931), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4139) );
  AOI22_X1 U4644 ( .A1(n3835), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U4645 ( .A1(n4650), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4137) );
  NAND4_X1 U4646 ( .A1(n4140), .A2(n4139), .A3(n4138), .A4(n4137), .ZN(n4141)
         );
  OAI21_X1 U4647 ( .B1(n4142), .B2(n4141), .A(n4154), .ZN(n4143) );
  NAND2_X1 U4648 ( .A1(n4144), .A2(n4143), .ZN(n5716) );
  XNOR2_X1 U4649 ( .A(n4145), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6199)
         );
  AOI22_X1 U4650 ( .A1(n3833), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U4651 ( .A1(n3826), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U4652 ( .A1(n3931), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U4653 ( .A1(n4177), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4146) );
  NAND4_X1 U4654 ( .A1(n4149), .A2(n4148), .A3(n4147), .A4(n4146), .ZN(n4156)
         );
  AOI22_X1 U4655 ( .A1(n4642), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U4656 ( .A1(n4649), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U4657 ( .A1(n3832), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U4658 ( .A1(n4650), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4150) );
  NAND4_X1 U4659 ( .A1(n4153), .A2(n4152), .A3(n4151), .A4(n4150), .ZN(n4155)
         );
  OAI21_X1 U4660 ( .B1(n4156), .B2(n4155), .A(n4154), .ZN(n4159) );
  NAND2_X1 U4661 ( .A1(n4668), .A2(EAX_REG_15__SCAN_IN), .ZN(n4158) );
  NAND2_X1 U4662 ( .A1(n4667), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4157)
         );
  NAND3_X1 U4663 ( .A1(n4159), .A2(n4158), .A3(n4157), .ZN(n4160) );
  AOI21_X1 U4664 ( .B1(n6199), .B2(n3544), .A(n4160), .ZN(n5730) );
  XOR2_X1 U4665 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n4162), .Z(n6949) );
  INV_X1 U4666 ( .A(n6949), .ZN(n6191) );
  AOI22_X1 U4667 ( .A1(n4642), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U4668 ( .A1(n4650), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U4669 ( .A1(n3833), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U4670 ( .A1(n3903), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4163) );
  NAND4_X1 U4671 ( .A1(n4166), .A2(n4165), .A3(n4164), .A4(n4163), .ZN(n4172)
         );
  AOI22_X1 U4672 ( .A1(n3931), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U4673 ( .A1(n3832), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U4674 ( .A1(n3557), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U4675 ( .A1(n4643), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4167) );
  NAND4_X1 U4676 ( .A1(n4170), .A2(n4169), .A3(n4168), .A4(n4167), .ZN(n4171)
         );
  NOR2_X1 U4677 ( .A1(n4172), .A2(n4171), .ZN(n4174) );
  AOI22_X1 U4678 ( .A1(n4668), .A2(EAX_REG_16__SCAN_IN), .B1(n4667), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4173) );
  OAI21_X1 U4679 ( .B1(n4323), .B2(n4174), .A(n4173), .ZN(n4175) );
  AOI21_X1 U4680 ( .B1(n6191), .B2(n3544), .A(n4175), .ZN(n6040) );
  XNOR2_X1 U4681 ( .A(n4176), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6182)
         );
  AOI22_X1 U4682 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n4650), .B1(n3833), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U4683 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n3826), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U4684 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n4649), .B1(n3835), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U4685 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n3557), .B1(n4651), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4178) );
  NAND4_X1 U4686 ( .A1(n4181), .A2(n4180), .A3(n4179), .A4(n4178), .ZN(n4187)
         );
  AOI22_X1 U4687 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n4642), .B1(n4648), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U4688 ( .A1(n3832), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4184) );
  AOI22_X1 U4689 ( .A1(n4273), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4183) );
  AOI22_X1 U4690 ( .A1(n3931), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4182) );
  NAND4_X1 U4691 ( .A1(n4185), .A2(n4184), .A3(n4183), .A4(n4182), .ZN(n4186)
         );
  OR2_X1 U4692 ( .A1(n4187), .A2(n4186), .ZN(n4191) );
  INV_X1 U4693 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4189) );
  NAND2_X1 U4694 ( .A1(n7128), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4188)
         );
  OAI211_X1 U4695 ( .C1(n4662), .C2(n4189), .A(n3690), .B(n4188), .ZN(n4190)
         );
  AOI21_X1 U4696 ( .B1(n4664), .B2(n4191), .A(n4190), .ZN(n4192) );
  AOI21_X1 U4697 ( .B1(n6182), .B2(n3544), .A(n4192), .ZN(n5777) );
  INV_X1 U4698 ( .A(n4193), .ZN(n4195) );
  INV_X1 U4699 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4194) );
  NAND2_X1 U4700 ( .A1(n4195), .A2(n4194), .ZN(n4196) );
  NAND2_X1 U4701 ( .A1(n4213), .A2(n4196), .ZN(n6966) );
  AOI22_X1 U4702 ( .A1(n4642), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U4703 ( .A1(n3832), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U4704 ( .A1(n4177), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U4705 ( .A1(n3931), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4197) );
  NAND4_X1 U4706 ( .A1(n4200), .A2(n4199), .A3(n4198), .A4(n4197), .ZN(n4206)
         );
  AOI22_X1 U4707 ( .A1(n3833), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U4708 ( .A1(n4650), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U4709 ( .A1(n3557), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U4710 ( .A1(n3903), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3867), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4201) );
  NAND4_X1 U4711 ( .A1(n4204), .A2(n4203), .A3(n4202), .A4(n4201), .ZN(n4205)
         );
  NOR2_X1 U4712 ( .A1(n4206), .A2(n4205), .ZN(n4209) );
  OAI21_X1 U4713 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n7126), .A(n7128), 
        .ZN(n4208) );
  NAND2_X1 U4714 ( .A1(n4668), .A2(EAX_REG_18__SCAN_IN), .ZN(n4207) );
  OAI211_X1 U4715 ( .C1(n4323), .C2(n4209), .A(n4208), .B(n4207), .ZN(n4210)
         );
  NAND2_X1 U4716 ( .A1(n4211), .A2(n4210), .ZN(n6030) );
  XNOR2_X1 U4717 ( .A(n4213), .B(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6168)
         );
  NAND2_X1 U4718 ( .A1(n6168), .A2(n4343), .ZN(n4228) );
  AOI22_X1 U4719 ( .A1(n4642), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4217) );
  AOI22_X1 U4720 ( .A1(n3832), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U4721 ( .A1(n4650), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4215) );
  AOI22_X1 U4722 ( .A1(n4273), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4214) );
  NAND4_X1 U4723 ( .A1(n4217), .A2(n4216), .A3(n4215), .A4(n4214), .ZN(n4223)
         );
  AOI22_X1 U4724 ( .A1(n3826), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U4725 ( .A1(n3931), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U4726 ( .A1(n4649), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U4727 ( .A1(n3557), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4218) );
  NAND4_X1 U4728 ( .A1(n4221), .A2(n4220), .A3(n4219), .A4(n4218), .ZN(n4222)
         );
  NOR2_X1 U4729 ( .A1(n4223), .A2(n4222), .ZN(n4226) );
  INV_X1 U4730 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6164) );
  AOI21_X1 U4731 ( .B1(n6164), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4224) );
  AOI21_X1 U4732 ( .B1(n4668), .B2(EAX_REG_19__SCAN_IN), .A(n4224), .ZN(n4225)
         );
  OAI21_X1 U4733 ( .B1(n4323), .B2(n4226), .A(n4225), .ZN(n4227) );
  NAND2_X1 U4734 ( .A1(n4228), .A2(n4227), .ZN(n5984) );
  INV_X1 U4735 ( .A(n4229), .ZN(n4231) );
  INV_X1 U4736 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4230) );
  NAND2_X1 U4737 ( .A1(n4231), .A2(n4230), .ZN(n4232) );
  NAND2_X1 U4738 ( .A1(n4249), .A2(n4232), .ZN(n6974) );
  AOI22_X1 U4739 ( .A1(n4642), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U4740 ( .A1(n3826), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U4741 ( .A1(n4649), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4234) );
  AOI22_X1 U4742 ( .A1(n3835), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4233) );
  NAND4_X1 U4743 ( .A1(n4236), .A2(n4235), .A3(n4234), .A4(n4233), .ZN(n4242)
         );
  AOI22_X1 U4744 ( .A1(n3832), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4240) );
  AOI22_X1 U4745 ( .A1(n3931), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4239) );
  AOI22_X1 U4746 ( .A1(n4650), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4238) );
  AOI22_X1 U4747 ( .A1(n3557), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4237) );
  NAND4_X1 U4748 ( .A1(n4240), .A2(n4239), .A3(n4238), .A4(n4237), .ZN(n4241)
         );
  NOR2_X1 U4749 ( .A1(n4242), .A2(n4241), .ZN(n4246) );
  NAND2_X1 U4750 ( .A1(n7128), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4243)
         );
  NAND2_X1 U4751 ( .A1(n3690), .A2(n4243), .ZN(n4244) );
  AOI21_X1 U4752 ( .B1(n3881), .B2(EAX_REG_20__SCAN_IN), .A(n4244), .ZN(n4245)
         );
  OAI21_X1 U4753 ( .B1(n4323), .B2(n4246), .A(n4245), .ZN(n4247) );
  XNOR2_X1 U4754 ( .A(n4249), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6153)
         );
  AOI22_X1 U4755 ( .A1(n3734), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4253) );
  AOI22_X1 U4756 ( .A1(n3826), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4252) );
  AOI22_X1 U4757 ( .A1(n4648), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U4758 ( .A1(n4650), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4250) );
  NAND4_X1 U4759 ( .A1(n4253), .A2(n4252), .A3(n4251), .A4(n4250), .ZN(n4259)
         );
  AOI22_X1 U4760 ( .A1(n3832), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4642), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4257) );
  AOI22_X1 U4761 ( .A1(n3825), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4256) );
  AOI22_X1 U4762 ( .A1(n3835), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4255) );
  AOI22_X1 U4763 ( .A1(n3557), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4254) );
  NAND4_X1 U4764 ( .A1(n4257), .A2(n4256), .A3(n4255), .A4(n4254), .ZN(n4258)
         );
  OR2_X1 U4765 ( .A1(n4259), .A2(n4258), .ZN(n4263) );
  INV_X1 U4766 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4261) );
  NAND2_X1 U4767 ( .A1(n7128), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4260)
         );
  OAI211_X1 U4768 ( .C1(n4662), .C2(n4261), .A(n3690), .B(n4260), .ZN(n4262)
         );
  AOI21_X1 U4769 ( .B1(n4664), .B2(n4263), .A(n4262), .ZN(n4264) );
  AOI21_X1 U4770 ( .B1(n6153), .B2(n3544), .A(n4264), .ZN(n5972) );
  INV_X1 U4771 ( .A(n4265), .ZN(n4267) );
  INV_X1 U4772 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4266) );
  NAND2_X1 U4773 ( .A1(n4267), .A2(n4266), .ZN(n4268) );
  NAND2_X1 U4774 ( .A1(n4287), .A2(n4268), .ZN(n6141) );
  AOI22_X1 U4775 ( .A1(n4642), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4648), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U4776 ( .A1(n3832), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3833), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U4777 ( .A1(n3734), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3903), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4270) );
  AOI22_X1 U4778 ( .A1(n4177), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3769), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4269) );
  NAND4_X1 U4779 ( .A1(n4272), .A2(n4271), .A3(n4270), .A4(n4269), .ZN(n4279)
         );
  AOI22_X1 U4780 ( .A1(n3835), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3557), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U4781 ( .A1(n3825), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U4782 ( .A1(n4650), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4643), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U4783 ( .A1(n4649), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4274) );
  NAND4_X1 U4784 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4278)
         );
  NOR2_X1 U4785 ( .A1(n4279), .A2(n4278), .ZN(n4283) );
  NAND2_X1 U4786 ( .A1(n7128), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4280)
         );
  NAND2_X1 U4787 ( .A1(n3690), .A2(n4280), .ZN(n4281) );
  AOI21_X1 U4788 ( .B1(n4668), .B2(EAX_REG_22__SCAN_IN), .A(n4281), .ZN(n4282)
         );
  OAI21_X1 U4789 ( .B1(n4323), .B2(n4283), .A(n4282), .ZN(n4284) );
  NAND2_X1 U4790 ( .A1(n4285), .A2(n4284), .ZN(n5953) );
  XNOR2_X1 U4791 ( .A(n4287), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6131)
         );
  NAND2_X1 U4792 ( .A1(n6131), .A2(n4343), .ZN(n4295) );
  XOR2_X1 U4793 ( .A(n4289), .B(n4288), .Z(n4290) );
  NAND2_X1 U4794 ( .A1(n4664), .A2(n4290), .ZN(n4293) );
  OAI21_X1 U4795 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6133), .A(n3690), .ZN(
        n4291) );
  AOI21_X1 U4796 ( .B1(n3881), .B2(EAX_REG_23__SCAN_IN), .A(n4291), .ZN(n4292)
         );
  NAND2_X1 U4797 ( .A1(n4293), .A2(n4292), .ZN(n4294) );
  NAND2_X1 U4798 ( .A1(n4295), .A2(n4294), .ZN(n5937) );
  XNOR2_X1 U4799 ( .A(n4296), .B(n4301), .ZN(n6122) );
  NAND2_X1 U4800 ( .A1(n6122), .A2(n4343), .ZN(n4306) );
  INV_X1 U4801 ( .A(n4297), .ZN(n4298) );
  XNOR2_X1 U4802 ( .A(n4299), .B(n4298), .ZN(n4304) );
  INV_X1 U4803 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4302) );
  OAI22_X1 U4804 ( .A1(n4662), .A2(n4302), .B1(n4301), .B2(n4300), .ZN(n4303)
         );
  AOI21_X1 U4805 ( .B1(n4304), .B2(n4664), .A(n4303), .ZN(n4305) );
  NAND2_X1 U4806 ( .A1(n4306), .A2(n4305), .ZN(n5924) );
  XNOR2_X1 U4807 ( .A(n4307), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5917)
         );
  NOR2_X1 U4808 ( .A1(n4308), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4309) );
  AOI211_X1 U4809 ( .C1(n4668), .C2(EAX_REG_25__SCAN_IN), .A(n4343), .B(n4309), 
        .ZN(n4314) );
  XOR2_X1 U4810 ( .A(n4311), .B(n4310), .Z(n4312) );
  NAND2_X1 U4811 ( .A1(n4312), .A2(n4664), .ZN(n4313) );
  AOI22_X1 U4812 ( .A1(n5917), .A2(n4343), .B1(n4314), .B2(n4313), .ZN(n5911)
         );
  INV_X1 U4813 ( .A(n4315), .ZN(n4317) );
  INV_X1 U4814 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4316) );
  NAND2_X1 U4815 ( .A1(n4317), .A2(n4316), .ZN(n4318) );
  NAND2_X1 U4816 ( .A1(n4326), .A2(n4318), .ZN(n6099) );
  XNOR2_X1 U4817 ( .A(n4320), .B(n4319), .ZN(n4324) );
  OAI21_X1 U4818 ( .B1(n7126), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n7128), 
        .ZN(n4322) );
  NAND2_X1 U4819 ( .A1(n3881), .A2(EAX_REG_26__SCAN_IN), .ZN(n4321) );
  OAI211_X1 U4820 ( .C1(n4324), .C2(n4323), .A(n4322), .B(n4321), .ZN(n4325)
         );
  XNOR2_X1 U4821 ( .A(n4326), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5888)
         );
  XOR2_X1 U4822 ( .A(n4328), .B(n4327), .Z(n4332) );
  INV_X1 U4823 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4330) );
  NAND2_X1 U4824 ( .A1(n7128), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4329)
         );
  OAI211_X1 U4825 ( .C1(n4662), .C2(n4330), .A(n3690), .B(n4329), .ZN(n4331)
         );
  AOI21_X1 U4826 ( .B1(n4332), .B2(n4664), .A(n4331), .ZN(n4333) );
  AOI21_X1 U4827 ( .B1(n5888), .B2(n3544), .A(n4333), .ZN(n5881) );
  INV_X1 U4828 ( .A(n4334), .ZN(n4335) );
  INV_X1 U4829 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U4830 ( .A1(n4335), .A2(n5874), .ZN(n4336) );
  NOR2_X1 U4831 ( .A1(n5874), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4337) );
  AOI211_X1 U4832 ( .C1(n4668), .C2(EAX_REG_28__SCAN_IN), .A(n4343), .B(n4337), 
        .ZN(n4342) );
  XOR2_X1 U4833 ( .A(n4339), .B(n4338), .Z(n4340) );
  NAND2_X1 U4834 ( .A1(n4340), .A2(n4664), .ZN(n4341) );
  AOI22_X1 U4835 ( .A1(n6081), .A2(n4343), .B1(n4342), .B2(n4341), .ZN(n5873)
         );
  INV_X1 U4836 ( .A(n4636), .ZN(n6051) );
  XNOR2_X1 U4837 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4356) );
  NAND2_X1 U4838 ( .A1(n4356), .A2(n4355), .ZN(n4347) );
  NAND2_X1 U4839 ( .A1(n7008), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4346) );
  NAND2_X1 U4840 ( .A1(n4347), .A2(n4346), .ZN(n4368) );
  XNOR2_X1 U4841 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4367) );
  NAND2_X1 U4842 ( .A1(n4368), .A2(n4367), .ZN(n4349) );
  NAND2_X1 U4843 ( .A1(n7012), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4348) );
  NAND2_X1 U4844 ( .A1(n4349), .A2(n4348), .ZN(n4376) );
  XNOR2_X1 U4845 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4375) );
  NAND2_X1 U4846 ( .A1(n4376), .A2(n4375), .ZN(n4351) );
  NAND2_X1 U4847 ( .A1(n5128), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4350) );
  NAND2_X1 U4848 ( .A1(n4351), .A2(n4350), .ZN(n4394) );
  NAND2_X1 U4849 ( .A1(n4397), .A2(n4418), .ZN(n4358) );
  XNOR2_X1 U4850 ( .A(n4356), .B(n4355), .ZN(n4674) );
  NAND2_X1 U4851 ( .A1(n4389), .A2(n4674), .ZN(n4357) );
  NAND3_X1 U4852 ( .A1(n4358), .A2(n4357), .A3(n4354), .ZN(n4372) );
  NOR2_X1 U4853 ( .A1(n4674), .A2(n7046), .ZN(n4384) );
  OAI21_X1 U4854 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7123), .A(n4359), 
        .ZN(n4360) );
  INV_X1 U4855 ( .A(n4360), .ZN(n4362) );
  OAI211_X1 U4856 ( .C1(n4372), .C2(n4384), .A(n4362), .B(n4397), .ZN(n4361)
         );
  NAND2_X1 U4857 ( .A1(n4361), .A2(n4401), .ZN(n4366) );
  AOI21_X1 U4858 ( .B1(n4627), .B2(n4362), .A(n4855), .ZN(n4364) );
  NAND2_X1 U4859 ( .A1(n5184), .A2(n4855), .ZN(n6714) );
  NAND2_X1 U4860 ( .A1(n5184), .A2(n4354), .ZN(n4363) );
  NAND2_X1 U4861 ( .A1(n6714), .A2(n4363), .ZN(n4373) );
  OR2_X1 U4862 ( .A1(n4364), .A2(n4373), .ZN(n4365) );
  NAND2_X1 U4863 ( .A1(n4366), .A2(n4365), .ZN(n4371) );
  XNOR2_X1 U4864 ( .A(n4368), .B(n4367), .ZN(n4673) );
  INV_X1 U4865 ( .A(n4673), .ZN(n4369) );
  NAND2_X1 U4866 ( .A1(n4374), .A2(n4373), .ZN(n4370) );
  NAND2_X1 U4867 ( .A1(n4371), .A2(n4370), .ZN(n4383) );
  NOR2_X1 U4868 ( .A1(n4383), .A2(n4372), .ZN(n4382) );
  INV_X1 U4869 ( .A(n4373), .ZN(n4378) );
  INV_X1 U4870 ( .A(n4374), .ZN(n4377) );
  XNOR2_X1 U4871 ( .A(n4376), .B(n4375), .ZN(n4675) );
  AOI21_X1 U4872 ( .B1(n4378), .B2(n4377), .A(n4675), .ZN(n4379) );
  AOI21_X1 U4873 ( .B1(n4389), .B2(n4673), .A(n4379), .ZN(n4381) );
  INV_X1 U4874 ( .A(n4675), .ZN(n4380) );
  OAI22_X1 U4875 ( .A1(n4382), .A2(n4381), .B1(n4380), .B2(n4401), .ZN(n4388)
         );
  INV_X1 U4876 ( .A(n4383), .ZN(n4386) );
  INV_X1 U4877 ( .A(n4384), .ZN(n4385) );
  NAND3_X1 U4878 ( .A1(n4386), .A2(n4401), .A3(n4385), .ZN(n4387) );
  OAI211_X1 U4879 ( .C1(n4389), .C2(n4678), .A(n4388), .B(n4387), .ZN(n4390)
         );
  OAI21_X1 U4880 ( .B1(n4678), .B2(n4401), .A(n4390), .ZN(n4391) );
  AOI21_X1 U4881 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7046), .A(n4391), 
        .ZN(n4399) );
  NAND2_X1 U4882 ( .A1(n4392), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4396) );
  NAND2_X1 U4883 ( .A1(n4394), .A2(n4393), .ZN(n4395) );
  NAND2_X1 U4884 ( .A1(n4396), .A2(n4395), .ZN(n4677) );
  NAND2_X1 U4885 ( .A1(n4397), .A2(n4677), .ZN(n4398) );
  NAND2_X1 U4886 ( .A1(n4399), .A2(n4398), .ZN(n4403) );
  INV_X1 U4887 ( .A(n4677), .ZN(n4400) );
  NOR2_X1 U4888 ( .A1(n3784), .A2(n5184), .ZN(n4740) );
  NAND2_X1 U4889 ( .A1(n6988), .A2(n4740), .ZN(n4729) );
  INV_X1 U4890 ( .A(n4406), .ZN(n4408) );
  AOI21_X1 U4891 ( .B1(n4408), .B2(n5169), .A(n4407), .ZN(n4409) );
  OR2_X1 U4892 ( .A1(n4410), .A2(n4409), .ZN(n4726) );
  NAND2_X1 U4893 ( .A1(n4863), .A2(n5169), .ZN(n4439) );
  INV_X1 U4894 ( .A(n5844), .ZN(n4411) );
  NAND2_X1 U4895 ( .A1(n4855), .A2(n4418), .ZN(n5173) );
  OR2_X1 U4896 ( .A1(n5173), .A2(n3795), .ZN(n4777) );
  NAND2_X1 U4897 ( .A1(n4411), .A2(n4777), .ZN(n4414) );
  INV_X1 U4898 ( .A(n4626), .ZN(n4413) );
  AOI22_X1 U4899 ( .A1(n4414), .A2(n4413), .B1(n4412), .B2(n3795), .ZN(n4415)
         );
  OAI211_X1 U4900 ( .C1(n3809), .C2(n4490), .A(n4726), .B(n4415), .ZN(n4748)
         );
  NOR2_X1 U4901 ( .A1(n4748), .A2(n4680), .ZN(n4416) );
  NAND2_X1 U4902 ( .A1(n3431), .A2(n4416), .ZN(n4784) );
  INV_X1 U4903 ( .A(n5837), .ZN(n5028) );
  NAND4_X1 U4904 ( .A1(n5028), .A2(n4871), .A3(n6992), .A4(n3428), .ZN(n4681)
         );
  NAND4_X1 U4905 ( .A1(n4833), .A2(n3750), .A3(n4867), .A4(n4863), .ZN(n4419)
         );
  INV_X1 U4906 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U4907 ( .A1(n4439), .A2(n5052), .ZN(n4423) );
  INV_X1 U4908 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4421) );
  NAND2_X1 U4909 ( .A1(n4833), .A2(n4421), .ZN(n4422) );
  NAND3_X1 U4910 ( .A1(n4423), .A2(n4490), .A3(n4422), .ZN(n4424) );
  NAND2_X1 U4911 ( .A1(n4439), .A2(EBX_REG_0__SCAN_IN), .ZN(n4428) );
  INV_X1 U4912 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U4913 ( .A1(n4490), .A2(n4426), .ZN(n4427) );
  NAND2_X1 U4914 ( .A1(n4428), .A2(n4427), .ZN(n4715) );
  XNOR2_X1 U4915 ( .A(n4429), .B(n4715), .ZN(n5177) );
  NAND2_X1 U4916 ( .A1(n5177), .A2(n4833), .ZN(n4430) );
  OR2_X1 U4917 ( .A1(n4431), .A2(EBX_REG_2__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U4918 ( .A1(n4439), .A2(n4542), .ZN(n4434) );
  INV_X1 U4919 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4432) );
  NAND2_X1 U4920 ( .A1(n4833), .A2(n4432), .ZN(n4433) );
  NAND3_X1 U4921 ( .A1(n4434), .A2(n4490), .A3(n4433), .ZN(n4435) );
  NAND2_X1 U4922 ( .A1(n4436), .A2(n4435), .ZN(n4812) );
  MUX2_X1 U4923 ( .A(n4513), .B(n4490), .S(EBX_REG_3__SCAN_IN), .Z(n4438) );
  OR2_X1 U4924 ( .A1(n5844), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4437)
         );
  AND2_X1 U4925 ( .A1(n4438), .A2(n4437), .ZN(n4912) );
  OR2_X1 U4926 ( .A1(n4431), .A2(EBX_REG_4__SCAN_IN), .ZN(n4444) );
  INV_X1 U4927 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U4928 ( .A1(n4439), .A2(n4904), .ZN(n4442) );
  INV_X1 U4929 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4440) );
  NAND2_X1 U4930 ( .A1(n4833), .A2(n4440), .ZN(n4441) );
  NAND3_X1 U4931 ( .A1(n4442), .A2(n4490), .A3(n4441), .ZN(n4443) );
  MUX2_X1 U4932 ( .A(n4513), .B(n4490), .S(EBX_REG_5__SCAN_IN), .Z(n4446) );
  OAI21_X1 U4933 ( .B1(n5844), .B2(INSTADDRPOINTER_REG_5__SCAN_IN), .A(n4446), 
        .ZN(n4770) );
  OR2_X1 U4934 ( .A1(n4431), .A2(EBX_REG_6__SCAN_IN), .ZN(n4450) );
  INV_X1 U4935 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U4936 ( .A1(n4439), .A2(n6773), .ZN(n4448) );
  INV_X1 U4937 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6882) );
  NAND2_X1 U4938 ( .A1(n4833), .A2(n6882), .ZN(n4447) );
  NAND3_X1 U4939 ( .A1(n4448), .A2(n4490), .A3(n4447), .ZN(n4449) );
  NAND2_X1 U4940 ( .A1(n4450), .A2(n4449), .ZN(n5023) );
  INV_X1 U4941 ( .A(n4513), .ZN(n4489) );
  INV_X1 U4942 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4451) );
  NAND2_X1 U4943 ( .A1(n4489), .A2(n4451), .ZN(n4454) );
  NAND2_X1 U4944 ( .A1(n4490), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4452)
         );
  OAI211_X1 U4945 ( .C1(n5843), .C2(EBX_REG_7__SCAN_IN), .A(n4439), .B(n4452), 
        .ZN(n4453) );
  OR2_X1 U4946 ( .A1(n4431), .A2(EBX_REG_8__SCAN_IN), .ZN(n4459) );
  INV_X1 U4947 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U4948 ( .A1(n4439), .A2(n4598), .ZN(n4457) );
  INV_X1 U4949 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4455) );
  NAND2_X1 U4950 ( .A1(n4833), .A2(n4455), .ZN(n4456) );
  NAND3_X1 U4951 ( .A1(n4457), .A2(n4490), .A3(n4456), .ZN(n4458) );
  NAND2_X1 U4952 ( .A1(n4490), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4460)
         );
  OAI211_X1 U4953 ( .C1(n5843), .C2(EBX_REG_9__SCAN_IN), .A(n4439), .B(n4460), 
        .ZN(n4461) );
  OAI21_X1 U4954 ( .B1(n4513), .B2(EBX_REG_9__SCAN_IN), .A(n4461), .ZN(n5307)
         );
  OR2_X1 U4955 ( .A1(n4431), .A2(EBX_REG_10__SCAN_IN), .ZN(n4465) );
  INV_X1 U4956 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6807) );
  NAND2_X1 U4957 ( .A1(n4439), .A2(n6807), .ZN(n4463) );
  INV_X1 U4958 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U4959 ( .A1(n4833), .A2(n5538), .ZN(n4462) );
  NAND3_X1 U4960 ( .A1(n4463), .A2(n4490), .A3(n4462), .ZN(n4464) );
  NAND2_X1 U4961 ( .A1(n4465), .A2(n4464), .ZN(n5535) );
  MUX2_X1 U4962 ( .A(n4513), .B(n4490), .S(EBX_REG_11__SCAN_IN), .Z(n4466) );
  OAI21_X1 U4963 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5844), .A(n4466), 
        .ZN(n5566) );
  MUX2_X1 U4964 ( .A(n4513), .B(n4490), .S(EBX_REG_13__SCAN_IN), .Z(n4467) );
  OAI21_X1 U4965 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5844), .A(n4467), 
        .ZN(n4468) );
  INV_X1 U4966 ( .A(n4468), .ZN(n5708) );
  OR2_X1 U4967 ( .A1(n4431), .A2(EBX_REG_12__SCAN_IN), .ZN(n4472) );
  NAND2_X1 U4968 ( .A1(n4490), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4469) );
  NAND2_X1 U4969 ( .A1(n4439), .A2(n4469), .ZN(n4470) );
  OAI21_X1 U4970 ( .B1(EBX_REG_12__SCAN_IN), .B2(n5843), .A(n4470), .ZN(n4471)
         );
  NAND2_X1 U4971 ( .A1(n4472), .A2(n4471), .ZN(n5709) );
  NAND2_X1 U4972 ( .A1(n5708), .A2(n5709), .ZN(n4473) );
  OR2_X1 U4973 ( .A1(n4431), .A2(EBX_REG_14__SCAN_IN), .ZN(n4477) );
  INV_X1 U4974 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U4975 ( .A1(n4439), .A2(n5769), .ZN(n4475) );
  INV_X1 U4976 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U4977 ( .A1(n4833), .A2(n6934), .ZN(n4474) );
  NAND3_X1 U4978 ( .A1(n4475), .A2(n4490), .A3(n4474), .ZN(n4476) );
  MUX2_X1 U4979 ( .A(n4513), .B(n4490), .S(EBX_REG_15__SCAN_IN), .Z(n4479) );
  OR2_X1 U4980 ( .A1(n5844), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4478)
         );
  OR2_X1 U4981 ( .A1(n4431), .A2(EBX_REG_16__SCAN_IN), .ZN(n4483) );
  NAND2_X1 U4982 ( .A1(n4490), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4480) );
  NAND2_X1 U4983 ( .A1(n4439), .A2(n4480), .ZN(n4481) );
  OAI21_X1 U4984 ( .B1(EBX_REG_16__SCAN_IN), .B2(n5843), .A(n4481), .ZN(n4482)
         );
  NAND2_X1 U4985 ( .A1(n4483), .A2(n4482), .ZN(n6041) );
  MUX2_X1 U4986 ( .A(n4513), .B(n4490), .S(EBX_REG_17__SCAN_IN), .Z(n4484) );
  OAI21_X1 U4987 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5844), .A(n4484), 
        .ZN(n5778) );
  OR2_X1 U4988 ( .A1(n4431), .A2(EBX_REG_18__SCAN_IN), .ZN(n4488) );
  INV_X1 U4989 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U4990 ( .A1(n4439), .A2(n6537), .ZN(n4486) );
  INV_X1 U4991 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U4992 ( .A1(n4833), .A2(n6035), .ZN(n4485) );
  NAND3_X1 U4993 ( .A1(n4486), .A2(n4490), .A3(n4485), .ZN(n4487) );
  INV_X1 U4994 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U4995 ( .A1(n4489), .A2(n6026), .ZN(n4493) );
  NAND2_X1 U4996 ( .A1(n4490), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4491) );
  OAI211_X1 U4997 ( .C1(n5843), .C2(EBX_REG_19__SCAN_IN), .A(n4439), .B(n4491), 
        .ZN(n4492) );
  AND2_X1 U4998 ( .A1(n4493), .A2(n4492), .ZN(n5987) );
  OR2_X1 U4999 ( .A1(n4431), .A2(EBX_REG_20__SCAN_IN), .ZN(n4497) );
  NAND2_X1 U5000 ( .A1(n4490), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4494) );
  NAND2_X1 U5001 ( .A1(n4439), .A2(n4494), .ZN(n4495) );
  OAI21_X1 U5002 ( .B1(EBX_REG_20__SCAN_IN), .B2(n5843), .A(n4495), .ZN(n4496)
         );
  NAND2_X1 U5003 ( .A1(n4497), .A2(n4496), .ZN(n6021) );
  NAND2_X1 U5004 ( .A1(n4490), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4498) );
  OAI211_X1 U5005 ( .C1(n5843), .C2(EBX_REG_21__SCAN_IN), .A(n4439), .B(n4498), 
        .ZN(n4499) );
  OAI21_X1 U5006 ( .B1(n4513), .B2(EBX_REG_21__SCAN_IN), .A(n4499), .ZN(n5973)
         );
  OR2_X1 U5007 ( .A1(n4431), .A2(EBX_REG_22__SCAN_IN), .ZN(n4502) );
  INV_X1 U5008 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U5009 ( .A1(n4439), .A2(n6289), .ZN(n4500) );
  OAI211_X1 U5010 ( .C1(EBX_REG_22__SCAN_IN), .C2(n5843), .A(n4500), .B(n4490), 
        .ZN(n4501) );
  AND2_X1 U5011 ( .A1(n4502), .A2(n4501), .ZN(n5954) );
  MUX2_X1 U5012 ( .A(n4513), .B(n4490), .S(EBX_REG_23__SCAN_IN), .Z(n4503) );
  OAI21_X1 U5013 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5844), .A(n4503), 
        .ZN(n5938) );
  OR2_X1 U5014 ( .A1(n4431), .A2(EBX_REG_24__SCAN_IN), .ZN(n4506) );
  INV_X1 U5015 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U5016 ( .A1(n4439), .A2(n6269), .ZN(n4504) );
  OAI211_X1 U5017 ( .C1(EBX_REG_24__SCAN_IN), .C2(n5843), .A(n4504), .B(n4490), 
        .ZN(n4505) );
  AND2_X1 U5018 ( .A1(n4506), .A2(n4505), .ZN(n5933) );
  MUX2_X1 U5019 ( .A(n4513), .B(n4490), .S(EBX_REG_25__SCAN_IN), .Z(n4508) );
  OR2_X1 U5020 ( .A1(n5844), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4507)
         );
  NAND2_X1 U5021 ( .A1(n4508), .A2(n4507), .ZN(n5914) );
  NOR2_X1 U5022 ( .A1(n5933), .A2(n5914), .ZN(n4509) );
  OR2_X1 U5023 ( .A1(n4431), .A2(EBX_REG_26__SCAN_IN), .ZN(n4512) );
  INV_X1 U5024 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U5025 ( .A1(n4439), .A2(n6252), .ZN(n4510) );
  OAI211_X1 U5026 ( .C1(EBX_REG_26__SCAN_IN), .C2(n5843), .A(n4510), .B(n4490), 
        .ZN(n4511) );
  NAND2_X1 U5027 ( .A1(n4512), .A2(n4511), .ZN(n5901) );
  MUX2_X1 U5028 ( .A(n4513), .B(n4490), .S(EBX_REG_27__SCAN_IN), .Z(n4514) );
  OAI21_X1 U5029 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5844), .A(n4514), 
        .ZN(n5885) );
  OR2_X1 U5030 ( .A1(n4431), .A2(EBX_REG_28__SCAN_IN), .ZN(n4517) );
  INV_X1 U5031 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4621) );
  NAND2_X1 U5032 ( .A1(n4439), .A2(n4621), .ZN(n4515) );
  OAI211_X1 U5033 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5843), .A(n4515), .B(n4490), 
        .ZN(n4516) );
  AND2_X1 U5034 ( .A1(n4517), .A2(n4516), .ZN(n5869) );
  OR2_X1 U5035 ( .A1(n5844), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4519)
         );
  INV_X1 U5036 ( .A(EBX_REG_29__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U5037 ( .A1(n4833), .A2(n4521), .ZN(n4518) );
  NAND2_X1 U5038 ( .A1(n4519), .A2(n4518), .ZN(n4706) );
  OAI22_X1 U5039 ( .A1(n4706), .A2(n4705), .B1(EBX_REG_29__SCAN_IN), .B2(n4431), .ZN(n4520) );
  NAND2_X1 U5040 ( .A1(n5870), .A2(n4520), .ZN(n5847) );
  OAI21_X1 U5041 ( .B1(n5870), .B2(n4520), .A(n5847), .ZN(n5861) );
  NAND2_X1 U5042 ( .A1(n6012), .A2(EBX_REG_29__SCAN_IN), .ZN(n4522) );
  NAND2_X1 U5043 ( .A1(n4525), .A2(n4572), .ZN(n4530) );
  NAND2_X1 U5044 ( .A1(n4526), .A2(n4532), .ZN(n4547) );
  OAI21_X1 U5045 ( .B1(n4532), .B2(n4526), .A(n4547), .ZN(n4527) );
  INV_X1 U5046 ( .A(n4407), .ZN(n4753) );
  OAI211_X1 U5047 ( .C1(n4527), .C2(n4753), .A(n4626), .B(n4354), .ZN(n4528)
         );
  INV_X1 U5048 ( .A(n4528), .ZN(n4529) );
  INV_X1 U5049 ( .A(n4572), .ZN(n4582) );
  NAND2_X1 U5050 ( .A1(n4855), .A2(n4531), .ZN(n4538) );
  OAI21_X1 U5051 ( .B1(n4753), .B2(n4532), .A(n4538), .ZN(n4533) );
  INV_X1 U5052 ( .A(n4533), .ZN(n4534) );
  NAND2_X1 U5053 ( .A1(n4535), .A2(n4534), .ZN(n4738) );
  NAND2_X1 U5054 ( .A1(n5055), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4536)
         );
  NAND2_X1 U5055 ( .A1(n4537), .A2(n4536), .ZN(n4541) );
  NAND2_X1 U5056 ( .A1(n4541), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4808)
         );
  XNOR2_X1 U5057 ( .A(n4547), .B(n4545), .ZN(n4539) );
  OAI21_X1 U5058 ( .B1(n4539), .B2(n4753), .A(n4538), .ZN(n4540) );
  NAND2_X1 U5059 ( .A1(n4808), .A2(n4811), .ZN(n4544) );
  NAND2_X1 U5060 ( .A1(n4544), .A2(n4809), .ZN(n4551) );
  NAND2_X1 U5061 ( .A1(n3437), .A2(n4544), .ZN(n5032) );
  INV_X1 U5062 ( .A(n4545), .ZN(n4546) );
  NAND2_X1 U5063 ( .A1(n4547), .A2(n4546), .ZN(n4555) );
  INV_X1 U5064 ( .A(n4554), .ZN(n4548) );
  XNOR2_X1 U5065 ( .A(n4555), .B(n4548), .ZN(n4549) );
  AND2_X1 U5066 ( .A1(n4549), .A2(n4407), .ZN(n4550) );
  AOI21_X1 U5067 ( .B1(n3445), .B2(n4572), .A(n4550), .ZN(n5034) );
  NAND2_X1 U5068 ( .A1(n5032), .A2(n5034), .ZN(n4552) );
  NAND2_X1 U5069 ( .A1(n4551), .A2(n6762), .ZN(n5033) );
  NAND2_X1 U5070 ( .A1(n4552), .A2(n5033), .ZN(n5379) );
  NAND2_X1 U5071 ( .A1(n4553), .A2(n4572), .ZN(n4558) );
  NAND2_X1 U5072 ( .A1(n4555), .A2(n4554), .ZN(n4563) );
  XNOR2_X1 U5073 ( .A(n4563), .B(n4561), .ZN(n4556) );
  NAND2_X1 U5074 ( .A1(n4556), .A2(n4407), .ZN(n4557) );
  NAND2_X1 U5075 ( .A1(n4558), .A2(n4557), .ZN(n4559) );
  XNOR2_X1 U5076 ( .A(n4559), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n5380)
         );
  NAND2_X1 U5077 ( .A1(n4559), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4560)
         );
  INV_X1 U5078 ( .A(n4561), .ZN(n4562) );
  NOR2_X1 U5079 ( .A1(n4563), .A2(n4562), .ZN(n4565) );
  NAND2_X1 U5080 ( .A1(n4565), .A2(n4564), .ZN(n4584) );
  OAI211_X1 U5081 ( .C1(n4565), .C2(n4564), .A(n4584), .B(n4407), .ZN(n4566)
         );
  INV_X1 U5082 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4568) );
  XNOR2_X1 U5083 ( .A(n4569), .B(n4568), .ZN(n4903) );
  NAND2_X1 U5084 ( .A1(n4902), .A2(n4903), .ZN(n4571) );
  NAND2_X1 U5085 ( .A1(n4569), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4570)
         );
  NAND2_X1 U5086 ( .A1(n4571), .A2(n4570), .ZN(n6692) );
  INV_X1 U5087 ( .A(n4574), .ZN(n4575) );
  OR2_X1 U5088 ( .A1(n4593), .A2(n4575), .ZN(n4578) );
  XNOR2_X1 U5089 ( .A(n4584), .B(n4585), .ZN(n4576) );
  NAND2_X1 U5090 ( .A1(n4576), .A2(n4407), .ZN(n4577) );
  NAND2_X1 U5091 ( .A1(n4578), .A2(n4577), .ZN(n4579) );
  NAND2_X1 U5092 ( .A1(n6692), .A2(n6694), .ZN(n4580) );
  NAND2_X1 U5093 ( .A1(n4579), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6693)
         );
  NAND2_X1 U5094 ( .A1(n4580), .A2(n6693), .ZN(n6699) );
  INV_X1 U5095 ( .A(n4581), .ZN(n4583) );
  INV_X1 U5096 ( .A(n4584), .ZN(n4586) );
  NAND2_X1 U5097 ( .A1(n4586), .A2(n4585), .ZN(n4594) );
  XNOR2_X1 U5098 ( .A(n4594), .B(n4595), .ZN(n4587) );
  NAND2_X1 U5099 ( .A1(n4587), .A2(n4407), .ZN(n4588) );
  INV_X1 U5100 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6793) );
  XNOR2_X1 U5101 ( .A(n4590), .B(n6793), .ZN(n6702) );
  NAND2_X1 U5102 ( .A1(n6699), .A2(n6702), .ZN(n6700) );
  NAND2_X1 U5103 ( .A1(n4590), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4591)
         );
  INV_X1 U5104 ( .A(n4594), .ZN(n4596) );
  NAND3_X1 U5105 ( .A1(n4596), .A2(n4407), .A3(n4595), .ZN(n4597) );
  NAND2_X1 U5106 ( .A1(n4614), .A2(n4597), .ZN(n4599) );
  XNOR2_X1 U5107 ( .A(n4599), .B(n4598), .ZN(n5478) );
  NAND2_X1 U5108 ( .A1(n4599), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4600)
         );
  INV_X2 U5109 ( .A(n6089), .ZN(n6137) );
  INV_X1 U5110 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4601) );
  OR2_X1 U5111 ( .A1(n6187), .A2(n4601), .ZN(n4602) );
  NAND2_X1 U5112 ( .A1(n6171), .A2(n6807), .ZN(n5678) );
  NAND2_X1 U5113 ( .A1(n5677), .A2(n5678), .ZN(n4604) );
  OR2_X1 U5114 ( .A1(n6171), .A2(n6807), .ZN(n5679) );
  INV_X1 U5115 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U5116 ( .A1(n6171), .A2(n5701), .ZN(n5689) );
  NAND2_X1 U5117 ( .A1(n5691), .A2(n5689), .ZN(n4605) );
  NAND2_X1 U5118 ( .A1(n4605), .A2(n5690), .ZN(n5720) );
  INV_X1 U5119 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4606) );
  NOR2_X1 U5120 ( .A1(n6187), .A2(n4606), .ZN(n5721) );
  OR2_X2 U5121 ( .A1(n5720), .A2(n5721), .ZN(n4607) );
  NAND2_X1 U5122 ( .A1(n6171), .A2(n4606), .ZN(n5722) );
  XNOR2_X1 U5123 ( .A(n6187), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5748)
         );
  INV_X1 U5124 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U5125 ( .A1(n6171), .A2(n5750), .ZN(n4608) );
  NAND2_X1 U5126 ( .A1(n6171), .A2(n5769), .ZN(n4609) );
  NAND2_X1 U5127 ( .A1(n4610), .A2(n4609), .ZN(n6196) );
  INV_X1 U5128 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U5129 ( .A1(n6196), .A2(n6195), .ZN(n4611) );
  NAND2_X1 U5130 ( .A1(n6171), .A2(n6832), .ZN(n6194) );
  NAND2_X1 U5131 ( .A1(n4611), .A2(n6194), .ZN(n6186) );
  INV_X1 U5132 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U5133 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5791) );
  INV_X1 U5134 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6532) );
  AND3_X1 U5135 ( .A1(n6532), .A2(n6841), .A3(n6537), .ZN(n4612) );
  NOR2_X1 U5136 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6307) );
  NOR2_X1 U5137 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6116) );
  INV_X1 U5138 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6275) );
  NAND4_X1 U5139 ( .A1(n6307), .A2(n6116), .A3(n6275), .A4(n6269), .ZN(n4615)
         );
  AND2_X1 U5140 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6308) );
  AND2_X1 U5141 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U5142 ( .A1(n6308), .A2(n5797), .ZN(n6127) );
  NAND2_X1 U5143 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5800) );
  NOR2_X1 U5144 ( .A1(n6127), .A2(n5800), .ZN(n5809) );
  INV_X1 U5145 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6251) );
  XNOR2_X1 U5146 ( .A(n6187), .B(n6251), .ZN(n6105) );
  NAND2_X1 U5147 ( .A1(n6171), .A2(n6251), .ZN(n4616) );
  INV_X1 U5148 ( .A(n6097), .ZN(n4617) );
  INV_X1 U5149 ( .A(n6087), .ZN(n4618) );
  INV_X1 U5150 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U5151 ( .A1(n4618), .A2(n3535), .ZN(n6078) );
  NOR2_X1 U5152 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4619) );
  OR2_X1 U5153 ( .A1(n6171), .A2(n4619), .ZN(n6077) );
  OR2_X1 U5154 ( .A1(n6171), .A2(n4621), .ZN(n4620) );
  INV_X1 U5155 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4622) );
  XNOR2_X1 U5156 ( .A(n6187), .B(n4622), .ZN(n4688) );
  OAI21_X1 U5157 ( .B1(n3815), .B2(n3750), .A(n4855), .ZN(n4625) );
  NAND3_X1 U5158 ( .A1(n3809), .A2(n4626), .A3(n4625), .ZN(n4725) );
  NOR2_X1 U5159 ( .A1(n4725), .A2(n4627), .ZN(n7021) );
  INV_X1 U5160 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n4629) );
  NAND2_X1 U5161 ( .A1(n7046), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5113) );
  INV_X1 U5162 ( .A(n5113), .ZN(n5157) );
  NAND2_X1 U5163 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n5157), .ZN(n6733) );
  NAND2_X1 U5164 ( .A1(n4630), .A2(n7139), .ZN(n6740) );
  NAND2_X1 U5165 ( .A1(n6740), .A2(n7046), .ZN(n4631) );
  AND2_X2 U5166 ( .A1(n6993), .A2(n4631), .ZN(n6691) );
  NAND2_X1 U5167 ( .A1(n7046), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4633) );
  NAND2_X1 U5168 ( .A1(n7126), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4632) );
  AND2_X1 U5169 ( .A1(n4633), .A2(n4632), .ZN(n4760) );
  INV_X2 U5170 ( .A(n6801), .ZN(n6843) );
  NAND2_X1 U5171 ( .A1(n6843), .A2(REIP_REG_29__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U5172 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4634)
         );
  OAI211_X1 U5173 ( .C1(n5863), .C2(n6707), .A(n6222), .B(n4634), .ZN(n4635)
         );
  AOI21_X1 U5174 ( .B1(n4636), .B2(n6710), .A(n4635), .ZN(n4637) );
  INV_X1 U5175 ( .A(n4638), .ZN(n4639) );
  NAND2_X1 U5176 ( .A1(n4639), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4696)
         );
  XNOR2_X1 U5177 ( .A(n4696), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5829)
         );
  NOR2_X1 U5178 ( .A1(n4641), .A2(n4640), .ZN(n4659) );
  AOI22_X1 U5179 ( .A1(n3832), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4642), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4647) );
  AOI22_X1 U5180 ( .A1(n3903), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4646) );
  AOI22_X1 U5181 ( .A1(n3734), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3835), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4645) );
  AOI22_X1 U5182 ( .A1(n4643), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3827), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4644) );
  NAND4_X1 U5183 ( .A1(n4647), .A2(n4646), .A3(n4645), .A4(n4644), .ZN(n4657)
         );
  AOI22_X1 U5184 ( .A1(n4648), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5185 ( .A1(n3833), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4649), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4654) );
  AOI22_X1 U5186 ( .A1(n4650), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4653) );
  AOI22_X1 U5187 ( .A1(n3557), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4651), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4652) );
  NAND4_X1 U5188 ( .A1(n4655), .A2(n4654), .A3(n4653), .A4(n4652), .ZN(n4656)
         );
  NOR2_X1 U5189 ( .A1(n4657), .A2(n4656), .ZN(n4658) );
  XNOR2_X1 U5190 ( .A(n4659), .B(n4658), .ZN(n4665) );
  INV_X1 U5191 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4661) );
  NAND2_X1 U5192 ( .A1(n7128), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4660)
         );
  OAI211_X1 U5193 ( .C1(n4662), .C2(n4661), .A(n4660), .B(n3690), .ZN(n4663)
         );
  AOI21_X1 U5194 ( .B1(n4665), .B2(n4664), .A(n4663), .ZN(n4666) );
  AOI21_X1 U5195 ( .B1(n5829), .B2(n3544), .A(n4666), .ZN(n4701) );
  AOI22_X1 U5196 ( .A1(n4668), .A2(EAX_REG_31__SCAN_IN), .B1(n4667), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4669) );
  INV_X1 U5197 ( .A(n4669), .ZN(n4670) );
  INV_X1 U5198 ( .A(READY_N), .ZN(n7028) );
  OR2_X1 U5199 ( .A1(n4725), .A2(n6714), .ZN(n4735) );
  NOR3_X1 U5200 ( .A1(n4675), .A2(n4674), .A3(n4673), .ZN(n4676) );
  OR2_X1 U5201 ( .A1(n4677), .A2(n4676), .ZN(n4679) );
  NAND2_X1 U5202 ( .A1(n4679), .A2(n4678), .ZN(n6715) );
  NAND2_X1 U5203 ( .A1(n7028), .A2(n6715), .ZN(n4720) );
  OAI22_X1 U5204 ( .A1(n6988), .A2(n4735), .B1(n4720), .B2(n4923), .ZN(n4780)
         );
  NOR2_X1 U5205 ( .A1(n4746), .A2(n4681), .ZN(n4682) );
  AOI21_X1 U5206 ( .B1(n4780), .B2(n6992), .A(n4682), .ZN(n4683) );
  AND2_X1 U5207 ( .A1(n5839), .A2(n5028), .ZN(n4684) );
  NAND2_X1 U5208 ( .A1(n7096), .A2(EAX_REG_31__SCAN_IN), .ZN(n4685) );
  NAND2_X1 U5209 ( .A1(n5839), .A2(n3854), .ZN(n5836) );
  INV_X1 U5210 ( .A(DATAI_31_), .ZN(n6424) );
  AND2_X1 U5211 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U5212 ( .A1(n6223), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5810) );
  AND2_X1 U5213 ( .A1(n6171), .A2(n5810), .ZN(n4690) );
  NAND2_X1 U5214 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4691) );
  NAND2_X1 U5215 ( .A1(n4691), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4692) );
  NAND3_X1 U5216 ( .A1(n4694), .A2(n4693), .A3(n4692), .ZN(n4695) );
  INV_X1 U5217 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6216) );
  XNOR2_X1 U5218 ( .A(n4695), .B(n6216), .ZN(n6221) );
  INV_X1 U5219 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5817) );
  INV_X1 U5220 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U5221 ( .A1(n6843), .A2(REIP_REG_31__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U5222 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4698)
         );
  OAI211_X1 U5223 ( .C1(n5179), .C2(n6707), .A(n6215), .B(n4698), .ZN(n4699)
         );
  OAI21_X1 U5224 ( .B1(n6221), .B2(n6993), .A(n4700), .ZN(U2955) );
  OAI22_X1 U5225 ( .A1(n5844), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n5843), .ZN(n5846) );
  INV_X1 U5226 ( .A(n5870), .ZN(n4707) );
  NAND2_X1 U5227 ( .A1(n5847), .A2(n4705), .ZN(n5845) );
  INV_X1 U5228 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4709) );
  OAI22_X1 U5229 ( .A1(n5834), .A2(n6045), .B1(n4709), .B2(n6047), .ZN(n4710)
         );
  INV_X1 U5230 ( .A(n4710), .ZN(n4711) );
  AND3_X1 U5231 ( .A1(n3438), .A2(n6992), .A3(n6715), .ZN(n5155) );
  INV_X1 U5232 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6476) );
  INV_X1 U5233 ( .A(n5156), .ZN(n4714) );
  OAI211_X1 U5234 ( .C1(n5155), .C2(n6476), .A(n4714), .B(n6726), .ZN(U2788)
         );
  OR2_X1 U5235 ( .A1(n5844), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4716)
         );
  AND2_X1 U5236 ( .A1(n4716), .A2(n4715), .ZN(n5469) );
  INV_X1 U5237 ( .A(n5469), .ZN(n4719) );
  XNOR2_X1 U5238 ( .A(n4718), .B(n4717), .ZN(n5476) );
  OAI222_X1 U5239 ( .A1(n4719), .A2(n6045), .B1(n6039), .B2(n5476), .C1(n4426), 
        .C2(n6047), .ZN(U2859) );
  NAND2_X1 U5240 ( .A1(n7067), .A2(n7075), .ZN(n6730) );
  AOI21_X1 U5241 ( .B1(n4418), .B2(n6730), .A(n4720), .ZN(n4723) );
  NOR2_X1 U5242 ( .A1(n3854), .A2(n4855), .ZN(n4721) );
  NOR2_X1 U5243 ( .A1(n6988), .A2(n4721), .ZN(n4722) );
  MUX2_X1 U5244 ( .A(n4723), .B(n4722), .S(n4867), .Z(n4731) );
  NAND2_X1 U5245 ( .A1(n5184), .A2(n6730), .ZN(n5165) );
  NAND2_X1 U5246 ( .A1(n5165), .A2(n7028), .ZN(n4724) );
  OR2_X1 U5247 ( .A1(n6988), .A2(n4724), .ZN(n4775) );
  INV_X1 U5248 ( .A(n3438), .ZN(n6716) );
  INV_X1 U5249 ( .A(n4725), .ZN(n4727) );
  NAND2_X1 U5250 ( .A1(n4727), .A2(n4726), .ZN(n4728) );
  NAND2_X1 U5251 ( .A1(n6716), .A2(n4728), .ZN(n4778) );
  OAI211_X1 U5252 ( .C1(n4775), .C2(n4786), .A(n4729), .B(n4778), .ZN(n4730)
         );
  OAI22_X1 U5253 ( .A1(n4672), .A2(n5184), .B1(n4871), .B2(n4733), .ZN(n4734)
         );
  INV_X1 U5254 ( .A(n4734), .ZN(n4736) );
  INV_X1 U5255 ( .A(n4735), .ZN(n4789) );
  NOR2_X1 U5256 ( .A1(n7021), .A2(n4789), .ZN(n6983) );
  NAND3_X1 U5257 ( .A1(n4736), .A2(n6983), .A3(n4923), .ZN(n4737) );
  NOR2_X1 U5258 ( .A1(n4738), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4739)
         );
  OR2_X1 U5259 ( .A1(n5053), .A2(n4739), .ZN(n4766) );
  AND2_X1 U5260 ( .A1(n3438), .A2(n4418), .ZN(n7000) );
  NAND2_X1 U5261 ( .A1(n4751), .A2(n7000), .ZN(n5753) );
  NAND2_X1 U5262 ( .A1(n4756), .A2(n6801), .ZN(n6542) );
  NAND2_X1 U5263 ( .A1(n5753), .A2(n6542), .ZN(n4752) );
  INV_X1 U5264 ( .A(n4740), .ZN(n4741) );
  NOR2_X1 U5265 ( .A1(n4784), .A2(n4741), .ZN(n6982) );
  INV_X1 U5266 ( .A(n4742), .ZN(n4743) );
  NAND2_X1 U5267 ( .A1(n4743), .A2(n4354), .ZN(n4938) );
  INV_X1 U5268 ( .A(n4785), .ZN(n4744) );
  NAND2_X1 U5269 ( .A1(n4744), .A2(n4855), .ZN(n4745) );
  OAI211_X1 U5270 ( .C1(n4746), .C2(n3428), .A(n4938), .B(n4745), .ZN(n4747)
         );
  NOR2_X1 U5271 ( .A1(n4748), .A2(n4747), .ZN(n4749) );
  NAND2_X1 U5272 ( .A1(n3431), .A2(n4749), .ZN(n4750) );
  NAND2_X1 U5273 ( .A1(n4751), .A2(n4750), .ZN(n5697) );
  NAND2_X1 U5274 ( .A1(n6744), .A2(n5697), .ZN(n5751) );
  INV_X1 U5275 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5696) );
  AND2_X1 U5276 ( .A1(n5751), .A2(n5696), .ZN(n6544) );
  AOI21_X1 U5277 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n4752), .A(n6544), 
        .ZN(n4758) );
  NAND2_X1 U5278 ( .A1(n3435), .A2(n4871), .ZN(n4754) );
  AND2_X1 U5279 ( .A1(n7030), .A2(n4754), .ZN(n4755) );
  AND2_X1 U5280 ( .A1(n6843), .A2(REIP_REG_0__SCAN_IN), .ZN(n4762) );
  AOI21_X1 U5281 ( .B1(n6846), .B2(n5469), .A(n4762), .ZN(n4757) );
  OAI211_X1 U5282 ( .C1(n6756), .C2(n4766), .A(n4758), .B(n4757), .ZN(U3018)
         );
  INV_X1 U5283 ( .A(n6691), .ZN(n6205) );
  INV_X1 U5284 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4759) );
  AOI21_X1 U5285 ( .B1(n6205), .B2(n4760), .A(n4759), .ZN(n4761) );
  INV_X1 U5286 ( .A(n4761), .ZN(n4765) );
  INV_X1 U5287 ( .A(n5476), .ZN(n4763) );
  AOI21_X1 U5288 ( .B1(n4763), .B2(n6710), .A(n4762), .ZN(n4764) );
  OAI211_X1 U5289 ( .C1(n4766), .C2(n6993), .A(n4765), .B(n4764), .ZN(U2986)
         );
  OAI21_X1 U5290 ( .B1(n4767), .B2(n4769), .A(n4768), .ZN(n5466) );
  AND2_X1 U5291 ( .A1(n4838), .A2(n4770), .ZN(n4771) );
  NOR2_X1 U5292 ( .A1(n5024), .A2(n4771), .ZN(n6867) );
  AOI22_X1 U5293 ( .A1(n6037), .A2(n6867), .B1(EBX_REG_5__SCAN_IN), .B2(n6012), 
        .ZN(n4772) );
  OAI21_X1 U5294 ( .B1(n5466), .B2(n6039), .A(n4772), .ZN(U2854) );
  NOR2_X1 U5295 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4629), .ZN(n4854) );
  INV_X1 U5296 ( .A(n6730), .ZN(n6736) );
  NAND2_X1 U5297 ( .A1(n7000), .A2(n6736), .ZN(n4773) );
  AND2_X1 U5298 ( .A1(n4773), .A2(n4672), .ZN(n4776) );
  OAI21_X1 U5299 ( .B1(n4776), .B2(n4775), .A(n4774), .ZN(n4782) );
  NAND2_X1 U5300 ( .A1(n4778), .A2(n4777), .ZN(n4779) );
  OR2_X1 U5301 ( .A1(n4780), .A2(n4779), .ZN(n4781) );
  INV_X1 U5302 ( .A(n4944), .ZN(n7003) );
  NAND2_X1 U5303 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n7040) );
  NOR2_X1 U5304 ( .A1(n7046), .A2(n7040), .ZN(n6735) );
  INV_X1 U5305 ( .A(n6735), .ZN(n7038) );
  INV_X1 U5306 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7024) );
  OAI22_X1 U5307 ( .A1(n7003), .A2(n7051), .B1(n7038), .B2(n7024), .ZN(n6997)
         );
  NOR2_X1 U5308 ( .A1(n4854), .A2(n6997), .ZN(n6995) );
  INV_X1 U5309 ( .A(n4784), .ZN(n4788) );
  AND3_X1 U5310 ( .A1(n4923), .A2(n4786), .A3(n4785), .ZN(n4787) );
  NAND2_X1 U5311 ( .A1(n4788), .A2(n4787), .ZN(n6559) );
  OR2_X1 U5312 ( .A1(n6982), .A2(n4789), .ZN(n4930) );
  XNOR2_X1 U5313 ( .A(n4790), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4791)
         );
  NAND2_X1 U5314 ( .A1(n4930), .A2(n4791), .ZN(n4795) );
  XNOR2_X1 U5315 ( .A(n6552), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4793)
         );
  NOR2_X1 U5316 ( .A1(n4938), .A2(n4791), .ZN(n4792) );
  AOI21_X1 U5317 ( .B1(n7000), .B2(n4793), .A(n4792), .ZN(n4794) );
  NAND2_X1 U5318 ( .A1(n4795), .A2(n4794), .ZN(n4796) );
  AOI21_X1 U5319 ( .B1(n3447), .B2(n6559), .A(n4796), .ZN(n4942) );
  INV_X1 U5320 ( .A(n4942), .ZN(n4799) );
  NOR2_X1 U5321 ( .A1(n6732), .A2(n5696), .ZN(n6562) );
  INV_X1 U5322 ( .A(n6562), .ZN(n4803) );
  AOI22_X1 U5323 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6216), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5052), .ZN(n6561) );
  NAND3_X1 U5324 ( .A1(n4790), .A2(n4847), .A3(n4927), .ZN(n4797) );
  OAI21_X1 U5325 ( .B1(n4803), .B2(n6561), .A(n4797), .ZN(n4798) );
  AOI21_X1 U5326 ( .B1(n4799), .B2(n6560), .A(n4798), .ZN(n4801) );
  INV_X1 U5327 ( .A(n4847), .ZN(n7047) );
  NOR2_X1 U5328 ( .A1(n4790), .A2(n7047), .ZN(n6564) );
  OAI21_X1 U5329 ( .B1(n6995), .B2(n6564), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4800) );
  OAI21_X1 U5330 ( .B1(n6995), .B2(n4801), .A(n4800), .ZN(U3459) );
  AOI21_X1 U5331 ( .B1(n7000), .B2(n6560), .A(n6995), .ZN(n4806) );
  NOR2_X1 U5332 ( .A1(n3784), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4802)
         );
  AOI21_X1 U5333 ( .B1(n3443), .B2(n6559), .A(n4802), .ZN(n7002) );
  OAI21_X1 U5334 ( .B1(n7002), .B2(STATE2_REG_3__SCAN_IN), .A(n6732), .ZN(
        n4804) );
  AOI22_X1 U5335 ( .A1(n4804), .A2(n4803), .B1(n4847), .B2(n3468), .ZN(n4805)
         );
  OAI22_X1 U5336 ( .A1(n4806), .A2(n3468), .B1(n6995), .B2(n4805), .ZN(U3461)
         );
  NAND2_X1 U5337 ( .A1(n5753), .A2(n5697), .ZN(n6525) );
  NAND2_X1 U5338 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6745) );
  OAI21_X1 U5339 ( .B1(n5697), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6542), 
        .ZN(n5788) );
  AOI21_X1 U5340 ( .B1(n6525), .B2(n6745), .A(n5788), .ZN(n6778) );
  NAND2_X1 U5341 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4807) );
  OAI21_X1 U5342 ( .B1(n5052), .B2(n5696), .A(n4542), .ZN(n6764) );
  OAI21_X1 U5343 ( .B1(n4542), .B2(n4807), .A(n6764), .ZN(n4818) );
  NAND2_X1 U5344 ( .A1(n4809), .A2(n4808), .ZN(n4810) );
  XNOR2_X1 U5345 ( .A(n4811), .B(n4810), .ZN(n6686) );
  NOR2_X1 U5346 ( .A1(n6756), .A2(n6686), .ZN(n4817) );
  NOR2_X1 U5347 ( .A1(n4813), .A2(n4812), .ZN(n4814) );
  OR2_X1 U5348 ( .A1(n4913), .A2(n4814), .ZN(n5521) );
  INV_X1 U5349 ( .A(REIP_REG_2__SCAN_IN), .ZN(n4815) );
  OAI22_X1 U5350 ( .A1(n6836), .A2(n5521), .B1(n6801), .B2(n4815), .ZN(n4816)
         );
  AOI211_X1 U5351 ( .C1(n6768), .C2(n4818), .A(n4817), .B(n4816), .ZN(n4820)
         );
  NAND2_X1 U5352 ( .A1(n5753), .A2(n5696), .ZN(n6548) );
  NAND2_X1 U5353 ( .A1(n6525), .A2(n6548), .ZN(n6746) );
  INV_X1 U5354 ( .A(n6746), .ZN(n6531) );
  NAND3_X1 U5355 ( .A1(n6531), .A2(n4542), .A3(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4819) );
  OAI211_X1 U5356 ( .C1(n6778), .C2(n4542), .A(n4820), .B(n4819), .ZN(U3016)
         );
  INV_X1 U5357 ( .A(n4822), .ZN(n4825) );
  INV_X1 U5358 ( .A(n4823), .ZN(n4824) );
  OR3_X1 U5359 ( .A1(n4826), .A2(n4825), .A3(n4824), .ZN(n4827) );
  NAND2_X1 U5360 ( .A1(n4821), .A2(n4827), .ZN(n6684) );
  INV_X1 U5361 ( .A(n5521), .ZN(n4828) );
  AOI22_X1 U5362 ( .A1(n6037), .A2(n4828), .B1(n6012), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4829) );
  OAI21_X1 U5363 ( .B1(n6039), .B2(n6684), .A(n4829), .ZN(U2857) );
  OR2_X1 U5364 ( .A1(n4831), .A2(n4830), .ZN(n4832) );
  AND2_X1 U5365 ( .A1(n4822), .A2(n4832), .ZN(n5181) );
  INV_X1 U5366 ( .A(n5181), .ZN(n5467) );
  XNOR2_X1 U5367 ( .A(n5177), .B(n4833), .ZN(n6547) );
  AOI22_X1 U5368 ( .A1(n6037), .A2(n6547), .B1(n6012), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4834) );
  OAI21_X1 U5369 ( .B1(n6039), .B2(n5467), .A(n4834), .ZN(U2858) );
  NOR2_X1 U5370 ( .A1(n4835), .A2(n4836), .ZN(n4837) );
  OR2_X1 U5371 ( .A1(n4767), .A2(n4837), .ZN(n6858) );
  INV_X1 U5372 ( .A(n4838), .ZN(n4839) );
  AOI21_X1 U5373 ( .B1(n4840), .B2(n4915), .A(n4839), .ZN(n6852) );
  AOI22_X1 U5374 ( .A1(n6037), .A2(n6852), .B1(n6012), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4841) );
  OAI21_X1 U5375 ( .B1(n6039), .B2(n6858), .A(n4841), .ZN(U2855) );
  AND2_X1 U5376 ( .A1(n3444), .A2(n3443), .ZN(n7124) );
  AND2_X1 U5377 ( .A1(n4843), .A2(n3447), .ZN(n7142) );
  NOR2_X1 U5378 ( .A1(n4844), .A2(n5128), .ZN(n5369) );
  AOI21_X1 U5379 ( .B1(n7124), .B2(n7142), .A(n5369), .ZN(n4851) );
  INV_X1 U5380 ( .A(n4851), .ZN(n4846) );
  INV_X1 U5381 ( .A(n7139), .ZN(n7152) );
  NAND3_X1 U5382 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5131) );
  INV_X1 U5383 ( .A(n5131), .ZN(n4845) );
  AOI22_X1 U5384 ( .A1(n4846), .A2(n7152), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4845), .ZN(n5372) );
  NAND2_X1 U5385 ( .A1(n7128), .A2(n6732), .ZN(n7048) );
  AOI21_X1 U5386 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7123), .A(n4953), .ZN(
        n7149) );
  OR2_X1 U5387 ( .A1(n5208), .A2(n5207), .ZN(n5089) );
  INV_X1 U5388 ( .A(n4849), .ZN(n4880) );
  NOR2_X1 U5389 ( .A1(n7139), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5280) );
  INV_X1 U5390 ( .A(n5280), .ZN(n5632) );
  OAI21_X1 U5391 ( .B1(n4856), .B2(n6685), .A(n5632), .ZN(n4850) );
  AOI22_X1 U5392 ( .A1(n4851), .A2(n4850), .B1(n7139), .B2(n5131), .ZN(n4852)
         );
  NAND2_X1 U5393 ( .A1(n7149), .A2(n4852), .ZN(n5367) );
  NAND2_X1 U5394 ( .A1(n5367), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4859)
         );
  NOR2_X2 U5395 ( .A1(n5193), .A2(n4855), .ZN(n7146) );
  NAND2_X1 U5396 ( .A1(n6710), .A2(DATAI_16_), .ZN(n7130) );
  NAND2_X1 U5397 ( .A1(n6710), .A2(DATAI_24_), .ZN(n5643) );
  OAI22_X1 U5398 ( .A1(n5603), .A2(n7130), .B1(n5393), .B2(n5643), .ZN(n4857)
         );
  AOI21_X1 U5399 ( .B1(n7146), .B2(n5369), .A(n4857), .ZN(n4858) );
  OAI211_X1 U5400 ( .C1(n5372), .C2(n7156), .A(n4859), .B(n4858), .ZN(U3140)
         );
  NAND2_X1 U5401 ( .A1(n5367), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4862)
         );
  NOR2_X2 U5402 ( .A1(n5193), .A2(n5028), .ZN(n7269) );
  NAND2_X1 U5403 ( .A1(n6710), .A2(DATAI_23_), .ZN(n7250) );
  NAND2_X1 U5404 ( .A1(n6710), .A2(DATAI_31_), .ZN(n5659) );
  OAI22_X1 U5405 ( .A1(n5603), .A2(n7250), .B1(n5393), .B2(n5659), .ZN(n4860)
         );
  AOI21_X1 U5406 ( .B1(n7269), .B2(n5369), .A(n4860), .ZN(n4861) );
  OAI211_X1 U5407 ( .C1(n5372), .C2(n7275), .A(n4862), .B(n4861), .ZN(U3147)
         );
  NAND2_X1 U5408 ( .A1(n5367), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4866)
         );
  NOR2_X2 U5409 ( .A1(n5193), .A2(n4863), .ZN(n7195) );
  NAND2_X1 U5410 ( .A1(n6710), .A2(DATAI_19_), .ZN(n7190) );
  NAND2_X1 U5411 ( .A1(n6710), .A2(DATAI_27_), .ZN(n5655) );
  OAI22_X1 U5412 ( .A1(n5603), .A2(n7190), .B1(n5393), .B2(n5655), .ZN(n4864)
         );
  AOI21_X1 U5413 ( .B1(n7195), .B2(n5369), .A(n4864), .ZN(n4865) );
  OAI211_X1 U5414 ( .C1(n5372), .C2(n7199), .A(n4866), .B(n4865), .ZN(U3143)
         );
  NAND2_X1 U5415 ( .A1(n5367), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4870)
         );
  NOR2_X2 U5416 ( .A1(n5193), .A2(n4867), .ZN(n7181) );
  NAND2_X1 U5417 ( .A1(n6710), .A2(DATAI_18_), .ZN(n7176) );
  NAND2_X1 U5418 ( .A1(n6710), .A2(DATAI_26_), .ZN(n5651) );
  OAI22_X1 U5419 ( .A1(n5603), .A2(n7176), .B1(n5393), .B2(n5651), .ZN(n4868)
         );
  AOI21_X1 U5420 ( .B1(n7181), .B2(n5369), .A(n4868), .ZN(n4869) );
  OAI211_X1 U5421 ( .C1(n5372), .C2(n7185), .A(n4870), .B(n4869), .ZN(U3142)
         );
  NAND2_X1 U5422 ( .A1(n5367), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4874)
         );
  NOR2_X2 U5423 ( .A1(n5193), .A2(n4871), .ZN(n7210) );
  NAND2_X1 U5424 ( .A1(n6710), .A2(DATAI_20_), .ZN(n7205) );
  NAND2_X1 U5425 ( .A1(n6710), .A2(DATAI_28_), .ZN(n5647) );
  OAI22_X1 U5426 ( .A1(n5603), .A2(n7205), .B1(n5393), .B2(n5647), .ZN(n4872)
         );
  AOI21_X1 U5427 ( .B1(n7210), .B2(n5369), .A(n4872), .ZN(n4873) );
  OAI211_X1 U5428 ( .C1(n5372), .C2(n7214), .A(n4874), .B(n4873), .ZN(U3144)
         );
  INV_X1 U5429 ( .A(n4843), .ZN(n5174) );
  AND2_X1 U5430 ( .A1(n3447), .A2(n5174), .ZN(n7101) );
  INV_X1 U5431 ( .A(n5129), .ZN(n4875) );
  OR2_X1 U5432 ( .A1(n4998), .A2(n4875), .ZN(n4876) );
  INV_X1 U5433 ( .A(n4876), .ZN(n5568) );
  NAND2_X1 U5434 ( .A1(n4877), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5286) );
  INV_X1 U5435 ( .A(n5286), .ZN(n5130) );
  AOI22_X1 U5436 ( .A1(n5569), .A2(n7101), .B1(n5568), .B2(n5130), .ZN(n5366)
         );
  NAND3_X1 U5437 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n5128), .A3(n7008), .ZN(n4967) );
  NOR2_X1 U5438 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4967), .ZN(n5363)
         );
  INV_X1 U5439 ( .A(n5363), .ZN(n4879) );
  AND2_X1 U5440 ( .A1(n4876), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5577) );
  INV_X1 U5441 ( .A(n4877), .ZN(n4878) );
  NAND2_X1 U5442 ( .A1(n4878), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U5443 ( .A1(n5285), .A2(n5278), .ZN(n5140) );
  AOI211_X1 U5444 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4879), .A(n5577), .B(
        n5140), .ZN(n4886) );
  NOR2_X1 U5445 ( .A1(n7101), .A2(n7139), .ZN(n5000) );
  NAND2_X1 U5446 ( .A1(n4960), .A2(n4880), .ZN(n4955) );
  INV_X1 U5447 ( .A(n4881), .ZN(n4882) );
  NAND2_X1 U5448 ( .A1(n4882), .A2(n3446), .ZN(n5062) );
  NOR2_X1 U5449 ( .A1(n5062), .A2(n7057), .ZN(n4999) );
  OAI21_X1 U5450 ( .B1(n5197), .B2(n5319), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4884) );
  OAI21_X1 U5451 ( .B1(n5000), .B2(n5571), .A(n4884), .ZN(n4885) );
  NAND2_X1 U5452 ( .A1(n4886), .A2(n4885), .ZN(n5359) );
  NAND2_X1 U5453 ( .A1(n5359), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4889) );
  OAI22_X1 U5454 ( .A1(n5361), .A2(n7250), .B1(n5659), .B2(n5360), .ZN(n4887)
         );
  AOI21_X1 U5455 ( .B1(n7269), .B2(n5363), .A(n4887), .ZN(n4888) );
  OAI211_X1 U5456 ( .C1(n5366), .C2(n7275), .A(n4889), .B(n4888), .ZN(U3059)
         );
  NAND2_X1 U5457 ( .A1(n5359), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4892) );
  OAI22_X1 U5458 ( .A1(n5361), .A2(n7130), .B1(n5643), .B2(n5360), .ZN(n4890)
         );
  AOI21_X1 U5459 ( .B1(n7146), .B2(n5363), .A(n4890), .ZN(n4891) );
  OAI211_X1 U5460 ( .C1(n5366), .C2(n7156), .A(n4892), .B(n4891), .ZN(U3052)
         );
  NAND2_X1 U5461 ( .A1(n5359), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4895) );
  OAI22_X1 U5462 ( .A1(n5361), .A2(n7205), .B1(n5647), .B2(n5360), .ZN(n4893)
         );
  AOI21_X1 U5463 ( .B1(n7210), .B2(n5363), .A(n4893), .ZN(n4894) );
  OAI211_X1 U5464 ( .C1(n5366), .C2(n7214), .A(n4895), .B(n4894), .ZN(U3056)
         );
  NAND2_X1 U5465 ( .A1(n5359), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4898) );
  OAI22_X1 U5466 ( .A1(n5361), .A2(n7176), .B1(n5651), .B2(n5360), .ZN(n4896)
         );
  AOI21_X1 U5467 ( .B1(n7181), .B2(n5363), .A(n4896), .ZN(n4897) );
  OAI211_X1 U5468 ( .C1(n5366), .C2(n7185), .A(n4898), .B(n4897), .ZN(U3054)
         );
  NAND2_X1 U5469 ( .A1(n5359), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4901) );
  OAI22_X1 U5470 ( .A1(n5361), .A2(n7190), .B1(n5655), .B2(n5360), .ZN(n4899)
         );
  AOI21_X1 U5471 ( .B1(n7195), .B2(n5363), .A(n4899), .ZN(n4900) );
  OAI211_X1 U5472 ( .C1(n5366), .C2(n7199), .A(n4901), .B(n4900), .ZN(U3055)
         );
  XNOR2_X1 U5473 ( .A(n4902), .B(n4903), .ZN(n5044) );
  INV_X1 U5474 ( .A(n6825), .ZN(n6779) );
  INV_X1 U5475 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6762) );
  NOR2_X1 U5476 ( .A1(n4904), .A2(n6762), .ZN(n6765) );
  INV_X1 U5477 ( .A(n6764), .ZN(n5693) );
  NAND2_X1 U5478 ( .A1(n6768), .A2(n5693), .ZN(n4905) );
  OAI21_X1 U5479 ( .B1(n6779), .B2(n6765), .A(n6781), .ZN(n6766) );
  INV_X1 U5480 ( .A(n6765), .ZN(n6747) );
  NOR4_X1 U5481 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6746), .A3(n6745), 
        .A4(n6747), .ZN(n6767) );
  AOI21_X1 U5482 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n6766), .A(n6767), 
        .ZN(n4909) );
  INV_X1 U5483 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6617) );
  NOR2_X1 U5484 ( .A1(n6801), .A2(n6617), .ZN(n4907) );
  NOR4_X1 U5485 ( .A1(n6744), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6747), 
        .A4(n5693), .ZN(n4906) );
  AOI211_X1 U5486 ( .C1(n6846), .C2(n6867), .A(n4907), .B(n4906), .ZN(n4908)
         );
  OAI211_X1 U5487 ( .C1(n6756), .C2(n5044), .A(n4909), .B(n4908), .ZN(U3013)
         );
  AND2_X1 U5488 ( .A1(n4821), .A2(n4910), .ZN(n4911) );
  NOR2_X1 U5489 ( .A1(n4835), .A2(n4911), .ZN(n5515) );
  INV_X1 U5490 ( .A(n5515), .ZN(n5031) );
  INV_X1 U5491 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4916) );
  OR2_X1 U5492 ( .A1(n4913), .A2(n4912), .ZN(n4914) );
  AND2_X1 U5493 ( .A1(n4915), .A2(n4914), .ZN(n6755) );
  INV_X1 U5494 ( .A(n6755), .ZN(n5513) );
  OAI222_X1 U5495 ( .A1(n5031), .A2(n6039), .B1(n6047), .B2(n4916), .C1(n5513), 
        .C2(n6045), .ZN(U2856) );
  NAND2_X1 U5496 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n7024), .ZN(n4948) );
  INV_X1 U5497 ( .A(n4917), .ZN(n4947) );
  MUX2_X1 U5498 ( .A(n4944), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n4918) );
  INV_X1 U5499 ( .A(n4918), .ZN(n4925) );
  INV_X1 U5500 ( .A(n4919), .ZN(n4920) );
  NOR2_X1 U5501 ( .A1(n4921), .A2(n4920), .ZN(n4922) );
  XNOR2_X1 U5502 ( .A(n4922), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6866)
         );
  OR2_X1 U5503 ( .A1(n4923), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4924) );
  NOR2_X1 U5504 ( .A1(n6866), .A2(n4924), .ZN(n6996) );
  AOI21_X1 U5505 ( .B1(n4925), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n6996), 
        .ZN(n4950) );
  NAND2_X1 U5506 ( .A1(n3444), .A2(n6559), .ZN(n4941) );
  AOI21_X1 U5507 ( .B1(n4790), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3921), 
        .ZN(n4926) );
  NOR2_X1 U5508 ( .A1(n3557), .A2(n4926), .ZN(n6568) );
  INV_X1 U5509 ( .A(n4790), .ZN(n4935) );
  NAND2_X1 U5510 ( .A1(n4935), .A2(n4927), .ZN(n4929) );
  NAND2_X1 U5511 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4931) );
  INV_X1 U5512 ( .A(n4931), .ZN(n4928) );
  AOI22_X1 U5513 ( .A1(n4930), .A2(n4929), .B1(n7000), .B2(n4928), .ZN(n4933)
         );
  NAND2_X1 U5514 ( .A1(n7000), .A2(n4931), .ZN(n4932) );
  MUX2_X1 U5515 ( .A(n4933), .B(n4932), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4937) );
  NAND2_X1 U5516 ( .A1(n4935), .A2(n4934), .ZN(n4936) );
  OAI211_X1 U5517 ( .C1(n6568), .C2(n4938), .A(n4937), .B(n4936), .ZN(n4939)
         );
  INV_X1 U5518 ( .A(n4939), .ZN(n4940) );
  NAND2_X1 U5519 ( .A1(n4941), .A2(n4940), .ZN(n6567) );
  MUX2_X1 U5520 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6567), .S(n4944), 
        .Z(n7014) );
  NAND2_X1 U5521 ( .A1(n4944), .A2(n4942), .ZN(n4943) );
  OAI21_X1 U5522 ( .B1(n4944), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4943), 
        .ZN(n7010) );
  NOR2_X1 U5523 ( .A1(n7010), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4945) );
  NAND2_X1 U5524 ( .A1(n7014), .A2(n4945), .ZN(n4946) );
  OAI211_X1 U5525 ( .C1(n4948), .C2(n4947), .A(n4950), .B(n4946), .ZN(n7020)
         );
  NAND2_X1 U5526 ( .A1(n4950), .A2(n4949), .ZN(n4951) );
  NAND2_X1 U5527 ( .A1(n7020), .A2(n4951), .ZN(n7042) );
  NAND2_X1 U5528 ( .A1(n7042), .A2(n7024), .ZN(n4952) );
  NAND2_X1 U5529 ( .A1(n4952), .A2(n6735), .ZN(n4954) );
  NAND2_X1 U5530 ( .A1(n4954), .A2(n4953), .ZN(n7061) );
  OAI21_X1 U5531 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6732), .A(n7061), .ZN(
        n7053) );
  NAND2_X1 U5532 ( .A1(n7061), .A2(n7152), .ZN(n7058) );
  NAND2_X1 U5533 ( .A1(n4960), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4956) );
  NAND2_X1 U5534 ( .A1(n3446), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4959) );
  NOR2_X1 U5535 ( .A1(n4955), .A2(n4959), .ZN(n7140) );
  NAND3_X1 U5536 ( .A1(n4960), .A2(n4849), .A3(n5207), .ZN(n5132) );
  NOR2_X1 U5537 ( .A1(n5132), .A2(n7126), .ZN(n7100) );
  AOI211_X1 U5538 ( .C1(n3445), .C2(n4956), .A(n7140), .B(n7100), .ZN(n4957)
         );
  OAI222_X1 U5539 ( .A1(n7061), .A2(n5128), .B1(n5282), .B2(n7053), .C1(n7058), 
        .C2(n4957), .ZN(U3462) );
  XNOR2_X1 U5540 ( .A(n3446), .B(STATEBS16_REG_SCAN_IN), .ZN(n4958) );
  OAI222_X1 U5541 ( .A1(n4958), .A2(n7058), .B1(n5174), .B2(n7053), .C1(n7008), 
        .C2(n7061), .ZN(U3464) );
  INV_X1 U5542 ( .A(n3447), .ZN(n4963) );
  OR2_X1 U5543 ( .A1(n5062), .A2(n7126), .ZN(n7111) );
  NAND2_X1 U5544 ( .A1(n4960), .A2(n4959), .ZN(n4961) );
  AND2_X1 U5545 ( .A1(n7111), .A2(n4961), .ZN(n4962) );
  OAI222_X1 U5546 ( .A1(n7061), .A2(n7012), .B1(n4963), .B2(n7053), .C1(n7058), 
        .C2(n4962), .ZN(U3463) );
  INV_X1 U5547 ( .A(n7269), .ZN(n4974) );
  NOR2_X1 U5548 ( .A1(n7123), .A2(n4967), .ZN(n4964) );
  INV_X1 U5549 ( .A(n4964), .ZN(n5201) );
  INV_X1 U5550 ( .A(n3443), .ZN(n5472) );
  NOR2_X1 U5551 ( .A1(n3444), .A2(n5472), .ZN(n7143) );
  AOI21_X1 U5552 ( .B1(n7143), .B2(n7101), .A(n4964), .ZN(n4969) );
  INV_X1 U5553 ( .A(n4969), .ZN(n4966) );
  OAI21_X1 U5554 ( .B1(n4971), .B2(n7126), .A(n7152), .ZN(n4968) );
  NAND2_X1 U5555 ( .A1(n7139), .A2(n4967), .ZN(n4965) );
  OAI211_X1 U5556 ( .C1(n4966), .C2(n4968), .A(n7149), .B(n4965), .ZN(n5196)
         );
  INV_X1 U5557 ( .A(n7275), .ZN(n4970) );
  OAI22_X1 U5558 ( .A1(n4969), .A2(n4968), .B1(n7128), .B2(n4967), .ZN(n5194)
         );
  AOI22_X1 U5559 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5196), .B1(n4970), 
        .B2(n5194), .ZN(n4973) );
  INV_X1 U5560 ( .A(n7250), .ZN(n7271) );
  INV_X1 U5561 ( .A(n5659), .ZN(n7267) );
  AOI22_X1 U5562 ( .A1(n7271), .A2(n5198), .B1(n5197), .B2(n7267), .ZN(n4972)
         );
  OAI211_X1 U5563 ( .C1(n4974), .C2(n5201), .A(n4973), .B(n4972), .ZN(U3067)
         );
  INV_X1 U5564 ( .A(n7146), .ZN(n4978) );
  INV_X1 U5565 ( .A(n7156), .ZN(n4975) );
  AOI22_X1 U5566 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5196), .B1(n4975), 
        .B2(n5194), .ZN(n4977) );
  INV_X1 U5567 ( .A(n5643), .ZN(n7145) );
  INV_X1 U5568 ( .A(n7130), .ZN(n7153) );
  AOI22_X1 U5569 ( .A1(n7145), .A2(n5197), .B1(n5198), .B2(n7153), .ZN(n4976)
         );
  OAI211_X1 U5570 ( .C1(n4978), .C2(n5201), .A(n4977), .B(n4976), .ZN(U3060)
         );
  INV_X1 U5571 ( .A(n7181), .ZN(n4982) );
  INV_X1 U5572 ( .A(n7185), .ZN(n4979) );
  AOI22_X1 U5573 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5196), .B1(n4979), 
        .B2(n5194), .ZN(n4981) );
  INV_X1 U5574 ( .A(n7176), .ZN(n7180) );
  INV_X1 U5575 ( .A(n5651), .ZN(n7182) );
  AOI22_X1 U5576 ( .A1(n7180), .A2(n5198), .B1(n5197), .B2(n7182), .ZN(n4980)
         );
  OAI211_X1 U5577 ( .C1(n4982), .C2(n5201), .A(n4981), .B(n4980), .ZN(U3062)
         );
  INV_X1 U5578 ( .A(n7195), .ZN(n4986) );
  INV_X1 U5579 ( .A(n7199), .ZN(n4983) );
  AOI22_X1 U5580 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5196), .B1(n4983), 
        .B2(n5194), .ZN(n4985) );
  INV_X1 U5581 ( .A(n5655), .ZN(n7194) );
  INV_X1 U5582 ( .A(n7190), .ZN(n7196) );
  AOI22_X1 U5583 ( .A1(n7194), .A2(n5197), .B1(n5198), .B2(n7196), .ZN(n4984)
         );
  OAI211_X1 U5584 ( .C1(n4986), .C2(n5201), .A(n4985), .B(n4984), .ZN(U3063)
         );
  INV_X1 U5585 ( .A(n7210), .ZN(n4990) );
  INV_X1 U5586 ( .A(n7214), .ZN(n4987) );
  AOI22_X1 U5587 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5196), .B1(n4987), 
        .B2(n5194), .ZN(n4989) );
  INV_X1 U5588 ( .A(n5647), .ZN(n7211) );
  INV_X1 U5589 ( .A(n7205), .ZN(n7209) );
  AOI22_X1 U5590 ( .A1(n7211), .A2(n5197), .B1(n5198), .B2(n7209), .ZN(n4988)
         );
  OAI211_X1 U5591 ( .C1(n4990), .C2(n5201), .A(n4989), .B(n4988), .ZN(U3064)
         );
  NAND2_X1 U5592 ( .A1(n5255), .A2(DATAI_11_), .ZN(n5264) );
  AOI22_X1 U5593 ( .A1(n5275), .A2(EAX_REG_27__SCAN_IN), .B1(n5230), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U5594 ( .A1(n5264), .A2(n4992), .ZN(U2935) );
  NAND2_X1 U5595 ( .A1(n5255), .A2(DATAI_10_), .ZN(n5232) );
  AOI22_X1 U5596 ( .A1(n5275), .A2(EAX_REG_26__SCAN_IN), .B1(n5230), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U5597 ( .A1(n5232), .A2(n4993), .ZN(U2934) );
  NAND2_X1 U5598 ( .A1(n5255), .A2(DATAI_6_), .ZN(n5239) );
  AOI22_X1 U5599 ( .A1(n5275), .A2(EAX_REG_22__SCAN_IN), .B1(n5230), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n4994) );
  NAND2_X1 U5600 ( .A1(n5239), .A2(n4994), .ZN(U2930) );
  NAND2_X1 U5601 ( .A1(n5255), .A2(DATAI_9_), .ZN(n5244) );
  AOI22_X1 U5602 ( .A1(n5275), .A2(EAX_REG_25__SCAN_IN), .B1(n5230), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U5603 ( .A1(n5244), .A2(n4995), .ZN(U2933) );
  NAND2_X1 U5604 ( .A1(n5255), .A2(DATAI_8_), .ZN(n5260) );
  AOI22_X1 U5605 ( .A1(n5275), .A2(EAX_REG_24__SCAN_IN), .B1(n5230), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n4996) );
  NAND2_X1 U5606 ( .A1(n5260), .A2(n4996), .ZN(U2932) );
  NAND2_X1 U5607 ( .A1(n5255), .A2(DATAI_7_), .ZN(n5273) );
  AOI22_X1 U5608 ( .A1(n5275), .A2(EAX_REG_23__SCAN_IN), .B1(n5230), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U5609 ( .A1(n5273), .A2(n4997), .ZN(U2931) );
  NAND2_X1 U5610 ( .A1(n4998), .A2(n5129), .ZN(n5001) );
  INV_X1 U5611 ( .A(n5001), .ZN(n5412) );
  AOI22_X1 U5612 ( .A1(n5571), .A2(n7101), .B1(n5130), .B2(n5412), .ZN(n5378)
         );
  NAND2_X1 U5613 ( .A1(n4999), .A2(n3445), .ZN(n7251) );
  AOI21_X1 U5614 ( .B1(n7251), .B2(n7108), .A(n7126), .ZN(n5004) );
  NOR2_X1 U5615 ( .A1(n5000), .A2(n5569), .ZN(n5003) );
  NAND3_X1 U5616 ( .A1(n7008), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7104) );
  INV_X1 U5617 ( .A(n7104), .ZN(n7103) );
  NAND2_X1 U5618 ( .A1(n7123), .A2(n7103), .ZN(n5005) );
  AND2_X1 U5619 ( .A1(n5001), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5413) );
  AOI211_X1 U5620 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5005), .A(n5413), .B(
        n5140), .ZN(n5002) );
  NAND2_X1 U5621 ( .A1(n5373), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5008)
         );
  INV_X1 U5622 ( .A(n5005), .ZN(n5375) );
  OAI22_X1 U5623 ( .A1(n7251), .A2(n5659), .B1(n7108), .B2(n7250), .ZN(n5006)
         );
  AOI21_X1 U5624 ( .B1(n7269), .B2(n5375), .A(n5006), .ZN(n5007) );
  OAI211_X1 U5625 ( .C1(n5378), .C2(n7275), .A(n5008), .B(n5007), .ZN(U3123)
         );
  NAND2_X1 U5626 ( .A1(n5373), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5011)
         );
  OAI22_X1 U5627 ( .A1(n7251), .A2(n5647), .B1(n7108), .B2(n7205), .ZN(n5009)
         );
  AOI21_X1 U5628 ( .B1(n7210), .B2(n5375), .A(n5009), .ZN(n5010) );
  OAI211_X1 U5629 ( .C1(n5378), .C2(n7214), .A(n5011), .B(n5010), .ZN(U3120)
         );
  NAND2_X1 U5630 ( .A1(n5373), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5014)
         );
  OAI22_X1 U5631 ( .A1(n7251), .A2(n5651), .B1(n7108), .B2(n7176), .ZN(n5012)
         );
  AOI21_X1 U5632 ( .B1(n7181), .B2(n5375), .A(n5012), .ZN(n5013) );
  OAI211_X1 U5633 ( .C1(n5378), .C2(n7185), .A(n5014), .B(n5013), .ZN(U3118)
         );
  NAND2_X1 U5634 ( .A1(n5373), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5017)
         );
  OAI22_X1 U5635 ( .A1(n7251), .A2(n5655), .B1(n7108), .B2(n7190), .ZN(n5015)
         );
  AOI21_X1 U5636 ( .B1(n7195), .B2(n5375), .A(n5015), .ZN(n5016) );
  OAI211_X1 U5637 ( .C1(n5378), .C2(n7199), .A(n5017), .B(n5016), .ZN(U3119)
         );
  NAND2_X1 U5638 ( .A1(n5373), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5020)
         );
  OAI22_X1 U5639 ( .A1(n7251), .A2(n5643), .B1(n7108), .B2(n7130), .ZN(n5018)
         );
  AOI21_X1 U5640 ( .B1(n7146), .B2(n5375), .A(n5018), .ZN(n5019) );
  OAI211_X1 U5641 ( .C1(n5378), .C2(n7156), .A(n5020), .B(n5019), .ZN(U3116)
         );
  AOI21_X1 U5642 ( .B1(n5022), .B2(n4768), .A(n4034), .ZN(n6696) );
  INV_X1 U5643 ( .A(n6696), .ZN(n6886) );
  NOR2_X1 U5644 ( .A1(n5024), .A2(n5023), .ZN(n5025) );
  OR2_X1 U5645 ( .A1(n5049), .A2(n5025), .ZN(n6881) );
  INV_X1 U5646 ( .A(n6881), .ZN(n5026) );
  AOI22_X1 U5647 ( .A1(n6037), .A2(n5026), .B1(n6012), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n5027) );
  OAI21_X1 U5648 ( .B1(n6886), .B2(n6039), .A(n5027), .ZN(U2853) );
  OR2_X1 U5649 ( .A1(n4406), .A2(n5028), .ZN(n5029) );
  INV_X1 U5650 ( .A(n5029), .ZN(n5030) );
  INV_X1 U5651 ( .A(DATAI_0_), .ZN(n5240) );
  INV_X1 U5652 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6579) );
  OAI222_X1 U5653 ( .A1(n7086), .A2(n5476), .B1(n5745), .B2(n5240), .C1(n5839), 
        .C2(n6579), .ZN(U2891) );
  INV_X1 U5654 ( .A(DATAI_3_), .ZN(n6470) );
  INV_X1 U5655 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6585) );
  OAI222_X1 U5656 ( .A1(n5031), .A2(n7086), .B1(n5745), .B2(n6470), .C1(n5839), 
        .C2(n6585), .ZN(U2888) );
  INV_X1 U5657 ( .A(DATAI_2_), .ZN(n5233) );
  INV_X1 U5658 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6583) );
  OAI222_X1 U5659 ( .A1(n6684), .A2(n7086), .B1(n5745), .B2(n5233), .C1(n5839), 
        .C2(n6583), .ZN(U2889) );
  INV_X1 U5660 ( .A(DATAI_6_), .ZN(n6463) );
  OAI222_X1 U5661 ( .A1(n6886), .A2(n7086), .B1(n5745), .B2(n6463), .C1(n6592), 
        .C2(n5839), .ZN(U2885) );
  NAND2_X1 U5662 ( .A1(n5032), .A2(n5033), .ZN(n5036) );
  INV_X1 U5663 ( .A(n5034), .ZN(n5035) );
  XNOR2_X1 U5664 ( .A(n5036), .B(n5035), .ZN(n6757) );
  INV_X1 U5665 ( .A(n6757), .ZN(n5040) );
  AOI22_X1 U5666 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6843), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n5037) );
  OAI21_X1 U5667 ( .B1(n6707), .B2(n5518), .A(n5037), .ZN(n5038) );
  AOI21_X1 U5668 ( .B1(n6710), .B2(n5515), .A(n5038), .ZN(n5039) );
  OAI21_X1 U5669 ( .B1(n5040), .B2(n6993), .A(n5039), .ZN(U2983) );
  INV_X1 U5670 ( .A(n5466), .ZN(n6870) );
  AOI22_X1 U5671 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6843), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n5041) );
  OAI21_X1 U5672 ( .B1(n6707), .B2(n6868), .A(n5041), .ZN(n5042) );
  AOI21_X1 U5673 ( .B1(n6870), .B2(n6710), .A(n5042), .ZN(n5043) );
  OAI21_X1 U5674 ( .B1(n5044), .B2(n6993), .A(n5043), .ZN(U2981) );
  NAND2_X1 U5675 ( .A1(n5021), .A2(n5046), .ZN(n5047) );
  AND2_X1 U5676 ( .A1(n5045), .A2(n5047), .ZN(n6893) );
  INV_X1 U5677 ( .A(n6893), .ZN(n5468) );
  OAI21_X1 U5678 ( .B1(n5049), .B2(n5048), .A(n5125), .ZN(n5050) );
  INV_X1 U5679 ( .A(n5050), .ZN(n6890) );
  AOI22_X1 U5680 ( .A1(n6037), .A2(n6890), .B1(n6012), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5051) );
  OAI21_X1 U5681 ( .B1(n5468), .B2(n6039), .A(n5051), .ZN(U2852) );
  XNOR2_X1 U5682 ( .A(n5053), .B(n5052), .ZN(n5054) );
  XNOR2_X1 U5683 ( .A(n5055), .B(n5054), .ZN(n6545) );
  INV_X1 U5684 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5058) );
  AOI22_X1 U5685 ( .A1(n5181), .A2(n6710), .B1(n6843), .B2(REIP_REG_1__SCAN_IN), .ZN(n5056) );
  OAI21_X1 U5686 ( .B1(n6205), .B2(n5058), .A(n5056), .ZN(n5057) );
  AOI21_X1 U5687 ( .B1(n6709), .B2(n5058), .A(n5057), .ZN(n5059) );
  OAI21_X1 U5688 ( .B1(n6545), .B2(n6993), .A(n5059), .ZN(U2985) );
  OAI21_X1 U5689 ( .B1(n7111), .B2(n3445), .A(n7152), .ZN(n5064) );
  NAND2_X1 U5690 ( .A1(n5128), .A2(n7012), .ZN(n5203) );
  NOR2_X1 U5691 ( .A1(n5060), .A2(n5203), .ZN(n5324) );
  AOI21_X1 U5692 ( .B1(n7143), .B2(n3537), .A(n5324), .ZN(n5065) );
  INV_X1 U5693 ( .A(n5203), .ZN(n5570) );
  NAND2_X1 U5694 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5570), .ZN(n5284) );
  OAI22_X1 U5695 ( .A1(n5064), .A2(n5065), .B1(n5284), .B2(n7128), .ZN(n5061)
         );
  NOR2_X1 U5696 ( .A1(n5062), .A2(n5629), .ZN(n5630) );
  NAND2_X1 U5697 ( .A1(n5319), .A2(n7180), .ZN(n5069) );
  INV_X1 U5698 ( .A(n5064), .ZN(n5066) );
  AOI22_X1 U5699 ( .A1(n5066), .A2(n5065), .B1(n5284), .B2(n7139), .ZN(n5067)
         );
  NAND2_X1 U5700 ( .A1(n7149), .A2(n5067), .ZN(n5320) );
  NAND2_X1 U5701 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n5320), .ZN(n5068) );
  OAI211_X1 U5702 ( .C1(n5443), .C2(n5651), .A(n5069), .B(n5068), .ZN(n5070)
         );
  AOI21_X1 U5703 ( .B1(n7181), .B2(n5324), .A(n5070), .ZN(n5071) );
  OAI21_X1 U5704 ( .B1(n7185), .B2(n5326), .A(n5071), .ZN(U3046) );
  NAND2_X1 U5705 ( .A1(n5319), .A2(n7271), .ZN(n5073) );
  NAND2_X1 U5706 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n5320), .ZN(n5072) );
  OAI211_X1 U5707 ( .C1(n5443), .C2(n5659), .A(n5073), .B(n5072), .ZN(n5074)
         );
  AOI21_X1 U5708 ( .B1(n7269), .B2(n5324), .A(n5074), .ZN(n5075) );
  OAI21_X1 U5709 ( .B1(n7275), .B2(n5326), .A(n5075), .ZN(U3051) );
  NAND2_X1 U5710 ( .A1(n5319), .A2(n7209), .ZN(n5077) );
  NAND2_X1 U5711 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n5320), .ZN(n5076) );
  OAI211_X1 U5712 ( .C1(n5443), .C2(n5647), .A(n5077), .B(n5076), .ZN(n5078)
         );
  AOI21_X1 U5713 ( .B1(n7210), .B2(n5324), .A(n5078), .ZN(n5079) );
  OAI21_X1 U5714 ( .B1(n7214), .B2(n5326), .A(n5079), .ZN(U3048) );
  NAND2_X1 U5715 ( .A1(n5319), .A2(n7196), .ZN(n5081) );
  NAND2_X1 U5716 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n5320), .ZN(n5080) );
  OAI211_X1 U5717 ( .C1(n5443), .C2(n5655), .A(n5081), .B(n5080), .ZN(n5082)
         );
  AOI21_X1 U5718 ( .B1(n7195), .B2(n5324), .A(n5082), .ZN(n5083) );
  OAI21_X1 U5719 ( .B1(n7199), .B2(n5326), .A(n5083), .ZN(U3047) );
  NAND2_X1 U5720 ( .A1(n5319), .A2(n7153), .ZN(n5085) );
  NAND2_X1 U5721 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n5320), .ZN(n5084) );
  OAI211_X1 U5722 ( .C1(n5443), .C2(n5643), .A(n5085), .B(n5084), .ZN(n5086)
         );
  AOI21_X1 U5723 ( .B1(n7146), .B2(n5324), .A(n5086), .ZN(n5087) );
  OAI21_X1 U5724 ( .B1(n7156), .B2(n5326), .A(n5087), .ZN(U3044) );
  OR2_X1 U5725 ( .A1(n5129), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5092)
         );
  INV_X1 U5726 ( .A(n5092), .ZN(n5279) );
  AOI22_X1 U5727 ( .A1(n5569), .A2(n7142), .B1(n5130), .B2(n5279), .ZN(n5340)
         );
  NOR2_X1 U5728 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5088), .ZN(n5336)
         );
  NOR2_X1 U5729 ( .A1(n5089), .A2(n4849), .ZN(n5417) );
  OAI22_X1 U5730 ( .A1(n5334), .A2(n5643), .B1(n5333), .B2(n7130), .ZN(n5090)
         );
  AOI21_X1 U5731 ( .B1(n7146), .B2(n5336), .A(n5090), .ZN(n5096) );
  NOR2_X1 U5732 ( .A1(n7142), .A2(n7139), .ZN(n5136) );
  OAI21_X1 U5733 ( .B1(n5198), .B2(n7266), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5091) );
  OAI21_X1 U5734 ( .B1(n5571), .B2(n5136), .A(n5091), .ZN(n5093) );
  NAND2_X1 U5735 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5092), .ZN(n5287) );
  OAI211_X1 U5736 ( .C1(n4629), .C2(n5336), .A(n5093), .B(n5287), .ZN(n5094)
         );
  NAND2_X1 U5737 ( .A1(n5337), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5095) );
  OAI211_X1 U5738 ( .C1(n7156), .C2(n5340), .A(n5096), .B(n5095), .ZN(U3068)
         );
  OAI22_X1 U5739 ( .A1(n5334), .A2(n5659), .B1(n5333), .B2(n7250), .ZN(n5097)
         );
  AOI21_X1 U5740 ( .B1(n7269), .B2(n5336), .A(n5097), .ZN(n5099) );
  NAND2_X1 U5741 ( .A1(n5337), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5098) );
  OAI211_X1 U5742 ( .C1(n7275), .C2(n5340), .A(n5099), .B(n5098), .ZN(U3075)
         );
  OAI22_X1 U5743 ( .A1(n5334), .A2(n5651), .B1(n5333), .B2(n7176), .ZN(n5100)
         );
  AOI21_X1 U5744 ( .B1(n7181), .B2(n5336), .A(n5100), .ZN(n5102) );
  NAND2_X1 U5745 ( .A1(n5337), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5101) );
  OAI211_X1 U5746 ( .C1(n7185), .C2(n5340), .A(n5102), .B(n5101), .ZN(U3070)
         );
  OAI22_X1 U5747 ( .A1(n5334), .A2(n5655), .B1(n5333), .B2(n7190), .ZN(n5103)
         );
  AOI21_X1 U5748 ( .B1(n7195), .B2(n5336), .A(n5103), .ZN(n5105) );
  NAND2_X1 U5749 ( .A1(n5337), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5104) );
  OAI211_X1 U5750 ( .C1(n7199), .C2(n5340), .A(n5105), .B(n5104), .ZN(U3071)
         );
  OAI22_X1 U5751 ( .A1(n5334), .A2(n5647), .B1(n5333), .B2(n7205), .ZN(n5106)
         );
  AOI21_X1 U5752 ( .B1(n7210), .B2(n5336), .A(n5106), .ZN(n5108) );
  NAND2_X1 U5753 ( .A1(n5337), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5107) );
  OAI211_X1 U5754 ( .C1(n7214), .C2(n5340), .A(n5108), .B(n5107), .ZN(U3072)
         );
  INV_X1 U5755 ( .A(EAX_REG_25__SCAN_IN), .ZN(n5115) );
  INV_X1 U5756 ( .A(n7000), .ZN(n5109) );
  NOR2_X1 U5757 ( .A1(n5110), .A2(n5109), .ZN(n5111) );
  NAND2_X1 U5758 ( .A1(n6577), .A2(n5169), .ZN(n5499) );
  OR2_X1 U5759 ( .A1(n7128), .A2(n5113), .ZN(n7027) );
  NOR2_X4 U5762 ( .A1(n6741), .A2(n6577), .ZN(n6590) );
  AOI22_X1 U5763 ( .A1(n6741), .A2(UWORD_REG_9__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n5114) );
  OAI21_X1 U5764 ( .B1(n5115), .B2(n5499), .A(n5114), .ZN(U2898) );
  INV_X1 U5765 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5117) );
  AOI22_X1 U5766 ( .A1(n6741), .A2(UWORD_REG_6__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5116) );
  OAI21_X1 U5767 ( .B1(n5117), .B2(n5499), .A(n5116), .ZN(U2901) );
  AOI22_X1 U5768 ( .A1(n6741), .A2(UWORD_REG_8__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n5118) );
  OAI21_X1 U5769 ( .B1(n4302), .B2(n5499), .A(n5118), .ZN(U2899) );
  AOI22_X1 U5770 ( .A1(n6741), .A2(UWORD_REG_5__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5119) );
  OAI21_X1 U5771 ( .B1(n4261), .B2(n5499), .A(n5119), .ZN(U2902) );
  INV_X1 U5772 ( .A(EAX_REG_23__SCAN_IN), .ZN(n5121) );
  AOI22_X1 U5773 ( .A1(n6741), .A2(UWORD_REG_7__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5120) );
  OAI21_X1 U5774 ( .B1(n5121), .B2(n5499), .A(n5120), .ZN(U2900) );
  AND2_X1 U5775 ( .A1(n5045), .A2(n5122), .ZN(n5124) );
  OR2_X1 U5776 ( .A1(n5124), .A2(n5123), .ZN(n5480) );
  AOI21_X1 U5777 ( .B1(n5126), .B2(n5125), .A(n3471), .ZN(n6777) );
  AOI22_X1 U5778 ( .A1(n6037), .A2(n6777), .B1(n6012), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5127) );
  OAI21_X1 U5779 ( .B1(n5480), .B2(n6039), .A(n5127), .ZN(U2851) );
  OR2_X1 U5780 ( .A1(n5129), .A2(n5128), .ZN(n5137) );
  INV_X1 U5781 ( .A(n5137), .ZN(n5634) );
  AOI22_X1 U5782 ( .A1(n5571), .A2(n7142), .B1(n5130), .B2(n5634), .ZN(n5399)
         );
  NOR2_X1 U5783 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5131), .ZN(n5395)
         );
  OAI22_X1 U5784 ( .A1(n5393), .A2(n7176), .B1(n5392), .B2(n5651), .ZN(n5133)
         );
  AOI21_X1 U5785 ( .B1(n7181), .B2(n5395), .A(n5133), .ZN(n5142) );
  INV_X1 U5786 ( .A(n5393), .ZN(n5134) );
  OAI21_X1 U5787 ( .B1(n5134), .B2(n7243), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5135) );
  OAI21_X1 U5788 ( .B1(n5569), .B2(n5136), .A(n5135), .ZN(n5138) );
  NAND2_X1 U5789 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5137), .ZN(n5639) );
  OAI211_X1 U5790 ( .C1(n4629), .C2(n5395), .A(n5138), .B(n5639), .ZN(n5139)
         );
  NAND2_X1 U5791 ( .A1(n5396), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5141)
         );
  OAI211_X1 U5792 ( .C1(n7185), .C2(n5399), .A(n5142), .B(n5141), .ZN(U3134)
         );
  OAI22_X1 U5793 ( .A1(n5393), .A2(n7250), .B1(n5392), .B2(n5659), .ZN(n5143)
         );
  AOI21_X1 U5794 ( .B1(n7269), .B2(n5395), .A(n5143), .ZN(n5145) );
  NAND2_X1 U5795 ( .A1(n5396), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5144)
         );
  OAI211_X1 U5796 ( .C1(n7275), .C2(n5399), .A(n5145), .B(n5144), .ZN(U3139)
         );
  OAI22_X1 U5797 ( .A1(n5393), .A2(n7205), .B1(n5392), .B2(n5647), .ZN(n5146)
         );
  AOI21_X1 U5798 ( .B1(n7210), .B2(n5395), .A(n5146), .ZN(n5148) );
  NAND2_X1 U5799 ( .A1(n5396), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5147)
         );
  OAI211_X1 U5800 ( .C1(n7214), .C2(n5399), .A(n5148), .B(n5147), .ZN(U3136)
         );
  OAI22_X1 U5801 ( .A1(n5393), .A2(n7130), .B1(n5392), .B2(n5643), .ZN(n5149)
         );
  AOI21_X1 U5802 ( .B1(n7146), .B2(n5395), .A(n5149), .ZN(n5151) );
  NAND2_X1 U5803 ( .A1(n5396), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5150)
         );
  OAI211_X1 U5804 ( .C1(n7156), .C2(n5399), .A(n5151), .B(n5150), .ZN(U3132)
         );
  OAI22_X1 U5805 ( .A1(n5393), .A2(n7190), .B1(n5392), .B2(n5655), .ZN(n5152)
         );
  AOI21_X1 U5806 ( .B1(n7195), .B2(n5395), .A(n5152), .ZN(n5154) );
  NAND2_X1 U5807 ( .A1(n5396), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5153)
         );
  OAI211_X1 U5808 ( .C1(n7199), .C2(n5399), .A(n5154), .B(n5153), .ZN(U3135)
         );
  INV_X1 U5809 ( .A(DATAI_8_), .ZN(n6460) );
  INV_X1 U5810 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6595) );
  OAI222_X1 U5811 ( .A1(n5480), .A2(n7086), .B1(n5745), .B2(n6460), .C1(n5839), 
        .C2(n6595), .ZN(U2883) );
  AND2_X1 U5812 ( .A1(n4343), .A2(n5157), .ZN(n7032) );
  NOR3_X1 U5813 ( .A1(n7046), .A2(n4629), .A3(n7048), .ZN(n7043) );
  OR2_X1 U5814 ( .A1(n7032), .A2(n7043), .ZN(n5158) );
  NOR2_X1 U5815 ( .A1(n6843), .A2(n5158), .ZN(n5159) );
  NAND2_X1 U5816 ( .A1(n6875), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5178) );
  INV_X1 U5817 ( .A(n5178), .ZN(n5161) );
  NAND2_X1 U5818 ( .A1(n7028), .A2(n7126), .ZN(n5168) );
  NAND2_X1 U5819 ( .A1(n5168), .A2(EBX_REG_31__SCAN_IN), .ZN(n5162) );
  NOR2_X1 U5820 ( .A1(n5843), .A2(n5162), .ZN(n5163) );
  INV_X1 U5821 ( .A(n5168), .ZN(n5164) );
  AND3_X1 U5822 ( .A1(n5165), .A2(n5164), .A3(n5169), .ZN(n5166) );
  INV_X1 U5823 ( .A(n6875), .ZN(n5523) );
  AOI22_X1 U5824 ( .A1(n6955), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5523), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n5167) );
  OAI21_X1 U5825 ( .B1(n6905), .B2(REIP_REG_1__SCAN_IN), .A(n5167), .ZN(n5176)
         );
  OR2_X1 U5826 ( .A1(n6730), .A2(n5168), .ZN(n7031) );
  AND2_X1 U5827 ( .A1(n4407), .A2(n7031), .ZN(n5851) );
  INV_X1 U5828 ( .A(n5851), .ZN(n5171) );
  INV_X1 U5829 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6007) );
  NAND3_X1 U5830 ( .A1(n5169), .A2(n6007), .A3(n5168), .ZN(n5170) );
  NAND2_X1 U5831 ( .A1(n5171), .A2(n5170), .ZN(n5172) );
  AND2_X2 U5832 ( .A1(n5852), .A2(n5172), .ZN(n6972) );
  INV_X1 U5833 ( .A(n6972), .ZN(n6933) );
  INV_X1 U5834 ( .A(n5173), .ZN(n6724) );
  NAND2_X1 U5835 ( .A1(n5852), .A2(n6724), .ZN(n6865) );
  OAI22_X1 U5836 ( .A1(n6933), .A2(n4421), .B1(n5174), .B2(n6865), .ZN(n5175)
         );
  AOI211_X1 U5837 ( .C1(n6930), .C2(n5177), .A(n5176), .B(n5175), .ZN(n5183)
         );
  INV_X1 U5838 ( .A(n5852), .ZN(n5180) );
  OAI21_X1 U5839 ( .B1(n5180), .B2(n6714), .A(n6961), .ZN(n6871) );
  NAND2_X1 U5840 ( .A1(n6871), .A2(n5181), .ZN(n5182) );
  OAI211_X1 U5841 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6973), .A(n5183), 
        .B(n5182), .ZN(U2826) );
  NOR2_X2 U5842 ( .A1(n5193), .A2(n5184), .ZN(n7166) );
  INV_X1 U5843 ( .A(n7166), .ZN(n5188) );
  INV_X1 U5844 ( .A(n7170), .ZN(n5185) );
  AOI22_X1 U5845 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5196), .B1(n5185), 
        .B2(n5194), .ZN(n5187) );
  NAND2_X1 U5846 ( .A1(n6710), .A2(DATAI_17_), .ZN(n7161) );
  INV_X1 U5847 ( .A(n7161), .ZN(n7167) );
  NAND2_X1 U5848 ( .A1(n6710), .A2(DATAI_25_), .ZN(n5663) );
  INV_X1 U5849 ( .A(n5663), .ZN(n7165) );
  AOI22_X1 U5850 ( .A1(n7167), .A2(n5198), .B1(n5197), .B2(n7165), .ZN(n5186)
         );
  OAI211_X1 U5851 ( .C1(n5188), .C2(n5201), .A(n5187), .B(n5186), .ZN(U3061)
         );
  NOR2_X2 U5852 ( .A1(n5193), .A2(n3793), .ZN(n7238) );
  INV_X1 U5853 ( .A(n7238), .ZN(n5192) );
  INV_X1 U5854 ( .A(n7242), .ZN(n5189) );
  AOI22_X1 U5855 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5196), .B1(n5189), 
        .B2(n5194), .ZN(n5191) );
  NAND2_X1 U5856 ( .A1(n6710), .A2(DATAI_30_), .ZN(n5667) );
  INV_X1 U5857 ( .A(n5667), .ZN(n7239) );
  NAND2_X1 U5858 ( .A1(n6710), .A2(DATAI_22_), .ZN(n7232) );
  INV_X1 U5859 ( .A(n7232), .ZN(n7237) );
  AOI22_X1 U5860 ( .A1(n7239), .A2(n5197), .B1(n5198), .B2(n7237), .ZN(n5190)
         );
  OAI211_X1 U5861 ( .C1(n5192), .C2(n5201), .A(n5191), .B(n5190), .ZN(U3066)
         );
  NOR2_X2 U5862 ( .A1(n5193), .A2(n3750), .ZN(n7222) );
  INV_X1 U5863 ( .A(n7222), .ZN(n5202) );
  INV_X1 U5864 ( .A(n7226), .ZN(n5195) );
  AOI22_X1 U5865 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5196), .B1(n5195), 
        .B2(n5194), .ZN(n5200) );
  NAND2_X1 U5866 ( .A1(n6710), .A2(DATAI_21_), .ZN(n5583) );
  INV_X1 U5867 ( .A(n5583), .ZN(n7221) );
  NAND2_X1 U5868 ( .A1(n6710), .A2(DATAI_29_), .ZN(n5672) );
  INV_X1 U5869 ( .A(n5672), .ZN(n7223) );
  AOI22_X1 U5870 ( .A1(n7221), .A2(n5198), .B1(n5197), .B2(n7223), .ZN(n5199)
         );
  OAI211_X1 U5871 ( .C1(n5202), .C2(n5201), .A(n5200), .B(n5199), .ZN(U3065)
         );
  NAND2_X1 U5872 ( .A1(n7143), .A2(n3538), .ZN(n5209) );
  NOR3_X2 U5873 ( .A1(n7123), .A2(n5203), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5460) );
  INV_X1 U5874 ( .A(n5460), .ZN(n5204) );
  AOI21_X1 U5875 ( .B1(n5209), .B2(n5204), .A(n7139), .ZN(n5206) );
  NAND3_X1 U5876 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5570), .A3(n7008), .ZN(
        n5212) );
  INV_X1 U5877 ( .A(n5212), .ZN(n5205) );
  NAND2_X1 U5878 ( .A1(n5208), .A2(n5207), .ZN(n5415) );
  INV_X1 U5879 ( .A(n5209), .ZN(n5210) );
  AOI21_X1 U5880 ( .B1(n5214), .B2(STATEBS16_REG_SCAN_IN), .A(n5210), .ZN(
        n5211) );
  OAI22_X1 U5881 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5212), .B1(n5211), .B2(
        n7139), .ZN(n5213) );
  OAI21_X1 U5882 ( .B1(n5460), .B2(n5213), .A(n5285), .ZN(n5457) );
  NAND2_X1 U5883 ( .A1(n5457), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5217) );
  OAI22_X1 U5884 ( .A1(n5604), .A2(n5659), .B1(n5458), .B2(n7250), .ZN(n5215)
         );
  AOI21_X1 U5885 ( .B1(n7269), .B2(n5460), .A(n5215), .ZN(n5216) );
  OAI211_X1 U5886 ( .C1(n5463), .C2(n7275), .A(n5217), .B(n5216), .ZN(U3035)
         );
  NAND2_X1 U5887 ( .A1(n5457), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5220) );
  OAI22_X1 U5888 ( .A1(n5604), .A2(n5647), .B1(n5458), .B2(n7205), .ZN(n5218)
         );
  AOI21_X1 U5889 ( .B1(n7210), .B2(n5460), .A(n5218), .ZN(n5219) );
  OAI211_X1 U5890 ( .C1(n5463), .C2(n7214), .A(n5220), .B(n5219), .ZN(U3032)
         );
  NAND2_X1 U5891 ( .A1(n5457), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5223) );
  OAI22_X1 U5892 ( .A1(n5604), .A2(n5655), .B1(n5458), .B2(n7190), .ZN(n5221)
         );
  AOI21_X1 U5893 ( .B1(n7195), .B2(n5460), .A(n5221), .ZN(n5222) );
  OAI211_X1 U5894 ( .C1(n5463), .C2(n7199), .A(n5223), .B(n5222), .ZN(U3031)
         );
  NAND2_X1 U5895 ( .A1(n5457), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n5226) );
  OAI22_X1 U5896 ( .A1(n5604), .A2(n5651), .B1(n5458), .B2(n7176), .ZN(n5224)
         );
  AOI21_X1 U5897 ( .B1(n7181), .B2(n5460), .A(n5224), .ZN(n5225) );
  OAI211_X1 U5898 ( .C1(n5463), .C2(n7185), .A(n5226), .B(n5225), .ZN(U3030)
         );
  NAND2_X1 U5899 ( .A1(n5457), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n5229) );
  OAI22_X1 U5900 ( .A1(n5604), .A2(n5643), .B1(n5458), .B2(n7130), .ZN(n5227)
         );
  AOI21_X1 U5901 ( .B1(n7146), .B2(n5460), .A(n5227), .ZN(n5228) );
  OAI211_X1 U5902 ( .C1(n5463), .C2(n7156), .A(n5229), .B(n5228), .ZN(U3028)
         );
  AOI22_X1 U5903 ( .A1(n5269), .A2(EAX_REG_10__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n5231) );
  NAND2_X1 U5904 ( .A1(n5232), .A2(n5231), .ZN(U2949) );
  OR2_X1 U5905 ( .A1(n5277), .A2(n5233), .ZN(n5246) );
  AOI22_X1 U5906 ( .A1(n5275), .A2(EAX_REG_2__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n5234) );
  NAND2_X1 U5907 ( .A1(n5246), .A2(n5234), .ZN(U2941) );
  NAND2_X1 U5908 ( .A1(n5255), .A2(DATAI_3_), .ZN(n5248) );
  AOI22_X1 U5909 ( .A1(n5275), .A2(EAX_REG_3__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U5910 ( .A1(n5248), .A2(n5235), .ZN(U2942) );
  INV_X1 U5911 ( .A(DATAI_4_), .ZN(n5464) );
  OR2_X1 U5912 ( .A1(n5277), .A2(n5464), .ZN(n5250) );
  AOI22_X1 U5913 ( .A1(n5275), .A2(EAX_REG_4__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U5914 ( .A1(n5250), .A2(n5236), .ZN(U2943) );
  INV_X1 U5915 ( .A(DATAI_5_), .ZN(n5465) );
  OR2_X1 U5916 ( .A1(n5277), .A2(n5465), .ZN(n5252) );
  AOI22_X1 U5917 ( .A1(n5275), .A2(EAX_REG_5__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U5918 ( .A1(n5252), .A2(n5237), .ZN(U2944) );
  AOI22_X1 U5919 ( .A1(n5275), .A2(EAX_REG_6__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U5920 ( .A1(n5239), .A2(n5238), .ZN(U2945) );
  OR2_X1 U5921 ( .A1(n5277), .A2(n5240), .ZN(n5258) );
  AOI22_X1 U5922 ( .A1(n5275), .A2(EAX_REG_16__SCAN_IN), .B1(n5274), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n5241) );
  NAND2_X1 U5923 ( .A1(n5258), .A2(n5241), .ZN(U2924) );
  NAND2_X1 U5924 ( .A1(n5255), .A2(DATAI_1_), .ZN(n5262) );
  AOI22_X1 U5925 ( .A1(n5275), .A2(EAX_REG_17__SCAN_IN), .B1(n5274), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U5926 ( .A1(n5262), .A2(n5242), .ZN(U2925) );
  AOI22_X1 U5927 ( .A1(n5275), .A2(EAX_REG_9__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n5243) );
  NAND2_X1 U5928 ( .A1(n5244), .A2(n5243), .ZN(U2948) );
  AOI22_X1 U5929 ( .A1(n5275), .A2(EAX_REG_18__SCAN_IN), .B1(n5274), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U5930 ( .A1(n5246), .A2(n5245), .ZN(U2926) );
  AOI22_X1 U5931 ( .A1(n5275), .A2(EAX_REG_19__SCAN_IN), .B1(n5274), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U5932 ( .A1(n5248), .A2(n5247), .ZN(U2927) );
  AOI22_X1 U5933 ( .A1(n5275), .A2(EAX_REG_20__SCAN_IN), .B1(n5274), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U5934 ( .A1(n5250), .A2(n5249), .ZN(U2928) );
  AOI22_X1 U5935 ( .A1(n5275), .A2(EAX_REG_21__SCAN_IN), .B1(n5274), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U5936 ( .A1(n5252), .A2(n5251), .ZN(U2929) );
  NAND2_X1 U5937 ( .A1(n5255), .A2(DATAI_12_), .ZN(n5266) );
  AOI22_X1 U5938 ( .A1(n5275), .A2(EAX_REG_28__SCAN_IN), .B1(n5274), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U5939 ( .A1(n5266), .A2(n5253), .ZN(U2936) );
  NAND2_X1 U5940 ( .A1(n5255), .A2(DATAI_13_), .ZN(n5268) );
  AOI22_X1 U5941 ( .A1(n5275), .A2(EAX_REG_29__SCAN_IN), .B1(n5274), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U5942 ( .A1(n5268), .A2(n5254), .ZN(U2937) );
  NAND2_X1 U5943 ( .A1(n5255), .A2(DATAI_14_), .ZN(n5271) );
  AOI22_X1 U5944 ( .A1(n5275), .A2(EAX_REG_30__SCAN_IN), .B1(n5274), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n5256) );
  NAND2_X1 U5945 ( .A1(n5271), .A2(n5256), .ZN(U2938) );
  AOI22_X1 U5946 ( .A1(n5275), .A2(EAX_REG_0__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U5947 ( .A1(n5258), .A2(n5257), .ZN(U2939) );
  AOI22_X1 U5948 ( .A1(n5275), .A2(EAX_REG_8__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U5949 ( .A1(n5260), .A2(n5259), .ZN(U2947) );
  AOI22_X1 U5950 ( .A1(n5275), .A2(EAX_REG_1__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U5951 ( .A1(n5262), .A2(n5261), .ZN(U2940) );
  AOI22_X1 U5952 ( .A1(n5269), .A2(EAX_REG_11__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n5263) );
  NAND2_X1 U5953 ( .A1(n5264), .A2(n5263), .ZN(U2950) );
  AOI22_X1 U5954 ( .A1(n5269), .A2(EAX_REG_12__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n5265) );
  NAND2_X1 U5955 ( .A1(n5266), .A2(n5265), .ZN(U2951) );
  AOI22_X1 U5956 ( .A1(n5269), .A2(EAX_REG_13__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U5957 ( .A1(n5268), .A2(n5267), .ZN(U2952) );
  AOI22_X1 U5958 ( .A1(n5269), .A2(EAX_REG_14__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U5959 ( .A1(n5271), .A2(n5270), .ZN(U2953) );
  AOI22_X1 U5960 ( .A1(n5275), .A2(EAX_REG_7__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U5961 ( .A1(n5273), .A2(n5272), .ZN(U2946) );
  INV_X1 U5962 ( .A(DATAI_15_), .ZN(n5744) );
  AOI22_X1 U5963 ( .A1(n5275), .A2(EAX_REG_15__SCAN_IN), .B1(n5274), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n5276) );
  OAI21_X1 U5964 ( .B1(n5277), .B2(n5744), .A(n5276), .ZN(U2954) );
  INV_X1 U5965 ( .A(n5278), .ZN(n5635) );
  AOI22_X1 U5966 ( .A1(n5569), .A2(n3537), .B1(n5635), .B2(n5279), .ZN(n5448)
         );
  AOI21_X1 U5967 ( .B1(n5458), .B2(n5443), .A(n5280), .ZN(n5281) );
  AOI21_X1 U5968 ( .B1(n5282), .B2(n3537), .A(n5281), .ZN(n5283) );
  NOR2_X1 U5969 ( .A1(n5283), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5288) );
  NOR2_X1 U5970 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5284), .ZN(n5445)
         );
  NAND2_X1 U5971 ( .A1(n5442), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5291) );
  OAI22_X1 U5972 ( .A1(n5458), .A2(n5655), .B1(n5443), .B2(n7190), .ZN(n5289)
         );
  AOI21_X1 U5973 ( .B1(n7195), .B2(n5445), .A(n5289), .ZN(n5290) );
  OAI211_X1 U5974 ( .C1(n5448), .C2(n7199), .A(n5291), .B(n5290), .ZN(U3039)
         );
  NAND2_X1 U5975 ( .A1(n5442), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5294) );
  OAI22_X1 U5976 ( .A1(n5458), .A2(n5651), .B1(n5443), .B2(n7176), .ZN(n5292)
         );
  AOI21_X1 U5977 ( .B1(n7181), .B2(n5445), .A(n5292), .ZN(n5293) );
  OAI211_X1 U5978 ( .C1(n5448), .C2(n7185), .A(n5294), .B(n5293), .ZN(U3038)
         );
  NAND2_X1 U5979 ( .A1(n5442), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5297) );
  OAI22_X1 U5980 ( .A1(n5458), .A2(n5643), .B1(n5443), .B2(n7130), .ZN(n5295)
         );
  AOI21_X1 U5981 ( .B1(n7146), .B2(n5445), .A(n5295), .ZN(n5296) );
  OAI211_X1 U5982 ( .C1(n5448), .C2(n7156), .A(n5297), .B(n5296), .ZN(U3036)
         );
  NAND2_X1 U5983 ( .A1(n5442), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5300) );
  OAI22_X1 U5984 ( .A1(n5458), .A2(n5659), .B1(n5443), .B2(n7250), .ZN(n5298)
         );
  AOI21_X1 U5985 ( .B1(n7269), .B2(n5445), .A(n5298), .ZN(n5299) );
  OAI211_X1 U5986 ( .C1(n5448), .C2(n7275), .A(n5300), .B(n5299), .ZN(U3043)
         );
  NAND2_X1 U5987 ( .A1(n5442), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5303) );
  OAI22_X1 U5988 ( .A1(n5458), .A2(n5647), .B1(n5443), .B2(n7205), .ZN(n5301)
         );
  AOI21_X1 U5989 ( .B1(n7210), .B2(n5445), .A(n5301), .ZN(n5302) );
  OAI211_X1 U5990 ( .C1(n5448), .C2(n7214), .A(n5303), .B(n5302), .ZN(U3040)
         );
  NOR2_X1 U5991 ( .A1(n5123), .A2(n5305), .ZN(n5306) );
  OR2_X1 U5992 ( .A1(n5304), .A2(n5306), .ZN(n5550) );
  INV_X1 U5993 ( .A(n5307), .ZN(n5308) );
  XNOR2_X1 U5994 ( .A(n5309), .B(n5308), .ZN(n6810) );
  AOI22_X1 U5995 ( .A1(n6037), .A2(n6810), .B1(n6012), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n5310) );
  OAI21_X1 U5996 ( .B1(n5550), .B2(n6039), .A(n5310), .ZN(U2850) );
  NAND2_X1 U5997 ( .A1(n5319), .A2(n7237), .ZN(n5312) );
  NAND2_X1 U5998 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n5320), .ZN(n5311) );
  OAI211_X1 U5999 ( .C1(n5443), .C2(n5667), .A(n5312), .B(n5311), .ZN(n5313)
         );
  AOI21_X1 U6000 ( .B1(n7238), .B2(n5324), .A(n5313), .ZN(n5314) );
  OAI21_X1 U6001 ( .B1(n7242), .B2(n5326), .A(n5314), .ZN(U3050) );
  NAND2_X1 U6002 ( .A1(n5319), .A2(n7167), .ZN(n5316) );
  NAND2_X1 U6003 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n5320), .ZN(n5315) );
  OAI211_X1 U6004 ( .C1(n5443), .C2(n5663), .A(n5316), .B(n5315), .ZN(n5317)
         );
  AOI21_X1 U6005 ( .B1(n7166), .B2(n5324), .A(n5317), .ZN(n5318) );
  OAI21_X1 U6006 ( .B1(n7170), .B2(n5326), .A(n5318), .ZN(U3045) );
  NAND2_X1 U6007 ( .A1(n5319), .A2(n7221), .ZN(n5322) );
  NAND2_X1 U6008 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n5320), .ZN(n5321) );
  OAI211_X1 U6009 ( .C1(n5443), .C2(n5672), .A(n5322), .B(n5321), .ZN(n5323)
         );
  AOI21_X1 U6010 ( .B1(n7222), .B2(n5324), .A(n5323), .ZN(n5325) );
  OAI21_X1 U6011 ( .B1(n7226), .B2(n5326), .A(n5325), .ZN(U3049) );
  OAI22_X1 U6012 ( .A1(n5334), .A2(n5667), .B1(n5333), .B2(n7232), .ZN(n5327)
         );
  AOI21_X1 U6013 ( .B1(n7238), .B2(n5336), .A(n5327), .ZN(n5329) );
  NAND2_X1 U6014 ( .A1(n5337), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5328) );
  OAI211_X1 U6015 ( .C1(n7242), .C2(n5340), .A(n5329), .B(n5328), .ZN(U3074)
         );
  OAI22_X1 U6016 ( .A1(n5334), .A2(n5663), .B1(n5333), .B2(n7161), .ZN(n5330)
         );
  AOI21_X1 U6017 ( .B1(n7166), .B2(n5336), .A(n5330), .ZN(n5332) );
  NAND2_X1 U6018 ( .A1(n5337), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5331) );
  OAI211_X1 U6019 ( .C1(n7170), .C2(n5340), .A(n5332), .B(n5331), .ZN(U3069)
         );
  OAI22_X1 U6020 ( .A1(n5334), .A2(n5672), .B1(n5333), .B2(n5583), .ZN(n5335)
         );
  AOI21_X1 U6021 ( .B1(n7222), .B2(n5336), .A(n5335), .ZN(n5339) );
  NAND2_X1 U6022 ( .A1(n5337), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5338) );
  OAI211_X1 U6023 ( .C1(n7226), .C2(n5340), .A(n5339), .B(n5338), .ZN(U3073)
         );
  NAND2_X1 U6024 ( .A1(n5373), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5343)
         );
  OAI22_X1 U6025 ( .A1(n7251), .A2(n5667), .B1(n7108), .B2(n7232), .ZN(n5341)
         );
  AOI21_X1 U6026 ( .B1(n7238), .B2(n5375), .A(n5341), .ZN(n5342) );
  OAI211_X1 U6027 ( .C1(n5378), .C2(n7242), .A(n5343), .B(n5342), .ZN(U3122)
         );
  NAND2_X1 U6028 ( .A1(n5367), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5346)
         );
  OAI22_X1 U6029 ( .A1(n7161), .A2(n5603), .B1(n5393), .B2(n5663), .ZN(n5344)
         );
  AOI21_X1 U6030 ( .B1(n7166), .B2(n5369), .A(n5344), .ZN(n5345) );
  OAI211_X1 U6031 ( .C1(n5372), .C2(n7170), .A(n5346), .B(n5345), .ZN(U3141)
         );
  NAND2_X1 U6032 ( .A1(n5359), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5349) );
  OAI22_X1 U6033 ( .A1(n5361), .A2(n7232), .B1(n5667), .B2(n5360), .ZN(n5347)
         );
  AOI21_X1 U6034 ( .B1(n7238), .B2(n5363), .A(n5347), .ZN(n5348) );
  OAI211_X1 U6035 ( .C1(n5366), .C2(n7242), .A(n5349), .B(n5348), .ZN(U3058)
         );
  NAND2_X1 U6036 ( .A1(n5373), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5352)
         );
  OAI22_X1 U6037 ( .A1(n7251), .A2(n5663), .B1(n7108), .B2(n7161), .ZN(n5350)
         );
  AOI21_X1 U6038 ( .B1(n7166), .B2(n5375), .A(n5350), .ZN(n5351) );
  OAI211_X1 U6039 ( .C1(n5378), .C2(n7170), .A(n5352), .B(n5351), .ZN(U3117)
         );
  NAND2_X1 U6040 ( .A1(n5359), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5355) );
  OAI22_X1 U6041 ( .A1(n5361), .A2(n7161), .B1(n5663), .B2(n5360), .ZN(n5353)
         );
  AOI21_X1 U6042 ( .B1(n7166), .B2(n5363), .A(n5353), .ZN(n5354) );
  OAI211_X1 U6043 ( .C1(n5366), .C2(n7170), .A(n5355), .B(n5354), .ZN(U3053)
         );
  NAND2_X1 U6044 ( .A1(n5367), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5358)
         );
  OAI22_X1 U6045 ( .A1(n5603), .A2(n7232), .B1(n5393), .B2(n5667), .ZN(n5356)
         );
  AOI21_X1 U6046 ( .B1(n7238), .B2(n5369), .A(n5356), .ZN(n5357) );
  OAI211_X1 U6047 ( .C1(n5372), .C2(n7242), .A(n5358), .B(n5357), .ZN(U3146)
         );
  NAND2_X1 U6048 ( .A1(n5359), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5365) );
  OAI22_X1 U6049 ( .A1(n5361), .A2(n5583), .B1(n5672), .B2(n5360), .ZN(n5362)
         );
  AOI21_X1 U6050 ( .B1(n7222), .B2(n5363), .A(n5362), .ZN(n5364) );
  OAI211_X1 U6051 ( .C1(n5366), .C2(n7226), .A(n5365), .B(n5364), .ZN(U3057)
         );
  NAND2_X1 U6052 ( .A1(n5367), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5371)
         );
  OAI22_X1 U6053 ( .A1(n5603), .A2(n5583), .B1(n5393), .B2(n5672), .ZN(n5368)
         );
  AOI21_X1 U6054 ( .B1(n7222), .B2(n5369), .A(n5368), .ZN(n5370) );
  OAI211_X1 U6055 ( .C1(n5372), .C2(n7226), .A(n5371), .B(n5370), .ZN(U3145)
         );
  NAND2_X1 U6056 ( .A1(n5373), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5377)
         );
  OAI22_X1 U6057 ( .A1(n7251), .A2(n5672), .B1(n7108), .B2(n5583), .ZN(n5374)
         );
  AOI21_X1 U6058 ( .B1(n7222), .B2(n5375), .A(n5374), .ZN(n5376) );
  OAI211_X1 U6059 ( .C1(n5378), .C2(n7226), .A(n5377), .B(n5376), .ZN(U3121)
         );
  XNOR2_X1 U6060 ( .A(n5379), .B(n5380), .ZN(n6750) );
  INV_X1 U6061 ( .A(n6858), .ZN(n5384) );
  NAND2_X1 U6062 ( .A1(n6843), .A2(REIP_REG_4__SCAN_IN), .ZN(n6749) );
  INV_X1 U6063 ( .A(n6749), .ZN(n5381) );
  AOI21_X1 U6064 ( .B1(n6691), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n5381), 
        .ZN(n5382) );
  OAI21_X1 U6065 ( .B1(n6707), .B2(n6857), .A(n5382), .ZN(n5383) );
  AOI21_X1 U6066 ( .B1(n6710), .B2(n5384), .A(n5383), .ZN(n5385) );
  OAI21_X1 U6067 ( .B1(n6750), .B2(n6993), .A(n5385), .ZN(U2982) );
  OAI22_X1 U6068 ( .A1(n5393), .A2(n7161), .B1(n5392), .B2(n5663), .ZN(n5386)
         );
  AOI21_X1 U6069 ( .B1(n7166), .B2(n5395), .A(n5386), .ZN(n5388) );
  NAND2_X1 U6070 ( .A1(n5396), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5387)
         );
  OAI211_X1 U6071 ( .C1(n7170), .C2(n5399), .A(n5388), .B(n5387), .ZN(U3133)
         );
  OAI22_X1 U6072 ( .A1(n5393), .A2(n7232), .B1(n5392), .B2(n5667), .ZN(n5389)
         );
  AOI21_X1 U6073 ( .B1(n7238), .B2(n5395), .A(n5389), .ZN(n5391) );
  NAND2_X1 U6074 ( .A1(n5396), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5390)
         );
  OAI211_X1 U6075 ( .C1(n7242), .C2(n5399), .A(n5391), .B(n5390), .ZN(U3138)
         );
  OAI22_X1 U6076 ( .A1(n5393), .A2(n5583), .B1(n5392), .B2(n5672), .ZN(n5394)
         );
  AOI21_X1 U6077 ( .B1(n7222), .B2(n5395), .A(n5394), .ZN(n5398) );
  NAND2_X1 U6078 ( .A1(n5396), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5397)
         );
  OAI211_X1 U6079 ( .C1(n7226), .C2(n5399), .A(n5398), .B(n5397), .ZN(U3137)
         );
  NAND2_X1 U6080 ( .A1(n5442), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5402) );
  OAI22_X1 U6081 ( .A1(n5458), .A2(n5667), .B1(n5443), .B2(n7232), .ZN(n5400)
         );
  AOI21_X1 U6082 ( .B1(n7238), .B2(n5445), .A(n5400), .ZN(n5401) );
  OAI211_X1 U6083 ( .C1(n5448), .C2(n7242), .A(n5402), .B(n5401), .ZN(U3042)
         );
  NAND2_X1 U6084 ( .A1(n5442), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5405) );
  OAI22_X1 U6085 ( .A1(n5458), .A2(n5663), .B1(n5443), .B2(n7161), .ZN(n5403)
         );
  AOI21_X1 U6086 ( .B1(n7166), .B2(n5445), .A(n5403), .ZN(n5404) );
  OAI211_X1 U6087 ( .C1(n5448), .C2(n7170), .A(n5405), .B(n5404), .ZN(U3037)
         );
  NAND2_X1 U6088 ( .A1(n5457), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n5408) );
  OAI22_X1 U6089 ( .A1(n7161), .A2(n5458), .B1(n5604), .B2(n5663), .ZN(n5406)
         );
  AOI21_X1 U6090 ( .B1(n7166), .B2(n5460), .A(n5406), .ZN(n5407) );
  OAI211_X1 U6091 ( .C1(n5463), .C2(n7170), .A(n5408), .B(n5407), .ZN(U3029)
         );
  NAND2_X1 U6092 ( .A1(n5457), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5411) );
  OAI22_X1 U6093 ( .A1(n5604), .A2(n5667), .B1(n5458), .B2(n7232), .ZN(n5409)
         );
  AOI21_X1 U6094 ( .B1(n7238), .B2(n5460), .A(n5409), .ZN(n5410) );
  OAI211_X1 U6095 ( .C1(n5463), .C2(n7242), .A(n5411), .B(n5410), .ZN(U3034)
         );
  AOI22_X1 U6096 ( .A1(n5571), .A2(n3538), .B1(n5635), .B2(n5412), .ZN(n5456)
         );
  NAND3_X1 U6097 ( .A1(n7012), .A2(n7008), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7133) );
  NOR2_X1 U6098 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7133), .ZN(n5453)
         );
  INV_X1 U6099 ( .A(n5453), .ZN(n5414) );
  AOI21_X1 U6100 ( .B1(n5414), .B2(STATE2_REG_3__SCAN_IN), .A(n5413), .ZN(
        n5420) );
  NOR2_X1 U6101 ( .A1(n3538), .A2(n7139), .ZN(n5572) );
  INV_X1 U6102 ( .A(n5415), .ZN(n5416) );
  OAI21_X1 U6103 ( .B1(n7259), .B2(n7270), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5418) );
  OAI21_X1 U6104 ( .B1(n5569), .B2(n5572), .A(n5418), .ZN(n5419) );
  NAND3_X1 U6105 ( .A1(n5641), .A2(n5420), .A3(n5419), .ZN(n5449) );
  NAND2_X1 U6106 ( .A1(n5449), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5423) );
  OAI22_X1 U6107 ( .A1(n5451), .A2(n7161), .B1(n5450), .B2(n5663), .ZN(n5421)
         );
  AOI21_X1 U6108 ( .B1(n7166), .B2(n5453), .A(n5421), .ZN(n5422) );
  OAI211_X1 U6109 ( .C1(n7170), .C2(n5456), .A(n5423), .B(n5422), .ZN(U3085)
         );
  NAND2_X1 U6110 ( .A1(n5449), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5426) );
  OAI22_X1 U6111 ( .A1(n5451), .A2(n7205), .B1(n5450), .B2(n5647), .ZN(n5424)
         );
  AOI21_X1 U6112 ( .B1(n7210), .B2(n5453), .A(n5424), .ZN(n5425) );
  OAI211_X1 U6113 ( .C1(n7214), .C2(n5456), .A(n5426), .B(n5425), .ZN(U3088)
         );
  NAND2_X1 U6114 ( .A1(n5449), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5429) );
  OAI22_X1 U6115 ( .A1(n5451), .A2(n7232), .B1(n5450), .B2(n5667), .ZN(n5427)
         );
  AOI21_X1 U6116 ( .B1(n7238), .B2(n5453), .A(n5427), .ZN(n5428) );
  OAI211_X1 U6117 ( .C1(n7242), .C2(n5456), .A(n5429), .B(n5428), .ZN(U3090)
         );
  NAND2_X1 U6118 ( .A1(n5449), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5432) );
  OAI22_X1 U6119 ( .A1(n5451), .A2(n7250), .B1(n5450), .B2(n5659), .ZN(n5430)
         );
  AOI21_X1 U6120 ( .B1(n7269), .B2(n5453), .A(n5430), .ZN(n5431) );
  OAI211_X1 U6121 ( .C1(n7275), .C2(n5456), .A(n5432), .B(n5431), .ZN(U3091)
         );
  NAND2_X1 U6122 ( .A1(n5449), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5435) );
  OAI22_X1 U6123 ( .A1(n5451), .A2(n7176), .B1(n5450), .B2(n5651), .ZN(n5433)
         );
  AOI21_X1 U6124 ( .B1(n7181), .B2(n5453), .A(n5433), .ZN(n5434) );
  OAI211_X1 U6125 ( .C1(n7185), .C2(n5456), .A(n5435), .B(n5434), .ZN(U3086)
         );
  NAND2_X1 U6126 ( .A1(n5449), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5438) );
  OAI22_X1 U6127 ( .A1(n5450), .A2(n5643), .B1(n7130), .B2(n5451), .ZN(n5436)
         );
  AOI21_X1 U6128 ( .B1(n7146), .B2(n5453), .A(n5436), .ZN(n5437) );
  OAI211_X1 U6129 ( .C1(n7156), .C2(n5456), .A(n5438), .B(n5437), .ZN(U3084)
         );
  NAND2_X1 U6130 ( .A1(n5449), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5441) );
  OAI22_X1 U6131 ( .A1(n5451), .A2(n7190), .B1(n5450), .B2(n5655), .ZN(n5439)
         );
  AOI21_X1 U6132 ( .B1(n7195), .B2(n5453), .A(n5439), .ZN(n5440) );
  OAI211_X1 U6133 ( .C1(n7199), .C2(n5456), .A(n5441), .B(n5440), .ZN(U3087)
         );
  NAND2_X1 U6134 ( .A1(n5442), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5447) );
  OAI22_X1 U6135 ( .A1(n5458), .A2(n5672), .B1(n5443), .B2(n5583), .ZN(n5444)
         );
  AOI21_X1 U6136 ( .B1(n7222), .B2(n5445), .A(n5444), .ZN(n5446) );
  OAI211_X1 U6137 ( .C1(n5448), .C2(n7226), .A(n5447), .B(n5446), .ZN(U3041)
         );
  NAND2_X1 U6138 ( .A1(n5449), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5455) );
  OAI22_X1 U6139 ( .A1(n5451), .A2(n5583), .B1(n5450), .B2(n5672), .ZN(n5452)
         );
  AOI21_X1 U6140 ( .B1(n7222), .B2(n5453), .A(n5452), .ZN(n5454) );
  OAI211_X1 U6141 ( .C1(n7226), .C2(n5456), .A(n5455), .B(n5454), .ZN(U3089)
         );
  NAND2_X1 U6142 ( .A1(n5457), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n5462) );
  OAI22_X1 U6143 ( .A1(n5604), .A2(n5672), .B1(n5458), .B2(n5583), .ZN(n5459)
         );
  AOI21_X1 U6144 ( .B1(n7222), .B2(n5460), .A(n5459), .ZN(n5461) );
  OAI211_X1 U6145 ( .C1(n5463), .C2(n7226), .A(n5462), .B(n5461), .ZN(U3033)
         );
  INV_X1 U6146 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6587) );
  OAI222_X1 U6147 ( .A1(n6858), .A2(n7086), .B1(n5745), .B2(n5464), .C1(n5839), 
        .C2(n6587), .ZN(U2887) );
  INV_X1 U6148 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6589) );
  OAI222_X1 U6149 ( .A1(n5466), .A2(n7086), .B1(n5745), .B2(n5465), .C1(n5839), 
        .C2(n6589), .ZN(U2886) );
  INV_X1 U6150 ( .A(DATAI_1_), .ZN(n6417) );
  INV_X1 U6151 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6581) );
  OAI222_X1 U6152 ( .A1(n5467), .A2(n7086), .B1(n5745), .B2(n6417), .C1(n5839), 
        .C2(n6581), .ZN(U2890) );
  INV_X1 U6153 ( .A(DATAI_9_), .ZN(n6457) );
  INV_X1 U6154 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6597) );
  OAI222_X1 U6155 ( .A1(n5550), .A2(n7086), .B1(n5745), .B2(n6457), .C1(n5839), 
        .C2(n6597), .ZN(U2882) );
  INV_X1 U6156 ( .A(DATAI_7_), .ZN(n6464) );
  OAI222_X1 U6157 ( .A1(n5468), .A2(n7086), .B1(n5745), .B2(n6464), .C1(n5839), 
        .C2(n4031), .ZN(U2884) );
  INV_X1 U6158 ( .A(n6871), .ZN(n6859) );
  NAND2_X1 U6159 ( .A1(n6905), .A2(n6875), .ZN(n5964) );
  NAND2_X1 U6160 ( .A1(n6972), .A2(EBX_REG_0__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U6161 ( .A1(n6930), .A2(n5469), .ZN(n5470) );
  OAI211_X1 U6162 ( .C1(n5472), .C2(n6865), .A(n5471), .B(n5470), .ZN(n5473)
         );
  AOI21_X1 U6163 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5964), .A(n5473), .ZN(n5475)
         );
  OAI21_X1 U6164 ( .B1(n6950), .B2(n6955), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5474) );
  OAI211_X1 U6165 ( .C1(n6859), .C2(n5476), .A(n5475), .B(n5474), .ZN(U2827)
         );
  OAI21_X1 U6166 ( .B1(n5479), .B2(n5478), .A(n5477), .ZN(n6782) );
  INV_X1 U6167 ( .A(n5480), .ZN(n5508) );
  NAND2_X1 U6168 ( .A1(n6843), .A2(REIP_REG_8__SCAN_IN), .ZN(n6775) );
  NAND2_X1 U6169 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5481)
         );
  OAI211_X1 U6170 ( .C1(n6707), .C2(n5502), .A(n6775), .B(n5481), .ZN(n5482)
         );
  AOI21_X1 U6171 ( .B1(n5508), .B2(n6710), .A(n5482), .ZN(n5483) );
  OAI21_X1 U6172 ( .B1(n6782), .B2(n6993), .A(n5483), .ZN(U2978) );
  INV_X1 U6173 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5485) );
  AOI22_X1 U6174 ( .A1(n6741), .A2(UWORD_REG_3__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5484) );
  OAI21_X1 U6175 ( .B1(n5485), .B2(n5499), .A(n5484), .ZN(U2904) );
  INV_X1 U6176 ( .A(EAX_REG_20__SCAN_IN), .ZN(n5487) );
  AOI22_X1 U6177 ( .A1(n6741), .A2(UWORD_REG_4__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5486) );
  OAI21_X1 U6178 ( .B1(n5487), .B2(n5499), .A(n5486), .ZN(U2903) );
  INV_X1 U6179 ( .A(EAX_REG_28__SCAN_IN), .ZN(n5489) );
  AOI22_X1 U6180 ( .A1(n6741), .A2(UWORD_REG_12__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n5488) );
  OAI21_X1 U6181 ( .B1(n5489), .B2(n5499), .A(n5488), .ZN(U2895) );
  AOI22_X1 U6182 ( .A1(n6741), .A2(UWORD_REG_1__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5490) );
  OAI21_X1 U6183 ( .B1(n4189), .B2(n5499), .A(n5490), .ZN(U2906) );
  AOI22_X1 U6184 ( .A1(n6741), .A2(UWORD_REG_13__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n5491) );
  OAI21_X1 U6185 ( .B1(n3693), .B2(n5499), .A(n5491), .ZN(U2894) );
  INV_X1 U6186 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5493) );
  AOI22_X1 U6187 ( .A1(n6741), .A2(UWORD_REG_2__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5492) );
  OAI21_X1 U6188 ( .B1(n5493), .B2(n5499), .A(n5492), .ZN(U2905) );
  AOI22_X1 U6189 ( .A1(n6741), .A2(UWORD_REG_11__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5494) );
  OAI21_X1 U6190 ( .B1(n4330), .B2(n5499), .A(n5494), .ZN(U2896) );
  INV_X1 U6191 ( .A(EAX_REG_16__SCAN_IN), .ZN(n5496) );
  AOI22_X1 U6192 ( .A1(n6741), .A2(UWORD_REG_0__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5495) );
  OAI21_X1 U6193 ( .B1(n5496), .B2(n5499), .A(n5495), .ZN(U2907) );
  AOI22_X1 U6194 ( .A1(n6741), .A2(UWORD_REG_14__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5497) );
  OAI21_X1 U6195 ( .B1(n4661), .B2(n5499), .A(n5497), .ZN(U2893) );
  INV_X1 U6196 ( .A(EAX_REG_26__SCAN_IN), .ZN(n5500) );
  AOI22_X1 U6197 ( .A1(n6741), .A2(UWORD_REG_10__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n5498) );
  OAI21_X1 U6198 ( .B1(n5500), .B2(n5499), .A(n5498), .ZN(U2897) );
  NAND3_X1 U6199 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n6853) );
  INV_X1 U6200 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6855) );
  NOR2_X1 U6201 ( .A1(n6853), .A2(n6855), .ZN(n6872) );
  NAND2_X1 U6202 ( .A1(n6872), .A2(REIP_REG_5__SCAN_IN), .ZN(n6874) );
  INV_X1 U6203 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6891) );
  INV_X1 U6204 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6620) );
  NOR3_X1 U6205 ( .A1(n6874), .A2(n6891), .A3(n6620), .ZN(n5501) );
  NAND2_X1 U6206 ( .A1(n5501), .A2(REIP_REG_8__SCAN_IN), .ZN(n5539) );
  INV_X1 U6207 ( .A(n5539), .ZN(n5552) );
  OAI21_X1 U6208 ( .B1(n6905), .B2(n5552), .A(n6875), .ZN(n5556) );
  INV_X1 U6209 ( .A(n5556), .ZN(n5534) );
  INV_X1 U6210 ( .A(n6905), .ZN(n5990) );
  AOI21_X1 U6211 ( .B1(n5990), .B2(n5501), .A(REIP_REG_8__SCAN_IN), .ZN(n5503)
         );
  OAI22_X1 U6212 ( .A1(n5534), .A2(n5503), .B1(n5502), .B2(n6973), .ZN(n5507)
         );
  AOI22_X1 U6213 ( .A1(EBX_REG_8__SCAN_IN), .A2(n6972), .B1(n6930), .B2(n6777), 
        .ZN(n5504) );
  INV_X1 U6214 ( .A(n6954), .ZN(n6912) );
  OAI211_X1 U6215 ( .C1(n6981), .C2(n5505), .A(n5504), .B(n6912), .ZN(n5506)
         );
  AOI211_X1 U6216 ( .C1(n5508), .C2(n6978), .A(n5507), .B(n5506), .ZN(n5509)
         );
  INV_X1 U6217 ( .A(n5509), .ZN(U2819) );
  INV_X1 U6218 ( .A(n6865), .ZN(n5529) );
  AOI22_X1 U6219 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6955), .B1(
        EBX_REG_3__SCAN_IN), .B2(n6972), .ZN(n5512) );
  INV_X1 U6220 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U6221 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n5519) );
  OAI21_X1 U6222 ( .B1(n5523), .B2(n6853), .A(n5964), .ZN(n6854) );
  AOI221_X1 U6223 ( .B1(n5523), .B2(n6614), .C1(n5519), .C2(n6614), .A(n6854), 
        .ZN(n5510) );
  INV_X1 U6224 ( .A(n5510), .ZN(n5511) );
  OAI211_X1 U6225 ( .C1(n6975), .C2(n5513), .A(n5512), .B(n5511), .ZN(n5514)
         );
  AOI21_X1 U6226 ( .B1(n5529), .B2(n3444), .A(n5514), .ZN(n5517) );
  NAND2_X1 U6227 ( .A1(n6871), .A2(n5515), .ZN(n5516) );
  OAI211_X1 U6228 ( .C1(n6973), .C2(n5518), .A(n5517), .B(n5516), .ZN(U2824)
         );
  NOR2_X1 U6229 ( .A1(n6973), .A2(n6690), .ZN(n5528) );
  NAND2_X1 U6230 ( .A1(n6972), .A2(EBX_REG_2__SCAN_IN), .ZN(n5525) );
  OAI211_X1 U6231 ( .C1(REIP_REG_2__SCAN_IN), .C2(REIP_REG_1__SCAN_IN), .A(
        n5990), .B(n5519), .ZN(n5520) );
  OAI21_X1 U6232 ( .B1(n5521), .B2(n6975), .A(n5520), .ZN(n5522) );
  AOI21_X1 U6233 ( .B1(n5523), .B2(REIP_REG_2__SCAN_IN), .A(n5522), .ZN(n5524)
         );
  OAI211_X1 U6234 ( .C1(n6981), .C2(n5526), .A(n5525), .B(n5524), .ZN(n5527)
         );
  AOI211_X1 U6235 ( .C1(n5529), .C2(n3447), .A(n5528), .B(n5527), .ZN(n5530)
         );
  OAI21_X1 U6236 ( .B1(n6859), .B2(n6684), .A(n5530), .ZN(U2825) );
  NOR2_X1 U6237 ( .A1(n5304), .A2(n5532), .ZN(n5533) );
  OR2_X1 U6238 ( .A1(n5531), .A2(n5533), .ZN(n5681) );
  OAI21_X1 U6239 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6905), .A(n5534), .ZN(n5546)
         );
  OR2_X1 U6240 ( .A1(n5536), .A2(n5535), .ZN(n5537) );
  NAND2_X1 U6241 ( .A1(n5565), .A2(n5537), .ZN(n5548) );
  OAI22_X1 U6242 ( .A1(n5538), .A2(n6933), .B1(n6975), .B2(n5548), .ZN(n5543)
         );
  INV_X1 U6243 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6802) );
  INV_X1 U6244 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6623) );
  NOR2_X1 U6245 ( .A1(n5539), .A2(n6623), .ZN(n5620) );
  NAND3_X1 U6246 ( .A1(n5990), .A2(n6802), .A3(n5620), .ZN(n5540) );
  OAI211_X1 U6247 ( .C1(n6981), .C2(n5541), .A(n6912), .B(n5540), .ZN(n5542)
         );
  NOR2_X1 U6248 ( .A1(n5543), .A2(n5542), .ZN(n5544) );
  OAI21_X1 U6249 ( .B1(n6973), .B2(n5683), .A(n5544), .ZN(n5545) );
  AOI21_X1 U6250 ( .B1(n5546), .B2(REIP_REG_10__SCAN_IN), .A(n5545), .ZN(n5547) );
  OAI21_X1 U6251 ( .B1(n5681), .B2(n6961), .A(n5547), .ZN(U2817) );
  INV_X1 U6252 ( .A(n5548), .ZN(n6799) );
  AOI22_X1 U6253 ( .A1(n6037), .A2(n6799), .B1(n6012), .B2(EBX_REG_10__SCAN_IN), .ZN(n5549) );
  OAI21_X1 U6254 ( .B1(n5681), .B2(n6039), .A(n5549), .ZN(U2849) );
  INV_X1 U6255 ( .A(n5550), .ZN(n5616) );
  INV_X1 U6256 ( .A(n5551), .ZN(n5614) );
  NAND2_X1 U6257 ( .A1(n6930), .A2(n6810), .ZN(n5555) );
  NAND2_X1 U6258 ( .A1(n5552), .A2(n6623), .ZN(n5553) );
  OR2_X1 U6259 ( .A1(n6905), .A2(n5553), .ZN(n5554) );
  OAI211_X1 U6260 ( .C1(n6973), .C2(n5614), .A(n5555), .B(n5554), .ZN(n5560)
         );
  INV_X1 U6261 ( .A(EBX_REG_9__SCAN_IN), .ZN(n5558) );
  AOI22_X1 U6262 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6955), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5556), .ZN(n5557) );
  OAI211_X1 U6263 ( .C1(n6933), .C2(n5558), .A(n5557), .B(n6912), .ZN(n5559)
         );
  AOI211_X1 U6264 ( .C1(n5616), .C2(n6978), .A(n5560), .B(n5559), .ZN(n5561)
         );
  INV_X1 U6265 ( .A(n5561), .ZN(U2818) );
  INV_X1 U6266 ( .A(DATAI_10_), .ZN(n6419) );
  INV_X1 U6267 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6599) );
  OAI222_X1 U6268 ( .A1(n5681), .A2(n7086), .B1(n5745), .B2(n6419), .C1(n5839), 
        .C2(n6599), .ZN(U2881) );
  OAI21_X1 U6269 ( .B1(n5531), .B2(n5563), .A(n5619), .ZN(n6708) );
  INV_X1 U6270 ( .A(n5564), .ZN(n5710) );
  AOI21_X1 U6271 ( .B1(n5566), .B2(n5565), .A(n5710), .ZN(n6903) );
  AOI22_X1 U6272 ( .A1(n6037), .A2(n6903), .B1(EBX_REG_11__SCAN_IN), .B2(n6012), .ZN(n5567) );
  OAI21_X1 U6273 ( .B1(n6708), .B2(n6039), .A(n5567), .ZN(U2848) );
  AOI22_X1 U6274 ( .A1(n5569), .A2(n3538), .B1(n5635), .B2(n5568), .ZN(n5609)
         );
  NAND3_X1 U6275 ( .A1(n7008), .A2(n7123), .A3(n5570), .ZN(n5579) );
  INV_X1 U6276 ( .A(n5571), .ZN(n5575) );
  INV_X1 U6277 ( .A(n5572), .ZN(n5574) );
  AOI21_X1 U6278 ( .B1(n5604), .B2(n5603), .A(n7126), .ZN(n5573) );
  AOI21_X1 U6279 ( .B1(n5575), .B2(n5574), .A(n5573), .ZN(n5576) );
  AOI211_X1 U6280 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5579), .A(n5577), .B(
        n5576), .ZN(n5578) );
  NAND2_X1 U6281 ( .A1(n5641), .A2(n5578), .ZN(n5602) );
  NAND2_X1 U6282 ( .A1(n5602), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5582) );
  INV_X1 U6283 ( .A(n5579), .ZN(n5606) );
  OAI22_X1 U6284 ( .A1(n5604), .A2(n7232), .B1(n5603), .B2(n5667), .ZN(n5580)
         );
  AOI21_X1 U6285 ( .B1(n7238), .B2(n5606), .A(n5580), .ZN(n5581) );
  OAI211_X1 U6286 ( .C1(n5609), .C2(n7242), .A(n5582), .B(n5581), .ZN(U3026)
         );
  NAND2_X1 U6287 ( .A1(n5602), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5586) );
  OAI22_X1 U6288 ( .A1(n5604), .A2(n5583), .B1(n5603), .B2(n5672), .ZN(n5584)
         );
  AOI21_X1 U6289 ( .B1(n7222), .B2(n5606), .A(n5584), .ZN(n5585) );
  OAI211_X1 U6290 ( .C1(n5609), .C2(n7226), .A(n5586), .B(n5585), .ZN(U3025)
         );
  NAND2_X1 U6291 ( .A1(n5602), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5589) );
  OAI22_X1 U6292 ( .A1(n5604), .A2(n7205), .B1(n5603), .B2(n5647), .ZN(n5587)
         );
  AOI21_X1 U6293 ( .B1(n7210), .B2(n5606), .A(n5587), .ZN(n5588) );
  OAI211_X1 U6294 ( .C1(n5609), .C2(n7214), .A(n5589), .B(n5588), .ZN(U3024)
         );
  NAND2_X1 U6295 ( .A1(n5602), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5592) );
  OAI22_X1 U6296 ( .A1(n5604), .A2(n7190), .B1(n5603), .B2(n5655), .ZN(n5590)
         );
  AOI21_X1 U6297 ( .B1(n7195), .B2(n5606), .A(n5590), .ZN(n5591) );
  OAI211_X1 U6298 ( .C1(n5609), .C2(n7199), .A(n5592), .B(n5591), .ZN(U3023)
         );
  NAND2_X1 U6299 ( .A1(n5602), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5595) );
  OAI22_X1 U6300 ( .A1(n5604), .A2(n7161), .B1(n5603), .B2(n5663), .ZN(n5593)
         );
  AOI21_X1 U6301 ( .B1(n7166), .B2(n5606), .A(n5593), .ZN(n5594) );
  OAI211_X1 U6302 ( .C1(n5609), .C2(n7170), .A(n5595), .B(n5594), .ZN(U3021)
         );
  NAND2_X1 U6303 ( .A1(n5602), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5598) );
  OAI22_X1 U6304 ( .A1(n5604), .A2(n7130), .B1(n5603), .B2(n5643), .ZN(n5596)
         );
  AOI21_X1 U6305 ( .B1(n7146), .B2(n5606), .A(n5596), .ZN(n5597) );
  OAI211_X1 U6306 ( .C1(n5609), .C2(n7156), .A(n5598), .B(n5597), .ZN(U3020)
         );
  NAND2_X1 U6307 ( .A1(n5602), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5601) );
  OAI22_X1 U6308 ( .A1(n5604), .A2(n7250), .B1(n5603), .B2(n5659), .ZN(n5599)
         );
  AOI21_X1 U6309 ( .B1(n7269), .B2(n5606), .A(n5599), .ZN(n5600) );
  OAI211_X1 U6310 ( .C1(n5609), .C2(n7275), .A(n5601), .B(n5600), .ZN(U3027)
         );
  NAND2_X1 U6311 ( .A1(n5602), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5608) );
  OAI22_X1 U6312 ( .A1(n5604), .A2(n7176), .B1(n5603), .B2(n5651), .ZN(n5605)
         );
  AOI21_X1 U6313 ( .B1(n7181), .B2(n5606), .A(n5605), .ZN(n5607) );
  OAI211_X1 U6314 ( .C1(n5609), .C2(n7185), .A(n5608), .B(n5607), .ZN(U3022)
         );
  OAI21_X1 U6315 ( .B1(n5612), .B2(n5611), .A(n5610), .ZN(n6808) );
  AOI22_X1 U6316 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n6843), 
        .B2(REIP_REG_9__SCAN_IN), .ZN(n5613) );
  OAI21_X1 U6317 ( .B1(n6707), .B2(n5614), .A(n5613), .ZN(n5615) );
  AOI21_X1 U6318 ( .B1(n5616), .B2(n6710), .A(n5615), .ZN(n5617) );
  OAI21_X1 U6319 ( .B1(n6808), .B2(n6993), .A(n5617), .ZN(U2977) );
  INV_X1 U6320 ( .A(DATAI_11_), .ZN(n6321) );
  INV_X1 U6321 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6601) );
  OAI222_X1 U6322 ( .A1(n6708), .A2(n7086), .B1(n5745), .B2(n6321), .C1(n5839), 
        .C2(n6601), .ZN(U2880) );
  XNOR2_X1 U6323 ( .A(n5619), .B(n5618), .ZN(n5729) );
  INV_X1 U6324 ( .A(n5725), .ZN(n5627) );
  XNOR2_X1 U6325 ( .A(n5710), .B(n5709), .ZN(n6814) );
  NAND2_X1 U6326 ( .A1(n5620), .A2(REIP_REG_10__SCAN_IN), .ZN(n6904) );
  INV_X1 U6327 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6907) );
  NOR2_X1 U6328 ( .A1(n6904), .A2(n6907), .ZN(n5737) );
  INV_X1 U6329 ( .A(n5737), .ZN(n5621) );
  OR2_X1 U6330 ( .A1(n6905), .A2(n5621), .ZN(n6931) );
  NOR2_X1 U6331 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6931), .ZN(n6924) );
  INV_X1 U6332 ( .A(n6924), .ZN(n5622) );
  OAI211_X1 U6333 ( .C1(n6975), .C2(n6814), .A(n6912), .B(n5622), .ZN(n5626)
         );
  OAI21_X1 U6334 ( .B1(n6905), .B2(n5737), .A(n6875), .ZN(n6923) );
  AOI22_X1 U6335 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6972), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6923), .ZN(n5623) );
  OAI21_X1 U6336 ( .B1(n5624), .B2(n6981), .A(n5623), .ZN(n5625) );
  AOI211_X1 U6337 ( .C1(n6950), .C2(n5627), .A(n5626), .B(n5625), .ZN(n5628)
         );
  OAI21_X1 U6338 ( .B1(n5729), .B2(n6961), .A(n5628), .ZN(U2815) );
  INV_X1 U6339 ( .A(n7254), .ZN(n5631) );
  NAND3_X1 U6340 ( .A1(n7233), .A2(n7152), .A3(n5631), .ZN(n5633) );
  NAND2_X1 U6341 ( .A1(n5633), .A2(n5632), .ZN(n5637) );
  NAND3_X1 U6342 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n7012), .ZN(n7113) );
  INV_X1 U6343 ( .A(n7113), .ZN(n7120) );
  NAND2_X1 U6344 ( .A1(n7123), .A2(n7120), .ZN(n5638) );
  INV_X1 U6345 ( .A(n5638), .ZN(n5674) );
  INV_X1 U6346 ( .A(n7114), .ZN(n5636) );
  AOI22_X1 U6347 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5638), .B1(n5637), .B2(
        n5636), .ZN(n5640) );
  NAND3_X1 U6348 ( .A1(n5641), .A2(n5640), .A3(n5639), .ZN(n5670) );
  AOI22_X1 U6349 ( .A1(n7254), .A2(n7153), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5670), .ZN(n5642) );
  OAI21_X1 U6350 ( .B1(n5643), .B2(n7233), .A(n5642), .ZN(n5644) );
  AOI21_X1 U6351 ( .B1(n7146), .B2(n5674), .A(n5644), .ZN(n5645) );
  OAI21_X1 U6352 ( .B1(n7156), .B2(n5676), .A(n5645), .ZN(U3100) );
  AOI22_X1 U6353 ( .A1(n7254), .A2(n7209), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5670), .ZN(n5646) );
  OAI21_X1 U6354 ( .B1(n5647), .B2(n7233), .A(n5646), .ZN(n5648) );
  AOI21_X1 U6355 ( .B1(n7210), .B2(n5674), .A(n5648), .ZN(n5649) );
  OAI21_X1 U6356 ( .B1(n7214), .B2(n5676), .A(n5649), .ZN(U3104) );
  AOI22_X1 U6357 ( .A1(n7254), .A2(n7180), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5670), .ZN(n5650) );
  OAI21_X1 U6358 ( .B1(n5651), .B2(n7233), .A(n5650), .ZN(n5652) );
  AOI21_X1 U6359 ( .B1(n7181), .B2(n5674), .A(n5652), .ZN(n5653) );
  OAI21_X1 U6360 ( .B1(n7185), .B2(n5676), .A(n5653), .ZN(U3102) );
  AOI22_X1 U6361 ( .A1(n7254), .A2(n7196), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5670), .ZN(n5654) );
  OAI21_X1 U6362 ( .B1(n5655), .B2(n7233), .A(n5654), .ZN(n5656) );
  AOI21_X1 U6363 ( .B1(n7195), .B2(n5674), .A(n5656), .ZN(n5657) );
  OAI21_X1 U6364 ( .B1(n7199), .B2(n5676), .A(n5657), .ZN(U3103) );
  AOI22_X1 U6365 ( .A1(n7254), .A2(n7271), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5670), .ZN(n5658) );
  OAI21_X1 U6366 ( .B1(n5659), .B2(n7233), .A(n5658), .ZN(n5660) );
  AOI21_X1 U6367 ( .B1(n7269), .B2(n5674), .A(n5660), .ZN(n5661) );
  OAI21_X1 U6368 ( .B1(n7275), .B2(n5676), .A(n5661), .ZN(U3107) );
  AOI22_X1 U6369 ( .A1(n7254), .A2(n7167), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5670), .ZN(n5662) );
  OAI21_X1 U6370 ( .B1(n5663), .B2(n7233), .A(n5662), .ZN(n5664) );
  AOI21_X1 U6371 ( .B1(n7166), .B2(n5674), .A(n5664), .ZN(n5665) );
  OAI21_X1 U6372 ( .B1(n7170), .B2(n5676), .A(n5665), .ZN(U3101) );
  AOI22_X1 U6373 ( .A1(n7254), .A2(n7237), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5670), .ZN(n5666) );
  OAI21_X1 U6374 ( .B1(n5667), .B2(n7233), .A(n5666), .ZN(n5668) );
  AOI21_X1 U6375 ( .B1(n7238), .B2(n5674), .A(n5668), .ZN(n5669) );
  OAI21_X1 U6376 ( .B1(n7242), .B2(n5676), .A(n5669), .ZN(U3106) );
  AOI22_X1 U6377 ( .A1(n7254), .A2(n7221), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5670), .ZN(n5671) );
  OAI21_X1 U6378 ( .B1(n5672), .B2(n7233), .A(n5671), .ZN(n5673) );
  AOI21_X1 U6379 ( .B1(n7222), .B2(n5674), .A(n5673), .ZN(n5675) );
  OAI21_X1 U6380 ( .B1(n7226), .B2(n5676), .A(n5675), .ZN(U3105) );
  NAND2_X1 U6381 ( .A1(n5679), .A2(n5678), .ZN(n5680) );
  XNOR2_X1 U6382 ( .A(n5677), .B(n5680), .ZN(n6798) );
  INV_X1 U6383 ( .A(n6798), .ZN(n5687) );
  INV_X1 U6384 ( .A(n5681), .ZN(n5685) );
  AOI22_X1 U6385 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6843), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5682) );
  OAI21_X1 U6386 ( .B1(n6707), .B2(n5683), .A(n5682), .ZN(n5684) );
  AOI21_X1 U6387 ( .B1(n5685), .B2(n6710), .A(n5684), .ZN(n5686) );
  OAI21_X1 U6388 ( .B1(n5687), .B2(n6993), .A(n5686), .ZN(U2976) );
  INV_X1 U6389 ( .A(DATAI_12_), .ZN(n6320) );
  OAI222_X1 U6390 ( .A1(n7086), .A2(n5729), .B1(n5745), .B2(n6320), .C1(n5839), 
        .C2(n4093), .ZN(U2879) );
  INV_X1 U6391 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5688) );
  OAI222_X1 U6392 ( .A1(n6047), .A2(n5688), .B1(n6045), .B2(n6814), .C1(n6039), 
        .C2(n5729), .ZN(U2847) );
  NAND2_X1 U6393 ( .A1(n5690), .A2(n5689), .ZN(n5692) );
  XOR2_X1 U6394 ( .A(n5692), .B(n3436), .Z(n6713) );
  NAND3_X1 U6395 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6765), .ZN(n6785) );
  INV_X1 U6396 ( .A(n6785), .ZN(n6780) );
  NAND2_X1 U6397 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6795) );
  INV_X1 U6398 ( .A(n6795), .ZN(n6797) );
  NAND4_X1 U6399 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6780), .A4(n6797), .ZN(n5694)
         );
  NOR2_X1 U6400 ( .A1(n5693), .A2(n5694), .ZN(n5790) );
  NOR2_X1 U6401 ( .A1(n6745), .A2(n5694), .ZN(n5786) );
  INV_X1 U6402 ( .A(n5786), .ZN(n5695) );
  AOI21_X1 U6403 ( .B1(n6525), .B2(n5695), .A(n5788), .ZN(n6528) );
  OAI21_X1 U6404 ( .B1(n6744), .B2(n5790), .A(n6528), .ZN(n6823) );
  INV_X1 U6405 ( .A(n5753), .ZN(n5700) );
  INV_X1 U6406 ( .A(n5790), .ZN(n5699) );
  OR3_X1 U6407 ( .A1(n5697), .A2(n5696), .A3(n5695), .ZN(n5698) );
  OAI21_X1 U6408 ( .B1(n5699), .B2(n6744), .A(n5698), .ZN(n5767) );
  AOI21_X1 U6409 ( .B1(n5700), .B2(n5786), .A(n5767), .ZN(n6304) );
  INV_X1 U6410 ( .A(n6304), .ZN(n6819) );
  AOI22_X1 U6411 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6823), .B1(n6819), .B2(n5701), .ZN(n5702) );
  OAI21_X1 U6412 ( .B1(n6801), .B2(n6907), .A(n5702), .ZN(n5703) );
  AOI21_X1 U6413 ( .B1(n6846), .B2(n6903), .A(n5703), .ZN(n5704) );
  OAI21_X1 U6414 ( .B1(n6713), .B2(n6756), .A(n5704), .ZN(U3007) );
  OAI21_X1 U6415 ( .B1(n5705), .B2(n5707), .A(n5706), .ZN(n6919) );
  AOI21_X1 U6416 ( .B1(n5710), .B2(n5709), .A(n5708), .ZN(n5712) );
  INV_X1 U6417 ( .A(n5717), .ZN(n5711) );
  NOR2_X1 U6418 ( .A1(n5712), .A2(n5711), .ZN(n6916) );
  AOI22_X1 U6419 ( .A1(n6037), .A2(n6916), .B1(EBX_REG_13__SCAN_IN), .B2(n6012), .ZN(n5713) );
  OAI21_X1 U6420 ( .B1(n6919), .B2(n6039), .A(n5713), .ZN(U2846) );
  OAI21_X1 U6421 ( .B1(n5714), .B2(n5716), .A(n5715), .ZN(n6937) );
  AOI21_X1 U6422 ( .B1(n5718), .B2(n5717), .A(n5734), .ZN(n6929) );
  AOI22_X1 U6423 ( .A1(n6037), .A2(n6929), .B1(n6012), .B2(EBX_REG_14__SCAN_IN), .ZN(n5719) );
  OAI21_X1 U6424 ( .B1(n6937), .B2(n6039), .A(n5719), .ZN(U2845) );
  INV_X1 U6425 ( .A(DATAI_14_), .ZN(n6449) );
  OAI222_X1 U6426 ( .A1(n6937), .A2(n7086), .B1(n5745), .B2(n6449), .C1(n5839), 
        .C2(n4130), .ZN(U2877) );
  INV_X1 U6427 ( .A(DATAI_13_), .ZN(n6452) );
  INV_X1 U6428 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6604) );
  OAI222_X1 U6429 ( .A1(n6919), .A2(n7086), .B1(n5745), .B2(n6452), .C1(n5839), 
        .C2(n6604), .ZN(U2878) );
  INV_X1 U6430 ( .A(n5721), .ZN(n5723) );
  NAND2_X1 U6431 ( .A1(n5723), .A2(n5722), .ZN(n5724) );
  XNOR2_X1 U6432 ( .A(n5720), .B(n5724), .ZN(n6817) );
  INV_X1 U6433 ( .A(n6993), .ZN(n6704) );
  NAND2_X1 U6434 ( .A1(n6817), .A2(n6704), .ZN(n5728) );
  AND2_X1 U6435 ( .A1(n6843), .A2(REIP_REG_12__SCAN_IN), .ZN(n6815) );
  NOR2_X1 U6436 ( .A1(n6707), .A2(n5725), .ZN(n5726) );
  AOI211_X1 U6437 ( .C1(n6691), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6815), 
        .B(n5726), .ZN(n5727) );
  OAI211_X1 U6438 ( .C1(n5729), .C2(n6685), .A(n5728), .B(n5727), .ZN(U2974)
         );
  INV_X1 U6439 ( .A(n5715), .ZN(n5732) );
  OAI21_X1 U6440 ( .B1(n5732), .B2(n4161), .A(n5731), .ZN(n6203) );
  INV_X1 U6441 ( .A(n6199), .ZN(n5742) );
  INV_X1 U6442 ( .A(n6042), .ZN(n5733) );
  OAI21_X1 U6443 ( .B1(n5735), .B2(n5734), .A(n5733), .ZN(n6826) );
  AOI21_X1 U6444 ( .B1(n6955), .B2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6954), 
        .ZN(n5736) );
  OAI21_X1 U6445 ( .B1(n6975), .B2(n6826), .A(n5736), .ZN(n5741) );
  NAND4_X1 U6446 ( .A1(n5737), .A2(REIP_REG_12__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_14__SCAN_IN), .ZN(n5822) );
  NOR2_X1 U6447 ( .A1(n6905), .A2(n5822), .ZN(n6945) );
  INV_X1 U6448 ( .A(n6945), .ZN(n5998) );
  INV_X1 U6449 ( .A(n5822), .ZN(n5738) );
  OAI21_X1 U6450 ( .B1(n6905), .B2(n5738), .A(n6875), .ZN(n6943) );
  AOI22_X1 U6451 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6972), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6943), .ZN(n5739) );
  OAI21_X1 U6452 ( .B1(REIP_REG_15__SCAN_IN), .B2(n5998), .A(n5739), .ZN(n5740) );
  AOI211_X1 U6453 ( .C1(n6950), .C2(n5742), .A(n5741), .B(n5740), .ZN(n5743)
         );
  OAI21_X1 U6454 ( .B1(n6203), .B2(n6961), .A(n5743), .ZN(U2812) );
  INV_X1 U6455 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6609) );
  OAI222_X1 U6456 ( .A1(n6203), .A2(n7086), .B1(n5745), .B2(n5744), .C1(n5839), 
        .C2(n6609), .ZN(U2876) );
  INV_X1 U6457 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5746) );
  OAI222_X1 U6458 ( .A1(n6203), .A2(n6039), .B1(n6047), .B2(n5746), .C1(n6045), 
        .C2(n6826), .ZN(U2844) );
  OAI21_X1 U6459 ( .B1(n5749), .B2(n5748), .A(n5747), .ZN(n5757) );
  INV_X1 U6460 ( .A(n5757), .ZN(n5756) );
  NAND2_X1 U6461 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6818) );
  NOR2_X1 U6462 ( .A1(n5750), .A2(n6818), .ZN(n5785) );
  AOI21_X1 U6463 ( .B1(n5751), .B2(n6818), .A(n6823), .ZN(n5752) );
  OAI21_X1 U6464 ( .B1(n5785), .B2(n5753), .A(n5752), .ZN(n5766) );
  NOR2_X1 U6465 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6818), .ZN(n5768)
         );
  AOI22_X1 U6466 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5766), .B1(n5768), .B2(n6819), .ZN(n5755) );
  AND2_X1 U6467 ( .A1(n6843), .A2(REIP_REG_13__SCAN_IN), .ZN(n5759) );
  AOI21_X1 U6468 ( .B1(n6846), .B2(n6916), .A(n5759), .ZN(n5754) );
  OAI211_X1 U6469 ( .C1(n5756), .C2(n6756), .A(n5755), .B(n5754), .ZN(U3005)
         );
  NAND2_X1 U6470 ( .A1(n5757), .A2(n6704), .ZN(n5761) );
  NOR2_X1 U6471 ( .A1(n6707), .A2(n6920), .ZN(n5758) );
  AOI211_X1 U6472 ( .C1(n6691), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5759), 
        .B(n5758), .ZN(n5760) );
  OAI211_X1 U6473 ( .C1(n6685), .C2(n6919), .A(n5761), .B(n5760), .ZN(U2973)
         );
  XNOR2_X1 U6474 ( .A(n6137), .B(n5769), .ZN(n5763) );
  XNOR2_X1 U6475 ( .A(n5762), .B(n5763), .ZN(n6209) );
  NAND2_X1 U6476 ( .A1(n6843), .A2(REIP_REG_14__SCAN_IN), .ZN(n6204) );
  NOR2_X1 U6477 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6304), .ZN(n5764)
         );
  NAND2_X1 U6478 ( .A1(n5785), .A2(n5764), .ZN(n5765) );
  NAND2_X1 U6479 ( .A1(n6204), .A2(n5765), .ZN(n5772) );
  AOI21_X1 U6480 ( .B1(n5768), .B2(n5767), .A(n5766), .ZN(n5770) );
  NOR2_X1 U6481 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  AOI211_X1 U6482 ( .C1(n6846), .C2(n6929), .A(n5772), .B(n5771), .ZN(n5773)
         );
  OAI21_X1 U6483 ( .B1(n6209), .B2(n6756), .A(n5773), .ZN(U3004) );
  OAI21_X1 U6484 ( .B1(n5775), .B2(n5777), .A(n5776), .ZN(n6185) );
  NAND2_X1 U6485 ( .A1(n6044), .A2(n5778), .ZN(n5779) );
  AND2_X1 U6486 ( .A1(n6032), .A2(n5779), .ZN(n6845) );
  AOI22_X1 U6487 ( .A1(n6845), .A2(n6037), .B1(n6012), .B2(EBX_REG_17__SCAN_IN), .ZN(n5780) );
  OAI21_X1 U6488 ( .B1(n6185), .B2(n6039), .A(n5780), .ZN(U2842) );
  NAND2_X1 U6489 ( .A1(n5783), .A2(n6171), .ZN(n5781) );
  OAI21_X1 U6490 ( .B1(n5783), .B2(n5782), .A(n5781), .ZN(n5784) );
  XNOR2_X1 U6491 ( .A(n5784), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5820)
         );
  INV_X1 U6492 ( .A(n5834), .ZN(n5813) );
  NOR2_X1 U6493 ( .A1(n6841), .A2(n6832), .ZN(n6305) );
  INV_X1 U6494 ( .A(n6305), .ZN(n6834) );
  NAND2_X1 U6495 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5785), .ZN(n6824) );
  NOR2_X1 U6496 ( .A1(n6834), .A2(n6824), .ZN(n6529) );
  AND2_X1 U6497 ( .A1(n5786), .A2(n6529), .ZN(n5787) );
  INV_X1 U6498 ( .A(n5791), .ZN(n6306) );
  NAND2_X1 U6499 ( .A1(n5787), .A2(n6306), .ZN(n5805) );
  AND2_X1 U6500 ( .A1(n6525), .A2(n5805), .ZN(n5789) );
  OR2_X1 U6501 ( .A1(n5789), .A2(n5788), .ZN(n5793) );
  NAND2_X1 U6502 ( .A1(n6529), .A2(n5790), .ZN(n6526) );
  NOR2_X1 U6503 ( .A1(n5791), .A2(n6526), .ZN(n5806) );
  NOR2_X1 U6504 ( .A1(n6744), .A2(n5806), .ZN(n5792) );
  NOR2_X1 U6505 ( .A1(n5793), .A2(n5792), .ZN(n6302) );
  NAND2_X1 U6506 ( .A1(n6302), .A2(n6308), .ZN(n5796) );
  INV_X1 U6507 ( .A(n5793), .ZN(n5794) );
  NAND2_X1 U6508 ( .A1(n5794), .A2(n6779), .ZN(n5795) );
  NAND2_X1 U6509 ( .A1(n5796), .A2(n5795), .ZN(n6294) );
  INV_X1 U6510 ( .A(n5797), .ZN(n5798) );
  NAND2_X1 U6511 ( .A1(n6825), .A2(n5798), .ZN(n5799) );
  NAND2_X1 U6512 ( .A1(n6294), .A2(n5799), .ZN(n6281) );
  INV_X1 U6513 ( .A(n5800), .ZN(n5801) );
  AOI21_X1 U6514 ( .B1(n6746), .B2(n6744), .A(n5801), .ZN(n5802) );
  NAND2_X1 U6515 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6249) );
  AND2_X1 U6516 ( .A1(n6825), .A2(n6249), .ZN(n5803) );
  NOR2_X1 U6517 ( .A1(n6266), .A2(n5803), .ZN(n6237) );
  NAND2_X1 U6518 ( .A1(n6825), .A2(n5810), .ZN(n5804) );
  NAND2_X1 U6519 ( .A1(n6237), .A2(n5804), .ZN(n6211) );
  INV_X1 U6520 ( .A(n6211), .ZN(n6225) );
  INV_X1 U6521 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U6522 ( .A1(n6843), .A2(REIP_REG_30__SCAN_IN), .ZN(n5815) );
  OR2_X1 U6523 ( .A1(n6746), .A2(n5805), .ZN(n5808) );
  NAND2_X1 U6524 ( .A1(n6768), .A2(n5806), .ZN(n5807) );
  NAND2_X1 U6525 ( .A1(n5808), .A2(n5807), .ZN(n6288) );
  NAND2_X1 U6526 ( .A1(n6288), .A2(n5809), .ZN(n6262) );
  NOR2_X1 U6527 ( .A1(n6262), .A2(n6249), .ZN(n6232) );
  INV_X1 U6528 ( .A(n5810), .ZN(n6213) );
  NAND3_X1 U6529 ( .A1(n6232), .A2(n6213), .A3(n6212), .ZN(n5811) );
  OAI211_X1 U6530 ( .C1(n6225), .C2(n6212), .A(n5815), .B(n5811), .ZN(n5812)
         );
  AOI21_X1 U6531 ( .B1(n5813), .B2(n6846), .A(n5812), .ZN(n5814) );
  OAI21_X1 U6532 ( .B1(n5820), .B2(n6756), .A(n5814), .ZN(U2988) );
  NAND2_X1 U6533 ( .A1(n5829), .A2(n6709), .ZN(n5816) );
  OAI211_X1 U6534 ( .C1(n5817), .C2(n6205), .A(n5816), .B(n5815), .ZN(n5818)
         );
  AOI21_X1 U6535 ( .B1(n5821), .B2(n6710), .A(n5818), .ZN(n5819) );
  OAI21_X1 U6536 ( .B1(n5820), .B2(n6993), .A(n5819), .ZN(U2956) );
  INV_X1 U6537 ( .A(REIP_REG_30__SCAN_IN), .ZN(n5855) );
  INV_X1 U6538 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6655) );
  NOR2_X1 U6539 ( .A1(n5855), .A2(n6655), .ZN(n5826) );
  AND2_X1 U6540 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5828) );
  INV_X1 U6541 ( .A(n5828), .ZN(n5823) );
  INV_X1 U6542 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6643) );
  INV_X1 U6543 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6641) );
  INV_X1 U6544 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6638) );
  NAND2_X1 U6545 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n6944) );
  INV_X1 U6546 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6633) );
  NOR3_X1 U6547 ( .A1(n5822), .A2(n6944), .A3(n6633), .ZN(n5991) );
  NAND4_X1 U6548 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_20__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5991), .ZN(n5962) );
  NOR2_X1 U6549 ( .A1(n6638), .A2(n5962), .ZN(n5956) );
  NAND2_X1 U6550 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5956), .ZN(n5941) );
  NOR2_X1 U6551 ( .A1(n6641), .A2(n5941), .ZN(n5927) );
  NAND2_X1 U6552 ( .A1(n5927), .A2(n6875), .ZN(n5926) );
  OR2_X1 U6553 ( .A1(n6643), .A2(n5926), .ZN(n5918) );
  NOR2_X1 U6554 ( .A1(n5823), .A2(n5918), .ZN(n5889) );
  AND2_X1 U6555 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5824) );
  NAND2_X1 U6556 ( .A1(n5889), .A2(n5824), .ZN(n5825) );
  NAND2_X1 U6557 ( .A1(n5964), .A2(n5825), .ZN(n5875) );
  OAI21_X1 U6558 ( .B1(n5826), .B2(n6905), .A(n5875), .ZN(n5858) );
  NAND2_X1 U6559 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5927), .ZN(n5827) );
  NOR2_X1 U6560 ( .A1(n6905), .A2(n5827), .ZN(n5903) );
  NAND2_X1 U6561 ( .A1(n5903), .A2(n5828), .ZN(n5891) );
  INV_X1 U6562 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6649) );
  INV_X1 U6563 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U6564 ( .A1(n5855), .A2(REIP_REG_29__SCAN_IN), .ZN(n5833) );
  AOI22_X1 U6565 ( .A1(n6972), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6955), .ZN(n5832) );
  INV_X1 U6566 ( .A(n5829), .ZN(n5830) );
  OR2_X1 U6567 ( .A1(n6973), .A2(n5830), .ZN(n5831) );
  OAI211_X1 U6568 ( .C1(n5862), .C2(n5833), .A(n5832), .B(n5831), .ZN(n5835)
         );
  AOI22_X1 U6569 ( .A1(n7093), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n7096), .ZN(n5841) );
  AND2_X1 U6570 ( .A1(n3750), .A2(n5837), .ZN(n5838) );
  NAND2_X1 U6571 ( .A1(n7097), .A2(DATAI_14_), .ZN(n5840) );
  OAI211_X1 U6572 ( .C1(n5842), .C2(n7086), .A(n5841), .B(n5840), .ZN(U2861)
         );
  OAI22_X1 U6573 ( .A1(n5844), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5843), .ZN(n5849) );
  OAI21_X1 U6574 ( .B1(n5847), .B2(n5846), .A(n5845), .ZN(n5848) );
  XOR2_X1 U6575 ( .A(n5849), .B(n5848), .Z(n6210) );
  NAND2_X1 U6576 ( .A1(n5850), .A2(n6978), .ZN(n5860) );
  NAND3_X1 U6577 ( .A1(n5852), .A2(EBX_REG_31__SCAN_IN), .A3(n5851), .ZN(n5853) );
  OAI21_X1 U6578 ( .B1(n6981), .B2(n5854), .A(n5853), .ZN(n5857) );
  NOR4_X1 U6579 ( .A1(n5862), .A2(REIP_REG_31__SCAN_IN), .A3(n5855), .A4(n6655), .ZN(n5856) );
  AOI211_X1 U6580 ( .C1(REIP_REG_31__SCAN_IN), .C2(n5858), .A(n5857), .B(n5856), .ZN(n5859) );
  OAI211_X1 U6581 ( .C1(n6210), .C2(n6975), .A(n5860), .B(n5859), .ZN(U2796)
         );
  INV_X1 U6582 ( .A(n5861), .ZN(n6228) );
  NOR2_X1 U6583 ( .A1(n5862), .A2(REIP_REG_29__SCAN_IN), .ZN(n5867) );
  AOI22_X1 U6584 ( .A1(n6972), .A2(EBX_REG_29__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6955), .ZN(n5865) );
  OR2_X1 U6585 ( .A1(n6973), .A2(n5863), .ZN(n5864) );
  OAI211_X1 U6586 ( .C1(n5875), .C2(n6655), .A(n5865), .B(n5864), .ZN(n5866)
         );
  AOI211_X1 U6587 ( .C1(n6228), .C2(n6930), .A(n5867), .B(n5866), .ZN(n5868)
         );
  OAI21_X1 U6588 ( .B1(n6051), .B2(n6961), .A(n5868), .ZN(U2798) );
  AND2_X1 U6589 ( .A1(n5887), .A2(n5869), .ZN(n5871) );
  OR2_X1 U6590 ( .A1(n5871), .A2(n5870), .ZN(n6231) );
  INV_X1 U6591 ( .A(n6054), .ZN(n6085) );
  NAND2_X1 U6592 ( .A1(n6085), .A2(n6978), .ZN(n5880) );
  INV_X1 U6593 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6008) );
  OAI22_X1 U6594 ( .A1(n6933), .A2(n6008), .B1(n5874), .B2(n6981), .ZN(n5878)
         );
  NAND2_X1 U6595 ( .A1(n6651), .A2(REIP_REG_27__SCAN_IN), .ZN(n5876) );
  OAI22_X1 U6596 ( .A1(n5891), .A2(n5876), .B1(n6651), .B2(n5875), .ZN(n5877)
         );
  AOI211_X1 U6597 ( .C1(n6081), .C2(n6950), .A(n5878), .B(n5877), .ZN(n5879)
         );
  OAI211_X1 U6598 ( .C1(n6975), .C2(n6231), .A(n5880), .B(n5879), .ZN(U2799)
         );
  INV_X1 U6599 ( .A(n5881), .ZN(n5884) );
  INV_X1 U6600 ( .A(n5882), .ZN(n5883) );
  INV_X1 U6601 ( .A(n6094), .ZN(n6057) );
  NAND2_X1 U6602 ( .A1(n3453), .A2(n5885), .ZN(n5886) );
  AND2_X1 U6603 ( .A1(n5887), .A2(n5886), .ZN(n6244) );
  INV_X1 U6604 ( .A(n5888), .ZN(n6092) );
  INV_X1 U6605 ( .A(n5964), .ZN(n5890) );
  NOR2_X1 U6606 ( .A1(n5890), .A2(n5889), .ZN(n5904) );
  NOR2_X1 U6607 ( .A1(n5891), .A2(REIP_REG_27__SCAN_IN), .ZN(n5892) );
  AOI21_X1 U6608 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5904), .A(n5892), .ZN(n5894) );
  AOI22_X1 U6609 ( .A1(n6972), .A2(EBX_REG_27__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6955), .ZN(n5893) );
  OAI211_X1 U6610 ( .C1(n6092), .C2(n6973), .A(n5894), .B(n5893), .ZN(n5895)
         );
  AOI21_X1 U6611 ( .B1(n6244), .B2(n6930), .A(n5895), .ZN(n5896) );
  OAI21_X1 U6612 ( .B1(n6057), .B2(n6961), .A(n5896), .ZN(U2800) );
  AOI21_X1 U6613 ( .B1(n5899), .B2(n5898), .A(n5882), .ZN(n6101) );
  INV_X1 U6614 ( .A(n6101), .ZN(n6060) );
  OR2_X1 U6615 ( .A1(n5900), .A2(n5901), .ZN(n5902) );
  AND2_X1 U6616 ( .A1(n5902), .A2(n3453), .ZN(n6255) );
  INV_X1 U6617 ( .A(n5903), .ZN(n5916) );
  INV_X1 U6618 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6504) );
  NOR2_X1 U6619 ( .A1(n5916), .A2(n6504), .ZN(n5905) );
  OAI21_X1 U6620 ( .B1(n5905), .B2(REIP_REG_26__SCAN_IN), .A(n5904), .ZN(n5907) );
  AOI22_X1 U6621 ( .A1(n6972), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6955), .ZN(n5906) );
  OAI211_X1 U6622 ( .C1(n6973), .C2(n6099), .A(n5907), .B(n5906), .ZN(n5908)
         );
  AOI21_X1 U6623 ( .B1(n6255), .B2(n6930), .A(n5908), .ZN(n5909) );
  OAI21_X1 U6624 ( .B1(n6060), .B2(n6961), .A(n5909), .ZN(U2801) );
  OAI21_X1 U6625 ( .B1(n5910), .B2(n5911), .A(n5898), .ZN(n6106) );
  INV_X1 U6626 ( .A(n5933), .ZN(n5912) );
  NAND2_X1 U6627 ( .A1(n5939), .A2(n5912), .ZN(n5913) );
  AOI21_X1 U6628 ( .B1(n5914), .B2(n5913), .A(n5900), .ZN(n6260) );
  AOI22_X1 U6629 ( .A1(n6972), .A2(EBX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6955), .ZN(n5915) );
  OAI21_X1 U6630 ( .B1(n5916), .B2(REIP_REG_25__SCAN_IN), .A(n5915), .ZN(n5921) );
  INV_X1 U6631 ( .A(n5917), .ZN(n6108) );
  NAND3_X1 U6632 ( .A1(n5964), .A2(REIP_REG_25__SCAN_IN), .A3(n5918), .ZN(
        n5919) );
  OAI21_X1 U6633 ( .B1(n6973), .B2(n6108), .A(n5919), .ZN(n5920) );
  AOI211_X1 U6634 ( .C1(n6260), .C2(n6930), .A(n5921), .B(n5920), .ZN(n5922)
         );
  OAI21_X1 U6635 ( .B1(n6106), .B2(n6961), .A(n5922), .ZN(U2802) );
  NOR2_X1 U6636 ( .A1(n5923), .A2(n5924), .ZN(n5925) );
  AND2_X1 U6637 ( .A1(n5964), .A2(n5926), .ZN(n5942) );
  NOR2_X1 U6638 ( .A1(n6973), .A2(n6122), .ZN(n5932) );
  NAND2_X1 U6639 ( .A1(n6643), .A2(n5927), .ZN(n5930) );
  NAND2_X1 U6640 ( .A1(n6972), .A2(EBX_REG_24__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U6641 ( .A1(n6955), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5928)
         );
  OAI211_X1 U6642 ( .C1(n6905), .C2(n5930), .A(n5929), .B(n5928), .ZN(n5931)
         );
  AOI211_X1 U6643 ( .C1(n5942), .C2(REIP_REG_24__SCAN_IN), .A(n5932), .B(n5931), .ZN(n5935) );
  XNOR2_X1 U6644 ( .A(n5939), .B(n5933), .ZN(n6272) );
  NAND2_X1 U6645 ( .A1(n6272), .A2(n6930), .ZN(n5934) );
  OAI211_X1 U6646 ( .C1(n6120), .C2(n6961), .A(n5935), .B(n5934), .ZN(U2803)
         );
  AOI21_X1 U6647 ( .B1(n5937), .B2(n5936), .A(n5923), .ZN(n6135) );
  INV_X1 U6648 ( .A(n6135), .ZN(n6067) );
  AND2_X1 U6649 ( .A1(n3459), .A2(n5938), .ZN(n5940) );
  OR2_X1 U6650 ( .A1(n5940), .A2(n5939), .ZN(n6279) );
  INV_X1 U6651 ( .A(n6279), .ZN(n5949) );
  INV_X1 U6652 ( .A(n6131), .ZN(n5947) );
  NOR2_X1 U6653 ( .A1(n6905), .A2(n5941), .ZN(n5943) );
  OAI21_X1 U6654 ( .B1(REIP_REG_23__SCAN_IN), .B2(n5943), .A(n5942), .ZN(n5946) );
  NOR2_X1 U6655 ( .A1(n6133), .A2(n6981), .ZN(n5944) );
  AOI21_X1 U6656 ( .B1(n6972), .B2(EBX_REG_23__SCAN_IN), .A(n5944), .ZN(n5945)
         );
  OAI211_X1 U6657 ( .C1(n6973), .C2(n5947), .A(n5946), .B(n5945), .ZN(n5948)
         );
  AOI21_X1 U6658 ( .B1(n5949), .B2(n6930), .A(n5948), .ZN(n5950) );
  OAI21_X1 U6659 ( .B1(n6067), .B2(n6961), .A(n5950), .ZN(U2804) );
  INV_X1 U6660 ( .A(n5936), .ZN(n5952) );
  AOI21_X1 U6661 ( .B1(n5953), .B2(n5951), .A(n5952), .ZN(n6143) );
  NAND2_X1 U6662 ( .A1(n5975), .A2(n5954), .ZN(n5955) );
  NAND2_X1 U6663 ( .A1(n3459), .A2(n5955), .ZN(n6286) );
  INV_X1 U6664 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U6665 ( .A1(n6401), .A2(n5956), .ZN(n5959) );
  NAND2_X1 U6666 ( .A1(n6972), .A2(EBX_REG_22__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U6667 ( .A1(n6955), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5957)
         );
  OAI211_X1 U6668 ( .C1(n6905), .C2(n5959), .A(n5958), .B(n5957), .ZN(n5961)
         );
  NOR2_X1 U6669 ( .A1(n6973), .A2(n6141), .ZN(n5960) );
  NOR2_X1 U6670 ( .A1(n5961), .A2(n5960), .ZN(n5968) );
  INV_X1 U6671 ( .A(n5962), .ZN(n5965) );
  NAND2_X1 U6672 ( .A1(n6875), .A2(n5965), .ZN(n5963) );
  AND2_X1 U6673 ( .A1(n5964), .A2(n5963), .ZN(n6971) );
  NAND2_X1 U6674 ( .A1(n6638), .A2(n5965), .ZN(n5966) );
  NOR2_X1 U6675 ( .A1(n6905), .A2(n5966), .ZN(n5977) );
  OAI21_X1 U6676 ( .B1(n6971), .B2(n5977), .A(REIP_REG_22__SCAN_IN), .ZN(n5967) );
  OAI211_X1 U6677 ( .C1(n6286), .C2(n6975), .A(n5968), .B(n5967), .ZN(n5969)
         );
  AOI21_X1 U6678 ( .B1(n6143), .B2(n6978), .A(n5969), .ZN(n5970) );
  INV_X1 U6679 ( .A(n5970), .ZN(U2805) );
  OAI21_X1 U6680 ( .B1(n5971), .B2(n5972), .A(n5951), .ZN(n6150) );
  INV_X1 U6681 ( .A(n6153), .ZN(n5980) );
  NAND2_X1 U6682 ( .A1(n6024), .A2(n5973), .ZN(n5974) );
  NAND2_X1 U6683 ( .A1(n5975), .A2(n5974), .ZN(n6297) );
  INV_X1 U6684 ( .A(n6297), .ZN(n5978) );
  INV_X1 U6685 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6149) );
  INV_X1 U6686 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6016) );
  OAI22_X1 U6687 ( .A1(n6149), .A2(n6981), .B1(n6016), .B2(n6933), .ZN(n5976)
         );
  AOI211_X1 U6688 ( .C1(n5978), .C2(n6930), .A(n5977), .B(n5976), .ZN(n5979)
         );
  OAI21_X1 U6689 ( .B1(n5980), .B2(n6973), .A(n5979), .ZN(n5981) );
  AOI21_X1 U6690 ( .B1(REIP_REG_21__SCAN_IN), .B2(n6971), .A(n5981), .ZN(n5982) );
  OAI21_X1 U6691 ( .B1(n6150), .B2(n6961), .A(n5982), .ZN(U2806) );
  AND2_X1 U6692 ( .A1(n5983), .A2(n5984), .ZN(n5986) );
  OR2_X1 U6693 ( .A1(n5986), .A2(n5985), .ZN(n6165) );
  NOR2_X1 U6694 ( .A1(n6034), .A2(n5987), .ZN(n5988) );
  OR2_X1 U6695 ( .A1(n6022), .A2(n5988), .ZN(n6516) );
  AOI21_X1 U6696 ( .B1(n6955), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6954), 
        .ZN(n5989) );
  OAI21_X1 U6697 ( .B1(n6975), .B2(n6516), .A(n5989), .ZN(n5996) );
  NAND2_X1 U6698 ( .A1(n5990), .A2(n5991), .ZN(n6968) );
  NAND2_X1 U6699 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n6969) );
  OAI21_X1 U6700 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n6969), .ZN(n5994) );
  OR2_X1 U6701 ( .A1(n6905), .A2(n5991), .ZN(n5992) );
  AND2_X1 U6702 ( .A1(n5992), .A2(n6875), .ZN(n6957) );
  INV_X1 U6703 ( .A(n6957), .ZN(n5999) );
  AOI22_X1 U6704 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6972), .B1(
        REIP_REG_19__SCAN_IN), .B2(n5999), .ZN(n5993) );
  OAI21_X1 U6705 ( .B1(n6968), .B2(n5994), .A(n5993), .ZN(n5995) );
  AOI211_X1 U6706 ( .C1(n6950), .C2(n6168), .A(n5996), .B(n5995), .ZN(n5997)
         );
  OAI21_X1 U6707 ( .B1(n6165), .B2(n6961), .A(n5997), .ZN(U2808) );
  OAI21_X1 U6708 ( .B1(n6944), .B2(n5998), .A(n6633), .ZN(n6000) );
  AOI22_X1 U6709 ( .A1(n6000), .A2(n5999), .B1(PHYADDRPOINTER_REG_17__SCAN_IN), 
        .B2(n6955), .ZN(n6006) );
  INV_X1 U6710 ( .A(n6182), .ZN(n6003) );
  AOI21_X1 U6711 ( .B1(n6972), .B2(EBX_REG_17__SCAN_IN), .A(n6954), .ZN(n6002)
         );
  NAND2_X1 U6712 ( .A1(n6930), .A2(n6845), .ZN(n6001) );
  OAI211_X1 U6713 ( .C1(n6003), .C2(n6973), .A(n6002), .B(n6001), .ZN(n6004)
         );
  INV_X1 U6714 ( .A(n6004), .ZN(n6005) );
  OAI211_X1 U6715 ( .C1(n6185), .C2(n6961), .A(n6006), .B(n6005), .ZN(U2810)
         );
  OAI22_X1 U6716 ( .A1(n6210), .A2(n6045), .B1(n6047), .B2(n6007), .ZN(U2828)
         );
  OAI222_X1 U6717 ( .A1(n6008), .A2(n6047), .B1(n6045), .B2(n6231), .C1(n6054), 
        .C2(n6039), .ZN(U2831) );
  AOI22_X1 U6718 ( .A1(n6244), .A2(n6037), .B1(n6012), .B2(EBX_REG_27__SCAN_IN), .ZN(n6009) );
  OAI21_X1 U6719 ( .B1(n6057), .B2(n6039), .A(n6009), .ZN(U2832) );
  AOI22_X1 U6720 ( .A1(n6255), .A2(n6037), .B1(n6012), .B2(EBX_REG_26__SCAN_IN), .ZN(n6010) );
  OAI21_X1 U6721 ( .B1(n6060), .B2(n6039), .A(n6010), .ZN(U2833) );
  AOI22_X1 U6722 ( .A1(n6260), .A2(n6037), .B1(n6012), .B2(EBX_REG_25__SCAN_IN), .ZN(n6011) );
  OAI21_X1 U6723 ( .B1(n6106), .B2(n6039), .A(n6011), .ZN(U2834) );
  AOI22_X1 U6724 ( .A1(n6272), .A2(n6037), .B1(EBX_REG_24__SCAN_IN), .B2(n6012), .ZN(n6013) );
  OAI21_X1 U6725 ( .B1(n6120), .B2(n6039), .A(n6013), .ZN(U2835) );
  INV_X1 U6726 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6014) );
  OAI222_X1 U6727 ( .A1(n6014), .A2(n6047), .B1(n6045), .B2(n6279), .C1(n6067), 
        .C2(n6039), .ZN(U2836) );
  INV_X1 U6728 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6015) );
  INV_X1 U6729 ( .A(n6143), .ZN(n6070) );
  OAI222_X1 U6730 ( .A1(n6015), .A2(n6047), .B1(n6045), .B2(n6286), .C1(n6070), 
        .C2(n6039), .ZN(U2837) );
  OAI22_X1 U6731 ( .A1(n6297), .A2(n6045), .B1(n6016), .B2(n6047), .ZN(n6017)
         );
  INV_X1 U6732 ( .A(n6017), .ZN(n6018) );
  OAI21_X1 U6733 ( .B1(n6150), .B2(n6039), .A(n6018), .ZN(U2838) );
  NOR2_X1 U6734 ( .A1(n5985), .A2(n6019), .ZN(n6020) );
  OR2_X1 U6735 ( .A1(n5971), .A2(n6020), .ZN(n6157) );
  INV_X1 U6736 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6025) );
  OR2_X1 U6737 ( .A1(n6022), .A2(n6021), .ZN(n6023) );
  NAND2_X1 U6738 ( .A1(n6024), .A2(n6023), .ZN(n6976) );
  OAI222_X1 U6739 ( .A1(n6039), .A2(n6157), .B1(n6047), .B2(n6025), .C1(n6976), 
        .C2(n6045), .ZN(U2839) );
  OAI22_X1 U6740 ( .A1(n6516), .A2(n6045), .B1(n6026), .B2(n6047), .ZN(n6027)
         );
  INV_X1 U6741 ( .A(n6027), .ZN(n6028) );
  OAI21_X1 U6742 ( .B1(n6165), .B2(n6039), .A(n6028), .ZN(U2840) );
  INV_X1 U6743 ( .A(n5983), .ZN(n6029) );
  AOI21_X1 U6744 ( .B1(n6030), .B2(n5776), .A(n6029), .ZN(n7090) );
  INV_X1 U6745 ( .A(n7090), .ZN(n6962) );
  AND2_X1 U6746 ( .A1(n6032), .A2(n6031), .ZN(n6033) );
  NOR2_X1 U6747 ( .A1(n6034), .A2(n6033), .ZN(n6959) );
  NOR2_X1 U6748 ( .A1(n6047), .A2(n6035), .ZN(n6036) );
  AOI21_X1 U6749 ( .B1(n6959), .B2(n6037), .A(n6036), .ZN(n6038) );
  OAI21_X1 U6750 ( .B1(n6962), .B2(n6039), .A(n6038), .ZN(U2841) );
  AOI21_X1 U6751 ( .B1(n6040), .B2(n5731), .A(n5775), .ZN(n7087) );
  INV_X1 U6752 ( .A(n7087), .ZN(n6048) );
  INV_X1 U6753 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6046) );
  OR2_X1 U6754 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  NAND2_X1 U6755 ( .A1(n6044), .A2(n6043), .ZN(n6953) );
  OAI222_X1 U6756 ( .A1(n6048), .A2(n6039), .B1(n6047), .B2(n6046), .C1(n6953), 
        .C2(n6045), .ZN(U2843) );
  AOI22_X1 U6757 ( .A1(n7093), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n7096), .ZN(n6050) );
  NAND2_X1 U6758 ( .A1(n7097), .A2(DATAI_13_), .ZN(n6049) );
  OAI211_X1 U6759 ( .C1(n6051), .C2(n7086), .A(n6050), .B(n6049), .ZN(U2862)
         );
  AOI22_X1 U6760 ( .A1(n7093), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n7096), .ZN(n6053) );
  NAND2_X1 U6761 ( .A1(n7097), .A2(DATAI_12_), .ZN(n6052) );
  OAI211_X1 U6762 ( .C1(n6054), .C2(n7086), .A(n6053), .B(n6052), .ZN(U2863)
         );
  AOI22_X1 U6763 ( .A1(n7093), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n7096), .ZN(n6056) );
  NAND2_X1 U6764 ( .A1(n7097), .A2(DATAI_11_), .ZN(n6055) );
  OAI211_X1 U6765 ( .C1(n6057), .C2(n7086), .A(n6056), .B(n6055), .ZN(U2864)
         );
  AOI22_X1 U6766 ( .A1(n7093), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n7096), .ZN(n6059) );
  NAND2_X1 U6767 ( .A1(n7097), .A2(DATAI_10_), .ZN(n6058) );
  OAI211_X1 U6768 ( .C1(n6060), .C2(n7086), .A(n6059), .B(n6058), .ZN(U2865)
         );
  AOI22_X1 U6769 ( .A1(n7093), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n7096), .ZN(n6062) );
  NAND2_X1 U6770 ( .A1(n7097), .A2(DATAI_9_), .ZN(n6061) );
  OAI211_X1 U6771 ( .C1(n6106), .C2(n7086), .A(n6062), .B(n6061), .ZN(U2866)
         );
  AOI22_X1 U6772 ( .A1(n7093), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n7096), .ZN(n6064) );
  NAND2_X1 U6773 ( .A1(n7097), .A2(DATAI_8_), .ZN(n6063) );
  OAI211_X1 U6774 ( .C1(n6120), .C2(n7086), .A(n6064), .B(n6063), .ZN(U2867)
         );
  AOI22_X1 U6775 ( .A1(n7093), .A2(DATAI_23_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n7096), .ZN(n6066) );
  NAND2_X1 U6776 ( .A1(n7097), .A2(DATAI_7_), .ZN(n6065) );
  OAI211_X1 U6777 ( .C1(n6067), .C2(n7086), .A(n6066), .B(n6065), .ZN(U2868)
         );
  AOI22_X1 U6778 ( .A1(n7093), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n7096), .ZN(n6069) );
  NAND2_X1 U6779 ( .A1(n7097), .A2(DATAI_6_), .ZN(n6068) );
  OAI211_X1 U6780 ( .C1(n6070), .C2(n7086), .A(n6069), .B(n6068), .ZN(U2869)
         );
  AOI22_X1 U6781 ( .A1(n7093), .A2(DATAI_21_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n7096), .ZN(n6072) );
  NAND2_X1 U6782 ( .A1(n7097), .A2(DATAI_5_), .ZN(n6071) );
  OAI211_X1 U6783 ( .C1(n6150), .C2(n7086), .A(n6072), .B(n6071), .ZN(U2870)
         );
  AOI22_X1 U6784 ( .A1(n7093), .A2(DATAI_19_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n7096), .ZN(n6074) );
  NAND2_X1 U6785 ( .A1(n7097), .A2(DATAI_3_), .ZN(n6073) );
  OAI211_X1 U6786 ( .C1(n6165), .C2(n7086), .A(n6074), .B(n6073), .ZN(U2872)
         );
  AOI22_X1 U6787 ( .A1(n7093), .A2(DATAI_17_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n7096), .ZN(n6076) );
  NAND2_X1 U6788 ( .A1(n7097), .A2(DATAI_1_), .ZN(n6075) );
  OAI211_X1 U6789 ( .C1(n6185), .C2(n7086), .A(n6076), .B(n6075), .ZN(U2874)
         );
  NAND2_X1 U6790 ( .A1(n6078), .A2(n6077), .ZN(n6080) );
  XNOR2_X1 U6791 ( .A(n6137), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n6079)
         );
  XNOR2_X1 U6792 ( .A(n6080), .B(n6079), .ZN(n6241) );
  INV_X1 U6793 ( .A(n6081), .ZN(n6083) );
  AND2_X1 U6794 ( .A1(n6843), .A2(REIP_REG_28__SCAN_IN), .ZN(n6235) );
  AOI21_X1 U6795 ( .B1(n6691), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n6235), 
        .ZN(n6082) );
  OAI21_X1 U6796 ( .B1(n6083), .B2(n6707), .A(n6082), .ZN(n6084) );
  AOI21_X1 U6797 ( .B1(n6085), .B2(n6710), .A(n6084), .ZN(n6086) );
  OAI21_X1 U6798 ( .B1(n6241), .B2(n6993), .A(n6086), .ZN(U2958) );
  NAND2_X1 U6799 ( .A1(n4603), .A2(n6252), .ZN(n6088) );
  MUX2_X1 U6800 ( .A(n6089), .B(n6088), .S(n6087), .Z(n6090) );
  XNOR2_X1 U6801 ( .A(n6090), .B(n6233), .ZN(n6248) );
  AND2_X1 U6802 ( .A1(n6843), .A2(REIP_REG_27__SCAN_IN), .ZN(n6242) );
  AOI21_X1 U6803 ( .B1(n6691), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n6242), 
        .ZN(n6091) );
  OAI21_X1 U6804 ( .B1(n6707), .B2(n6092), .A(n6091), .ZN(n6093) );
  AOI21_X1 U6805 ( .B1(n6094), .B2(n6710), .A(n6093), .ZN(n6095) );
  OAI21_X1 U6806 ( .B1(n6248), .B2(n6993), .A(n6095), .ZN(U2959) );
  XNOR2_X1 U6807 ( .A(n6137), .B(n6252), .ZN(n6096) );
  XNOR2_X1 U6808 ( .A(n6097), .B(n6096), .ZN(n6258) );
  AND2_X1 U6809 ( .A1(n6843), .A2(REIP_REG_26__SCAN_IN), .ZN(n6254) );
  AOI21_X1 U6810 ( .B1(n6691), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6254), 
        .ZN(n6098) );
  OAI21_X1 U6811 ( .B1(n6707), .B2(n6099), .A(n6098), .ZN(n6100) );
  AOI21_X1 U6812 ( .B1(n6101), .B2(n6710), .A(n6100), .ZN(n6102) );
  OAI21_X1 U6813 ( .B1(n6993), .B2(n6258), .A(n6102), .ZN(U2960) );
  AOI21_X1 U6814 ( .B1(n6105), .B2(n6103), .A(n6104), .ZN(n6265) );
  INV_X1 U6815 ( .A(n6106), .ZN(n6110) );
  AND2_X1 U6816 ( .A1(n6843), .A2(REIP_REG_25__SCAN_IN), .ZN(n6259) );
  AOI21_X1 U6817 ( .B1(n6691), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n6259), 
        .ZN(n6107) );
  OAI21_X1 U6818 ( .B1(n6707), .B2(n6108), .A(n6107), .ZN(n6109) );
  AOI21_X1 U6819 ( .B1(n6110), .B2(n6710), .A(n6109), .ZN(n6111) );
  OAI21_X1 U6820 ( .B1(n6265), .B2(n6993), .A(n6111), .ZN(U2961) );
  INV_X1 U6821 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6113) );
  XNOR2_X1 U6822 ( .A(n6137), .B(n6113), .ZN(n6163) );
  OR2_X2 U6823 ( .A1(n6112), .A2(n6163), .ZN(n6161) );
  INV_X1 U6824 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6114) );
  NOR2_X1 U6825 ( .A1(n6187), .A2(n6114), .ZN(n6115) );
  NAND3_X1 U6826 ( .A1(n6146), .A2(n6089), .A3(n6116), .ZN(n6128) );
  XNOR2_X1 U6827 ( .A(n6137), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6147)
         );
  NOR2_X1 U6828 ( .A1(n6089), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6117)
         );
  NOR2_X1 U6829 ( .A1(n6089), .A2(n6308), .ZN(n6145) );
  NAND4_X1 U6830 ( .A1(n6139), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n6187), .ZN(n6118) );
  OAI21_X1 U6831 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n6128), .A(n6118), 
        .ZN(n6119) );
  XNOR2_X1 U6832 ( .A(n6119), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6274)
         );
  INV_X1 U6833 ( .A(n6120), .ZN(n6124) );
  NOR2_X1 U6834 ( .A1(n6801), .A2(n6643), .ZN(n6271) );
  AOI21_X1 U6835 ( .B1(n6691), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n6271), 
        .ZN(n6121) );
  OAI21_X1 U6836 ( .B1(n6707), .B2(n6122), .A(n6121), .ZN(n6123) );
  AOI21_X1 U6837 ( .B1(n6124), .B2(n6710), .A(n6123), .ZN(n6125) );
  OAI21_X1 U6838 ( .B1(n6274), .B2(n6993), .A(n6125), .ZN(U2962) );
  INV_X1 U6839 ( .A(n6127), .ZN(n6276) );
  NAND2_X1 U6840 ( .A1(n6171), .A2(n6276), .ZN(n6129) );
  OAI21_X1 U6841 ( .B1(n6126), .B2(n6129), .A(n6128), .ZN(n6130) );
  XNOR2_X1 U6842 ( .A(n6130), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6283)
         );
  NAND2_X1 U6843 ( .A1(n6709), .A2(n6131), .ZN(n6132) );
  NAND2_X1 U6844 ( .A1(n6843), .A2(REIP_REG_23__SCAN_IN), .ZN(n6278) );
  OAI211_X1 U6845 ( .C1(n6205), .C2(n6133), .A(n6132), .B(n6278), .ZN(n6134)
         );
  AOI21_X1 U6846 ( .B1(n6135), .B2(n6710), .A(n6134), .ZN(n6136) );
  OAI21_X1 U6847 ( .B1(n6283), .B2(n6993), .A(n6136), .ZN(U2963) );
  XNOR2_X1 U6848 ( .A(n6137), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6138)
         );
  XNOR2_X1 U6849 ( .A(n6139), .B(n6138), .ZN(n6293) );
  NAND2_X1 U6850 ( .A1(n6843), .A2(REIP_REG_22__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U6851 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6140)
         );
  OAI211_X1 U6852 ( .C1(n6707), .C2(n6141), .A(n6285), .B(n6140), .ZN(n6142)
         );
  AOI21_X1 U6853 ( .B1(n6143), .B2(n6710), .A(n6142), .ZN(n6144) );
  OAI21_X1 U6854 ( .B1(n6293), .B2(n6993), .A(n6144), .ZN(U2964) );
  NOR2_X1 U6855 ( .A1(n6146), .A2(n6145), .ZN(n6148) );
  XNOR2_X1 U6856 ( .A(n6148), .B(n6147), .ZN(n6301) );
  NAND2_X1 U6857 ( .A1(n6843), .A2(REIP_REG_21__SCAN_IN), .ZN(n6296) );
  OAI21_X1 U6858 ( .B1(n6205), .B2(n6149), .A(n6296), .ZN(n6152) );
  NOR2_X1 U6859 ( .A1(n6150), .A2(n6685), .ZN(n6151) );
  AOI211_X1 U6860 ( .C1(n6709), .C2(n6153), .A(n6152), .B(n6151), .ZN(n6154)
         );
  OAI21_X1 U6861 ( .B1(n6301), .B2(n6993), .A(n6154), .ZN(U2965) );
  NAND2_X1 U6862 ( .A1(n6161), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6155) );
  MUX2_X1 U6863 ( .A(n6161), .B(n6155), .S(n6171), .Z(n6156) );
  XOR2_X1 U6864 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .B(n6156), .Z(n6312) );
  NAND2_X1 U6865 ( .A1(n6843), .A2(REIP_REG_20__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U6866 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6158)
         );
  OAI211_X1 U6867 ( .C1(n6707), .C2(n6974), .A(n6303), .B(n6158), .ZN(n6159)
         );
  AOI21_X1 U6868 ( .B1(n7095), .B2(n6710), .A(n6159), .ZN(n6160) );
  OAI21_X1 U6869 ( .B1(n6312), .B2(n6993), .A(n6160), .ZN(U2966) );
  INV_X1 U6870 ( .A(n6161), .ZN(n6162) );
  AOI21_X1 U6871 ( .B1(n6112), .B2(n6163), .A(n6162), .ZN(n6522) );
  NAND2_X1 U6872 ( .A1(n6843), .A2(REIP_REG_19__SCAN_IN), .ZN(n6515) );
  OAI21_X1 U6873 ( .B1(n6205), .B2(n6164), .A(n6515), .ZN(n6167) );
  NOR2_X1 U6874 ( .A1(n6165), .A2(n6685), .ZN(n6166) );
  AOI211_X1 U6875 ( .C1(n6709), .C2(n6168), .A(n6167), .B(n6166), .ZN(n6169)
         );
  OAI21_X1 U6876 ( .B1(n6522), .B2(n6993), .A(n6169), .ZN(U2967) );
  OAI21_X1 U6877 ( .B1(n6171), .B2(n6841), .A(n6170), .ZN(n6179) );
  NAND2_X1 U6878 ( .A1(n4603), .A2(n6532), .ZN(n6173) );
  NAND2_X1 U6879 ( .A1(n6187), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6172) );
  OAI22_X1 U6880 ( .A1(n6179), .A2(n6173), .B1(n6170), .B2(n6172), .ZN(n6174)
         );
  XNOR2_X1 U6881 ( .A(n6174), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6541)
         );
  AND2_X1 U6882 ( .A1(n6843), .A2(REIP_REG_18__SCAN_IN), .ZN(n6536) );
  AOI21_X1 U6883 ( .B1(n6691), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6536), 
        .ZN(n6175) );
  OAI21_X1 U6884 ( .B1(n6707), .B2(n6966), .A(n6175), .ZN(n6176) );
  AOI21_X1 U6885 ( .B1(n7090), .B2(n6710), .A(n6176), .ZN(n6177) );
  OAI21_X1 U6886 ( .B1(n6541), .B2(n6993), .A(n6177), .ZN(U2968) );
  XNOR2_X1 U6887 ( .A(n6187), .B(n6532), .ZN(n6178) );
  XNOR2_X1 U6888 ( .A(n6179), .B(n6178), .ZN(n6848) );
  NAND2_X1 U6889 ( .A1(n6848), .A2(n6704), .ZN(n6184) );
  OAI22_X1 U6890 ( .A1(n6205), .A2(n6180), .B1(n6801), .B2(n6633), .ZN(n6181)
         );
  AOI21_X1 U6891 ( .B1(n6709), .B2(n6182), .A(n6181), .ZN(n6183) );
  OAI211_X1 U6892 ( .C1(n6685), .C2(n6185), .A(n6184), .B(n6183), .ZN(U2969)
         );
  XNOR2_X1 U6893 ( .A(n6187), .B(n6841), .ZN(n6188) );
  XNOR2_X1 U6894 ( .A(n6189), .B(n6188), .ZN(n6837) );
  AOI22_X1 U6895 ( .A1(n6691), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6843), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n6190) );
  OAI21_X1 U6896 ( .B1(n6707), .B2(n6191), .A(n6190), .ZN(n6192) );
  AOI21_X1 U6897 ( .B1(n7087), .B2(n6710), .A(n6192), .ZN(n6193) );
  OAI21_X1 U6898 ( .B1(n6837), .B2(n6993), .A(n6193), .ZN(U2970) );
  NAND2_X1 U6899 ( .A1(n6195), .A2(n6194), .ZN(n6197) );
  XOR2_X1 U6900 ( .A(n6197), .B(n6196), .Z(n6829) );
  NAND2_X1 U6901 ( .A1(n6829), .A2(n6704), .ZN(n6202) );
  INV_X1 U6902 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6198) );
  NOR2_X1 U6903 ( .A1(n6801), .A2(n6198), .ZN(n6827) );
  NOR2_X1 U6904 ( .A1(n6707), .A2(n6199), .ZN(n6200) );
  AOI211_X1 U6905 ( .C1(n6691), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6827), 
        .B(n6200), .ZN(n6201) );
  OAI211_X1 U6906 ( .C1(n6685), .C2(n6203), .A(n6202), .B(n6201), .ZN(U2971)
         );
  OAI21_X1 U6907 ( .B1(n6205), .B2(n4128), .A(n6204), .ZN(n6207) );
  NOR2_X1 U6908 ( .A1(n6937), .A2(n6685), .ZN(n6206) );
  AOI211_X1 U6909 ( .C1(n6709), .C2(n6938), .A(n6207), .B(n6206), .ZN(n6208)
         );
  OAI21_X1 U6910 ( .B1(n6993), .B2(n6209), .A(n6208), .ZN(U2972) );
  INV_X1 U6911 ( .A(n6210), .ZN(n6219) );
  AOI21_X1 U6912 ( .B1(n6212), .B2(n6825), .A(n6211), .ZN(n6217) );
  NAND4_X1 U6913 ( .A1(n6232), .A2(n6213), .A3(INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n6216), .ZN(n6214) );
  OAI211_X1 U6914 ( .C1(n6217), .C2(n6216), .A(n6215), .B(n6214), .ZN(n6218)
         );
  AOI21_X1 U6915 ( .B1(n6219), .B2(n6846), .A(n6218), .ZN(n6220) );
  OAI21_X1 U6916 ( .B1(n6221), .B2(n6756), .A(n6220), .ZN(U2987) );
  INV_X1 U6917 ( .A(n6222), .ZN(n6227) );
  AOI21_X1 U6918 ( .B1(n6232), .B2(n6223), .A(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n6224) );
  NOR2_X1 U6919 ( .A1(n6225), .A2(n6224), .ZN(n6226) );
  AOI211_X1 U6920 ( .C1(n6228), .C2(n6846), .A(n6227), .B(n6226), .ZN(n6229)
         );
  OAI21_X1 U6921 ( .B1(n6230), .B2(n6756), .A(n6229), .ZN(U2989) );
  INV_X1 U6922 ( .A(n6231), .ZN(n6236) );
  INV_X1 U6923 ( .A(n6232), .ZN(n6238) );
  NOR3_X1 U6924 ( .A1(n6238), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n6233), 
        .ZN(n6234) );
  AOI211_X1 U6925 ( .C1(n6236), .C2(n6846), .A(n6235), .B(n6234), .ZN(n6240)
         );
  INV_X1 U6926 ( .A(n6237), .ZN(n6245) );
  NOR2_X1 U6927 ( .A1(n6238), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6243)
         );
  OAI21_X1 U6928 ( .B1(n6245), .B2(n6243), .A(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n6239) );
  OAI211_X1 U6929 ( .C1(n6241), .C2(n6756), .A(n6240), .B(n6239), .ZN(U2990)
         );
  AOI211_X1 U6930 ( .C1(n6244), .C2(n6846), .A(n6243), .B(n6242), .ZN(n6247)
         );
  NAND2_X1 U6931 ( .A1(n6245), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6246) );
  OAI211_X1 U6932 ( .C1(n6248), .C2(n6756), .A(n6247), .B(n6246), .ZN(U2991)
         );
  INV_X1 U6933 ( .A(n6249), .ZN(n6250) );
  AOI211_X1 U6934 ( .C1(n6252), .C2(n6251), .A(n6250), .B(n6262), .ZN(n6253)
         );
  AOI211_X1 U6935 ( .C1(n6255), .C2(n6846), .A(n6254), .B(n6253), .ZN(n6257)
         );
  NAND2_X1 U6936 ( .A1(n6266), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6256) );
  OAI211_X1 U6937 ( .C1(n6258), .C2(n6756), .A(n6257), .B(n6256), .ZN(U2992)
         );
  AOI21_X1 U6938 ( .B1(n6260), .B2(n6846), .A(n6259), .ZN(n6261) );
  OAI21_X1 U6939 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n6262), .A(n6261), 
        .ZN(n6263) );
  AOI21_X1 U6940 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n6266), .A(n6263), 
        .ZN(n6264) );
  OAI21_X1 U6941 ( .B1(n6265), .B2(n6756), .A(n6264), .ZN(U2993) );
  NAND3_X1 U6942 ( .A1(n6288), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n6276), .ZN(n6268) );
  INV_X1 U6943 ( .A(n6266), .ZN(n6267) );
  AOI21_X1 U6944 ( .B1(n6269), .B2(n6268), .A(n6267), .ZN(n6270) );
  AOI211_X1 U6945 ( .C1(n6846), .C2(n6272), .A(n6271), .B(n6270), .ZN(n6273)
         );
  OAI21_X1 U6946 ( .B1(n6274), .B2(n6756), .A(n6273), .ZN(U2994) );
  NAND3_X1 U6947 ( .A1(n6288), .A2(n6276), .A3(n6275), .ZN(n6277) );
  OAI211_X1 U6948 ( .C1(n6279), .C2(n6836), .A(n6278), .B(n6277), .ZN(n6280)
         );
  AOI21_X1 U6949 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n6281), .A(n6280), 
        .ZN(n6282) );
  OAI21_X1 U6950 ( .B1(n6283), .B2(n6756), .A(n6282), .ZN(U2995) );
  NAND4_X1 U6951 ( .A1(n6288), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n6308), .A4(n6289), .ZN(n6284) );
  OAI211_X1 U6952 ( .C1(n6286), .C2(n6836), .A(n6285), .B(n6284), .ZN(n6291)
         );
  INV_X1 U6953 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6287) );
  NAND3_X1 U6954 ( .A1(n6288), .A2(n6308), .A3(n6287), .ZN(n6295) );
  AOI21_X1 U6955 ( .B1(n6294), .B2(n6295), .A(n6289), .ZN(n6290) );
  NOR2_X1 U6956 ( .A1(n6291), .A2(n6290), .ZN(n6292) );
  OAI21_X1 U6957 ( .B1(n6293), .B2(n6756), .A(n6292), .ZN(U2996) );
  INV_X1 U6958 ( .A(n6294), .ZN(n6299) );
  OAI211_X1 U6959 ( .C1(n6297), .C2(n6836), .A(n6296), .B(n6295), .ZN(n6298)
         );
  AOI21_X1 U6960 ( .B1(n6299), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6298), 
        .ZN(n6300) );
  OAI21_X1 U6961 ( .B1(n6301), .B2(n6756), .A(n6300), .ZN(U2997) );
  INV_X1 U6962 ( .A(n6302), .ZN(n6520) );
  OAI21_X1 U6963 ( .B1(n6976), .B2(n6836), .A(n6303), .ZN(n6310) );
  NOR2_X1 U6964 ( .A1(n6304), .A2(n6824), .ZN(n6833) );
  NAND2_X1 U6965 ( .A1(n6833), .A2(n6305), .ZN(n6851) );
  INV_X1 U6966 ( .A(n6851), .ZN(n6538) );
  NAND2_X1 U6967 ( .A1(n6538), .A2(n6306), .ZN(n6517) );
  NOR3_X1 U6968 ( .A1(n6517), .A2(n6308), .A3(n6307), .ZN(n6309) );
  AOI211_X1 U6969 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n6520), .A(n6310), .B(n6309), .ZN(n6311) );
  OAI21_X1 U6970 ( .B1(n6312), .B2(n6756), .A(n6311), .ZN(U2998) );
  INV_X1 U6971 ( .A(keyinput_62), .ZN(n6405) );
  INV_X1 U6972 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6967) );
  INV_X1 U6973 ( .A(keyinput_61), .ZN(n6403) );
  OAI22_X1 U6974 ( .A1(n6643), .A2(keyinput_58), .B1(n6641), .B2(keyinput_59), 
        .ZN(n6313) );
  AOI221_X1 U6975 ( .B1(n6643), .B2(keyinput_58), .C1(keyinput_59), .C2(n6641), 
        .A(n6313), .ZN(n6399) );
  OAI22_X1 U6976 ( .A1(n6649), .A2(keyinput_55), .B1(keyinput_56), .B2(
        REIP_REG_26__SCAN_IN), .ZN(n6314) );
  AOI221_X1 U6977 ( .B1(n6649), .B2(keyinput_55), .C1(REIP_REG_26__SCAN_IN), 
        .C2(keyinput_56), .A(n6314), .ZN(n6396) );
  INV_X1 U6978 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6728) );
  AOI22_X1 U6979 ( .A1(n7024), .A2(keyinput_45), .B1(keyinput_46), .B2(n6728), 
        .ZN(n6315) );
  OAI221_X1 U6980 ( .B1(n7024), .B2(keyinput_45), .C1(n6728), .C2(keyinput_46), 
        .A(n6315), .ZN(n6384) );
  INV_X1 U6981 ( .A(keyinput_44), .ZN(n6382) );
  INV_X1 U6982 ( .A(MORE_REG_SCAN_IN), .ZN(n7025) );
  INV_X1 U6983 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6729) );
  OAI22_X1 U6984 ( .A1(n7126), .A2(keyinput_43), .B1(D_C_N_REG_SCAN_IN), .B2(
        keyinput_41), .ZN(n6316) );
  AOI221_X1 U6985 ( .B1(n7126), .B2(keyinput_43), .C1(keyinput_41), .C2(
        D_C_N_REG_SCAN_IN), .A(n6316), .ZN(n6379) );
  OAI22_X1 U6986 ( .A1(BS16_N), .A2(keyinput_34), .B1(NA_N), .B2(keyinput_33), 
        .ZN(n6317) );
  AOI221_X1 U6987 ( .B1(BS16_N), .B2(keyinput_34), .C1(keyinput_33), .C2(NA_N), 
        .A(n6317), .ZN(n6372) );
  INV_X1 U6988 ( .A(keyinput_32), .ZN(n6368) );
  OAI22_X1 U6989 ( .A1(n6417), .A2(keyinput_30), .B1(DATAI_2_), .B2(
        keyinput_29), .ZN(n6318) );
  AOI221_X1 U6990 ( .B1(n6417), .B2(keyinput_30), .C1(keyinput_29), .C2(
        DATAI_2_), .A(n6318), .ZN(n6365) );
  INV_X1 U6991 ( .A(keyinput_28), .ZN(n6363) );
  INV_X1 U6992 ( .A(keyinput_23), .ZN(n6356) );
  INV_X1 U6993 ( .A(keyinput_22), .ZN(n6354) );
  OAI22_X1 U6994 ( .A1(n6321), .A2(keyinput_20), .B1(n6320), .B2(keyinput_19), 
        .ZN(n6319) );
  AOI221_X1 U6995 ( .B1(n6321), .B2(keyinput_20), .C1(keyinput_19), .C2(n6320), 
        .A(n6319), .ZN(n6351) );
  INV_X1 U6996 ( .A(keyinput_18), .ZN(n6349) );
  INV_X1 U6997 ( .A(DATAI_16_), .ZN(n6323) );
  OAI22_X1 U6998 ( .A1(n6323), .A2(keyinput_15), .B1(DATAI_15_), .B2(
        keyinput_16), .ZN(n6322) );
  AOI221_X1 U6999 ( .B1(n6323), .B2(keyinput_15), .C1(keyinput_16), .C2(
        DATAI_15_), .A(n6322), .ZN(n6346) );
  INV_X1 U7000 ( .A(DATAI_17_), .ZN(n6444) );
  INV_X1 U7001 ( .A(keyinput_14), .ZN(n6344) );
  XNOR2_X1 U7002 ( .A(DATAI_27_), .B(keyinput_4), .ZN(n6335) );
  INV_X1 U7003 ( .A(DATAI_28_), .ZN(n6426) );
  INV_X1 U7004 ( .A(keyinput_3), .ZN(n6328) );
  INV_X1 U7005 ( .A(keyinput_0), .ZN(n6326) );
  OAI22_X1 U7006 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(DATAI_29_), .B2(
        keyinput_2), .ZN(n6324) );
  AOI221_X1 U7007 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(keyinput_2), .C2(
        DATAI_29_), .A(n6324), .ZN(n6325) );
  OAI221_X1 U7008 ( .B1(DATAI_31_), .B2(keyinput_0), .C1(n6424), .C2(n6326), 
        .A(n6325), .ZN(n6327) );
  OAI221_X1 U7009 ( .B1(DATAI_28_), .B2(keyinput_3), .C1(n6426), .C2(n6328), 
        .A(n6327), .ZN(n6334) );
  INV_X1 U7010 ( .A(DATAI_23_), .ZN(n6330) );
  AOI22_X1 U7011 ( .A1(keyinput_6), .A2(DATAI_25_), .B1(n6330), .B2(keyinput_8), .ZN(n6329) );
  OAI221_X1 U7012 ( .B1(keyinput_6), .B2(DATAI_25_), .C1(n6330), .C2(
        keyinput_8), .A(n6329), .ZN(n6333) );
  AOI22_X1 U7013 ( .A1(DATAI_24_), .A2(keyinput_7), .B1(DATAI_26_), .B2(
        keyinput_5), .ZN(n6331) );
  OAI221_X1 U7014 ( .B1(DATAI_24_), .B2(keyinput_7), .C1(DATAI_26_), .C2(
        keyinput_5), .A(n6331), .ZN(n6332) );
  AOI211_X1 U7015 ( .C1(n6335), .C2(n6334), .A(n6333), .B(n6332), .ZN(n6342)
         );
  XOR2_X1 U7016 ( .A(DATAI_22_), .B(keyinput_9), .Z(n6341) );
  INV_X1 U7017 ( .A(DATAI_21_), .ZN(n6337) );
  INV_X1 U7018 ( .A(DATAI_20_), .ZN(n6437) );
  OAI22_X1 U7019 ( .A1(n6337), .A2(keyinput_10), .B1(n6437), .B2(keyinput_11), 
        .ZN(n6336) );
  AOI221_X1 U7020 ( .B1(n6337), .B2(keyinput_10), .C1(keyinput_11), .C2(n6437), 
        .A(n6336), .ZN(n6340) );
  OAI22_X1 U7021 ( .A1(DATAI_19_), .A2(keyinput_12), .B1(DATAI_18_), .B2(
        keyinput_13), .ZN(n6338) );
  AOI221_X1 U7022 ( .B1(DATAI_19_), .B2(keyinput_12), .C1(keyinput_13), .C2(
        DATAI_18_), .A(n6338), .ZN(n6339) );
  OAI211_X1 U7023 ( .C1(n6342), .C2(n6341), .A(n6340), .B(n6339), .ZN(n6343)
         );
  OAI221_X1 U7024 ( .B1(DATAI_17_), .B2(keyinput_14), .C1(n6444), .C2(n6344), 
        .A(n6343), .ZN(n6345) );
  AOI22_X1 U7025 ( .A1(keyinput_17), .A2(n6449), .B1(n6346), .B2(n6345), .ZN(
        n6347) );
  OAI21_X1 U7026 ( .B1(n6449), .B2(keyinput_17), .A(n6347), .ZN(n6348) );
  OAI221_X1 U7027 ( .B1(DATAI_13_), .B2(keyinput_18), .C1(n6452), .C2(n6349), 
        .A(n6348), .ZN(n6350) );
  OAI211_X1 U7028 ( .C1(DATAI_10_), .C2(keyinput_21), .A(n6351), .B(n6350), 
        .ZN(n6352) );
  AOI21_X1 U7029 ( .B1(DATAI_10_), .B2(keyinput_21), .A(n6352), .ZN(n6353) );
  AOI221_X1 U7030 ( .B1(DATAI_9_), .B2(keyinput_22), .C1(n6457), .C2(n6354), 
        .A(n6353), .ZN(n6355) );
  AOI221_X1 U7031 ( .B1(DATAI_8_), .B2(n6356), .C1(n6460), .C2(keyinput_23), 
        .A(n6355), .ZN(n6361) );
  AOI22_X1 U7032 ( .A1(DATAI_6_), .A2(keyinput_25), .B1(DATAI_7_), .B2(
        keyinput_24), .ZN(n6357) );
  OAI221_X1 U7033 ( .B1(DATAI_6_), .B2(keyinput_25), .C1(DATAI_7_), .C2(
        keyinput_24), .A(n6357), .ZN(n6360) );
  OAI22_X1 U7034 ( .A1(DATAI_4_), .A2(keyinput_27), .B1(DATAI_5_), .B2(
        keyinput_26), .ZN(n6358) );
  AOI221_X1 U7035 ( .B1(DATAI_4_), .B2(keyinput_27), .C1(keyinput_26), .C2(
        DATAI_5_), .A(n6358), .ZN(n6359) );
  OAI21_X1 U7036 ( .B1(n6361), .B2(n6360), .A(n6359), .ZN(n6362) );
  OAI221_X1 U7037 ( .B1(DATAI_3_), .B2(n6363), .C1(n6470), .C2(keyinput_28), 
        .A(n6362), .ZN(n6364) );
  AOI22_X1 U7038 ( .A1(n6365), .A2(n6364), .B1(keyinput_31), .B2(DATAI_0_), 
        .ZN(n6366) );
  OAI21_X1 U7039 ( .B1(keyinput_31), .B2(DATAI_0_), .A(n6366), .ZN(n6367) );
  OAI221_X1 U7040 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n6368), .C1(n6476), .C2(
        keyinput_32), .A(n6367), .ZN(n6371) );
  INV_X1 U7041 ( .A(HOLD), .ZN(n7072) );
  AOI22_X1 U7042 ( .A1(keyinput_35), .A2(READY_N), .B1(n7072), .B2(keyinput_36), .ZN(n6369) );
  OAI221_X1 U7043 ( .B1(keyinput_35), .B2(READY_N), .C1(n7072), .C2(
        keyinput_36), .A(n6369), .ZN(n6370) );
  AOI21_X1 U7044 ( .B1(n6372), .B2(n6371), .A(n6370), .ZN(n6377) );
  INV_X1 U7045 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6727) );
  XOR2_X1 U7046 ( .A(n6727), .B(keyinput_37), .Z(n6376) );
  INV_X1 U7047 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6720) );
  OAI22_X1 U7048 ( .A1(n6720), .A2(keyinput_39), .B1(keyinput_38), .B2(
        ADS_N_REG_SCAN_IN), .ZN(n6373) );
  AOI221_X1 U7049 ( .B1(n6720), .B2(keyinput_39), .C1(ADS_N_REG_SCAN_IN), .C2(
        keyinput_38), .A(n6373), .ZN(n6375) );
  XNOR2_X1 U7050 ( .A(M_IO_N_REG_SCAN_IN), .B(keyinput_40), .ZN(n6374) );
  OAI211_X1 U7051 ( .C1(n6377), .C2(n6376), .A(n6375), .B(n6374), .ZN(n6378)
         );
  OAI211_X1 U7052 ( .C1(n6729), .C2(keyinput_42), .A(n6379), .B(n6378), .ZN(
        n6380) );
  AOI21_X1 U7053 ( .B1(n6729), .B2(keyinput_42), .A(n6380), .ZN(n6381) );
  AOI221_X1 U7054 ( .B1(MORE_REG_SCAN_IN), .B2(n6382), .C1(n7025), .C2(
        keyinput_44), .A(n6381), .ZN(n6383) );
  OAI22_X1 U7055 ( .A1(n6384), .A2(n6383), .B1(keyinput_47), .B2(
        BYTEENABLE_REG_0__SCAN_IN), .ZN(n6385) );
  AOI21_X1 U7056 ( .B1(keyinput_47), .B2(BYTEENABLE_REG_0__SCAN_IN), .A(n6385), 
        .ZN(n6392) );
  AOI22_X1 U7057 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_48), .B1(
        BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_49), .ZN(n6386) );
  OAI221_X1 U7058 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_48), .C1(
        BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_49), .A(n6386), .ZN(n6391) );
  OAI22_X1 U7059 ( .A1(REIP_REG_30__SCAN_IN), .A2(keyinput_52), .B1(
        BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_50), .ZN(n6387) );
  AOI221_X1 U7060 ( .B1(REIP_REG_30__SCAN_IN), .B2(keyinput_52), .C1(
        keyinput_50), .C2(BYTEENABLE_REG_3__SCAN_IN), .A(n6387), .ZN(n6390) );
  OAI22_X1 U7061 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_51), .B1(
        keyinput_53), .B2(REIP_REG_29__SCAN_IN), .ZN(n6388) );
  AOI221_X1 U7062 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_51), .C1(
        REIP_REG_29__SCAN_IN), .C2(keyinput_53), .A(n6388), .ZN(n6389) );
  OAI211_X1 U7063 ( .C1(n6392), .C2(n6391), .A(n6390), .B(n6389), .ZN(n6393)
         );
  AOI21_X1 U7064 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_54), .A(n6393), 
        .ZN(n6394) );
  OAI21_X1 U7065 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_54), .A(n6394), 
        .ZN(n6395) );
  AOI22_X1 U7066 ( .A1(keyinput_57), .A2(n6504), .B1(n6396), .B2(n6395), .ZN(
        n6397) );
  OAI21_X1 U7067 ( .B1(n6504), .B2(keyinput_57), .A(n6397), .ZN(n6398) );
  AOI22_X1 U7068 ( .A1(keyinput_60), .A2(n6401), .B1(n6399), .B2(n6398), .ZN(
        n6400) );
  OAI21_X1 U7069 ( .B1(n6401), .B2(keyinput_60), .A(n6400), .ZN(n6402) );
  OAI221_X1 U7070 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_61), .C1(n6638), 
        .C2(n6403), .A(n6402), .ZN(n6404) );
  OAI221_X1 U7071 ( .B1(REIP_REG_20__SCAN_IN), .B2(n6405), .C1(n6967), .C2(
        keyinput_62), .A(n6404), .ZN(n6407) );
  AOI21_X1 U7072 ( .B1(keyinput_63), .B2(n6407), .A(keyinput_127), .ZN(n6409)
         );
  INV_X1 U7073 ( .A(keyinput_63), .ZN(n6406) );
  AOI21_X1 U7074 ( .B1(n6407), .B2(n6406), .A(REIP_REG_19__SCAN_IN), .ZN(n6408) );
  AOI22_X1 U7075 ( .A1(n6409), .A2(REIP_REG_19__SCAN_IN), .B1(n6408), .B2(
        keyinput_127), .ZN(n6514) );
  OAI22_X1 U7076 ( .A1(n6643), .A2(keyinput_122), .B1(n6641), .B2(keyinput_123), .ZN(n6410) );
  AOI221_X1 U7077 ( .B1(n6643), .B2(keyinput_122), .C1(keyinput_123), .C2(
        n6641), .A(n6410), .ZN(n6508) );
  INV_X1 U7078 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6646) );
  AOI22_X1 U7079 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput_119), .B1(n6646), 
        .B2(keyinput_120), .ZN(n6411) );
  OAI221_X1 U7080 ( .B1(REIP_REG_27__SCAN_IN), .B2(keyinput_119), .C1(n6646), 
        .C2(keyinput_120), .A(n6411), .ZN(n6506) );
  INV_X1 U7081 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6679) );
  OAI22_X1 U7082 ( .A1(n6679), .A2(keyinput_112), .B1(
        BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_113), .ZN(n6412) );
  AOI221_X1 U7083 ( .B1(n6679), .B2(keyinput_112), .C1(keyinput_113), .C2(
        BYTEENABLE_REG_2__SCAN_IN), .A(n6412), .ZN(n6500) );
  AOI22_X1 U7084 ( .A1(n6728), .A2(keyinput_110), .B1(n7024), .B2(keyinput_109), .ZN(n6413) );
  OAI221_X1 U7085 ( .B1(n6728), .B2(keyinput_110), .C1(n7024), .C2(
        keyinput_109), .A(n6413), .ZN(n6494) );
  INV_X1 U7086 ( .A(keyinput_108), .ZN(n6491) );
  OAI22_X1 U7087 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_106), .B1(
        D_C_N_REG_SCAN_IN), .B2(keyinput_105), .ZN(n6414) );
  AOI221_X1 U7088 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_106), .C1(
        keyinput_105), .C2(D_C_N_REG_SCAN_IN), .A(n6414), .ZN(n6488) );
  INV_X1 U7089 ( .A(BS16_N), .ZN(n6572) );
  OAI22_X1 U7090 ( .A1(n6572), .A2(keyinput_98), .B1(NA_N), .B2(keyinput_97), 
        .ZN(n6415) );
  AOI221_X1 U7091 ( .B1(n6572), .B2(keyinput_98), .C1(keyinput_97), .C2(NA_N), 
        .A(n6415), .ZN(n6481) );
  INV_X1 U7092 ( .A(keyinput_96), .ZN(n6477) );
  OAI22_X1 U7093 ( .A1(n6417), .A2(keyinput_94), .B1(DATAI_2_), .B2(
        keyinput_93), .ZN(n6416) );
  AOI221_X1 U7094 ( .B1(n6417), .B2(keyinput_94), .C1(keyinput_93), .C2(
        DATAI_2_), .A(n6416), .ZN(n6473) );
  INV_X1 U7095 ( .A(keyinput_92), .ZN(n6471) );
  INV_X1 U7096 ( .A(keyinput_87), .ZN(n6461) );
  INV_X1 U7097 ( .A(keyinput_86), .ZN(n6458) );
  OAI22_X1 U7098 ( .A1(n6419), .A2(keyinput_85), .B1(keyinput_83), .B2(
        DATAI_12_), .ZN(n6418) );
  AOI221_X1 U7099 ( .B1(n6419), .B2(keyinput_85), .C1(DATAI_12_), .C2(
        keyinput_83), .A(n6418), .ZN(n6454) );
  INV_X1 U7100 ( .A(keyinput_82), .ZN(n6451) );
  OAI22_X1 U7101 ( .A1(DATAI_16_), .A2(keyinput_79), .B1(keyinput_80), .B2(
        DATAI_15_), .ZN(n6420) );
  AOI221_X1 U7102 ( .B1(DATAI_16_), .B2(keyinput_79), .C1(DATAI_15_), .C2(
        keyinput_80), .A(n6420), .ZN(n6447) );
  INV_X1 U7103 ( .A(keyinput_78), .ZN(n6445) );
  XNOR2_X1 U7104 ( .A(DATAI_27_), .B(keyinput_68), .ZN(n6435) );
  INV_X1 U7105 ( .A(keyinput_67), .ZN(n6427) );
  INV_X1 U7106 ( .A(keyinput_64), .ZN(n6423) );
  OAI22_X1 U7107 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(DATAI_29_), .B2(
        keyinput_66), .ZN(n6421) );
  AOI221_X1 U7108 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(keyinput_66), .C2(
        DATAI_29_), .A(n6421), .ZN(n6422) );
  OAI221_X1 U7109 ( .B1(DATAI_31_), .B2(keyinput_64), .C1(n6424), .C2(n6423), 
        .A(n6422), .ZN(n6425) );
  OAI221_X1 U7110 ( .B1(DATAI_28_), .B2(n6427), .C1(n6426), .C2(keyinput_67), 
        .A(n6425), .ZN(n6434) );
  INV_X1 U7111 ( .A(DATAI_25_), .ZN(n6430) );
  INV_X1 U7112 ( .A(DATAI_26_), .ZN(n6429) );
  AOI22_X1 U7113 ( .A1(n6430), .A2(keyinput_70), .B1(n6429), .B2(keyinput_69), 
        .ZN(n6428) );
  OAI221_X1 U7114 ( .B1(n6430), .B2(keyinput_70), .C1(n6429), .C2(keyinput_69), 
        .A(n6428), .ZN(n6433) );
  AOI22_X1 U7115 ( .A1(DATAI_23_), .A2(keyinput_72), .B1(DATAI_24_), .B2(
        keyinput_71), .ZN(n6431) );
  OAI221_X1 U7116 ( .B1(DATAI_23_), .B2(keyinput_72), .C1(DATAI_24_), .C2(
        keyinput_71), .A(n6431), .ZN(n6432) );
  AOI211_X1 U7117 ( .C1(n6435), .C2(n6434), .A(n6433), .B(n6432), .ZN(n6442)
         );
  XNOR2_X1 U7118 ( .A(DATAI_22_), .B(keyinput_73), .ZN(n6441) );
  OAI22_X1 U7119 ( .A1(n6437), .A2(keyinput_75), .B1(keyinput_76), .B2(
        DATAI_19_), .ZN(n6436) );
  AOI221_X1 U7120 ( .B1(n6437), .B2(keyinput_75), .C1(DATAI_19_), .C2(
        keyinput_76), .A(n6436), .ZN(n6440) );
  OAI22_X1 U7121 ( .A1(DATAI_18_), .A2(keyinput_77), .B1(keyinput_74), .B2(
        DATAI_21_), .ZN(n6438) );
  AOI221_X1 U7122 ( .B1(DATAI_18_), .B2(keyinput_77), .C1(DATAI_21_), .C2(
        keyinput_74), .A(n6438), .ZN(n6439) );
  OAI211_X1 U7123 ( .C1(n6442), .C2(n6441), .A(n6440), .B(n6439), .ZN(n6443)
         );
  OAI221_X1 U7124 ( .B1(DATAI_17_), .B2(n6445), .C1(n6444), .C2(keyinput_78), 
        .A(n6443), .ZN(n6446) );
  AOI22_X1 U7125 ( .A1(keyinput_81), .A2(n6449), .B1(n6447), .B2(n6446), .ZN(
        n6448) );
  OAI21_X1 U7126 ( .B1(n6449), .B2(keyinput_81), .A(n6448), .ZN(n6450) );
  OAI221_X1 U7127 ( .B1(DATAI_13_), .B2(keyinput_82), .C1(n6452), .C2(n6451), 
        .A(n6450), .ZN(n6453) );
  OAI211_X1 U7128 ( .C1(DATAI_11_), .C2(keyinput_84), .A(n6454), .B(n6453), 
        .ZN(n6455) );
  AOI21_X1 U7129 ( .B1(DATAI_11_), .B2(keyinput_84), .A(n6455), .ZN(n6456) );
  AOI221_X1 U7130 ( .B1(DATAI_9_), .B2(n6458), .C1(n6457), .C2(keyinput_86), 
        .A(n6456), .ZN(n6459) );
  AOI221_X1 U7131 ( .B1(DATAI_8_), .B2(n6461), .C1(n6460), .C2(keyinput_87), 
        .A(n6459), .ZN(n6468) );
  AOI22_X1 U7132 ( .A1(n6464), .A2(keyinput_88), .B1(keyinput_89), .B2(n6463), 
        .ZN(n6462) );
  OAI221_X1 U7133 ( .B1(n6464), .B2(keyinput_88), .C1(n6463), .C2(keyinput_89), 
        .A(n6462), .ZN(n6467) );
  OAI22_X1 U7134 ( .A1(DATAI_4_), .A2(keyinput_91), .B1(keyinput_90), .B2(
        DATAI_5_), .ZN(n6465) );
  AOI221_X1 U7135 ( .B1(DATAI_4_), .B2(keyinput_91), .C1(DATAI_5_), .C2(
        keyinput_90), .A(n6465), .ZN(n6466) );
  OAI21_X1 U7136 ( .B1(n6468), .B2(n6467), .A(n6466), .ZN(n6469) );
  OAI221_X1 U7137 ( .B1(DATAI_3_), .B2(n6471), .C1(n6470), .C2(keyinput_92), 
        .A(n6469), .ZN(n6472) );
  AOI22_X1 U7138 ( .A1(n6473), .A2(n6472), .B1(keyinput_95), .B2(DATAI_0_), 
        .ZN(n6474) );
  OAI21_X1 U7139 ( .B1(keyinput_95), .B2(DATAI_0_), .A(n6474), .ZN(n6475) );
  OAI221_X1 U7140 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n6477), .C1(n6476), .C2(
        keyinput_96), .A(n6475), .ZN(n6480) );
  AOI22_X1 U7141 ( .A1(HOLD), .A2(keyinput_100), .B1(READY_N), .B2(keyinput_99), .ZN(n6478) );
  OAI221_X1 U7142 ( .B1(HOLD), .B2(keyinput_100), .C1(READY_N), .C2(
        keyinput_99), .A(n6478), .ZN(n6479) );
  AOI21_X1 U7143 ( .B1(n6481), .B2(n6480), .A(n6479), .ZN(n6486) );
  XNOR2_X1 U7144 ( .A(n6727), .B(keyinput_101), .ZN(n6485) );
  OAI22_X1 U7145 ( .A1(n6720), .A2(keyinput_103), .B1(ADS_N_REG_SCAN_IN), .B2(
        keyinput_102), .ZN(n6482) );
  AOI221_X1 U7146 ( .B1(n6720), .B2(keyinput_103), .C1(keyinput_102), .C2(
        ADS_N_REG_SCAN_IN), .A(n6482), .ZN(n6484) );
  XNOR2_X1 U7147 ( .A(M_IO_N_REG_SCAN_IN), .B(keyinput_104), .ZN(n6483) );
  OAI211_X1 U7148 ( .C1(n6486), .C2(n6485), .A(n6484), .B(n6483), .ZN(n6487)
         );
  OAI211_X1 U7149 ( .C1(STATEBS16_REG_SCAN_IN), .C2(keyinput_107), .A(n6488), 
        .B(n6487), .ZN(n6489) );
  AOI21_X1 U7150 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_107), .A(n6489), 
        .ZN(n6490) );
  AOI221_X1 U7151 ( .B1(MORE_REG_SCAN_IN), .B2(n6491), .C1(n7025), .C2(
        keyinput_108), .A(n6490), .ZN(n6493) );
  NAND2_X1 U7152 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_111), .ZN(
        n6492) );
  OAI221_X1 U7153 ( .B1(n6494), .B2(n6493), .C1(BYTEENABLE_REG_0__SCAN_IN), 
        .C2(keyinput_111), .A(n6492), .ZN(n6499) );
  INV_X1 U7154 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6671) );
  AOI22_X1 U7155 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_117), .B1(n6671), 
        .B2(keyinput_114), .ZN(n6495) );
  OAI221_X1 U7156 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_117), .C1(n6671), 
        .C2(keyinput_114), .A(n6495), .ZN(n6498) );
  AOI22_X1 U7157 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_115), .B1(
        REIP_REG_30__SCAN_IN), .B2(keyinput_116), .ZN(n6496) );
  OAI221_X1 U7158 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_115), .C1(
        REIP_REG_30__SCAN_IN), .C2(keyinput_116), .A(n6496), .ZN(n6497) );
  AOI211_X1 U7159 ( .C1(n6500), .C2(n6499), .A(n6498), .B(n6497), .ZN(n6501)
         );
  OAI21_X1 U7160 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_118), .A(n6501), 
        .ZN(n6502) );
  AOI21_X1 U7161 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_118), .A(n6502), 
        .ZN(n6505) );
  NAND2_X1 U7162 ( .A1(n6504), .A2(keyinput_121), .ZN(n6503) );
  OAI221_X1 U7163 ( .B1(n6506), .B2(n6505), .C1(n6504), .C2(keyinput_121), .A(
        n6503), .ZN(n6507) );
  AOI22_X1 U7164 ( .A1(n6508), .A2(n6507), .B1(keyinput_124), .B2(
        REIP_REG_22__SCAN_IN), .ZN(n6509) );
  OAI21_X1 U7165 ( .B1(keyinput_124), .B2(REIP_REG_22__SCAN_IN), .A(n6509), 
        .ZN(n6512) );
  XOR2_X1 U7166 ( .A(REIP_REG_21__SCAN_IN), .B(keyinput_125), .Z(n6511) );
  XOR2_X1 U7167 ( .A(REIP_REG_20__SCAN_IN), .B(keyinput_126), .Z(n6510) );
  AOI21_X1 U7168 ( .B1(n6512), .B2(n6511), .A(n6510), .ZN(n6513) );
  NOR2_X1 U7169 ( .A1(n6514), .A2(n6513), .ZN(n6524) );
  OAI21_X1 U7170 ( .B1(n6516), .B2(n6836), .A(n6515), .ZN(n6519) );
  NOR2_X1 U7171 ( .A1(n6517), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6518)
         );
  AOI211_X1 U7172 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6520), .A(n6519), .B(n6518), .ZN(n6521) );
  OAI21_X1 U7173 ( .B1(n6522), .B2(n6756), .A(n6521), .ZN(n6523) );
  XOR2_X1 U7174 ( .A(n6524), .B(n6523), .Z(U2999) );
  INV_X1 U7175 ( .A(n6525), .ZN(n6530) );
  OAI21_X1 U7176 ( .B1(n6532), .B2(n6526), .A(n6768), .ZN(n6527) );
  OAI211_X1 U7177 ( .C1(n6530), .C2(n6529), .A(n6528), .B(n6527), .ZN(n6844)
         );
  INV_X1 U7178 ( .A(n6844), .ZN(n6534) );
  NAND2_X1 U7179 ( .A1(n6532), .A2(n6531), .ZN(n6533) );
  AOI21_X1 U7180 ( .B1(n6534), .B2(n6533), .A(n6537), .ZN(n6535) );
  AOI211_X1 U7181 ( .C1(n6846), .C2(n6959), .A(n6536), .B(n6535), .ZN(n6540)
         );
  NAND3_X1 U7182 ( .A1(n6538), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n6537), .ZN(n6539) );
  OAI211_X1 U7183 ( .C1(n6541), .C2(n6756), .A(n6540), .B(n6539), .ZN(U3000)
         );
  INV_X1 U7184 ( .A(n6542), .ZN(n6543) );
  OAI21_X1 U7185 ( .B1(n6544), .B2(n6543), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n6551) );
  INV_X1 U7186 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6611) );
  OAI22_X1 U7187 ( .A1(n6756), .A2(n6545), .B1(n6611), .B2(n6801), .ZN(n6546)
         );
  AOI21_X1 U7188 ( .B1(n6846), .B2(n6547), .A(n6546), .ZN(n6550) );
  NAND3_X1 U7189 ( .A1(n6825), .A2(n5052), .A3(n6548), .ZN(n6549) );
  NAND3_X1 U7190 ( .A1(n6551), .A2(n6550), .A3(n6549), .ZN(U3017) );
  NAND2_X1 U7191 ( .A1(n7000), .A2(n6552), .ZN(n6557) );
  OAI21_X1 U7192 ( .B1(n6555), .B2(n6554), .A(n6553), .ZN(n6556) );
  NAND2_X1 U7193 ( .A1(n6557), .A2(n6556), .ZN(n6558) );
  AOI21_X1 U7194 ( .B1(n4843), .B2(n6559), .A(n6558), .ZN(n7004) );
  INV_X1 U7195 ( .A(n6560), .ZN(n6569) );
  INV_X1 U7196 ( .A(n4949), .ZN(n6563) );
  AOI22_X1 U7197 ( .A1(n6564), .A2(n6563), .B1(n6562), .B2(n6561), .ZN(n6565)
         );
  OAI21_X1 U7198 ( .B1(n7004), .B2(n6569), .A(n6565), .ZN(n6566) );
  MUX2_X1 U7199 ( .A(n6566), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(n6995), 
        .Z(U3460) );
  INV_X1 U7200 ( .A(n6567), .ZN(n6570) );
  OAI22_X1 U7201 ( .A1(n6570), .A2(n6569), .B1(n6568), .B2(n7047), .ZN(n6571)
         );
  MUX2_X1 U7202 ( .A(n6571), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6995), 
        .Z(U3456) );
  INV_X1 U7203 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U7204 ( .A1(STATE_REG_1__SCAN_IN), .A2(n7075), .ZN(n6644) );
  NAND2_X1 U7205 ( .A1(STATE_REG_0__SCAN_IN), .A2(n7071), .ZN(n6575) );
  NAND2_X1 U7206 ( .A1(n6644), .A2(n6575), .ZN(n6573) );
  CLKBUF_X1 U7207 ( .A(n6573), .Z(n7064) );
  NAND2_X1 U7208 ( .A1(n7074), .A2(n7075), .ZN(n6723) );
  AOI21_X1 U7209 ( .B1(n6572), .B2(n6723), .A(n7064), .ZN(n7063) );
  AOI21_X1 U7210 ( .B1(n6673), .B2(n7064), .A(n7063), .ZN(U3451) );
  AND2_X1 U7211 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n7064), .ZN(U3180) );
  AND2_X1 U7212 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6573), .ZN(U3179) );
  AND2_X1 U7213 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6573), .ZN(U3178) );
  AND2_X1 U7214 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6573), .ZN(U3177) );
  AND2_X1 U7215 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6573), .ZN(U3176) );
  AND2_X1 U7216 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n7064), .ZN(U3175) );
  AND2_X1 U7217 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n7064), .ZN(U3174) );
  AND2_X1 U7218 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n7064), .ZN(U3173) );
  AND2_X1 U7219 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n7064), .ZN(U3172) );
  AND2_X1 U7220 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n7064), .ZN(U3171) );
  AND2_X1 U7221 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6573), .ZN(U3170) );
  AND2_X1 U7222 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6573), .ZN(U3169) );
  AND2_X1 U7223 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6573), .ZN(U3168) );
  AND2_X1 U7224 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6573), .ZN(U3167) );
  AND2_X1 U7225 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6573), .ZN(U3166) );
  AND2_X1 U7226 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6573), .ZN(U3165) );
  AND2_X1 U7227 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6573), .ZN(U3164) );
  AND2_X1 U7228 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6573), .ZN(U3163) );
  AND2_X1 U7229 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6573), .ZN(U3162) );
  AND2_X1 U7230 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6573), .ZN(U3161) );
  AND2_X1 U7231 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n7064), .ZN(U3160) );
  AND2_X1 U7232 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n7064), .ZN(U3159) );
  AND2_X1 U7233 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n7064), .ZN(U3158) );
  AND2_X1 U7234 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6573), .ZN(U3157) );
  AND2_X1 U7235 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n7064), .ZN(U3156) );
  AND2_X1 U7236 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n7064), .ZN(U3155) );
  AND2_X1 U7237 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n7064), .ZN(U3154) );
  AND2_X1 U7238 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n7064), .ZN(U3153) );
  AND2_X1 U7239 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n7064), .ZN(U3152) );
  AND2_X1 U7240 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n7064), .ZN(U3151) );
  INV_X1 U7241 ( .A(n7061), .ZN(n6574) );
  AND2_X1 U7242 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6574), .ZN(U3019)
         );
  AND2_X1 U7243 ( .A1(n6590), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U7244 ( .A(n6644), .ZN(n7083) );
  INV_X1 U7245 ( .A(n7083), .ZN(n7084) );
  OAI21_X1 U7246 ( .B1(n6575), .B2(ADS_N_REG_SCAN_IN), .A(n7084), .ZN(n6576)
         );
  INV_X1 U7247 ( .A(n6576), .ZN(U2789) );
  AOI22_X1 U7248 ( .A1(n6741), .A2(LWORD_REG_0__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6578) );
  OAI21_X1 U7249 ( .B1(n6579), .B2(n6608), .A(n6578), .ZN(U2923) );
  AOI22_X1 U7250 ( .A1(n6741), .A2(LWORD_REG_1__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6580) );
  OAI21_X1 U7251 ( .B1(n6581), .B2(n6608), .A(n6580), .ZN(U2922) );
  AOI22_X1 U7252 ( .A1(n6741), .A2(LWORD_REG_2__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6582) );
  OAI21_X1 U7253 ( .B1(n6583), .B2(n6608), .A(n6582), .ZN(U2921) );
  AOI22_X1 U7254 ( .A1(n6741), .A2(LWORD_REG_3__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6584) );
  OAI21_X1 U7255 ( .B1(n6585), .B2(n6608), .A(n6584), .ZN(U2920) );
  AOI22_X1 U7256 ( .A1(n6741), .A2(LWORD_REG_4__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6586) );
  OAI21_X1 U7257 ( .B1(n6587), .B2(n6608), .A(n6586), .ZN(U2919) );
  AOI22_X1 U7258 ( .A1(n6741), .A2(LWORD_REG_5__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6588) );
  OAI21_X1 U7259 ( .B1(n6589), .B2(n6608), .A(n6588), .ZN(U2918) );
  AOI22_X1 U7260 ( .A1(n6741), .A2(LWORD_REG_6__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6591) );
  OAI21_X1 U7261 ( .B1(n6592), .B2(n6608), .A(n6591), .ZN(U2917) );
  AOI22_X1 U7262 ( .A1(n6741), .A2(LWORD_REG_7__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6593) );
  OAI21_X1 U7263 ( .B1(n4031), .B2(n6608), .A(n6593), .ZN(U2916) );
  AOI22_X1 U7264 ( .A1(n6741), .A2(LWORD_REG_8__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6594) );
  OAI21_X1 U7265 ( .B1(n6595), .B2(n6608), .A(n6594), .ZN(U2915) );
  AOI22_X1 U7266 ( .A1(n6741), .A2(LWORD_REG_9__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6596) );
  OAI21_X1 U7267 ( .B1(n6597), .B2(n6608), .A(n6596), .ZN(U2914) );
  AOI22_X1 U7268 ( .A1(n6741), .A2(LWORD_REG_10__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6598) );
  OAI21_X1 U7269 ( .B1(n6599), .B2(n6608), .A(n6598), .ZN(U2913) );
  AOI22_X1 U7270 ( .A1(n6741), .A2(LWORD_REG_11__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6600) );
  OAI21_X1 U7271 ( .B1(n6601), .B2(n6608), .A(n6600), .ZN(U2912) );
  AOI22_X1 U7272 ( .A1(n6741), .A2(LWORD_REG_12__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6602) );
  OAI21_X1 U7273 ( .B1(n4093), .B2(n6608), .A(n6602), .ZN(U2911) );
  AOI22_X1 U7274 ( .A1(n6741), .A2(LWORD_REG_13__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6603) );
  OAI21_X1 U7275 ( .B1(n6604), .B2(n6608), .A(n6603), .ZN(U2910) );
  AOI22_X1 U7276 ( .A1(n6741), .A2(LWORD_REG_14__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6605) );
  OAI21_X1 U7277 ( .B1(n4130), .B2(n6608), .A(n6605), .ZN(U2909) );
  AOI22_X1 U7278 ( .A1(n6741), .A2(LWORD_REG_15__SCAN_IN), .B1(n6590), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6607) );
  OAI21_X1 U7279 ( .B1(n6609), .B2(n6608), .A(n6607), .ZN(U2908) );
  NOR2_X2 U7280 ( .A1(n7074), .A2(n7084), .ZN(n6656) );
  NAND2_X1 U7281 ( .A1(n7074), .A2(n7083), .ZN(n6658) );
  INV_X1 U7282 ( .A(n6658), .ZN(n6652) );
  AOI22_X1 U7283 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6644), .ZN(n6610) );
  OAI21_X1 U7284 ( .B1(n6611), .B2(n6654), .A(n6610), .ZN(U3184) );
  AOI22_X1 U7285 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6644), .ZN(n6612) );
  OAI21_X1 U7286 ( .B1(n6614), .B2(n6658), .A(n6612), .ZN(U3185) );
  AOI22_X1 U7287 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6644), .ZN(n6613) );
  OAI21_X1 U7288 ( .B1(n6614), .B2(n6654), .A(n6613), .ZN(U3186) );
  AOI22_X1 U7289 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6644), .ZN(n6615) );
  OAI21_X1 U7290 ( .B1(n6855), .B2(n6654), .A(n6615), .ZN(U3187) );
  AOI22_X1 U7291 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6644), .ZN(n6616) );
  OAI21_X1 U7292 ( .B1(n6617), .B2(n6654), .A(n6616), .ZN(U3188) );
  AOI22_X1 U7293 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6644), .ZN(n6618) );
  OAI21_X1 U7294 ( .B1(n6620), .B2(n6658), .A(n6618), .ZN(U3189) );
  AOI22_X1 U7295 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6644), .ZN(n6619) );
  OAI21_X1 U7296 ( .B1(n6620), .B2(n6654), .A(n6619), .ZN(U3190) );
  AOI22_X1 U7297 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6644), .ZN(n6621) );
  OAI21_X1 U7298 ( .B1(n6623), .B2(n6658), .A(n6621), .ZN(U3191) );
  AOI22_X1 U7299 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6644), .ZN(n6622) );
  OAI21_X1 U7300 ( .B1(n6623), .B2(n6654), .A(n6622), .ZN(U3192) );
  AOI22_X1 U7301 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6644), .ZN(n6624) );
  OAI21_X1 U7302 ( .B1(n6907), .B2(n6658), .A(n6624), .ZN(U3193) );
  INV_X1 U7303 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6917) );
  AOI22_X1 U7304 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6644), .ZN(n6625) );
  OAI21_X1 U7305 ( .B1(n6917), .B2(n6658), .A(n6625), .ZN(U3194) );
  AOI22_X1 U7306 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6644), .ZN(n6626) );
  OAI21_X1 U7307 ( .B1(n6917), .B2(n6654), .A(n6626), .ZN(U3195) );
  INV_X1 U7308 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U7309 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6644), .ZN(n6627) );
  OAI21_X1 U7310 ( .B1(n6629), .B2(n6658), .A(n6627), .ZN(U3196) );
  AOI22_X1 U7311 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n7084), .ZN(n6628) );
  OAI21_X1 U7312 ( .B1(n6629), .B2(n6654), .A(n6628), .ZN(U3197) );
  AOI22_X1 U7313 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6644), .ZN(n6630) );
  OAI21_X1 U7314 ( .B1(n6198), .B2(n6654), .A(n6630), .ZN(U3198) );
  AOI22_X1 U7315 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6644), .ZN(n6631) );
  OAI21_X1 U7316 ( .B1(n6633), .B2(n6658), .A(n6631), .ZN(U3199) );
  AOI22_X1 U7317 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6644), .ZN(n6632) );
  OAI21_X1 U7318 ( .B1(n6633), .B2(n6654), .A(n6632), .ZN(U3200) );
  INV_X1 U7319 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6958) );
  AOI22_X1 U7320 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6644), .ZN(n6634) );
  OAI21_X1 U7321 ( .B1(n6958), .B2(n6654), .A(n6634), .ZN(U3201) );
  AOI22_X1 U7322 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6644), .ZN(n6635) );
  OAI21_X1 U7323 ( .B1(n6967), .B2(n6658), .A(n6635), .ZN(U3202) );
  AOI22_X1 U7324 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n7084), .ZN(n6636) );
  OAI21_X1 U7325 ( .B1(n6638), .B2(n6658), .A(n6636), .ZN(U3203) );
  AOI22_X1 U7326 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6644), .ZN(n6637) );
  OAI21_X1 U7327 ( .B1(n6638), .B2(n6654), .A(n6637), .ZN(U3204) );
  AOI22_X1 U7328 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n7084), .ZN(n6639) );
  OAI21_X1 U7329 ( .B1(n6641), .B2(n6658), .A(n6639), .ZN(U3205) );
  AOI22_X1 U7330 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6644), .ZN(n6640) );
  OAI21_X1 U7331 ( .B1(n6641), .B2(n6654), .A(n6640), .ZN(U3206) );
  AOI22_X1 U7332 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6644), .ZN(n6642) );
  OAI21_X1 U7333 ( .B1(n6643), .B2(n6654), .A(n6642), .ZN(U3207) );
  AOI22_X1 U7334 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6644), .ZN(n6645) );
  OAI21_X1 U7335 ( .B1(n6646), .B2(n6658), .A(n6645), .ZN(U3208) );
  AOI22_X1 U7336 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n7084), .ZN(n6647) );
  OAI21_X1 U7337 ( .B1(n6649), .B2(n6658), .A(n6647), .ZN(U3209) );
  AOI22_X1 U7338 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n7084), .ZN(n6648) );
  OAI21_X1 U7339 ( .B1(n6649), .B2(n6654), .A(n6648), .ZN(U3210) );
  AOI22_X1 U7340 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n7084), .ZN(n6650) );
  OAI21_X1 U7341 ( .B1(n6651), .B2(n6654), .A(n6650), .ZN(U3211) );
  AOI22_X1 U7342 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6652), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n7084), .ZN(n6653) );
  OAI21_X1 U7343 ( .B1(n6655), .B2(n6654), .A(n6653), .ZN(U3212) );
  INV_X1 U7344 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6659) );
  AOI22_X1 U7345 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6656), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n7084), .ZN(n6657) );
  OAI21_X1 U7346 ( .B1(n6659), .B2(n6658), .A(n6657), .ZN(U3213) );
  MUX2_X1 U7347 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n7084), .Z(U3445) );
  NOR4_X1 U7348 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6663) );
  NOR4_X1 U7349 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6662) );
  NOR4_X1 U7350 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(
        n6661) );
  NOR4_X1 U7351 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6660) );
  NAND4_X1 U7352 ( .A1(n6663), .A2(n6662), .A3(n6661), .A4(n6660), .ZN(n6669)
         );
  NOR4_X1 U7353 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6667) );
  AOI211_X1 U7354 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_31__SCAN_IN), .B(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6666) );
  NOR4_X1 U7355 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6665) );
  NOR4_X1 U7356 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6664) );
  NAND4_X1 U7357 ( .A1(n6667), .A2(n6666), .A3(n6665), .A4(n6664), .ZN(n6668)
         );
  NOR2_X1 U7358 ( .A1(n6669), .A2(n6668), .ZN(n6683) );
  NOR3_X1 U7359 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6677) );
  NOR2_X1 U7360 ( .A1(REIP_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .ZN(n6674) );
  OAI21_X1 U7361 ( .B1(n6677), .B2(n6674), .A(n6683), .ZN(n6670) );
  OAI21_X1 U7362 ( .B1(n6683), .B2(n6671), .A(n6670), .ZN(U2795) );
  MUX2_X1 U7363 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n7084), .Z(U3446) );
  NOR3_X1 U7364 ( .A1(n6673), .A2(REIP_REG_0__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n6672) );
  AOI221_X1 U7365 ( .B1(n6674), .B2(n6673), .C1(REIP_REG_1__SCAN_IN), .C2(
        REIP_REG_0__SCAN_IN), .A(n6672), .ZN(n6676) );
  INV_X1 U7366 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6675) );
  INV_X1 U7367 ( .A(n6683), .ZN(n6680) );
  AOI22_X1 U7368 ( .A1(n6683), .A2(n6676), .B1(n6675), .B2(n6680), .ZN(U3468)
         );
  MUX2_X1 U7369 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n7084), .Z(U3447) );
  OAI21_X1 U7370 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6677), .A(n6683), .ZN(n6678)
         );
  OAI21_X1 U7371 ( .B1(n6683), .B2(n6679), .A(n6678), .ZN(U2794) );
  MUX2_X1 U7372 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n7084), .Z(U3448) );
  NOR2_X1 U7373 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6682) );
  INV_X1 U7374 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6681) );
  AOI22_X1 U7375 ( .A1(n6683), .A2(n6682), .B1(n6681), .B2(n6680), .ZN(U3469)
         );
  AOI22_X1 U7376 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6691), .B1(n6843), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6689) );
  OAI22_X1 U7377 ( .A1(n6686), .A2(n6993), .B1(n6685), .B2(n6684), .ZN(n6687)
         );
  INV_X1 U7378 ( .A(n6687), .ZN(n6688) );
  OAI211_X1 U7379 ( .C1(n6707), .C2(n6690), .A(n6689), .B(n6688), .ZN(U2984)
         );
  AOI22_X1 U7380 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6691), .B1(n6843), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U7381 ( .A1(n6694), .A2(n6693), .ZN(n6695) );
  XNOR2_X1 U7382 ( .A(n6692), .B(n6695), .ZN(n6770) );
  AOI22_X1 U7383 ( .A1(n6704), .A2(n6770), .B1(n6696), .B2(n6710), .ZN(n6697)
         );
  OAI211_X1 U7384 ( .C1(n6707), .C2(n6885), .A(n6698), .B(n6697), .ZN(U2980)
         );
  AOI22_X1 U7385 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n6691), .B1(n6843), 
        .B2(REIP_REG_7__SCAN_IN), .ZN(n6706) );
  OAI21_X1 U7386 ( .B1(n6699), .B2(n6702), .A(n6700), .ZN(n6703) );
  INV_X1 U7387 ( .A(n6703), .ZN(n6789) );
  AOI22_X1 U7388 ( .A1(n6789), .A2(n6704), .B1(n6710), .B2(n6893), .ZN(n6705)
         );
  OAI211_X1 U7389 ( .C1(n6707), .C2(n6902), .A(n6706), .B(n6705), .ZN(U2979)
         );
  AOI22_X1 U7390 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6691), .B1(n6843), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n6712) );
  INV_X1 U7391 ( .A(n6708), .ZN(n6911) );
  AOI22_X1 U7392 ( .A1(n6911), .A2(n6710), .B1(n6709), .B2(n6910), .ZN(n6711)
         );
  OAI211_X1 U7393 ( .C1(n6713), .C2(n6993), .A(n6712), .B(n6711), .ZN(U2975)
         );
  INV_X1 U7394 ( .A(n6988), .ZN(n6719) );
  INV_X1 U7395 ( .A(n6714), .ZN(n6718) );
  INV_X1 U7396 ( .A(n6715), .ZN(n6984) );
  OAI21_X1 U7397 ( .B1(n6716), .B2(n6984), .A(n4672), .ZN(n6717) );
  OAI21_X1 U7398 ( .B1(n6719), .B2(n6718), .A(n6717), .ZN(n6989) );
  NOR2_X1 U7399 ( .A1(n6989), .A2(n7051), .ZN(n6721) );
  OAI22_X1 U7400 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7034), .B1(n6721), .B2(
        n6720), .ZN(U2790) );
  NOR2_X1 U7401 ( .A1(n7083), .A2(D_C_N_REG_SCAN_IN), .ZN(n6722) );
  AOI22_X1 U7402 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7083), .B1(n6723), .B2(
        n6722), .ZN(U2791) );
  NOR2_X1 U7403 ( .A1(n6724), .A2(n4407), .ZN(n6737) );
  NAND2_X1 U7404 ( .A1(n6739), .A2(n6737), .ZN(n6725) );
  OAI211_X1 U7405 ( .C1(n6739), .C2(n6727), .A(n6726), .B(n6725), .ZN(U3474)
         );
  AOI22_X1 U7406 ( .A1(n7083), .A2(READREQUEST_REG_SCAN_IN), .B1(n6728), .B2(
        n7084), .ZN(U3470) );
  NOR2_X1 U7407 ( .A1(n7074), .A2(n7072), .ZN(n7066) );
  NOR2_X1 U7408 ( .A1(n7075), .A2(n6729), .ZN(n7078) );
  AOI21_X1 U7409 ( .B1(HOLD), .B2(STATE_REG_1__SCAN_IN), .A(n7078), .ZN(n6731)
         );
  NAND2_X1 U7410 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n7079) );
  OAI211_X1 U7411 ( .C1(n7066), .C2(n6731), .A(n6730), .B(n7079), .ZN(U3182)
         );
  NOR2_X1 U7412 ( .A1(n7046), .A2(n6732), .ZN(n7033) );
  AOI21_X1 U7413 ( .B1(n7033), .B2(n7028), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6734) );
  OAI21_X1 U7414 ( .B1(n6735), .B2(n6734), .A(n6733), .ZN(U3150) );
  OAI21_X1 U7415 ( .B1(n6737), .B2(n6736), .A(n7028), .ZN(n6990) );
  AOI211_X1 U7416 ( .C1(n4407), .C2(n7126), .A(n7128), .B(n6990), .ZN(n6738)
         );
  OAI21_X1 U7417 ( .B1(n6738), .B2(n7046), .A(n7048), .ZN(n6743) );
  AOI211_X1 U7418 ( .C1(n6741), .C2(n7028), .A(n6740), .B(n6739), .ZN(n6742)
         );
  MUX2_X1 U7419 ( .A(n6743), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6742), .Z(
        U3472) );
  OAI21_X1 U7420 ( .B1(n6746), .B2(n6745), .A(n6744), .ZN(n6763) );
  NAND2_X1 U7421 ( .A1(n6764), .A2(n6763), .ZN(n6784) );
  OAI21_X1 U7422 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6747), .ZN(n6754) );
  INV_X1 U7423 ( .A(n6781), .ZN(n6752) );
  NAND2_X1 U7424 ( .A1(n6846), .A2(n6852), .ZN(n6748) );
  OAI211_X1 U7425 ( .C1(n6750), .C2(n6756), .A(n6749), .B(n6748), .ZN(n6751)
         );
  AOI21_X1 U7426 ( .B1(n6752), .B2(INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6751), 
        .ZN(n6753) );
  OAI21_X1 U7427 ( .B1(n6784), .B2(n6754), .A(n6753), .ZN(U3014) );
  AOI22_X1 U7428 ( .A1(n6846), .A2(n6755), .B1(n6843), .B2(REIP_REG_3__SCAN_IN), .ZN(n6759) );
  NAND2_X1 U7429 ( .A1(n6847), .A2(n6757), .ZN(n6758) );
  OAI211_X1 U7430 ( .C1(n6784), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6759), 
        .B(n6758), .ZN(n6760) );
  INV_X1 U7431 ( .A(n6760), .ZN(n6761) );
  OAI21_X1 U7432 ( .B1(n6781), .B2(n6762), .A(n6761), .ZN(U3015) );
  NAND4_X1 U7433 ( .A1(n6765), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6764), 
        .A4(n6763), .ZN(n6774) );
  AOI211_X1 U7434 ( .C1(n6768), .C2(n4568), .A(n6767), .B(n6766), .ZN(n6772)
         );
  OAI22_X1 U7435 ( .A1(n6836), .A2(n6881), .B1(n6891), .B2(n6801), .ZN(n6769)
         );
  AOI21_X1 U7436 ( .B1(n6770), .B2(n6847), .A(n6769), .ZN(n6771) );
  OAI221_X1 U7437 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6774), .C1(n6773), .C2(n6772), .A(n6771), .ZN(U3012) );
  INV_X1 U7438 ( .A(n6775), .ZN(n6776) );
  AOI21_X1 U7439 ( .B1(n6846), .B2(n6777), .A(n6776), .ZN(n6788) );
  AOI22_X1 U7440 ( .A1(n6781), .A2(n6780), .B1(n6779), .B2(n6778), .ZN(n6794)
         );
  INV_X1 U7441 ( .A(n6782), .ZN(n6783) );
  AOI22_X1 U7442 ( .A1(n6794), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .B1(n6847), 
        .B2(n6783), .ZN(n6787) );
  NOR2_X1 U7443 ( .A1(n6785), .A2(n6784), .ZN(n6796) );
  OAI211_X1 U7444 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6796), .B(n6795), .ZN(n6786) );
  NAND3_X1 U7445 ( .A1(n6788), .A2(n6787), .A3(n6786), .ZN(U3010) );
  INV_X1 U7446 ( .A(n6794), .ZN(n6792) );
  AOI22_X1 U7447 ( .A1(n6846), .A2(n6890), .B1(n6843), .B2(REIP_REG_7__SCAN_IN), .ZN(n6791) );
  AOI22_X1 U7448 ( .A1(n6796), .A2(n6793), .B1(n6847), .B2(n6789), .ZN(n6790)
         );
  OAI211_X1 U7449 ( .C1(n6793), .C2(n6792), .A(n6791), .B(n6790), .ZN(U3011)
         );
  AOI21_X1 U7450 ( .B1(n6825), .B2(n6795), .A(n6794), .ZN(n6812) );
  NAND2_X1 U7451 ( .A1(n6797), .A2(n6796), .ZN(n6813) );
  AOI221_X1 U7452 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n4601), .C2(n6807), .A(n6813), 
        .ZN(n6805) );
  AND2_X1 U7453 ( .A1(n6798), .A2(n6847), .ZN(n6804) );
  NAND2_X1 U7454 ( .A1(n6846), .A2(n6799), .ZN(n6800) );
  OAI21_X1 U7455 ( .B1(n6802), .B2(n6801), .A(n6800), .ZN(n6803) );
  NOR3_X1 U7456 ( .A1(n6805), .A2(n6804), .A3(n6803), .ZN(n6806) );
  OAI21_X1 U7457 ( .B1(n6812), .B2(n6807), .A(n6806), .ZN(U3008) );
  INV_X1 U7458 ( .A(n6808), .ZN(n6809) );
  AOI222_X1 U7459 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6843), .B1(n6846), .B2(
        n6810), .C1(n6847), .C2(n6809), .ZN(n6811) );
  OAI221_X1 U7460 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n6813), .C1(n4601), .C2(n6812), .A(n6811), .ZN(U3009) );
  INV_X1 U7461 ( .A(n6814), .ZN(n6816) );
  AOI21_X1 U7462 ( .B1(n6846), .B2(n6816), .A(n6815), .ZN(n6822) );
  AOI22_X1 U7463 ( .A1(n6817), .A2(n6847), .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6823), .ZN(n6821) );
  OAI211_X1 U7464 ( .C1(INSTADDRPOINTER_REG_12__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .A(n6819), .B(n6818), .ZN(n6820) );
  NAND3_X1 U7465 ( .A1(n6822), .A2(n6821), .A3(n6820), .ZN(U3006) );
  AOI21_X1 U7466 ( .B1(n6825), .B2(n6824), .A(n6823), .ZN(n6842) );
  INV_X1 U7467 ( .A(n6826), .ZN(n6828) );
  AOI21_X1 U7468 ( .B1(n6828), .B2(n6846), .A(n6827), .ZN(n6831) );
  AOI22_X1 U7469 ( .A1(n6829), .A2(n6847), .B1(n6833), .B2(n6832), .ZN(n6830)
         );
  OAI211_X1 U7470 ( .C1(n6842), .C2(n6832), .A(n6831), .B(n6830), .ZN(U3003)
         );
  OAI211_X1 U7471 ( .C1(INSTADDRPOINTER_REG_16__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A(n6834), .B(n6833), .ZN(n6835) );
  INV_X1 U7472 ( .A(n6835), .ZN(n6839) );
  OAI22_X1 U7473 ( .A1(n6837), .A2(n6756), .B1(n6836), .B2(n6953), .ZN(n6838)
         );
  AOI211_X1 U7474 ( .C1(REIP_REG_16__SCAN_IN), .C2(n6843), .A(n6839), .B(n6838), .ZN(n6840) );
  OAI21_X1 U7475 ( .B1(n6842), .B2(n6841), .A(n6840), .ZN(U3002) );
  AOI22_X1 U7476 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6844), .B1(n6843), .B2(REIP_REG_17__SCAN_IN), .ZN(n6850) );
  AOI22_X1 U7477 ( .A1(n6848), .A2(n6847), .B1(n6846), .B2(n6845), .ZN(n6849)
         );
  OAI211_X1 U7478 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n6851), .A(n6850), .B(n6849), .ZN(U3001) );
  AOI22_X1 U7479 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6972), .B1(n6930), .B2(n6852), 
        .ZN(n6864) );
  NOR3_X1 U7480 ( .A1(n6905), .A2(n6853), .A3(REIP_REG_4__SCAN_IN), .ZN(n6862)
         );
  INV_X1 U7481 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6856) );
  OAI22_X1 U7482 ( .A1(n6856), .A2(n6981), .B1(n6855), .B2(n6854), .ZN(n6861)
         );
  OAI22_X1 U7483 ( .A1(n6859), .A2(n6858), .B1(n6857), .B2(n6973), .ZN(n6860)
         );
  NOR4_X1 U7484 ( .A1(n6954), .A2(n6862), .A3(n6861), .A4(n6860), .ZN(n6863)
         );
  OAI211_X1 U7485 ( .C1(n6866), .C2(n6865), .A(n6864), .B(n6863), .ZN(U2823)
         );
  AOI22_X1 U7486 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n6955), .B1(
        EBX_REG_5__SCAN_IN), .B2(n6972), .ZN(n6880) );
  AOI21_X1 U7487 ( .B1(n6930), .B2(n6867), .A(n6954), .ZN(n6879) );
  INV_X1 U7488 ( .A(n6868), .ZN(n6869) );
  AOI22_X1 U7489 ( .A1(n6871), .A2(n6870), .B1(n6950), .B2(n6869), .ZN(n6878)
         );
  INV_X1 U7490 ( .A(n6872), .ZN(n6873) );
  NOR2_X1 U7491 ( .A1(n6905), .A2(n6873), .ZN(n6884) );
  INV_X1 U7492 ( .A(n6874), .ZN(n6876) );
  OAI21_X1 U7493 ( .B1(n6905), .B2(n6876), .A(n6875), .ZN(n6898) );
  OAI21_X1 U7494 ( .B1(n6884), .B2(REIP_REG_5__SCAN_IN), .A(n6898), .ZN(n6877)
         );
  NAND4_X1 U7495 ( .A1(n6880), .A2(n6879), .A3(n6878), .A4(n6877), .ZN(U2822)
         );
  OAI22_X1 U7496 ( .A1(n6882), .A2(n6933), .B1(n6975), .B2(n6881), .ZN(n6883)
         );
  AOI211_X1 U7497 ( .C1(n6955), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6954), 
        .B(n6883), .ZN(n6889) );
  NAND2_X1 U7498 ( .A1(n6884), .A2(REIP_REG_5__SCAN_IN), .ZN(n6892) );
  NOR2_X1 U7499 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6892), .ZN(n6899) );
  OAI22_X1 U7500 ( .A1(n6886), .A2(n6961), .B1(n6885), .B2(n6973), .ZN(n6887)
         );
  AOI211_X1 U7501 ( .C1(REIP_REG_6__SCAN_IN), .C2(n6898), .A(n6899), .B(n6887), 
        .ZN(n6888) );
  NAND2_X1 U7502 ( .A1(n6889), .A2(n6888), .ZN(U2821) );
  AOI22_X1 U7503 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6972), .B1(n6930), .B2(n6890), 
        .ZN(n6897) );
  AOI21_X1 U7504 ( .B1(n6955), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6954), 
        .ZN(n6896) );
  OR3_X1 U7505 ( .A1(n6892), .A2(n6891), .A3(REIP_REG_7__SCAN_IN), .ZN(n6895)
         );
  NAND2_X1 U7506 ( .A1(n6978), .A2(n6893), .ZN(n6894) );
  AND4_X1 U7507 ( .A1(n6897), .A2(n6896), .A3(n6895), .A4(n6894), .ZN(n6901)
         );
  OAI21_X1 U7508 ( .B1(n6899), .B2(n6898), .A(REIP_REG_7__SCAN_IN), .ZN(n6900)
         );
  OAI211_X1 U7509 ( .C1(n6973), .C2(n6902), .A(n6901), .B(n6900), .ZN(U2820)
         );
  AOI22_X1 U7510 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n6955), .B1(n6930), 
        .B2(n6903), .ZN(n6915) );
  INV_X1 U7511 ( .A(n6923), .ZN(n6908) );
  OR3_X1 U7512 ( .A1(n6905), .A2(REIP_REG_11__SCAN_IN), .A3(n6904), .ZN(n6906)
         );
  OAI21_X1 U7513 ( .B1(n6908), .B2(n6907), .A(n6906), .ZN(n6909) );
  AOI21_X1 U7514 ( .B1(EBX_REG_11__SCAN_IN), .B2(n6972), .A(n6909), .ZN(n6914)
         );
  AOI22_X1 U7515 ( .A1(n6911), .A2(n6978), .B1(n6950), .B2(n6910), .ZN(n6913)
         );
  NAND4_X1 U7516 ( .A1(n6915), .A2(n6914), .A3(n6913), .A4(n6912), .ZN(U2816)
         );
  AOI22_X1 U7517 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6972), .B1(n6930), .B2(n6916), .ZN(n6928) );
  NOR3_X1 U7518 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6917), .A3(n6931), .ZN(n6918) );
  AOI211_X1 U7519 ( .C1(n6955), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6954), 
        .B(n6918), .ZN(n6927) );
  INV_X1 U7520 ( .A(n6919), .ZN(n6922) );
  INV_X1 U7521 ( .A(n6920), .ZN(n6921) );
  AOI22_X1 U7522 ( .A1(n6922), .A2(n6978), .B1(n6921), .B2(n6950), .ZN(n6926)
         );
  OAI21_X1 U7523 ( .B1(n6924), .B2(n6923), .A(REIP_REG_13__SCAN_IN), .ZN(n6925) );
  NAND4_X1 U7524 ( .A1(n6928), .A2(n6927), .A3(n6926), .A4(n6925), .ZN(U2814)
         );
  AOI22_X1 U7525 ( .A1(n6930), .A2(n6929), .B1(REIP_REG_14__SCAN_IN), .B2(
        n6943), .ZN(n6942) );
  INV_X1 U7526 ( .A(n6931), .ZN(n6932) );
  NAND3_X1 U7527 ( .A1(n6932), .A2(REIP_REG_12__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .ZN(n6935) );
  OAI22_X1 U7528 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6935), .B1(n6934), .B2(
        n6933), .ZN(n6936) );
  AOI211_X1 U7529 ( .C1(n6955), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6954), 
        .B(n6936), .ZN(n6941) );
  INV_X1 U7530 ( .A(n6937), .ZN(n6939) );
  AOI22_X1 U7531 ( .A1(n6939), .A2(n6978), .B1(n6938), .B2(n6950), .ZN(n6940)
         );
  NAND3_X1 U7532 ( .A1(n6942), .A2(n6941), .A3(n6940), .ZN(U2813) );
  AOI22_X1 U7533 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6972), .B1(
        REIP_REG_16__SCAN_IN), .B2(n6943), .ZN(n6947) );
  OAI211_X1 U7534 ( .C1(REIP_REG_15__SCAN_IN), .C2(REIP_REG_16__SCAN_IN), .A(
        n6945), .B(n6944), .ZN(n6946) );
  NAND2_X1 U7535 ( .A1(n6947), .A2(n6946), .ZN(n6948) );
  AOI211_X1 U7536 ( .C1(n6955), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6954), 
        .B(n6948), .ZN(n6952) );
  AOI22_X1 U7537 ( .A1(n7087), .A2(n6978), .B1(n6950), .B2(n6949), .ZN(n6951)
         );
  OAI211_X1 U7538 ( .C1(n6975), .C2(n6953), .A(n6952), .B(n6951), .ZN(U2811)
         );
  AOI21_X1 U7539 ( .B1(n6955), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6954), 
        .ZN(n6956) );
  OAI221_X1 U7540 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6968), .C1(n6958), .C2(
        n6957), .A(n6956), .ZN(n6964) );
  INV_X1 U7541 ( .A(n6959), .ZN(n6960) );
  OAI22_X1 U7542 ( .A1(n6962), .A2(n6961), .B1(n6975), .B2(n6960), .ZN(n6963)
         );
  AOI211_X1 U7543 ( .C1(EBX_REG_18__SCAN_IN), .C2(n6972), .A(n6964), .B(n6963), 
        .ZN(n6965) );
  OAI21_X1 U7544 ( .B1(n6966), .B2(n6973), .A(n6965), .ZN(U2809) );
  OAI21_X1 U7545 ( .B1(n6969), .B2(n6968), .A(n6967), .ZN(n6970) );
  AOI22_X1 U7546 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6972), .B1(n6971), .B2(n6970), .ZN(n6980) );
  OAI22_X1 U7547 ( .A1(n6976), .A2(n6975), .B1(n6974), .B2(n6973), .ZN(n6977)
         );
  AOI21_X1 U7548 ( .B1(n7095), .B2(n6978), .A(n6977), .ZN(n6979) );
  OAI211_X1 U7549 ( .C1(n4230), .C2(n6981), .A(n6980), .B(n6979), .ZN(U2807)
         );
  INV_X1 U7550 ( .A(n6982), .ZN(n6987) );
  NAND2_X1 U7551 ( .A1(n6983), .A2(n4672), .ZN(n6985) );
  AOI22_X1 U7552 ( .A1(n6988), .A2(n6985), .B1(n3438), .B2(n6984), .ZN(n6986)
         );
  OAI21_X1 U7553 ( .B1(n6988), .B2(n6987), .A(n6986), .ZN(n7019) );
  INV_X1 U7554 ( .A(n6989), .ZN(n6991) );
  NAND2_X1 U7555 ( .A1(n6991), .A2(n6990), .ZN(n7026) );
  AND2_X1 U7556 ( .A1(n6992), .A2(n7026), .ZN(n6994) );
  MUX2_X1 U7557 ( .A(MORE_REG_SCAN_IN), .B(n7019), .S(n6994), .Z(U3471) );
  OAI21_X1 U7558 ( .B1(n6994), .B2(n7024), .A(n6993), .ZN(U2793) );
  INV_X1 U7559 ( .A(n6995), .ZN(n6999) );
  NAND3_X1 U7560 ( .A1(n6997), .A2(n4629), .A3(n6996), .ZN(n6998) );
  OAI21_X1 U7561 ( .B1(n6999), .B2(n4352), .A(n6998), .ZN(U3455) );
  INV_X1 U7562 ( .A(n7010), .ZN(n7013) );
  AOI21_X1 U7563 ( .B1(n7000), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n7123), 
        .ZN(n7001) );
  AND2_X1 U7564 ( .A1(n7002), .A2(n7001), .ZN(n7005) );
  INV_X1 U7565 ( .A(n7005), .ZN(n7007) );
  AOI211_X1 U7566 ( .C1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n7005), .A(n7004), .B(n7003), .ZN(n7006) );
  AOI21_X1 U7567 ( .B1(n7008), .B2(n7007), .A(n7006), .ZN(n7009) );
  OAI21_X1 U7568 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n7010), .A(n7009), 
        .ZN(n7011) );
  OAI21_X1 U7569 ( .B1(n7013), .B2(n7012), .A(n7011), .ZN(n7018) );
  INV_X1 U7570 ( .A(n7014), .ZN(n7016) );
  OR2_X1 U7571 ( .A1(n7018), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n7015)
         );
  AND2_X1 U7572 ( .A1(n7016), .A2(n7015), .ZN(n7017) );
  AOI211_X1 U7573 ( .C1(n7018), .C2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n7017), .ZN(n7022) );
  NOR4_X1 U7574 ( .A1(n7022), .A2(n7021), .A3(n7020), .A4(n7019), .ZN(n7023)
         );
  OAI221_X1 U7575 ( .B1(n7026), .B2(n7025), .C1(n7026), .C2(n7024), .A(n7023), 
        .ZN(n7039) );
  OAI22_X1 U7576 ( .A1(n7039), .A2(n7051), .B1(n7028), .B2(n7027), .ZN(n7029)
         );
  OAI21_X1 U7577 ( .B1(n7031), .B2(n7030), .A(n7029), .ZN(n7045) );
  OAI21_X1 U7578 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n7028), .A(n7045), .ZN(
        n7044) );
  AOI21_X1 U7579 ( .B1(n7033), .B2(n7044), .A(n7032), .ZN(n7037) );
  OAI21_X1 U7580 ( .B1(READY_N), .B2(n7034), .A(n7051), .ZN(n7035) );
  NAND2_X1 U7581 ( .A1(n7045), .A2(n7035), .ZN(n7036) );
  OAI211_X1 U7582 ( .C1(n7040), .C2(n7045), .A(n7037), .B(n7036), .ZN(U3149)
         );
  OAI221_X1 U7583 ( .B1(n4629), .B2(STATE2_REG_0__SCAN_IN), .C1(n4629), .C2(
        n7045), .A(n7038), .ZN(U3453) );
  INV_X1 U7584 ( .A(n7039), .ZN(n7052) );
  INV_X1 U7585 ( .A(n7040), .ZN(n7041) );
  AND2_X1 U7586 ( .A1(n7042), .A2(n7041), .ZN(n7055) );
  AOI221_X1 U7587 ( .B1(n7055), .B2(STATE2_REG_0__SCAN_IN), .C1(n7044), .C2(
        STATE2_REG_0__SCAN_IN), .A(n7043), .ZN(n7050) );
  OAI211_X1 U7588 ( .C1(n7048), .C2(n7047), .A(n7046), .B(n7045), .ZN(n7049)
         );
  OAI211_X1 U7589 ( .C1(n7052), .C2(n7051), .A(n7050), .B(n7049), .ZN(U3148)
         );
  INV_X1 U7590 ( .A(n7053), .ZN(n7054) );
  AOI22_X1 U7591 ( .A1(n7061), .A2(n7055), .B1(n3443), .B2(n7054), .ZN(n7056)
         );
  OAI21_X1 U7592 ( .B1(n7058), .B2(n7057), .A(n7056), .ZN(n7059) );
  INV_X1 U7593 ( .A(n7059), .ZN(n7060) );
  OAI21_X1 U7594 ( .B1(n7123), .B2(n7061), .A(n7060), .ZN(U3465) );
  AOI21_X1 U7595 ( .B1(n7064), .B2(STATEBS16_REG_SCAN_IN), .A(n7063), .ZN(
        n7062) );
  INV_X1 U7596 ( .A(n7062), .ZN(U2792) );
  AOI21_X1 U7597 ( .B1(n7064), .B2(DATAWIDTH_REG_1__SCAN_IN), .A(n7063), .ZN(
        n7065) );
  INV_X1 U7598 ( .A(n7065), .ZN(U3452) );
  NAND2_X1 U7599 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n7070) );
  INV_X1 U7600 ( .A(n7079), .ZN(n7068) );
  INV_X1 U7601 ( .A(NA_N), .ZN(n7077) );
  AOI221_X1 U7602 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7077), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7081) );
  AOI221_X1 U7603 ( .B1(n7068), .B2(n7067), .C1(n7066), .C2(n7067), .A(n7081), 
        .ZN(n7069) );
  OAI221_X1 U7604 ( .B1(n7083), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n7083), 
        .C2(n7070), .A(n7069), .ZN(U3181) );
  AOI21_X1 U7605 ( .B1(READY_N), .B2(n7077), .A(n7071), .ZN(n7073) );
  AOI211_X1 U7606 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n7074), .A(n7073), 
        .B(n7072), .ZN(n7076) );
  NOR2_X1 U7607 ( .A1(n7076), .A2(n7075), .ZN(n7082) );
  AOI21_X1 U7608 ( .B1(n7078), .B2(n7077), .A(STATE_REG_2__SCAN_IN), .ZN(n7080) );
  OAI22_X1 U7609 ( .A1(n7082), .A2(n7081), .B1(n7080), .B2(n7079), .ZN(U3183)
         );
  OAI22_X1 U7610 ( .A1(n7084), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        M_IO_N_REG_SCAN_IN), .B2(n7083), .ZN(n7085) );
  INV_X1 U7611 ( .A(n7085), .ZN(U3473) );
  INV_X1 U7612 ( .A(n7086), .ZN(n7094) );
  AOI22_X1 U7613 ( .A1(n7087), .A2(n7094), .B1(n7093), .B2(DATAI_16_), .ZN(
        n7089) );
  AOI22_X1 U7614 ( .A1(n7097), .A2(DATAI_0_), .B1(n7096), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n7088) );
  NAND2_X1 U7615 ( .A1(n7089), .A2(n7088), .ZN(U2875) );
  AOI22_X1 U7616 ( .A1(n7090), .A2(n7094), .B1(n7093), .B2(DATAI_18_), .ZN(
        n7092) );
  AOI22_X1 U7617 ( .A1(n7097), .A2(DATAI_2_), .B1(n7096), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n7091) );
  NAND2_X1 U7618 ( .A1(n7092), .A2(n7091), .ZN(U2873) );
  AOI22_X1 U7619 ( .A1(n7095), .A2(n7094), .B1(n7093), .B2(DATAI_20_), .ZN(
        n7099) );
  AOI22_X1 U7620 ( .A1(n7097), .A2(DATAI_4_), .B1(n7096), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n7098) );
  NAND2_X1 U7621 ( .A1(n7099), .A2(n7098), .ZN(U2871) );
  NOR2_X1 U7622 ( .A1(n7100), .A2(n7139), .ZN(n7106) );
  NOR2_X1 U7623 ( .A1(n7123), .A2(n7104), .ZN(n7244) );
  AOI21_X1 U7624 ( .B1(n7124), .B2(n7101), .A(n7244), .ZN(n7105) );
  INV_X1 U7625 ( .A(n7105), .ZN(n7102) );
  AOI22_X1 U7626 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7103), .B1(n7106), .B2(
        n7102), .ZN(n7249) );
  AOI22_X1 U7627 ( .A1(n7146), .A2(n7244), .B1(n7153), .B2(n7243), .ZN(n7110)
         );
  AOI22_X1 U7628 ( .A1(n7106), .A2(n7105), .B1(n7139), .B2(n7104), .ZN(n7107)
         );
  NAND2_X1 U7629 ( .A1(n7149), .A2(n7107), .ZN(n7246) );
  AOI22_X1 U7630 ( .A1(n7246), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n7145), 
        .B2(n7245), .ZN(n7109) );
  OAI211_X1 U7631 ( .C1(n7249), .C2(n7156), .A(n7110), .B(n7109), .ZN(U3124)
         );
  INV_X1 U7632 ( .A(n7111), .ZN(n7112) );
  AOI21_X1 U7633 ( .B1(n7112), .B2(n3445), .A(n7139), .ZN(n7118) );
  NOR2_X1 U7634 ( .A1(n7123), .A2(n7113), .ZN(n7253) );
  AOI21_X1 U7635 ( .B1(n7114), .B2(n3443), .A(n7253), .ZN(n7117) );
  INV_X1 U7636 ( .A(n7117), .ZN(n7115) );
  AOI22_X1 U7637 ( .A1(n7118), .A2(n7115), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7120), .ZN(n7258) );
  NOR2_X1 U7638 ( .A1(n7251), .A2(n7130), .ZN(n7116) );
  AOI21_X1 U7639 ( .B1(n7146), .B2(n7253), .A(n7116), .ZN(n7122) );
  NAND2_X1 U7640 ( .A1(n7118), .A2(n7117), .ZN(n7119) );
  OAI211_X1 U7641 ( .C1(n7152), .C2(n7120), .A(n7119), .B(n7149), .ZN(n7255)
         );
  AOI22_X1 U7642 ( .A1(n7255), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n7145), 
        .B2(n7254), .ZN(n7121) );
  OAI211_X1 U7643 ( .C1(n7258), .C2(n7156), .A(n7122), .B(n7121), .ZN(U3108)
         );
  NOR2_X1 U7644 ( .A1(n7123), .A2(n7133), .ZN(n7260) );
  AOI21_X1 U7645 ( .B1(n7124), .B2(n3538), .A(n7260), .ZN(n7132) );
  INV_X1 U7646 ( .A(n7125), .ZN(n7127) );
  OAI21_X1 U7647 ( .B1(n7127), .B2(n7126), .A(n7152), .ZN(n7136) );
  OAI22_X1 U7648 ( .A1(n7128), .A2(n7133), .B1(n7132), .B2(n7136), .ZN(n7129)
         );
  NOR2_X1 U7649 ( .A1(n7233), .A2(n7130), .ZN(n7131) );
  AOI21_X1 U7650 ( .B1(n7146), .B2(n7260), .A(n7131), .ZN(n7138) );
  INV_X1 U7651 ( .A(n7132), .ZN(n7135) );
  NAND2_X1 U7652 ( .A1(n7139), .A2(n7133), .ZN(n7134) );
  OAI211_X1 U7653 ( .C1(n7136), .C2(n7135), .A(n7149), .B(n7134), .ZN(n7262)
         );
  AOI22_X1 U7654 ( .A1(n7262), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n7145), 
        .B2(n7259), .ZN(n7137) );
  OAI211_X1 U7655 ( .C1(n7265), .C2(n7156), .A(n7138), .B(n7137), .ZN(U3092)
         );
  NOR2_X1 U7656 ( .A1(n7140), .A2(n7139), .ZN(n7148) );
  INV_X1 U7657 ( .A(n7141), .ZN(n7268) );
  AOI21_X1 U7658 ( .B1(n7143), .B2(n7142), .A(n7268), .ZN(n7147) );
  INV_X1 U7659 ( .A(n7147), .ZN(n7144) );
  AOI22_X1 U7660 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7151), .B1(n7148), .B2(
        n7144), .ZN(n7276) );
  AOI22_X1 U7661 ( .A1(n7146), .A2(n7268), .B1(n7145), .B2(n7266), .ZN(n7155)
         );
  NAND2_X1 U7662 ( .A1(n7148), .A2(n7147), .ZN(n7150) );
  OAI211_X1 U7663 ( .C1(n7152), .C2(n7151), .A(n7150), .B(n7149), .ZN(n7272)
         );
  AOI22_X1 U7664 ( .A1(n7272), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n7153), 
        .B2(n7270), .ZN(n7154) );
  OAI211_X1 U7665 ( .C1(n7276), .C2(n7156), .A(n7155), .B(n7154), .ZN(U3076)
         );
  AOI22_X1 U7666 ( .A1(n7166), .A2(n7244), .B1(n7167), .B2(n7243), .ZN(n7158)
         );
  AOI22_X1 U7667 ( .A1(n7246), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n7165), 
        .B2(n7245), .ZN(n7157) );
  OAI211_X1 U7668 ( .C1(n7249), .C2(n7170), .A(n7158), .B(n7157), .ZN(U3125)
         );
  AOI22_X1 U7669 ( .A1(n7166), .A2(n7253), .B1(n7165), .B2(n7254), .ZN(n7160)
         );
  INV_X1 U7670 ( .A(n7251), .ZN(n7229) );
  AOI22_X1 U7671 ( .A1(n7255), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n7167), 
        .B2(n7229), .ZN(n7159) );
  OAI211_X1 U7672 ( .C1(n7258), .C2(n7170), .A(n7160), .B(n7159), .ZN(U3109)
         );
  NOR2_X1 U7673 ( .A1(n7233), .A2(n7161), .ZN(n7162) );
  AOI21_X1 U7674 ( .B1(n7166), .B2(n7260), .A(n7162), .ZN(n7164) );
  AOI22_X1 U7675 ( .A1(n7262), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n7165), 
        .B2(n7259), .ZN(n7163) );
  OAI211_X1 U7676 ( .C1(n7265), .C2(n7170), .A(n7164), .B(n7163), .ZN(U3093)
         );
  AOI22_X1 U7677 ( .A1(n7166), .A2(n7268), .B1(n7165), .B2(n7266), .ZN(n7169)
         );
  AOI22_X1 U7678 ( .A1(n7272), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n7167), 
        .B2(n7270), .ZN(n7168) );
  OAI211_X1 U7679 ( .C1(n7276), .C2(n7170), .A(n7169), .B(n7168), .ZN(U3077)
         );
  AOI22_X1 U7680 ( .A1(n7181), .A2(n7244), .B1(n7180), .B2(n7243), .ZN(n7172)
         );
  AOI22_X1 U7681 ( .A1(n7246), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n7182), 
        .B2(n7245), .ZN(n7171) );
  OAI211_X1 U7682 ( .C1(n7249), .C2(n7185), .A(n7172), .B(n7171), .ZN(U3126)
         );
  NOR2_X1 U7683 ( .A1(n7251), .A2(n7176), .ZN(n7173) );
  AOI21_X1 U7684 ( .B1(n7181), .B2(n7253), .A(n7173), .ZN(n7175) );
  AOI22_X1 U7685 ( .A1(n7255), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n7182), 
        .B2(n7254), .ZN(n7174) );
  OAI211_X1 U7686 ( .C1(n7258), .C2(n7185), .A(n7175), .B(n7174), .ZN(U3110)
         );
  NOR2_X1 U7687 ( .A1(n7233), .A2(n7176), .ZN(n7177) );
  AOI21_X1 U7688 ( .B1(n7181), .B2(n7260), .A(n7177), .ZN(n7179) );
  AOI22_X1 U7689 ( .A1(n7262), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n7182), 
        .B2(n7259), .ZN(n7178) );
  OAI211_X1 U7690 ( .C1(n7265), .C2(n7185), .A(n7179), .B(n7178), .ZN(U3094)
         );
  AOI22_X1 U7691 ( .A1(n7181), .A2(n7268), .B1(n7180), .B2(n7270), .ZN(n7184)
         );
  AOI22_X1 U7692 ( .A1(n7272), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n7182), 
        .B2(n7266), .ZN(n7183) );
  OAI211_X1 U7693 ( .C1(n7276), .C2(n7185), .A(n7184), .B(n7183), .ZN(U3078)
         );
  AOI22_X1 U7694 ( .A1(n7195), .A2(n7244), .B1(n7194), .B2(n7245), .ZN(n7187)
         );
  AOI22_X1 U7695 ( .A1(n7246), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n7196), 
        .B2(n7243), .ZN(n7186) );
  OAI211_X1 U7696 ( .C1(n7249), .C2(n7199), .A(n7187), .B(n7186), .ZN(U3127)
         );
  AOI22_X1 U7697 ( .A1(n7195), .A2(n7253), .B1(n7194), .B2(n7254), .ZN(n7189)
         );
  AOI22_X1 U7698 ( .A1(n7255), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n7196), 
        .B2(n7229), .ZN(n7188) );
  OAI211_X1 U7699 ( .C1(n7258), .C2(n7199), .A(n7189), .B(n7188), .ZN(U3111)
         );
  NOR2_X1 U7700 ( .A1(n7233), .A2(n7190), .ZN(n7191) );
  AOI21_X1 U7701 ( .B1(n7195), .B2(n7260), .A(n7191), .ZN(n7193) );
  AOI22_X1 U7702 ( .A1(n7262), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n7194), 
        .B2(n7259), .ZN(n7192) );
  OAI211_X1 U7703 ( .C1(n7265), .C2(n7199), .A(n7193), .B(n7192), .ZN(U3095)
         );
  AOI22_X1 U7704 ( .A1(n7195), .A2(n7268), .B1(n7194), .B2(n7266), .ZN(n7198)
         );
  AOI22_X1 U7705 ( .A1(n7272), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n7196), 
        .B2(n7270), .ZN(n7197) );
  OAI211_X1 U7706 ( .C1(n7276), .C2(n7199), .A(n7198), .B(n7197), .ZN(U3079)
         );
  AOI22_X1 U7707 ( .A1(n7210), .A2(n7244), .B1(n7211), .B2(n7245), .ZN(n7201)
         );
  AOI22_X1 U7708 ( .A1(n7246), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n7209), 
        .B2(n7243), .ZN(n7200) );
  OAI211_X1 U7709 ( .C1(n7249), .C2(n7214), .A(n7201), .B(n7200), .ZN(U3128)
         );
  NOR2_X1 U7710 ( .A1(n7251), .A2(n7205), .ZN(n7202) );
  AOI21_X1 U7711 ( .B1(n7210), .B2(n7253), .A(n7202), .ZN(n7204) );
  AOI22_X1 U7712 ( .A1(n7255), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n7211), 
        .B2(n7254), .ZN(n7203) );
  OAI211_X1 U7713 ( .C1(n7258), .C2(n7214), .A(n7204), .B(n7203), .ZN(U3112)
         );
  NOR2_X1 U7714 ( .A1(n7233), .A2(n7205), .ZN(n7206) );
  AOI21_X1 U7715 ( .B1(n7210), .B2(n7260), .A(n7206), .ZN(n7208) );
  AOI22_X1 U7716 ( .A1(n7262), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n7211), 
        .B2(n7259), .ZN(n7207) );
  OAI211_X1 U7717 ( .C1(n7265), .C2(n7214), .A(n7208), .B(n7207), .ZN(U3096)
         );
  AOI22_X1 U7718 ( .A1(n7210), .A2(n7268), .B1(n7209), .B2(n7270), .ZN(n7213)
         );
  AOI22_X1 U7719 ( .A1(n7272), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n7211), 
        .B2(n7266), .ZN(n7212) );
  OAI211_X1 U7720 ( .C1(n7276), .C2(n7214), .A(n7213), .B(n7212), .ZN(U3080)
         );
  AOI22_X1 U7721 ( .A1(n7222), .A2(n7244), .B1(n7221), .B2(n7243), .ZN(n7216)
         );
  AOI22_X1 U7722 ( .A1(n7246), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n7223), 
        .B2(n7245), .ZN(n7215) );
  OAI211_X1 U7723 ( .C1(n7249), .C2(n7226), .A(n7216), .B(n7215), .ZN(U3129)
         );
  AOI22_X1 U7724 ( .A1(n7222), .A2(n7253), .B1(n7223), .B2(n7254), .ZN(n7218)
         );
  AOI22_X1 U7725 ( .A1(n7255), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n7221), 
        .B2(n7229), .ZN(n7217) );
  OAI211_X1 U7726 ( .C1(n7258), .C2(n7226), .A(n7218), .B(n7217), .ZN(U3113)
         );
  AOI22_X1 U7727 ( .A1(n7222), .A2(n7260), .B1(n7223), .B2(n7259), .ZN(n7220)
         );
  INV_X1 U7728 ( .A(n7233), .ZN(n7261) );
  AOI22_X1 U7729 ( .A1(n7262), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n7221), 
        .B2(n7261), .ZN(n7219) );
  OAI211_X1 U7730 ( .C1(n7265), .C2(n7226), .A(n7220), .B(n7219), .ZN(U3097)
         );
  AOI22_X1 U7731 ( .A1(n7222), .A2(n7268), .B1(n7221), .B2(n7270), .ZN(n7225)
         );
  AOI22_X1 U7732 ( .A1(n7272), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n7223), 
        .B2(n7266), .ZN(n7224) );
  OAI211_X1 U7733 ( .C1(n7276), .C2(n7226), .A(n7225), .B(n7224), .ZN(U3081)
         );
  AOI22_X1 U7734 ( .A1(n7238), .A2(n7244), .B1(n7239), .B2(n7245), .ZN(n7228)
         );
  AOI22_X1 U7735 ( .A1(n7246), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n7237), 
        .B2(n7243), .ZN(n7227) );
  OAI211_X1 U7736 ( .C1(n7249), .C2(n7242), .A(n7228), .B(n7227), .ZN(U3130)
         );
  AOI22_X1 U7737 ( .A1(n7238), .A2(n7253), .B1(n7239), .B2(n7254), .ZN(n7231)
         );
  AOI22_X1 U7738 ( .A1(n7255), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n7237), 
        .B2(n7229), .ZN(n7230) );
  OAI211_X1 U7739 ( .C1(n7258), .C2(n7242), .A(n7231), .B(n7230), .ZN(U3114)
         );
  NOR2_X1 U7740 ( .A1(n7233), .A2(n7232), .ZN(n7234) );
  AOI21_X1 U7741 ( .B1(n7238), .B2(n7260), .A(n7234), .ZN(n7236) );
  AOI22_X1 U7742 ( .A1(n7262), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n7239), 
        .B2(n7259), .ZN(n7235) );
  OAI211_X1 U7743 ( .C1(n7265), .C2(n7242), .A(n7236), .B(n7235), .ZN(U3098)
         );
  AOI22_X1 U7744 ( .A1(n7238), .A2(n7268), .B1(n7237), .B2(n7270), .ZN(n7241)
         );
  AOI22_X1 U7745 ( .A1(n7272), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n7239), 
        .B2(n7266), .ZN(n7240) );
  OAI211_X1 U7746 ( .C1(n7276), .C2(n7242), .A(n7241), .B(n7240), .ZN(U3082)
         );
  AOI22_X1 U7747 ( .A1(n7269), .A2(n7244), .B1(n7271), .B2(n7243), .ZN(n7248)
         );
  AOI22_X1 U7748 ( .A1(n7246), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n7267), 
        .B2(n7245), .ZN(n7247) );
  OAI211_X1 U7749 ( .C1(n7249), .C2(n7275), .A(n7248), .B(n7247), .ZN(U3131)
         );
  NOR2_X1 U7750 ( .A1(n7251), .A2(n7250), .ZN(n7252) );
  AOI21_X1 U7751 ( .B1(n7269), .B2(n7253), .A(n7252), .ZN(n7257) );
  AOI22_X1 U7752 ( .A1(n7255), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n7267), 
        .B2(n7254), .ZN(n7256) );
  OAI211_X1 U7753 ( .C1(n7258), .C2(n7275), .A(n7257), .B(n7256), .ZN(U3115)
         );
  AOI22_X1 U7754 ( .A1(n7269), .A2(n7260), .B1(n7267), .B2(n7259), .ZN(n7264)
         );
  AOI22_X1 U7755 ( .A1(n7262), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n7271), 
        .B2(n7261), .ZN(n7263) );
  OAI211_X1 U7756 ( .C1(n7265), .C2(n7275), .A(n7264), .B(n7263), .ZN(U3099)
         );
  AOI22_X1 U7757 ( .A1(n7269), .A2(n7268), .B1(n7267), .B2(n7266), .ZN(n7274)
         );
  AOI22_X1 U7758 ( .A1(n7272), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n7271), 
        .B2(n7270), .ZN(n7273) );
  OAI211_X1 U7759 ( .C1(n7276), .C2(n7275), .A(n7274), .B(n7273), .ZN(U3083)
         );
  INV_X2 U3498 ( .A(n4603), .ZN(n6171) );
  CLKBUF_X1 U3487 ( .A(n3827), .Z(n3867) );
  CLKBUF_X1 U3491 ( .A(n3880), .Z(n3443) );
  AOI21_X1 U3505 ( .B1(n6078), .B2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n4688), 
        .ZN(n4694) );
  CLKBUF_X1 U3506 ( .A(n4713), .Z(n3438) );
  CLKBUF_X1 U3842 ( .A(n5230), .Z(n5274) );
  CLKBUF_X1 U4033 ( .A(n6186), .Z(n6189) );
  INV_X2 U4125 ( .A(n7027), .ZN(n6741) );
  CLKBUF_X1 U4353 ( .A(n3734), .Z(n3931) );
endmodule

