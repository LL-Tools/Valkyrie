

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047,
         n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057,
         n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067,
         n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077,
         n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087,
         n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097,
         n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107,
         n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
         n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127,
         n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137,
         n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147,
         n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157,
         n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167,
         n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177,
         n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187,
         n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197,
         n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207,
         n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217,
         n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227,
         n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237,
         n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247,
         n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257,
         n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267,
         n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277,
         n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
         n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
         n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
         n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
         n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
         n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
         n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
         n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
         n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
         n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397,
         n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407,
         n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417,
         n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427,
         n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
         n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447,
         n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457,
         n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
         n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
         n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
         n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
         n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507,
         n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517,
         n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527,
         n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537,
         n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557,
         n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567,
         n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577,
         n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587,
         n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597,
         n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607,
         n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617,
         n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627,
         n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637,
         n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647,
         n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657,
         n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667,
         n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677,
         n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687,
         n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697,
         n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707,
         n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717,
         n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727,
         n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737,
         n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747,
         n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757,
         n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777,
         n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787,
         n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797,
         n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807,
         n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837,
         n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847,
         n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054;

  INV_X4 U5093 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  OAI21_X1 U5094 ( .B1(n6400), .B2(n5211), .A(n5209), .ZN(n6412) );
  NAND2_X1 U5095 ( .A1(n8445), .A2(n5169), .ZN(n10308) );
  NAND2_X1 U5096 ( .A1(n5879), .A2(n5878), .ZN(n10863) );
  XNOR2_X1 U5097 ( .A(n5226), .B(n5225), .ZN(n10229) );
  NAND4_X2 U5098 ( .A1(n6865), .A2(n6863), .A3(n5661), .A4(n6864), .ZN(n7107)
         );
  CLKBUF_X2 U5099 ( .A(n5800), .Z(n8030) );
  NAND2_X2 U5100 ( .A1(n6482), .A2(n6481), .ZN(n10512) );
  INV_X1 U5101 ( .A(n8186), .ZN(n8155) );
  INV_X1 U5102 ( .A(n5825), .ZN(n6072) );
  INV_X4 U5103 ( .A(n9187), .ZN(n9181) );
  BUF_X1 U5104 ( .A(n7058), .Z(n5030) );
  INV_X1 U5105 ( .A(n6634), .ZN(n6583) );
  INV_X2 U5106 ( .A(n6350), .ZN(n6696) );
  INV_X1 U5107 ( .A(n6252), .ZN(n8029) );
  INV_X1 U5108 ( .A(n9182), .ZN(n8396) );
  OR2_X1 U5109 ( .A1(n9592), .A2(n10229), .ZN(n5309) );
  INV_X1 U5110 ( .A(n7016), .ZN(n7753) );
  AND2_X1 U5111 ( .A1(n8518), .A2(n10447), .ZN(n7712) );
  OR2_X1 U5112 ( .A1(n10909), .A2(n7773), .ZN(n7789) );
  NAND2_X1 U5113 ( .A1(n9402), .A2(n9404), .ZN(n7290) );
  INV_X1 U5114 ( .A(n6223), .ZN(n10815) );
  NAND2_X1 U5115 ( .A1(n7822), .A2(n7821), .ZN(n10398) );
  NAND2_X2 U5116 ( .A1(n10512), .A2(n10510), .ZN(n6895) );
  OAI22_X1 U5117 ( .A1(n10308), .A2(n8446), .B1(n9533), .B2(n11022), .ZN(
        n10283) );
  AND2_X1 U5118 ( .A1(n6498), .A2(n6497), .ZN(n9595) );
  INV_X1 U5119 ( .A(n8665), .ZN(P2_U3966) );
  INV_X2 U5120 ( .A(n10942), .ZN(n10296) );
  INV_X2 U5121 ( .A(n6692), .ZN(n6675) );
  AND2_X2 U5122 ( .A1(n5214), .A2(n6508), .ZN(n6510) );
  BUF_X2 U5123 ( .A(n6227), .Z(n5028) );
  AND2_X1 U5124 ( .A1(n5772), .A2(n9138), .ZN(n5800) );
  AND2_X1 U5125 ( .A1(n5772), .A2(n5771), .ZN(n5901) );
  INV_X2 U5126 ( .A(n5772), .ZN(n8499) );
  NAND2_X1 U5127 ( .A1(n6895), .A2(n8021), .ZN(n5029) );
  OAI22_X2 U5128 ( .A1(n8831), .A2(n8835), .B1(n9052), .B2(n8655), .ZN(n8814)
         );
  AOI22_X2 U5129 ( .A1(n8846), .A2(n8852), .B1(n8851), .B2(n8861), .ZN(n8831)
         );
  AOI21_X1 U5130 ( .B1(n5322), .B2(n11024), .A(n5188), .ZN(n5187) );
  XNOR2_X1 U5131 ( .A(n6412), .B(n6410), .ZN(n8597) );
  NAND2_X1 U5132 ( .A1(n5477), .A2(n5063), .ZN(n8865) );
  INV_X1 U5133 ( .A(n5482), .ZN(n8892) );
  OAI21_X1 U5134 ( .B1(n8454), .B2(n5172), .A(n5170), .ZN(n5376) );
  NAND2_X1 U5135 ( .A1(n5609), .A2(n8296), .ZN(n9307) );
  NAND2_X1 U5136 ( .A1(n9308), .A2(n9306), .ZN(n9312) );
  OAI211_X1 U5137 ( .C1(n5460), .C2(n5464), .A(n5461), .B(n5459), .ZN(n10275)
         );
  NAND2_X1 U5138 ( .A1(n7870), .A2(n7869), .ZN(n8267) );
  OR2_X1 U5139 ( .A1(n7788), .A2(n9429), .ZN(n7786) );
  OR2_X1 U5140 ( .A1(n9109), .A2(n7942), .ZN(n8999) );
  OR2_X1 U5141 ( .A1(n9100), .A2(n8627), .ZN(n8123) );
  NAND2_X1 U5142 ( .A1(n7322), .A2(n7321), .ZN(n7320) );
  NAND2_X1 U5143 ( .A1(n10888), .A2(n6330), .ZN(n7322) );
  AOI21_X1 U5144 ( .B1(n10912), .B2(n7543), .A(n9326), .ZN(n7544) );
  NAND2_X1 U5145 ( .A1(n5976), .A2(n5975), .ZN(n8107) );
  NAND2_X1 U5146 ( .A1(n7086), .A2(n7087), .ZN(n7085) );
  NAND2_X1 U5147 ( .A1(n7967), .A2(n7966), .ZN(n10316) );
  NAND3_X1 U5148 ( .A1(n9021), .A2(n5896), .A3(n5880), .ZN(n5135) );
  NAND2_X1 U5149 ( .A1(n5918), .A2(n5917), .ZN(n10962) );
  NAND2_X1 U5150 ( .A1(n5965), .A2(n5964), .ZN(n7737) );
  NAND2_X2 U5151 ( .A1(n7159), .A2(n8987), .ZN(n10818) );
  XNOR2_X1 U5152 ( .A(n5911), .B(n5910), .ZN(n7522) );
  OR2_X1 U5153 ( .A1(n7413), .A2(n6128), .ZN(n5888) );
  NAND2_X1 U5154 ( .A1(n5871), .A2(n5146), .ZN(n7331) );
  INV_X1 U5155 ( .A(n7263), .ZN(n10784) );
  AND2_X1 U5156 ( .A1(n7021), .A2(n5667), .ZN(n7292) );
  NAND2_X1 U5157 ( .A1(n5836), .A2(n5057), .ZN(n8542) );
  AND4_X1 U5158 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(n6323)
         );
  INV_X4 U5159 ( .A(n8418), .ZN(n9185) );
  INV_X1 U5160 ( .A(n10766), .ZN(n6304) );
  NAND2_X2 U5161 ( .A1(n6462), .A2(n10621), .ZN(n8665) );
  OAI211_X1 U5162 ( .C1(n6895), .C2(n10016), .A(n7005), .B(n7004), .ZN(n7213)
         );
  OAI211_X1 U5163 ( .C1(n6634), .C2(n6776), .A(n5832), .B(n5831), .ZN(n10766)
         );
  NAND2_X2 U5164 ( .A1(n10923), .A2(n7111), .ZN(n8418) );
  NAND3_X1 U5165 ( .A1(n5213), .A2(n8237), .A3(n5212), .ZN(n6303) );
  AND3_X1 U5166 ( .A1(n6899), .A2(n6897), .A3(n6898), .ZN(n10713) );
  NOR2_X2 U5167 ( .A1(n8382), .A2(n6894), .ZN(n9182) );
  NAND3_X1 U5168 ( .A1(n6891), .A2(n6890), .A3(n7124), .ZN(n10923) );
  NAND4_X1 U5169 ( .A1(n5792), .A2(n5789), .A3(n5790), .A4(n5791), .ZN(n7469)
         );
  CLKBUF_X1 U5170 ( .A(n5035), .Z(n8412) );
  INV_X1 U5171 ( .A(n7108), .ZN(n10712) );
  OR2_X2 U5172 ( .A1(n6223), .A2(n8035), .ZN(n8186) );
  BUF_X2 U5173 ( .A(n7712), .Z(n5035) );
  AND2_X1 U5174 ( .A1(n5695), .A2(n5869), .ZN(n5696) );
  AND2_X1 U5175 ( .A1(n5664), .A2(n5872), .ZN(n5693) );
  INV_X1 U5176 ( .A(n5771), .ZN(n9138) );
  OR2_X1 U5177 ( .A1(n5694), .A2(n5867), .ZN(n5869) );
  XNOR2_X1 U5178 ( .A(n5144), .B(n5768), .ZN(n5772) );
  XNOR2_X1 U5179 ( .A(n5653), .B(n6601), .ZN(n8518) );
  XNOR2_X1 U5180 ( .A(n5770), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U5181 ( .A1(n5769), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5770) );
  AND2_X1 U5182 ( .A1(n5165), .A2(n5685), .ZN(n5844) );
  OR2_X1 U5183 ( .A1(n10438), .A2(n10439), .ZN(n5653) );
  XNOR2_X1 U5184 ( .A(n6604), .B(n6603), .ZN(n10447) );
  NAND2_X1 U5185 ( .A1(n6477), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n6482) );
  XNOR2_X1 U5186 ( .A(n5762), .B(n5761), .ZN(n6253) );
  OR2_X1 U5187 ( .A1(n5763), .A2(n5354), .ZN(n5353) );
  NAND2_X1 U5188 ( .A1(n5766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5762) );
  BUF_X4 U5189 ( .A(n6507), .Z(n6881) );
  OR2_X1 U5190 ( .A1(n5903), .A2(n5902), .ZN(n5920) );
  AND2_X1 U5191 ( .A1(n5760), .A2(n5607), .ZN(n5606) );
  INV_X2 U5192 ( .A(n8021), .ZN(n6507) );
  AND2_X1 U5193 ( .A1(n6271), .A2(n5759), .ZN(n5760) );
  AND3_X1 U5194 ( .A1(n5152), .A2(n6274), .A3(n6278), .ZN(n6271) );
  AND2_X1 U5195 ( .A1(n5471), .A2(n6474), .ZN(n5470) );
  INV_X1 U5196 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6016) );
  INV_X1 U5197 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5961) );
  INV_X1 U5198 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5960) );
  NOR2_X1 U5199 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5752) );
  INV_X1 U5200 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6495) );
  NOR2_X1 U5201 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5757) );
  INV_X1 U5202 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6831) );
  INV_X4 U5203 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5204 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n6537) );
  INV_X1 U5205 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5122) );
  INV_X1 U5206 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5124) );
  INV_X1 U5207 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5123) );
  NOR2_X1 U5208 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5355) );
  NOR2_X2 U5209 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5564) );
  OAI211_X1 U5210 ( .C1(n5346), .C2(n5345), .A(n8092), .B(n8093), .ZN(n5344)
         );
  NOR2_X2 U5211 ( .A1(n7466), .A2(n10766), .ZN(n7260) );
  OAI21_X2 U5212 ( .B1(n5911), .B2(n5711), .A(n5710), .ZN(n5929) );
  NOR3_X2 U5213 ( .A1(n7789), .A2(n10398), .A3(n5326), .ZN(n5324) );
  NAND2_X1 U5214 ( .A1(n6607), .A2(n6605), .ZN(n5031) );
  NAND2_X2 U5215 ( .A1(n6607), .A2(n6605), .ZN(n5032) );
  INV_X1 U5216 ( .A(n5032), .ZN(n5033) );
  NAND2_X1 U5217 ( .A1(n6607), .A2(n6605), .ZN(n8432) );
  NAND4_X2 U5218 ( .A1(n6880), .A2(n6879), .A3(n6878), .A4(n6877), .ZN(n6949)
         );
  BUF_X4 U5219 ( .A(n7017), .Z(n5034) );
  NAND2_X1 U5220 ( .A1(n6605), .A2(n8518), .ZN(n7017) );
  AND2_X1 U5221 ( .A1(n8995), .A2(n8117), .ZN(n8118) );
  NAND2_X1 U5222 ( .A1(n8166), .A2(n8186), .ZN(n5539) );
  OR2_X1 U5223 ( .A1(n10323), .A2(n9467), .ZN(n9388) );
  AND2_X1 U5224 ( .A1(n5509), .A2(n5203), .ZN(n5202) );
  NAND2_X1 U5225 ( .A1(n5511), .A2(n5204), .ZN(n5203) );
  AOI21_X1 U5226 ( .B1(n5511), .B2(n5513), .A(n5061), .ZN(n5509) );
  INV_X1 U5227 ( .A(n6418), .ZN(n5204) );
  INV_X1 U5228 ( .A(n7924), .ZN(n5984) );
  NOR2_X1 U5229 ( .A1(n5897), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5962) );
  AND2_X1 U5230 ( .A1(n6464), .A2(n6463), .ZN(n5215) );
  INV_X1 U5231 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U5232 ( .A1(n6889), .A2(n7502), .ZN(n7124) );
  NAND2_X1 U5233 ( .A1(n8126), .A2(n8125), .ZN(n8133) );
  OR2_X1 U5234 ( .A1(n8172), .A2(n8155), .ZN(n5341) );
  INV_X1 U5235 ( .A(n8066), .ZN(n5486) );
  INV_X1 U5236 ( .A(SI_20_), .ZN(n5744) );
  INV_X1 U5237 ( .A(SI_19_), .ZN(n9627) );
  INV_X1 U5238 ( .A(n5727), .ZN(n5289) );
  NAND2_X1 U5239 ( .A1(n5202), .A2(n5199), .ZN(n5198) );
  NAND2_X1 U5240 ( .A1(n5205), .A2(n5200), .ZN(n5199) );
  NOR2_X1 U5241 ( .A1(n9057), .A2(n9062), .ZN(n5272) );
  INV_X1 U5242 ( .A(n8859), .ZN(n6247) );
  OR2_X1 U5243 ( .A1(n9079), .A2(n8934), .ZN(n8144) );
  OR2_X1 U5244 ( .A1(n7908), .A2(n8646), .ZN(n8112) );
  OR2_X1 U5245 ( .A1(n7737), .A2(n7915), .ZN(n8097) );
  AND2_X1 U5246 ( .A1(n5153), .A2(n5909), .ZN(n5134) );
  NAND2_X1 U5247 ( .A1(n5052), .A2(n5752), .ZN(n5141) );
  NAND2_X1 U5248 ( .A1(n5521), .A2(n5520), .ZN(n5519) );
  INV_X1 U5249 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5520) );
  INV_X1 U5250 ( .A(n5522), .ZN(n5521) );
  NAND2_X1 U5251 ( .A1(n8352), .A2(n9250), .ZN(n5645) );
  AND2_X1 U5252 ( .A1(n7223), .A2(n7224), .ZN(n7232) );
  OR2_X1 U5253 ( .A1(n6911), .A2(n6887), .ZN(n8382) );
  NOR2_X1 U5254 ( .A1(n9582), .A2(n5298), .ZN(n5297) );
  AOI21_X1 U5255 ( .B1(n5173), .B2(n5171), .A(n5380), .ZN(n5170) );
  INV_X1 U5256 ( .A(n5175), .ZN(n5171) );
  AND2_X1 U5257 ( .A1(n5388), .A2(n8456), .ZN(n5387) );
  NAND2_X1 U5258 ( .A1(n10191), .A2(n8455), .ZN(n5388) );
  AND2_X1 U5259 ( .A1(n5384), .A2(n5177), .ZN(n5173) );
  OR2_X1 U5260 ( .A1(n10378), .A2(n10251), .ZN(n9561) );
  OR2_X1 U5261 ( .A1(n10393), .A2(n10304), .ZN(n9546) );
  AND2_X1 U5262 ( .A1(n7492), .A2(n10229), .ZN(n6893) );
  NAND2_X1 U5263 ( .A1(n9422), .A2(n9388), .ZN(n9582) );
  AND2_X1 U5264 ( .A1(n6467), .A2(n5225), .ZN(n5652) );
  NAND2_X1 U5265 ( .A1(n8002), .A2(n8001), .ZN(n8018) );
  NAND2_X1 U5266 ( .A1(n6189), .A2(n6188), .ZN(n6200) );
  AOI21_X1 U5267 ( .B1(n5292), .B2(n5294), .A(n5555), .ZN(n5290) );
  INV_X1 U5268 ( .A(n5748), .ZN(n5747) );
  XNOR2_X1 U5269 ( .A(n5743), .B(n5744), .ZN(n6080) );
  INV_X1 U5270 ( .A(n5558), .ZN(n5281) );
  AOI21_X1 U5271 ( .B1(n5561), .B2(n5560), .A(n5559), .ZN(n5558) );
  INV_X1 U5272 ( .A(n5735), .ZN(n5559) );
  INV_X1 U5273 ( .A(n6012), .ZN(n5560) );
  NAND2_X1 U5274 ( .A1(n5734), .A2(SI_17_), .ZN(n5735) );
  INV_X1 U5275 ( .A(SI_16_), .ZN(n9625) );
  NAND2_X1 U5276 ( .A1(n5284), .A2(n5285), .ZN(n6013) );
  NAND2_X1 U5277 ( .A1(n5986), .A2(n5288), .ZN(n5284) );
  AOI21_X1 U5278 ( .B1(n5547), .B2(n5549), .A(n5546), .ZN(n5545) );
  INV_X1 U5279 ( .A(n5716), .ZN(n5546) );
  INV_X1 U5280 ( .A(n5928), .ZN(n5547) );
  INV_X1 U5281 ( .A(n5549), .ZN(n5548) );
  OR2_X1 U5282 ( .A1(n5709), .A2(n5708), .ZN(n5710) );
  OR2_X1 U5283 ( .A1(n5910), .A2(n5709), .ZN(n5711) );
  NAND2_X1 U5284 ( .A1(n5884), .A2(n5701), .ZN(n5911) );
  INV_X1 U5285 ( .A(n5793), .ZN(n6252) );
  OR2_X1 U5286 ( .A1(n9057), .A2(n8861), .ZN(n8833) );
  NAND2_X1 U5287 ( .A1(n9005), .A2(n5492), .ZN(n8975) );
  AND2_X1 U5288 ( .A1(n6045), .A2(n6031), .ZN(n5492) );
  NAND2_X1 U5289 ( .A1(n9007), .A2(n9006), .ZN(n9005) );
  NAND2_X1 U5290 ( .A1(n7731), .A2(n5972), .ZN(n7924) );
  INV_X1 U5291 ( .A(n6128), .ZN(n8036) );
  NAND2_X1 U5292 ( .A1(n5133), .A2(n5131), .ZN(n7401) );
  OR2_X1 U5293 ( .A1(n7373), .A2(n5132), .ZN(n5131) );
  NAND2_X1 U5294 ( .A1(n5135), .A2(n5134), .ZN(n5133) );
  INV_X1 U5295 ( .A(n5909), .ZN(n5132) );
  NOR2_X1 U5297 ( .A1(n9032), .A2(n9038), .ZN(n5261) );
  AND2_X1 U5298 ( .A1(n8240), .A2(n8189), .ZN(n10864) );
  NOR2_X1 U5299 ( .A1(n5974), .A2(n5523), .ZN(n6021) );
  AND4_X1 U5300 ( .A1(n8436), .A2(n8435), .A3(n8434), .A4(n8433), .ZN(n9188)
         );
  NAND2_X1 U5301 ( .A1(n10117), .A2(n10096), .ZN(n10090) );
  NOR2_X1 U5302 ( .A1(n8463), .A2(n5186), .ZN(n5185) );
  INV_X1 U5303 ( .A(n8461), .ZN(n5186) );
  AND2_X1 U5304 ( .A1(n5317), .A2(n5316), .ZN(n5315) );
  OAI21_X1 U5305 ( .B1(n10219), .B2(n8451), .A(n8452), .ZN(n10207) );
  AOI21_X1 U5306 ( .B1(n5360), .B2(n5362), .A(n5094), .ZN(n5358) );
  AND4_X1 U5307 ( .A1(n7769), .A2(n7768), .A3(n7767), .A4(n7766), .ZN(n10303)
         );
  INV_X1 U5308 ( .A(n5030), .ZN(n9390) );
  INV_X1 U5309 ( .A(n6893), .ZN(n7123) );
  INV_X1 U5310 ( .A(n10915), .ZN(n10843) );
  INV_X1 U5311 ( .A(n10917), .ZN(n10842) );
  INV_X1 U5312 ( .A(n9582), .ZN(n5368) );
  INV_X1 U5313 ( .A(n8500), .ZN(n8466) );
  NAND2_X1 U5314 ( .A1(n6465), .A2(n6516), .ZN(n6466) );
  INV_X1 U5315 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U5316 ( .A1(n5882), .A2(n5881), .ZN(n5884) );
  NAND2_X1 U5317 ( .A1(n5229), .A2(n5231), .ZN(n9192) );
  NAND2_X1 U5318 ( .A1(n5253), .A2(n5252), .ZN(n5251) );
  INV_X1 U5319 ( .A(n10082), .ZN(n5253) );
  NAND2_X1 U5320 ( .A1(n10664), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U5321 ( .A1(n10942), .A2(n7131), .ZN(n10300) );
  INV_X1 U5322 ( .A(n9628), .ZN(n5394) );
  AND2_X1 U5323 ( .A1(n5393), .A2(n5392), .ZN(n5391) );
  NAND2_X1 U5324 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_128), .ZN(n5393) );
  NAND2_X1 U5325 ( .A1(keyinput_129), .A2(SI_31_), .ZN(n5392) );
  NAND2_X1 U5326 ( .A1(n9631), .A2(keyinput_131), .ZN(n9634) );
  OAI21_X1 U5327 ( .B1(n9656), .B2(n5413), .A(n5410), .ZN(n5409) );
  AND2_X1 U5328 ( .A1(n5412), .A2(n5411), .ZN(n5410) );
  AND2_X1 U5329 ( .A1(n9657), .A2(keyinput_142), .ZN(n5413) );
  INV_X1 U5330 ( .A(n9660), .ZN(n5408) );
  XNOR2_X1 U5331 ( .A(SI_14_), .B(keyinput_146), .ZN(n5407) );
  AOI21_X1 U5332 ( .B1(n5416), .B2(n5415), .A(n5414), .ZN(n9685) );
  XNOR2_X1 U5333 ( .A(keyinput_160), .B(SI_0_), .ZN(n5414) );
  INV_X1 U5334 ( .A(n9676), .ZN(n5415) );
  OAI21_X1 U5335 ( .B1(n9667), .B2(n5418), .A(n5417), .ZN(n5416) );
  OAI21_X1 U5336 ( .B1(n5351), .B2(n8048), .A(n8155), .ZN(n5350) );
  NOR2_X1 U5337 ( .A1(n8195), .A2(n8049), .ZN(n5351) );
  NAND2_X1 U5338 ( .A1(n8050), .A2(n8186), .ZN(n5349) );
  OAI21_X1 U5339 ( .B1(n9741), .B2(n5430), .A(n5429), .ZN(n5428) );
  INV_X1 U5340 ( .A(n9742), .ZN(n5429) );
  INV_X1 U5341 ( .A(n5431), .ZN(n5430) );
  AND2_X1 U5342 ( .A1(n8161), .A2(n8160), .ZN(n5332) );
  INV_X1 U5343 ( .A(n5335), .ZN(n5334) );
  OAI21_X1 U5344 ( .B1(n8148), .B2(n8147), .A(n5336), .ZN(n5335) );
  INV_X1 U5345 ( .A(n5337), .ZN(n5333) );
  AND2_X1 U5346 ( .A1(n10191), .A2(n10206), .ZN(n5158) );
  NAND2_X1 U5347 ( .A1(n5404), .A2(n5402), .ZN(n9783) );
  XNOR2_X1 U5348 ( .A(n6830), .B(n5403), .ZN(n5402) );
  NAND2_X1 U5349 ( .A1(n5405), .A2(n9782), .ZN(n5404) );
  INV_X1 U5350 ( .A(keyinput_232), .ZN(n5403) );
  NAND2_X1 U5351 ( .A1(n5398), .A2(n9799), .ZN(n5397) );
  NAND2_X1 U5352 ( .A1(n5400), .A2(n5399), .ZN(n5398) );
  INV_X1 U5353 ( .A(n6429), .ZN(n5200) );
  INV_X1 U5354 ( .A(n8088), .ZN(n5603) );
  INV_X1 U5355 ( .A(n5602), .ZN(n5601) );
  OAI21_X1 U5356 ( .B1(n5049), .B2(n5603), .A(n8204), .ZN(n5602) );
  NOR2_X1 U5357 ( .A1(n9274), .A2(n5643), .ZN(n5642) );
  INV_X1 U5358 ( .A(n9203), .ZN(n5643) );
  OAI21_X1 U5359 ( .B1(n9274), .B2(n5104), .A(n9272), .ZN(n5641) );
  INV_X1 U5360 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5356) );
  AND2_X1 U5361 ( .A1(n5202), .A2(n5200), .ZN(n5196) );
  OR2_X1 U5362 ( .A1(n8633), .A2(n5513), .ZN(n5512) );
  INV_X1 U5363 ( .A(n5526), .ZN(n5210) );
  NOR2_X1 U5364 ( .A1(n8614), .A2(n5527), .ZN(n5526) );
  INV_X1 U5365 ( .A(n6399), .ZN(n5527) );
  NOR2_X1 U5366 ( .A1(n10957), .A2(n5508), .ZN(n5507) );
  INV_X1 U5367 ( .A(n6334), .ZN(n5508) );
  INV_X1 U5368 ( .A(n6303), .ZN(n6390) );
  AOI21_X1 U5370 ( .B1(n8234), .B2(n8233), .A(n8232), .ZN(n8235) );
  OR2_X1 U5371 ( .A1(n6228), .A2(n6977), .ZN(n8223) );
  AND2_X1 U5372 ( .A1(n5272), .A2(n8832), .ZN(n5271) );
  NOR2_X1 U5373 ( .A1(n9052), .A2(n8824), .ZN(n8169) );
  AND2_X1 U5374 ( .A1(n9052), .A2(n8824), .ZN(n8172) );
  NAND2_X1 U5375 ( .A1(n8845), .A2(n5579), .ZN(n5578) );
  NAND2_X1 U5376 ( .A1(n8866), .A2(n8164), .ZN(n5579) );
  OR2_X1 U5377 ( .A1(n9074), .A2(n8534), .ZN(n8145) );
  NOR2_X1 U5378 ( .A1(n9079), .A2(n5484), .ZN(n5483) );
  INV_X1 U5379 ( .A(n8934), .ZN(n5484) );
  NAND2_X1 U5380 ( .A1(n5601), .A2(n7393), .ZN(n5116) );
  NAND2_X1 U5381 ( .A1(n5601), .A2(n5603), .ZN(n5115) );
  NAND2_X1 U5382 ( .A1(n8089), .A2(n8088), .ZN(n5942) );
  OR2_X1 U5383 ( .A1(n10962), .A2(n7507), .ZN(n8086) );
  NAND2_X1 U5384 ( .A1(n8071), .A2(n8070), .ZN(n5895) );
  NAND2_X1 U5385 ( .A1(n6229), .A2(n8227), .ZN(n8237) );
  NOR2_X1 U5386 ( .A1(n6230), .A2(n7160), .ZN(n6671) );
  INV_X1 U5387 ( .A(n6445), .ZN(n7156) );
  INV_X1 U5388 ( .A(n5587), .ZN(n5586) );
  OAI21_X1 U5389 ( .B1(n5048), .B2(n5588), .A(n5589), .ZN(n5587) );
  NOR2_X1 U5390 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5605) );
  INV_X1 U5391 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5607) );
  INV_X1 U5392 ( .A(n7445), .ZN(n5224) );
  NOR2_X1 U5393 ( .A1(n7707), .A2(n7709), .ZN(n5629) );
  NAND2_X1 U5394 ( .A1(n7707), .A2(n7709), .ZN(n5631) );
  NOR2_X1 U5395 ( .A1(n5629), .A2(n5625), .ZN(n5624) );
  INV_X1 U5396 ( .A(n7689), .ZN(n5625) );
  AND2_X1 U5397 ( .A1(n5241), .A2(n9231), .ZN(n5240) );
  NAND2_X1 U5398 ( .A1(n5243), .A2(n5242), .ZN(n5241) );
  INV_X1 U5399 ( .A(n5613), .ZN(n8292) );
  OAI21_X1 U5400 ( .B1(n8267), .B2(n5069), .A(n5612), .ZN(n5613) );
  OR2_X1 U5401 ( .A1(n5617), .A2(n9152), .ZN(n5612) );
  NAND2_X1 U5402 ( .A1(n9588), .A2(n9589), .ZN(n5160) );
  AND2_X1 U5403 ( .A1(n9460), .A2(n9426), .ZN(n9449) );
  AND2_X1 U5404 ( .A1(n10322), .A2(n9607), .ZN(n9450) );
  INV_X1 U5405 ( .A(n5173), .ZN(n5172) );
  NOR2_X1 U5406 ( .A1(n9445), .A2(n5177), .ZN(n5446) );
  INV_X1 U5407 ( .A(n9478), .ZN(n5448) );
  NAND2_X1 U5408 ( .A1(n8459), .A2(n5382), .ZN(n5381) );
  INV_X1 U5409 ( .A(n8458), .ZN(n5382) );
  NOR2_X1 U5410 ( .A1(n5386), .A2(n5176), .ZN(n5175) );
  INV_X1 U5411 ( .A(n8453), .ZN(n5176) );
  INV_X1 U5412 ( .A(n5387), .ZN(n5386) );
  NOR2_X1 U5413 ( .A1(n5444), .A2(n9444), .ZN(n5441) );
  NOR2_X1 U5414 ( .A1(n10358), .A2(n10364), .ZN(n5319) );
  INV_X1 U5415 ( .A(n9546), .ZN(n5462) );
  OAI21_X1 U5416 ( .B1(n5038), .B2(n5466), .A(n5465), .ZN(n5464) );
  OR2_X1 U5417 ( .A1(n10389), .A2(n10250), .ZN(n9551) );
  INV_X1 U5418 ( .A(n5455), .ZN(n5454) );
  OR2_X1 U5419 ( .A1(n7886), .A2(n9264), .ZN(n9526) );
  NOR2_X1 U5420 ( .A1(n10406), .A2(n10412), .ZN(n5327) );
  NAND2_X1 U5421 ( .A1(n7287), .A2(n5043), .ZN(n7418) );
  INV_X1 U5422 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U5423 ( .A1(n6204), .A2(n6203), .ZN(n8000) );
  NAND2_X1 U5424 ( .A1(n6157), .A2(n6156), .ZN(n6167) );
  INV_X1 U5425 ( .A(n6105), .ZN(n5556) );
  AOI21_X1 U5426 ( .B1(n5295), .B2(n5293), .A(n5098), .ZN(n5292) );
  INV_X1 U5427 ( .A(n5742), .ZN(n5293) );
  INV_X1 U5428 ( .A(n5295), .ZN(n5294) );
  NAND2_X1 U5429 ( .A1(n5050), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U5430 ( .A1(n6051), .A2(n5739), .ZN(n6064) );
  AOI21_X1 U5431 ( .B1(n5286), .B2(n5288), .A(n5075), .ZN(n5285) );
  NAND2_X1 U5432 ( .A1(n5736), .A2(SI_18_), .ZN(n5739) );
  NAND2_X1 U5433 ( .A1(n5723), .A2(SI_14_), .ZN(n5727) );
  NAND2_X1 U5434 ( .A1(n5722), .A2(n5721), .ZN(n5986) );
  AOI21_X1 U5435 ( .B1(n5545), .B2(n5548), .A(n5076), .ZN(n5303) );
  NAND2_X1 U5436 ( .A1(n5717), .A2(SI_12_), .ZN(n5304) );
  NAND2_X1 U5437 ( .A1(n5715), .A2(SI_11_), .ZN(n5716) );
  INV_X1 U5438 ( .A(SI_10_), .ZN(n9662) );
  NAND2_X1 U5439 ( .A1(n5495), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U5440 ( .A1(n5121), .A2(n5122), .ZN(n5668) );
  NAND2_X1 U5441 ( .A1(n5497), .A2(SI_2_), .ZN(n5676) );
  NAND2_X1 U5442 ( .A1(n5194), .A2(n5192), .ZN(n5191) );
  NAND2_X1 U5443 ( .A1(n8641), .A2(n6369), .ZN(n8575) );
  OR2_X1 U5444 ( .A1(n5966), .A2(n9700), .ZN(n5978) );
  NAND2_X1 U5445 ( .A1(n5952), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U5446 ( .A1(n8575), .A2(n8576), .ZN(n8574) );
  INV_X1 U5447 ( .A(n6221), .ZN(n6222) );
  NAND2_X1 U5448 ( .A1(n5329), .A2(n5541), .ZN(n5565) );
  NOR2_X1 U5449 ( .A1(n6229), .A2(n8189), .ZN(n5541) );
  INV_X1 U5450 ( .A(n8188), .ZN(n5542) );
  NAND2_X1 U5451 ( .A1(n5028), .A2(n6223), .ZN(n8240) );
  AND4_X1 U5452 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), .ZN(n7562)
         );
  OR2_X1 U5453 ( .A1(n7890), .A2(n6284), .ZN(n6633) );
  NOR2_X1 U5454 ( .A1(n5974), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6018) );
  AND2_X1 U5455 ( .A1(n8241), .A2(n8227), .ZN(n6585) );
  XNOR2_X1 U5456 ( .A(n9041), .B(n8823), .ZN(n8805) );
  NAND2_X1 U5457 ( .A1(n6183), .A2(n6182), .ZN(n8799) );
  NAND2_X1 U5458 ( .A1(n8865), .A2(n6139), .ZN(n8846) );
  AND2_X1 U5459 ( .A1(n9068), .A2(n5536), .ZN(n6116) );
  NAND2_X1 U5460 ( .A1(n5581), .A2(n5583), .ZN(n8859) );
  AOI21_X1 U5461 ( .B1(n8153), .B2(n5585), .A(n5584), .ZN(n5583) );
  INV_X1 U5462 ( .A(n8157), .ZN(n5584) );
  NOR2_X1 U5463 ( .A1(n9068), .A2(n8894), .ZN(n8885) );
  NAND2_X1 U5464 ( .A1(n8893), .A2(n8897), .ZN(n8894) );
  AND2_X1 U5465 ( .A1(n8144), .A2(n8149), .ZN(n8916) );
  NOR2_X1 U5466 ( .A1(n8916), .A2(n5481), .ZN(n5480) );
  INV_X1 U5467 ( .A(n8141), .ZN(n5481) );
  OR2_X1 U5468 ( .A1(n6079), .A2(n8935), .ZN(n5663) );
  NAND2_X1 U5469 ( .A1(n8926), .A2(n8933), .ZN(n8925) );
  NAND2_X1 U5470 ( .A1(n8982), .A2(n5039), .ZN(n8957) );
  AND2_X1 U5471 ( .A1(n8123), .A2(n8124), .ZN(n8978) );
  AOI21_X1 U5472 ( .B1(n5490), .B2(n8208), .A(n5067), .ZN(n5489) );
  AND2_X1 U5473 ( .A1(n8206), .A2(n5958), .ZN(n5136) );
  NAND2_X1 U5474 ( .A1(n7399), .A2(n5488), .ZN(n5130) );
  AND2_X1 U5475 ( .A1(n5942), .A2(n5927), .ZN(n5488) );
  INV_X1 U5476 ( .A(n5942), .ZN(n8192) );
  NAND2_X1 U5477 ( .A1(n7393), .A2(n5049), .ZN(n7505) );
  INV_X1 U5478 ( .A(n9014), .ZN(n10792) );
  NAND2_X1 U5479 ( .A1(n7394), .A2(n8203), .ZN(n7393) );
  NAND2_X1 U5480 ( .A1(n5900), .A2(n5899), .ZN(n8077) );
  XNOR2_X1 U5481 ( .A(n8077), .B(n8076), .ZN(n7373) );
  AND2_X1 U5482 ( .A1(n6237), .A2(n8070), .ZN(n5599) );
  NAND2_X1 U5483 ( .A1(n5151), .A2(n9017), .ZN(n8071) );
  CLKBUF_X1 U5484 ( .A(n5895), .Z(n5145) );
  AND2_X1 U5485 ( .A1(n9020), .A2(n8200), .ZN(n5880) );
  OAI21_X1 U5486 ( .B1(n10806), .B2(n8062), .A(n8060), .ZN(n9013) );
  OAI21_X1 U5487 ( .B1(n7469), .B2(n6692), .A(n6686), .ZN(n5143) );
  OR2_X1 U5488 ( .A1(n10743), .A2(n8227), .ZN(n7157) );
  NAND2_X1 U5489 ( .A1(n6004), .A2(n6003), .ZN(n9109) );
  NAND2_X1 U5490 ( .A1(n5984), .A2(n8103), .ZN(n11014) );
  OR2_X1 U5491 ( .A1(n7331), .A2(n6128), .ZN(n5879) );
  OR2_X1 U5492 ( .A1(n10469), .A2(n6281), .ZN(n6282) );
  AND2_X1 U5493 ( .A1(n6633), .A2(n10621), .ZN(n10471) );
  INV_X1 U5494 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U5495 ( .A1(n5873), .A2(n5752), .ZN(n5897) );
  AOI21_X1 U5496 ( .B1(n5217), .B2(n7344), .A(n5224), .ZN(n5223) );
  INV_X1 U5497 ( .A(n7236), .ZN(n5217) );
  NOR2_X1 U5498 ( .A1(n5224), .A2(n5222), .ZN(n5221) );
  INV_X1 U5499 ( .A(n7327), .ZN(n5222) );
  OAI21_X1 U5500 ( .B1(n8267), .B2(n5068), .A(n5617), .ZN(n9151) );
  INV_X1 U5501 ( .A(n5103), .ZN(n5614) );
  OR2_X1 U5502 ( .A1(n7546), .A2(n7721), .ZN(n7715) );
  NAND2_X1 U5503 ( .A1(n7690), .A2(n7689), .ZN(n5632) );
  AND2_X1 U5504 ( .A1(n5232), .A2(n5647), .ZN(n5231) );
  NOR2_X1 U5505 ( .A1(n5649), .A2(n5648), .ZN(n5647) );
  NAND2_X1 U5506 ( .A1(n5236), .A2(n5233), .ZN(n5232) );
  NAND2_X1 U5507 ( .A1(n5080), .A2(n5645), .ZN(n5637) );
  AND2_X1 U5508 ( .A1(n8279), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8281) );
  OAI21_X1 U5509 ( .B1(n7231), .B2(n7232), .A(n7229), .ZN(n7328) );
  XNOR2_X1 U5510 ( .A(n5216), .B(n8418), .ZN(n7055) );
  INV_X1 U5511 ( .A(n7007), .ZN(n5216) );
  AND3_X1 U5512 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n7241) );
  INV_X1 U5513 ( .A(n9449), .ZN(n9456) );
  INV_X1 U5514 ( .A(n9450), .ZN(n9594) );
  AND4_X1 U5515 ( .A1(n8381), .A2(n8380), .A3(n8379), .A4(n8378), .ZN(n8457)
         );
  AND4_X1 U5516 ( .A1(n7720), .A2(n7719), .A3(n7718), .A4(n7717), .ZN(n7880)
         );
  XNOR2_X1 U5517 ( .A(n10607), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n10604) );
  OR2_X1 U5518 ( .A1(n6549), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6833) );
  NOR2_X1 U5519 ( .A1(n10545), .A2(n5090), .ZN(n10565) );
  NOR2_X1 U5520 ( .A1(n10031), .A2(n5100), .ZN(n10040) );
  AOI21_X1 U5521 ( .B1(n5435), .B2(n5437), .A(n9383), .ZN(n5433) );
  INV_X1 U5522 ( .A(n5180), .ZN(n5179) );
  NAND2_X1 U5523 ( .A1(n5184), .A2(n8464), .ZN(n5183) );
  OAI21_X1 U5524 ( .B1(n5181), .B2(n10098), .A(n8465), .ZN(n5180) );
  AND4_X1 U5525 ( .A1(n8471), .A2(n8470), .A3(n8469), .A4(n8468), .ZN(n9467)
         );
  OAI21_X1 U5526 ( .B1(n10109), .B2(n5437), .A(n5435), .ZN(n8503) );
  NAND2_X1 U5527 ( .A1(n5434), .A2(n5438), .ZN(n8504) );
  AND4_X1 U5528 ( .A1(n8250), .A2(n8249), .A3(n8248), .A4(n8247), .ZN(n10111)
         );
  INV_X1 U5529 ( .A(n8459), .ZN(n5383) );
  NAND2_X1 U5530 ( .A1(n10162), .A2(n10163), .ZN(n10161) );
  AOI21_X1 U5531 ( .B1(n5387), .B2(n5385), .A(n5059), .ZN(n5384) );
  INV_X1 U5532 ( .A(n8455), .ZN(n5385) );
  NAND2_X1 U5533 ( .A1(n8454), .A2(n5175), .ZN(n5174) );
  NAND2_X1 U5534 ( .A1(n5174), .A2(n5173), .ZN(n10152) );
  AND2_X1 U5535 ( .A1(n9482), .A2(n9483), .ZN(n10178) );
  NAND2_X1 U5536 ( .A1(n8454), .A2(n8453), .ZN(n10185) );
  OR2_X1 U5537 ( .A1(n10185), .A2(n10191), .ZN(n10186) );
  NAND2_X1 U5538 ( .A1(n10203), .A2(n10206), .ZN(n10202) );
  NAND2_X1 U5539 ( .A1(n5167), .A2(n8450), .ZN(n10219) );
  AOI21_X1 U5540 ( .B1(n10275), .B2(n9549), .A(n9335), .ZN(n10249) );
  INV_X1 U5541 ( .A(n8447), .ZN(n5362) );
  INV_X1 U5542 ( .A(n9528), .ZN(n5466) );
  AND2_X1 U5543 ( .A1(n8443), .A2(n8444), .ZN(n5169) );
  AND2_X1 U5544 ( .A1(n9528), .A2(n9524), .ZN(n10307) );
  NAND2_X1 U5545 ( .A1(n9526), .A2(n9530), .ZN(n9438) );
  NAND2_X1 U5546 ( .A1(n7794), .A2(n9429), .ZN(n7850) );
  NOR2_X1 U5547 ( .A1(n7789), .A2(n10412), .ZN(n7856) );
  NAND2_X1 U5548 ( .A1(n10908), .A2(n7531), .ZN(n7772) );
  NAND2_X1 U5549 ( .A1(n10512), .A2(n9591), .ZN(n10917) );
  OR2_X1 U5550 ( .A1(n6871), .A2(n7123), .ZN(n6890) );
  NAND2_X1 U5551 ( .A1(n8008), .A2(n8007), .ZN(n11047) );
  AOI21_X1 U5552 ( .B1(n10324), .B2(n10711), .A(n5323), .ZN(n10325) );
  AND2_X1 U5553 ( .A1(n10323), .A2(n11048), .ZN(n5323) );
  INV_X1 U5554 ( .A(n5475), .ZN(n10326) );
  NAND2_X1 U5555 ( .A1(n7971), .A2(n7970), .ZN(n10393) );
  NAND2_X1 U5556 ( .A1(n7983), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6886) );
  OAI211_X1 U5557 ( .C1(P1_B_REG_SCAN_IN), .C2(n7891), .A(n6840), .B(n6530), 
        .ZN(n6925) );
  XNOR2_X1 U5558 ( .A(n8025), .B(n8024), .ZN(n9391) );
  NAND2_X1 U5559 ( .A1(n8020), .A2(n8019), .ZN(n8025) );
  NOR2_X1 U5560 ( .A1(n5650), .A2(n5469), .ZN(n5468) );
  NAND2_X1 U5561 ( .A1(n5651), .A2(n6483), .ZN(n5650) );
  INV_X1 U5562 ( .A(n5470), .ZN(n5469) );
  NAND2_X1 U5563 ( .A1(n6091), .A2(n6090), .ZN(n6106) );
  OR2_X1 U5564 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  NAND2_X1 U5565 ( .A1(n6049), .A2(n6048), .ZN(n6051) );
  INV_X1 U5566 ( .A(n6032), .ZN(n5562) );
  XNOR2_X1 U5567 ( .A(n5306), .B(n5150), .ZN(n7749) );
  XNOR2_X1 U5568 ( .A(n5717), .B(SI_12_), .ZN(n5150) );
  NOR2_X1 U5569 ( .A1(n5550), .A2(n5944), .ZN(n5549) );
  INV_X1 U5570 ( .A(n5714), .ZN(n5550) );
  NAND2_X1 U5571 ( .A1(n5929), .A2(n5928), .ZN(n5551) );
  XNOR2_X1 U5572 ( .A(n5929), .B(n5928), .ZN(n7700) );
  OR2_X1 U5573 ( .A1(n5911), .A2(n5910), .ZN(n5913) );
  NAND2_X1 U5574 ( .A1(n5870), .A2(n5696), .ZN(n5882) );
  AND2_X1 U5575 ( .A1(n5701), .A2(n5700), .ZN(n5881) );
  INV_X1 U5576 ( .A(n5867), .ZN(n5148) );
  OAI21_X1 U5577 ( .B1(n5497), .B2(SI_2_), .A(n5676), .ZN(n5809) );
  NAND2_X1 U5578 ( .A1(n5537), .A2(n6107), .ZN(n9068) );
  NAND2_X1 U5579 ( .A1(n6144), .A2(n6143), .ZN(n9057) );
  NAND2_X1 U5580 ( .A1(n6024), .A2(n6023), .ZN(n9105) );
  OAI211_X1 U5581 ( .C1(n7218), .C2(n6128), .A(n5859), .B(n5066), .ZN(n10810)
         );
  INV_X1 U5582 ( .A(n10964), .ZN(n10890) );
  XNOR2_X1 U5583 ( .A(n6275), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8241) );
  NAND2_X1 U5584 ( .A1(n6038), .A2(n6037), .ZN(n9100) );
  OR2_X1 U5585 ( .A1(n7975), .A2(n6128), .ZN(n6038) );
  OR2_X1 U5586 ( .A1(n6128), .A2(n7059), .ZN(n5849) );
  NAND2_X1 U5587 ( .A1(n5262), .A2(n5260), .ZN(n9034) );
  OR2_X1 U5588 ( .A1(n8781), .A2(n5263), .ZN(n5262) );
  INV_X1 U5589 ( .A(n9032), .ZN(n5263) );
  AND2_X1 U5590 ( .A1(n6257), .A2(n8797), .ZN(n6258) );
  NOR2_X1 U5591 ( .A1(n5767), .A2(n5258), .ZN(n5257) );
  NOR2_X1 U5592 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5258) );
  AND2_X1 U5593 ( .A1(n6840), .A2(n6490), .ZN(n6911) );
  NAND2_X1 U5594 ( .A1(n7952), .A2(n7951), .ZN(n10333) );
  INV_X1 U5595 ( .A(n5236), .ZN(n5234) );
  NOR2_X1 U5596 ( .A1(n5238), .A2(n5228), .ZN(n5227) );
  OR2_X1 U5597 ( .A1(n9197), .A2(n9309), .ZN(n5238) );
  INV_X1 U5598 ( .A(n5231), .ZN(n5228) );
  NAND2_X1 U5599 ( .A1(n7950), .A2(n7949), .ZN(n10328) );
  NAND2_X1 U5600 ( .A1(n7977), .A2(n7976), .ZN(n10383) );
  NAND2_X1 U5601 ( .A1(n7988), .A2(n7987), .ZN(n10368) );
  OAI21_X1 U5602 ( .B1(n6936), .B2(n6938), .A(n10937), .ZN(n9220) );
  AND4_X1 U5603 ( .A1(n6730), .A2(n6729), .A3(n6728), .A4(n6727), .ZN(n10110)
         );
  INV_X1 U5604 ( .A(n9309), .ZN(n9295) );
  INV_X1 U5605 ( .A(n10293), .ZN(n9533) );
  INV_X1 U5606 ( .A(n10303), .ZN(n10007) );
  INV_X1 U5607 ( .A(n7880), .ZN(n10009) );
  OR2_X1 U5608 ( .A1(n5031), .A2(n6862), .ZN(n6865) );
  XNOR2_X1 U5609 ( .A(n10040), .B(n10047), .ZN(n10033) );
  NOR2_X1 U5610 ( .A1(n10033), .A2(n10032), .ZN(n10041) );
  XNOR2_X1 U5611 ( .A(n5255), .B(n5110), .ZN(n5254) );
  NOR2_X1 U5612 ( .A1(n10581), .A2(n5256), .ZN(n5255) );
  AND2_X1 U5613 ( .A1(n10586), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5256) );
  AND2_X1 U5614 ( .A1(n10104), .A2(n10103), .ZN(n10336) );
  NAND2_X1 U5615 ( .A1(n10100), .A2(n10920), .ZN(n10104) );
  NAND2_X1 U5616 ( .A1(n5178), .A2(n8464), .ZN(n10089) );
  NAND2_X1 U5617 ( .A1(n8462), .A2(n5185), .ZN(n5178) );
  OAI21_X1 U5618 ( .B1(n7413), .B2(n5030), .A(n7414), .ZN(n7450) );
  AND2_X1 U5619 ( .A1(n10942), .A2(n7125), .ZN(n10932) );
  NAND2_X1 U5620 ( .A1(n10326), .A2(n10325), .ZN(n5188) );
  OAI211_X1 U5621 ( .C1(n5374), .C2(n5368), .A(n5367), .B(n5365), .ZN(n10327)
         );
  OR2_X1 U5622 ( .A1(n8502), .A2(n5368), .ZN(n5367) );
  NAND2_X1 U5623 ( .A1(n8502), .A2(n5366), .ZN(n5365) );
  OAI21_X1 U5624 ( .B1(n10326), .B2(n11051), .A(n5372), .ZN(n5370) );
  OR2_X1 U5625 ( .A1(n11054), .A2(n5373), .ZN(n5372) );
  INV_X1 U5626 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5373) );
  NAND2_X1 U5627 ( .A1(n6844), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U5628 ( .A1(n6522), .A2(n6473), .ZN(n6844) );
  AOI21_X1 U5629 ( .B1(n9637), .B2(n5390), .A(n5096), .ZN(n9641) );
  NOR2_X1 U5630 ( .A1(n9636), .A2(n9635), .ZN(n9637) );
  NAND2_X1 U5631 ( .A1(SI_27_), .A2(n9639), .ZN(n9640) );
  NAND2_X1 U5632 ( .A1(n9658), .A2(keyinput_143), .ZN(n5412) );
  NAND2_X1 U5633 ( .A1(n9659), .A2(SI_17_), .ZN(n5411) );
  AOI21_X1 U5634 ( .B1(n5409), .B2(n5408), .A(n5407), .ZN(n9666) );
  NOR2_X1 U5635 ( .A1(n9674), .A2(n9675), .ZN(n5417) );
  NAND2_X1 U5636 ( .A1(n5420), .A2(n5419), .ZN(n5418) );
  NAND2_X1 U5637 ( .A1(n9669), .A2(SI_9_), .ZN(n5420) );
  NAND2_X1 U5638 ( .A1(n9668), .A2(keyinput_151), .ZN(n5419) );
  AOI211_X1 U5639 ( .C1(n9685), .C2(n9684), .A(n9683), .B(n9682), .ZN(n9692)
         );
  NAND2_X1 U5640 ( .A1(n5347), .A2(n8053), .ZN(n8055) );
  NAND2_X1 U5641 ( .A1(n9716), .A2(n9713), .ZN(n5424) );
  NAND2_X1 U5642 ( .A1(n8736), .A2(n9714), .ZN(n5425) );
  NOR2_X1 U5643 ( .A1(n5423), .A2(n5421), .ZN(n9724) );
  NAND2_X1 U5644 ( .A1(n5105), .A2(n5422), .ZN(n5421) );
  AOI21_X1 U5645 ( .B1(n9708), .B2(n5425), .A(n5424), .ZN(n5423) );
  NAND2_X1 U5646 ( .A1(n9715), .A2(keyinput_183), .ZN(n5422) );
  NAND2_X1 U5647 ( .A1(n8087), .A2(n8089), .ZN(n5345) );
  MUX2_X1 U5648 ( .A(n8091), .B(n8090), .S(n8186), .Z(n8093) );
  NOR3_X1 U5649 ( .A1(n8083), .A2(n8082), .A3(n8081), .ZN(n5346) );
  INV_X1 U5650 ( .A(n8102), .ZN(n8104) );
  AOI21_X1 U5651 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput_201), .A(n9740), 
        .ZN(n5431) );
  INV_X1 U5652 ( .A(keyinput_205), .ZN(n5427) );
  INV_X1 U5653 ( .A(n8151), .ZN(n5336) );
  INV_X1 U5654 ( .A(n8131), .ZN(n8127) );
  NAND2_X1 U5655 ( .A1(n9522), .A2(n9521), .ZN(n9531) );
  AOI21_X1 U5656 ( .B1(n5428), .B2(n5426), .A(n5046), .ZN(n9748) );
  XNOR2_X1 U5657 ( .A(n9743), .B(n5427), .ZN(n5426) );
  OAI21_X1 U5658 ( .B1(n5337), .B2(n5334), .A(n5332), .ZN(n5331) );
  OAI21_X1 U5659 ( .B1(n9774), .B2(n5111), .A(n5406), .ZN(n5405) );
  AND2_X1 U5660 ( .A1(n9778), .A2(n5112), .ZN(n5406) );
  INV_X1 U5661 ( .A(n8173), .ZN(n5343) );
  NOR2_X1 U5662 ( .A1(n8169), .A2(n8186), .ZN(n5340) );
  OAI21_X1 U5663 ( .B1(n5045), .B2(n5155), .A(n5070), .ZN(n9573) );
  NAND2_X1 U5664 ( .A1(n9571), .A2(n10163), .ZN(n5155) );
  NAND2_X1 U5665 ( .A1(n9788), .A2(n5401), .ZN(n5400) );
  AND2_X1 U5666 ( .A1(n9787), .A2(n9786), .ZN(n5401) );
  INV_X1 U5667 ( .A(n9790), .ZN(n5399) );
  NOR2_X1 U5668 ( .A1(n5657), .A2(n5396), .ZN(n5395) );
  NOR2_X1 U5669 ( .A1(keyinput_245), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n5396) );
  INV_X1 U5670 ( .A(n6423), .ZN(n5513) );
  NAND2_X1 U5671 ( .A1(n8219), .A2(n8186), .ZN(n5543) );
  AOI21_X1 U5672 ( .B1(n8226), .B2(n8225), .A(n8224), .ZN(n8230) );
  NAND2_X1 U5673 ( .A1(n8116), .A2(n8112), .ZN(n5588) );
  NOR2_X1 U5674 ( .A1(n5591), .A2(n5590), .ZN(n5589) );
  INV_X1 U5675 ( .A(n8994), .ZN(n5590) );
  INV_X1 U5676 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5525) );
  AND3_X1 U5677 ( .A1(n6016), .A2(n6015), .A3(n6014), .ZN(n6017) );
  NAND2_X1 U5678 ( .A1(n5524), .A2(n6020), .ZN(n5522) );
  INV_X1 U5679 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6020) );
  INV_X1 U5680 ( .A(n9233), .ZN(n5243) );
  INV_X1 U5681 ( .A(n5610), .ZN(n5242) );
  NOR2_X1 U5682 ( .A1(n9233), .A2(n9225), .ZN(n5244) );
  NAND2_X1 U5683 ( .A1(n5103), .A2(n8274), .ZN(n5615) );
  NAND2_X1 U5684 ( .A1(n5397), .A2(n5395), .ZN(n9802) );
  NOR2_X1 U5685 ( .A1(n5456), .A2(n5452), .ZN(n5451) );
  OAI21_X1 U5686 ( .B1(n7748), .B2(n5456), .A(n9521), .ZN(n5455) );
  OR2_X1 U5687 ( .A1(n10328), .A2(n9188), .ZN(n9468) );
  INV_X1 U5688 ( .A(SI_28_), .ZN(n9632) );
  NOR2_X1 U5689 ( .A1(n6152), .A2(n5311), .ZN(n5310) );
  INV_X1 U5690 ( .A(n6140), .ZN(n5311) );
  AOI21_X1 U5691 ( .B1(n6063), .B2(n5742), .A(n5296), .ZN(n5295) );
  INV_X1 U5692 ( .A(n6080), .ZN(n5296) );
  INV_X1 U5693 ( .A(n5303), .ZN(n5302) );
  AOI21_X1 U5694 ( .B1(n5303), .B2(n5301), .A(n5079), .ZN(n5300) );
  INV_X1 U5695 ( .A(n5545), .ZN(n5301) );
  INV_X1 U5696 ( .A(SI_9_), .ZN(n9668) );
  NAND2_X1 U5697 ( .A1(n5124), .A2(n5123), .ZN(n5121) );
  NAND2_X1 U5698 ( .A1(n5120), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5669) );
  NAND2_X1 U5699 ( .A1(n5356), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5120) );
  NAND2_X1 U5700 ( .A1(n5537), .A2(n5534), .ZN(n8154) );
  NOR2_X1 U5701 ( .A1(n8860), .A2(n5535), .ZN(n5534) );
  INV_X1 U5702 ( .A(n6107), .ZN(n5535) );
  NOR2_X1 U5703 ( .A1(n5573), .A2(n5570), .ZN(n5569) );
  INV_X1 U5704 ( .A(n6244), .ZN(n5570) );
  INV_X1 U5705 ( .A(n8129), .ZN(n5573) );
  OR2_X1 U5706 ( .A1(n6025), .A2(n8579), .ZN(n6039) );
  NOR2_X1 U5707 ( .A1(n5279), .A2(n7621), .ZN(n5278) );
  OR2_X1 U5708 ( .A1(n7516), .A2(n10962), .ZN(n5279) );
  NOR2_X1 U5709 ( .A1(n5597), .A2(n7373), .ZN(n5596) );
  INV_X1 U5710 ( .A(n8071), .ZN(n5597) );
  INV_X1 U5711 ( .A(n5599), .ZN(n5594) );
  INV_X1 U5712 ( .A(n8078), .ZN(n5593) );
  NAND2_X1 U5713 ( .A1(n5896), .A2(n5486), .ZN(n5485) );
  NAND2_X1 U5714 ( .A1(n5816), .A2(n7463), .ZN(n6232) );
  NAND2_X1 U5715 ( .A1(n5270), .A2(n5269), .ZN(n7466) );
  INV_X1 U5716 ( .A(n7464), .ZN(n5270) );
  NAND2_X1 U5717 ( .A1(n6675), .A2(n7160), .ZN(n7464) );
  AOI21_X1 U5718 ( .B1(n5077), .B2(n9261), .A(n5618), .ZN(n5617) );
  AND2_X1 U5719 ( .A1(n5619), .A2(n9260), .ZN(n5618) );
  NOR2_X1 U5720 ( .A1(n9260), .A2(n9261), .ZN(n5620) );
  NAND2_X1 U5721 ( .A1(n5636), .A2(n5634), .ZN(n8385) );
  AOI21_X1 U5722 ( .B1(n5642), .B2(n5635), .A(n5641), .ZN(n5634) );
  INV_X1 U5723 ( .A(n5637), .ZN(n5635) );
  INV_X1 U5724 ( .A(n9213), .ZN(n5233) );
  INV_X1 U5725 ( .A(n8424), .ZN(n5648) );
  OR2_X1 U5726 ( .A1(n5185), .A2(n5182), .ZN(n5181) );
  INV_X1 U5727 ( .A(n8464), .ZN(n5182) );
  AND2_X1 U5728 ( .A1(n9473), .A2(n10112), .ZN(n5439) );
  NAND2_X1 U5729 ( .A1(n5078), .A2(n9473), .ZN(n5438) );
  AOI21_X1 U5730 ( .B1(n5438), .B2(n5436), .A(n9447), .ZN(n5435) );
  INV_X1 U5731 ( .A(n5439), .ZN(n5436) );
  INV_X1 U5732 ( .A(n5438), .ZN(n5437) );
  NOR2_X1 U5733 ( .A1(n5318), .A2(n10353), .ZN(n5317) );
  INV_X1 U5734 ( .A(n5319), .ZN(n5318) );
  OR2_X1 U5735 ( .A1(n10383), .A2(n8479), .ZN(n9555) );
  AND2_X1 U5736 ( .A1(n10274), .A2(n5361), .ZN(n5360) );
  NAND2_X1 U5737 ( .A1(n5465), .A2(n8447), .ZN(n5361) );
  NAND2_X1 U5738 ( .A1(n5327), .A2(n10996), .ZN(n5326) );
  NAND2_X1 U5739 ( .A1(n7521), .A2(n5047), .ZN(n10905) );
  NAND2_X1 U5740 ( .A1(n7418), .A2(n7416), .ZN(n10912) );
  XNOR2_X1 U5741 ( .A(n10736), .B(n6949), .ZN(n9434) );
  NAND2_X1 U5742 ( .A1(n6889), .A2(n10730), .ZN(n9559) );
  AND2_X1 U5743 ( .A1(n8001), .A2(n6207), .ZN(n7999) );
  INV_X1 U5744 ( .A(n6476), .ZN(n5651) );
  INV_X1 U5745 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6474) );
  INV_X1 U5746 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6485) );
  INV_X1 U5747 ( .A(SI_23_), .ZN(n6120) );
  NAND2_X1 U5748 ( .A1(n6492), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6496) );
  INV_X1 U5749 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6467) );
  INV_X1 U5750 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6516) );
  INV_X1 U5751 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6463) );
  INV_X1 U5752 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U5753 ( .A1(n7957), .A2(n8036), .ZN(n5537) );
  NAND2_X1 U5754 ( .A1(n5511), .A2(n6429), .ZN(n5201) );
  OAI21_X1 U5755 ( .B1(n5202), .B2(n6429), .A(n5198), .ZN(n5197) );
  NAND2_X1 U5756 ( .A1(n7085), .A2(n5514), .ZN(n10888) );
  AND2_X1 U5757 ( .A1(n6329), .A2(n6322), .ZN(n5514) );
  NAND2_X1 U5758 ( .A1(n10815), .A2(n8034), .ZN(n5212) );
  NOR2_X1 U5759 ( .A1(n5500), .A2(n5036), .ZN(n5499) );
  INV_X1 U5760 ( .A(n5507), .ZN(n5500) );
  INV_X1 U5761 ( .A(n5503), .ZN(n5502) );
  OAI21_X1 U5762 ( .B1(n5504), .B2(n5036), .A(n7560), .ZN(n5503) );
  INV_X1 U5763 ( .A(n8542), .ZN(n10793) );
  INV_X1 U5764 ( .A(n6407), .ZN(n5211) );
  AOI21_X1 U5765 ( .B1(n5210), .B2(n6407), .A(n5074), .ZN(n5209) );
  NOR2_X1 U5766 ( .A1(n5920), .A2(n8682), .ZN(n5936) );
  AOI21_X1 U5767 ( .B1(n8548), .B2(n5193), .A(n5062), .ZN(n5192) );
  INV_X1 U5768 ( .A(n8622), .ZN(n5193) );
  NAND2_X1 U5769 ( .A1(n5529), .A2(n5528), .ZN(n7892) );
  AND2_X1 U5770 ( .A1(n6356), .A2(n6349), .ZN(n5528) );
  NAND2_X1 U5771 ( .A1(n7681), .A2(n7682), .ZN(n5529) );
  OR2_X1 U5772 ( .A1(n5978), .A2(n5977), .ZN(n5992) );
  NAND2_X1 U5773 ( .A1(n6400), .A2(n5526), .ZN(n8612) );
  AND2_X1 U5774 ( .A1(n5505), .A2(n10958), .ZN(n5504) );
  INV_X1 U5775 ( .A(n7493), .ZN(n5505) );
  INV_X1 U5776 ( .A(n6592), .ZN(n6825) );
  NOR2_X1 U5777 ( .A1(n6039), .A2(n8736), .ZN(n6055) );
  NOR2_X1 U5778 ( .A1(n5860), .A2(n9726), .ZN(n5889) );
  NOR2_X1 U5779 ( .A1(n5992), .A2(n5991), .ZN(n6005) );
  INV_X1 U5780 ( .A(n8237), .ZN(n5567) );
  AND4_X1 U5781 ( .A1(n6010), .A2(n6009), .A3(n6008), .A4(n6007), .ZN(n8578)
         );
  AND4_X1 U5782 ( .A1(n5908), .A2(n5907), .A3(n5906), .A4(n5905), .ZN(n8076)
         );
  AND4_X1 U5783 ( .A1(n5855), .A2(n5854), .A3(n5853), .A4(n5852), .ZN(n7091)
         );
  AND2_X1 U5784 ( .A1(n7181), .A2(n7180), .ZN(n7182) );
  INV_X1 U5785 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U5786 ( .A1(n8808), .A2(n5117), .ZN(n8226) );
  NAND2_X1 U5787 ( .A1(n8654), .A2(n8803), .ZN(n5117) );
  NAND2_X1 U5788 ( .A1(n8826), .A2(n8175), .ZN(n8804) );
  NAND2_X1 U5789 ( .A1(n8804), .A2(n8798), .ZN(n8808) );
  AND4_X1 U5790 ( .A1(n6165), .A2(n6164), .A3(n6163), .A4(n6162), .ZN(n8824)
         );
  AOI21_X1 U5791 ( .B1(n8859), .B2(n5575), .A(n5574), .ZN(n8820) );
  AND2_X1 U5792 ( .A1(n8173), .A2(n8164), .ZN(n5575) );
  INV_X1 U5793 ( .A(n5576), .ZN(n5574) );
  AOI21_X1 U5794 ( .B1(n5578), .B2(n8173), .A(n8172), .ZN(n5576) );
  NAND2_X1 U5795 ( .A1(n8885), .A2(n5095), .ZN(n8815) );
  NAND2_X1 U5796 ( .A1(n8885), .A2(n5271), .ZN(n8838) );
  AND2_X1 U5797 ( .A1(n6175), .A2(n6161), .ZN(n8840) );
  NOR2_X1 U5798 ( .A1(n8172), .A2(n8169), .ZN(n8835) );
  NAND2_X1 U5799 ( .A1(n8833), .A2(n8170), .ZN(n8852) );
  OAI21_X1 U5800 ( .B1(n6247), .B2(n5580), .A(n5577), .ZN(n8854) );
  INV_X1 U5801 ( .A(n5578), .ZN(n5577) );
  INV_X1 U5802 ( .A(n6116), .ZN(n5476) );
  NAND2_X1 U5803 ( .A1(n6247), .A2(n6246), .ZN(n8863) );
  NAND2_X1 U5804 ( .A1(n8898), .A2(n8899), .ZN(n8875) );
  NAND2_X1 U5805 ( .A1(n8915), .A2(n8144), .ZN(n8898) );
  INV_X1 U5806 ( .A(n5480), .ZN(n5479) );
  AOI21_X1 U5807 ( .B1(n5480), .B2(n8213), .A(n5483), .ZN(n5478) );
  NAND2_X1 U5808 ( .A1(n5129), .A2(n5571), .ZN(n8937) );
  AND2_X1 U5809 ( .A1(n5572), .A2(n8213), .ZN(n5571) );
  NAND2_X1 U5810 ( .A1(n8965), .A2(n5569), .ZN(n5129) );
  NAND2_X1 U5811 ( .A1(n8943), .A2(n8129), .ZN(n5572) );
  OR2_X1 U5812 ( .A1(n9091), .A2(n8935), .ZN(n8129) );
  NAND2_X1 U5813 ( .A1(n8982), .A2(n5274), .ZN(n8927) );
  AND2_X1 U5814 ( .A1(n5041), .A2(n8931), .ZN(n5274) );
  AND2_X1 U5815 ( .A1(n6055), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6075) );
  AND2_X1 U5816 ( .A1(n6075), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U5817 ( .A1(n8965), .A2(n6244), .ZN(n8947) );
  NAND2_X1 U5818 ( .A1(n8947), .A2(n8946), .ZN(n8945) );
  NAND2_X1 U5819 ( .A1(n6243), .A2(n8123), .ZN(n8967) );
  NAND2_X1 U5820 ( .A1(n8967), .A2(n8966), .ZN(n8965) );
  INV_X1 U5821 ( .A(n8212), .ZN(n8966) );
  NAND2_X1 U5822 ( .A1(n8975), .A2(n6047), .ZN(n8956) );
  NAND2_X1 U5823 ( .A1(n5990), .A2(n5989), .ZN(n7908) );
  NAND2_X1 U5824 ( .A1(n6240), .A2(n5048), .ZN(n7902) );
  AND2_X1 U5825 ( .A1(n11010), .A2(n7916), .ZN(n7917) );
  AND2_X1 U5826 ( .A1(n5114), .A2(n5113), .ZN(n7913) );
  NAND2_X1 U5827 ( .A1(n8206), .A2(n8098), .ZN(n5113) );
  AND3_X1 U5828 ( .A1(n5278), .A2(n5277), .A3(n5276), .ZN(n7916) );
  NAND2_X1 U5829 ( .A1(n5278), .A2(n5277), .ZN(n7733) );
  NOR2_X1 U5830 ( .A1(n7402), .A2(n5279), .ZN(n7616) );
  AND2_X1 U5831 ( .A1(n7393), .A2(n8086), .ZN(n7506) );
  AND4_X1 U5832 ( .A1(n5926), .A2(n5925), .A3(n5924), .A4(n5923), .ZN(n7507)
         );
  NAND2_X1 U5833 ( .A1(n6253), .A2(n6585), .ZN(n10794) );
  NOR2_X1 U5834 ( .A1(n7402), .A2(n10962), .ZN(n7512) );
  INV_X1 U5835 ( .A(n5600), .ZN(n7394) );
  OAI21_X1 U5836 ( .B1(n6238), .B2(n5595), .A(n5592), .ZN(n5600) );
  AOI21_X1 U5837 ( .B1(n5596), .B2(n5594), .A(n5593), .ZN(n5592) );
  INV_X1 U5838 ( .A(n5596), .ZN(n5595) );
  NAND2_X1 U5839 ( .A1(n5135), .A2(n5153), .ZN(n7374) );
  INV_X1 U5840 ( .A(n5145), .ZN(n8074) );
  NOR2_X1 U5841 ( .A1(n9025), .A2(n10863), .ZN(n9027) );
  XNOR2_X1 U5842 ( .A(n8664), .B(n10863), .ZN(n9022) );
  NAND2_X1 U5843 ( .A1(n6232), .A2(n8043), .ZN(n8049) );
  AND2_X1 U5844 ( .A1(n6255), .A2(n6585), .ZN(n9014) );
  AND2_X1 U5845 ( .A1(n8793), .A2(n8800), .ZN(n8781) );
  NAND2_X1 U5846 ( .A1(n6209), .A2(n6208), .ZN(n6228) );
  INV_X1 U5847 ( .A(n10810), .ZN(n10824) );
  INV_X1 U5848 ( .A(n6456), .ZN(n7152) );
  NOR2_X1 U5849 ( .A1(n6289), .A2(n6288), .ZN(n6457) );
  AND2_X1 U5850 ( .A1(n5605), .A2(n5752), .ZN(n5138) );
  AND2_X1 U5851 ( .A1(n6218), .A2(n5604), .ZN(n5763) );
  AND2_X1 U5852 ( .A1(n5606), .A2(n5758), .ZN(n5604) );
  NAND2_X1 U5853 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n5354) );
  INV_X1 U5854 ( .A(n6218), .ZN(n6219) );
  INV_X1 U5855 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5959) );
  INV_X1 U5856 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5751) );
  INV_X1 U5857 ( .A(n8367), .ZN(n8377) );
  NAND2_X1 U5858 ( .A1(n5632), .A2(n7699), .ZN(n7708) );
  NAND2_X1 U5859 ( .A1(n8299), .A2(n8298), .ZN(n5610) );
  XNOR2_X1 U5860 ( .A(n7064), .B(n9185), .ZN(n7223) );
  OAI21_X1 U5861 ( .B1(n7292), .B2(n9187), .A(n7063), .ZN(n7064) );
  AOI21_X1 U5862 ( .B1(n10014), .B2(n9182), .A(n7065), .ZN(n7224) );
  OR2_X1 U5863 ( .A1(n7536), .A2(n7535), .ZN(n7546) );
  AND2_X1 U5864 ( .A1(n6914), .A2(n6913), .ZN(n6980) );
  AOI21_X1 U5865 ( .B1(n9181), .B2(n7108), .A(n6912), .ZN(n6913) );
  OR2_X1 U5866 ( .A1(n6905), .A2(n10611), .ZN(n5659) );
  OR2_X1 U5867 ( .A1(n5630), .A2(n5629), .ZN(n5622) );
  AND2_X1 U5868 ( .A1(n7699), .A2(n5631), .ZN(n5630) );
  XNOR2_X1 U5869 ( .A(n6892), .B(n8418), .ZN(n7011) );
  NAND2_X1 U5870 ( .A1(n7107), .A2(n9181), .ZN(n6901) );
  AND2_X1 U5871 ( .A1(n8301), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8313) );
  OR2_X1 U5872 ( .A1(n6911), .A2(n7111), .ZN(n9187) );
  NAND2_X1 U5873 ( .A1(n5106), .A2(n5646), .ZN(n7446) );
  NAND2_X1 U5874 ( .A1(n7328), .A2(n7327), .ZN(n5646) );
  NAND2_X1 U5875 ( .A1(n7237), .A2(n7236), .ZN(n7329) );
  AND2_X1 U5876 ( .A1(n9297), .A2(n5237), .ZN(n5236) );
  NAND2_X1 U5877 ( .A1(n9212), .A2(n9213), .ZN(n5237) );
  AND2_X1 U5878 ( .A1(n6937), .A2(n9600), .ZN(n6932) );
  AND2_X1 U5879 ( .A1(n8292), .A2(n8294), .ZN(n8289) );
  AND2_X1 U5880 ( .A1(n8297), .A2(n8295), .ZN(n5609) );
  OR2_X1 U5881 ( .A1(n6911), .A2(n6531), .ZN(n6939) );
  NAND2_X1 U5882 ( .A1(n6496), .A2(n6495), .ZN(n6498) );
  AOI211_X1 U5883 ( .C1(n9813), .C2(n9812), .A(n9811), .B(n9810), .ZN(n9816)
         );
  OR2_X1 U5884 ( .A1(n8432), .A2(n7120), .ZN(n6880) );
  NOR2_X1 U5885 ( .A1(n10666), .A2(n5051), .ZN(n10021) );
  OR2_X1 U5886 ( .A1(n10021), .A2(n10020), .ZN(n5247) );
  AND2_X1 U5887 ( .A1(n5247), .A2(n5246), .ZN(n10684) );
  NAND2_X1 U5888 ( .A1(n6568), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U5889 ( .A1(n10684), .A2(n10685), .ZN(n10683) );
  NAND2_X1 U5890 ( .A1(n7998), .A2(n7997), .ZN(n10323) );
  INV_X1 U5891 ( .A(n8509), .ZN(n8473) );
  AND2_X1 U5892 ( .A1(n5378), .A2(n8483), .ZN(n5377) );
  NAND2_X1 U5893 ( .A1(n5379), .A2(n5383), .ZN(n5378) );
  AND2_X1 U5894 ( .A1(n9475), .A2(n10097), .ZN(n10112) );
  NAND2_X1 U5895 ( .A1(n5445), .A2(n5447), .ZN(n10133) );
  AOI21_X1 U5896 ( .B1(n10143), .B2(n5449), .A(n5448), .ZN(n5447) );
  INV_X1 U5897 ( .A(n9481), .ZN(n5449) );
  NAND2_X1 U5898 ( .A1(n10211), .A2(n5317), .ZN(n10155) );
  NAND2_X1 U5899 ( .A1(n5440), .A2(n5442), .ZN(n10177) );
  AOI21_X1 U5900 ( .B1(n10191), .B2(n9360), .A(n5443), .ZN(n5442) );
  INV_X1 U5901 ( .A(n9484), .ZN(n5443) );
  NAND2_X1 U5902 ( .A1(n10211), .A2(n10188), .ZN(n10194) );
  AND3_X1 U5903 ( .A1(n8359), .A2(n8358), .A3(n8357), .ZN(n10205) );
  AND2_X1 U5904 ( .A1(n9565), .A2(n9566), .ZN(n10222) );
  NAND2_X1 U5905 ( .A1(n5168), .A2(n8449), .ZN(n10235) );
  INV_X1 U5906 ( .A(n10223), .ZN(n10251) );
  NAND2_X1 U5907 ( .A1(n5463), .A2(n7836), .ZN(n5459) );
  AOI21_X1 U5908 ( .B1(n5463), .B2(n5466), .A(n5462), .ZN(n5461) );
  NOR2_X1 U5909 ( .A1(n7765), .A2(n7277), .ZN(n8279) );
  AND4_X1 U5910 ( .A1(n8285), .A2(n8284), .A3(n8283), .A4(n8282), .ZN(n10304)
         );
  OR2_X1 U5911 ( .A1(n7826), .A2(n7827), .ZN(n7829) );
  NAND2_X1 U5912 ( .A1(n7824), .A2(n7823), .ZN(n8445) );
  NAND2_X1 U5913 ( .A1(n5389), .A2(n7836), .ZN(n8443) );
  INV_X1 U5914 ( .A(n7829), .ZN(n5389) );
  NOR2_X1 U5915 ( .A1(n7715), .A2(n7714), .ZN(n7755) );
  AND2_X1 U5916 ( .A1(n9438), .A2(n7777), .ZN(n7826) );
  NOR2_X1 U5917 ( .A1(n7789), .A2(n5325), .ZN(n7857) );
  INV_X1 U5918 ( .A(n5327), .ZN(n5325) );
  AND4_X1 U5919 ( .A1(n7760), .A2(n7759), .A3(n7758), .A4(n7757), .ZN(n9264)
         );
  AND2_X1 U5920 ( .A1(n9325), .A2(n9506), .ZN(n9503) );
  NAND2_X1 U5921 ( .A1(n10910), .A2(n10936), .ZN(n10909) );
  AND2_X1 U5922 ( .A1(n9501), .A2(n9500), .ZN(n10913) );
  AND4_X1 U5923 ( .A1(n7245), .A2(n7244), .A3(n7243), .A4(n7242), .ZN(n7428)
         );
  AND4_X1 U5924 ( .A1(n7427), .A2(n7426), .A3(n7425), .A4(n7424), .ZN(n7602)
         );
  NAND2_X1 U5925 ( .A1(n5314), .A2(n10855), .ZN(n10834) );
  AND2_X1 U5926 ( .A1(n9493), .A2(n9349), .ZN(n10838) );
  AND2_X1 U5927 ( .A1(n10835), .A2(n10837), .ZN(n9488) );
  AND4_X1 U5928 ( .A1(n7075), .A2(n7074), .A3(n7073), .A4(n7072), .ZN(n7356)
         );
  OAI22_X1 U5929 ( .A1(n10709), .A2(n10708), .B1(n7107), .B2(n10726), .ZN(
        n7132) );
  NAND2_X1 U5930 ( .A1(n8356), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6928) );
  NAND2_X1 U5931 ( .A1(n10713), .A2(n10712), .ZN(n10710) );
  OR2_X1 U5932 ( .A1(n10707), .A2(n9595), .ZN(n6934) );
  INV_X1 U5933 ( .A(n7124), .ZN(n7144) );
  NOR2_X1 U5934 ( .A1(n9582), .A2(n5375), .ZN(n5366) );
  NAND2_X1 U5935 ( .A1(n7954), .A2(n7953), .ZN(n10338) );
  OR2_X1 U5936 ( .A1(n7993), .A2(n5030), .ZN(n7996) );
  INV_X1 U5937 ( .A(n7450), .ZN(n10876) );
  AND2_X1 U5938 ( .A1(n7144), .A2(n7123), .ZN(n11048) );
  INV_X1 U5939 ( .A(n10711), .ZN(n11043) );
  INV_X1 U5940 ( .A(n11048), .ZN(n11021) );
  XNOR2_X1 U5941 ( .A(n8018), .B(n8017), .ZN(n8497) );
  XNOR2_X1 U5942 ( .A(n8000), .B(n7999), .ZN(n9136) );
  XNOR2_X1 U5943 ( .A(n6200), .B(n6199), .ZN(n8495) );
  NAND2_X1 U5944 ( .A1(n6172), .A2(n6171), .ZN(n6185) );
  XNOR2_X1 U5945 ( .A(n6167), .B(n6166), .ZN(n9142) );
  AND2_X1 U5946 ( .A1(n5313), .A2(n6122), .ZN(n5312) );
  INV_X1 U5947 ( .A(n6125), .ZN(n5313) );
  INV_X1 U5948 ( .A(n5554), .ZN(n5553) );
  NAND2_X1 U5949 ( .A1(n5291), .A2(n5290), .ZN(n5552) );
  OAI21_X1 U5950 ( .B1(n5747), .B2(n5555), .A(n6104), .ZN(n5554) );
  XNOR2_X1 U5951 ( .A(n6500), .B(n5471), .ZN(n7799) );
  OAI21_X1 U5952 ( .B1(n6064), .B2(n5294), .A(n5292), .ZN(n5749) );
  NAND2_X1 U5953 ( .A1(n5557), .A2(n5747), .ZN(n6091) );
  INV_X1 U5954 ( .A(n5749), .ZN(n5557) );
  OAI21_X1 U5955 ( .B1(n6064), .B2(n6063), .A(n5742), .ZN(n6081) );
  INV_X1 U5956 ( .A(n5283), .ZN(n5282) );
  AOI21_X1 U5957 ( .B1(n5283), .B2(n5287), .A(n5281), .ZN(n5280) );
  AND2_X1 U5958 ( .A1(n5561), .A2(n5285), .ZN(n5283) );
  AND2_X1 U5959 ( .A1(n5739), .A2(n5738), .ZN(n6048) );
  OAI21_X1 U5960 ( .B1(n5986), .B2(n5286), .A(n5727), .ZN(n5999) );
  NAND2_X1 U5961 ( .A1(n5299), .A2(n5303), .ZN(n5305) );
  NAND2_X1 U5962 ( .A1(n5929), .A2(n5545), .ZN(n5299) );
  OR2_X1 U5963 ( .A1(n6539), .A2(n6538), .ZN(n6549) );
  NOR2_X1 U5964 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10484), .ZN(n7635) );
  NAND2_X1 U5965 ( .A1(n7085), .A2(n6322), .ZN(n10891) );
  NAND2_X1 U5966 ( .A1(n5510), .A2(n6423), .ZN(n8519) );
  NAND2_X1 U5967 ( .A1(n8632), .A2(n8633), .ZN(n5510) );
  AND4_X1 U5968 ( .A1(n6101), .A2(n6100), .A3(n6099), .A4(n6098), .ZN(n8534)
         );
  NAND2_X1 U5969 ( .A1(n5506), .A2(n10958), .ZN(n7494) );
  INV_X1 U5970 ( .A(n8539), .ZN(n5208) );
  AND4_X1 U5971 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n7685)
         );
  NAND2_X1 U5972 ( .A1(n8574), .A2(n6375), .ZN(n8588) );
  NAND2_X1 U5973 ( .A1(n7320), .A2(n6334), .ZN(n10961) );
  NOR2_X1 U5974 ( .A1(n6445), .A2(n6444), .ZN(n10955) );
  NAND2_X1 U5975 ( .A1(n5190), .A2(n5192), .ZN(n8604) );
  OR2_X1 U5976 ( .A1(n6386), .A2(n5194), .ZN(n5190) );
  AND4_X1 U5977 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .ZN(n7915)
         );
  NAND2_X1 U5978 ( .A1(n5529), .A2(n6349), .ZN(n7894) );
  NAND2_X1 U5979 ( .A1(n6400), .A2(n6399), .ZN(n8615) );
  NAND2_X1 U5980 ( .A1(n6093), .A2(n6092), .ZN(n9074) );
  INV_X1 U5981 ( .A(n5501), .ZN(n7561) );
  AOI21_X1 U5982 ( .B1(n5506), .B2(n5504), .A(n5036), .ZN(n5501) );
  NOR2_X1 U5983 ( .A1(n8585), .A2(n5517), .ZN(n5516) );
  INV_X1 U5984 ( .A(n6375), .ZN(n5517) );
  NAND2_X1 U5985 ( .A1(n6419), .A2(n6418), .ZN(n8632) );
  AND4_X1 U5986 ( .A1(n5997), .A2(n5996), .A3(n5995), .A4(n5994), .ZN(n8646)
         );
  AND2_X1 U5987 ( .A1(n6434), .A2(n6433), .ZN(n10964) );
  AND4_X1 U5988 ( .A1(n6151), .A2(n6150), .A3(n6149), .A4(n6148), .ZN(n8861)
         );
  INV_X1 U5989 ( .A(n8534), .ZN(n8918) );
  AND4_X1 U5990 ( .A1(n5778), .A2(n5777), .A3(n5776), .A4(n5775), .ZN(n8934)
         );
  NAND2_X1 U5991 ( .A1(n5901), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U5992 ( .A1(n5800), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U5993 ( .A1(n5793), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5794) );
  INV_X1 U5994 ( .A(n6633), .ZN(n6462) );
  NAND2_X1 U5995 ( .A1(n8028), .A2(n8027), .ZN(n9032) );
  INV_X1 U5996 ( .A(n8987), .ZN(n10813) );
  XNOR2_X1 U5997 ( .A(n5137), .B(n8217), .ZN(n8795) );
  NAND2_X1 U5998 ( .A1(n8885), .A2(n8162), .ZN(n8848) );
  NAND2_X1 U5999 ( .A1(n8925), .A2(n8141), .ZN(n8910) );
  AND2_X1 U6000 ( .A1(n8925), .A2(n5480), .ZN(n8909) );
  NAND2_X1 U6001 ( .A1(n8982), .A2(n6046), .ZN(n8959) );
  NAND2_X1 U6002 ( .A1(n9005), .A2(n6031), .ZN(n8976) );
  NAND2_X1 U6003 ( .A1(n11014), .A2(n5490), .ZN(n7905) );
  AND2_X1 U6004 ( .A1(n7612), .A2(n5958), .ZN(n7732) );
  NAND2_X1 U6005 ( .A1(n7505), .A2(n8088), .ZN(n7608) );
  NAND2_X1 U6006 ( .A1(n7399), .A2(n5927), .ZN(n7503) );
  NAND2_X1 U6007 ( .A1(n8071), .A2(n5598), .ZN(n7364) );
  NAND2_X1 U6008 ( .A1(n6238), .A2(n5599), .ZN(n5598) );
  AND2_X1 U6009 ( .A1(n10868), .A2(n8066), .ZN(n7385) );
  NAND2_X1 U6010 ( .A1(n9021), .A2(n5880), .ZN(n10868) );
  NAND2_X1 U6011 ( .A1(n10818), .A2(n10811), .ZN(n8963) );
  INV_X1 U6012 ( .A(n9024), .ZN(n9008) );
  OR2_X1 U6013 ( .A1(n7157), .A2(n8239), .ZN(n8987) );
  AND2_X1 U6014 ( .A1(n10818), .A2(n10817), .ZN(n9024) );
  INV_X1 U6015 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n5268) );
  OR2_X1 U6016 ( .A1(n9035), .A2(n11030), .ZN(n9040) );
  XNOR2_X1 U6017 ( .A(n6270), .B(P2_IR_REG_26__SCAN_IN), .ZN(n10468) );
  XNOR2_X1 U6018 ( .A(n6273), .B(P2_IR_REG_25__SCAN_IN), .ZN(n10469) );
  NAND2_X1 U6019 ( .A1(n6271), .A2(n6221), .ZN(n6272) );
  INV_X1 U6020 ( .A(n8241), .ZN(n7678) );
  OAI21_X1 U6021 ( .B1(n6067), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U6022 ( .A1(n6070), .A2(n6069), .ZN(n6216) );
  AND2_X1 U6023 ( .A1(n5948), .A2(n5933), .ZN(n6807) );
  NAND2_X1 U6024 ( .A1(n5897), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U6025 ( .A1(n7328), .A2(n5221), .ZN(n5220) );
  NAND2_X1 U6026 ( .A1(n5223), .A2(n7346), .ZN(n5218) );
  NAND2_X1 U6027 ( .A1(n7446), .A2(n7445), .ZN(n7447) );
  NAND2_X1 U6028 ( .A1(n7708), .A2(n7707), .ZN(n7807) );
  NAND2_X1 U6029 ( .A1(n5632), .A2(n5627), .ZN(n5626) );
  AND2_X1 U6030 ( .A1(n7699), .A2(n5628), .ZN(n5627) );
  INV_X1 U6031 ( .A(n7707), .ZN(n5628) );
  NAND2_X1 U6032 ( .A1(n7702), .A2(n7701), .ZN(n10412) );
  INV_X1 U6033 ( .A(n7578), .ZN(n10936) );
  NAND2_X1 U6034 ( .A1(n5633), .A2(n5637), .ZN(n9205) );
  OR2_X1 U6035 ( .A1(n5639), .A2(n5638), .ZN(n5633) );
  INV_X1 U6036 ( .A(n9172), .ZN(n5639) );
  NAND2_X1 U6037 ( .A1(n7956), .A2(n7955), .ZN(n10343) );
  NAND2_X1 U6038 ( .A1(n9312), .A2(n9307), .ZN(n9224) );
  NAND2_X1 U6039 ( .A1(n7974), .A2(n7973), .ZN(n10389) );
  AND2_X1 U6040 ( .A1(n5611), .A2(n5610), .ZN(n9235) );
  NAND2_X1 U6041 ( .A1(n7534), .A2(n7533), .ZN(n7773) );
  NOR2_X1 U6042 ( .A1(n5055), .A2(n5040), .ZN(n9253) );
  NAND2_X1 U6043 ( .A1(n5621), .A2(n8266), .ZN(n9263) );
  NAND2_X1 U6044 ( .A1(n5616), .A2(n5103), .ZN(n5621) );
  INV_X1 U6045 ( .A(n8267), .ZN(n5616) );
  AOI21_X1 U6046 ( .B1(n9205), .B2(n9203), .A(n5640), .ZN(n9276) );
  INV_X1 U6047 ( .A(n5104), .ZN(n5640) );
  NAND2_X1 U6048 ( .A1(n7964), .A2(n7963), .ZN(n10358) );
  AND4_X1 U6049 ( .A1(n7551), .A2(n7550), .A3(n7549), .A4(n7548), .ZN(n7853)
         );
  INV_X1 U6050 ( .A(n9314), .ZN(n9289) );
  NAND2_X1 U6051 ( .A1(n7980), .A2(n7979), .ZN(n10378) );
  INV_X1 U6052 ( .A(n9321), .ZN(n9292) );
  AND2_X1 U6053 ( .A1(n7027), .A2(n7026), .ZN(n9315) );
  NAND2_X1 U6054 ( .A1(n5230), .A2(n5236), .ZN(n9296) );
  NAND2_X1 U6055 ( .A1(n9216), .A2(n9213), .ZN(n5230) );
  NAND2_X1 U6056 ( .A1(n5235), .A2(n9213), .ZN(n9298) );
  OR2_X1 U6057 ( .A1(n9216), .A2(n9212), .ZN(n5235) );
  INV_X1 U6058 ( .A(n9220), .ZN(n9321) );
  NOR2_X1 U6059 ( .A1(n6936), .A2(n6933), .ZN(n9318) );
  INV_X1 U6060 ( .A(n6939), .ZN(n9600) );
  NAND2_X1 U6061 ( .A1(n5054), .A2(n5309), .ZN(n5161) );
  NAND2_X1 U6062 ( .A1(n9599), .A2(n7492), .ZN(n5307) );
  XNOR2_X1 U6063 ( .A(n6494), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9603) );
  NAND2_X1 U6064 ( .A1(n6498), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6494) );
  INV_X1 U6065 ( .A(n10111), .ZN(n9610) );
  INV_X1 U6066 ( .A(n10304), .ZN(n10276) );
  INV_X1 U6067 ( .A(n7853), .ZN(n10010) );
  INV_X1 U6068 ( .A(n7602), .ZN(n10012) );
  INV_X1 U6069 ( .A(n7428), .ZN(n10013) );
  INV_X1 U6070 ( .A(n7356), .ZN(n10844) );
  INV_X1 U6071 ( .A(P1_U4006), .ZN(n10671) );
  NOR2_X1 U6072 ( .A1(n10565), .A2(n10564), .ZN(n10562) );
  AOI21_X1 U6073 ( .B1(n10545), .B2(n5250), .A(n5248), .ZN(n6972) );
  INV_X1 U6074 ( .A(n5249), .ZN(n5248) );
  AOI21_X1 U6075 ( .B1(n5090), .B2(n5250), .A(n10563), .ZN(n5249) );
  NOR2_X1 U6076 ( .A1(n10041), .A2(n10042), .ZN(n10045) );
  AND2_X1 U6077 ( .A1(n9394), .A2(n9393), .ZN(n10322) );
  INV_X1 U6078 ( .A(n11047), .ZN(n8014) );
  NAND2_X1 U6079 ( .A1(n8493), .A2(n8492), .ZN(n5475) );
  INV_X1 U6080 ( .A(n8508), .ZN(n10331) );
  OAI21_X1 U6081 ( .B1(n10332), .B2(n10923), .A(n8507), .ZN(n8508) );
  AOI21_X1 U6082 ( .B1(n8506), .B2(n10920), .A(n8505), .ZN(n8507) );
  OAI21_X1 U6083 ( .B1(n10152), .B2(n5383), .A(n5379), .ZN(n10124) );
  NAND2_X1 U6084 ( .A1(n10142), .A2(n10143), .ZN(n10141) );
  NAND2_X1 U6085 ( .A1(n10161), .A2(n9481), .ZN(n10142) );
  NAND2_X1 U6086 ( .A1(n10152), .A2(n8458), .ZN(n10140) );
  NAND2_X1 U6087 ( .A1(n5174), .A2(n5384), .ZN(n10154) );
  NAND2_X1 U6088 ( .A1(n10186), .A2(n8455), .ZN(n10170) );
  NAND2_X1 U6089 ( .A1(n10190), .A2(n10191), .ZN(n10189) );
  NAND2_X1 U6090 ( .A1(n10202), .A2(n9359), .ZN(n10190) );
  NAND2_X1 U6091 ( .A1(n7985), .A2(n7984), .ZN(n10374) );
  INV_X1 U6092 ( .A(n5359), .ZN(n10268) );
  AOI21_X1 U6093 ( .B1(n10283), .B2(n10292), .A(n5362), .ZN(n5359) );
  AOI21_X1 U6094 ( .B1(n5467), .B2(n5038), .A(n5466), .ZN(n10291) );
  INV_X1 U6095 ( .A(n5453), .ZN(n7834) );
  AOI21_X1 U6096 ( .B1(n7850), .B2(n7748), .A(n5456), .ZN(n5453) );
  NAND2_X1 U6097 ( .A1(n7752), .A2(n7751), .ZN(n7886) );
  INV_X1 U6098 ( .A(n10935), .ZN(n10317) );
  XNOR2_X1 U6099 ( .A(n6489), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6839) );
  NAND2_X1 U6100 ( .A1(n9600), .A2(n6925), .ZN(n10467) );
  INV_X1 U6101 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6603) );
  XNOR2_X1 U6102 ( .A(n6185), .B(n6184), .ZN(n10451) );
  INV_X1 U6103 ( .A(n9595), .ZN(n7502) );
  NAND2_X1 U6104 ( .A1(n5563), .A2(n5561), .ZN(n6035) );
  NAND2_X1 U6105 ( .A1(n5551), .A2(n5549), .ZN(n5947) );
  NAND2_X1 U6106 ( .A1(n5551), .A2(n5714), .ZN(n5945) );
  OR2_X1 U6107 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  NAND2_X1 U6108 ( .A1(n5868), .A2(n5147), .ZN(n5146) );
  AND2_X1 U6109 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  NOR2_X1 U6110 ( .A1(n5872), .A2(n5148), .ZN(n5147) );
  NAND2_X1 U6111 ( .A1(n5858), .A2(n5868), .ZN(n7218) );
  NAND2_X1 U6112 ( .A1(n5847), .A2(n5846), .ZN(n7059) );
  INV_X1 U6113 ( .A(n5531), .ZN(n5810) );
  NAND2_X1 U6114 ( .A1(n6511), .A2(n5245), .ZN(n10607) );
  NOR2_X1 U6115 ( .A1(n7655), .A2(n7654), .ZN(n10500) );
  NOR2_X1 U6116 ( .A1(n10498), .A2(n10497), .ZN(n7654) );
  NAND2_X1 U6117 ( .A1(n5125), .A2(n5566), .ZN(P2_U3244) );
  OR2_X1 U6118 ( .A1(n8243), .A2(n8242), .ZN(n5566) );
  NAND2_X1 U6119 ( .A1(n5259), .A2(n5091), .ZN(n9114) );
  OR2_X1 U6120 ( .A1(n9034), .A2(n11030), .ZN(n5259) );
  OAI21_X1 U6121 ( .B1(n9034), .B2(n5266), .A(n5264), .ZN(P2_U3519) );
  NAND2_X1 U6122 ( .A1(n11041), .A2(n10865), .ZN(n5266) );
  INV_X1 U6123 ( .A(n5265), .ZN(n5264) );
  OAI21_X1 U6124 ( .B1(n5091), .B2(n11038), .A(n5267), .ZN(n5265) );
  NAND2_X1 U6125 ( .A1(n5229), .A2(n5227), .ZN(n9201) );
  AOI21_X1 U6126 ( .B1(n5254), .B2(n10687), .A(n5251), .ZN(n10083) );
  OAI211_X1 U6127 ( .C1(n10327), .C2(n10300), .A(n5474), .B(n5473), .ZN(
        P1_U3355) );
  NAND2_X1 U6128 ( .A1(n5475), .A2(n10942), .ZN(n5474) );
  AOI21_X1 U6129 ( .B1(n10324), .B2(n10932), .A(n8494), .ZN(n5473) );
  NOR2_X1 U6130 ( .A1(n10336), .A2(n10296), .ZN(n10105) );
  OAI21_X1 U6131 ( .B1(n5187), .B2(n11049), .A(n5321), .ZN(P1_U3552) );
  OR2_X1 U6132 ( .A1(n11050), .A2(n8467), .ZN(n5321) );
  INV_X1 U6133 ( .A(n10327), .ZN(n5322) );
  NAND2_X1 U6134 ( .A1(n11054), .A2(n11024), .ZN(n5371) );
  INV_X1 U6135 ( .A(n5370), .ZN(n5369) );
  NAND2_X1 U6136 ( .A1(n5364), .A2(n11054), .ZN(n5363) );
  AND2_X1 U6137 ( .A1(n6339), .A2(n6340), .ZN(n5036) );
  NAND2_X2 U6138 ( .A1(n6071), .A2(n6216), .ZN(n6223) );
  OAI211_X1 U6139 ( .C1(n6634), .C2(n10637), .A(n5787), .B(n5788), .ZN(n6692)
         );
  CLKBUF_X3 U6140 ( .A(n5901), .Z(n5919) );
  AND4_X1 U6141 ( .A1(n5753), .A2(n5755), .A3(n5756), .A4(n5754), .ZN(n5037)
         );
  AND2_X1 U6142 ( .A1(n10307), .A2(n9523), .ZN(n5038) );
  NOR2_X1 U6143 ( .A1(n5998), .A2(n5289), .ZN(n5288) );
  AND2_X1 U6144 ( .A1(n6046), .A2(n8964), .ZN(n5039) );
  OR2_X1 U6145 ( .A1(n10333), .A2(n10111), .ZN(n9473) );
  INV_X1 U6146 ( .A(n9429), .ZN(n5452) );
  AND2_X1 U6147 ( .A1(n8339), .A2(n8338), .ZN(n5040) );
  AND2_X1 U6148 ( .A1(n6607), .A2(n10447), .ZN(n7421) );
  INV_X1 U6149 ( .A(n7016), .ZN(n7239) );
  AND2_X1 U6150 ( .A1(n5039), .A2(n6079), .ZN(n5041) );
  AND4_X1 U6151 ( .A1(n10112), .A2(n10134), .A3(n10163), .A4(n9446), .ZN(n5042) );
  NOR2_X1 U6152 ( .A1(n9401), .A2(n5457), .ZN(n5043) );
  AND2_X1 U6153 ( .A1(n9527), .A2(n9523), .ZN(n9440) );
  OR2_X1 U6154 ( .A1(n8236), .A2(n6350), .ZN(n5044) );
  INV_X1 U6155 ( .A(n9444), .ZN(n10206) );
  AND3_X1 U6156 ( .A1(n10178), .A2(n9570), .A3(n9569), .ZN(n5045) );
  INV_X1 U6157 ( .A(n5092), .ZN(n5286) );
  INV_X1 U6158 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U6159 ( .A1(n8052), .A2(n8051), .ZN(n8054) );
  INV_X1 U6160 ( .A(n8054), .ZN(n5348) );
  INV_X1 U6161 ( .A(n5491), .ZN(n5490) );
  NAND2_X1 U6162 ( .A1(n8207), .A2(n5985), .ZN(n5491) );
  NAND2_X1 U6163 ( .A1(n10865), .A2(n6223), .ZN(n6350) );
  INV_X1 U6164 ( .A(n10564), .ZN(n5250) );
  NAND2_X1 U6165 ( .A1(n6191), .A2(n6190), .ZN(n9041) );
  INV_X1 U6166 ( .A(n5518), .ZN(n6052) );
  INV_X1 U6167 ( .A(n7737), .ZN(n5276) );
  OR2_X1 U6168 ( .A1(n9747), .A2(n5108), .ZN(n5046) );
  INV_X1 U6169 ( .A(n5034), .ZN(n8356) );
  OR2_X1 U6170 ( .A1(n10316), .A2(n9533), .ZN(n9528) );
  NOR2_X1 U6171 ( .A1(n5142), .A2(n5141), .ZN(n6218) );
  INV_X1 U6172 ( .A(n9603), .ZN(n6889) );
  INV_X1 U6173 ( .A(n7463), .ZN(n5269) );
  INV_X1 U6174 ( .A(n10292), .ZN(n5465) );
  INV_X1 U6175 ( .A(n9038), .ZN(n8784) );
  NAND2_X1 U6176 ( .A1(n8038), .A2(n8037), .ZN(n9038) );
  NOR2_X1 U6177 ( .A1(n10838), .A2(n7529), .ZN(n5047) );
  NAND2_X1 U6178 ( .A1(n5765), .A2(n5764), .ZN(n9079) );
  AND2_X1 U6179 ( .A1(n6241), .A2(n6239), .ZN(n5048) );
  AND2_X1 U6180 ( .A1(n8192), .A2(n8086), .ZN(n5049) );
  AND2_X1 U6181 ( .A1(n6525), .A2(n6467), .ZN(n6522) );
  NAND2_X2 U6182 ( .A1(n6895), .A2(n8021), .ZN(n7060) );
  NAND3_X1 U6183 ( .A1(n6525), .A2(n5652), .A3(n6473), .ZN(n5050) );
  NAND2_X1 U6184 ( .A1(n5888), .A2(n5887), .ZN(n10895) );
  INV_X1 U6185 ( .A(n10895), .ZN(n5151) );
  AND2_X1 U6186 ( .A1(n10663), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5051) );
  AND4_X1 U6187 ( .A1(n5757), .A2(n5961), .A3(n5960), .A4(n6016), .ZN(n5052)
         );
  INV_X1 U6188 ( .A(n5815), .ZN(n5816) );
  INV_X1 U6189 ( .A(n8227), .ZN(n8034) );
  XNOR2_X1 U6190 ( .A(n6220), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8227) );
  AND2_X1 U6191 ( .A1(n9251), .A2(n8351), .ZN(n5053) );
  AND3_X1 U6192 ( .A1(n9597), .A2(n9598), .A3(n5308), .ZN(n5054) );
  AND4_X1 U6193 ( .A1(n6473), .A2(n6525), .A3(n5472), .A4(n5468), .ZN(n6479)
         );
  INV_X1 U6194 ( .A(n8266), .ZN(n5619) );
  NAND2_X1 U6195 ( .A1(n6123), .A2(n5312), .ZN(n6141) );
  AND2_X1 U6196 ( .A1(n9172), .A2(n9173), .ZN(n5055) );
  AND3_X1 U6197 ( .A1(n9585), .A2(n9586), .A3(n9587), .ZN(n5056) );
  NAND2_X1 U6198 ( .A1(n5215), .A2(n6510), .ZN(n6514) );
  AND3_X1 U6199 ( .A1(n5838), .A2(n5839), .A3(n5837), .ZN(n5057) );
  AND2_X1 U6200 ( .A1(n8138), .A2(n8141), .ZN(n8933) );
  AND3_X1 U6201 ( .A1(n9554), .A2(n10248), .A3(n9553), .ZN(n5058) );
  AND2_X1 U6202 ( .A1(n9479), .A2(n9478), .ZN(n10143) );
  NAND2_X1 U6203 ( .A1(n5806), .A2(n5564), .ZN(n5840) );
  NAND2_X1 U6204 ( .A1(n6510), .A2(n6463), .ZN(n6505) );
  AND2_X1 U6205 ( .A1(n10358), .A2(n10192), .ZN(n5059) );
  NAND4_X1 U6206 ( .A1(n6473), .A2(n6525), .A3(n5472), .A4(n5471), .ZN(n5060)
         );
  AND2_X1 U6207 ( .A1(n6426), .A2(n6425), .ZN(n5061) );
  AND2_X1 U6208 ( .A1(n6389), .A2(n6388), .ZN(n5062) );
  NAND2_X1 U6209 ( .A1(n7746), .A2(n7745), .ZN(n10406) );
  INV_X1 U6210 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10439) );
  NAND2_X1 U6211 ( .A1(n7992), .A2(n7991), .ZN(n10364) );
  INV_X1 U6212 ( .A(n9225), .ZN(n5608) );
  AND2_X1 U6213 ( .A1(n8866), .A2(n5476), .ZN(n5063) );
  OR2_X1 U6214 ( .A1(n10736), .A2(n8382), .ZN(n5064) );
  NAND2_X1 U6215 ( .A1(n8885), .A2(n5272), .ZN(n5273) );
  NAND2_X1 U6216 ( .A1(n10211), .A2(n5319), .ZN(n5320) );
  NAND2_X1 U6217 ( .A1(n7960), .A2(n7959), .ZN(n10353) );
  INV_X1 U6218 ( .A(n7346), .ZN(n7344) );
  AND2_X1 U6219 ( .A1(n8863), .A2(n8164), .ZN(n5065) );
  INV_X1 U6220 ( .A(n5288), .ZN(n5287) );
  NAND2_X1 U6221 ( .A1(n6083), .A2(n6082), .ZN(n9084) );
  OR2_X1 U6222 ( .A1(n6634), .A2(n6670), .ZN(n5066) );
  NOR2_X1 U6223 ( .A1(n7908), .A2(n8659), .ZN(n5067) );
  INV_X1 U6224 ( .A(n5644), .ZN(n5638) );
  AND2_X1 U6225 ( .A1(n5645), .A2(n9173), .ZN(n5644) );
  OR2_X1 U6226 ( .A1(n5620), .A2(n5614), .ZN(n5068) );
  OR2_X1 U6227 ( .A1(n5620), .A2(n5615), .ZN(n5069) );
  AND2_X1 U6228 ( .A1(n9572), .A2(n10143), .ZN(n5070) );
  AND2_X1 U6229 ( .A1(n5565), .A2(n5127), .ZN(n5071) );
  OR2_X1 U6230 ( .A1(n8172), .A2(n8168), .ZN(n5072) );
  AND2_X1 U6231 ( .A1(n9473), .A2(n9474), .ZN(n10098) );
  INV_X1 U6232 ( .A(n10098), .ZN(n5184) );
  AND2_X1 U6233 ( .A1(n6314), .A2(n6313), .ZN(n5073) );
  NAND2_X1 U6234 ( .A1(n8097), .A2(n8098), .ZN(n8206) );
  AND2_X1 U6235 ( .A1(n6409), .A2(n6408), .ZN(n5074) );
  AND2_X1 U6236 ( .A1(n5730), .A2(n5729), .ZN(n5075) );
  INV_X1 U6237 ( .A(n8866), .ZN(n6246) );
  NAND2_X1 U6238 ( .A1(n8164), .A2(n8158), .ZN(n8866) );
  NOR2_X1 U6239 ( .A1(n5717), .A2(SI_12_), .ZN(n5076) );
  INV_X1 U6240 ( .A(n5380), .ZN(n5379) );
  NAND2_X1 U6241 ( .A1(n8460), .A2(n5381), .ZN(n5380) );
  OR2_X1 U6242 ( .A1(n9260), .A2(n5619), .ZN(n5077) );
  INV_X1 U6243 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9131) );
  OR2_X1 U6244 ( .A1(n5184), .A2(n9385), .ZN(n5078) );
  NAND2_X1 U6245 ( .A1(n5973), .A2(n5304), .ZN(n5079) );
  AND2_X1 U6246 ( .A1(n9480), .A2(n9481), .ZN(n10163) );
  INV_X1 U6247 ( .A(n10163), .ZN(n5177) );
  INV_X1 U6248 ( .A(n5464), .ZN(n5463) );
  OR2_X1 U6249 ( .A1(n5053), .A2(n5040), .ZN(n5080) );
  INV_X1 U6250 ( .A(n5524), .ZN(n5523) );
  AND2_X1 U6251 ( .A1(n6017), .A2(n5525), .ZN(n5524) );
  NAND2_X1 U6252 ( .A1(n9466), .A2(n9468), .ZN(n9447) );
  INV_X1 U6253 ( .A(n9447), .ZN(n9581) );
  NAND2_X1 U6254 ( .A1(n8175), .A2(n8174), .ZN(n8821) );
  INV_X1 U6255 ( .A(n8821), .ZN(n8813) );
  AND2_X1 U6256 ( .A1(n5305), .A2(n5304), .ZN(n5081) );
  AND2_X1 U6257 ( .A1(n5191), .A2(n8603), .ZN(n5082) );
  AND2_X1 U6258 ( .A1(n8798), .A2(n8176), .ZN(n5083) );
  AND2_X1 U6259 ( .A1(n5642), .A2(n5644), .ZN(n5084) );
  AND2_X1 U6260 ( .A1(n9032), .A2(n9038), .ZN(n5085) );
  INV_X1 U6261 ( .A(n8164), .ZN(n5580) );
  OR2_X1 U6262 ( .A1(n9062), .A2(n8568), .ZN(n8164) );
  AND2_X1 U6263 ( .A1(n8210), .A2(n8114), .ZN(n5086) );
  AND2_X1 U6264 ( .A1(n9503), .A2(n9502), .ZN(n5087) );
  NAND2_X1 U6265 ( .A1(n5139), .A2(n5606), .ZN(n5766) );
  INV_X1 U6266 ( .A(n5766), .ZN(n5767) );
  AND2_X1 U6267 ( .A1(n8150), .A2(n8916), .ZN(n5088) );
  AND2_X1 U6268 ( .A1(n5562), .A2(n5733), .ZN(n5561) );
  INV_X1 U6269 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5225) );
  INV_X1 U6270 ( .A(n8876), .ZN(n8882) );
  NAND2_X1 U6271 ( .A1(n8157), .A2(n8154), .ZN(n8876) );
  NAND2_X1 U6272 ( .A1(n8187), .A2(n8186), .ZN(n5089) );
  INV_X1 U6273 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U6274 ( .A1(n7902), .A2(n8112), .ZN(n7939) );
  AND2_X1 U6275 ( .A1(n10550), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5090) );
  AND2_X1 U6276 ( .A1(n9033), .A2(n9036), .ZN(n5091) );
  AND4_X1 U6277 ( .A1(n6115), .A2(n6114), .A3(n6113), .A4(n6112), .ZN(n8860)
         );
  INV_X1 U6278 ( .A(n8860), .ZN(n5536) );
  INV_X1 U6279 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5496) );
  OAI21_X1 U6280 ( .B1(n5974), .B2(n5519), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6066) );
  AND2_X1 U6281 ( .A1(n5727), .A2(n5726), .ZN(n5092) );
  NAND2_X1 U6282 ( .A1(n6054), .A2(n6053), .ZN(n9094) );
  NAND2_X1 U6283 ( .A1(n6074), .A2(n6073), .ZN(n9091) );
  AND2_X1 U6284 ( .A1(n8223), .A2(n8225), .ZN(n8217) );
  NAND2_X1 U6285 ( .A1(n7786), .A2(n7776), .ZN(n7824) );
  AND2_X1 U6286 ( .A1(n9369), .A2(n9484), .ZN(n10191) );
  INV_X1 U6287 ( .A(n10191), .ZN(n5444) );
  NAND2_X1 U6288 ( .A1(n9603), .A2(n9595), .ZN(n6871) );
  AND2_X1 U6289 ( .A1(n8145), .A2(n8150), .ZN(n8899) );
  INV_X1 U6290 ( .A(n8899), .ZN(n5585) );
  OR2_X1 U6291 ( .A1(n10406), .A2(n7880), .ZN(n9517) );
  INV_X1 U6292 ( .A(n9517), .ZN(n5456) );
  NAND2_X1 U6293 ( .A1(n6130), .A2(n6129), .ZN(n9062) );
  NOR2_X1 U6294 ( .A1(n5974), .A2(n5522), .ZN(n5518) );
  INV_X1 U6295 ( .A(n8819), .ZN(n9046) );
  AND2_X1 U6296 ( .A1(n6174), .A2(n6173), .ZN(n8819) );
  NAND2_X1 U6297 ( .A1(n8982), .A2(n5041), .ZN(n5275) );
  AND2_X1 U6298 ( .A1(n8945), .A2(n8129), .ZN(n5093) );
  AND2_X1 U6299 ( .A1(n10389), .A2(n10294), .ZN(n5094) );
  INV_X1 U6300 ( .A(n8893), .ZN(n8911) );
  NOR2_X1 U6301 ( .A1(n8927), .A2(n9079), .ZN(n8893) );
  AND2_X1 U6302 ( .A1(n5271), .A2(n8819), .ZN(n5095) );
  NOR2_X1 U6303 ( .A1(n7837), .A2(n7836), .ZN(n8478) );
  INV_X1 U6304 ( .A(n8478), .ZN(n5467) );
  INV_X1 U6305 ( .A(n5375), .ZN(n5374) );
  NOR2_X1 U6306 ( .A1(n8512), .A2(n9188), .ZN(n5375) );
  AND4_X1 U6307 ( .A1(n6198), .A2(n6197), .A3(n6196), .A4(n6195), .ZN(n8823)
         );
  INV_X1 U6308 ( .A(n8823), .ZN(n8654) );
  AND2_X1 U6309 ( .A1(n9638), .A2(keyinput_133), .ZN(n5096) );
  AND2_X1 U6310 ( .A1(n8803), .A2(n8823), .ZN(n5097) );
  AND2_X1 U6311 ( .A1(n5745), .A2(n5744), .ZN(n5098) );
  INV_X1 U6312 ( .A(n5477), .ZN(n9073) );
  OR2_X1 U6313 ( .A1(n8883), .A2(n8882), .ZN(n5477) );
  NAND2_X1 U6314 ( .A1(n5556), .A2(n6090), .ZN(n5555) );
  INV_X1 U6315 ( .A(n5511), .ZN(n5205) );
  AND2_X1 U6316 ( .A1(n8520), .A2(n5512), .ZN(n5511) );
  NAND2_X1 U6317 ( .A1(n7996), .A2(n7995), .ZN(n10349) );
  INV_X1 U6318 ( .A(n10349), .ZN(n5316) );
  AND2_X1 U6319 ( .A1(n6240), .A2(n6239), .ZN(n5099) );
  NAND2_X1 U6320 ( .A1(n6159), .A2(n6158), .ZN(n9052) );
  INV_X1 U6321 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U6322 ( .A1(n7320), .A2(n5507), .ZN(n5506) );
  XNOR2_X1 U6323 ( .A(n5515), .B(n6217), .ZN(n6227) );
  AND2_X2 U6324 ( .A1(n6457), .A2(n7152), .ZN(n11041) );
  NAND2_X1 U6325 ( .A1(n7374), .A2(n7373), .ZN(n7375) );
  AND3_X2 U6326 ( .A1(n7481), .A2(n7480), .A3(n7479), .ZN(n11050) );
  INV_X1 U6327 ( .A(n9402), .ZN(n5457) );
  NAND2_X1 U6328 ( .A1(n7057), .A2(n7056), .ZN(n7231) );
  AND2_X1 U6329 ( .A1(n10035), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5100) );
  INV_X1 U6330 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5152) );
  AND2_X1 U6331 ( .A1(n5626), .A2(n7709), .ZN(n5101) );
  NAND2_X1 U6332 ( .A1(n7612), .A2(n5136), .ZN(n7731) );
  NAND2_X1 U6333 ( .A1(n5646), .A2(n7329), .ZN(n7343) );
  OR2_X1 U6334 ( .A1(n7789), .A2(n5326), .ZN(n5102) );
  NAND2_X1 U6335 ( .A1(n5760), .A2(n6221), .ZN(n6269) );
  INV_X1 U6336 ( .A(n5314), .ZN(n10833) );
  NOR2_X1 U6337 ( .A1(n7299), .A2(n7483), .ZN(n5314) );
  NAND2_X1 U6338 ( .A1(n5623), .A2(n5622), .ZN(n7808) );
  OR2_X1 U6339 ( .A1(n7386), .A2(n8077), .ZN(n7402) );
  INV_X1 U6340 ( .A(n7402), .ZN(n5277) );
  NAND2_X1 U6341 ( .A1(n7875), .A2(n7876), .ZN(n5103) );
  NAND2_X1 U6342 ( .A1(n8365), .A2(n8364), .ZN(n5104) );
  OR2_X1 U6343 ( .A1(n9715), .A2(keyinput_183), .ZN(n5105) );
  AND2_X1 U6344 ( .A1(n7329), .A2(n7344), .ZN(n5106) );
  AND2_X1 U6345 ( .A1(n11014), .A2(n5985), .ZN(n5107) );
  NOR2_X1 U6346 ( .A1(n8241), .A2(n8227), .ZN(n8189) );
  INV_X1 U6347 ( .A(n8189), .ZN(n5213) );
  INV_X1 U6348 ( .A(n10865), .ZN(n11030) );
  NAND4_X1 U6349 ( .A1(n5821), .A2(n5820), .A3(n5819), .A4(n5818), .ZN(n6592)
         );
  AND2_X1 U6350 ( .A1(n10923), .A2(n10707), .ZN(n10415) );
  AND2_X1 U6351 ( .A1(keyinput_207), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n5108)
         );
  AND2_X1 U6352 ( .A1(n8540), .A2(n6311), .ZN(n5109) );
  NAND2_X1 U6353 ( .A1(n5353), .A2(n5257), .ZN(n9140) );
  XNOR2_X1 U6354 ( .A(n6843), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9598) );
  INV_X1 U6355 ( .A(n9598), .ZN(n7492) );
  INV_X1 U6356 ( .A(n10229), .ZN(n10730) );
  XOR2_X1 U6357 ( .A(n10730), .B(P1_REG2_REG_19__SCAN_IN), .Z(n5110) );
  NOR2_X1 U6358 ( .A1(n5769), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n9130) );
  NOR2_X1 U6359 ( .A1(n6602), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n10438) );
  OR2_X1 U6360 ( .A1(n9772), .A2(n9773), .ZN(n5111) );
  AND2_X1 U6361 ( .A1(n9776), .A2(n9777), .ZN(n5112) );
  INV_X1 U6362 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5214) );
  INV_X1 U6363 ( .A(n10808), .ZN(n8932) );
  NAND3_X1 U6364 ( .A1(n5116), .A2(n5115), .A3(n8094), .ZN(n7727) );
  NAND4_X1 U6365 ( .A1(n5116), .A2(n8098), .A3(n5115), .A4(n8094), .ZN(n5114)
         );
  NAND3_X1 U6366 ( .A1(n5119), .A2(n5533), .A3(n5118), .ZN(n5532) );
  AND2_X2 U6367 ( .A1(n5119), .A2(n5118), .ZN(n8021) );
  NAND3_X1 U6368 ( .A1(n5356), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5118) );
  NAND3_X1 U6369 ( .A1(n5122), .A2(n5124), .A3(n5123), .ZN(n5119) );
  NAND2_X1 U6370 ( .A1(n5126), .A2(n6584), .ZN(n5125) );
  NAND3_X1 U6371 ( .A1(n5128), .A2(n5071), .A3(n5044), .ZN(n5126) );
  INV_X1 U6372 ( .A(n8238), .ZN(n5127) );
  NAND2_X1 U6373 ( .A1(n5568), .A2(n5567), .ZN(n5128) );
  NAND2_X1 U6374 ( .A1(n5130), .A2(n5943), .ZN(n7614) );
  NAND2_X1 U6375 ( .A1(n7504), .A2(n5130), .ZN(n10978) );
  AOI21_X2 U6376 ( .B1(n8799), .B2(n8805), .A(n5097), .ZN(n5137) );
  NAND4_X1 U6377 ( .A1(n5873), .A2(n5037), .A3(n5138), .A4(n5052), .ZN(n5140)
         );
  NAND2_X1 U6378 ( .A1(n5037), .A2(n5873), .ZN(n5142) );
  INV_X1 U6379 ( .A(n5140), .ZN(n5139) );
  AOI21_X2 U6380 ( .B1(n8956), .B2(n8212), .A(n5662), .ZN(n8944) );
  NAND2_X1 U6381 ( .A1(n7462), .A2(n8049), .ZN(n7461) );
  AND2_X1 U6382 ( .A1(n5799), .A2(n5143), .ZN(n7462) );
  AND2_X2 U6383 ( .A1(n6230), .A2(n6690), .ZN(n6686) );
  NOR2_X1 U6384 ( .A1(n9130), .A2(n9131), .ZN(n5144) );
  NAND2_X2 U6385 ( .A1(n10802), .A2(n10805), .ZN(n9021) );
  OAI22_X1 U6386 ( .A1(n8892), .A2(n8899), .B1(n9074), .B2(n8918), .ZN(n8883)
         );
  OAI21_X1 U6387 ( .B1(n8926), .B2(n5479), .A(n5478), .ZN(n5482) );
  OAI21_X1 U6388 ( .B1(n5984), .B2(n5491), .A(n5489), .ZN(n7944) );
  NAND2_X1 U6389 ( .A1(n7401), .A2(n7400), .ZN(n7399) );
  NAND4_X1 U6390 ( .A1(n5796), .A2(n5795), .A3(n5797), .A4(n5794), .ZN(n6230)
         );
  INV_X1 U6391 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U6392 ( .A1(n7250), .A2(n5850), .ZN(n10802) );
  INV_X4 U6393 ( .A(n5862), .ZN(n6131) );
  NAND2_X1 U6394 ( .A1(n7614), .A2(n7613), .ZN(n7612) );
  NAND2_X1 U6395 ( .A1(n10784), .A2(n8542), .ZN(n8057) );
  NAND2_X1 U6396 ( .A1(n5847), .A2(n5685), .ZN(n5857) );
  INV_X1 U6397 ( .A(n5154), .ZN(n5153) );
  NAND3_X1 U6398 ( .A1(n5149), .A2(n8135), .A3(n5352), .ZN(n8139) );
  OAI21_X1 U6399 ( .B1(n5654), .B2(n8127), .A(n8186), .ZN(n5149) );
  OAI21_X1 U6400 ( .B1(n5538), .B2(n8167), .A(n5539), .ZN(n8171) );
  NAND2_X1 U6401 ( .A1(n5163), .A2(n5330), .ZN(n8165) );
  NAND2_X1 U6402 ( .A1(n5166), .A2(n5089), .ZN(n8222) );
  XNOR2_X1 U6403 ( .A(n8190), .B(n5542), .ZN(n5329) );
  NAND2_X1 U6404 ( .A1(n5338), .A2(n5083), .ZN(n8179) );
  OAI211_X1 U6405 ( .C1(n8021), .C2(P2_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n5532), .ZN(n5672) );
  OAI21_X1 U6406 ( .B1(n5895), .B2(n5487), .A(n5485), .ZN(n5154) );
  NAND2_X1 U6407 ( .A1(n5781), .A2(n5782), .ZN(n5786) );
  NAND2_X1 U6408 ( .A1(n7251), .A2(n7253), .ZN(n7250) );
  INV_X1 U6409 ( .A(n5896), .ZN(n5487) );
  NAND2_X1 U6410 ( .A1(n5828), .A2(n5829), .ZN(n7003) );
  NAND2_X1 U6411 ( .A1(n5884), .A2(n5883), .ZN(n7413) );
  NAND2_X1 U6412 ( .A1(n5670), .A2(SI_1_), .ZN(n5674) );
  NAND2_X1 U6413 ( .A1(n5156), .A2(n9509), .ZN(n9513) );
  OAI21_X1 U6414 ( .B1(n9505), .B2(n9504), .A(n5087), .ZN(n5156) );
  OAI21_X1 U6415 ( .B1(n5058), .B2(n5157), .A(n9562), .ZN(n9563) );
  NAND2_X1 U6416 ( .A1(n9557), .A2(n9558), .ZN(n5157) );
  NAND2_X1 U6417 ( .A1(n5159), .A2(n5158), .ZN(n9569) );
  NAND2_X1 U6418 ( .A1(n9568), .A2(n9567), .ZN(n5159) );
  NAND2_X2 U6419 ( .A1(n7138), .A2(n9339), .ZN(n9400) );
  AOI21_X2 U6420 ( .B1(n9584), .B2(n5056), .A(n5160), .ZN(n9593) );
  OR4_X2 U6421 ( .A1(n9545), .A2(n9544), .A3(n10292), .A4(n9543), .ZN(n9550)
         );
  NAND2_X1 U6422 ( .A1(n5161), .A2(n5307), .ZN(n9606) );
  NOR2_X2 U6423 ( .A1(n5162), .A2(n6472), .ZN(n6473) );
  NAND4_X1 U6424 ( .A1(n6469), .A2(n6470), .A3(n6471), .A4(n6468), .ZN(n5162)
         );
  NAND3_X1 U6425 ( .A1(n8143), .A2(n5333), .A3(n5088), .ZN(n5163) );
  NAND2_X1 U6426 ( .A1(n5164), .A2(n8118), .ZN(n8122) );
  NAND2_X1 U6427 ( .A1(n8115), .A2(n5086), .ZN(n5164) );
  OR3_X1 U6428 ( .A1(n8943), .A2(n8134), .A3(n8133), .ZN(n8135) );
  INV_X1 U6429 ( .A(n8222), .ZN(n8190) );
  INV_X1 U6430 ( .A(n8139), .ZN(n8142) );
  NAND2_X1 U6431 ( .A1(n5544), .A2(n5543), .ZN(n5166) );
  OAI211_X1 U6432 ( .C1(n5342), .C2(n5341), .A(n5339), .B(n8813), .ZN(n5338)
         );
  NAND2_X1 U6433 ( .A1(n5684), .A2(n5683), .ZN(n5165) );
  AND3_X1 U6434 ( .A1(n8128), .A2(n8129), .A3(n9094), .ZN(n5654) );
  NAND2_X1 U6435 ( .A1(n5786), .A2(n5674), .ZN(n5531) );
  AND2_X2 U6436 ( .A1(n8499), .A2(n5771), .ZN(n5793) );
  NAND2_X1 U6437 ( .A1(n8105), .A2(n5344), .ZN(n8111) );
  AOI21_X1 U6438 ( .B1(n8171), .B2(n8170), .A(n5343), .ZN(n5342) );
  NAND2_X1 U6439 ( .A1(n10235), .A2(n10241), .ZN(n5167) );
  NAND2_X1 U6440 ( .A1(n10253), .A2(n8448), .ZN(n5168) );
  OAI21_X1 U6441 ( .B1(n8462), .B2(n5183), .A(n5179), .ZN(n8500) );
  NAND2_X1 U6442 ( .A1(n8462), .A2(n8461), .ZN(n10113) );
  NAND2_X1 U6443 ( .A1(n5189), .A2(n5082), .ZN(n6395) );
  NAND2_X1 U6444 ( .A1(n6386), .A2(n5192), .ZN(n5189) );
  NAND2_X1 U6445 ( .A1(n6386), .A2(n8622), .ZN(n8549) );
  INV_X1 U6446 ( .A(n8548), .ZN(n5194) );
  NAND2_X1 U6447 ( .A1(n6419), .A2(n5196), .ZN(n5195) );
  OAI211_X1 U6448 ( .C1(n6419), .C2(n5201), .A(n5197), .B(n5195), .ZN(n6437)
         );
  NAND2_X1 U6449 ( .A1(n8574), .A2(n5516), .ZN(n6381) );
  NAND2_X1 U6450 ( .A1(n8642), .A2(n8643), .ZN(n8641) );
  NAND2_X1 U6451 ( .A1(n5206), .A2(n5207), .ZN(n10796) );
  AOI21_X1 U6452 ( .B1(n5530), .B2(n8538), .A(n5073), .ZN(n5206) );
  NAND2_X1 U6453 ( .A1(n8539), .A2(n5530), .ZN(n5207) );
  NAND2_X1 U6454 ( .A1(n8540), .A2(n5530), .ZN(n6820) );
  NAND2_X1 U6455 ( .A1(n5208), .A2(n6310), .ZN(n8540) );
  NOR2_X4 U6456 ( .A1(n6514), .A2(n6466), .ZN(n6525) );
  XNOR2_X1 U6457 ( .A(n7053), .B(n7055), .ZN(n7051) );
  NAND2_X1 U6458 ( .A1(n7237), .A2(n5223), .ZN(n5219) );
  NAND4_X1 U6459 ( .A1(n5220), .A2(n5219), .A3(n5218), .A4(n7448), .ZN(n7574)
         );
  OR2_X1 U6460 ( .A1(n9216), .A2(n5234), .ZN(n5229) );
  NAND2_X1 U6461 ( .A1(n5239), .A2(n5240), .ZN(n8323) );
  NAND3_X1 U6462 ( .A1(n9312), .A2(n9307), .A3(n5244), .ZN(n5239) );
  NAND3_X1 U6463 ( .A1(n9312), .A2(n9307), .A3(n5608), .ZN(n5611) );
  NOR2_X1 U6464 ( .A1(n8323), .A2(n8322), .ZN(n9284) );
  MUX2_X1 U6465 ( .A(n6509), .B(P1_IR_REG_31__SCAN_IN), .S(n6508), .Z(n5245)
         );
  INV_X1 U6466 ( .A(n5247), .ZN(n10019) );
  AOI21_X1 U6467 ( .B1(n8781), .B2(n5261), .A(n5085), .ZN(n5260) );
  NAND2_X1 U6468 ( .A1(n8781), .A2(n8784), .ZN(n8783) );
  OR2_X1 U6469 ( .A1(n11041), .A2(n5268), .ZN(n5267) );
  INV_X1 U6470 ( .A(n5273), .ZN(n8847) );
  INV_X1 U6471 ( .A(n5275), .ZN(n8950) );
  OAI21_X1 U6472 ( .B1(n5986), .B2(n5282), .A(n5280), .ZN(n6049) );
  NAND2_X1 U6473 ( .A1(n6064), .A2(n5292), .ZN(n5291) );
  NAND3_X1 U6474 ( .A1(n9459), .A2(n9448), .A3(n5297), .ZN(n9451) );
  NAND3_X1 U6475 ( .A1(n9581), .A2(n10098), .A3(n5042), .ZN(n5298) );
  OAI21_X1 U6476 ( .B1(n5929), .B2(n5302), .A(n5300), .ZN(n5722) );
  OAI21_X1 U6477 ( .B1(n5929), .B2(n5548), .A(n5545), .ZN(n5306) );
  NAND3_X1 U6478 ( .A1(n9453), .A2(n9454), .A3(n10229), .ZN(n5308) );
  NAND2_X1 U6479 ( .A1(n6141), .A2(n6140), .ZN(n6153) );
  NAND2_X1 U6480 ( .A1(n6141), .A2(n5310), .ZN(n6157) );
  NAND2_X1 U6481 ( .A1(n6123), .A2(n6122), .ZN(n6126) );
  NOR2_X2 U6482 ( .A1(n10090), .A2(n10328), .ZN(n8509) );
  NOR2_X2 U6483 ( .A1(n10125), .A2(n10338), .ZN(n10117) );
  NOR2_X2 U6484 ( .A1(n10834), .A2(n7450), .ZN(n10910) );
  AND2_X2 U6485 ( .A1(n10211), .A2(n5315), .ZN(n10146) );
  INV_X1 U6486 ( .A(n5320), .ZN(n10171) );
  INV_X1 U6487 ( .A(n5324), .ZN(n10311) );
  XNOR2_X2 U6488 ( .A(n5328), .B(n6483), .ZN(n10510) );
  OAI21_X2 U6489 ( .B1(n6484), .B2(n6476), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5328) );
  INV_X2 U6490 ( .A(n10713), .ZN(n10726) );
  NOR2_X2 U6491 ( .A1(n9341), .A2(n10710), .ZN(n7209) );
  INV_X1 U6492 ( .A(n5331), .ZN(n5330) );
  NOR2_X1 U6493 ( .A1(n8153), .A2(n8152), .ZN(n5337) );
  OAI21_X1 U6494 ( .B1(n8171), .B2(n5072), .A(n5340), .ZN(n5339) );
  NAND3_X1 U6495 ( .A1(n5350), .A2(n5349), .A3(n5348), .ZN(n5347) );
  NAND3_X1 U6496 ( .A1(n8132), .A2(n8155), .A3(n8131), .ZN(n5352) );
  NAND2_X2 U6497 ( .A1(n6253), .A2(n9140), .ZN(n6634) );
  AND3_X2 U6498 ( .A1(n5806), .A2(n5564), .A3(n5355), .ZN(n5873) );
  NAND2_X1 U6499 ( .A1(n10283), .A2(n5360), .ZN(n5357) );
  NAND2_X1 U6500 ( .A1(n5357), .A2(n5358), .ZN(n10253) );
  INV_X1 U6501 ( .A(n10325), .ZN(n5364) );
  OAI211_X1 U6502 ( .C1(n10327), .C2(n5371), .A(n5363), .B(n5369), .ZN(
        P1_U3520) );
  NAND2_X1 U6503 ( .A1(n5376), .A2(n5377), .ZN(n8462) );
  NAND3_X1 U6504 ( .A1(n9630), .A2(n5394), .A3(n5391), .ZN(n5390) );
  AOI211_X1 U6505 ( .C1(n9757), .C2(n9756), .A(n9755), .B(n9754), .ZN(n9764)
         );
  OR2_X1 U6506 ( .A1(n9705), .A2(n5655), .ZN(n9706) );
  AOI21_X1 U6507 ( .B1(n9653), .B2(n9652), .A(n9651), .ZN(n9654) );
  AOI22_X1 U6508 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_178), .B1(n9707), 
        .B2(n9706), .ZN(n9708) );
  NAND2_X1 U6509 ( .A1(n8133), .A2(n8134), .ZN(n8128) );
  NAND2_X1 U6510 ( .A1(n8185), .A2(n8231), .ZN(n5544) );
  NAND2_X1 U6511 ( .A1(n5563), .A2(n5733), .ZN(n6033) );
  NOR2_X1 U6512 ( .A1(n8166), .A2(n5540), .ZN(n5538) );
  OAI21_X1 U6513 ( .B1(n8142), .B2(n8141), .A(n8140), .ZN(n8143) );
  NOR3_X1 U6514 ( .A1(n9666), .A2(n9665), .A3(n9664), .ZN(n9667) );
  AOI211_X1 U6515 ( .C1(n9735), .C2(n9734), .A(n9733), .B(n9732), .ZN(n9736)
         );
  NAND2_X1 U6516 ( .A1(n9641), .A2(n9640), .ZN(n9653) );
  NAND2_X1 U6517 ( .A1(n10109), .A2(n5435), .ZN(n5432) );
  NAND2_X1 U6518 ( .A1(n5432), .A2(n5433), .ZN(n8485) );
  NAND2_X1 U6519 ( .A1(n10109), .A2(n5439), .ZN(n5434) );
  NAND2_X1 U6520 ( .A1(n10109), .A2(n10112), .ZN(n10108) );
  NAND2_X1 U6521 ( .A1(n10203), .A2(n5441), .ZN(n5440) );
  NAND2_X1 U6522 ( .A1(n10162), .A2(n5446), .ZN(n5445) );
  NAND2_X1 U6523 ( .A1(n5450), .A2(n5454), .ZN(n7835) );
  NAND2_X1 U6524 ( .A1(n7794), .A2(n5451), .ZN(n5450) );
  NAND2_X2 U6525 ( .A1(n7287), .A2(n9402), .ZN(n5458) );
  AOI21_X1 U6526 ( .B1(n5458), .B2(n10837), .A(n10836), .ZN(n10839) );
  XNOR2_X1 U6527 ( .A(n5458), .B(n9564), .ZN(n9489) );
  XNOR2_X1 U6528 ( .A(n5458), .B(n9488), .ZN(n7289) );
  INV_X1 U6529 ( .A(n7837), .ZN(n5460) );
  NOR2_X1 U6530 ( .A1(n8478), .A2(n8477), .ZN(n10302) );
  NAND4_X1 U6531 ( .A1(n6473), .A2(n6525), .A3(n5472), .A4(n5470), .ZN(n6484)
         );
  NAND3_X1 U6532 ( .A1(n6473), .A2(n6525), .A3(n5472), .ZN(n6499) );
  AND2_X1 U6533 ( .A1(n5658), .A2(n5652), .ZN(n5472) );
  NOR2_X1 U6534 ( .A1(n9073), .A2(n6116), .ZN(n8867) );
  NAND3_X1 U6535 ( .A1(n10868), .A2(n8066), .A3(n5145), .ZN(n7384) );
  OAI211_X1 U6536 ( .C1(n5668), .C2(n5496), .A(n5494), .B(n5493), .ZN(n5497)
         );
  NAND3_X1 U6537 ( .A1(n5668), .A2(n5669), .A3(P2_DATAO_REG_2__SCAN_IN), .ZN(
        n5493) );
  INV_X1 U6538 ( .A(n5669), .ZN(n5495) );
  NAND2_X1 U6539 ( .A1(n5498), .A2(n5502), .ZN(n6345) );
  NAND2_X1 U6540 ( .A1(n7320), .A2(n5499), .ZN(n5498) );
  NAND3_X1 U6541 ( .A1(n5806), .A2(n5564), .A3(n5751), .ZN(n5842) );
  NAND2_X1 U6542 ( .A1(n6067), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6070) );
  AND2_X1 U6543 ( .A1(n6821), .A2(n6311), .ZN(n5530) );
  NAND2_X1 U6544 ( .A1(n5531), .A2(n5675), .ZN(n5811) );
  INV_X1 U6545 ( .A(n5672), .ZN(n5670) );
  AND2_X1 U6546 ( .A1(n8568), .A2(n8155), .ZN(n5540) );
  NAND2_X1 U6547 ( .A1(n5552), .A2(n5553), .ZN(n6118) );
  NAND2_X1 U6548 ( .A1(n6013), .A2(n6012), .ZN(n5563) );
  NOR2_X4 U6549 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5806) );
  XNOR2_X1 U6550 ( .A(n8235), .B(n6223), .ZN(n5568) );
  NAND2_X1 U6551 ( .A1(n8915), .A2(n5582), .ZN(n5581) );
  AND2_X1 U6552 ( .A1(n8153), .A2(n8144), .ZN(n5582) );
  NAND2_X1 U6553 ( .A1(n8875), .A2(n8153), .ZN(n8878) );
  OAI21_X1 U6554 ( .B1(n6240), .B2(n5588), .A(n5586), .ZN(n6242) );
  INV_X1 U6555 ( .A(n8120), .ZN(n5591) );
  NAND2_X1 U6556 ( .A1(n6238), .A2(n6237), .ZN(n7380) );
  AND2_X1 U6557 ( .A1(n6218), .A2(n5758), .ZN(n6221) );
  INV_X1 U6558 ( .A(n5611), .ZN(n9223) );
  NAND2_X1 U6559 ( .A1(n7690), .A2(n5624), .ZN(n5623) );
  NAND2_X1 U6560 ( .A1(n9172), .A2(n5084), .ZN(n5636) );
  NAND2_X1 U6561 ( .A1(n9296), .A2(n8424), .ZN(n9179) );
  INV_X1 U6562 ( .A(n9180), .ZN(n5649) );
  NAND2_X1 U6563 ( .A1(n6167), .A2(n6166), .ZN(n6172) );
  NAND2_X1 U6564 ( .A1(n6200), .A2(n6199), .ZN(n6204) );
  NAND2_X1 U6565 ( .A1(n6185), .A2(n6184), .ZN(n6189) );
  XNOR2_X1 U6566 ( .A(n6153), .B(n6152), .ZN(n9145) );
  NOR2_X2 U6567 ( .A1(n10226), .A2(n10368), .ZN(n10211) );
  XNOR2_X1 U6568 ( .A(n6118), .B(n6117), .ZN(n7957) );
  NAND2_X1 U6569 ( .A1(n8237), .A2(n8188), .ZN(n10808) );
  NOR2_X2 U6570 ( .A1(n10285), .A2(n10389), .ZN(n10269) );
  OR2_X1 U6571 ( .A1(n5034), .A2(n6876), .ZN(n6879) );
  OR2_X1 U6572 ( .A1(n5034), .A2(n10611), .ZN(n6869) );
  XNOR2_X1 U6573 ( .A(n6902), .B(n8418), .ZN(n6917) );
  NAND2_X2 U6574 ( .A1(n6634), .A2(n6881), .ZN(n5825) );
  OAI21_X2 U6575 ( .B1(n9284), .B2(n9285), .A(n9282), .ZN(n9172) );
  NOR2_X2 U6576 ( .A1(n6910), .A2(n10712), .ZN(n10714) );
  AND2_X1 U6577 ( .A1(n6677), .A2(n10864), .ZN(n10963) );
  INV_X1 U6578 ( .A(n10963), .ZN(n6439) );
  AND4_X1 U6579 ( .A1(n6044), .A2(n6043), .A3(n6042), .A4(n6041), .ZN(n8627)
         );
  OR2_X1 U6580 ( .A1(n9704), .A2(n9703), .ZN(n5655) );
  AND2_X1 U6581 ( .A1(n10439), .A2(n6478), .ZN(n5656) );
  AND2_X1 U6582 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_245), .ZN(n5657) );
  AND3_X1 U6583 ( .A1(n6491), .A2(n6493), .A3(n6495), .ZN(n5658) );
  AND3_X1 U6584 ( .A1(n5961), .A2(n5960), .A3(n5959), .ZN(n5660) );
  OR2_X1 U6585 ( .A1(n7017), .A2(n10721), .ZN(n5661) );
  AND2_X1 U6586 ( .A1(n8964), .A2(n8591), .ZN(n5662) );
  AND2_X1 U6587 ( .A1(n6210), .A2(n6194), .ZN(n8801) );
  INV_X1 U6588 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U6589 ( .A1(n7411), .A2(n7410), .ZN(n10830) );
  AND2_X1 U6590 ( .A1(n5867), .A2(n5689), .ZN(n5664) );
  INV_X1 U6591 ( .A(n8217), .ZN(n6215) );
  INV_X1 U6592 ( .A(n9100), .ZN(n6046) );
  AND2_X1 U6593 ( .A1(n8978), .A2(n8121), .ZN(n5665) );
  AND2_X1 U6594 ( .A1(n7294), .A2(n7293), .ZN(n5666) );
  NAND2_X1 U6595 ( .A1(n7145), .A2(n10937), .ZN(n10942) );
  AND3_X1 U6596 ( .A1(n7020), .A2(n7019), .A3(n7018), .ZN(n5667) );
  NAND2_X1 U6597 ( .A1(n9632), .A2(keyinput_132), .ZN(n9633) );
  NAND2_X1 U6598 ( .A1(n9634), .A2(n9633), .ZN(n9635) );
  INV_X1 U6599 ( .A(keyinput_133), .ZN(n9639) );
  INV_X1 U6600 ( .A(n9645), .ZN(n9648) );
  AND2_X1 U6601 ( .A1(n9648), .A2(n9647), .ZN(n9652) );
  XNOR2_X1 U6602 ( .A(n9702), .B(keyinput_175), .ZN(n9703) );
  AOI21_X1 U6603 ( .B1(n8059), .B2(n8058), .A(n10805), .ZN(n8065) );
  INV_X1 U6604 ( .A(n8208), .ZN(n8103) );
  NOR2_X1 U6605 ( .A1(n8104), .A2(n8103), .ZN(n8105) );
  NAND2_X1 U6606 ( .A1(n8122), .A2(n5665), .ZN(n8126) );
  NAND2_X1 U6607 ( .A1(n8159), .A2(n8186), .ZN(n8160) );
  NAND2_X1 U6608 ( .A1(n8156), .A2(n8155), .ZN(n8161) );
  NAND2_X1 U6609 ( .A1(n8163), .A2(n8833), .ZN(n8167) );
  INV_X1 U6610 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5759) );
  INV_X1 U6611 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6475) );
  OR2_X1 U6612 ( .A1(n6160), .A2(n9730), .ZN(n6175) );
  INV_X1 U6613 ( .A(n8207), .ZN(n6241) );
  NAND2_X1 U6614 ( .A1(n6901), .A2(n6900), .ZN(n6902) );
  INV_X1 U6615 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7714) );
  INV_X1 U6616 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7535) );
  INV_X1 U6617 ( .A(n9440), .ZN(n7836) );
  INV_X1 U6618 ( .A(n9488), .ZN(n7295) );
  INV_X1 U6619 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n7080) );
  NOR2_X1 U6620 ( .A1(n5704), .A2(n5914), .ZN(n5709) );
  OR2_X1 U6621 ( .A1(n6175), .A2(n9679), .ZN(n6193) );
  NAND2_X1 U6622 ( .A1(n6634), .A2(n8021), .ZN(n5830) );
  XNOR2_X1 U6623 ( .A(n6675), .B(n6303), .ZN(n6295) );
  INV_X1 U6624 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5902) );
  AND2_X1 U6625 ( .A1(n5936), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5952) );
  INV_X1 U6626 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9726) );
  AND2_X1 U6627 ( .A1(n8240), .A2(n6585), .ZN(n7154) );
  INV_X1 U6628 ( .A(n8421), .ZN(n8422) );
  NAND2_X1 U6629 ( .A1(n6895), .A2(n6881), .ZN(n7058) );
  AND2_X1 U6630 ( .A1(n8281), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8301) );
  AND2_X1 U6631 ( .A1(n6906), .A2(n5659), .ZN(n6907) );
  OR2_X1 U6632 ( .A1(n7763), .A2(n7762), .ZN(n7765) );
  NAND2_X1 U6633 ( .A1(n8313), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8326) );
  INV_X1 U6634 ( .A(n8354), .ZN(n8368) );
  OR2_X1 U6635 ( .A1(n8326), .A2(n8325), .ZN(n8340) );
  NAND2_X1 U6636 ( .A1(n8000), .A2(n7999), .ZN(n8002) );
  INV_X1 U6637 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U6638 ( .A1(n6118), .A2(n6117), .ZN(n6123) );
  INV_X1 U6639 ( .A(SI_13_), .ZN(n5719) );
  INV_X1 U6640 ( .A(n8538), .ZN(n6310) );
  INV_X1 U6641 ( .A(n10968), .ZN(n6450) );
  OR2_X1 U6642 ( .A1(n6431), .A2(n6430), .ZN(n6445) );
  NAND2_X1 U6643 ( .A1(n6084), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6085) );
  INV_X1 U6644 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8682) );
  INV_X1 U6645 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9700) );
  NAND2_X1 U6646 ( .A1(n8820), .A2(n8813), .ZN(n8826) );
  AOI21_X1 U6647 ( .B1(n7944), .B2(n7945), .A(n6011), .ZN(n9007) );
  INV_X1 U6648 ( .A(n10864), .ZN(n11028) );
  OR2_X1 U6649 ( .A1(n6431), .A2(n7154), .ZN(n6289) );
  NAND2_X1 U6650 ( .A1(n8423), .A2(n8422), .ZN(n8424) );
  NOR2_X1 U6651 ( .A1(n8385), .A2(n8384), .ZN(n9164) );
  NAND2_X1 U6652 ( .A1(n7982), .A2(n6565), .ZN(n6898) );
  INV_X1 U6653 ( .A(n6871), .ZN(n9591) );
  INV_X1 U6654 ( .A(n6932), .ZN(n6936) );
  NOR2_X1 U6655 ( .A1(n8340), .A2(n9254), .ZN(n8353) );
  INV_X1 U6656 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7721) );
  INV_X1 U6657 ( .A(n10353), .ZN(n10160) );
  NAND2_X1 U6658 ( .A1(n8486), .A2(n10920), .ZN(n8493) );
  AND2_X1 U6659 ( .A1(n7144), .A2(n7492), .ZN(n10711) );
  OR2_X1 U6660 ( .A1(n10512), .A2(n6871), .ZN(n10915) );
  OR3_X1 U6661 ( .A1(n10458), .A2(n6839), .A3(n8012), .ZN(n6530) );
  XNOR2_X1 U6662 ( .A(n5712), .B(n9662), .ZN(n5928) );
  AND2_X1 U6663 ( .A1(n10955), .A2(n9016), .ZN(n10884) );
  AND2_X1 U6664 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5851) );
  AND3_X1 U6665 ( .A1(n8033), .A2(n8032), .A3(n8031), .ZN(n8652) );
  AND4_X1 U6666 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .ZN(n8568)
         );
  AND4_X1 U6667 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n8590)
         );
  OR2_X1 U6668 ( .A1(n8670), .A2(n8669), .ZN(n8672) );
  AND2_X1 U6669 ( .A1(n6998), .A2(n6997), .ZN(n6999) );
  INV_X1 U6670 ( .A(n10624), .ZN(n10656) );
  INV_X1 U6671 ( .A(n10648), .ZN(n10622) );
  INV_X1 U6672 ( .A(n8805), .ZN(n8798) );
  INV_X1 U6673 ( .A(n8852), .ZN(n8845) );
  INV_X1 U6674 ( .A(n10794), .ZN(n9016) );
  INV_X1 U6675 ( .A(n8963), .ZN(n10767) );
  AND2_X1 U6676 ( .A1(n6290), .A2(n10617), .ZN(n6456) );
  INV_X1 U6677 ( .A(n11034), .ZN(n11008) );
  NAND2_X1 U6678 ( .A1(n8985), .A2(n10743), .ZN(n11034) );
  NAND2_X1 U6679 ( .A1(n10468), .A2(n6282), .ZN(n10470) );
  AND2_X1 U6680 ( .A1(n5877), .A2(n5885), .ZN(n6740) );
  AND2_X1 U6681 ( .A1(n10458), .A2(n6839), .ZN(n6490) );
  INV_X1 U6682 ( .A(n10110), .ZN(n10144) );
  AND4_X1 U6683 ( .A1(n8264), .A2(n8263), .A3(n8262), .A4(n8261), .ZN(n10250)
         );
  AND2_X1 U6684 ( .A1(n6957), .A2(n6956), .ZN(n10572) );
  OR2_X1 U6685 ( .A1(n10559), .A2(n6574), .ZN(n10691) );
  OR2_X1 U6686 ( .A1(n10559), .A2(n10512), .ZN(n10665) );
  INV_X1 U6687 ( .A(n10700), .ZN(n10664) );
  INV_X1 U6688 ( .A(n8483), .ZN(n10134) );
  AND2_X1 U6689 ( .A1(n9510), .A2(n9511), .ZN(n9429) );
  INV_X1 U6690 ( .A(n10736), .ZN(n9341) );
  INV_X1 U6691 ( .A(n6934), .ZN(n6935) );
  AND2_X1 U6692 ( .A1(n6842), .A2(n6841), .ZN(n7479) );
  OR2_X1 U6693 ( .A1(n9559), .A2(n9598), .ZN(n10707) );
  AND3_X1 U6694 ( .A1(n6858), .A2(n6934), .A3(n6857), .ZN(n7481) );
  NOR2_X1 U6695 ( .A1(n7022), .A2(P1_U3084), .ZN(n7480) );
  AND2_X1 U6696 ( .A1(n6629), .A2(n6703), .ZN(n7750) );
  NOR2_X1 U6697 ( .A1(n10485), .A2(n7635), .ZN(n7636) );
  NOR2_X1 U6698 ( .A1(n10496), .A2(n10495), .ZN(n7652) );
  NAND2_X1 U6699 ( .A1(n6587), .A2(n6586), .ZN(n10647) );
  INV_X1 U6700 ( .A(n7908), .ZN(n11029) );
  NAND2_X1 U6701 ( .A1(n6449), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10968) );
  AND4_X1 U6702 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6211), .ZN(n6977)
         );
  NAND2_X1 U6703 ( .A1(n6652), .A2(n6253), .ZN(n10638) );
  AND2_X1 U6704 ( .A1(n8975), .A2(n8977), .ZN(n9103) );
  INV_X1 U6705 ( .A(n11037), .ZN(n11036) );
  AND2_X2 U6706 ( .A1(n6457), .A2(n6456), .ZN(n11037) );
  INV_X1 U6707 ( .A(n11041), .ZN(n11038) );
  NAND2_X1 U6708 ( .A1(n10471), .A2(n10470), .ZN(n10618) );
  AND2_X1 U6709 ( .A1(n6582), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10621) );
  XNOR2_X1 U6710 ( .A(n6279), .B(n6278), .ZN(n7890) );
  INV_X1 U6711 ( .A(n9134), .ZN(n9146) );
  INV_X1 U6712 ( .A(n9188), .ZN(n10102) );
  INV_X1 U6713 ( .A(n8457), .ZN(n10180) );
  INV_X1 U6714 ( .A(n10250), .ZN(n10294) );
  OR2_X1 U6715 ( .A1(P1_U3083), .A2(n6578), .ZN(n10700) );
  NAND2_X1 U6716 ( .A1(n10942), .A2(n10725), .ZN(n10935) );
  NAND2_X1 U6717 ( .A1(n9600), .A2(n6935), .ZN(n10937) );
  INV_X1 U6718 ( .A(n11050), .ZN(n11049) );
  AND2_X1 U6719 ( .A1(n10880), .A2(n10879), .ZN(n10882) );
  INV_X1 U6720 ( .A(n11054), .ZN(n11051) );
  AND3_X2 U6721 ( .A1(n7110), .A2(n7480), .A3(n7481), .ZN(n11054) );
  AND2_X1 U6722 ( .A1(n7799), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6534) );
  NOR2_X1 U6723 ( .A1(n7653), .A2(n7652), .ZN(n10498) );
  AND2_X1 U6724 ( .A1(n6911), .A2(n6534), .ZN(P1_U4006) );
  INV_X1 U6725 ( .A(SI_0_), .ZN(n6859) );
  INV_X1 U6726 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6860) );
  INV_X1 U6727 ( .A(SI_1_), .ZN(n5671) );
  NAND2_X1 U6728 ( .A1(n5672), .A2(n5671), .ZN(n5673) );
  AND2_X1 U6729 ( .A1(n5674), .A2(n5673), .ZN(n5781) );
  MUX2_X1 U6730 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6507), .Z(n5782) );
  INV_X1 U6731 ( .A(n5809), .ZN(n5675) );
  NAND2_X1 U6732 ( .A1(n5811), .A2(n5676), .ZN(n5827) );
  MUX2_X1 U6733 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6507), .Z(n5677) );
  NAND2_X1 U6734 ( .A1(n5677), .A2(SI_3_), .ZN(n5681) );
  INV_X1 U6735 ( .A(n5677), .ZN(n5679) );
  INV_X1 U6736 ( .A(SI_3_), .ZN(n5678) );
  NAND2_X1 U6737 ( .A1(n5679), .A2(n5678), .ZN(n5680) );
  AND2_X1 U6738 ( .A1(n5681), .A2(n5680), .ZN(n5826) );
  NAND2_X1 U6739 ( .A1(n5827), .A2(n5826), .ZN(n5829) );
  NAND2_X1 U6740 ( .A1(n5829), .A2(n5681), .ZN(n5845) );
  MUX2_X1 U6741 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6881), .Z(n5682) );
  NAND2_X1 U6742 ( .A1(n5682), .A2(SI_4_), .ZN(n5685) );
  INV_X1 U6743 ( .A(n5682), .ZN(n5684) );
  INV_X1 U6744 ( .A(SI_4_), .ZN(n5683) );
  NAND2_X1 U6745 ( .A1(n5845), .A2(n5844), .ZN(n5847) );
  MUX2_X1 U6746 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6881), .Z(n5686) );
  NAND2_X1 U6747 ( .A1(n5686), .A2(SI_5_), .ZN(n5867) );
  INV_X1 U6748 ( .A(n5686), .ZN(n5688) );
  INV_X1 U6749 ( .A(SI_5_), .ZN(n5687) );
  NAND2_X1 U6750 ( .A1(n5688), .A2(n5687), .ZN(n5689) );
  MUX2_X1 U6751 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6881), .Z(n5690) );
  NAND2_X1 U6752 ( .A1(n5690), .A2(SI_6_), .ZN(n5695) );
  INV_X1 U6753 ( .A(n5690), .ZN(n5691) );
  INV_X1 U6754 ( .A(SI_6_), .ZN(n9671) );
  NAND2_X1 U6755 ( .A1(n5691), .A2(n9671), .ZN(n5692) );
  NAND2_X1 U6756 ( .A1(n5695), .A2(n5692), .ZN(n5694) );
  INV_X1 U6757 ( .A(n5694), .ZN(n5872) );
  NAND2_X1 U6758 ( .A1(n5857), .A2(n5693), .ZN(n5870) );
  MUX2_X1 U6759 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6881), .Z(n5697) );
  NAND2_X1 U6760 ( .A1(n5697), .A2(SI_7_), .ZN(n5701) );
  INV_X1 U6761 ( .A(n5697), .ZN(n5699) );
  INV_X1 U6762 ( .A(SI_7_), .ZN(n5698) );
  NAND2_X1 U6763 ( .A1(n5699), .A2(n5698), .ZN(n5700) );
  MUX2_X1 U6764 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6881), .Z(n5705) );
  XNOR2_X1 U6765 ( .A(n5705), .B(SI_8_), .ZN(n5910) );
  MUX2_X1 U6766 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n6881), .Z(n5703) );
  INV_X1 U6767 ( .A(n5703), .ZN(n5702) );
  NAND2_X1 U6768 ( .A1(n5702), .A2(n9668), .ZN(n5707) );
  INV_X1 U6769 ( .A(n5707), .ZN(n5704) );
  XNOR2_X1 U6770 ( .A(n5703), .B(n9668), .ZN(n5914) );
  INV_X1 U6771 ( .A(n5705), .ZN(n5706) );
  INV_X1 U6772 ( .A(SI_8_), .ZN(n9672) );
  NAND2_X1 U6773 ( .A1(n5706), .A2(n9672), .ZN(n5912) );
  AND2_X1 U6774 ( .A1(n5912), .A2(n5707), .ZN(n5708) );
  MUX2_X1 U6775 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6881), .Z(n5712) );
  INV_X1 U6776 ( .A(n5712), .ZN(n5713) );
  NAND2_X1 U6777 ( .A1(n5713), .A2(n9662), .ZN(n5714) );
  MUX2_X1 U6778 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6881), .Z(n5715) );
  OAI21_X1 U6779 ( .B1(n5715), .B2(SI_11_), .A(n5716), .ZN(n5944) );
  MUX2_X1 U6780 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6507), .Z(n5717) );
  MUX2_X1 U6781 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6881), .Z(n5718) );
  XNOR2_X1 U6782 ( .A(n5718), .B(n5719), .ZN(n5973) );
  INV_X1 U6783 ( .A(n5718), .ZN(n5720) );
  NAND2_X1 U6784 ( .A1(n5720), .A2(n5719), .ZN(n5721) );
  MUX2_X1 U6785 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6881), .Z(n5723) );
  INV_X1 U6786 ( .A(n5723), .ZN(n5725) );
  INV_X1 U6787 ( .A(SI_14_), .ZN(n5724) );
  NAND2_X1 U6788 ( .A1(n5725), .A2(n5724), .ZN(n5726) );
  MUX2_X1 U6789 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6881), .Z(n5728) );
  XNOR2_X1 U6790 ( .A(n5728), .B(SI_15_), .ZN(n5998) );
  INV_X1 U6791 ( .A(n5728), .ZN(n5730) );
  INV_X1 U6792 ( .A(SI_15_), .ZN(n5729) );
  MUX2_X1 U6793 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6881), .Z(n5731) );
  XNOR2_X1 U6794 ( .A(n5731), .B(n9625), .ZN(n6012) );
  INV_X1 U6795 ( .A(n5731), .ZN(n5732) );
  NAND2_X1 U6796 ( .A1(n5732), .A2(n9625), .ZN(n5733) );
  MUX2_X1 U6797 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6881), .Z(n5734) );
  OAI21_X1 U6798 ( .B1(n5734), .B2(SI_17_), .A(n5735), .ZN(n6032) );
  MUX2_X1 U6799 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6881), .Z(n5736) );
  INV_X1 U6800 ( .A(n5736), .ZN(n5737) );
  INV_X1 U6801 ( .A(SI_18_), .ZN(n9657) );
  NAND2_X1 U6802 ( .A1(n5737), .A2(n9657), .ZN(n5738) );
  MUX2_X1 U6803 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n6881), .Z(n5740) );
  XNOR2_X1 U6804 ( .A(n5740), .B(SI_19_), .ZN(n6063) );
  INV_X1 U6805 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U6806 ( .A1(n5741), .A2(n9627), .ZN(n5742) );
  MUX2_X1 U6807 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6881), .Z(n5743) );
  INV_X1 U6808 ( .A(n5743), .ZN(n5745) );
  MUX2_X1 U6809 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6881), .Z(n5746) );
  NAND2_X1 U6810 ( .A1(n5746), .A2(SI_21_), .ZN(n6090) );
  OAI21_X1 U6811 ( .B1(n5746), .B2(SI_21_), .A(n6090), .ZN(n5748) );
  NAND2_X1 U6812 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U6813 ( .A1(n6091), .A2(n5750), .ZN(n7989) );
  NOR2_X1 U6814 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5756) );
  NOR2_X1 U6815 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5755) );
  NOR2_X1 U6816 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5754) );
  NOR2_X1 U6817 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5753) );
  OR2_X1 U6818 ( .A1(n7989), .A2(n6128), .ZN(n5765) );
  INV_X1 U6819 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7501) );
  OR2_X1 U6820 ( .A1(n5825), .A2(n7501), .ZN(n5764) );
  INV_X1 U6821 ( .A(n9079), .ZN(n8914) );
  NAND2_X1 U6822 ( .A1(n5767), .A2(n5761), .ZN(n5769) );
  INV_X1 U6823 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U6824 ( .A1(n8030), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U6825 ( .A1(n8029), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5777) );
  INV_X1 U6826 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9701) );
  NAND2_X1 U6827 ( .A1(n5851), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U6828 ( .A1(n5889), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5903) );
  INV_X1 U6829 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5977) );
  INV_X1 U6830 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U6831 ( .A1(n6005), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6025) );
  INV_X1 U6832 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8579) );
  INV_X1 U6833 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U6834 ( .A1(n9701), .A2(n6085), .ZN(n5774) );
  INV_X1 U6835 ( .A(n6085), .ZN(n5773) );
  NAND2_X1 U6836 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(n5773), .ZN(n6095) );
  AND2_X1 U6837 ( .A1(n5774), .A2(n6095), .ZN(n8912) );
  NAND2_X1 U6838 ( .A1(n5919), .A2(n8912), .ZN(n5776) );
  AND2_X2 U6839 ( .A1(n8499), .A2(n9138), .ZN(n5801) );
  INV_X1 U6840 ( .A(n5801), .ZN(n5862) );
  NAND2_X1 U6841 ( .A1(n6131), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5775) );
  INV_X1 U6842 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U6843 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5779) );
  XNOR2_X1 U6844 ( .A(n5780), .B(n5779), .ZN(n10637) );
  INV_X1 U6845 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6503) );
  OR2_X1 U6846 ( .A1(n5825), .A2(n6503), .ZN(n5788) );
  INV_X1 U6847 ( .A(n5781), .ZN(n5784) );
  INV_X1 U6848 ( .A(n5782), .ZN(n5783) );
  NAND2_X1 U6849 ( .A1(n5784), .A2(n5783), .ZN(n5785) );
  NAND2_X1 U6850 ( .A1(n5786), .A2(n5785), .ZN(n6896) );
  OR2_X1 U6851 ( .A1(n5830), .A2(n6896), .ZN(n5787) );
  NAND2_X1 U6852 ( .A1(n5793), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U6853 ( .A1(n5801), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U6854 ( .A1(n5801), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U6855 ( .A1(n5901), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U6856 ( .A1(n5800), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U6857 ( .A1(n8021), .A2(SI_0_), .ZN(n5798) );
  XNOR2_X1 U6858 ( .A(n5798), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9150) );
  MUX2_X1 U6859 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9150), .S(n6634), .Z(n6690) );
  NAND2_X1 U6860 ( .A1(n7469), .A2(n6692), .ZN(n5799) );
  NAND2_X1 U6861 ( .A1(n5793), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U6862 ( .A1(n5901), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U6863 ( .A1(n5800), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U6864 ( .A1(n5801), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5802) );
  NAND4_X1 U6865 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n5815)
         );
  OR2_X1 U6866 ( .A1(n5806), .A2(n9131), .ZN(n5808) );
  INV_X1 U6867 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U6868 ( .A1(n5808), .A2(n5807), .ZN(n5822) );
  OAI21_X1 U6869 ( .B1(n5808), .B2(n5807), .A(n5822), .ZN(n6646) );
  OR2_X1 U6870 ( .A1(n5825), .A2(n5496), .ZN(n5814) );
  NAND2_X1 U6871 ( .A1(n5810), .A2(n5809), .ZN(n5812) );
  NAND2_X1 U6872 ( .A1(n5812), .A2(n5811), .ZN(n6882) );
  OR2_X1 U6873 ( .A1(n5830), .A2(n6882), .ZN(n5813) );
  OAI211_X1 U6874 ( .C1(n6634), .C2(n6646), .A(n5814), .B(n5813), .ZN(n7463)
         );
  NAND2_X1 U6875 ( .A1(n5815), .A2(n5269), .ZN(n8043) );
  CLKBUF_X1 U6876 ( .A(n5269), .Z(n10744) );
  NAND2_X1 U6877 ( .A1(n5816), .A2(n10744), .ZN(n5817) );
  NAND2_X1 U6878 ( .A1(n7461), .A2(n5817), .ZN(n7041) );
  NAND2_X1 U6879 ( .A1(n5793), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U6880 ( .A1(n5800), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5820) );
  INV_X1 U6881 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10763) );
  NAND2_X1 U6882 ( .A1(n5901), .A2(n10763), .ZN(n5819) );
  NAND2_X1 U6883 ( .A1(n5801), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U6884 ( .A1(n5822), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5824) );
  INV_X1 U6885 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5823) );
  XNOR2_X1 U6886 ( .A(n5824), .B(n5823), .ZN(n6776) );
  INV_X1 U6887 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6504) );
  OR2_X1 U6888 ( .A1(n5825), .A2(n6504), .ZN(n5832) );
  OR2_X1 U6889 ( .A1(n5827), .A2(n5826), .ZN(n5828) );
  OR2_X1 U6890 ( .A1(n5830), .A2(n7003), .ZN(n5831) );
  NAND2_X1 U6891 ( .A1(n6592), .A2(n6304), .ZN(n8052) );
  NAND2_X1 U6892 ( .A1(n6825), .A2(n10766), .ZN(n8051) );
  NAND2_X1 U6893 ( .A1(n7041), .A2(n8054), .ZN(n7040) );
  NAND2_X1 U6894 ( .A1(n6825), .A2(n6304), .ZN(n5833) );
  NAND2_X1 U6895 ( .A1(n7040), .A2(n5833), .ZN(n7251) );
  INV_X1 U6896 ( .A(n5851), .ZN(n5835) );
  INV_X1 U6897 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9710) );
  NAND2_X1 U6898 ( .A1(n9710), .A2(n10763), .ZN(n5834) );
  NAND2_X1 U6899 ( .A1(n5835), .A2(n5834), .ZN(n7259) );
  INV_X1 U6900 ( .A(n7259), .ZN(n6827) );
  NAND2_X1 U6901 ( .A1(n5919), .A2(n6827), .ZN(n5839) );
  NAND2_X1 U6902 ( .A1(n5793), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U6903 ( .A1(n6131), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U6904 ( .A1(n8030), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U6905 ( .A1(n5840), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5841) );
  MUX2_X1 U6906 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5841), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5843) );
  NAND2_X1 U6907 ( .A1(n5843), .A2(n5842), .ZN(n6665) );
  OR2_X1 U6908 ( .A1(n5845), .A2(n5844), .ZN(n5846) );
  INV_X1 U6909 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6513) );
  OR2_X1 U6910 ( .A1(n5825), .A2(n6513), .ZN(n5848) );
  OAI211_X1 U6911 ( .C1(n6634), .C2(n6665), .A(n5849), .B(n5848), .ZN(n7263)
         );
  NAND2_X1 U6912 ( .A1(n10793), .A2(n7263), .ZN(n8056) );
  NAND2_X1 U6913 ( .A1(n8056), .A2(n8057), .ZN(n7253) );
  NAND2_X1 U6914 ( .A1(n10793), .A2(n10784), .ZN(n5850) );
  NAND2_X1 U6915 ( .A1(n8030), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U6916 ( .A1(n5793), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5854) );
  OAI21_X1 U6917 ( .B1(n5851), .B2(P2_REG3_REG_5__SCAN_IN), .A(n5860), .ZN(
        n10801) );
  INV_X1 U6918 ( .A(n10801), .ZN(n10812) );
  NAND2_X1 U6919 ( .A1(n5919), .A2(n10812), .ZN(n5853) );
  NAND2_X1 U6920 ( .A1(n6131), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U6921 ( .A1(n5842), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5856) );
  XNOR2_X1 U6922 ( .A(n5856), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6741) );
  INV_X1 U6923 ( .A(n6741), .ZN(n6670) );
  NAND2_X1 U6924 ( .A1(n5857), .A2(n5664), .ZN(n5868) );
  OR2_X1 U6925 ( .A1(n5857), .A2(n5664), .ZN(n5858) );
  INV_X1 U6926 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6515) );
  OR2_X1 U6927 ( .A1(n5825), .A2(n6515), .ZN(n5859) );
  NAND2_X1 U6928 ( .A1(n7091), .A2(n10810), .ZN(n8060) );
  INV_X1 U6929 ( .A(n7091), .ZN(n9015) );
  NAND2_X1 U6930 ( .A1(n9015), .A2(n10824), .ZN(n6235) );
  NAND2_X1 U6931 ( .A1(n8060), .A2(n6235), .ZN(n10805) );
  NAND2_X1 U6932 ( .A1(n7091), .A2(n10824), .ZN(n9020) );
  NAND2_X1 U6933 ( .A1(n8030), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5866) );
  NAND2_X1 U6934 ( .A1(n5793), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5865) );
  AND2_X1 U6935 ( .A1(n5860), .A2(n9726), .ZN(n5861) );
  NOR2_X1 U6936 ( .A1(n5889), .A2(n5861), .ZN(n9019) );
  NAND2_X1 U6937 ( .A1(n5919), .A2(n9019), .ZN(n5864) );
  NAND2_X1 U6938 ( .A1(n6131), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5863) );
  NAND4_X1 U6939 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n8664)
         );
  OR2_X1 U6940 ( .A1(n5873), .A2(n9131), .ZN(n5876) );
  INV_X1 U6941 ( .A(n5876), .ZN(n5874) );
  NAND2_X1 U6942 ( .A1(n5874), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5877) );
  INV_X1 U6943 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U6944 ( .A1(n5876), .A2(n5875), .ZN(n5885) );
  AOI22_X1 U6945 ( .A1(n6072), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6583), .B2(
        n6740), .ZN(n5878) );
  INV_X1 U6946 ( .A(n9022), .ZN(n8200) );
  NAND2_X1 U6947 ( .A1(n10863), .A2(n8664), .ZN(n8066) );
  NAND2_X1 U6948 ( .A1(n5885), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5886) );
  XNOR2_X1 U6949 ( .A(n5886), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6785) );
  AOI22_X1 U6950 ( .A1(n6072), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6583), .B2(
        n6785), .ZN(n5887) );
  NAND2_X1 U6951 ( .A1(n8030), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U6952 ( .A1(n5793), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5893) );
  OR2_X1 U6953 ( .A1(n5889), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U6954 ( .A1(n5903), .A2(n5890), .ZN(n10897) );
  INV_X1 U6955 ( .A(n10897), .ZN(n7387) );
  NAND2_X1 U6956 ( .A1(n5919), .A2(n7387), .ZN(n5892) );
  NAND2_X1 U6957 ( .A1(n6131), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U6958 ( .A1(n10895), .A2(n6323), .ZN(n8070) );
  INV_X1 U6959 ( .A(n6323), .ZN(n9017) );
  OR2_X1 U6960 ( .A1(n10895), .A2(n9017), .ZN(n5896) );
  NAND2_X1 U6961 ( .A1(n7522), .A2(n8036), .ZN(n5900) );
  XNOR2_X1 U6962 ( .A(n5898), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6788) );
  AOI22_X1 U6963 ( .A1(n6072), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6583), .B2(
        n6788), .ZN(n5899) );
  NAND2_X1 U6964 ( .A1(n8030), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U6965 ( .A1(n8029), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U6966 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  AND2_X1 U6967 ( .A1(n5920), .A2(n5904), .ZN(n7368) );
  NAND2_X1 U6968 ( .A1(n5919), .A2(n7368), .ZN(n5906) );
  NAND2_X1 U6969 ( .A1(n6131), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5905) );
  INV_X1 U6970 ( .A(n8076), .ZN(n10883) );
  NAND2_X1 U6971 ( .A1(n8077), .A2(n10883), .ZN(n5909) );
  NAND2_X1 U6972 ( .A1(n5913), .A2(n5912), .ZN(n5915) );
  XNOR2_X1 U6973 ( .A(n5915), .B(n5914), .ZN(n7532) );
  NAND2_X1 U6974 ( .A1(n7532), .A2(n8036), .ZN(n5918) );
  INV_X1 U6975 ( .A(n5962), .ZN(n5916) );
  NAND2_X1 U6976 ( .A1(n5916), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5930) );
  XNOR2_X1 U6977 ( .A(n5930), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8687) );
  AOI22_X1 U6978 ( .A1(n6072), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6583), .B2(
        n8687), .ZN(n5917) );
  NAND2_X1 U6979 ( .A1(n8030), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U6980 ( .A1(n8029), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5925) );
  AND2_X1 U6981 ( .A1(n5920), .A2(n8682), .ZN(n5921) );
  OR2_X1 U6982 ( .A1(n5921), .A2(n5936), .ZN(n10969) );
  INV_X1 U6983 ( .A(n10969), .ZN(n5922) );
  NAND2_X1 U6984 ( .A1(n5919), .A2(n5922), .ZN(n5924) );
  NAND2_X1 U6985 ( .A1(n6131), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U6986 ( .A1(n10962), .A2(n7507), .ZN(n8084) );
  NAND2_X1 U6987 ( .A1(n8086), .A2(n8084), .ZN(n7400) );
  INV_X1 U6988 ( .A(n7507), .ZN(n7323) );
  OR2_X1 U6989 ( .A1(n10962), .A2(n7323), .ZN(n5927) );
  NAND2_X1 U6990 ( .A1(n7700), .A2(n8036), .ZN(n5935) );
  NAND2_X1 U6991 ( .A1(n5930), .A2(n5961), .ZN(n5931) );
  NAND2_X1 U6992 ( .A1(n5931), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U6993 ( .A1(n5932), .A2(n5960), .ZN(n5948) );
  OR2_X1 U6994 ( .A1(n5932), .A2(n5960), .ZN(n5933) );
  AOI22_X1 U6995 ( .A1(n6072), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6583), .B2(
        n6807), .ZN(n5934) );
  NAND2_X1 U6996 ( .A1(n5935), .A2(n5934), .ZN(n7516) );
  NAND2_X1 U6997 ( .A1(n8029), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U6998 ( .A1(n6131), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5940) );
  NOR2_X1 U6999 ( .A1(n5936), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5937) );
  OR2_X1 U7000 ( .A1(n5952), .A2(n5937), .ZN(n7511) );
  INV_X1 U7001 ( .A(n7511), .ZN(n7497) );
  NAND2_X1 U7002 ( .A1(n5919), .A2(n7497), .ZN(n5939) );
  NAND2_X1 U7003 ( .A1(n8030), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5938) );
  OR2_X1 U7004 ( .A1(n7516), .A2(n7562), .ZN(n8089) );
  NAND2_X1 U7005 ( .A1(n7516), .A2(n7562), .ZN(n8088) );
  INV_X1 U7006 ( .A(n7562), .ZN(n8663) );
  NAND2_X1 U7007 ( .A1(n7516), .A2(n8663), .ZN(n5943) );
  NAND2_X1 U7008 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  NAND2_X1 U7009 ( .A1(n5947), .A2(n5946), .ZN(n7744) );
  OR2_X1 U7010 ( .A1(n7744), .A2(n6128), .ZN(n5951) );
  NAND2_X1 U7011 ( .A1(n5948), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5949) );
  XNOR2_X1 U7012 ( .A(n5949), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6996) );
  AOI22_X1 U7013 ( .A1(n6072), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6583), .B2(
        n6996), .ZN(n5950) );
  NAND2_X1 U7014 ( .A1(n5951), .A2(n5950), .ZN(n7621) );
  NAND2_X1 U7015 ( .A1(n8030), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7016 ( .A1(n8029), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5956) );
  OR2_X1 U7017 ( .A1(n5952), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5953) );
  AND2_X1 U7018 ( .A1(n5966), .A2(n5953), .ZN(n7617) );
  NAND2_X1 U7019 ( .A1(n5919), .A2(n7617), .ZN(n5955) );
  NAND2_X1 U7020 ( .A1(n6131), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5954) );
  OR2_X1 U7021 ( .A1(n7621), .A2(n7685), .ZN(n8096) );
  NAND2_X1 U7022 ( .A1(n7621), .A2(n7685), .ZN(n8094) );
  NAND2_X1 U7023 ( .A1(n8096), .A2(n8094), .ZN(n7613) );
  INV_X1 U7024 ( .A(n7685), .ZN(n8662) );
  NAND2_X1 U7025 ( .A1(n7621), .A2(n8662), .ZN(n5958) );
  NAND2_X1 U7026 ( .A1(n7749), .A2(n8036), .ZN(n5965) );
  NAND2_X1 U7027 ( .A1(n5962), .A2(n5660), .ZN(n5974) );
  NAND2_X1 U7028 ( .A1(n5974), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U7029 ( .A(n5963), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7179) );
  AOI22_X1 U7030 ( .A1(n6072), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6583), .B2(
        n7179), .ZN(n5964) );
  NAND2_X1 U7031 ( .A1(n8029), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7032 ( .A1(n6131), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7033 ( .A1(n5966), .A2(n9700), .ZN(n5967) );
  AND2_X1 U7034 ( .A1(n5978), .A2(n5967), .ZN(n7736) );
  NAND2_X1 U7035 ( .A1(n5919), .A2(n7736), .ZN(n5969) );
  NAND2_X1 U7036 ( .A1(n8030), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7037 ( .A1(n7737), .A2(n7915), .ZN(n8098) );
  INV_X1 U7038 ( .A(n7915), .ZN(n8661) );
  OR2_X1 U7039 ( .A1(n7737), .A2(n8661), .ZN(n5972) );
  XNOR2_X1 U7040 ( .A(n5081), .B(n5973), .ZN(n7819) );
  NAND2_X1 U7041 ( .A1(n7819), .A2(n8036), .ZN(n5976) );
  OR2_X1 U7042 ( .A1(n6018), .A2(n9131), .ZN(n5987) );
  XNOR2_X1 U7043 ( .A(n5987), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7314) );
  AOI22_X1 U7044 ( .A1(n6072), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6583), .B2(
        n7314), .ZN(n5975) );
  NAND2_X1 U7045 ( .A1(n8030), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5983) );
  NAND2_X1 U7046 ( .A1(n8029), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7047 ( .A1(n5978), .A2(n5977), .ZN(n5979) );
  AND2_X1 U7048 ( .A1(n5992), .A2(n5979), .ZN(n7919) );
  NAND2_X1 U7049 ( .A1(n5919), .A2(n7919), .ZN(n5981) );
  NAND2_X1 U7050 ( .A1(n6131), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5980) );
  NAND4_X1 U7051 ( .A1(n5983), .A2(n5982), .A3(n5981), .A4(n5980), .ZN(n8660)
         );
  XNOR2_X1 U7052 ( .A(n8107), .B(n8660), .ZN(n8208) );
  NAND2_X1 U7053 ( .A1(n8107), .A2(n8660), .ZN(n5985) );
  XNOR2_X1 U7054 ( .A(n5986), .B(n5092), .ZN(n7965) );
  NAND2_X1 U7055 ( .A1(n7965), .A2(n8036), .ZN(n5990) );
  NAND2_X1 U7056 ( .A1(n5987), .A2(n6016), .ZN(n5988) );
  NAND2_X1 U7057 ( .A1(n5988), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6000) );
  XNOR2_X1 U7058 ( .A(n6000), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8693) );
  AOI22_X1 U7059 ( .A1(n6072), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6583), .B2(
        n8693), .ZN(n5989) );
  NAND2_X1 U7060 ( .A1(n8030), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7061 ( .A1(n8029), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5996) );
  AND2_X1 U7062 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  NOR2_X1 U7063 ( .A1(n6005), .A2(n5993), .ZN(n7936) );
  NAND2_X1 U7064 ( .A1(n5919), .A2(n7936), .ZN(n5995) );
  NAND2_X1 U7065 ( .A1(n6131), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7066 ( .A1(n7908), .A2(n8646), .ZN(n8113) );
  NAND2_X1 U7067 ( .A1(n8112), .A2(n8113), .ZN(n8207) );
  INV_X1 U7068 ( .A(n8646), .ZN(n8659) );
  XNOR2_X1 U7069 ( .A(n5999), .B(n5998), .ZN(n7968) );
  NAND2_X1 U7070 ( .A1(n7968), .A2(n8036), .ZN(n6004) );
  NAND2_X1 U7071 ( .A1(n6000), .A2(n6015), .ZN(n6001) );
  NAND2_X1 U7072 ( .A1(n6001), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6002) );
  XNOR2_X1 U7073 ( .A(n6002), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8714) );
  AOI22_X1 U7074 ( .A1(n6072), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6583), .B2(
        n8714), .ZN(n6003) );
  NAND2_X1 U7075 ( .A1(n8030), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7076 ( .A1(n8029), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6009) );
  OR2_X1 U7077 ( .A1(n6005), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6006) );
  AND2_X1 U7078 ( .A1(n6006), .A2(n6025), .ZN(n8648) );
  NAND2_X1 U7079 ( .A1(n5919), .A2(n8648), .ZN(n6008) );
  NAND2_X1 U7080 ( .A1(n6131), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6007) );
  OR2_X1 U7081 ( .A1(n9109), .A2(n8578), .ZN(n8116) );
  NAND2_X1 U7082 ( .A1(n9109), .A2(n8578), .ZN(n8994) );
  NAND2_X1 U7083 ( .A1(n8116), .A2(n8994), .ZN(n7945) );
  INV_X1 U7084 ( .A(n8578), .ZN(n8658) );
  NOR2_X1 U7085 ( .A1(n9109), .A2(n8658), .ZN(n6011) );
  XNOR2_X1 U7086 ( .A(n6013), .B(n6012), .ZN(n7972) );
  NAND2_X1 U7087 ( .A1(n7972), .A2(n8036), .ZN(n6024) );
  INV_X1 U7088 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6014) );
  NOR2_X1 U7089 ( .A1(n6021), .A2(n9131), .ZN(n6019) );
  MUX2_X1 U7090 ( .A(n9131), .B(n6019), .S(P2_IR_REG_16__SCAN_IN), .Z(n6022)
         );
  NOR2_X1 U7091 ( .A1(n6022), .A2(n5518), .ZN(n8726) );
  AOI22_X1 U7092 ( .A1(n6072), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6583), .B2(
        n8726), .ZN(n6023) );
  NAND2_X1 U7093 ( .A1(n8029), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7094 ( .A1(n6131), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7095 ( .A1(n6025), .A2(n8579), .ZN(n6026) );
  AND2_X1 U7096 ( .A1(n6039), .A2(n6026), .ZN(n9002) );
  NAND2_X1 U7097 ( .A1(n5919), .A2(n9002), .ZN(n6028) );
  NAND2_X1 U7098 ( .A1(n8030), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6027) );
  OR2_X1 U7099 ( .A1(n9105), .A2(n8590), .ZN(n8119) );
  NAND2_X1 U7100 ( .A1(n9105), .A2(n8590), .ZN(n8120) );
  NAND2_X1 U7101 ( .A1(n8119), .A2(n8120), .ZN(n9006) );
  INV_X1 U7102 ( .A(n8590), .ZN(n8657) );
  NAND2_X1 U7103 ( .A1(n9105), .A2(n8657), .ZN(n6031) );
  NAND2_X1 U7104 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  NAND2_X1 U7105 ( .A1(n6035), .A2(n6034), .ZN(n7975) );
  NAND2_X1 U7106 ( .A1(n6052), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6036) );
  XNOR2_X1 U7107 ( .A(n6036), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8753) );
  AOI22_X1 U7108 ( .A1(n6072), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6583), .B2(
        n8753), .ZN(n6037) );
  NAND2_X1 U7109 ( .A1(n8029), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7110 ( .A1(n8030), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6043) );
  AND2_X1 U7111 ( .A1(n6039), .A2(n8736), .ZN(n6040) );
  NOR2_X1 U7112 ( .A1(n6055), .A2(n6040), .ZN(n8589) );
  NAND2_X1 U7113 ( .A1(n5919), .A2(n8589), .ZN(n6042) );
  NAND2_X1 U7114 ( .A1(n6131), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7115 ( .A1(n9100), .A2(n8627), .ZN(n8124) );
  INV_X1 U7116 ( .A(n8978), .ZN(n6045) );
  INV_X1 U7117 ( .A(n8627), .ZN(n8969) );
  NAND2_X1 U7118 ( .A1(n6046), .A2(n8627), .ZN(n6047) );
  OR2_X1 U7119 ( .A1(n6049), .A2(n6048), .ZN(n6050) );
  NAND2_X1 U7120 ( .A1(n6051), .A2(n6050), .ZN(n7978) );
  OR2_X1 U7121 ( .A1(n7978), .A2(n6128), .ZN(n6054) );
  XNOR2_X1 U7122 ( .A(n6066), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8762) );
  AOI22_X1 U7123 ( .A1(n6072), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6583), .B2(
        n8762), .ZN(n6053) );
  NOR2_X1 U7124 ( .A1(n6055), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6056) );
  OR2_X1 U7125 ( .A1(n6075), .A2(n6056), .ZN(n8960) );
  INV_X1 U7126 ( .A(n5919), .ZN(n6089) );
  NAND2_X1 U7127 ( .A1(n6131), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6057) );
  OAI21_X1 U7128 ( .B1(n8960), .B2(n6089), .A(n6057), .ZN(n6061) );
  NAND2_X1 U7129 ( .A1(n8030), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6059) );
  NAND2_X1 U7130 ( .A1(n8029), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7131 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  NOR2_X1 U7132 ( .A1(n6061), .A2(n6060), .ZN(n8591) );
  OR2_X1 U7133 ( .A1(n9094), .A2(n8591), .ZN(n6244) );
  NAND2_X1 U7134 ( .A1(n9094), .A2(n8591), .ZN(n6062) );
  NAND2_X1 U7135 ( .A1(n6244), .A2(n6062), .ZN(n8212) );
  INV_X1 U7136 ( .A(n9094), .ZN(n8964) );
  XNOR2_X1 U7137 ( .A(n6064), .B(n6063), .ZN(n7981) );
  NAND2_X1 U7138 ( .A1(n7981), .A2(n8036), .ZN(n6074) );
  NAND2_X1 U7139 ( .A1(n6066), .A2(n6065), .ZN(n6067) );
  INV_X1 U7140 ( .A(n6070), .ZN(n6068) );
  NAND2_X1 U7141 ( .A1(n6068), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n6071) );
  INV_X1 U7142 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6069) );
  AOI22_X1 U7143 ( .A1(n6072), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10815), 
        .B2(n6583), .ZN(n6073) );
  NOR2_X1 U7144 ( .A1(n6075), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6076) );
  OR2_X1 U7145 ( .A1(n6084), .A2(n6076), .ZN(n8951) );
  AOI22_X1 U7146 ( .A1(n8029), .A2(P2_REG1_REG_19__SCAN_IN), .B1(n8030), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7147 ( .A1(n5801), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6077) );
  OAI211_X1 U7148 ( .C1(n8951), .C2(n6089), .A(n6078), .B(n6077), .ZN(n8968)
         );
  INV_X1 U7149 ( .A(n8968), .ZN(n8935) );
  NAND2_X1 U7150 ( .A1(n9091), .A2(n8935), .ZN(n8131) );
  NAND2_X1 U7151 ( .A1(n8129), .A2(n8131), .ZN(n8943) );
  NAND2_X1 U7152 ( .A1(n8944), .A2(n8943), .ZN(n8942) );
  INV_X1 U7153 ( .A(n9091), .ZN(n6079) );
  NAND2_X1 U7154 ( .A1(n8942), .A2(n5663), .ZN(n8926) );
  XNOR2_X1 U7155 ( .A(n6081), .B(n6080), .ZN(n7986) );
  NAND2_X1 U7156 ( .A1(n7986), .A2(n8036), .ZN(n6083) );
  INV_X1 U7157 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7478) );
  OR2_X1 U7158 ( .A1(n5825), .A2(n7478), .ZN(n6082) );
  OR2_X1 U7159 ( .A1(n6084), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7160 ( .A1(n6086), .A2(n6085), .ZN(n8605) );
  AOI22_X1 U7161 ( .A1(n8029), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6131), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7162 ( .A1(n8030), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6087) );
  OAI211_X1 U7163 ( .C1(n8605), .C2(n6089), .A(n6088), .B(n6087), .ZN(n8919)
         );
  OR2_X1 U7164 ( .A1(n9084), .A2(n8919), .ZN(n8138) );
  NAND2_X1 U7165 ( .A1(n9084), .A2(n8919), .ZN(n8141) );
  NAND2_X1 U7166 ( .A1(n9079), .A2(n8934), .ZN(n8149) );
  MUX2_X1 U7167 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n6881), .Z(n6102) );
  XNOR2_X1 U7168 ( .A(n6102), .B(SI_22_), .ZN(n6105) );
  XNOR2_X1 U7169 ( .A(n6106), .B(n6105), .ZN(n7961) );
  NAND2_X1 U7170 ( .A1(n7961), .A2(n8036), .ZN(n6093) );
  INV_X1 U7171 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7680) );
  OR2_X1 U7172 ( .A1(n5825), .A2(n7680), .ZN(n6092) );
  NAND2_X1 U7173 ( .A1(n8030), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7174 ( .A1(n8029), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6100) );
  INV_X1 U7175 ( .A(n6095), .ZN(n6094) );
  NAND2_X1 U7176 ( .A1(n6094), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6110) );
  INV_X1 U7177 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7178 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  AND2_X1 U7179 ( .A1(n6110), .A2(n6097), .ZN(n8904) );
  NAND2_X1 U7180 ( .A1(n5919), .A2(n8904), .ZN(n6099) );
  NAND2_X1 U7181 ( .A1(n5801), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7182 ( .A1(n9074), .A2(n8534), .ZN(n8150) );
  INV_X1 U7183 ( .A(n6102), .ZN(n6103) );
  INV_X1 U7184 ( .A(SI_22_), .ZN(n9650) );
  NAND2_X1 U7185 ( .A1(n6103), .A2(n9650), .ZN(n6104) );
  MUX2_X1 U7186 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n6881), .Z(n6119) );
  XNOR2_X1 U7187 ( .A(n6119), .B(n6120), .ZN(n6117) );
  INV_X1 U7188 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7818) );
  OR2_X1 U7189 ( .A1(n5825), .A2(n7818), .ZN(n6107) );
  NAND2_X1 U7190 ( .A1(n8029), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7191 ( .A1(n6131), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6114) );
  INV_X1 U7192 ( .A(n6110), .ZN(n6108) );
  NAND2_X1 U7193 ( .A1(n6108), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6133) );
  INV_X1 U7194 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7195 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  AND2_X1 U7196 ( .A1(n6133), .A2(n6111), .ZN(n8886) );
  NAND2_X1 U7197 ( .A1(n5919), .A2(n8886), .ZN(n6113) );
  NAND2_X1 U7198 ( .A1(n8030), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7199 ( .A1(n9068), .A2(n8860), .ZN(n8157) );
  INV_X1 U7200 ( .A(n6119), .ZN(n6121) );
  NAND2_X1 U7201 ( .A1(n6121), .A2(n6120), .ZN(n6122) );
  MUX2_X1 U7202 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n6881), .Z(n6124) );
  NAND2_X1 U7203 ( .A1(n6124), .A2(SI_24_), .ZN(n6140) );
  OAI21_X1 U7204 ( .B1(n6124), .B2(SI_24_), .A(n6140), .ZN(n6125) );
  NAND2_X1 U7205 ( .A1(n6126), .A2(n6125), .ZN(n6127) );
  NAND2_X1 U7206 ( .A1(n6141), .A2(n6127), .ZN(n7993) );
  OR2_X1 U7207 ( .A1(n7993), .A2(n6128), .ZN(n6130) );
  INV_X1 U7208 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7889) );
  OR2_X1 U7209 ( .A1(n5825), .A2(n7889), .ZN(n6129) );
  NAND2_X1 U7210 ( .A1(n8029), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7211 ( .A1(n6131), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6137) );
  INV_X1 U7212 ( .A(n6133), .ZN(n6132) );
  NAND2_X1 U7213 ( .A1(n6132), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6146) );
  INV_X1 U7214 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9711) );
  NAND2_X1 U7215 ( .A1(n6133), .A2(n9711), .ZN(n6134) );
  AND2_X1 U7216 ( .A1(n6146), .A2(n6134), .ZN(n8868) );
  NAND2_X1 U7217 ( .A1(n5919), .A2(n8868), .ZN(n6136) );
  NAND2_X1 U7218 ( .A1(n8030), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7219 ( .A1(n9062), .A2(n8568), .ZN(n8158) );
  INV_X1 U7220 ( .A(n8568), .ZN(n8880) );
  NAND2_X1 U7221 ( .A1(n8162), .A2(n8568), .ZN(n6139) );
  MUX2_X1 U7222 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n6881), .Z(n6154) );
  XNOR2_X1 U7223 ( .A(n6154), .B(SI_25_), .ZN(n6152) );
  NAND2_X1 U7224 ( .A1(n9145), .A2(n8036), .ZN(n6144) );
  INV_X1 U7225 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n6142) );
  OR2_X1 U7226 ( .A1(n5825), .A2(n6142), .ZN(n6143) );
  NAND2_X1 U7227 ( .A1(n8030), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7228 ( .A1(n8029), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6150) );
  INV_X1 U7229 ( .A(n6146), .ZN(n6145) );
  NAND2_X1 U7230 ( .A1(n6145), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6160) );
  INV_X1 U7231 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9702) );
  NAND2_X1 U7232 ( .A1(n6146), .A2(n9702), .ZN(n6147) );
  AND2_X1 U7233 ( .A1(n6160), .A2(n6147), .ZN(n8849) );
  NAND2_X1 U7234 ( .A1(n5919), .A2(n8849), .ZN(n6149) );
  NAND2_X1 U7235 ( .A1(n5801), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7236 ( .A1(n9057), .A2(n8861), .ZN(n8170) );
  INV_X1 U7237 ( .A(n9057), .ZN(n8851) );
  INV_X1 U7238 ( .A(n6154), .ZN(n6155) );
  INV_X1 U7239 ( .A(SI_25_), .ZN(n9643) );
  NAND2_X1 U7240 ( .A1(n6155), .A2(n9643), .ZN(n6156) );
  MUX2_X1 U7241 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n6881), .Z(n6168) );
  INV_X1 U7242 ( .A(SI_26_), .ZN(n6169) );
  XNOR2_X1 U7243 ( .A(n6168), .B(n6169), .ZN(n6166) );
  NAND2_X1 U7244 ( .A1(n9142), .A2(n8036), .ZN(n6159) );
  INV_X1 U7245 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9143) );
  OR2_X1 U7246 ( .A1(n5825), .A2(n9143), .ZN(n6158) );
  NAND2_X1 U7247 ( .A1(n8029), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7248 ( .A1(n5801), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6164) );
  INV_X1 U7249 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U7250 ( .A1(n6160), .A2(n9730), .ZN(n6161) );
  NAND2_X1 U7251 ( .A1(n5919), .A2(n8840), .ZN(n6163) );
  NAND2_X1 U7252 ( .A1(n8030), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6162) );
  INV_X1 U7253 ( .A(n8824), .ZN(n8655) );
  INV_X1 U7254 ( .A(n6168), .ZN(n6170) );
  NAND2_X1 U7255 ( .A1(n6170), .A2(n6169), .ZN(n6171) );
  MUX2_X1 U7256 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n6881), .Z(n6186) );
  INV_X1 U7257 ( .A(SI_27_), .ZN(n9638) );
  XNOR2_X1 U7258 ( .A(n6186), .B(n9638), .ZN(n6184) );
  NAND2_X1 U7259 ( .A1(n10451), .A2(n8036), .ZN(n6174) );
  INV_X1 U7260 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9139) );
  OR2_X1 U7261 ( .A1(n5825), .A2(n9139), .ZN(n6173) );
  NAND2_X1 U7262 ( .A1(n8029), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7263 ( .A1(n5801), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6179) );
  INV_X1 U7264 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9679) );
  NAND2_X1 U7265 ( .A1(n6175), .A2(n9679), .ZN(n6176) );
  NAND2_X1 U7266 ( .A1(n6193), .A2(n6176), .ZN(n8521) );
  INV_X1 U7267 ( .A(n8521), .ZN(n8817) );
  NAND2_X1 U7268 ( .A1(n5919), .A2(n8817), .ZN(n6178) );
  NAND2_X1 U7269 ( .A1(n8030), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6177) );
  NAND4_X1 U7270 ( .A1(n6180), .A2(n6179), .A3(n6178), .A4(n6177), .ZN(n8634)
         );
  NAND2_X1 U7271 ( .A1(n8819), .A2(n8634), .ZN(n8175) );
  INV_X1 U7272 ( .A(n8634), .ZN(n6181) );
  NAND2_X1 U7273 ( .A1(n9046), .A2(n6181), .ZN(n8174) );
  NAND2_X1 U7274 ( .A1(n8814), .A2(n8821), .ZN(n6183) );
  NAND2_X1 U7275 ( .A1(n8819), .A2(n6181), .ZN(n6182) );
  INV_X1 U7276 ( .A(n6186), .ZN(n6187) );
  NAND2_X1 U7277 ( .A1(n6187), .A2(n9638), .ZN(n6188) );
  MUX2_X1 U7278 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6881), .Z(n6201) );
  XNOR2_X1 U7279 ( .A(n6201), .B(n9632), .ZN(n6199) );
  NAND2_X1 U7280 ( .A1(n8495), .A2(n8036), .ZN(n6191) );
  INV_X1 U7281 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8496) );
  OR2_X1 U7282 ( .A1(n5825), .A2(n8496), .ZN(n6190) );
  NAND2_X1 U7283 ( .A1(n8029), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7284 ( .A1(n5801), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6197) );
  INV_X1 U7285 ( .A(n6193), .ZN(n6192) );
  NAND2_X1 U7286 ( .A1(n6192), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6210) );
  INV_X1 U7287 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9694) );
  NAND2_X1 U7288 ( .A1(n6193), .A2(n9694), .ZN(n6194) );
  NAND2_X1 U7289 ( .A1(n5919), .A2(n8801), .ZN(n6196) );
  NAND2_X1 U7290 ( .A1(n8030), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6195) );
  INV_X1 U7291 ( .A(n9041), .ZN(n8803) );
  INV_X1 U7292 ( .A(n6201), .ZN(n6202) );
  NAND2_X1 U7293 ( .A1(n6202), .A2(n9632), .ZN(n6203) );
  INV_X1 U7294 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9137) );
  INV_X1 U7295 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10445) );
  MUX2_X1 U7296 ( .A(n9137), .B(n10445), .S(n6507), .Z(n6205) );
  INV_X1 U7297 ( .A(SI_29_), .ZN(n9631) );
  NAND2_X1 U7298 ( .A1(n6205), .A2(n9631), .ZN(n8001) );
  INV_X1 U7299 ( .A(n6205), .ZN(n6206) );
  NAND2_X1 U7300 ( .A1(n6206), .A2(SI_29_), .ZN(n6207) );
  NAND2_X1 U7301 ( .A1(n9136), .A2(n8036), .ZN(n6209) );
  OR2_X1 U7302 ( .A1(n5825), .A2(n9137), .ZN(n6208) );
  NAND2_X1 U7303 ( .A1(n8029), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7304 ( .A1(n5801), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6213) );
  INV_X1 U7305 ( .A(n6210), .ZN(n8790) );
  NAND2_X1 U7306 ( .A1(n5919), .A2(n8790), .ZN(n6212) );
  NAND2_X1 U7307 ( .A1(n8030), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7308 ( .A1(n6228), .A2(n6977), .ZN(n8225) );
  INV_X1 U7309 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6217) );
  INV_X1 U7310 ( .A(n5028), .ZN(n6229) );
  NAND2_X1 U7311 ( .A1(n6219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7312 ( .A1(n5028), .A2(n8227), .ZN(n7158) );
  NAND2_X1 U7313 ( .A1(n6222), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6275) );
  XNOR2_X1 U7314 ( .A(n7158), .B(n8241), .ZN(n6224) );
  NAND2_X1 U7315 ( .A1(n6224), .A2(n6223), .ZN(n8985) );
  NOR2_X1 U7316 ( .A1(n6223), .A2(n8241), .ZN(n6225) );
  NAND2_X1 U7317 ( .A1(n5028), .A2(n6225), .ZN(n10743) );
  NAND2_X1 U7318 ( .A1(n8795), .A2(n11034), .ZN(n6259) );
  INV_X1 U7319 ( .A(n9084), .ZN(n8931) );
  INV_X1 U7320 ( .A(n8107), .ZN(n11010) );
  NAND2_X1 U7321 ( .A1(n7260), .A2(n10784), .ZN(n10803) );
  OR2_X1 U7322 ( .A1(n10803), .A2(n10810), .ZN(n9025) );
  NAND2_X1 U7323 ( .A1(n9027), .A2(n5151), .ZN(n7386) );
  INV_X1 U7324 ( .A(n7516), .ZN(n10979) );
  INV_X1 U7325 ( .A(n7621), .ZN(n10988) );
  NAND2_X1 U7326 ( .A1(n11029), .A2(n7917), .ZN(n7942) );
  NOR2_X2 U7327 ( .A1(n8999), .A2(n9105), .ZN(n8982) );
  INV_X1 U7328 ( .A(n9062), .ZN(n8162) );
  INV_X1 U7329 ( .A(n9052), .ZN(n8832) );
  NOR2_X2 U7330 ( .A1(n9041), .A2(n8815), .ZN(n8800) );
  INV_X1 U7331 ( .A(n8800), .ZN(n6226) );
  INV_X1 U7332 ( .A(n6228), .ZN(n8793) );
  AOI21_X1 U7333 ( .B1(n6228), .B2(n6226), .A(n8781), .ZN(n8789) );
  AND2_X4 U7334 ( .A1(n5028), .A2(n8189), .ZN(n10865) );
  AOI22_X1 U7335 ( .A1(n8789), .A2(n10865), .B1(n10864), .B2(n6228), .ZN(n6257) );
  OR2_X1 U7336 ( .A1(n6223), .A2(n7678), .ZN(n8188) );
  INV_X1 U7337 ( .A(n6690), .ZN(n7160) );
  NAND2_X1 U7338 ( .A1(n7469), .A2(n6675), .ZN(n8041) );
  NAND2_X1 U7339 ( .A1(n6671), .A2(n8041), .ZN(n6231) );
  INV_X1 U7340 ( .A(n7469), .ZN(n6711) );
  NAND2_X1 U7341 ( .A1(n6711), .A2(n6692), .ZN(n6685) );
  NAND2_X1 U7342 ( .A1(n6231), .A2(n6685), .ZN(n8044) );
  INV_X1 U7343 ( .A(n8049), .ZN(n8193) );
  NAND2_X1 U7344 ( .A1(n8044), .A2(n8193), .ZN(n7470) );
  NAND2_X1 U7345 ( .A1(n7470), .A2(n6232), .ZN(n8048) );
  NAND2_X1 U7346 ( .A1(n8048), .A2(n5348), .ZN(n7254) );
  INV_X1 U7347 ( .A(n8051), .ZN(n6233) );
  NOR2_X1 U7348 ( .A1(n7253), .A2(n6233), .ZN(n6234) );
  NAND2_X1 U7349 ( .A1(n7254), .A2(n6234), .ZN(n7252) );
  NAND2_X1 U7350 ( .A1(n7252), .A2(n8057), .ZN(n10806) );
  INV_X1 U7351 ( .A(n6235), .ZN(n8062) );
  INV_X1 U7352 ( .A(n10863), .ZN(n7095) );
  NAND2_X1 U7353 ( .A1(n7095), .A2(n8664), .ZN(n6236) );
  NAND2_X1 U7354 ( .A1(n9013), .A2(n6236), .ZN(n6238) );
  INV_X1 U7355 ( .A(n8664), .ZN(n10887) );
  NAND2_X1 U7356 ( .A1(n10887), .A2(n10863), .ZN(n6237) );
  NAND2_X1 U7357 ( .A1(n8077), .A2(n8076), .ZN(n8078) );
  INV_X1 U7358 ( .A(n7400), .ZN(n8203) );
  INV_X1 U7359 ( .A(n7613), .ZN(n8204) );
  INV_X1 U7360 ( .A(n8206), .ZN(n8092) );
  NAND2_X1 U7361 ( .A1(n7913), .A2(n8208), .ZN(n6240) );
  INV_X1 U7362 ( .A(n8660), .ZN(n8106) );
  NAND2_X1 U7363 ( .A1(n8107), .A2(n8106), .ZN(n6239) );
  INV_X1 U7364 ( .A(n8116), .ZN(n8993) );
  NAND2_X1 U7365 ( .A1(n6242), .A2(n8119), .ZN(n8979) );
  NAND2_X1 U7366 ( .A1(n8979), .A2(n8978), .ZN(n6243) );
  INV_X1 U7367 ( .A(n8943), .ZN(n8946) );
  INV_X1 U7368 ( .A(n8933), .ZN(n8213) );
  INV_X1 U7369 ( .A(n8919), .ZN(n8561) );
  OR2_X1 U7370 ( .A1(n8561), .A2(n9084), .ZN(n6245) );
  NAND2_X1 U7371 ( .A1(n8937), .A2(n6245), .ZN(n8917) );
  NAND2_X1 U7372 ( .A1(n8917), .A2(n8916), .ZN(n8915) );
  INV_X1 U7373 ( .A(n8145), .ZN(n8877) );
  NOR2_X1 U7374 ( .A1(n8876), .A2(n8877), .ZN(n8153) );
  INV_X1 U7375 ( .A(n8833), .ZN(n6248) );
  NOR2_X1 U7376 ( .A1(n8169), .A2(n6248), .ZN(n8173) );
  XNOR2_X1 U7377 ( .A(n8226), .B(n6215), .ZN(n6256) );
  INV_X1 U7378 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7379 ( .A1(n8030), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7380 ( .A1(n5801), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6249) );
  OAI211_X1 U7381 ( .C1(n6252), .C2(n6251), .A(n6250), .B(n6249), .ZN(n8653)
         );
  INV_X1 U7382 ( .A(P2_B_REG_SCAN_IN), .ZN(n9616) );
  NOR2_X1 U7383 ( .A1(n9140), .A2(n9616), .ZN(n6254) );
  NOR2_X1 U7384 ( .A1(n10794), .A2(n6254), .ZN(n8777) );
  INV_X1 U7385 ( .A(n6253), .ZN(n6255) );
  AOI222_X1 U7386 ( .A1(n10808), .A2(n6256), .B1(n8653), .B2(n8777), .C1(n8654), .C2(n9014), .ZN(n8797) );
  NAND2_X1 U7387 ( .A1(n6259), .A2(n6258), .ZN(n6458) );
  NOR4_X1 U7388 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6268) );
  NOR4_X1 U7389 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6267) );
  OR4_X1 U7390 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6265) );
  NOR4_X1 U7391 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6263) );
  NOR4_X1 U7392 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6262) );
  NOR4_X1 U7393 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6261) );
  NOR4_X1 U7394 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6260) );
  NAND4_X1 U7395 ( .A1(n6263), .A2(n6262), .A3(n6261), .A4(n6260), .ZN(n6264)
         );
  NOR4_X1 U7396 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6265), .A4(n6264), .ZN(n6266) );
  AND3_X1 U7397 ( .A1(n6268), .A2(n6267), .A3(n6266), .ZN(n6283) );
  NAND2_X1 U7398 ( .A1(n6269), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7399 ( .A1(n6272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6273) );
  INV_X1 U7400 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7401 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  NAND2_X1 U7402 ( .A1(n6276), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7403 ( .A1(n6285), .A2(n5152), .ZN(n6277) );
  NAND2_X1 U7404 ( .A1(n6277), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6279) );
  INV_X1 U7405 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6278) );
  INV_X1 U7406 ( .A(n7890), .ZN(n6280) );
  AOI22_X1 U7407 ( .A1(P2_B_REG_SCAN_IN), .A2(n7890), .B1(n6280), .B2(n9616), 
        .ZN(n6281) );
  NOR2_X1 U7408 ( .A1(n6283), .A2(n10470), .ZN(n6431) );
  NAND2_X1 U7409 ( .A1(n10468), .A2(n10469), .ZN(n6284) );
  XNOR2_X1 U7410 ( .A(n6285), .B(n5152), .ZN(n6582) );
  OR2_X1 U7411 ( .A1(n10470), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6287) );
  OR2_X1 U7412 ( .A1(n10468), .A2(n10469), .ZN(n6286) );
  NAND2_X1 U7413 ( .A1(n6287), .A2(n6286), .ZN(n6430) );
  NAND3_X1 U7414 ( .A1(n7157), .A2(n10471), .A3(n6430), .ZN(n6288) );
  OR2_X1 U7415 ( .A1(n10470), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6290) );
  INV_X1 U7416 ( .A(n10468), .ZN(n9144) );
  NAND2_X1 U7417 ( .A1(n7890), .A2(n9144), .ZN(n10617) );
  NAND2_X1 U7418 ( .A1(n6458), .A2(n11037), .ZN(n6293) );
  INV_X1 U7419 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6291) );
  OR2_X1 U7420 ( .A1(n11037), .A2(n6291), .ZN(n6292) );
  NAND2_X1 U7421 ( .A1(n6293), .A2(n6292), .ZN(P2_U3549) );
  NAND2_X1 U7422 ( .A1(n6686), .A2(n6350), .ZN(n6699) );
  NAND2_X1 U7423 ( .A1(n7160), .A2(n6303), .ZN(n6294) );
  AND2_X1 U7424 ( .A1(n6699), .A2(n6294), .ZN(n6679) );
  NAND2_X1 U7425 ( .A1(n7469), .A2(n6350), .ZN(n6296) );
  XNOR2_X1 U7426 ( .A(n6295), .B(n6296), .ZN(n6680) );
  NAND2_X1 U7427 ( .A1(n6679), .A2(n6680), .ZN(n6678) );
  INV_X1 U7428 ( .A(n6295), .ZN(n6297) );
  NAND2_X1 U7429 ( .A1(n6297), .A2(n6296), .ZN(n6298) );
  NAND2_X1 U7430 ( .A1(n6678), .A2(n6298), .ZN(n6707) );
  NAND2_X1 U7431 ( .A1(n6350), .A2(n5815), .ZN(n6301) );
  XNOR2_X1 U7432 ( .A(n10744), .B(n6303), .ZN(n6299) );
  XNOR2_X1 U7433 ( .A(n6301), .B(n6299), .ZN(n6709) );
  NAND2_X1 U7434 ( .A1(n6707), .A2(n6709), .ZN(n6708) );
  INV_X1 U7435 ( .A(n6299), .ZN(n6300) );
  NAND2_X1 U7436 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  NAND2_X1 U7437 ( .A1(n6708), .A2(n6302), .ZN(n8539) );
  NOR2_X1 U7438 ( .A1(n6825), .A2(n6696), .ZN(n6305) );
  XNOR2_X1 U7439 ( .A(n6304), .B(n6303), .ZN(n6306) );
  NAND2_X1 U7440 ( .A1(n6305), .A2(n6306), .ZN(n6311) );
  INV_X1 U7441 ( .A(n6305), .ZN(n6308) );
  INV_X1 U7442 ( .A(n6306), .ZN(n6307) );
  NAND2_X1 U7443 ( .A1(n6308), .A2(n6307), .ZN(n6309) );
  NAND2_X1 U7444 ( .A1(n6311), .A2(n6309), .ZN(n8538) );
  OR2_X1 U7445 ( .A1(n10793), .A2(n6696), .ZN(n6314) );
  XNOR2_X1 U7446 ( .A(n10784), .B(n6303), .ZN(n6312) );
  XNOR2_X1 U7447 ( .A(n6314), .B(n6312), .ZN(n6821) );
  INV_X1 U7448 ( .A(n6312), .ZN(n6313) );
  OR2_X1 U7449 ( .A1(n7091), .A2(n6696), .ZN(n6317) );
  XNOR2_X1 U7450 ( .A(n6390), .B(n10810), .ZN(n6315) );
  XNOR2_X1 U7451 ( .A(n6317), .B(n6315), .ZN(n10797) );
  NAND2_X1 U7452 ( .A1(n10796), .A2(n10797), .ZN(n10795) );
  INV_X1 U7453 ( .A(n6315), .ZN(n6316) );
  NAND2_X1 U7454 ( .A1(n6317), .A2(n6316), .ZN(n6318) );
  NAND2_X1 U7455 ( .A1(n10795), .A2(n6318), .ZN(n7086) );
  XNOR2_X1 U7456 ( .A(n10863), .B(n6390), .ZN(n6319) );
  NAND2_X1 U7457 ( .A1(n8664), .A2(n6350), .ZN(n6320) );
  XNOR2_X1 U7458 ( .A(n6319), .B(n6320), .ZN(n7087) );
  INV_X1 U7459 ( .A(n6319), .ZN(n6321) );
  NAND2_X1 U7460 ( .A1(n6321), .A2(n6320), .ZN(n6322) );
  XNOR2_X1 U7461 ( .A(n10895), .B(n6390), .ZN(n6324) );
  NOR2_X1 U7462 ( .A1(n6323), .A2(n6696), .ZN(n6325) );
  NAND2_X1 U7463 ( .A1(n6324), .A2(n6325), .ZN(n6330) );
  INV_X1 U7464 ( .A(n6324), .ZN(n6327) );
  INV_X1 U7465 ( .A(n6325), .ZN(n6326) );
  NAND2_X1 U7466 ( .A1(n6327), .A2(n6326), .ZN(n6328) );
  NAND2_X1 U7467 ( .A1(n6330), .A2(n6328), .ZN(n10892) );
  INV_X1 U7468 ( .A(n10892), .ZN(n6329) );
  XNOR2_X1 U7469 ( .A(n8077), .B(n6303), .ZN(n6331) );
  NOR2_X1 U7470 ( .A1(n8076), .A2(n6696), .ZN(n6332) );
  XNOR2_X1 U7471 ( .A(n6331), .B(n6332), .ZN(n7321) );
  INV_X1 U7472 ( .A(n6331), .ZN(n6333) );
  NAND2_X1 U7473 ( .A1(n6333), .A2(n6332), .ZN(n6334) );
  XNOR2_X1 U7474 ( .A(n10962), .B(n6390), .ZN(n6335) );
  NOR2_X1 U7475 ( .A1(n7507), .A2(n6696), .ZN(n6336) );
  AND2_X1 U7476 ( .A1(n6335), .A2(n6336), .ZN(n10957) );
  INV_X1 U7477 ( .A(n6335), .ZN(n6338) );
  INV_X1 U7478 ( .A(n6336), .ZN(n6337) );
  NAND2_X1 U7479 ( .A1(n6338), .A2(n6337), .ZN(n10958) );
  XNOR2_X1 U7480 ( .A(n7516), .B(n6390), .ZN(n6339) );
  NOR2_X1 U7481 ( .A1(n7562), .A2(n6696), .ZN(n6340) );
  XNOR2_X1 U7482 ( .A(n6339), .B(n6340), .ZN(n7493) );
  XNOR2_X1 U7483 ( .A(n7621), .B(n6303), .ZN(n6341) );
  NOR2_X1 U7484 ( .A1(n7685), .A2(n6696), .ZN(n6342) );
  XNOR2_X1 U7485 ( .A(n6341), .B(n6342), .ZN(n7560) );
  INV_X1 U7486 ( .A(n6341), .ZN(n6343) );
  NAND2_X1 U7487 ( .A1(n6343), .A2(n6342), .ZN(n6344) );
  NAND2_X1 U7488 ( .A1(n6345), .A2(n6344), .ZN(n7681) );
  XNOR2_X1 U7489 ( .A(n7737), .B(n6427), .ZN(n6346) );
  NOR2_X1 U7490 ( .A1(n7915), .A2(n6696), .ZN(n6347) );
  XNOR2_X1 U7491 ( .A(n6346), .B(n6347), .ZN(n7682) );
  INV_X1 U7492 ( .A(n6346), .ZN(n6348) );
  NAND2_X1 U7493 ( .A1(n6348), .A2(n6347), .ZN(n6349) );
  XNOR2_X1 U7494 ( .A(n8107), .B(n6427), .ZN(n6351) );
  NAND2_X1 U7495 ( .A1(n8660), .A2(n6350), .ZN(n6352) );
  NAND2_X1 U7496 ( .A1(n6351), .A2(n6352), .ZN(n6357) );
  INV_X1 U7497 ( .A(n6351), .ZN(n6354) );
  INV_X1 U7498 ( .A(n6352), .ZN(n6353) );
  NAND2_X1 U7499 ( .A1(n6354), .A2(n6353), .ZN(n6355) );
  NAND2_X1 U7500 ( .A1(n6357), .A2(n6355), .ZN(n7895) );
  INV_X1 U7501 ( .A(n7895), .ZN(n6356) );
  NAND2_X1 U7502 ( .A1(n7892), .A2(n6357), .ZN(n7929) );
  XNOR2_X1 U7503 ( .A(n7908), .B(n6427), .ZN(n6358) );
  OR2_X1 U7504 ( .A1(n8646), .A2(n6696), .ZN(n6359) );
  NAND2_X1 U7505 ( .A1(n6358), .A2(n6359), .ZN(n6363) );
  INV_X1 U7506 ( .A(n6358), .ZN(n6361) );
  INV_X1 U7507 ( .A(n6359), .ZN(n6360) );
  NAND2_X1 U7508 ( .A1(n6361), .A2(n6360), .ZN(n6362) );
  AND2_X1 U7509 ( .A1(n6363), .A2(n6362), .ZN(n7931) );
  NAND2_X1 U7510 ( .A1(n7929), .A2(n7931), .ZN(n7930) );
  NAND2_X1 U7511 ( .A1(n7930), .A2(n6363), .ZN(n8642) );
  XNOR2_X1 U7512 ( .A(n9109), .B(n6427), .ZN(n6364) );
  OR2_X1 U7513 ( .A1(n8578), .A2(n6696), .ZN(n6365) );
  NAND2_X1 U7514 ( .A1(n6364), .A2(n6365), .ZN(n6369) );
  INV_X1 U7515 ( .A(n6364), .ZN(n6367) );
  INV_X1 U7516 ( .A(n6365), .ZN(n6366) );
  NAND2_X1 U7517 ( .A1(n6367), .A2(n6366), .ZN(n6368) );
  AND2_X1 U7518 ( .A1(n6369), .A2(n6368), .ZN(n8643) );
  XNOR2_X1 U7519 ( .A(n9105), .B(n6427), .ZN(n6370) );
  OR2_X1 U7520 ( .A1(n8590), .A2(n6696), .ZN(n6371) );
  NAND2_X1 U7521 ( .A1(n6370), .A2(n6371), .ZN(n6375) );
  INV_X1 U7522 ( .A(n6370), .ZN(n6373) );
  INV_X1 U7523 ( .A(n6371), .ZN(n6372) );
  NAND2_X1 U7524 ( .A1(n6373), .A2(n6372), .ZN(n6374) );
  AND2_X1 U7525 ( .A1(n6375), .A2(n6374), .ZN(n8576) );
  XNOR2_X1 U7526 ( .A(n9100), .B(n6427), .ZN(n6377) );
  OR2_X1 U7527 ( .A1(n8627), .A2(n6696), .ZN(n6378) );
  AND2_X1 U7528 ( .A1(n6377), .A2(n6378), .ZN(n8585) );
  INV_X1 U7529 ( .A(n8585), .ZN(n6376) );
  INV_X1 U7530 ( .A(n6377), .ZN(n6380) );
  INV_X1 U7531 ( .A(n6378), .ZN(n6379) );
  NAND2_X1 U7532 ( .A1(n6380), .A2(n6379), .ZN(n8586) );
  NAND2_X1 U7533 ( .A1(n6381), .A2(n8586), .ZN(n8624) );
  XNOR2_X1 U7534 ( .A(n9094), .B(n6427), .ZN(n6382) );
  OR2_X1 U7535 ( .A1(n8591), .A2(n6696), .ZN(n6383) );
  NAND2_X1 U7536 ( .A1(n6382), .A2(n6383), .ZN(n8623) );
  NAND2_X1 U7537 ( .A1(n8624), .A2(n8623), .ZN(n6386) );
  INV_X1 U7538 ( .A(n6382), .ZN(n6385) );
  INV_X1 U7539 ( .A(n6383), .ZN(n6384) );
  NAND2_X1 U7540 ( .A1(n6385), .A2(n6384), .ZN(n8622) );
  XNOR2_X1 U7541 ( .A(n9091), .B(n6390), .ZN(n6389) );
  NAND2_X1 U7542 ( .A1(n8968), .A2(n6350), .ZN(n6387) );
  XNOR2_X1 U7543 ( .A(n6389), .B(n6387), .ZN(n8548) );
  INV_X1 U7544 ( .A(n6387), .ZN(n6388) );
  XNOR2_X1 U7545 ( .A(n9084), .B(n6390), .ZN(n6393) );
  NAND2_X1 U7546 ( .A1(n8919), .A2(n6350), .ZN(n6391) );
  XNOR2_X1 U7547 ( .A(n6393), .B(n6391), .ZN(n8603) );
  INV_X1 U7548 ( .A(n6391), .ZN(n6392) );
  NAND2_X1 U7549 ( .A1(n6393), .A2(n6392), .ZN(n6394) );
  NAND2_X1 U7550 ( .A1(n6395), .A2(n6394), .ZN(n8558) );
  XNOR2_X1 U7551 ( .A(n9079), .B(n6427), .ZN(n6396) );
  NOR2_X1 U7552 ( .A1(n8934), .A2(n6696), .ZN(n6397) );
  XNOR2_X1 U7553 ( .A(n6396), .B(n6397), .ZN(n8557) );
  NAND2_X1 U7554 ( .A1(n8558), .A2(n8557), .ZN(n6400) );
  INV_X1 U7555 ( .A(n6396), .ZN(n6398) );
  NAND2_X1 U7556 ( .A1(n6398), .A2(n6397), .ZN(n6399) );
  XNOR2_X1 U7557 ( .A(n9074), .B(n6427), .ZN(n6401) );
  OR2_X1 U7558 ( .A1(n8534), .A2(n6696), .ZN(n6402) );
  NAND2_X1 U7559 ( .A1(n6401), .A2(n6402), .ZN(n8527) );
  INV_X1 U7560 ( .A(n6401), .ZN(n6404) );
  INV_X1 U7561 ( .A(n6402), .ZN(n6403) );
  NAND2_X1 U7562 ( .A1(n6404), .A2(n6403), .ZN(n6405) );
  NAND2_X1 U7563 ( .A1(n8527), .A2(n6405), .ZN(n8614) );
  XNOR2_X1 U7564 ( .A(n9068), .B(n6427), .ZN(n8529) );
  OR2_X1 U7565 ( .A1(n8860), .A2(n6696), .ZN(n8528) );
  INV_X1 U7566 ( .A(n8527), .ZN(n6406) );
  AOI21_X1 U7567 ( .B1(n8529), .B2(n8528), .A(n6406), .ZN(n6407) );
  INV_X1 U7568 ( .A(n8529), .ZN(n6409) );
  INV_X1 U7569 ( .A(n8528), .ZN(n6408) );
  XNOR2_X1 U7570 ( .A(n9062), .B(n6427), .ZN(n6410) );
  NOR2_X1 U7571 ( .A1(n8568), .A2(n6696), .ZN(n8596) );
  NAND2_X1 U7572 ( .A1(n8597), .A2(n8596), .ZN(n6414) );
  INV_X1 U7573 ( .A(n6410), .ZN(n6411) );
  NAND2_X1 U7574 ( .A1(n6412), .A2(n6411), .ZN(n6413) );
  NAND2_X1 U7575 ( .A1(n6414), .A2(n6413), .ZN(n8566) );
  XNOR2_X1 U7576 ( .A(n9057), .B(n6427), .ZN(n6415) );
  NOR2_X1 U7577 ( .A1(n8861), .A2(n6696), .ZN(n6416) );
  XNOR2_X1 U7578 ( .A(n6415), .B(n6416), .ZN(n8565) );
  NAND2_X1 U7579 ( .A1(n8566), .A2(n8565), .ZN(n6419) );
  INV_X1 U7580 ( .A(n6415), .ZN(n6417) );
  NAND2_X1 U7581 ( .A1(n6417), .A2(n6416), .ZN(n6418) );
  XNOR2_X1 U7582 ( .A(n9052), .B(n6427), .ZN(n6420) );
  NOR2_X1 U7583 ( .A1(n8824), .A2(n6696), .ZN(n6421) );
  XNOR2_X1 U7584 ( .A(n6420), .B(n6421), .ZN(n8633) );
  INV_X1 U7585 ( .A(n6420), .ZN(n6422) );
  NAND2_X1 U7586 ( .A1(n6422), .A2(n6421), .ZN(n6423) );
  XNOR2_X1 U7587 ( .A(n8819), .B(n6427), .ZN(n6426) );
  NAND2_X1 U7588 ( .A1(n8634), .A2(n6350), .ZN(n6424) );
  XNOR2_X1 U7589 ( .A(n6426), .B(n6424), .ZN(n8520) );
  INV_X1 U7590 ( .A(n6424), .ZN(n6425) );
  NAND2_X1 U7591 ( .A1(n8654), .A2(n6350), .ZN(n6428) );
  MUX2_X1 U7592 ( .A(n8654), .B(n6428), .S(n6427), .Z(n6429) );
  INV_X1 U7593 ( .A(n6437), .ZN(n6435) );
  NAND2_X1 U7594 ( .A1(n7156), .A2(n6456), .ZN(n6438) );
  INV_X1 U7595 ( .A(n6438), .ZN(n6434) );
  INV_X1 U7596 ( .A(n6585), .ZN(n6432) );
  NAND2_X1 U7597 ( .A1(n10471), .A2(n6432), .ZN(n6632) );
  NOR2_X1 U7598 ( .A1(n10864), .A2(n6632), .ZN(n6433) );
  NAND2_X1 U7599 ( .A1(n6435), .A2(n10964), .ZN(n6436) );
  OR2_X2 U7600 ( .A1(n6436), .A2(n9041), .ZN(n6455) );
  NAND2_X1 U7601 ( .A1(n6437), .A2(n10964), .ZN(n6440) );
  NAND2_X1 U7602 ( .A1(n6438), .A2(n7157), .ZN(n6448) );
  AND2_X1 U7603 ( .A1(n6448), .A2(n10471), .ZN(n6677) );
  NAND2_X1 U7604 ( .A1(n6440), .A2(n6439), .ZN(n6441) );
  NAND2_X1 U7605 ( .A1(n6441), .A2(n9041), .ZN(n6454) );
  NAND2_X1 U7606 ( .A1(n8634), .A2(n9014), .ZN(n6442) );
  OAI21_X1 U7607 ( .B1(n6977), .B2(n10794), .A(n6442), .ZN(n8807) );
  NAND2_X1 U7608 ( .A1(n10471), .A2(n6456), .ZN(n6443) );
  OR2_X1 U7609 ( .A1(n8240), .A2(n6443), .ZN(n6444) );
  AOI22_X1 U7610 ( .A1(n8807), .A2(n10955), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6452) );
  NAND2_X1 U7611 ( .A1(n6633), .A2(n6582), .ZN(n6446) );
  NOR2_X1 U7612 ( .A1(n7154), .A2(n6446), .ZN(n6447) );
  NAND2_X1 U7613 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  NAND2_X1 U7614 ( .A1(n8801), .A2(n6450), .ZN(n6451) );
  AND2_X1 U7615 ( .A1(n6452), .A2(n6451), .ZN(n6453) );
  NAND3_X1 U7616 ( .A1(n6455), .A2(n6454), .A3(n6453), .ZN(P2_U3222) );
  NAND2_X1 U7617 ( .A1(n6458), .A2(n11041), .ZN(n6461) );
  INV_X1 U7618 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6459) );
  OR2_X1 U7619 ( .A1(n11041), .A2(n6459), .ZN(n6460) );
  NAND2_X1 U7620 ( .A1(n6461), .A2(n6460), .ZN(P2_U3517) );
  NAND3_X1 U7621 ( .A1(n6537), .A2(n6831), .A3(n7080), .ZN(n6472) );
  NOR2_X1 U7622 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6471) );
  NOR2_X1 U7623 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6470) );
  NOR2_X1 U7624 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6469) );
  NOR2_X1 U7625 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6468) );
  NAND2_X1 U7626 ( .A1(n6475), .A2(n6485), .ZN(n6476) );
  NOR2_X1 U7627 ( .A1(n6479), .A2(n10439), .ZN(n6477) );
  NAND2_X1 U7628 ( .A1(n6479), .A2(n6478), .ZN(n6602) );
  INV_X1 U7629 ( .A(n6602), .ZN(n6480) );
  NOR2_X1 U7630 ( .A1(n6480), .A2(n5656), .ZN(n6481) );
  NAND2_X1 U7631 ( .A1(n6484), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U7632 ( .A1(n6488), .A2(n6485), .ZN(n6486) );
  NAND2_X1 U7633 ( .A1(n6486), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6487) );
  XNOR2_X1 U7634 ( .A(n6487), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6840) );
  XNOR2_X1 U7635 ( .A(n6488), .B(P1_IR_REG_25__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U7636 ( .A1(n5060), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U7637 ( .A1(n6843), .A2(n6491), .ZN(n6492) );
  OR2_X1 U7638 ( .A1(n6911), .A2(n9591), .ZN(n6501) );
  NAND2_X1 U7639 ( .A1(n6499), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U7640 ( .A1(n6501), .A2(n7799), .ZN(n6560) );
  NAND2_X1 U7641 ( .A1(n6895), .A2(n6560), .ZN(n6502) );
  NAND2_X1 U7642 ( .A1(n6502), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X1 U7643 ( .A1(n8021), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9134) );
  AND2_X1 U7644 ( .A1(n8021), .A2(P2_U3152), .ZN(n7816) );
  INV_X2 U7645 ( .A(n7816), .ZN(n9147) );
  OAI222_X1 U7646 ( .A1(n9146), .A2(n6503), .B1(n10637), .B2(P2_U3152), .C1(
        n9147), .C2(n6896), .ZN(P2_U3357) );
  OAI222_X1 U7647 ( .A1(n9146), .A2(n5496), .B1(n6646), .B2(P2_U3152), .C1(
        n9147), .C2(n6882), .ZN(P2_U3356) );
  OAI222_X1 U7648 ( .A1(n9146), .A2(n6504), .B1(n6776), .B2(P2_U3152), .C1(
        n9147), .C2(n7003), .ZN(P2_U3355) );
  NAND2_X1 U7649 ( .A1(n6505), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6506) );
  XNOR2_X1 U7650 ( .A(n6506), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6568) );
  INV_X1 U7651 ( .A(n6568), .ZN(n10016) );
  AND2_X1 U7652 ( .A1(n8021), .A2(P1_U3084), .ZN(n10442) );
  INV_X2 U7653 ( .A(n10442), .ZN(n10454) );
  INV_X1 U7654 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6594) );
  AND2_X1 U7655 ( .A1(n6881), .A2(P1_U3084), .ZN(n10450) );
  INV_X2 U7656 ( .A(n10450), .ZN(n10461) );
  OAI222_X1 U7657 ( .A1(n10016), .A2(P1_U3084), .B1(n10454), .B2(n6594), .C1(
        n7003), .C2(n10461), .ZN(P1_U3350) );
  NAND2_X1 U7658 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6509) );
  INV_X1 U7659 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6508) );
  INV_X1 U7660 ( .A(n6510), .ZN(n6511) );
  INV_X1 U7661 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6589) );
  OAI222_X1 U7662 ( .A1(n10607), .A2(P1_U3084), .B1(n10454), .B2(n6589), .C1(
        n6896), .C2(n10461), .ZN(P1_U3352) );
  OR2_X1 U7663 ( .A1(n6510), .A2(n10439), .ZN(n6512) );
  XNOR2_X1 U7664 ( .A(n6512), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10663) );
  INV_X1 U7665 ( .A(n10663), .ZN(n6883) );
  INV_X1 U7666 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6591) );
  OAI222_X1 U7667 ( .A1(n6883), .A2(P1_U3084), .B1(n10454), .B2(n6591), .C1(
        n6882), .C2(n10461), .ZN(P1_U3351) );
  OAI222_X1 U7668 ( .A1(n9147), .A2(n7059), .B1(n6665), .B2(P2_U3152), .C1(
        n6513), .C2(n9146), .ZN(P2_U3354) );
  NAND2_X1 U7669 ( .A1(n6514), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6517) );
  XNOR2_X1 U7670 ( .A(n6517), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6570) );
  INV_X1 U7671 ( .A(n6570), .ZN(n10692) );
  INV_X1 U7672 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6596) );
  OAI222_X1 U7673 ( .A1(n10692), .A2(P1_U3084), .B1(n10454), .B2(n6596), .C1(
        n7059), .C2(n10461), .ZN(P1_U3349) );
  OAI222_X1 U7674 ( .A1(n9147), .A2(n7218), .B1(n6670), .B2(P2_U3152), .C1(
        n6515), .C2(n9146), .ZN(P2_U3353) );
  NAND2_X1 U7675 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  NAND2_X1 U7676 ( .A1(n6518), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6519) );
  XNOR2_X1 U7677 ( .A(n6519), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6571) );
  INV_X1 U7678 ( .A(n6571), .ZN(n10592) );
  INV_X1 U7679 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7219) );
  OAI222_X1 U7680 ( .A1(P1_U3084), .A2(n10592), .B1(n10461), .B2(n7218), .C1(
        n7219), .C2(n10454), .ZN(P1_U3348) );
  INV_X1 U7681 ( .A(n6785), .ZN(n6752) );
  INV_X1 U7682 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6520) );
  OAI222_X1 U7683 ( .A1(n9147), .A2(n7413), .B1(n6752), .B2(P2_U3152), .C1(
        n6520), .C2(n9146), .ZN(P2_U3351) );
  INV_X1 U7684 ( .A(n6740), .ZN(n6764) );
  INV_X1 U7685 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6521) );
  OAI222_X1 U7686 ( .A1(n9147), .A2(n7331), .B1(n6764), .B2(P2_U3152), .C1(
        n6521), .C2(n9146), .ZN(P2_U3352) );
  OR2_X1 U7687 ( .A1(n6522), .A2(n10439), .ZN(n6523) );
  XNOR2_X1 U7688 ( .A(n6523), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7412) );
  INV_X1 U7689 ( .A(n7412), .ZN(n6575) );
  INV_X1 U7690 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6524) );
  OAI222_X1 U7691 ( .A1(P1_U3084), .A2(n6575), .B1(n10461), .B2(n7413), .C1(
        n6524), .C2(n10454), .ZN(P1_U3346) );
  INV_X1 U7692 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7330) );
  OR2_X1 U7693 ( .A1(n6525), .A2(n10439), .ZN(n6526) );
  XNOR2_X1 U7694 ( .A(n6526), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10525) );
  INV_X1 U7695 ( .A(n10525), .ZN(n7334) );
  OAI222_X1 U7696 ( .A1(n10454), .A2(n7330), .B1(n10461), .B2(n7331), .C1(
        P1_U3084), .C2(n7334), .ZN(P1_U3347) );
  INV_X1 U7697 ( .A(n7522), .ZN(n6529) );
  AOI22_X1 U7698 ( .A1(n6788), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n9134), .ZN(n6527) );
  OAI21_X1 U7699 ( .B1(n6529), .B2(n9147), .A(n6527), .ZN(P2_U3350) );
  INV_X1 U7700 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U7701 ( .A1(n6522), .A2(n6528), .ZN(n6539) );
  NAND2_X1 U7702 ( .A1(n6539), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6544) );
  XNOR2_X1 U7703 ( .A(n6544), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7523) );
  INV_X1 U7704 ( .A(n7523), .ZN(n6624) );
  INV_X1 U7705 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9759) );
  OAI222_X1 U7706 ( .A1(n6624), .A2(P1_U3084), .B1(n10461), .B2(n6529), .C1(
        n9759), .C2(n10454), .ZN(P1_U3345) );
  INV_X1 U7707 ( .A(n6534), .ZN(n6531) );
  INV_X1 U7708 ( .A(n6839), .ZN(n7891) );
  INV_X1 U7709 ( .A(P1_B_REG_SCAN_IN), .ZN(n8012) );
  INV_X1 U7710 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6838) );
  NOR2_X1 U7711 ( .A1(n6531), .A2(n6839), .ZN(n6532) );
  INV_X1 U7712 ( .A(n6840), .ZN(n10457) );
  AOI22_X1 U7713 ( .A1(n10467), .A2(n6838), .B1(n6532), .B2(n10457), .ZN(
        P1_U3440) );
  INV_X1 U7714 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6921) );
  OR2_X1 U7715 ( .A1(n6840), .A2(n10458), .ZN(n6923) );
  INV_X1 U7716 ( .A(n6923), .ZN(n6533) );
  AOI22_X1 U7717 ( .A1(n10467), .A2(n6921), .B1(n6534), .B2(n6533), .ZN(
        P1_U3441) );
  INV_X1 U7718 ( .A(n7532), .ZN(n6547) );
  AOI22_X1 U7719 ( .A1(n8687), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9134), .ZN(n6535) );
  OAI21_X1 U7720 ( .B1(n6547), .B2(n9147), .A(n6535), .ZN(P2_U3349) );
  INV_X1 U7721 ( .A(n7700), .ZN(n6542) );
  AOI22_X1 U7722 ( .A1(n6807), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9134), .ZN(n6536) );
  OAI21_X1 U7723 ( .B1(n6542), .B2(n9147), .A(n6536), .ZN(P2_U3348) );
  INV_X1 U7724 ( .A(n6537), .ZN(n6538) );
  NAND2_X1 U7725 ( .A1(n6549), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6540) );
  XNOR2_X1 U7726 ( .A(n6540), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10550) );
  AOI22_X1 U7727 ( .A1(n10550), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10442), .ZN(n6541) );
  OAI21_X1 U7728 ( .B1(n6542), .B2(n10461), .A(n6541), .ZN(P1_U3343) );
  INV_X1 U7729 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U7730 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  NAND2_X1 U7731 ( .A1(n6545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6546) );
  XNOR2_X1 U7732 ( .A(n6546), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10537) );
  INV_X1 U7733 ( .A(n10537), .ZN(n6955) );
  INV_X1 U7734 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6599) );
  OAI222_X1 U7735 ( .A1(n6955), .A2(P1_U3084), .B1(n10454), .B2(n6599), .C1(
        n6547), .C2(n10461), .ZN(P1_U3344) );
  AOI22_X1 U7736 ( .A1(n6996), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9134), .ZN(n6548) );
  OAI21_X1 U7737 ( .B1(n7744), .B2(n9147), .A(n6548), .ZN(P2_U3347) );
  NAND2_X1 U7738 ( .A1(n6833), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6550) );
  XNOR2_X1 U7739 ( .A(n6550), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10568) );
  INV_X1 U7740 ( .A(n10568), .ZN(n6958) );
  INV_X1 U7741 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9751) );
  OAI222_X1 U7742 ( .A1(P1_U3084), .A2(n6958), .B1(n10461), .B2(n7744), .C1(
        n9751), .C2(n10454), .ZN(P1_U3342) );
  NAND2_X1 U7743 ( .A1(n10525), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6556) );
  INV_X1 U7744 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7240) );
  MUX2_X1 U7745 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n7240), .S(n10525), .Z(n10527) );
  NAND2_X1 U7746 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6571), .ZN(n6555) );
  INV_X1 U7747 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7067) );
  MUX2_X1 U7748 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n7067), .S(n6571), .Z(n10597)
         );
  NOR2_X1 U7749 ( .A1(n6570), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U7750 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n6568), .ZN(n6553) );
  INV_X1 U7751 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6551) );
  MUX2_X1 U7752 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6551), .S(n6568), .Z(n10024)
         );
  INV_X1 U7753 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10721) );
  XNOR2_X1 U7754 ( .A(n10607), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n10614) );
  NAND3_X1 U7755 ( .A1(n10614), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n10612) );
  OAI21_X1 U7756 ( .B1(n10721), .B2(n10607), .A(n10612), .ZN(n10679) );
  INV_X1 U7757 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6876) );
  MUX2_X1 U7758 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6876), .S(n10663), .Z(n10678) );
  NAND2_X1 U7759 ( .A1(n10679), .A2(n10678), .ZN(n10676) );
  NAND2_X1 U7760 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(n10663), .ZN(n6552) );
  NAND2_X1 U7761 ( .A1(n10676), .A2(n6552), .ZN(n10025) );
  NAND2_X1 U7762 ( .A1(n10024), .A2(n10025), .ZN(n10023) );
  NAND2_X1 U7763 ( .A1(n6553), .A2(n10023), .ZN(n10690) );
  INV_X1 U7764 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10781) );
  AOI22_X1 U7765 ( .A1(n6570), .A2(n10781), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n10692), .ZN(n10689) );
  NOR2_X1 U7766 ( .A1(n10690), .A2(n10689), .ZN(n10688) );
  NOR2_X1 U7767 ( .A1(n6554), .A2(n10688), .ZN(n10598) );
  NAND2_X1 U7768 ( .A1(n10597), .A2(n10598), .ZN(n10596) );
  NAND2_X1 U7769 ( .A1(n6555), .A2(n10596), .ZN(n10528) );
  NAND2_X1 U7770 ( .A1(n10527), .A2(n10528), .ZN(n10526) );
  NAND2_X1 U7771 ( .A1(n6556), .A2(n10526), .ZN(n6558) );
  INV_X1 U7772 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7347) );
  MUX2_X1 U7773 ( .A(n7347), .B(P1_REG1_REG_7__SCAN_IN), .S(n7412), .Z(n6557)
         );
  NOR2_X1 U7774 ( .A1(n6558), .A2(n6557), .ZN(n6614) );
  AOI21_X1 U7775 ( .B1(n6558), .B2(n6557), .A(n6614), .ZN(n6581) );
  NAND3_X1 U7776 ( .A1(n6895), .A2(P1_STATE_REG_SCAN_IN), .A3(n6560), .ZN(
        n10519) );
  INV_X1 U7777 ( .A(n10510), .ZN(n10669) );
  OR2_X1 U7778 ( .A1(n10519), .A2(n10669), .ZN(n10694) );
  NAND2_X1 U7779 ( .A1(n10669), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10452) );
  INV_X1 U7780 ( .A(n10452), .ZN(n6559) );
  NAND2_X1 U7781 ( .A1(n6560), .A2(n6559), .ZN(n10559) );
  INV_X1 U7782 ( .A(n10665), .ZN(n10687) );
  NOR2_X1 U7783 ( .A1(n7412), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6561) );
  AOI21_X1 U7784 ( .B1(n7412), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6561), .ZN(
        n6573) );
  NAND2_X1 U7785 ( .A1(n10525), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6562) );
  OAI21_X1 U7786 ( .B1(n10525), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6562), .ZN(
        n10521) );
  NOR2_X1 U7787 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6571), .ZN(n6563) );
  AOI21_X1 U7788 ( .B1(n6571), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6563), .ZN(
        n10591) );
  INV_X1 U7789 ( .A(n10607), .ZN(n6565) );
  AND2_X1 U7790 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n10603) );
  NAND2_X1 U7791 ( .A1(n10604), .A2(n10603), .ZN(n10602) );
  INV_X1 U7792 ( .A(n10602), .ZN(n6564) );
  AOI21_X1 U7793 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n6565), .A(n6564), .ZN(
        n10668) );
  NAND2_X1 U7794 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n10663), .ZN(n6566) );
  OAI21_X1 U7795 ( .B1(n10663), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6566), .ZN(
        n10667) );
  NOR2_X1 U7796 ( .A1(n10668), .A2(n10667), .ZN(n10666) );
  NAND2_X1 U7797 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n6568), .ZN(n6567) );
  OAI21_X1 U7798 ( .B1(n6568), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6567), .ZN(
        n10020) );
  NOR2_X1 U7799 ( .A1(n6570), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6569) );
  AOI21_X1 U7800 ( .B1(n6570), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6569), .ZN(
        n10685) );
  OAI21_X1 U7801 ( .B1(n6570), .B2(P1_REG2_REG_4__SCAN_IN), .A(n10683), .ZN(
        n10590) );
  NAND2_X1 U7802 ( .A1(n10591), .A2(n10590), .ZN(n10589) );
  OAI21_X1 U7803 ( .B1(n6571), .B2(P1_REG2_REG_5__SCAN_IN), .A(n10589), .ZN(
        n10522) );
  NOR2_X1 U7804 ( .A1(n10521), .A2(n10522), .ZN(n10520) );
  AOI21_X1 U7805 ( .B1(n10525), .B2(P1_REG2_REG_6__SCAN_IN), .A(n10520), .ZN(
        n6572) );
  NAND2_X1 U7806 ( .A1(n6572), .A2(n6573), .ZN(n6619) );
  OAI21_X1 U7807 ( .B1(n6573), .B2(n6572), .A(n6619), .ZN(n6577) );
  AND2_X1 U7808 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7449) );
  INV_X1 U7809 ( .A(n10512), .ZN(n6574) );
  NOR2_X1 U7810 ( .A1(n10691), .A2(n6575), .ZN(n6576) );
  AOI211_X1 U7811 ( .C1(n10687), .C2(n6577), .A(n7449), .B(n6576), .ZN(n6580)
         );
  AND2_X1 U7812 ( .A1(n6911), .A2(n7799), .ZN(n6578) );
  NAND2_X1 U7813 ( .A1(n10664), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n6579) );
  OAI211_X1 U7814 ( .C1(n6581), .C2(n10694), .A(n6580), .B(n6579), .ZN(
        P1_U3248) );
  OR2_X1 U7815 ( .A1(n6582), .A2(P2_U3152), .ZN(n8244) );
  INV_X1 U7816 ( .A(n8244), .ZN(n6584) );
  OAI21_X1 U7817 ( .B1(n10471), .B2(n6584), .A(n6583), .ZN(n6587) );
  NAND2_X1 U7818 ( .A1(n10471), .A2(n6585), .ZN(n6586) );
  NOR2_X1 U7819 ( .A1(n10647), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U7820 ( .A1(n7469), .A2(P2_U3966), .ZN(n6588) );
  OAI21_X1 U7821 ( .B1(n6589), .B2(P2_U3966), .A(n6588), .ZN(P2_U3553) );
  NAND2_X1 U7822 ( .A1(n5815), .A2(P2_U3966), .ZN(n6590) );
  OAI21_X1 U7823 ( .B1(n6591), .B2(P2_U3966), .A(n6590), .ZN(P2_U3554) );
  NAND2_X1 U7824 ( .A1(n6592), .A2(P2_U3966), .ZN(n6593) );
  OAI21_X1 U7825 ( .B1(n6594), .B2(P2_U3966), .A(n6593), .ZN(P2_U3555) );
  NAND2_X1 U7826 ( .A1(n8542), .A2(P2_U3966), .ZN(n6595) );
  OAI21_X1 U7827 ( .B1(n6596), .B2(P2_U3966), .A(n6595), .ZN(P2_U3556) );
  INV_X1 U7828 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U7829 ( .A1(n8969), .A2(P2_U3966), .ZN(n6597) );
  OAI21_X1 U7830 ( .B1(n7083), .B2(P2_U3966), .A(n6597), .ZN(P2_U3569) );
  NAND2_X1 U7831 ( .A1(n7323), .A2(P2_U3966), .ZN(n6598) );
  OAI21_X1 U7832 ( .B1(n6599), .B2(P2_U3966), .A(n6598), .ZN(P2_U3561) );
  NAND2_X1 U7833 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n8665), .ZN(n6600) );
  OAI21_X1 U7834 ( .B1(n8934), .B2(n8665), .A(n6600), .ZN(P2_U3573) );
  INV_X1 U7835 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6716) );
  INV_X1 U7836 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U7837 ( .A1(n6602), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6604) );
  INV_X1 U7838 ( .A(n10447), .ZN(n6605) );
  INV_X1 U7839 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7267) );
  OR2_X1 U7840 ( .A1(n5034), .A2(n7267), .ZN(n6611) );
  INV_X1 U7841 ( .A(n8518), .ZN(n6607) );
  NAND2_X1 U7842 ( .A1(n7241), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7349) );
  INV_X1 U7843 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7348) );
  NOR2_X1 U7844 ( .A1(n7349), .A2(n7348), .ZN(n7422) );
  NAND2_X1 U7845 ( .A1(n7422), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7536) );
  NAND2_X1 U7846 ( .A1(n7755), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7763) );
  INV_X1 U7847 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7762) );
  INV_X1 U7848 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7277) );
  AND2_X1 U7849 ( .A1(n7765), .A2(n7277), .ZN(n6606) );
  OR2_X1 U7850 ( .A1(n6606), .A2(n8279), .ZN(n10310) );
  OR2_X1 U7851 ( .A1(n5032), .A2(n10310), .ZN(n6610) );
  NAND2_X1 U7852 ( .A1(n8412), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6609) );
  NAND2_X1 U7853 ( .A1(n7753), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6608) );
  NAND4_X1 U7854 ( .A1(n6611), .A2(n6610), .A3(n6609), .A4(n6608), .ZN(n10293)
         );
  NAND2_X1 U7855 ( .A1(n10293), .A2(P1_U4006), .ZN(n6612) );
  OAI21_X1 U7856 ( .B1(P1_U4006), .B2(n6716), .A(n6612), .ZN(P1_U3569) );
  INV_X1 U7857 ( .A(n7749), .ZN(n6631) );
  AOI22_X1 U7858 ( .A1(n7179), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n9134), .ZN(n6613) );
  OAI21_X1 U7859 ( .B1(n6631), .B2(n9147), .A(n6613), .ZN(P2_U3346) );
  NOR2_X1 U7860 ( .A1(n7412), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6615) );
  NOR2_X1 U7861 ( .A1(n6615), .A2(n6614), .ZN(n6617) );
  INV_X1 U7862 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U7863 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n6624), .B1(n7523), .B2(
        n10927), .ZN(n6616) );
  NOR2_X1 U7864 ( .A1(n6617), .A2(n6616), .ZN(n6953) );
  AOI21_X1 U7865 ( .B1(n6617), .B2(n6616), .A(n6953), .ZN(n6628) );
  NOR2_X1 U7866 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n7523), .ZN(n6618) );
  AOI21_X1 U7867 ( .B1(n7523), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6618), .ZN(
        n6621) );
  OAI21_X1 U7868 ( .B1(n7412), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6619), .ZN(
        n6620) );
  NAND2_X1 U7869 ( .A1(n6621), .A2(n6620), .ZN(n6967) );
  OAI21_X1 U7870 ( .B1(n6621), .B2(n6620), .A(n6967), .ZN(n6626) );
  NAND2_X1 U7871 ( .A1(n10664), .A2(P1_ADDR_REG_8__SCAN_IN), .ZN(n6623) );
  INV_X1 U7872 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6622) );
  OR2_X1 U7873 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6622), .ZN(n7587) );
  OAI211_X1 U7874 ( .C1(n10691), .C2(n6624), .A(n6623), .B(n7587), .ZN(n6625)
         );
  AOI21_X1 U7875 ( .B1(n10687), .B2(n6626), .A(n6625), .ZN(n6627) );
  OAI21_X1 U7876 ( .B1(n6628), .B2(n10694), .A(n6627), .ZN(P1_U3249) );
  OAI21_X1 U7877 ( .B1(n6833), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6719) );
  OR2_X1 U7878 ( .A1(n6719), .A2(n6831), .ZN(n6629) );
  NAND2_X1 U7879 ( .A1(n6719), .A2(n6831), .ZN(n6703) );
  INV_X1 U7880 ( .A(n7750), .ZN(n6965) );
  INV_X1 U7881 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6630) );
  OAI222_X1 U7882 ( .A1(n6965), .A2(P1_U3084), .B1(n10461), .B2(n6631), .C1(
        n6630), .C2(n10454), .ZN(P1_U3341) );
  OAI211_X1 U7883 ( .C1(n6633), .C2(P2_U3152), .A(n6632), .B(n8244), .ZN(n6635) );
  NAND2_X1 U7884 ( .A1(n6635), .A2(n6634), .ZN(n6638) );
  NAND2_X1 U7885 ( .A1(n6638), .A2(n8665), .ZN(n6652) );
  NAND2_X1 U7886 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6823) );
  INV_X1 U7887 ( .A(n6823), .ZN(n6643) );
  INV_X1 U7888 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7047) );
  MUX2_X1 U7889 ( .A(n7047), .B(P2_REG1_REG_3__SCAN_IN), .S(n6776), .Z(n6771)
         );
  INV_X1 U7890 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10749) );
  MUX2_X1 U7891 ( .A(n10749), .B(P2_REG1_REG_2__SCAN_IN), .S(n6646), .Z(n10657) );
  INV_X1 U7892 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6695) );
  MUX2_X1 U7893 ( .A(n6695), .B(P2_REG1_REG_1__SCAN_IN), .S(n10637), .Z(n10643) );
  NAND3_X1 U7894 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n10643), .ZN(n10642) );
  OAI21_X1 U7895 ( .B1(n10637), .B2(n6695), .A(n10642), .ZN(n10658) );
  NAND2_X1 U7896 ( .A1(n10657), .A2(n10658), .ZN(n10655) );
  OAI21_X1 U7897 ( .B1(n6646), .B2(n10749), .A(n10655), .ZN(n6772) );
  NAND2_X1 U7898 ( .A1(n6771), .A2(n6772), .ZN(n6770) );
  OAI21_X1 U7899 ( .B1(n6776), .B2(n7047), .A(n6770), .ZN(n6637) );
  INV_X1 U7900 ( .A(n6637), .ZN(n6641) );
  INV_X1 U7901 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10789) );
  MUX2_X1 U7902 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10789), .S(n6665), .Z(n6640)
         );
  MUX2_X1 U7903 ( .A(n10789), .B(P2_REG1_REG_4__SCAN_IN), .S(n6665), .Z(n6636)
         );
  AND2_X1 U7904 ( .A1(n6637), .A2(n6636), .ZN(n6657) );
  INV_X1 U7905 ( .A(n6638), .ZN(n6639) );
  NAND2_X1 U7906 ( .A1(n6639), .A2(n9140), .ZN(n10624) );
  AOI211_X1 U7907 ( .C1(n6641), .C2(n6640), .A(n6657), .B(n10624), .ZN(n6642)
         );
  AOI211_X1 U7908 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n10647), .A(n6643), .B(
        n6642), .ZN(n6656) );
  INV_X1 U7909 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7258) );
  MUX2_X1 U7910 ( .A(n7258), .B(P2_REG2_REG_4__SCAN_IN), .S(n6665), .Z(n6654)
         );
  INV_X1 U7911 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6650) );
  INV_X1 U7912 ( .A(n6646), .ZN(n10653) );
  INV_X1 U7913 ( .A(n10637), .ZN(n6645) );
  INV_X1 U7914 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10641) );
  INV_X1 U7915 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7167) );
  INV_X1 U7916 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6644) );
  MUX2_X1 U7917 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n6644), .S(n10637), .Z(n10630) );
  NOR3_X1 U7918 ( .A1(n10641), .A2(n7167), .A3(n10630), .ZN(n10631) );
  AOI21_X1 U7919 ( .B1(n6645), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10631), .ZN(
        n10651) );
  INV_X1 U7920 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6647) );
  MUX2_X1 U7921 ( .A(n6647), .B(P2_REG2_REG_2__SCAN_IN), .S(n6646), .Z(n6648)
         );
  INV_X1 U7922 ( .A(n6648), .ZN(n10650) );
  NOR2_X1 U7923 ( .A1(n10651), .A2(n10650), .ZN(n10649) );
  AOI21_X1 U7924 ( .B1(n10653), .B2(P2_REG2_REG_2__SCAN_IN), .A(n10649), .ZN(
        n6769) );
  MUX2_X1 U7925 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6650), .S(n6776), .Z(n6768)
         );
  NOR2_X1 U7926 ( .A1(n6769), .A2(n6768), .ZN(n6767) );
  INV_X1 U7927 ( .A(n6767), .ZN(n6649) );
  OAI21_X1 U7928 ( .B1(n6776), .B2(n6650), .A(n6649), .ZN(n6653) );
  NOR2_X1 U7929 ( .A1(n6253), .A2(n9140), .ZN(n6651) );
  NAND2_X1 U7930 ( .A1(n6652), .A2(n6651), .ZN(n10648) );
  NAND2_X1 U7931 ( .A1(n6654), .A2(n6653), .ZN(n6664) );
  OAI211_X1 U7932 ( .C1(n6654), .C2(n6653), .A(n10622), .B(n6664), .ZN(n6655)
         );
  OAI211_X1 U7933 ( .C1(n10638), .C2(n6665), .A(n6656), .B(n6655), .ZN(
        P2_U3249) );
  INV_X1 U7934 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9622) );
  NOR2_X1 U7935 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9622), .ZN(n6661) );
  INV_X1 U7936 ( .A(n6665), .ZN(n6658) );
  AOI21_X1 U7937 ( .B1(n6658), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6657), .ZN(
        n6743) );
  INV_X1 U7938 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10827) );
  MUX2_X1 U7939 ( .A(n10827), .B(P2_REG1_REG_5__SCAN_IN), .S(n6741), .Z(n6742)
         );
  XNOR2_X1 U7940 ( .A(n6743), .B(n6742), .ZN(n6659) );
  NOR2_X1 U7941 ( .A1(n10624), .A2(n6659), .ZN(n6660) );
  AOI211_X1 U7942 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n10647), .A(n6661), .B(
        n6660), .ZN(n6669) );
  NAND2_X1 U7943 ( .A1(n6741), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6662) );
  OAI21_X1 U7944 ( .B1(n6741), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6662), .ZN(
        n6663) );
  INV_X1 U7945 ( .A(n6663), .ZN(n6667) );
  OAI21_X1 U7946 ( .B1(n6665), .B2(n7258), .A(n6664), .ZN(n6666) );
  NAND2_X1 U7947 ( .A1(n6666), .A2(n6667), .ZN(n6733) );
  OAI211_X1 U7948 ( .C1(n6667), .C2(n6666), .A(n10622), .B(n6733), .ZN(n6668)
         );
  OAI211_X1 U7949 ( .C1(n10638), .C2(n6670), .A(n6669), .B(n6668), .ZN(
        P2_U3250) );
  INV_X1 U7950 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10640) );
  INV_X1 U7951 ( .A(n6671), .ZN(n6687) );
  NAND2_X1 U7952 ( .A1(n6230), .A2(n7160), .ZN(n8040) );
  NAND2_X1 U7953 ( .A1(n6687), .A2(n8040), .ZN(n8047) );
  AND2_X1 U7954 ( .A1(n7469), .A2(n9016), .ZN(n6672) );
  AOI21_X1 U7955 ( .B1(n8047), .B2(n10808), .A(n6672), .ZN(n7162) );
  NAND2_X1 U7956 ( .A1(n8047), .A2(n11034), .ZN(n6673) );
  OAI211_X1 U7957 ( .C1(n5213), .C2(n7160), .A(n7162), .B(n6673), .ZN(n6802)
         );
  NAND2_X1 U7958 ( .A1(n6802), .A2(n11037), .ZN(n6674) );
  OAI21_X1 U7959 ( .B1(n11037), .B2(n10640), .A(n6674), .ZN(P2_U3520) );
  INV_X1 U7960 ( .A(n7154), .ZN(n6676) );
  NAND2_X1 U7961 ( .A1(n6677), .A2(n6676), .ZN(n6713) );
  INV_X1 U7962 ( .A(n6230), .ZN(n6697) );
  OAI22_X1 U7963 ( .A1(n6697), .A2(n10792), .B1(n5816), .B2(n10794), .ZN(n6688) );
  AOI22_X1 U7964 ( .A1(n6713), .A2(P2_REG3_REG_1__SCAN_IN), .B1(n10955), .B2(
        n6688), .ZN(n6683) );
  OAI21_X1 U7965 ( .B1(n6680), .B2(n6679), .A(n6678), .ZN(n6681) );
  NAND2_X1 U7966 ( .A1(n6681), .A2(n10964), .ZN(n6682) );
  OAI211_X1 U7967 ( .C1(n6439), .C2(n6675), .A(n6683), .B(n6682), .ZN(P2_U3224) );
  INV_X1 U7968 ( .A(n7819), .ZN(n6705) );
  INV_X1 U7969 ( .A(n7314), .ZN(n7307) );
  INV_X1 U7970 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6684) );
  OAI222_X1 U7971 ( .A1(n9147), .A2(n6705), .B1(n7307), .B2(P2_U3152), .C1(
        n6684), .C2(n9146), .ZN(P2_U3345) );
  NAND2_X1 U7972 ( .A1(n6685), .A2(n8041), .ZN(n8046) );
  XNOR2_X1 U7973 ( .A(n6686), .B(n8046), .ZN(n7197) );
  XNOR2_X1 U7974 ( .A(n6687), .B(n8046), .ZN(n6689) );
  AOI21_X1 U7975 ( .B1(n6689), .B2(n10808), .A(n6688), .ZN(n7200) );
  NAND2_X1 U7976 ( .A1(n6692), .A2(n6690), .ZN(n6691) );
  AND2_X1 U7977 ( .A1(n7464), .A2(n6691), .ZN(n7192) );
  AOI22_X1 U7978 ( .A1(n7192), .A2(n10865), .B1(n10864), .B2(n6692), .ZN(n6693) );
  OAI211_X1 U7979 ( .C1(n11008), .C2(n7197), .A(n7200), .B(n6693), .ZN(n6799)
         );
  NAND2_X1 U7980 ( .A1(n6799), .A2(n11037), .ZN(n6694) );
  OAI21_X1 U7981 ( .B1(n11037), .B2(n6695), .A(n6694), .ZN(P2_U3521) );
  INV_X1 U7982 ( .A(n10884), .ZN(n8606) );
  OAI21_X1 U7983 ( .B1(n6697), .B2(n6696), .A(n7160), .ZN(n6698) );
  NAND3_X1 U7984 ( .A1(n10964), .A2(n6699), .A3(n6698), .ZN(n6700) );
  OAI21_X1 U7985 ( .B1(n8606), .B2(n6711), .A(n6700), .ZN(n6701) );
  AOI21_X1 U7986 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n6713), .A(n6701), .ZN(
        n6702) );
  OAI21_X1 U7987 ( .B1(n7160), .B2(n6439), .A(n6702), .ZN(P2_U3234) );
  NAND2_X1 U7988 ( .A1(n6703), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6704) );
  XNOR2_X1 U7989 ( .A(n6704), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7820) );
  INV_X1 U7990 ( .A(n7820), .ZN(n6706) );
  INV_X1 U7991 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9753) );
  OAI222_X1 U7992 ( .A1(P1_U3084), .A2(n6706), .B1(n10461), .B2(n6705), .C1(
        n9753), .C2(n10454), .ZN(P1_U3340) );
  OAI21_X1 U7993 ( .B1(n6709), .B2(n6707), .A(n6708), .ZN(n6710) );
  NAND2_X1 U7994 ( .A1(n6710), .A2(n10964), .ZN(n6715) );
  NAND2_X1 U7995 ( .A1(n10955), .A2(n9014), .ZN(n10886) );
  OAI22_X1 U7996 ( .A1(n8606), .A2(n6825), .B1(n6711), .B2(n10886), .ZN(n6712)
         );
  AOI21_X1 U7997 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6713), .A(n6712), .ZN(
        n6714) );
  OAI211_X1 U7998 ( .C1(n10744), .C2(n6439), .A(n6715), .B(n6714), .ZN(
        P2_U3239) );
  INV_X1 U7999 ( .A(n7965), .ZN(n6721) );
  INV_X1 U8000 ( .A(n8693), .ZN(n8700) );
  OAI222_X1 U8001 ( .A1(n9147), .A2(n6721), .B1(n9146), .B2(n6716), .C1(
        P2_U3152), .C2(n8700), .ZN(P2_U3344) );
  INV_X1 U8002 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9750) );
  OR2_X1 U8003 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6717) );
  NAND2_X1 U8004 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n6717), .ZN(n6718) );
  NAND2_X1 U8005 ( .A1(n6719), .A2(n6718), .ZN(n6720) );
  INV_X1 U8006 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9968) );
  XNOR2_X1 U8007 ( .A(n6720), .B(n9968), .ZN(n10035) );
  INV_X1 U8008 ( .A(n10035), .ZN(n7280) );
  OAI222_X1 U8009 ( .A1(n10454), .A2(n9750), .B1(P1_U3084), .B2(n7280), .C1(
        n6721), .C2(n10461), .ZN(P1_U3339) );
  NAND2_X1 U8010 ( .A1(n7712), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6730) );
  NAND2_X1 U8011 ( .A1(n7753), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6729) );
  INV_X1 U8012 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6722) );
  OR2_X1 U8013 ( .A1(n5034), .A2(n6722), .ZN(n6728) );
  INV_X1 U8014 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8325) );
  INV_X1 U8015 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9254) );
  NAND2_X1 U8016 ( .A1(n8353), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U8017 ( .A1(n8368), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8367) );
  NAND2_X1 U8018 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n8377), .ZN(n8388) );
  INV_X1 U8019 ( .A(n8388), .ZN(n6723) );
  NAND2_X1 U8020 ( .A1(n6723), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8390) );
  INV_X1 U8021 ( .A(n8390), .ZN(n6724) );
  NAND2_X1 U8022 ( .A1(n6724), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8410) );
  INV_X1 U8023 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U8024 ( .A1(n8390), .A2(n6725), .ZN(n6726) );
  NAND2_X1 U8025 ( .A1(n8410), .A2(n6726), .ZN(n10128) );
  OR2_X1 U8026 ( .A1(n8432), .A2(n10128), .ZN(n6727) );
  NAND2_X1 U8027 ( .A1(n10144), .A2(P1_U4006), .ZN(n6731) );
  OAI21_X1 U8028 ( .B1(P1_U4006), .B2(n6142), .A(n6731), .ZN(P1_U3580) );
  NAND2_X1 U8029 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n8665), .ZN(n6732) );
  OAI21_X1 U8030 ( .B1(n8861), .B2(n8665), .A(n6732), .ZN(P2_U3577) );
  INV_X1 U8031 ( .A(n6733), .ZN(n6734) );
  AOI21_X1 U8032 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n6741), .A(n6734), .ZN(
        n6757) );
  INV_X1 U8033 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6735) );
  MUX2_X1 U8034 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6735), .S(n6740), .Z(n6736)
         );
  INV_X1 U8035 ( .A(n6736), .ZN(n6756) );
  NOR2_X1 U8036 ( .A1(n6757), .A2(n6756), .ZN(n6755) );
  AOI21_X1 U8037 ( .B1(n6740), .B2(P2_REG2_REG_6__SCAN_IN), .A(n6755), .ZN(
        n6739) );
  NAND2_X1 U8038 ( .A1(n6785), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6737) );
  OAI21_X1 U8039 ( .B1(n6785), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6737), .ZN(
        n6738) );
  NOR2_X1 U8040 ( .A1(n6739), .A2(n6738), .ZN(n6779) );
  AOI211_X1 U8041 ( .C1(n6739), .C2(n6738), .A(n6779), .B(n10648), .ZN(n6754)
         );
  INV_X1 U8042 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10872) );
  MUX2_X1 U8043 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10872), .S(n6740), .Z(n6759)
         );
  NAND2_X1 U8044 ( .A1(n6741), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6745) );
  OR2_X1 U8045 ( .A1(n6743), .A2(n6742), .ZN(n6744) );
  NAND2_X1 U8046 ( .A1(n6745), .A2(n6744), .ZN(n6760) );
  NAND2_X1 U8047 ( .A1(n6759), .A2(n6760), .ZN(n6758) );
  OAI21_X1 U8048 ( .B1(n6764), .B2(n10872), .A(n6758), .ZN(n6748) );
  INV_X1 U8049 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6746) );
  MUX2_X1 U8050 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6746), .S(n6785), .Z(n6747)
         );
  NAND2_X1 U8051 ( .A1(n6747), .A2(n6748), .ZN(n6786) );
  OAI211_X1 U8052 ( .C1(n6748), .C2(n6747), .A(n10656), .B(n6786), .ZN(n6751)
         );
  INV_X1 U8053 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9681) );
  NOR2_X1 U8054 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9681), .ZN(n6749) );
  AOI21_X1 U8055 ( .B1(n10647), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n6749), .ZN(
        n6750) );
  OAI211_X1 U8056 ( .C1(n10638), .C2(n6752), .A(n6751), .B(n6750), .ZN(n6753)
         );
  OR2_X1 U8057 ( .A1(n6754), .A2(n6753), .ZN(P2_U3252) );
  AOI211_X1 U8058 ( .C1(n6757), .C2(n6756), .A(n6755), .B(n10648), .ZN(n6766)
         );
  OAI211_X1 U8059 ( .C1(n6760), .C2(n6759), .A(n10656), .B(n6758), .ZN(n6763)
         );
  NAND2_X1 U8060 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7089) );
  INV_X1 U8061 ( .A(n7089), .ZN(n6761) );
  AOI21_X1 U8062 ( .B1(n10647), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6761), .ZN(
        n6762) );
  OAI211_X1 U8063 ( .C1(n10638), .C2(n6764), .A(n6763), .B(n6762), .ZN(n6765)
         );
  OR2_X1 U8064 ( .A1(n6766), .A2(n6765), .ZN(P2_U3251) );
  AOI211_X1 U8065 ( .C1(n6769), .C2(n6768), .A(n6767), .B(n10648), .ZN(n6778)
         );
  OAI211_X1 U8066 ( .C1(n6772), .C2(n6771), .A(n10656), .B(n6770), .ZN(n6775)
         );
  NOR2_X1 U8067 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10763), .ZN(n6773) );
  AOI21_X1 U8068 ( .B1(n10647), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n6773), .ZN(
        n6774) );
  OAI211_X1 U8069 ( .C1(n10638), .C2(n6776), .A(n6775), .B(n6774), .ZN(n6777)
         );
  OR2_X1 U8070 ( .A1(n6778), .A2(n6777), .ZN(P2_U3248) );
  INV_X1 U8071 ( .A(n6788), .ZN(n8666) );
  INV_X1 U8072 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7370) );
  AOI21_X1 U8073 ( .B1(n6785), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6779), .ZN(
        n8670) );
  XNOR2_X1 U8074 ( .A(n6788), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n8669) );
  OAI21_X1 U8075 ( .B1(n8666), .B2(n7370), .A(n8672), .ZN(n8685) );
  INV_X1 U8076 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7404) );
  MUX2_X1 U8077 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7404), .S(n8687), .Z(n8686)
         );
  NAND2_X1 U8078 ( .A1(n8685), .A2(n8686), .ZN(n8684) );
  INV_X1 U8079 ( .A(n8684), .ZN(n6780) );
  AOI21_X1 U8080 ( .B1(n8687), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6780), .ZN(
        n6784) );
  INV_X1 U8081 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6781) );
  MUX2_X1 U8082 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n6781), .S(n6807), .Z(n6782)
         );
  INV_X1 U8083 ( .A(n6782), .ZN(n6783) );
  NOR2_X1 U8084 ( .A1(n6784), .A2(n6783), .ZN(n6806) );
  AOI211_X1 U8085 ( .C1(n6784), .C2(n6783), .A(n6806), .B(n10648), .ZN(n6798)
         );
  INV_X1 U8086 ( .A(n6807), .ZN(n6811) );
  INV_X1 U8087 ( .A(n8687), .ZN(n6790) );
  INV_X1 U8088 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10975) );
  MUX2_X1 U8089 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10975), .S(n8687), .Z(n8680)
         );
  INV_X1 U8090 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U8091 ( .A1(n6785), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6787) );
  NAND2_X1 U8092 ( .A1(n6787), .A2(n6786), .ZN(n8675) );
  MUX2_X1 U8093 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6789), .S(n6788), .Z(n8674)
         );
  NAND2_X1 U8094 ( .A1(n8675), .A2(n8674), .ZN(n8673) );
  OAI21_X1 U8095 ( .B1(n8666), .B2(n6789), .A(n8673), .ZN(n8681) );
  NAND2_X1 U8096 ( .A1(n8680), .A2(n8681), .ZN(n8679) );
  OAI21_X1 U8097 ( .B1(n6790), .B2(n10975), .A(n8679), .ZN(n6793) );
  INV_X1 U8098 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6791) );
  MUX2_X1 U8099 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6791), .S(n6807), .Z(n6792)
         );
  NAND2_X1 U8100 ( .A1(n6792), .A2(n6793), .ZN(n6810) );
  OAI211_X1 U8101 ( .C1(n6793), .C2(n6792), .A(n10656), .B(n6810), .ZN(n6796)
         );
  INV_X1 U8102 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9687) );
  NOR2_X1 U8103 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9687), .ZN(n6794) );
  AOI21_X1 U8104 ( .B1(n10647), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6794), .ZN(
        n6795) );
  OAI211_X1 U8105 ( .C1(n10638), .C2(n6811), .A(n6796), .B(n6795), .ZN(n6797)
         );
  OR2_X1 U8106 ( .A1(n6798), .A2(n6797), .ZN(P2_U3255) );
  INV_X1 U8107 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6801) );
  NAND2_X1 U8108 ( .A1(n6799), .A2(n11041), .ZN(n6800) );
  OAI21_X1 U8109 ( .B1(n11041), .B2(n6801), .A(n6800), .ZN(P2_U3454) );
  INV_X1 U8110 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U8111 ( .A1(n6802), .A2(n11041), .ZN(n6803) );
  OAI21_X1 U8112 ( .B1(n11041), .B2(n6804), .A(n6803), .ZN(P2_U3451) );
  NOR2_X1 U8113 ( .A1(n6996), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6805) );
  AOI21_X1 U8114 ( .B1(n6996), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6805), .ZN(
        n6809) );
  AOI21_X1 U8115 ( .B1(n6807), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6806), .ZN(
        n6808) );
  NAND2_X1 U8116 ( .A1(n6808), .A2(n6809), .ZN(n6997) );
  OAI21_X1 U8117 ( .B1(n6809), .B2(n6808), .A(n6997), .ZN(n6818) );
  INV_X1 U8118 ( .A(n6996), .ZN(n6987) );
  OAI21_X1 U8119 ( .B1(n6811), .B2(n6791), .A(n6810), .ZN(n6814) );
  INV_X1 U8120 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6812) );
  MUX2_X1 U8121 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6812), .S(n6996), .Z(n6813)
         );
  NAND2_X1 U8122 ( .A1(n6813), .A2(n6814), .ZN(n6986) );
  OAI211_X1 U8123 ( .C1(n6814), .C2(n6813), .A(n10656), .B(n6986), .ZN(n6816)
         );
  INV_X1 U8124 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9719) );
  NOR2_X1 U8125 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9719), .ZN(n7566) );
  AOI21_X1 U8126 ( .B1(n10647), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7566), .ZN(
        n6815) );
  OAI211_X1 U8127 ( .C1(n10638), .C2(n6987), .A(n6816), .B(n6815), .ZN(n6817)
         );
  AOI21_X1 U8128 ( .B1(n10622), .B2(n6818), .A(n6817), .ZN(n6819) );
  INV_X1 U8129 ( .A(n6819), .ZN(P2_U3256) );
  OAI21_X1 U8130 ( .B1(n6821), .B2(n5109), .A(n6820), .ZN(n6822) );
  NAND2_X1 U8131 ( .A1(n6822), .A2(n10964), .ZN(n6829) );
  NAND2_X1 U8132 ( .A1(n10884), .A2(n9015), .ZN(n6824) );
  OAI211_X1 U8133 ( .C1(n6825), .C2(n10886), .A(n6824), .B(n6823), .ZN(n6826)
         );
  AOI21_X1 U8134 ( .B1(n6827), .B2(n6450), .A(n6826), .ZN(n6828) );
  OAI211_X1 U8135 ( .C1(n10784), .C2(n6439), .A(n6829), .B(n6828), .ZN(
        P2_U3232) );
  INV_X1 U8136 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6830) );
  INV_X1 U8137 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9779) );
  NAND4_X1 U8138 ( .A1(n6831), .A2(n6830), .A3(n9968), .A4(n9779), .ZN(n6832)
         );
  NOR2_X1 U8139 ( .A1(n6833), .A2(n6832), .ZN(n7036) );
  OR2_X1 U8140 ( .A1(n7036), .A2(n10439), .ZN(n6834) );
  INV_X1 U8141 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7035) );
  XNOR2_X1 U8142 ( .A(n6834), .B(n7035), .ZN(n10047) );
  INV_X1 U8143 ( .A(n7968), .ZN(n6836) );
  INV_X1 U8144 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6835) );
  OAI222_X1 U8145 ( .A1(n10047), .A2(P1_U3084), .B1(n10461), .B2(n6836), .C1(
        n6835), .C2(n10454), .ZN(P1_U3338) );
  INV_X1 U8146 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6837) );
  INV_X1 U8147 ( .A(n8714), .ZN(n8706) );
  OAI222_X1 U8148 ( .A1(n9146), .A2(n6837), .B1(n9147), .B2(n6836), .C1(
        P2_U3152), .C2(n8706), .ZN(P2_U3343) );
  INV_X1 U8149 ( .A(n6925), .ZN(n6856) );
  NAND2_X1 U8150 ( .A1(n6856), .A2(n6838), .ZN(n6842) );
  OR2_X1 U8151 ( .A1(n6840), .A2(n6839), .ZN(n6841) );
  INV_X1 U8152 ( .A(n7479), .ZN(n7110) );
  OAI21_X1 U8153 ( .B1(n6871), .B2(n6893), .A(n7799), .ZN(n6845) );
  OR2_X1 U8154 ( .A1(n6911), .A2(n6845), .ZN(n7022) );
  OAI21_X1 U8155 ( .B1(n6925), .B2(P1_D_REG_1__SCAN_IN), .A(n6923), .ZN(n6858)
         );
  NOR4_X1 U8156 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6849) );
  NOR4_X1 U8157 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6848) );
  NOR4_X1 U8158 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6847) );
  NOR4_X1 U8159 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6846) );
  AND4_X1 U8160 ( .A1(n6849), .A2(n6848), .A3(n6847), .A4(n6846), .ZN(n6855)
         );
  NOR2_X1 U8161 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n6853) );
  NOR4_X1 U8162 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6852) );
  NOR4_X1 U8163 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6851) );
  NOR4_X1 U8164 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6850) );
  AND4_X1 U8165 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n6850), .ZN(n6854)
         );
  NAND2_X1 U8166 ( .A1(n6855), .A2(n6854), .ZN(n6922) );
  NAND2_X1 U8167 ( .A1(n6856), .A2(n6922), .ZN(n6857) );
  INV_X1 U8168 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6875) );
  NOR2_X1 U8169 ( .A1(n8021), .A2(n6859), .ZN(n6861) );
  XNOR2_X1 U8170 ( .A(n6861), .B(n6860), .ZN(n10463) );
  MUX2_X1 U8171 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10463), .S(n6895), .Z(n7108)
         );
  INV_X1 U8172 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6862) );
  NAND2_X1 U8173 ( .A1(n7712), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6864) );
  NAND2_X1 U8174 ( .A1(n7421), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6863) );
  INV_X1 U8175 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6866) );
  OR2_X1 U8176 ( .A1(n8432), .A2(n6866), .ZN(n6870) );
  INV_X1 U8177 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10611) );
  NAND2_X1 U8178 ( .A1(n7421), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U8179 ( .A1(n5035), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6867) );
  NAND4_X2 U8180 ( .A1(n6870), .A2(n6869), .A3(n6868), .A4(n6867), .ZN(n6910)
         );
  AND2_X1 U8181 ( .A1(n10712), .A2(n6910), .ZN(n9336) );
  NOR2_X1 U8182 ( .A1(n10714), .A2(n9336), .ZN(n9432) );
  INV_X1 U8183 ( .A(n6890), .ZN(n6872) );
  NOR3_X1 U8184 ( .A1(n9432), .A2(n6872), .A3(n7144), .ZN(n6873) );
  AOI21_X1 U8185 ( .B1(n10842), .B2(n7107), .A(n6873), .ZN(n10703) );
  OAI21_X1 U8186 ( .B1(n10712), .B2(n7124), .A(n10703), .ZN(n10417) );
  NAND2_X1 U8187 ( .A1(n10417), .A2(n11054), .ZN(n6874) );
  OAI21_X1 U8188 ( .B1(n11054), .B2(n6875), .A(n6874), .ZN(P1_U3454) );
  INV_X1 U8189 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7120) );
  NAND2_X1 U8190 ( .A1(n7712), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6878) );
  NAND2_X1 U8191 ( .A1(n7421), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6877) );
  NAND2_X1 U8192 ( .A1(n9595), .A2(n7492), .ZN(n7111) );
  NAND2_X1 U8193 ( .A1(n6949), .A2(n9181), .ZN(n6888) );
  OR2_X1 U8194 ( .A1(n5030), .A2(n6882), .ZN(n6885) );
  OR2_X1 U8195 ( .A1(n6895), .A2(n6883), .ZN(n6884) );
  AND3_X2 U8196 ( .A1(n6886), .A2(n6885), .A3(n6884), .ZN(n10736) );
  INV_X1 U8197 ( .A(n7111), .ZN(n6887) );
  NAND2_X1 U8198 ( .A1(n6888), .A2(n5064), .ZN(n6892) );
  AOI21_X1 U8199 ( .B1(n6889), .B2(n9598), .A(n10730), .ZN(n6891) );
  AND2_X1 U8200 ( .A1(n6889), .A2(n6893), .ZN(n6894) );
  AOI22_X1 U8201 ( .A1(n9341), .A2(n9181), .B1(n9182), .B2(n6949), .ZN(n7012)
         );
  XNOR2_X1 U8202 ( .A(n7011), .B(n7012), .ZN(n7009) );
  OR2_X1 U8203 ( .A1(n5029), .A2(n6589), .ZN(n6899) );
  OR2_X1 U8204 ( .A1(n7058), .A2(n6896), .ZN(n6897) );
  INV_X2 U8205 ( .A(n8382), .ZN(n7802) );
  NAND2_X1 U8206 ( .A1(n10726), .A2(n7802), .ZN(n6900) );
  NAND2_X1 U8207 ( .A1(n7107), .A2(n9182), .ZN(n6904) );
  NAND2_X1 U8208 ( .A1(n10726), .A2(n9181), .ZN(n6903) );
  NAND2_X1 U8209 ( .A1(n6904), .A2(n6903), .ZN(n6918) );
  NAND2_X1 U8210 ( .A1(n6917), .A2(n6918), .ZN(n6916) );
  NAND2_X1 U8211 ( .A1(n6910), .A2(n9181), .ZN(n6908) );
  NAND2_X1 U8212 ( .A1(n7108), .A2(n7802), .ZN(n6906) );
  INV_X1 U8213 ( .A(n6911), .ZN(n6905) );
  NAND2_X1 U8214 ( .A1(n6908), .A2(n6907), .ZN(n6979) );
  INV_X1 U8215 ( .A(n6979), .ZN(n6909) );
  NAND2_X1 U8216 ( .A1(n6909), .A2(n8418), .ZN(n6915) );
  NAND2_X1 U8217 ( .A1(n6910), .A2(n9182), .ZN(n6914) );
  AND2_X1 U8218 ( .A1(n6911), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6912) );
  NAND2_X1 U8219 ( .A1(n6980), .A2(n6979), .ZN(n6978) );
  NAND2_X1 U8220 ( .A1(n6915), .A2(n6978), .ZN(n6946) );
  NAND2_X1 U8221 ( .A1(n6916), .A2(n6946), .ZN(n6920) );
  INV_X1 U8222 ( .A(n6917), .ZN(n6945) );
  INV_X1 U8223 ( .A(n6918), .ZN(n6947) );
  NAND2_X1 U8224 ( .A1(n6945), .A2(n6947), .ZN(n6919) );
  NAND2_X1 U8225 ( .A1(n6920), .A2(n6919), .ZN(n7010) );
  XOR2_X1 U8226 ( .A(n7009), .B(n7010), .Z(n6944) );
  NOR2_X1 U8227 ( .A1(n6922), .A2(n6921), .ZN(n6924) );
  OAI21_X1 U8228 ( .B1(n6925), .B2(n6924), .A(n6923), .ZN(n6926) );
  INV_X1 U8229 ( .A(n6926), .ZN(n7109) );
  AND2_X1 U8230 ( .A1(n7109), .A2(n7479), .ZN(n6937) );
  NOR2_X1 U8231 ( .A1(n11048), .A2(n9591), .ZN(n6927) );
  NAND2_X2 U8232 ( .A1(n6932), .A2(n6927), .ZN(n9309) );
  NOR2_X1 U8233 ( .A1(n10915), .A2(n7123), .ZN(n9601) );
  NAND2_X1 U8234 ( .A1(n6932), .A2(n9601), .ZN(n9314) );
  NAND2_X1 U8235 ( .A1(n7239), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U8236 ( .A1(n5035), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6930) );
  OR2_X1 U8237 ( .A1(n5032), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6929) );
  AND4_X2 U8238 ( .A1(n6931), .A2(n6930), .A3(n6929), .A4(n6928), .ZN(n7140)
         );
  INV_X1 U8239 ( .A(n7140), .ZN(n10015) );
  OR2_X1 U8240 ( .A1(n10917), .A2(n7123), .ZN(n6933) );
  CLKBUF_X1 U8241 ( .A(n9318), .Z(n9300) );
  AOI22_X1 U8242 ( .A1(n9289), .A2(n7107), .B1(n10015), .B2(n9300), .ZN(n6943)
         );
  NOR2_X1 U8243 ( .A1(n7124), .A2(n7492), .ZN(n10725) );
  INV_X1 U8244 ( .A(n10725), .ZN(n6938) );
  INV_X1 U8245 ( .A(n6937), .ZN(n6941) );
  NOR2_X1 U8246 ( .A1(n6939), .A2(n6938), .ZN(n6940) );
  NAND2_X1 U8247 ( .A1(n6941), .A2(n6940), .ZN(n7026) );
  NAND2_X1 U8248 ( .A1(n6941), .A2(n11021), .ZN(n7024) );
  NAND3_X1 U8249 ( .A1(n7026), .A2(n7024), .A3(n7480), .ZN(n6982) );
  AOI22_X1 U8250 ( .A1(n9220), .A2(n9341), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n6982), .ZN(n6942) );
  OAI211_X1 U8251 ( .C1(n6944), .C2(n9309), .A(n6943), .B(n6942), .ZN(P1_U3235) );
  XNOR2_X1 U8252 ( .A(n6947), .B(n6946), .ZN(n6948) );
  XNOR2_X1 U8253 ( .A(n6945), .B(n6948), .ZN(n6952) );
  AOI22_X1 U8254 ( .A1(n9289), .A2(n6910), .B1(n9300), .B2(n6949), .ZN(n6951)
         );
  AOI22_X1 U8255 ( .A1(n9220), .A2(n10726), .B1(n6982), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6950) );
  OAI211_X1 U8256 ( .C1(n6952), .C2(n9309), .A(n6951), .B(n6950), .ZN(P1_U3220) );
  INV_X1 U8257 ( .A(n10694), .ZN(n10677) );
  INV_X1 U8258 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7713) );
  NOR2_X1 U8259 ( .A1(n6958), .A2(n7713), .ZN(n6959) );
  INV_X1 U8260 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7545) );
  OR2_X1 U8261 ( .A1(n10550), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6957) );
  INV_X1 U8262 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7556) );
  NOR2_X1 U8263 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n7523), .ZN(n6954) );
  NOR2_X1 U8264 ( .A1(n6954), .A2(n6953), .ZN(n10540) );
  MUX2_X1 U8265 ( .A(n7556), .B(P1_REG1_REG_9__SCAN_IN), .S(n10537), .Z(n10539) );
  NOR2_X1 U8266 ( .A1(n10540), .A2(n10539), .ZN(n10538) );
  AOI21_X1 U8267 ( .B1(n6955), .B2(n7556), .A(n10538), .ZN(n10553) );
  MUX2_X1 U8268 ( .A(n7545), .B(P1_REG1_REG_10__SCAN_IN), .S(n10550), .Z(
        n10552) );
  NOR2_X1 U8269 ( .A1(n10553), .A2(n10552), .ZN(n10551) );
  INV_X1 U8270 ( .A(n10551), .ZN(n6956) );
  NAND2_X1 U8271 ( .A1(n6958), .A2(n7713), .ZN(n10571) );
  OAI21_X1 U8272 ( .B1(n6959), .B2(n10572), .A(n10571), .ZN(n10570) );
  INV_X1 U8273 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7754) );
  MUX2_X1 U8274 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7754), .S(n7750), .Z(n6960)
         );
  NAND2_X1 U8275 ( .A1(n6960), .A2(n10570), .ZN(n7096) );
  OAI21_X1 U8276 ( .B1(n10570), .B2(n6960), .A(n7096), .ZN(n6961) );
  NAND2_X1 U8277 ( .A1(n10677), .A2(n6961), .ZN(n6964) );
  INV_X1 U8278 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6962) );
  NOR2_X1 U8279 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6962), .ZN(n7882) );
  INV_X1 U8280 ( .A(n7882), .ZN(n6963) );
  OAI211_X1 U8281 ( .C1(n10691), .C2(n6965), .A(n6964), .B(n6963), .ZN(n6974)
         );
  NOR2_X1 U8282 ( .A1(n10568), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10564) );
  NAND2_X1 U8283 ( .A1(n10537), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6966) );
  OAI21_X1 U8284 ( .B1(n10537), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6966), .ZN(
        n10533) );
  OAI21_X1 U8285 ( .B1(n7523), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6967), .ZN(
        n10534) );
  NOR2_X1 U8286 ( .A1(n10533), .A2(n10534), .ZN(n10532) );
  AOI21_X1 U8287 ( .B1(n10537), .B2(P1_REG2_REG_9__SCAN_IN), .A(n10532), .ZN(
        n10547) );
  INV_X1 U8288 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6968) );
  MUX2_X1 U8289 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n6968), .S(n10550), .Z(n6969) );
  INV_X1 U8290 ( .A(n6969), .ZN(n10546) );
  NOR2_X1 U8291 ( .A1(n10547), .A2(n10546), .ZN(n10545) );
  AND2_X1 U8292 ( .A1(n10568), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10563) );
  NAND2_X1 U8293 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7750), .ZN(n6970) );
  OAI21_X1 U8294 ( .B1(n7750), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6970), .ZN(
        n6971) );
  NOR2_X1 U8295 ( .A1(n6972), .A2(n6971), .ZN(n7099) );
  AOI211_X1 U8296 ( .C1(n6972), .C2(n6971), .A(n7099), .B(n10665), .ZN(n6973)
         );
  AOI211_X1 U8297 ( .C1(n10664), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n6974), .B(
        n6973), .ZN(n6975) );
  INV_X1 U8298 ( .A(n6975), .ZN(P1_U3253) );
  NAND2_X1 U8299 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8665), .ZN(n6976) );
  OAI21_X1 U8300 ( .B1(n6977), .B2(n8665), .A(n6976), .ZN(P2_U3581) );
  OAI21_X1 U8301 ( .B1(n6980), .B2(n6979), .A(n6978), .ZN(n6981) );
  INV_X1 U8302 ( .A(n6981), .ZN(n10670) );
  INV_X1 U8303 ( .A(n9318), .ZN(n9287) );
  INV_X1 U8304 ( .A(n7107), .ZN(n9338) );
  INV_X1 U8305 ( .A(n6982), .ZN(n6983) );
  OAI22_X1 U8306 ( .A1(n9287), .A2(n9338), .B1(n6983), .B2(n6866), .ZN(n6984)
         );
  AOI21_X1 U8307 ( .B1(n7108), .B2(n9292), .A(n6984), .ZN(n6985) );
  OAI21_X1 U8308 ( .B1(n10670), .B2(n9309), .A(n6985), .ZN(P1_U3230) );
  INV_X1 U8309 ( .A(n7179), .ZN(n7172) );
  NOR2_X1 U8310 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9700), .ZN(n6994) );
  OAI21_X1 U8311 ( .B1(n6987), .B2(n6812), .A(n6986), .ZN(n6991) );
  INV_X1 U8312 ( .A(n6991), .ZN(n6989) );
  INV_X1 U8313 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n11005) );
  MUX2_X1 U8314 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n11005), .S(n7179), .Z(n6988) );
  NAND2_X1 U8315 ( .A1(n6989), .A2(n6988), .ZN(n7170) );
  MUX2_X1 U8316 ( .A(n11005), .B(P2_REG1_REG_12__SCAN_IN), .S(n7179), .Z(n6990) );
  NAND2_X1 U8317 ( .A1(n6991), .A2(n6990), .ZN(n6992) );
  AOI21_X1 U8318 ( .B1(n7170), .B2(n6992), .A(n10624), .ZN(n6993) );
  AOI211_X1 U8319 ( .C1(P2_ADDR_REG_12__SCAN_IN), .C2(n10647), .A(n6994), .B(
        n6993), .ZN(n7002) );
  INV_X1 U8320 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6995) );
  MUX2_X1 U8321 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n6995), .S(n7179), .Z(n7000)
         );
  OR2_X1 U8322 ( .A1(n6996), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6998) );
  NAND2_X1 U8323 ( .A1(n6999), .A2(n7000), .ZN(n7181) );
  OAI211_X1 U8324 ( .C1(n7000), .C2(n6999), .A(n10622), .B(n7181), .ZN(n7001)
         );
  OAI211_X1 U8325 ( .C1(n10638), .C2(n7172), .A(n7002), .B(n7001), .ZN(
        P2_U3257) );
  OR2_X1 U8326 ( .A1(n5030), .A2(n7003), .ZN(n7005) );
  OR2_X1 U8327 ( .A1(n7060), .A2(n6594), .ZN(n7004) );
  NAND2_X1 U8328 ( .A1(n7213), .A2(n7802), .ZN(n7006) );
  OAI21_X1 U8329 ( .B1(n7140), .B2(n9187), .A(n7006), .ZN(n7007) );
  NAND2_X1 U8330 ( .A1(n7213), .A2(n9181), .ZN(n7008) );
  OAI21_X1 U8331 ( .B1(n7140), .B2(n8396), .A(n7008), .ZN(n7053) );
  NAND2_X1 U8332 ( .A1(n7010), .A2(n7009), .ZN(n7015) );
  INV_X1 U8333 ( .A(n7011), .ZN(n7013) );
  NAND2_X1 U8334 ( .A1(n7013), .A2(n7012), .ZN(n7014) );
  NAND2_X1 U8335 ( .A1(n7015), .A2(n7014), .ZN(n7052) );
  XOR2_X1 U8336 ( .A(n7051), .B(n7052), .Z(n7031) );
  XNOR2_X1 U8337 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7142) );
  OR2_X1 U8338 ( .A1(n5032), .A2(n7142), .ZN(n7021) );
  INV_X1 U8339 ( .A(n7421), .ZN(n7016) );
  NAND2_X1 U8340 ( .A1(n7239), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n7020) );
  OR2_X1 U8341 ( .A1(n5034), .A2(n10781), .ZN(n7019) );
  NAND2_X1 U8342 ( .A1(n5035), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n7018) );
  INV_X2 U8343 ( .A(n7292), .ZN(n10014) );
  AOI22_X1 U8344 ( .A1(n9318), .A2(n10014), .B1(n9220), .B2(n7213), .ZN(n7030)
         );
  INV_X1 U8345 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7212) );
  INV_X1 U8346 ( .A(n7022), .ZN(n7023) );
  NAND2_X1 U8347 ( .A1(n7024), .A2(n7023), .ZN(n7025) );
  NAND2_X1 U8348 ( .A1(n7025), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7027) );
  INV_X1 U8349 ( .A(n9315), .ZN(n9303) );
  AND2_X1 U8350 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10018) );
  INV_X1 U8351 ( .A(n6949), .ZN(n9342) );
  NOR2_X1 U8352 ( .A1(n9314), .A2(n9342), .ZN(n7028) );
  AOI211_X1 U8353 ( .C1(n7212), .C2(n9303), .A(n10018), .B(n7028), .ZN(n7029)
         );
  OAI211_X1 U8354 ( .C1(n7031), .C2(n9309), .A(n7030), .B(n7029), .ZN(P1_U3216) );
  INV_X1 U8355 ( .A(n7972), .ZN(n7038) );
  INV_X1 U8356 ( .A(n8726), .ZN(n8733) );
  INV_X1 U8357 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7032) );
  OAI222_X1 U8358 ( .A1(n9147), .A2(n7038), .B1(n8733), .B2(P2_U3152), .C1(
        n7032), .C2(n9146), .ZN(P2_U3342) );
  INV_X1 U8359 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7034) );
  NAND2_X1 U8360 ( .A1(n8634), .A2(P2_U3966), .ZN(n7033) );
  OAI21_X1 U8361 ( .B1(n7034), .B2(P2_U3966), .A(n7033), .ZN(P2_U3579) );
  NAND2_X1 U8362 ( .A1(n7036), .A2(n7035), .ZN(n7037) );
  NAND2_X1 U8363 ( .A1(n7037), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7081) );
  XNOR2_X1 U8364 ( .A(n7081), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10066) );
  INV_X1 U8365 ( .A(n10066), .ZN(n10054) );
  INV_X1 U8366 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9745) );
  OAI222_X1 U8367 ( .A1(P1_U3084), .A2(n10054), .B1(n10461), .B2(n7038), .C1(
        n9745), .C2(n10454), .ZN(P1_U3337) );
  INV_X1 U8368 ( .A(n8753), .ZN(n8744) );
  INV_X1 U8369 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7039) );
  OAI222_X1 U8370 ( .A1(n9147), .A2(n7975), .B1(n8744), .B2(P2_U3152), .C1(
        n7039), .C2(n9146), .ZN(P2_U3341) );
  OAI21_X1 U8371 ( .B1(n7041), .B2(n8054), .A(n7040), .ZN(n10772) );
  INV_X1 U8372 ( .A(n10772), .ZN(n7045) );
  OAI21_X1 U8373 ( .B1(n5348), .B2(n8048), .A(n7254), .ZN(n7042) );
  AOI222_X1 U8374 ( .A1(n10808), .A2(n7042), .B1(n8542), .B2(n9016), .C1(n5815), .C2(n9014), .ZN(n10760) );
  AND2_X1 U8375 ( .A1(n7466), .A2(n10766), .ZN(n7043) );
  NOR2_X1 U8376 ( .A1(n7260), .A2(n7043), .ZN(n10765) );
  AOI22_X1 U8377 ( .A1(n10765), .A2(n10865), .B1(n10864), .B2(n10766), .ZN(
        n7044) );
  OAI211_X1 U8378 ( .C1(n11008), .C2(n7045), .A(n10760), .B(n7044), .ZN(n7048)
         );
  NAND2_X1 U8379 ( .A1(n7048), .A2(n11037), .ZN(n7046) );
  OAI21_X1 U8380 ( .B1(n11037), .B2(n7047), .A(n7046), .ZN(P2_U3523) );
  INV_X1 U8381 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7050) );
  NAND2_X1 U8382 ( .A1(n7048), .A2(n11041), .ZN(n7049) );
  OAI21_X1 U8383 ( .B1(n11041), .B2(n7050), .A(n7049), .ZN(P2_U3460) );
  NAND2_X1 U8384 ( .A1(n7052), .A2(n7051), .ZN(n7057) );
  INV_X1 U8385 ( .A(n7053), .ZN(n7054) );
  NAND2_X1 U8386 ( .A1(n7055), .A2(n7054), .ZN(n7056) );
  OR2_X1 U8387 ( .A1(n5030), .A2(n7059), .ZN(n7062) );
  OR2_X1 U8388 ( .A1(n7060), .A2(n6596), .ZN(n7061) );
  OAI211_X1 U8389 ( .C1(n6895), .C2(n10692), .A(n7062), .B(n7061), .ZN(n7148)
         );
  NAND2_X1 U8390 ( .A1(n7148), .A2(n7802), .ZN(n7063) );
  AND2_X1 U8391 ( .A1(n7148), .A2(n9181), .ZN(n7065) );
  XNOR2_X1 U8392 ( .A(n7223), .B(n7224), .ZN(n7066) );
  XNOR2_X1 U8393 ( .A(n7231), .B(n7066), .ZN(n7079) );
  AOI22_X1 U8394 ( .A1(n9289), .A2(n10015), .B1(n9220), .B2(n7148), .ZN(n7078)
         );
  NAND2_X1 U8395 ( .A1(n7239), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7075) );
  NAND2_X1 U8396 ( .A1(n7712), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n7074) );
  OR2_X1 U8397 ( .A1(n5034), .A2(n7067), .ZN(n7073) );
  INV_X1 U8398 ( .A(n7241), .ZN(n7071) );
  INV_X1 U8399 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7069) );
  NAND2_X1 U8400 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7068) );
  NAND2_X1 U8401 ( .A1(n7069), .A2(n7068), .ZN(n7070) );
  NAND2_X1 U8402 ( .A1(n7071), .A2(n7070), .ZN(n7296) );
  OR2_X1 U8403 ( .A1(n5032), .A2(n7296), .ZN(n7072) );
  AND2_X1 U8404 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n10698) );
  NOR2_X1 U8405 ( .A1(n9315), .A2(n7142), .ZN(n7076) );
  AOI211_X1 U8406 ( .C1(n9300), .C2(n10844), .A(n10698), .B(n7076), .ZN(n7077)
         );
  OAI211_X1 U8407 ( .C1(n7079), .C2(n9309), .A(n7078), .B(n7077), .ZN(P1_U3228) );
  NAND2_X1 U8408 ( .A1(n7081), .A2(n7080), .ZN(n7082) );
  NAND2_X1 U8409 ( .A1(n7082), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7188) );
  XNOR2_X1 U8410 ( .A(n7188), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10078) );
  INV_X1 U8411 ( .A(n10078), .ZN(n7084) );
  OAI222_X1 U8412 ( .A1(n7084), .A2(P1_U3084), .B1(n10454), .B2(n7083), .C1(
        n7975), .C2(n10461), .ZN(P1_U3336) );
  OAI21_X1 U8413 ( .B1(n7087), .B2(n7086), .A(n7085), .ZN(n7088) );
  NAND2_X1 U8414 ( .A1(n7088), .A2(n10964), .ZN(n7094) );
  NAND2_X1 U8415 ( .A1(n10884), .A2(n9017), .ZN(n7090) );
  OAI211_X1 U8416 ( .C1(n7091), .C2(n10886), .A(n7090), .B(n7089), .ZN(n7092)
         );
  AOI21_X1 U8417 ( .B1(n9019), .B2(n6450), .A(n7092), .ZN(n7093) );
  OAI211_X1 U8418 ( .C1(n7095), .C2(n6439), .A(n7094), .B(n7093), .ZN(P2_U3241) );
  INV_X1 U8419 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7106) );
  INV_X1 U8420 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7761) );
  MUX2_X1 U8421 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7761), .S(n7820), .Z(n7098)
         );
  OAI21_X1 U8422 ( .B1(n7750), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7096), .ZN(
        n7097) );
  NAND2_X1 U8423 ( .A1(n7098), .A2(n7097), .ZN(n7269) );
  OAI21_X1 U8424 ( .B1(n7098), .B2(n7097), .A(n7269), .ZN(n7103) );
  AOI21_X1 U8425 ( .B1(n7750), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7099), .ZN(
        n7101) );
  MUX2_X1 U8426 ( .A(n7843), .B(P1_REG2_REG_13__SCAN_IN), .S(n7820), .Z(n7100)
         );
  NOR2_X1 U8427 ( .A1(n7101), .A2(n7100), .ZN(n7274) );
  AOI211_X1 U8428 ( .C1(n7101), .C2(n7100), .A(n7274), .B(n10665), .ZN(n7102)
         );
  AOI21_X1 U8429 ( .B1(n10677), .B2(n7103), .A(n7102), .ZN(n7105) );
  INV_X1 U8430 ( .A(n10691), .ZN(n10662) );
  AND2_X1 U8431 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9266) );
  AOI21_X1 U8432 ( .B1(n10662), .B2(n7820), .A(n9266), .ZN(n7104) );
  OAI211_X1 U8433 ( .C1(n10700), .C2(n7106), .A(n7105), .B(n7104), .ZN(
        P1_U3254) );
  XNOR2_X2 U8434 ( .A(n7107), .B(n10726), .ZN(n10709) );
  AND2_X1 U8435 ( .A1(n6910), .A2(n7108), .ZN(n10708) );
  INV_X1 U8436 ( .A(n9434), .ZN(n7137) );
  XNOR2_X1 U8437 ( .A(n7132), .B(n7137), .ZN(n10735) );
  NAND3_X1 U8438 ( .A1(n7110), .A2(n7480), .A3(n7109), .ZN(n7145) );
  NOR2_X1 U8439 ( .A1(n7111), .A2(n10229), .ZN(n7112) );
  NAND2_X1 U8440 ( .A1(n10942), .A2(n7112), .ZN(n10264) );
  NAND2_X1 U8441 ( .A1(n10709), .A2(n10714), .ZN(n7114) );
  NAND2_X1 U8442 ( .A1(n9338), .A2(n10726), .ZN(n7113) );
  NAND2_X1 U8443 ( .A1(n7114), .A2(n7113), .ZN(n9344) );
  XNOR2_X1 U8444 ( .A(n9344), .B(n7137), .ZN(n7118) );
  NAND2_X1 U8445 ( .A1(n9603), .A2(n10730), .ZN(n7116) );
  NAND2_X1 U8446 ( .A1(n9595), .A2(n9598), .ZN(n7115) );
  NAND2_X2 U8447 ( .A1(n7116), .A2(n7115), .ZN(n10920) );
  OAI22_X1 U8448 ( .A1(n9338), .A2(n10915), .B1(n7140), .B2(n10917), .ZN(n7117) );
  AOI21_X1 U8449 ( .B1(n7118), .B2(n10920), .A(n7117), .ZN(n7119) );
  OAI21_X1 U8450 ( .B1(n10735), .B2(n10923), .A(n7119), .ZN(n10738) );
  NAND2_X1 U8451 ( .A1(n10738), .A2(n10942), .ZN(n7129) );
  INV_X1 U8452 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7121) );
  OAI22_X1 U8453 ( .A1(n10942), .A2(n7121), .B1(n7120), .B2(n10937), .ZN(n7127) );
  AND2_X1 U8454 ( .A1(n10710), .A2(n9341), .ZN(n7122) );
  OR2_X1 U8455 ( .A1(n7209), .A2(n7122), .ZN(n10737) );
  NOR2_X1 U8456 ( .A1(n7124), .A2(n7123), .ZN(n7125) );
  INV_X1 U8457 ( .A(n10932), .ZN(n10702) );
  NOR2_X1 U8458 ( .A1(n10737), .A2(n10702), .ZN(n7126) );
  AOI211_X1 U8459 ( .C1(n10317), .C2(n9341), .A(n7127), .B(n7126), .ZN(n7128)
         );
  OAI211_X1 U8460 ( .C1(n10735), .C2(n10264), .A(n7129), .B(n7128), .ZN(
        P1_U3289) );
  NAND2_X1 U8461 ( .A1(n10923), .A2(n10229), .ZN(n7130) );
  AND2_X1 U8462 ( .A1(n8418), .A2(n7130), .ZN(n7131) );
  NAND2_X1 U8463 ( .A1(n7132), .A2(n9434), .ZN(n7134) );
  NAND2_X1 U8464 ( .A1(n9342), .A2(n10736), .ZN(n7133) );
  NAND2_X1 U8465 ( .A1(n7134), .A2(n7133), .ZN(n7202) );
  NAND2_X1 U8466 ( .A1(n7140), .A2(n7213), .ZN(n9403) );
  INV_X1 U8467 ( .A(n7213), .ZN(n10752) );
  NAND2_X1 U8468 ( .A1(n10752), .A2(n10015), .ZN(n9345) );
  NAND2_X1 U8469 ( .A1(n9403), .A2(n9345), .ZN(n7201) );
  NAND2_X1 U8470 ( .A1(n7202), .A2(n7201), .ZN(n7136) );
  NAND2_X1 U8471 ( .A1(n7140), .A2(n10752), .ZN(n7135) );
  NAND2_X1 U8472 ( .A1(n7136), .A2(n7135), .ZN(n7291) );
  NAND2_X1 U8473 ( .A1(n7292), .A2(n7148), .ZN(n9402) );
  INV_X1 U8474 ( .A(n7148), .ZN(n10777) );
  NAND2_X1 U8475 ( .A1(n10777), .A2(n10014), .ZN(n9404) );
  XNOR2_X1 U8476 ( .A(n7291), .B(n7290), .ZN(n10780) );
  INV_X1 U8477 ( .A(n10780), .ZN(n7151) );
  NAND2_X1 U8478 ( .A1(n9344), .A2(n7137), .ZN(n7138) );
  NAND2_X1 U8479 ( .A1(n9342), .A2(n9341), .ZN(n9339) );
  INV_X1 U8480 ( .A(n7201), .ZN(n7203) );
  NAND2_X1 U8481 ( .A1(n9400), .A2(n7203), .ZN(n7139) );
  NAND2_X1 U8482 ( .A1(n7139), .A2(n9403), .ZN(n7286) );
  XNOR2_X1 U8483 ( .A(n7286), .B(n7290), .ZN(n7141) );
  INV_X1 U8484 ( .A(n10920), .ZN(n10848) );
  OAI222_X1 U8485 ( .A1(n10917), .A2(n7356), .B1(n7141), .B2(n10848), .C1(
        n10915), .C2(n7140), .ZN(n10778) );
  NAND2_X1 U8486 ( .A1(n10778), .A2(n10942), .ZN(n7150) );
  INV_X1 U8487 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7143) );
  OAI22_X1 U8488 ( .A1(n10942), .A2(n7143), .B1(n7142), .B2(n10937), .ZN(n7147) );
  AND2_X1 U8489 ( .A1(n7209), .A2(n10752), .ZN(n7211) );
  NAND2_X1 U8490 ( .A1(n7211), .A2(n10777), .ZN(n7299) );
  OAI211_X1 U8491 ( .C1(n7211), .C2(n10777), .A(n10711), .B(n7299), .ZN(n10775) );
  NOR2_X1 U8492 ( .A1(n7145), .A2(n10730), .ZN(n10281) );
  INV_X1 U8493 ( .A(n10281), .ZN(n10313) );
  NOR2_X1 U8494 ( .A1(n10775), .A2(n10313), .ZN(n7146) );
  AOI211_X1 U8495 ( .C1(n10317), .C2(n7148), .A(n7147), .B(n7146), .ZN(n7149)
         );
  OAI211_X1 U8496 ( .C1(n10300), .C2(n7151), .A(n7150), .B(n7149), .ZN(
        P1_U3287) );
  NAND2_X1 U8497 ( .A1(n7152), .A2(n10471), .ZN(n7153) );
  NOR2_X1 U8498 ( .A1(n7154), .A2(n7153), .ZN(n7155) );
  NAND2_X1 U8499 ( .A1(n7156), .A2(n7155), .ZN(n7159) );
  INV_X1 U8500 ( .A(n10471), .ZN(n8239) );
  OR2_X1 U8501 ( .A1(n7158), .A2(n6223), .ZN(n7459) );
  NAND2_X1 U8502 ( .A1(n8985), .A2(n7459), .ZN(n10817) );
  NOR2_X2 U8503 ( .A1(n7159), .A2(n6350), .ZN(n10764) );
  INV_X1 U8504 ( .A(n10764), .ZN(n8788) );
  NOR2_X1 U8505 ( .A1(n5028), .A2(n5213), .ZN(n10811) );
  AOI21_X1 U8506 ( .B1(n8788), .B2(n8963), .A(n7160), .ZN(n7161) );
  AOI21_X1 U8507 ( .B1(n9024), .B2(n8047), .A(n7161), .ZN(n7166) );
  INV_X1 U8508 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7163) );
  OAI21_X1 U8509 ( .B1(n7163), .B2(n8987), .A(n7162), .ZN(n7164) );
  NAND2_X1 U8510 ( .A1(n7164), .A2(n10818), .ZN(n7165) );
  OAI211_X1 U8511 ( .C1(n7167), .C2(n10818), .A(n7166), .B(n7165), .ZN(
        P2_U3296) );
  INV_X1 U8512 ( .A(n10638), .ZN(n10654) );
  INV_X1 U8513 ( .A(n10647), .ZN(n7169) );
  INV_X1 U8514 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7168) );
  NAND2_X1 U8515 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3152), .ZN(n7896) );
  OAI21_X1 U8516 ( .B1(n7169), .B2(n7168), .A(n7896), .ZN(n7177) );
  INV_X1 U8517 ( .A(n7170), .ZN(n7171) );
  AOI21_X1 U8518 ( .B1(n11005), .B2(n7172), .A(n7171), .ZN(n7174) );
  INV_X1 U8519 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U8520 ( .A1(n7314), .A2(n11016), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7307), .ZN(n7173) );
  NOR2_X1 U8521 ( .A1(n7174), .A2(n7173), .ZN(n7306) );
  AOI21_X1 U8522 ( .B1(n7174), .B2(n7173), .A(n7306), .ZN(n7175) );
  NOR2_X1 U8523 ( .A1(n7175), .A2(n10624), .ZN(n7176) );
  AOI211_X1 U8524 ( .C1(n10654), .C2(n7314), .A(n7177), .B(n7176), .ZN(n7186)
         );
  NOR2_X1 U8525 ( .A1(n7314), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7178) );
  AOI21_X1 U8526 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n7314), .A(n7178), .ZN(
        n7183) );
  NAND2_X1 U8527 ( .A1(n7179), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7180) );
  NAND2_X1 U8528 ( .A1(n7182), .A2(n7183), .ZN(n7313) );
  OAI21_X1 U8529 ( .B1(n7183), .B2(n7182), .A(n7313), .ZN(n7184) );
  NAND2_X1 U8530 ( .A1(n10622), .A2(n7184), .ZN(n7185) );
  NAND2_X1 U8531 ( .A1(n7186), .A2(n7185), .ZN(P2_U3258) );
  INV_X1 U8532 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7187) );
  NAND2_X1 U8533 ( .A1(n7188), .A2(n7187), .ZN(n7189) );
  NAND2_X1 U8534 ( .A1(n7189), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7190) );
  XNOR2_X1 U8535 ( .A(n7190), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10586) );
  INV_X1 U8536 ( .A(n10586), .ZN(n10073) );
  INV_X1 U8537 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9746) );
  OAI222_X1 U8538 ( .A1(P1_U3084), .A2(n10073), .B1(n10461), .B2(n7978), .C1(
        n9746), .C2(n10454), .ZN(P1_U3335) );
  INV_X1 U8539 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7191) );
  INV_X1 U8540 ( .A(n8762), .ZN(n8760) );
  OAI222_X1 U8541 ( .A1(n9146), .A2(n7191), .B1(n8760), .B2(P2_U3152), .C1(
        n9147), .C2(n7978), .ZN(P2_U3340) );
  INV_X2 U8542 ( .A(n10818), .ZN(n10821) );
  NAND2_X1 U8543 ( .A1(n10764), .A2(n7192), .ZN(n7194) );
  NAND2_X1 U8544 ( .A1(n10813), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7193) );
  OAI211_X1 U8545 ( .C1(n6644), .C2(n10818), .A(n7194), .B(n7193), .ZN(n7196)
         );
  NOR2_X1 U8546 ( .A1(n8963), .A2(n6675), .ZN(n7195) );
  NOR2_X1 U8547 ( .A1(n7196), .A2(n7195), .ZN(n7199) );
  OR2_X1 U8548 ( .A1(n9008), .A2(n7197), .ZN(n7198) );
  OAI211_X1 U8549 ( .C1(n7200), .C2(n10821), .A(n7199), .B(n7198), .ZN(
        P2_U3295) );
  XNOR2_X1 U8550 ( .A(n7202), .B(n7201), .ZN(n10755) );
  INV_X1 U8551 ( .A(n10923), .ZN(n10840) );
  NAND2_X1 U8552 ( .A1(n10755), .A2(n10840), .ZN(n7208) );
  XNOR2_X1 U8553 ( .A(n9400), .B(n7203), .ZN(n7206) );
  NAND2_X1 U8554 ( .A1(n6949), .A2(n10843), .ZN(n7204) );
  OAI21_X1 U8555 ( .B1(n7292), .B2(n10917), .A(n7204), .ZN(n7205) );
  AOI21_X1 U8556 ( .B1(n7206), .B2(n10920), .A(n7205), .ZN(n7207) );
  AND2_X1 U8557 ( .A1(n7208), .A2(n7207), .ZN(n10757) );
  INV_X1 U8558 ( .A(n10264), .ZN(n10933) );
  NOR2_X1 U8559 ( .A1(n7209), .A2(n10752), .ZN(n7210) );
  OR2_X1 U8560 ( .A1(n7211), .A2(n7210), .ZN(n10753) );
  INV_X1 U8561 ( .A(n10937), .ZN(n10724) );
  AOI22_X1 U8562 ( .A1(n10296), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10724), .B2(
        n7212), .ZN(n7215) );
  NAND2_X1 U8563 ( .A1(n10317), .A2(n7213), .ZN(n7214) );
  OAI211_X1 U8564 ( .C1(n10753), .C2(n10702), .A(n7215), .B(n7214), .ZN(n7216)
         );
  AOI21_X1 U8565 ( .B1(n10755), .B2(n10933), .A(n7216), .ZN(n7217) );
  OAI21_X1 U8566 ( .B1(n10757), .B2(n10296), .A(n7217), .ZN(P1_U3288) );
  OR2_X1 U8567 ( .A1(n5030), .A2(n7218), .ZN(n7221) );
  OR2_X1 U8568 ( .A1(n7060), .A2(n7219), .ZN(n7220) );
  OAI211_X1 U8569 ( .C1(n6895), .C2(n10592), .A(n7221), .B(n7220), .ZN(n7483)
         );
  NAND2_X1 U8570 ( .A1(n7483), .A2(n9181), .ZN(n7222) );
  OAI21_X1 U8571 ( .B1(n7356), .B2(n8396), .A(n7222), .ZN(n7327) );
  INV_X1 U8572 ( .A(n7223), .ZN(n7226) );
  INV_X1 U8573 ( .A(n7224), .ZN(n7225) );
  NAND2_X1 U8574 ( .A1(n7226), .A2(n7225), .ZN(n7230) );
  NAND2_X1 U8575 ( .A1(n7483), .A2(n7802), .ZN(n7227) );
  OAI21_X1 U8576 ( .B1(n7356), .B2(n9187), .A(n7227), .ZN(n7228) );
  XNOR2_X1 U8577 ( .A(n7228), .B(n9185), .ZN(n7233) );
  AND2_X1 U8578 ( .A1(n7230), .A2(n7233), .ZN(n7229) );
  NAND2_X1 U8579 ( .A1(n7231), .A2(n7230), .ZN(n7237) );
  INV_X1 U8580 ( .A(n7232), .ZN(n7235) );
  INV_X1 U8581 ( .A(n7233), .ZN(n7234) );
  AND2_X1 U8582 ( .A1(n7235), .A2(n7234), .ZN(n7236) );
  NAND2_X1 U8583 ( .A1(n7328), .A2(n7329), .ZN(n7238) );
  XOR2_X1 U8584 ( .A(n7327), .B(n7238), .Z(n7249) );
  AOI22_X1 U8585 ( .A1(n9289), .A2(n10014), .B1(n9292), .B2(n7483), .ZN(n7248)
         );
  NAND2_X1 U8586 ( .A1(n5035), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n7245) );
  NAND2_X1 U8587 ( .A1(n7239), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7244) );
  OR2_X1 U8588 ( .A1(n5034), .A2(n7240), .ZN(n7243) );
  OAI21_X1 U8589 ( .B1(n7241), .B2(P1_REG3_REG_6__SCAN_IN), .A(n7349), .ZN(
        n10856) );
  OR2_X1 U8590 ( .A1(n5032), .A2(n10856), .ZN(n7242) );
  AND2_X1 U8591 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10594) );
  NOR2_X1 U8592 ( .A1(n9315), .A2(n7296), .ZN(n7246) );
  AOI211_X1 U8593 ( .C1(n9318), .C2(n10013), .A(n10594), .B(n7246), .ZN(n7247)
         );
  OAI211_X1 U8594 ( .C1(n7249), .C2(n9309), .A(n7248), .B(n7247), .ZN(P1_U3225) );
  OAI21_X1 U8595 ( .B1(n7251), .B2(n7253), .A(n7250), .ZN(n10788) );
  INV_X1 U8596 ( .A(n10788), .ZN(n7266) );
  NAND2_X1 U8597 ( .A1(n7252), .A2(n10808), .ZN(n7257) );
  INV_X1 U8598 ( .A(n7253), .ZN(n8194) );
  AOI21_X1 U8599 ( .B1(n7254), .B2(n8051), .A(n8194), .ZN(n7256) );
  AOI22_X1 U8600 ( .A1(n9014), .A2(n6592), .B1(n9015), .B2(n9016), .ZN(n7255)
         );
  OAI21_X1 U8601 ( .B1(n7257), .B2(n7256), .A(n7255), .ZN(n10786) );
  NAND2_X1 U8602 ( .A1(n10786), .A2(n10818), .ZN(n7265) );
  OAI22_X1 U8603 ( .A1(n7259), .A2(n8987), .B1(n7258), .B2(n10818), .ZN(n7262)
         );
  OAI21_X1 U8604 ( .B1(n7260), .B2(n10784), .A(n10803), .ZN(n10785) );
  NOR2_X1 U8605 ( .A1(n8788), .A2(n10785), .ZN(n7261) );
  AOI211_X1 U8606 ( .C1(n10767), .C2(n7263), .A(n7262), .B(n7261), .ZN(n7264)
         );
  OAI211_X1 U8607 ( .C1(n7266), .C2(n9008), .A(n7265), .B(n7264), .ZN(P2_U3292) );
  NOR2_X1 U8608 ( .A1(n7280), .A2(n7267), .ZN(n7268) );
  AOI21_X1 U8609 ( .B1(n7280), .B2(n7267), .A(n7268), .ZN(n7271) );
  OAI21_X1 U8610 ( .B1(n7820), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7269), .ZN(
        n7270) );
  NAND2_X1 U8611 ( .A1(n7271), .A2(n7270), .ZN(n10034) );
  OAI21_X1 U8612 ( .B1(n7271), .B2(n7270), .A(n10034), .ZN(n7283) );
  INV_X1 U8613 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7273) );
  NOR2_X1 U8614 ( .A1(n10035), .A2(n7273), .ZN(n7272) );
  AOI21_X1 U8615 ( .B1(n7273), .B2(n10035), .A(n7272), .ZN(n7276) );
  AOI21_X1 U8616 ( .B1(n7820), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7274), .ZN(
        n7275) );
  NOR2_X1 U8617 ( .A1(n7275), .A2(n7276), .ZN(n10031) );
  AOI211_X1 U8618 ( .C1(n7276), .C2(n7275), .A(n10031), .B(n10665), .ZN(n7282)
         );
  NAND2_X1 U8619 ( .A1(n10664), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n7279) );
  NOR2_X1 U8620 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7277), .ZN(n9157) );
  INV_X1 U8621 ( .A(n9157), .ZN(n7278) );
  OAI211_X1 U8622 ( .C1(n7280), .C2(n10691), .A(n7279), .B(n7278), .ZN(n7281)
         );
  AOI211_X1 U8623 ( .C1(n10677), .C2(n7283), .A(n7282), .B(n7281), .ZN(n7284)
         );
  INV_X1 U8624 ( .A(n7284), .ZN(P1_U3255) );
  INV_X1 U8625 ( .A(n7290), .ZN(n7285) );
  NAND2_X1 U8626 ( .A1(n7286), .A2(n7285), .ZN(n7287) );
  NAND2_X1 U8627 ( .A1(n7356), .A2(n7483), .ZN(n10835) );
  INV_X1 U8628 ( .A(n7483), .ZN(n7288) );
  NAND2_X1 U8629 ( .A1(n7288), .A2(n10844), .ZN(n10837) );
  AOI222_X1 U8630 ( .A1(n10014), .A2(n10843), .B1(n10013), .B2(n10842), .C1(
        n10920), .C2(n7289), .ZN(n7485) );
  NAND2_X1 U8631 ( .A1(n7291), .A2(n7290), .ZN(n7294) );
  NAND2_X1 U8632 ( .A1(n7292), .A2(n10777), .ZN(n7293) );
  NAND2_X1 U8633 ( .A1(n5666), .A2(n7295), .ZN(n7411) );
  OAI21_X1 U8634 ( .B1(n5666), .B2(n7295), .A(n7411), .ZN(n7486) );
  INV_X1 U8635 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7297) );
  OAI22_X1 U8636 ( .A1(n10942), .A2(n7297), .B1(n7296), .B2(n10937), .ZN(n7298) );
  AOI21_X1 U8637 ( .B1(n10317), .B2(n7483), .A(n7298), .ZN(n7302) );
  AOI21_X1 U8638 ( .B1(n7299), .B2(n7483), .A(n11043), .ZN(n7300) );
  AND2_X1 U8639 ( .A1(n7300), .A2(n10833), .ZN(n7482) );
  NAND2_X1 U8640 ( .A1(n7482), .A2(n10281), .ZN(n7301) );
  OAI211_X1 U8641 ( .C1(n7486), .C2(n10300), .A(n7302), .B(n7301), .ZN(n7303)
         );
  INV_X1 U8642 ( .A(n7303), .ZN(n7304) );
  OAI21_X1 U8643 ( .B1(n7485), .B2(n10296), .A(n7304), .ZN(P1_U3286) );
  NOR2_X1 U8644 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5991), .ZN(n7933) );
  INV_X1 U8645 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7305) );
  MUX2_X1 U8646 ( .A(n7305), .B(P2_REG1_REG_14__SCAN_IN), .S(n8693), .Z(n7309)
         );
  AOI21_X1 U8647 ( .B1(n7307), .B2(n11016), .A(n7306), .ZN(n7308) );
  NOR2_X1 U8648 ( .A1(n7308), .A2(n7309), .ZN(n8699) );
  AOI21_X1 U8649 ( .B1(n7309), .B2(n7308), .A(n8699), .ZN(n7310) );
  NOR2_X1 U8650 ( .A1(n10624), .A2(n7310), .ZN(n7311) );
  AOI211_X1 U8651 ( .C1(P2_ADDR_REG_14__SCAN_IN), .C2(n10647), .A(n7933), .B(
        n7311), .ZN(n7319) );
  INV_X1 U8652 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7312) );
  MUX2_X1 U8653 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n7312), .S(n8693), .Z(n7316)
         );
  OAI21_X1 U8654 ( .B1(n7314), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7313), .ZN(
        n7315) );
  NAND2_X1 U8655 ( .A1(n7316), .A2(n7315), .ZN(n8692) );
  OAI21_X1 U8656 ( .B1(n7316), .B2(n7315), .A(n8692), .ZN(n7317) );
  NAND2_X1 U8657 ( .A1(n10622), .A2(n7317), .ZN(n7318) );
  OAI211_X1 U8658 ( .C1(n10638), .C2(n8700), .A(n7319), .B(n7318), .ZN(
        P2_U3259) );
  INV_X1 U8659 ( .A(n8077), .ZN(n10948) );
  OAI211_X1 U8660 ( .C1(n7322), .C2(n7321), .A(n7320), .B(n10964), .ZN(n7326)
         );
  AND2_X1 U8661 ( .A1(P2_U3152), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8668) );
  AOI22_X1 U8662 ( .A1(n9014), .A2(n9017), .B1(n7323), .B2(n9016), .ZN(n7365)
         );
  INV_X1 U8663 ( .A(n10955), .ZN(n8552) );
  NOR2_X1 U8664 ( .A1(n7365), .A2(n8552), .ZN(n7324) );
  AOI211_X1 U8665 ( .C1(n6450), .C2(n7368), .A(n8668), .B(n7324), .ZN(n7325)
         );
  OAI211_X1 U8666 ( .C1(n10948), .C2(n6439), .A(n7326), .B(n7325), .ZN(
        P2_U3223) );
  OR2_X1 U8667 ( .A1(n7060), .A2(n7330), .ZN(n7333) );
  OR2_X1 U8668 ( .A1(n5030), .A2(n7331), .ZN(n7332) );
  OAI211_X1 U8669 ( .C1(n6895), .C2(n7334), .A(n7333), .B(n7332), .ZN(n7433)
         );
  NAND2_X1 U8670 ( .A1(n7433), .A2(n7802), .ZN(n7335) );
  OAI21_X1 U8671 ( .B1(n7428), .B2(n9187), .A(n7335), .ZN(n7336) );
  XNOR2_X1 U8672 ( .A(n7336), .B(n9185), .ZN(n7338) );
  AND2_X1 U8673 ( .A1(n7433), .A2(n9181), .ZN(n7337) );
  AOI21_X1 U8674 ( .B1(n10013), .B2(n9182), .A(n7337), .ZN(n7339) );
  NAND2_X1 U8675 ( .A1(n7338), .A2(n7339), .ZN(n7445) );
  INV_X1 U8676 ( .A(n7338), .ZN(n7341) );
  INV_X1 U8677 ( .A(n7339), .ZN(n7340) );
  NAND2_X1 U8678 ( .A1(n7341), .A2(n7340), .ZN(n7342) );
  NAND2_X1 U8679 ( .A1(n7445), .A2(n7342), .ZN(n7346) );
  INV_X1 U8680 ( .A(n7446), .ZN(n7345) );
  AOI21_X1 U8681 ( .B1(n7343), .B2(n7346), .A(n7345), .ZN(n7361) );
  OR2_X1 U8682 ( .A1(n5034), .A2(n7347), .ZN(n7354) );
  AND2_X1 U8683 ( .A1(n7349), .A2(n7348), .ZN(n7350) );
  OR2_X1 U8684 ( .A1(n7350), .A2(n7422), .ZN(n7451) );
  OR2_X1 U8685 ( .A1(n5032), .A2(n7451), .ZN(n7353) );
  NAND2_X1 U8686 ( .A1(n7753), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7352) );
  NAND2_X1 U8687 ( .A1(n7712), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n7351) );
  NAND4_X1 U8688 ( .A1(n7354), .A2(n7353), .A3(n7352), .A4(n7351), .ZN(n10841)
         );
  INV_X1 U8689 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7355) );
  NOR2_X1 U8690 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7355), .ZN(n10524) );
  NOR2_X1 U8691 ( .A1(n9314), .A2(n7356), .ZN(n7357) );
  AOI211_X1 U8692 ( .C1(n9300), .C2(n10841), .A(n10524), .B(n7357), .ZN(n7358)
         );
  OAI21_X1 U8693 ( .B1(n9315), .B2(n10856), .A(n7358), .ZN(n7359) );
  AOI21_X1 U8694 ( .B1(n7433), .B2(n9220), .A(n7359), .ZN(n7360) );
  OAI21_X1 U8695 ( .B1(n7361), .B2(n9309), .A(n7360), .ZN(P1_U3237) );
  INV_X1 U8696 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7362) );
  INV_X1 U8697 ( .A(n7981), .ZN(n7363) );
  OAI222_X1 U8698 ( .A1(n9146), .A2(n7362), .B1(n9147), .B2(n7363), .C1(n6223), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  INV_X1 U8699 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9743) );
  OAI222_X1 U8700 ( .A1(P1_U3084), .A2(n10229), .B1(n10461), .B2(n7363), .C1(
        n9743), .C2(n10454), .ZN(P1_U3334) );
  INV_X1 U8701 ( .A(n7373), .ZN(n8201) );
  XNOR2_X1 U8702 ( .A(n7364), .B(n8201), .ZN(n7366) );
  OAI21_X1 U8703 ( .B1(n7366), .B2(n8932), .A(n7365), .ZN(n10949) );
  AOI21_X1 U8704 ( .B1(n7386), .B2(n8077), .A(n11030), .ZN(n7367) );
  NAND2_X1 U8705 ( .A1(n7367), .A2(n7402), .ZN(n10947) );
  AND2_X1 U8706 ( .A1(n10818), .A2(n6223), .ZN(n9011) );
  INV_X1 U8707 ( .A(n9011), .ZN(n7623) );
  INV_X1 U8708 ( .A(n7368), .ZN(n7369) );
  OAI22_X1 U8709 ( .A1(n10818), .A2(n7370), .B1(n7369), .B2(n8987), .ZN(n7371)
         );
  AOI21_X1 U8710 ( .B1(n10767), .B2(n8077), .A(n7371), .ZN(n7372) );
  OAI21_X1 U8711 ( .B1(n10947), .B2(n7623), .A(n7372), .ZN(n7378) );
  NOR2_X1 U8712 ( .A1(n7374), .A2(n7373), .ZN(n10946) );
  INV_X1 U8713 ( .A(n7375), .ZN(n7376) );
  NOR3_X1 U8714 ( .A1(n10946), .A2(n7376), .A3(n9008), .ZN(n7377) );
  AOI211_X1 U8715 ( .C1(n10818), .C2(n10949), .A(n7378), .B(n7377), .ZN(n7379)
         );
  INV_X1 U8716 ( .A(n7379), .ZN(P2_U3288) );
  XNOR2_X1 U8717 ( .A(n7380), .B(n8074), .ZN(n7381) );
  NAND2_X1 U8718 ( .A1(n7381), .A2(n10808), .ZN(n7383) );
  AOI22_X1 U8719 ( .A1(n10883), .A2(n9016), .B1(n9014), .B2(n8664), .ZN(n7382)
         );
  NAND2_X1 U8720 ( .A1(n7383), .A2(n7382), .ZN(n10899) );
  INV_X1 U8721 ( .A(n10899), .ZN(n7392) );
  OAI21_X1 U8722 ( .B1(n7385), .B2(n5145), .A(n7384), .ZN(n10901) );
  OAI21_X1 U8723 ( .B1(n9027), .B2(n5151), .A(n7386), .ZN(n10898) );
  AOI22_X1 U8724 ( .A1(n10821), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7387), .B2(
        n10813), .ZN(n7389) );
  NAND2_X1 U8725 ( .A1(n10767), .A2(n10895), .ZN(n7388) );
  OAI211_X1 U8726 ( .C1(n10898), .C2(n8788), .A(n7389), .B(n7388), .ZN(n7390)
         );
  AOI21_X1 U8727 ( .B1(n10901), .B2(n9024), .A(n7390), .ZN(n7391) );
  OAI21_X1 U8728 ( .B1(n10821), .B2(n7392), .A(n7391), .ZN(P2_U3289) );
  OAI211_X1 U8729 ( .C1(n7394), .C2(n8203), .A(n7393), .B(n10808), .ZN(n7398)
         );
  OR2_X1 U8730 ( .A1(n7562), .A2(n10794), .ZN(n7396) );
  OR2_X1 U8731 ( .A1(n8076), .A2(n10792), .ZN(n7395) );
  NAND2_X1 U8732 ( .A1(n7396), .A2(n7395), .ZN(n10956) );
  INV_X1 U8733 ( .A(n10956), .ZN(n7397) );
  NAND2_X1 U8734 ( .A1(n7398), .A2(n7397), .ZN(n10972) );
  INV_X1 U8735 ( .A(n10972), .ZN(n7409) );
  OAI21_X1 U8736 ( .B1(n7401), .B2(n7400), .A(n7399), .ZN(n10974) );
  INV_X1 U8737 ( .A(n10962), .ZN(n10970) );
  INV_X1 U8738 ( .A(n7512), .ZN(n7403) );
  OAI21_X1 U8739 ( .B1(n10970), .B2(n5277), .A(n7403), .ZN(n10971) );
  OAI22_X1 U8740 ( .A1(n10818), .A2(n7404), .B1(n10969), .B2(n8987), .ZN(n7405) );
  AOI21_X1 U8741 ( .B1(n10962), .B2(n10767), .A(n7405), .ZN(n7406) );
  OAI21_X1 U8742 ( .B1(n10971), .B2(n8788), .A(n7406), .ZN(n7407) );
  AOI21_X1 U8743 ( .B1(n10974), .B2(n9024), .A(n7407), .ZN(n7408) );
  OAI21_X1 U8744 ( .B1(n10821), .B2(n7409), .A(n7408), .ZN(P2_U3287) );
  NAND2_X1 U8745 ( .A1(n10844), .A2(n7483), .ZN(n7410) );
  NAND2_X1 U8746 ( .A1(n7428), .A2(n7433), .ZN(n9493) );
  INV_X1 U8747 ( .A(n7433), .ZN(n10855) );
  NAND2_X1 U8748 ( .A1(n10855), .A2(n10013), .ZN(n9349) );
  OR2_X1 U8749 ( .A1(n10830), .A2(n10838), .ZN(n10831) );
  NAND2_X1 U8750 ( .A1(n7428), .A2(n10855), .ZN(n7527) );
  NAND2_X1 U8751 ( .A1(n10831), .A2(n7527), .ZN(n7415) );
  INV_X2 U8752 ( .A(n7060), .ZN(n7983) );
  INV_X2 U8753 ( .A(n6895), .ZN(n7982) );
  AOI22_X1 U8754 ( .A1(n7983), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7982), .B2(
        n7412), .ZN(n7414) );
  NAND2_X1 U8755 ( .A1(n10876), .A2(n10841), .ZN(n9496) );
  INV_X1 U8756 ( .A(n10841), .ZN(n10916) );
  NAND2_X1 U8757 ( .A1(n10916), .A2(n7450), .ZN(n10911) );
  NAND2_X1 U8758 ( .A1(n9496), .A2(n10911), .ZN(n7519) );
  XNOR2_X1 U8759 ( .A(n7415), .B(n7519), .ZN(n10878) );
  NAND2_X1 U8760 ( .A1(n10878), .A2(n10840), .ZN(n7432) );
  NAND2_X1 U8761 ( .A1(n9493), .A2(n10835), .ZN(n9401) );
  INV_X1 U8762 ( .A(n7519), .ZN(n9435) );
  INV_X1 U8763 ( .A(n10837), .ZN(n9494) );
  NAND2_X1 U8764 ( .A1(n9493), .A2(n9494), .ZN(n9399) );
  AND2_X1 U8765 ( .A1(n9399), .A2(n9349), .ZN(n7417) );
  AND2_X1 U8766 ( .A1(n9435), .A2(n7417), .ZN(n7416) );
  NAND2_X1 U8767 ( .A1(n7418), .A2(n7417), .ZN(n7419) );
  NAND2_X1 U8768 ( .A1(n7419), .A2(n7519), .ZN(n7420) );
  NAND2_X1 U8769 ( .A1(n10912), .A2(n7420), .ZN(n7430) );
  NAND2_X1 U8770 ( .A1(n8412), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7427) );
  NAND2_X1 U8771 ( .A1(n7753), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7426) );
  OR2_X1 U8772 ( .A1(n5034), .A2(n10927), .ZN(n7425) );
  OR2_X1 U8773 ( .A1(n7422), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7423) );
  NAND2_X1 U8774 ( .A1(n7536), .A2(n7423), .ZN(n10938) );
  OR2_X1 U8775 ( .A1(n5032), .A2(n10938), .ZN(n7424) );
  OAI22_X1 U8776 ( .A1(n7602), .A2(n10917), .B1(n7428), .B2(n10915), .ZN(n7429) );
  AOI21_X1 U8777 ( .B1(n7430), .B2(n10920), .A(n7429), .ZN(n7431) );
  AND2_X1 U8778 ( .A1(n7432), .A2(n7431), .ZN(n10880) );
  NAND2_X1 U8779 ( .A1(n10834), .A2(n7450), .ZN(n7434) );
  NAND2_X1 U8780 ( .A1(n7434), .A2(n10711), .ZN(n7435) );
  OR2_X1 U8781 ( .A1(n7435), .A2(n10910), .ZN(n10875) );
  INV_X1 U8782 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7436) );
  OAI22_X1 U8783 ( .A1(n10942), .A2(n7436), .B1(n7451), .B2(n10937), .ZN(n7437) );
  AOI21_X1 U8784 ( .B1(n10317), .B2(n7450), .A(n7437), .ZN(n7438) );
  OAI21_X1 U8785 ( .B1(n10875), .B2(n10313), .A(n7438), .ZN(n7439) );
  AOI21_X1 U8786 ( .B1(n10878), .B2(n10933), .A(n7439), .ZN(n7440) );
  OAI21_X1 U8787 ( .B1(n10880), .B2(n10296), .A(n7440), .ZN(P1_U3284) );
  NAND2_X1 U8788 ( .A1(n10841), .A2(n9181), .ZN(n7441) );
  OAI21_X1 U8789 ( .B1(n10876), .B2(n8382), .A(n7441), .ZN(n7442) );
  XNOR2_X1 U8790 ( .A(n7442), .B(n9185), .ZN(n7572) );
  OR2_X1 U8791 ( .A1(n10876), .A2(n9187), .ZN(n7444) );
  NAND2_X1 U8792 ( .A1(n10841), .A2(n9182), .ZN(n7443) );
  NAND2_X1 U8793 ( .A1(n7444), .A2(n7443), .ZN(n7570) );
  XNOR2_X1 U8794 ( .A(n7572), .B(n7570), .ZN(n7448) );
  OAI21_X1 U8795 ( .B1(n7448), .B2(n7447), .A(n7574), .ZN(n7457) );
  AOI21_X1 U8796 ( .B1(n9289), .B2(n10013), .A(n7449), .ZN(n7455) );
  NAND2_X1 U8797 ( .A1(n7450), .A2(n9292), .ZN(n7454) );
  OR2_X1 U8798 ( .A1(n9315), .A2(n7451), .ZN(n7453) );
  NAND2_X1 U8799 ( .A1(n10012), .A2(n9300), .ZN(n7452) );
  NAND4_X1 U8800 ( .A1(n7455), .A2(n7454), .A3(n7453), .A4(n7452), .ZN(n7456)
         );
  AOI21_X1 U8801 ( .B1(n7457), .B2(n9295), .A(n7456), .ZN(n7458) );
  INV_X1 U8802 ( .A(n7458), .ZN(P1_U3211) );
  INV_X1 U8803 ( .A(n7459), .ZN(n7460) );
  NAND2_X1 U8804 ( .A1(n10818), .A2(n7460), .ZN(n8992) );
  INV_X1 U8805 ( .A(n8992), .ZN(n10771) );
  OAI21_X1 U8806 ( .B1(n7462), .B2(n8049), .A(n7461), .ZN(n10748) );
  NAND2_X1 U8807 ( .A1(n7464), .A2(n7463), .ZN(n7465) );
  NAND2_X1 U8808 ( .A1(n7466), .A2(n7465), .ZN(n10745) );
  INV_X1 U8809 ( .A(n10745), .ZN(n7467) );
  AOI22_X1 U8810 ( .A1(n10764), .A2(n7467), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n10813), .ZN(n7468) );
  OAI21_X1 U8811 ( .B1(n10744), .B2(n8963), .A(n7468), .ZN(n7476) );
  INV_X1 U8812 ( .A(n8985), .ZN(n10762) );
  NAND2_X1 U8813 ( .A1(n10748), .A2(n10762), .ZN(n7474) );
  AOI22_X1 U8814 ( .A1(n6592), .A2(n9016), .B1(n9014), .B2(n7469), .ZN(n7473)
         );
  OAI21_X1 U8815 ( .B1(n8193), .B2(n8044), .A(n7470), .ZN(n7471) );
  NAND2_X1 U8816 ( .A1(n7471), .A2(n10808), .ZN(n7472) );
  NAND3_X1 U8817 ( .A1(n7474), .A2(n7473), .A3(n7472), .ZN(n10746) );
  MUX2_X1 U8818 ( .A(n10746), .B(P2_REG2_REG_2__SCAN_IN), .S(n10821), .Z(n7475) );
  AOI211_X1 U8819 ( .C1(n10771), .C2(n10748), .A(n7476), .B(n7475), .ZN(n7477)
         );
  INV_X1 U8820 ( .A(n7477), .ZN(P2_U3294) );
  INV_X1 U8821 ( .A(n7986), .ZN(n7491) );
  OAI222_X1 U8822 ( .A1(n9147), .A2(n7491), .B1(P2_U3152), .B2(n5028), .C1(
        n7478), .C2(n9146), .ZN(P2_U3338) );
  AOI21_X1 U8823 ( .B1(n11048), .B2(n7483), .A(n7482), .ZN(n7484) );
  OAI211_X1 U8824 ( .C1(n10415), .C2(n7486), .A(n7485), .B(n7484), .ZN(n7488)
         );
  NAND2_X1 U8825 ( .A1(n7488), .A2(n11050), .ZN(n7487) );
  OAI21_X1 U8826 ( .B1(n11050), .B2(n7067), .A(n7487), .ZN(P1_U3528) );
  INV_X1 U8827 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7490) );
  NAND2_X1 U8828 ( .A1(n7488), .A2(n11054), .ZN(n7489) );
  OAI21_X1 U8829 ( .B1(n11054), .B2(n7490), .A(n7489), .ZN(P1_U3469) );
  INV_X1 U8830 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n9612) );
  OAI222_X1 U8831 ( .A1(n7492), .A2(P1_U3084), .B1(n10461), .B2(n7491), .C1(
        n9612), .C2(n10454), .ZN(P1_U3333) );
  XNOR2_X1 U8832 ( .A(n7494), .B(n7493), .ZN(n7500) );
  NOR2_X1 U8833 ( .A1(n10886), .A2(n7507), .ZN(n7496) );
  OAI22_X1 U8834 ( .A1(n8606), .A2(n7685), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9687), .ZN(n7495) );
  AOI211_X1 U8835 ( .C1(n6450), .C2(n7497), .A(n7496), .B(n7495), .ZN(n7499)
         );
  NAND2_X1 U8836 ( .A1(n7516), .A2(n10963), .ZN(n7498) );
  OAI211_X1 U8837 ( .C1(n7500), .C2(n10890), .A(n7499), .B(n7498), .ZN(
        P2_U3219) );
  OAI222_X1 U8838 ( .A1(n9147), .A2(n7989), .B1(n8034), .B2(P2_U3152), .C1(
        n7501), .C2(n9146), .ZN(P2_U3337) );
  INV_X1 U8839 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7990) );
  OAI222_X1 U8840 ( .A1(n7502), .A2(P1_U3084), .B1(n10461), .B2(n7989), .C1(
        n7990), .C2(n10454), .ZN(P1_U3332) );
  NAND2_X1 U8841 ( .A1(n7503), .A2(n8192), .ZN(n7504) );
  OAI21_X1 U8842 ( .B1(n8192), .B2(n7506), .A(n7505), .ZN(n7509) );
  OAI22_X1 U8843 ( .A1(n7685), .A2(n10794), .B1(n7507), .B2(n10792), .ZN(n7508) );
  AOI21_X1 U8844 ( .B1(n7509), .B2(n10808), .A(n7508), .ZN(n7510) );
  OAI21_X1 U8845 ( .B1(n10978), .B2(n8985), .A(n7510), .ZN(n10981) );
  NAND2_X1 U8846 ( .A1(n10981), .A2(n10818), .ZN(n7518) );
  OAI22_X1 U8847 ( .A1(n10818), .A2(n6781), .B1(n7511), .B2(n8987), .ZN(n7515)
         );
  NOR2_X1 U8848 ( .A1(n7512), .A2(n10979), .ZN(n7513) );
  OR2_X1 U8849 ( .A1(n7616), .A2(n7513), .ZN(n10980) );
  NOR2_X1 U8850 ( .A1(n10980), .A2(n8788), .ZN(n7514) );
  AOI211_X1 U8851 ( .C1(n10767), .C2(n7516), .A(n7515), .B(n7514), .ZN(n7517)
         );
  OAI211_X1 U8852 ( .C1(n10978), .C2(n8992), .A(n7518), .B(n7517), .ZN(
        P2_U3286) );
  INV_X1 U8853 ( .A(n10830), .ZN(n7521) );
  NAND2_X1 U8854 ( .A1(n10876), .A2(n10916), .ZN(n7526) );
  INV_X1 U8855 ( .A(n7526), .ZN(n7520) );
  NOR2_X1 U8856 ( .A1(n7520), .A2(n7519), .ZN(n7529) );
  NAND2_X1 U8857 ( .A1(n7522), .A2(n9390), .ZN(n7525) );
  AOI22_X1 U8858 ( .A1(n7983), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7982), .B2(
        n7523), .ZN(n7524) );
  NAND2_X1 U8859 ( .A1(n7525), .A2(n7524), .ZN(n7578) );
  OR2_X1 U8860 ( .A1(n7578), .A2(n7602), .ZN(n9501) );
  NAND2_X1 U8861 ( .A1(n7578), .A2(n7602), .ZN(n9500) );
  INV_X1 U8862 ( .A(n10913), .ZN(n9504) );
  AND2_X1 U8863 ( .A1(n7527), .A2(n7526), .ZN(n7528) );
  OR2_X1 U8864 ( .A1(n7529), .A2(n7528), .ZN(n10904) );
  AND2_X1 U8865 ( .A1(n9504), .A2(n10904), .ZN(n7530) );
  NAND2_X1 U8866 ( .A1(n10905), .A2(n7530), .ZN(n10908) );
  NAND2_X1 U8867 ( .A1(n7578), .A2(n10012), .ZN(n7531) );
  NAND2_X1 U8868 ( .A1(n7532), .A2(n9390), .ZN(n7534) );
  AOI22_X1 U8869 ( .A1(n7983), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7982), .B2(
        n10537), .ZN(n7533) );
  OR2_X1 U8870 ( .A1(n5034), .A2(n7556), .ZN(n7541) );
  NAND2_X1 U8871 ( .A1(n7536), .A2(n7535), .ZN(n7537) );
  NAND2_X1 U8872 ( .A1(n7546), .A2(n7537), .ZN(n7668) );
  OR2_X1 U8873 ( .A1(n5032), .A2(n7668), .ZN(n7540) );
  NAND2_X1 U8874 ( .A1(n5035), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7539) );
  NAND2_X1 U8875 ( .A1(n7753), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n7538) );
  NAND4_X1 U8876 ( .A1(n7541), .A2(n7540), .A3(n7539), .A4(n7538), .ZN(n10011)
         );
  INV_X1 U8877 ( .A(n10011), .ZN(n10918) );
  OR2_X1 U8878 ( .A1(n7773), .A2(n10918), .ZN(n9325) );
  NAND2_X1 U8879 ( .A1(n7773), .A2(n10918), .ZN(n9506) );
  XOR2_X1 U8880 ( .A(n7772), .B(n9503), .Z(n7677) );
  INV_X1 U8881 ( .A(n10911), .ZN(n7542) );
  NOR2_X1 U8882 ( .A1(n9504), .A2(n7542), .ZN(n7543) );
  INV_X1 U8883 ( .A(n9501), .ZN(n9326) );
  NAND2_X1 U8884 ( .A1(n7544), .A2(n9503), .ZN(n7743) );
  OAI21_X1 U8885 ( .B1(n9503), .B2(n7544), .A(n7743), .ZN(n7552) );
  NAND2_X1 U8886 ( .A1(n8412), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7551) );
  NAND2_X1 U8887 ( .A1(n7753), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7550) );
  OR2_X1 U8888 ( .A1(n5034), .A2(n7545), .ZN(n7549) );
  NAND2_X1 U8889 ( .A1(n7546), .A2(n7721), .ZN(n7547) );
  NAND2_X1 U8890 ( .A1(n7715), .A2(n7547), .ZN(n7790) );
  OR2_X1 U8891 ( .A1(n5032), .A2(n7790), .ZN(n7548) );
  AOI222_X1 U8892 ( .A1(n10920), .A2(n7552), .B1(n10010), .B2(n10842), .C1(
        n10012), .C2(n10843), .ZN(n7672) );
  INV_X1 U8893 ( .A(n7789), .ZN(n7553) );
  AOI21_X1 U8894 ( .B1(n7773), .B2(n10909), .A(n7553), .ZN(n7675) );
  AOI22_X1 U8895 ( .A1(n7675), .A2(n10711), .B1(n11048), .B2(n7773), .ZN(n7554) );
  OAI211_X1 U8896 ( .C1(n7677), .C2(n10415), .A(n7672), .B(n7554), .ZN(n7557)
         );
  NAND2_X1 U8897 ( .A1(n7557), .A2(n11050), .ZN(n7555) );
  OAI21_X1 U8898 ( .B1(n11050), .B2(n7556), .A(n7555), .ZN(P1_U3532) );
  INV_X1 U8899 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7559) );
  NAND2_X1 U8900 ( .A1(n7557), .A2(n11054), .ZN(n7558) );
  OAI21_X1 U8901 ( .B1(n11054), .B2(n7559), .A(n7558), .ZN(P1_U3481) );
  XNOR2_X1 U8902 ( .A(n7561), .B(n7560), .ZN(n7569) );
  OR2_X1 U8903 ( .A1(n7915), .A2(n10794), .ZN(n7564) );
  OR2_X1 U8904 ( .A1(n7562), .A2(n10792), .ZN(n7563) );
  AND2_X1 U8905 ( .A1(n7564), .A2(n7563), .ZN(n7610) );
  NOR2_X1 U8906 ( .A1(n7610), .A2(n8552), .ZN(n7565) );
  AOI211_X1 U8907 ( .C1(n6450), .C2(n7617), .A(n7566), .B(n7565), .ZN(n7568)
         );
  NAND2_X1 U8908 ( .A1(n7621), .A2(n10963), .ZN(n7567) );
  OAI211_X1 U8909 ( .C1(n7569), .C2(n10890), .A(n7568), .B(n7567), .ZN(
        P2_U3238) );
  INV_X1 U8910 ( .A(n7570), .ZN(n7571) );
  NAND2_X1 U8911 ( .A1(n7572), .A2(n7571), .ZN(n7573) );
  NAND2_X1 U8912 ( .A1(n7574), .A2(n7573), .ZN(n7690) );
  INV_X1 U8913 ( .A(n7690), .ZN(n7577) );
  NAND2_X1 U8914 ( .A1(n7578), .A2(n9181), .ZN(n7576) );
  NAND2_X1 U8915 ( .A1(n10012), .A2(n9182), .ZN(n7575) );
  NAND2_X1 U8916 ( .A1(n7576), .A2(n7575), .ZN(n7693) );
  NAND2_X1 U8917 ( .A1(n7577), .A2(n7693), .ZN(n7584) );
  NAND2_X1 U8918 ( .A1(n7578), .A2(n7802), .ZN(n7580) );
  NAND2_X1 U8919 ( .A1(n10012), .A2(n9181), .ZN(n7579) );
  NAND2_X1 U8920 ( .A1(n7580), .A2(n7579), .ZN(n7581) );
  XNOR2_X1 U8921 ( .A(n7581), .B(n8418), .ZN(n7692) );
  INV_X1 U8922 ( .A(n7692), .ZN(n7695) );
  NAND2_X1 U8923 ( .A1(n7584), .A2(n7695), .ZN(n7594) );
  INV_X1 U8924 ( .A(n7693), .ZN(n7582) );
  NAND2_X1 U8925 ( .A1(n7690), .A2(n7582), .ZN(n7593) );
  INV_X1 U8926 ( .A(n7593), .ZN(n7583) );
  NOR2_X1 U8927 ( .A1(n7594), .A2(n7583), .ZN(n7586) );
  AOI21_X1 U8928 ( .B1(n7584), .B2(n7593), .A(n7695), .ZN(n7585) );
  OAI21_X1 U8929 ( .B1(n7586), .B2(n7585), .A(n9295), .ZN(n7592) );
  NOR2_X1 U8930 ( .A1(n9315), .A2(n10938), .ZN(n7590) );
  NAND2_X1 U8931 ( .A1(n9300), .A2(n10011), .ZN(n7588) );
  OAI211_X1 U8932 ( .C1(n9314), .C2(n10916), .A(n7588), .B(n7587), .ZN(n7589)
         );
  NOR2_X1 U8933 ( .A1(n7590), .A2(n7589), .ZN(n7591) );
  OAI211_X1 U8934 ( .C1(n10936), .C2(n9321), .A(n7592), .B(n7591), .ZN(
        P1_U3219) );
  NAND2_X1 U8935 ( .A1(n7594), .A2(n7593), .ZN(n7601) );
  NAND2_X1 U8936 ( .A1(n7773), .A2(n7802), .ZN(n7596) );
  NAND2_X1 U8937 ( .A1(n10011), .A2(n9181), .ZN(n7595) );
  NAND2_X1 U8938 ( .A1(n7596), .A2(n7595), .ZN(n7597) );
  XNOR2_X1 U8939 ( .A(n7597), .B(n8418), .ZN(n7691) );
  NAND2_X1 U8940 ( .A1(n7773), .A2(n9181), .ZN(n7599) );
  NAND2_X1 U8941 ( .A1(n10011), .A2(n9182), .ZN(n7598) );
  NAND2_X1 U8942 ( .A1(n7599), .A2(n7598), .ZN(n7694) );
  XNOR2_X1 U8943 ( .A(n7691), .B(n7694), .ZN(n7600) );
  XNOR2_X1 U8944 ( .A(n7601), .B(n7600), .ZN(n7607) );
  AND2_X1 U8945 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n10536) );
  NOR2_X1 U8946 ( .A1(n9314), .A2(n7602), .ZN(n7603) );
  AOI211_X1 U8947 ( .C1(n9300), .C2(n10010), .A(n10536), .B(n7603), .ZN(n7604)
         );
  OAI21_X1 U8948 ( .B1(n9315), .B2(n7668), .A(n7604), .ZN(n7605) );
  AOI21_X1 U8949 ( .B1(n7773), .B2(n9292), .A(n7605), .ZN(n7606) );
  OAI21_X1 U8950 ( .B1(n7607), .B2(n9309), .A(n7606), .ZN(P1_U3229) );
  XNOR2_X1 U8951 ( .A(n7608), .B(n8204), .ZN(n7609) );
  NAND2_X1 U8952 ( .A1(n7609), .A2(n10808), .ZN(n7611) );
  NAND2_X1 U8953 ( .A1(n7611), .A2(n7610), .ZN(n10989) );
  INV_X1 U8954 ( .A(n10989), .ZN(n7626) );
  OAI21_X1 U8955 ( .B1(n7614), .B2(n7613), .A(n7612), .ZN(n7615) );
  INV_X1 U8956 ( .A(n7615), .ZN(n10991) );
  OAI211_X1 U8957 ( .C1(n7616), .C2(n10988), .A(n10865), .B(n7733), .ZN(n10987) );
  INV_X1 U8958 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7619) );
  INV_X1 U8959 ( .A(n7617), .ZN(n7618) );
  OAI22_X1 U8960 ( .A1(n10818), .A2(n7619), .B1(n7618), .B2(n8987), .ZN(n7620)
         );
  AOI21_X1 U8961 ( .B1(n7621), .B2(n10767), .A(n7620), .ZN(n7622) );
  OAI21_X1 U8962 ( .B1(n10987), .B2(n7623), .A(n7622), .ZN(n7624) );
  AOI21_X1 U8963 ( .B1(n10991), .B2(n9024), .A(n7624), .ZN(n7625) );
  OAI21_X1 U8964 ( .B1(n10821), .B2(n7626), .A(n7625), .ZN(P2_U3285) );
  NOR2_X1 U8965 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7663) );
  NOR2_X1 U8966 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7661) );
  NOR2_X1 U8967 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7659) );
  NOR2_X1 U8968 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7657) );
  NOR2_X1 U8969 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7655) );
  NOR2_X1 U8970 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7653) );
  NAND2_X1 U8971 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7651) );
  XOR2_X1 U8972 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10494) );
  NAND2_X1 U8973 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7649) );
  XOR2_X1 U8974 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10492) );
  NOR2_X1 U8975 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7633) );
  XNOR2_X1 U8976 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10483) );
  NAND2_X1 U8977 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7631) );
  XOR2_X1 U8978 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10481) );
  NAND2_X1 U8979 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7629) );
  XOR2_X1 U8980 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10479) );
  AOI21_X1 U8981 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10474) );
  INV_X1 U8982 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7627) );
  NAND3_X1 U8983 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10476) );
  OAI21_X1 U8984 ( .B1(n10474), .B2(n7627), .A(n10476), .ZN(n10478) );
  NAND2_X1 U8985 ( .A1(n10479), .A2(n10478), .ZN(n7628) );
  NAND2_X1 U8986 ( .A1(n7629), .A2(n7628), .ZN(n10480) );
  NAND2_X1 U8987 ( .A1(n10481), .A2(n10480), .ZN(n7630) );
  NAND2_X1 U8988 ( .A1(n7631), .A2(n7630), .ZN(n10482) );
  NOR2_X1 U8989 ( .A1(n10483), .A2(n10482), .ZN(n7632) );
  NOR2_X1 U8990 ( .A1(n7633), .A2(n7632), .ZN(n7634) );
  NOR2_X1 U8991 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7634), .ZN(n10485) );
  AND2_X1 U8992 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7634), .ZN(n10484) );
  NAND2_X1 U8993 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7636), .ZN(n7638) );
  XOR2_X1 U8994 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7636), .Z(n10487) );
  NAND2_X1 U8995 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10487), .ZN(n7637) );
  NAND2_X1 U8996 ( .A1(n7638), .A2(n7637), .ZN(n7639) );
  NAND2_X1 U8997 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7639), .ZN(n7641) );
  XOR2_X1 U8998 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7639), .Z(n10488) );
  NAND2_X1 U8999 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10488), .ZN(n7640) );
  NAND2_X1 U9000 ( .A1(n7641), .A2(n7640), .ZN(n7642) );
  NAND2_X1 U9001 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7642), .ZN(n7644) );
  XOR2_X1 U9002 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7642), .Z(n10489) );
  NAND2_X1 U9003 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10489), .ZN(n7643) );
  NAND2_X1 U9004 ( .A1(n7644), .A2(n7643), .ZN(n7645) );
  NAND2_X1 U9005 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7645), .ZN(n7647) );
  XOR2_X1 U9006 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7645), .Z(n10490) );
  NAND2_X1 U9007 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10490), .ZN(n7646) );
  NAND2_X1 U9008 ( .A1(n7647), .A2(n7646), .ZN(n10491) );
  NAND2_X1 U9009 ( .A1(n10492), .A2(n10491), .ZN(n7648) );
  NAND2_X1 U9010 ( .A1(n7649), .A2(n7648), .ZN(n10493) );
  NAND2_X1 U9011 ( .A1(n10494), .A2(n10493), .ZN(n7650) );
  NAND2_X1 U9012 ( .A1(n7651), .A2(n7650), .ZN(n10496) );
  XNOR2_X1 U9013 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10495) );
  XNOR2_X1 U9014 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10497) );
  XNOR2_X1 U9015 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10499) );
  NOR2_X1 U9016 ( .A1(n10500), .A2(n10499), .ZN(n7656) );
  NOR2_X1 U9017 ( .A1(n7657), .A2(n7656), .ZN(n10502) );
  XNOR2_X1 U9018 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10501) );
  NOR2_X1 U9019 ( .A1(n10502), .A2(n10501), .ZN(n7658) );
  NOR2_X1 U9020 ( .A1(n7659), .A2(n7658), .ZN(n10504) );
  XNOR2_X1 U9021 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10503) );
  NOR2_X1 U9022 ( .A1(n10504), .A2(n10503), .ZN(n7660) );
  NOR2_X1 U9023 ( .A1(n7661), .A2(n7660), .ZN(n10506) );
  XNOR2_X1 U9024 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10505) );
  NOR2_X1 U9025 ( .A1(n10506), .A2(n10505), .ZN(n7662) );
  NOR2_X1 U9026 ( .A1(n7663), .A2(n7662), .ZN(n7664) );
  AND2_X1 U9027 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7664), .ZN(n10507) );
  NOR2_X1 U9028 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10507), .ZN(n7665) );
  NOR2_X1 U9029 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n7664), .ZN(n10508) );
  NOR2_X1 U9030 ( .A1(n7665), .A2(n10508), .ZN(n7667) );
  XNOR2_X1 U9031 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7666) );
  XNOR2_X1 U9032 ( .A(n7667), .B(n7666), .ZN(ADD_1071_U4) );
  INV_X1 U9033 ( .A(n7773), .ZN(n7671) );
  INV_X1 U9034 ( .A(n7668), .ZN(n7669) );
  AOI22_X1 U9035 ( .A1(n10296), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7669), .B2(
        n10724), .ZN(n7670) );
  OAI21_X1 U9036 ( .B1(n7671), .B2(n10935), .A(n7670), .ZN(n7674) );
  NOR2_X1 U9037 ( .A1(n7672), .A2(n10296), .ZN(n7673) );
  AOI211_X1 U9038 ( .C1(n7675), .C2(n10932), .A(n7674), .B(n7673), .ZN(n7676)
         );
  OAI21_X1 U9039 ( .B1(n10300), .B2(n7677), .A(n7676), .ZN(P1_U3282) );
  INV_X1 U9040 ( .A(n7961), .ZN(n7679) );
  INV_X1 U9041 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7962) );
  OAI222_X1 U9042 ( .A1(P1_U3084), .A2(n6889), .B1(n10461), .B2(n7679), .C1(
        n7962), .C2(n10454), .ZN(P1_U3331) );
  OAI222_X1 U9043 ( .A1(n9146), .A2(n7680), .B1(n9147), .B2(n7679), .C1(
        P2_U3152), .C2(n7678), .ZN(P2_U3336) );
  XNOR2_X1 U9044 ( .A(n7681), .B(n7682), .ZN(n7688) );
  NAND2_X1 U9045 ( .A1(n6450), .A2(n7736), .ZN(n7684) );
  AOI22_X1 U9046 ( .A1(n10884), .A2(n8660), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n7683) );
  OAI211_X1 U9047 ( .C1(n7685), .C2(n10886), .A(n7684), .B(n7683), .ZN(n7686)
         );
  AOI21_X1 U9048 ( .B1(n7737), .B2(n10963), .A(n7686), .ZN(n7687) );
  OAI21_X1 U9049 ( .B1(n7688), .B2(n10890), .A(n7687), .ZN(P2_U3226) );
  AOI22_X1 U9050 ( .A1(n7691), .A2(n7694), .B1(n7693), .B2(n7692), .ZN(n7689)
         );
  INV_X1 U9051 ( .A(n7691), .ZN(n7698) );
  OAI21_X1 U9052 ( .B1(n7692), .B2(n7693), .A(n7694), .ZN(n7697) );
  NOR2_X1 U9053 ( .A1(n7694), .A2(n7693), .ZN(n7696) );
  AOI22_X1 U9054 ( .A1(n7698), .A2(n7697), .B1(n7696), .B2(n7695), .ZN(n7699)
         );
  NAND2_X1 U9055 ( .A1(n7700), .A2(n9390), .ZN(n7702) );
  AOI22_X1 U9056 ( .A1(n7983), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7982), .B2(
        n10550), .ZN(n7701) );
  NAND2_X1 U9057 ( .A1(n10412), .A2(n7802), .ZN(n7704) );
  NAND2_X1 U9058 ( .A1(n10010), .A2(n9181), .ZN(n7703) );
  NAND2_X1 U9059 ( .A1(n7704), .A2(n7703), .ZN(n7705) );
  XNOR2_X1 U9060 ( .A(n7705), .B(n9185), .ZN(n7707) );
  NOR2_X1 U9061 ( .A1(n7853), .A2(n8396), .ZN(n7706) );
  AOI21_X1 U9062 ( .B1(n10412), .B2(n9181), .A(n7706), .ZN(n7709) );
  OR2_X1 U9063 ( .A1(n7708), .A2(n7707), .ZN(n7710) );
  AOI21_X1 U9064 ( .B1(n7710), .B2(n7807), .A(n7709), .ZN(n7711) );
  AOI21_X1 U9065 ( .B1(n5101), .B2(n7807), .A(n7711), .ZN(n7726) );
  NAND2_X1 U9066 ( .A1(n5035), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U9067 ( .A1(n7753), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n7719) );
  OR2_X1 U9068 ( .A1(n5034), .A2(n7713), .ZN(n7718) );
  AND2_X1 U9069 ( .A1(n7715), .A2(n7714), .ZN(n7716) );
  OR2_X1 U9070 ( .A1(n7716), .A2(n7755), .ZN(n7811) );
  OR2_X1 U9071 ( .A1(n5032), .A2(n7811), .ZN(n7717) );
  NOR2_X1 U9072 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7721), .ZN(n10549) );
  NOR2_X1 U9073 ( .A1(n9314), .A2(n10918), .ZN(n7722) );
  AOI211_X1 U9074 ( .C1(n9300), .C2(n10009), .A(n10549), .B(n7722), .ZN(n7723)
         );
  OAI21_X1 U9075 ( .B1(n9315), .B2(n7790), .A(n7723), .ZN(n7724) );
  AOI21_X1 U9076 ( .B1(n10412), .B2(n9220), .A(n7724), .ZN(n7725) );
  OAI21_X1 U9077 ( .B1(n7726), .B2(n9309), .A(n7725), .ZN(P1_U3215) );
  XNOR2_X1 U9078 ( .A(n7727), .B(n8092), .ZN(n7728) );
  NAND2_X1 U9079 ( .A1(n7728), .A2(n10808), .ZN(n7730) );
  AOI22_X1 U9080 ( .A1(n8662), .A2(n9014), .B1(n9016), .B2(n8660), .ZN(n7729)
         );
  NAND2_X1 U9081 ( .A1(n7730), .A2(n7729), .ZN(n11002) );
  INV_X1 U9082 ( .A(n11002), .ZN(n7742) );
  OAI21_X1 U9083 ( .B1(n7732), .B2(n8206), .A(n7731), .ZN(n11004) );
  INV_X1 U9084 ( .A(n7733), .ZN(n7735) );
  INV_X1 U9085 ( .A(n7916), .ZN(n7734) );
  OAI21_X1 U9086 ( .B1(n5276), .B2(n7735), .A(n7734), .ZN(n11001) );
  AOI22_X1 U9087 ( .A1(n10821), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7736), .B2(
        n10813), .ZN(n7739) );
  NAND2_X1 U9088 ( .A1(n7737), .A2(n10767), .ZN(n7738) );
  OAI211_X1 U9089 ( .C1(n11001), .C2(n8788), .A(n7739), .B(n7738), .ZN(n7740)
         );
  AOI21_X1 U9090 ( .B1(n11004), .B2(n9024), .A(n7740), .ZN(n7741) );
  OAI21_X1 U9091 ( .B1(n10821), .B2(n7742), .A(n7741), .ZN(P2_U3284) );
  NAND2_X1 U9092 ( .A1(n7743), .A2(n9506), .ZN(n7794) );
  OR2_X1 U9093 ( .A1(n10412), .A2(n7853), .ZN(n9510) );
  NAND2_X1 U9094 ( .A1(n10412), .A2(n7853), .ZN(n9511) );
  OR2_X1 U9095 ( .A1(n7744), .A2(n5030), .ZN(n7746) );
  AOI22_X1 U9096 ( .A1(n7983), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7982), .B2(
        n10568), .ZN(n7745) );
  NAND2_X1 U9097 ( .A1(n10406), .A2(n7880), .ZN(n9518) );
  NAND2_X1 U9098 ( .A1(n9517), .A2(n9518), .ZN(n9514) );
  INV_X1 U9099 ( .A(n9511), .ZN(n7747) );
  NOR2_X1 U9100 ( .A1(n9514), .A2(n7747), .ZN(n7748) );
  NAND2_X1 U9101 ( .A1(n7749), .A2(n9390), .ZN(n7752) );
  AOI22_X1 U9102 ( .A1(n7983), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7982), .B2(
        n7750), .ZN(n7751) );
  NAND2_X1 U9103 ( .A1(n8412), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7760) );
  NAND2_X1 U9104 ( .A1(n7753), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7759) );
  OR2_X1 U9105 ( .A1(n5034), .A2(n7754), .ZN(n7758) );
  OR2_X1 U9106 ( .A1(n7755), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U9107 ( .A1(n7763), .A2(n7756), .ZN(n7884) );
  OR2_X1 U9108 ( .A1(n5032), .A2(n7884), .ZN(n7757) );
  NAND2_X1 U9109 ( .A1(n7886), .A2(n9264), .ZN(n9530) );
  XNOR2_X1 U9110 ( .A(n7834), .B(n9438), .ZN(n7770) );
  NAND2_X1 U9111 ( .A1(n8412), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U9112 ( .A1(n7239), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7768) );
  OR2_X1 U9113 ( .A1(n5034), .A2(n7761), .ZN(n7767) );
  NAND2_X1 U9114 ( .A1(n7763), .A2(n7762), .ZN(n7764) );
  NAND2_X1 U9115 ( .A1(n7765), .A2(n7764), .ZN(n9268) );
  OR2_X1 U9116 ( .A1(n5032), .A2(n9268), .ZN(n7766) );
  AOI222_X1 U9117 ( .A1(n10920), .A2(n7770), .B1(n10007), .B2(n10842), .C1(
        n10009), .C2(n10843), .ZN(n10995) );
  OR2_X1 U9118 ( .A1(n7773), .A2(n10011), .ZN(n7771) );
  NAND2_X1 U9119 ( .A1(n7772), .A2(n7771), .ZN(n7775) );
  NAND2_X1 U9120 ( .A1(n7773), .A2(n10011), .ZN(n7774) );
  NAND2_X1 U9121 ( .A1(n7775), .A2(n7774), .ZN(n7788) );
  OR2_X1 U9122 ( .A1(n10412), .A2(n10010), .ZN(n7776) );
  NAND2_X1 U9123 ( .A1(n7824), .A2(n9514), .ZN(n7849) );
  OR2_X1 U9124 ( .A1(n10406), .A2(n10009), .ZN(n7777) );
  AND2_X1 U9125 ( .A1(n7849), .A2(n7777), .ZN(n7779) );
  NAND2_X1 U9126 ( .A1(n7849), .A2(n7826), .ZN(n7778) );
  OAI21_X1 U9127 ( .B1(n7779), .B2(n9438), .A(n7778), .ZN(n7780) );
  INV_X1 U9128 ( .A(n7780), .ZN(n10998) );
  INV_X1 U9129 ( .A(n10300), .ZN(n10309) );
  NAND2_X1 U9130 ( .A1(n10998), .A2(n10309), .ZN(n7785) );
  INV_X1 U9131 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7781) );
  OAI22_X1 U9132 ( .A1(n10942), .A2(n7781), .B1(n7884), .B2(n10937), .ZN(n7783) );
  INV_X1 U9133 ( .A(n10406), .ZN(n7861) );
  INV_X1 U9134 ( .A(n7886), .ZN(n10996) );
  OAI211_X1 U9135 ( .C1(n7857), .C2(n10996), .A(n10711), .B(n5102), .ZN(n10994) );
  NOR2_X1 U9136 ( .A1(n10994), .A2(n10313), .ZN(n7782) );
  AOI211_X1 U9137 ( .C1(n10317), .C2(n7886), .A(n7783), .B(n7782), .ZN(n7784)
         );
  OAI211_X1 U9138 ( .C1(n10296), .C2(n10995), .A(n7785), .B(n7784), .ZN(
        P1_U3279) );
  INV_X1 U9139 ( .A(n7786), .ZN(n7787) );
  AOI21_X1 U9140 ( .B1(n9429), .B2(n7788), .A(n7787), .ZN(n10416) );
  AOI211_X1 U9141 ( .C1(n10412), .C2(n7789), .A(n11043), .B(n7856), .ZN(n10411) );
  INV_X1 U9142 ( .A(n10412), .ZN(n7793) );
  INV_X1 U9143 ( .A(n7790), .ZN(n7791) );
  AOI22_X1 U9144 ( .A1(n10296), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7791), .B2(
        n10724), .ZN(n7792) );
  OAI21_X1 U9145 ( .B1(n7793), .B2(n10935), .A(n7792), .ZN(n7797) );
  OAI21_X1 U9146 ( .B1(n9429), .B2(n7794), .A(n7850), .ZN(n7795) );
  AOI222_X1 U9147 ( .A1(n10920), .A2(n7795), .B1(n10009), .B2(n10842), .C1(
        n10011), .C2(n10843), .ZN(n10414) );
  NOR2_X1 U9148 ( .A1(n10414), .A2(n10296), .ZN(n7796) );
  AOI211_X1 U9149 ( .C1(n10411), .C2(n10281), .A(n7797), .B(n7796), .ZN(n7798)
         );
  OAI21_X1 U9150 ( .B1(n10416), .B2(n10300), .A(n7798), .ZN(P1_U3281) );
  INV_X1 U9151 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U9152 ( .A1(n7957), .A2(n10450), .ZN(n7801) );
  INV_X1 U9153 ( .A(n7799), .ZN(n7800) );
  NAND2_X1 U9154 ( .A1(n7800), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9605) );
  OAI211_X1 U9155 ( .C1(n7958), .C2(n10454), .A(n7801), .B(n9605), .ZN(
        P1_U3330) );
  NAND2_X1 U9156 ( .A1(n10406), .A2(n7802), .ZN(n7804) );
  NAND2_X1 U9157 ( .A1(n10009), .A2(n9181), .ZN(n7803) );
  NAND2_X1 U9158 ( .A1(n7804), .A2(n7803), .ZN(n7805) );
  XNOR2_X1 U9159 ( .A(n7805), .B(n8418), .ZN(n7866) );
  NOR2_X1 U9160 ( .A1(n7880), .A2(n8396), .ZN(n7806) );
  AOI21_X1 U9161 ( .B1(n10406), .B2(n9181), .A(n7806), .ZN(n7867) );
  XNOR2_X1 U9162 ( .A(n7866), .B(n7867), .ZN(n7809) );
  NAND2_X1 U9163 ( .A1(n7808), .A2(n7809), .ZN(n7870) );
  OAI21_X1 U9164 ( .B1(n7809), .B2(n7808), .A(n7870), .ZN(n7810) );
  NAND2_X1 U9165 ( .A1(n7810), .A2(n9295), .ZN(n7815) );
  INV_X1 U9166 ( .A(n7811), .ZN(n7859) );
  INV_X1 U9167 ( .A(n9264), .ZN(n10008) );
  AND2_X1 U9168 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10561) );
  AOI21_X1 U9169 ( .B1(n10008), .B2(n9318), .A(n10561), .ZN(n7812) );
  OAI21_X1 U9170 ( .B1(n7853), .B2(n9314), .A(n7812), .ZN(n7813) );
  AOI21_X1 U9171 ( .B1(n7859), .B2(n9303), .A(n7813), .ZN(n7814) );
  OAI211_X1 U9172 ( .C1(n7861), .C2(n9321), .A(n7815), .B(n7814), .ZN(P1_U3234) );
  NAND2_X1 U9173 ( .A1(n7957), .A2(n7816), .ZN(n7817) );
  OAI211_X1 U9174 ( .C1(n7818), .C2(n9146), .A(n7817), .B(n8244), .ZN(P2_U3335) );
  NAND2_X1 U9175 ( .A1(n7886), .A2(n10008), .ZN(n7825) );
  AND2_X1 U9176 ( .A1(n9514), .A2(n7825), .ZN(n7828) );
  NAND2_X1 U9177 ( .A1(n7819), .A2(n9390), .ZN(n7822) );
  AOI22_X1 U9178 ( .A1(n7983), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7982), .B2(
        n7820), .ZN(n7821) );
  OR2_X1 U9179 ( .A1(n10398), .A2(n10303), .ZN(n9527) );
  NAND2_X1 U9180 ( .A1(n10398), .A2(n10303), .ZN(n9523) );
  AND2_X1 U9181 ( .A1(n7828), .A2(n7836), .ZN(n7823) );
  INV_X1 U9182 ( .A(n7825), .ZN(n7827) );
  AND2_X1 U9183 ( .A1(n8445), .A2(n8443), .ZN(n7833) );
  NAND2_X1 U9184 ( .A1(n7824), .A2(n7828), .ZN(n7830) );
  AND2_X1 U9185 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  NAND2_X1 U9186 ( .A1(n7831), .A2(n9440), .ZN(n7832) );
  NAND2_X1 U9187 ( .A1(n7833), .A2(n7832), .ZN(n10404) );
  INV_X1 U9188 ( .A(n10404), .ZN(n7848) );
  INV_X1 U9189 ( .A(n9438), .ZN(n9521) );
  NAND2_X1 U9190 ( .A1(n7835), .A2(n9526), .ZN(n7837) );
  NAND2_X1 U9191 ( .A1(n7837), .A2(n7836), .ZN(n7838) );
  NAND2_X1 U9192 ( .A1(n5467), .A2(n7838), .ZN(n7839) );
  NAND2_X1 U9193 ( .A1(n7839), .A2(n10920), .ZN(n7841) );
  AOI22_X1 U9194 ( .A1(n10008), .A2(n10843), .B1(n10842), .B2(n10293), .ZN(
        n7840) );
  NAND2_X1 U9195 ( .A1(n7841), .A2(n7840), .ZN(n10402) );
  AOI21_X1 U9196 ( .B1(n5102), .B2(n10398), .A(n11043), .ZN(n7842) );
  NAND2_X1 U9197 ( .A1(n7842), .A2(n10311), .ZN(n10399) );
  INV_X1 U9198 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7843) );
  OAI22_X1 U9199 ( .A1(n10942), .A2(n7843), .B1(n9268), .B2(n10937), .ZN(n7844) );
  AOI21_X1 U9200 ( .B1(n10398), .B2(n10317), .A(n7844), .ZN(n7845) );
  OAI21_X1 U9201 ( .B1(n10399), .B2(n10313), .A(n7845), .ZN(n7846) );
  AOI21_X1 U9202 ( .B1(n10402), .B2(n10942), .A(n7846), .ZN(n7847) );
  OAI21_X1 U9203 ( .B1(n7848), .B2(n10300), .A(n7847), .ZN(P1_U3278) );
  OAI21_X1 U9204 ( .B1(n7824), .B2(n9514), .A(n7849), .ZN(n7862) );
  NAND2_X1 U9205 ( .A1(n7850), .A2(n9511), .ZN(n7851) );
  XNOR2_X1 U9206 ( .A(n7851), .B(n9514), .ZN(n7852) );
  NOR2_X1 U9207 ( .A1(n7852), .A2(n10848), .ZN(n7855) );
  OAI22_X1 U9208 ( .A1(n7853), .A2(n10915), .B1(n9264), .B2(n10917), .ZN(n7854) );
  AOI211_X1 U9209 ( .C1(n7862), .C2(n10840), .A(n7855), .B(n7854), .ZN(n10409)
         );
  INV_X1 U9210 ( .A(n7856), .ZN(n7858) );
  AOI21_X1 U9211 ( .B1(n10406), .B2(n7858), .A(n7857), .ZN(n10407) );
  AOI22_X1 U9212 ( .A1(n10296), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7859), .B2(
        n10724), .ZN(n7860) );
  OAI21_X1 U9213 ( .B1(n7861), .B2(n10935), .A(n7860), .ZN(n7864) );
  INV_X1 U9214 ( .A(n7862), .ZN(n10410) );
  NOR2_X1 U9215 ( .A1(n10410), .A2(n10264), .ZN(n7863) );
  AOI211_X1 U9216 ( .C1(n10407), .C2(n10932), .A(n7864), .B(n7863), .ZN(n7865)
         );
  OAI21_X1 U9217 ( .B1(n10296), .B2(n10409), .A(n7865), .ZN(P1_U3280) );
  INV_X1 U9218 ( .A(n7866), .ZN(n7868) );
  NAND2_X1 U9219 ( .A1(n7868), .A2(n7867), .ZN(n7869) );
  NAND2_X1 U9220 ( .A1(n7886), .A2(n7802), .ZN(n7872) );
  NAND2_X1 U9221 ( .A1(n10008), .A2(n9181), .ZN(n7871) );
  NAND2_X1 U9222 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  XNOR2_X1 U9223 ( .A(n7873), .B(n9185), .ZN(n7875) );
  NOR2_X1 U9224 ( .A1(n9264), .A2(n8396), .ZN(n7874) );
  AOI21_X1 U9225 ( .B1(n7886), .B2(n9181), .A(n7874), .ZN(n7876) );
  INV_X1 U9226 ( .A(n7875), .ZN(n7878) );
  INV_X1 U9227 ( .A(n7876), .ZN(n7877) );
  NAND2_X1 U9228 ( .A1(n7878), .A2(n7877), .ZN(n8266) );
  NAND2_X1 U9229 ( .A1(n5103), .A2(n8266), .ZN(n7879) );
  XNOR2_X1 U9230 ( .A(n8267), .B(n7879), .ZN(n7888) );
  NOR2_X1 U9231 ( .A1(n9314), .A2(n7880), .ZN(n7881) );
  AOI211_X1 U9232 ( .C1(n9318), .C2(n10007), .A(n7882), .B(n7881), .ZN(n7883)
         );
  OAI21_X1 U9233 ( .B1(n9315), .B2(n7884), .A(n7883), .ZN(n7885) );
  AOI21_X1 U9234 ( .B1(n7886), .B2(n9220), .A(n7885), .ZN(n7887) );
  OAI21_X1 U9235 ( .B1(n7888), .B2(n9309), .A(n7887), .ZN(P1_U3222) );
  OAI222_X1 U9236 ( .A1(n9147), .A2(n7993), .B1(P2_U3152), .B2(n7890), .C1(
        n7889), .C2(n9146), .ZN(P2_U3334) );
  INV_X1 U9237 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7994) );
  OAI222_X1 U9238 ( .A1(n7891), .A2(P1_U3084), .B1(n10461), .B2(n7993), .C1(
        n7994), .C2(n10454), .ZN(P1_U3329) );
  INV_X1 U9239 ( .A(n7892), .ZN(n7893) );
  AOI21_X1 U9240 ( .B1(n7895), .B2(n7894), .A(n7893), .ZN(n7901) );
  NAND2_X1 U9241 ( .A1(n10884), .A2(n8659), .ZN(n7897) );
  OAI211_X1 U9242 ( .C1(n7915), .C2(n10886), .A(n7897), .B(n7896), .ZN(n7899)
         );
  NOR2_X1 U9243 ( .A1(n11010), .A2(n6439), .ZN(n7898) );
  AOI211_X1 U9244 ( .C1(n6450), .C2(n7919), .A(n7899), .B(n7898), .ZN(n7900)
         );
  OAI21_X1 U9245 ( .B1(n7901), .B2(n10890), .A(n7900), .ZN(P2_U3236) );
  OAI211_X1 U9246 ( .C1(n5099), .C2(n6241), .A(n10808), .B(n7902), .ZN(n7904)
         );
  AOI22_X1 U9247 ( .A1(n8658), .A2(n9016), .B1(n9014), .B2(n8660), .ZN(n7903)
         );
  NAND2_X1 U9248 ( .A1(n7904), .A2(n7903), .ZN(n11033) );
  INV_X1 U9249 ( .A(n11033), .ZN(n7912) );
  OAI21_X1 U9250 ( .B1(n5107), .B2(n8207), .A(n7905), .ZN(n11035) );
  XNOR2_X1 U9251 ( .A(n11029), .B(n7917), .ZN(n11031) );
  INV_X1 U9252 ( .A(n7936), .ZN(n7906) );
  OAI22_X1 U9253 ( .A1(n10818), .A2(n7312), .B1(n7906), .B2(n8987), .ZN(n7907)
         );
  AOI21_X1 U9254 ( .B1(n7908), .B2(n10767), .A(n7907), .ZN(n7909) );
  OAI21_X1 U9255 ( .B1(n11031), .B2(n8788), .A(n7909), .ZN(n7910) );
  AOI21_X1 U9256 ( .B1(n11035), .B2(n9024), .A(n7910), .ZN(n7911) );
  OAI21_X1 U9257 ( .B1(n10821), .B2(n7912), .A(n7911), .ZN(P2_U3282) );
  XOR2_X1 U9258 ( .A(n7913), .B(n8208), .Z(n7914) );
  OAI222_X1 U9259 ( .A1(n10794), .A2(n8646), .B1(n10792), .B2(n7915), .C1(
        n8932), .C2(n7914), .ZN(n11012) );
  NOR2_X1 U9260 ( .A1(n11010), .A2(n7916), .ZN(n7918) );
  OR2_X1 U9261 ( .A1(n7918), .A2(n7917), .ZN(n11011) );
  INV_X1 U9262 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7921) );
  INV_X1 U9263 ( .A(n7919), .ZN(n7920) );
  OAI22_X1 U9264 ( .A1(n10818), .A2(n7921), .B1(n7920), .B2(n8987), .ZN(n7922)
         );
  AOI21_X1 U9265 ( .B1(n8107), .B2(n10767), .A(n7922), .ZN(n7923) );
  OAI21_X1 U9266 ( .B1(n11011), .B2(n8788), .A(n7923), .ZN(n7927) );
  INV_X1 U9267 ( .A(n11014), .ZN(n7925) );
  AND2_X1 U9268 ( .A1(n7924), .A2(n8208), .ZN(n11009) );
  NOR3_X1 U9269 ( .A1(n7925), .A2(n11009), .A3(n9008), .ZN(n7926) );
  AOI211_X1 U9270 ( .C1(n10818), .C2(n11012), .A(n7927), .B(n7926), .ZN(n7928)
         );
  INV_X1 U9271 ( .A(n7928), .ZN(P2_U3283) );
  OAI21_X1 U9272 ( .B1(n7931), .B2(n7929), .A(n7930), .ZN(n7932) );
  NAND2_X1 U9273 ( .A1(n7932), .A2(n10964), .ZN(n7938) );
  AOI21_X1 U9274 ( .B1(n10884), .B2(n8658), .A(n7933), .ZN(n7934) );
  OAI21_X1 U9275 ( .B1(n8106), .B2(n10886), .A(n7934), .ZN(n7935) );
  AOI21_X1 U9276 ( .B1(n7936), .B2(n6450), .A(n7935), .ZN(n7937) );
  OAI211_X1 U9277 ( .C1(n11029), .C2(n6439), .A(n7938), .B(n7937), .ZN(
        P2_U3217) );
  XNOR2_X1 U9278 ( .A(n7939), .B(n7945), .ZN(n7940) );
  AOI222_X1 U9279 ( .A1(n10808), .A2(n7940), .B1(n8657), .B2(n9016), .C1(n8659), .C2(n9014), .ZN(n9112) );
  INV_X1 U9280 ( .A(n8999), .ZN(n7941) );
  AOI21_X1 U9281 ( .B1(n9109), .B2(n7942), .A(n7941), .ZN(n9110) );
  INV_X1 U9282 ( .A(n9109), .ZN(n8651) );
  AOI22_X1 U9283 ( .A1(n10821), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8648), .B2(
        n10813), .ZN(n7943) );
  OAI21_X1 U9284 ( .B1(n8651), .B2(n8963), .A(n7943), .ZN(n7947) );
  INV_X1 U9285 ( .A(n7945), .ZN(n8210) );
  XNOR2_X1 U9286 ( .A(n7944), .B(n8210), .ZN(n9113) );
  NOR2_X1 U9287 ( .A1(n9113), .A2(n9008), .ZN(n7946) );
  AOI211_X1 U9288 ( .C1(n9110), .C2(n10764), .A(n7947), .B(n7946), .ZN(n7948)
         );
  OAI21_X1 U9289 ( .B1(n10821), .B2(n9112), .A(n7948), .ZN(P2_U3281) );
  NAND2_X1 U9290 ( .A1(n8495), .A2(n9390), .ZN(n7950) );
  INV_X1 U9291 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10448) );
  OR2_X1 U9292 ( .A1(n7060), .A2(n10448), .ZN(n7949) );
  NAND2_X1 U9293 ( .A1(n10451), .A2(n9390), .ZN(n7952) );
  OR2_X1 U9294 ( .A1(n7060), .A2(n7034), .ZN(n7951) );
  INV_X1 U9295 ( .A(n10333), .ZN(n10096) );
  NAND2_X1 U9296 ( .A1(n9142), .A2(n9390), .ZN(n7954) );
  INV_X1 U9297 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10455) );
  OR2_X1 U9298 ( .A1(n7060), .A2(n10455), .ZN(n7953) );
  NAND2_X1 U9299 ( .A1(n9145), .A2(n9390), .ZN(n7956) );
  INV_X1 U9300 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10459) );
  OR2_X1 U9301 ( .A1(n7060), .A2(n10459), .ZN(n7955) );
  INV_X1 U9302 ( .A(n10343), .ZN(n10131) );
  NAND2_X1 U9303 ( .A1(n7957), .A2(n9390), .ZN(n7960) );
  OR2_X1 U9304 ( .A1(n7060), .A2(n7958), .ZN(n7959) );
  NAND2_X1 U9305 ( .A1(n7961), .A2(n9390), .ZN(n7964) );
  OR2_X1 U9306 ( .A1(n7060), .A2(n7962), .ZN(n7963) );
  NAND2_X1 U9307 ( .A1(n7965), .A2(n9390), .ZN(n7967) );
  AOI22_X1 U9308 ( .A1(n7983), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7982), .B2(
        n10035), .ZN(n7966) );
  NOR2_X1 U9309 ( .A1(n10311), .A2(n10316), .ZN(n10284) );
  NAND2_X1 U9310 ( .A1(n7968), .A2(n9390), .ZN(n7971) );
  INV_X1 U9311 ( .A(n10047), .ZN(n7969) );
  AOI22_X1 U9312 ( .A1(n7983), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7982), .B2(
        n7969), .ZN(n7970) );
  INV_X1 U9313 ( .A(n10393), .ZN(n10290) );
  NAND2_X1 U9314 ( .A1(n10284), .A2(n10290), .ZN(n10285) );
  NAND2_X1 U9315 ( .A1(n7972), .A2(n9390), .ZN(n7974) );
  AOI22_X1 U9316 ( .A1(n7983), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7982), .B2(
        n10066), .ZN(n7973) );
  OR2_X1 U9317 ( .A1(n7975), .A2(n5030), .ZN(n7977) );
  AOI22_X1 U9318 ( .A1(n7983), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7982), .B2(
        n10078), .ZN(n7976) );
  INV_X1 U9319 ( .A(n10383), .ZN(n10263) );
  NAND2_X1 U9320 ( .A1(n10269), .A2(n10263), .ZN(n10257) );
  OR2_X1 U9321 ( .A1(n7978), .A2(n5030), .ZN(n7980) );
  AOI22_X1 U9322 ( .A1(n7983), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7982), .B2(
        n10586), .ZN(n7979) );
  NOR2_X1 U9323 ( .A1(n10257), .A2(n10378), .ZN(n10236) );
  NAND2_X1 U9324 ( .A1(n7981), .A2(n9390), .ZN(n7985) );
  AOI22_X1 U9325 ( .A1(n7983), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10730), 
        .B2(n7982), .ZN(n7984) );
  INV_X1 U9326 ( .A(n10374), .ZN(n8332) );
  NAND2_X1 U9327 ( .A1(n10236), .A2(n8332), .ZN(n10226) );
  NAND2_X1 U9328 ( .A1(n7986), .A2(n9390), .ZN(n7988) );
  OR2_X1 U9329 ( .A1(n7060), .A2(n9612), .ZN(n7987) );
  OR2_X1 U9330 ( .A1(n7989), .A2(n5030), .ZN(n7992) );
  OR2_X1 U9331 ( .A1(n7060), .A2(n7990), .ZN(n7991) );
  INV_X1 U9332 ( .A(n10364), .ZN(n10188) );
  OR2_X1 U9333 ( .A1(n7060), .A2(n7994), .ZN(n7995) );
  NAND2_X1 U9334 ( .A1(n10131), .A2(n10146), .ZN(n10125) );
  NAND2_X1 U9335 ( .A1(n9136), .A2(n9390), .ZN(n7998) );
  OR2_X1 U9336 ( .A1(n7060), .A2(n10445), .ZN(n7997) );
  NOR2_X2 U9337 ( .A1(n8473), .A2(n10323), .ZN(n8472) );
  INV_X1 U9338 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8516) );
  INV_X1 U9339 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8498) );
  MUX2_X1 U9340 ( .A(n8516), .B(n8498), .S(n8021), .Z(n8004) );
  INV_X1 U9341 ( .A(SI_30_), .ZN(n8003) );
  NAND2_X1 U9342 ( .A1(n8004), .A2(n8003), .ZN(n8019) );
  INV_X1 U9343 ( .A(n8004), .ZN(n8005) );
  NAND2_X1 U9344 ( .A1(n8005), .A2(SI_30_), .ZN(n8006) );
  AND2_X1 U9345 ( .A1(n8019), .A2(n8006), .ZN(n8017) );
  NAND2_X1 U9346 ( .A1(n8497), .A2(n9390), .ZN(n8008) );
  OR2_X1 U9347 ( .A1(n7060), .A2(n8516), .ZN(n8007) );
  NAND2_X1 U9348 ( .A1(n8472), .A2(n8014), .ZN(n10085) );
  OAI21_X1 U9349 ( .B1(n8472), .B2(n8014), .A(n10085), .ZN(n11044) );
  INV_X1 U9350 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n8011) );
  NAND2_X1 U9351 ( .A1(n7753), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8010) );
  NAND2_X1 U9352 ( .A1(n8412), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8009) );
  OAI211_X1 U9353 ( .C1(n5034), .C2(n8011), .A(n8010), .B(n8009), .ZN(n9607)
         );
  NOR2_X1 U9354 ( .A1(n10510), .A2(n8012), .ZN(n8013) );
  NOR2_X1 U9355 ( .A1(n10917), .A2(n8013), .ZN(n8490) );
  NAND2_X1 U9356 ( .A1(n9607), .A2(n8490), .ZN(n11042) );
  NOR2_X1 U9357 ( .A1(n10296), .A2(n11042), .ZN(n10086) );
  NOR2_X1 U9358 ( .A1(n8014), .A2(n10935), .ZN(n8015) );
  AOI211_X1 U9359 ( .C1(n10296), .C2(P1_REG2_REG_30__SCAN_IN), .A(n10086), .B(
        n8015), .ZN(n8016) );
  OAI21_X1 U9360 ( .B1(n10702), .B2(n11044), .A(n8016), .ZN(P1_U3262) );
  NAND2_X1 U9361 ( .A1(n8018), .A2(n8017), .ZN(n8020) );
  MUX2_X1 U9362 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n8021), .Z(n8023) );
  INV_X1 U9363 ( .A(SI_31_), .ZN(n8022) );
  XNOR2_X1 U9364 ( .A(n8023), .B(n8022), .ZN(n8024) );
  NAND2_X1 U9365 ( .A1(n9391), .A2(n8036), .ZN(n8028) );
  INV_X1 U9366 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8026) );
  OR2_X1 U9367 ( .A1(n5825), .A2(n8026), .ZN(n8027) );
  NAND2_X1 U9368 ( .A1(n8029), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U9369 ( .A1(n8030), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8032) );
  NAND2_X1 U9370 ( .A1(n5801), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8031) );
  OR2_X1 U9371 ( .A1(n9032), .A2(n8652), .ZN(n8039) );
  INV_X1 U9372 ( .A(n8039), .ZN(n8187) );
  OR2_X1 U9373 ( .A1(n8241), .A2(n8034), .ZN(n8035) );
  NAND2_X1 U9374 ( .A1(n8497), .A2(n8036), .ZN(n8038) );
  OR2_X1 U9375 ( .A1(n5825), .A2(n8498), .ZN(n8037) );
  INV_X1 U9376 ( .A(n8653), .ZN(n8180) );
  NAND2_X1 U9377 ( .A1(n9038), .A2(n8180), .ZN(n8182) );
  AND2_X1 U9378 ( .A1(n8039), .A2(n8182), .ZN(n8191) );
  AND2_X1 U9379 ( .A1(n8157), .A2(n8155), .ZN(n8152) );
  NAND3_X1 U9380 ( .A1(n8041), .A2(n8040), .A3(n8227), .ZN(n8042) );
  NAND2_X1 U9381 ( .A1(n8193), .A2(n8042), .ZN(n8045) );
  OAI21_X1 U9382 ( .B1(n8045), .B2(n8044), .A(n8043), .ZN(n8050) );
  OR2_X1 U9383 ( .A1(n8047), .A2(n8046), .ZN(n8195) );
  MUX2_X1 U9384 ( .A(n8052), .B(n8051), .S(n8186), .Z(n8053) );
  NAND2_X1 U9385 ( .A1(n8055), .A2(n8194), .ZN(n8059) );
  MUX2_X1 U9386 ( .A(n8057), .B(n8056), .S(n8186), .Z(n8058) );
  INV_X1 U9387 ( .A(n8060), .ZN(n8061) );
  MUX2_X1 U9388 ( .A(n8062), .B(n8061), .S(n8186), .Z(n8064) );
  NOR2_X1 U9389 ( .A1(n8664), .A2(n10863), .ZN(n8063) );
  MUX2_X1 U9390 ( .A(n8664), .B(n10863), .S(n8186), .Z(n8067) );
  OAI22_X1 U9391 ( .A1(n8065), .A2(n8064), .B1(n8063), .B2(n8067), .ZN(n8069)
         );
  NAND2_X1 U9392 ( .A1(n8067), .A2(n8066), .ZN(n8068) );
  NAND2_X1 U9393 ( .A1(n8069), .A2(n8068), .ZN(n8075) );
  MUX2_X1 U9394 ( .A(n8071), .B(n8070), .S(n8186), .Z(n8072) );
  NAND2_X1 U9395 ( .A1(n8201), .A2(n8072), .ZN(n8073) );
  AOI21_X1 U9396 ( .B1(n8075), .B2(n8074), .A(n8073), .ZN(n8083) );
  INV_X1 U9397 ( .A(n8086), .ZN(n8082) );
  NOR2_X1 U9398 ( .A1(n8077), .A2(n8076), .ZN(n8080) );
  NAND2_X1 U9399 ( .A1(n8084), .A2(n8078), .ZN(n8079) );
  MUX2_X1 U9400 ( .A(n8080), .B(n8079), .S(n8155), .Z(n8081) );
  AND2_X1 U9401 ( .A1(n8088), .A2(n8084), .ZN(n8085) );
  MUX2_X1 U9402 ( .A(n8086), .B(n8085), .S(n8186), .Z(n8087) );
  AND2_X1 U9403 ( .A1(n8094), .A2(n8088), .ZN(n8091) );
  AND2_X1 U9404 ( .A1(n8096), .A2(n8089), .ZN(n8090) );
  NAND2_X1 U9405 ( .A1(n8098), .A2(n8094), .ZN(n8095) );
  NAND2_X1 U9406 ( .A1(n8095), .A2(n8097), .ZN(n8101) );
  NAND2_X1 U9407 ( .A1(n8097), .A2(n8096), .ZN(n8099) );
  NAND2_X1 U9408 ( .A1(n8099), .A2(n8098), .ZN(n8100) );
  MUX2_X1 U9409 ( .A(n8101), .B(n8100), .S(n8155), .Z(n8102) );
  NAND2_X1 U9410 ( .A1(n8660), .A2(n8186), .ZN(n8109) );
  NAND2_X1 U9411 ( .A1(n8106), .A2(n8155), .ZN(n8108) );
  MUX2_X1 U9412 ( .A(n8109), .B(n8108), .S(n8107), .Z(n8110) );
  NAND3_X1 U9413 ( .A1(n6241), .A2(n8111), .A3(n8110), .ZN(n8115) );
  MUX2_X1 U9414 ( .A(n8113), .B(n8112), .S(n8155), .Z(n8114) );
  INV_X1 U9415 ( .A(n9006), .ZN(n8995) );
  MUX2_X1 U9416 ( .A(n8994), .B(n8116), .S(n8186), .Z(n8117) );
  MUX2_X1 U9417 ( .A(n8120), .B(n8119), .S(n8155), .Z(n8121) );
  MUX2_X1 U9418 ( .A(n8124), .B(n8123), .S(n8186), .Z(n8125) );
  INV_X1 U9419 ( .A(n8591), .ZN(n8656) );
  MUX2_X1 U9420 ( .A(n8656), .B(n9094), .S(n8155), .Z(n8134) );
  NAND2_X1 U9421 ( .A1(n8128), .A2(n8656), .ZN(n8130) );
  NAND2_X1 U9422 ( .A1(n8130), .A2(n8129), .ZN(n8132) );
  MUX2_X1 U9423 ( .A(n8919), .B(n9084), .S(n8155), .Z(n8136) );
  INV_X1 U9424 ( .A(n8136), .ZN(n8137) );
  OAI21_X1 U9425 ( .B1(n8139), .B2(n8138), .A(n8137), .ZN(n8140) );
  NAND2_X1 U9426 ( .A1(n8145), .A2(n8144), .ZN(n8146) );
  NAND2_X1 U9427 ( .A1(n8146), .A2(n8155), .ZN(n8148) );
  INV_X1 U9428 ( .A(n8150), .ZN(n8147) );
  AOI21_X1 U9429 ( .B1(n8150), .B2(n8149), .A(n8155), .ZN(n8151) );
  NAND2_X1 U9430 ( .A1(n8164), .A2(n8154), .ZN(n8156) );
  NAND2_X1 U9431 ( .A1(n8158), .A2(n8157), .ZN(n8159) );
  NAND2_X1 U9432 ( .A1(n8165), .A2(n8162), .ZN(n8163) );
  NAND2_X1 U9433 ( .A1(n8165), .A2(n8164), .ZN(n8166) );
  INV_X1 U9434 ( .A(n8170), .ZN(n8168) );
  MUX2_X1 U9435 ( .A(n8175), .B(n8174), .S(n8186), .Z(n8176) );
  NAND3_X1 U9436 ( .A1(n8803), .A2(n8186), .A3(n8654), .ZN(n8178) );
  NAND3_X1 U9437 ( .A1(n9041), .A2(n8823), .A3(n8155), .ZN(n8177) );
  NAND4_X1 U9438 ( .A1(n8179), .A2(n8217), .A3(n8178), .A4(n8177), .ZN(n8183)
         );
  OR2_X1 U9439 ( .A1(n9038), .A2(n8180), .ZN(n8229) );
  MUX2_X1 U9440 ( .A(n8223), .B(n8225), .S(n8186), .Z(n8181) );
  NAND4_X1 U9441 ( .A1(n8183), .A2(n8229), .A3(n8182), .A4(n8181), .ZN(n8184)
         );
  OAI21_X1 U9442 ( .B1(n8191), .B2(n8186), .A(n8184), .ZN(n8185) );
  NAND2_X1 U9443 ( .A1(n9032), .A2(n8652), .ZN(n8231) );
  NAND2_X1 U9444 ( .A1(n8231), .A2(n8229), .ZN(n8219) );
  INV_X1 U9445 ( .A(n8191), .ZN(n8228) );
  NAND4_X1 U9446 ( .A1(n8194), .A2(n5348), .A3(n8193), .A4(n6229), .ZN(n8199)
         );
  INV_X1 U9447 ( .A(n8195), .ZN(n8197) );
  INV_X1 U9448 ( .A(n10805), .ZN(n8196) );
  NAND2_X1 U9449 ( .A1(n8197), .A2(n8196), .ZN(n8198) );
  NOR4_X1 U9450 ( .A1(n8200), .A2(n8199), .A3(n5145), .A4(n8198), .ZN(n8202)
         );
  NAND4_X1 U9451 ( .A1(n8204), .A2(n8203), .A3(n8202), .A4(n8201), .ZN(n8205)
         );
  NOR4_X1 U9452 ( .A1(n8207), .A2(n8206), .A3(n5942), .A4(n8205), .ZN(n8209)
         );
  NAND4_X1 U9453 ( .A1(n8978), .A2(n8210), .A3(n8209), .A4(n8208), .ZN(n8211)
         );
  NOR4_X1 U9454 ( .A1(n8943), .A2(n9006), .A3(n8212), .A4(n8211), .ZN(n8214)
         );
  NAND4_X1 U9455 ( .A1(n8916), .A2(n8899), .A3(n8214), .A4(n8213), .ZN(n8215)
         );
  NOR4_X1 U9456 ( .A1(n8866), .A2(n8876), .A3(n8852), .A4(n8215), .ZN(n8216)
         );
  NAND4_X1 U9457 ( .A1(n8217), .A2(n8813), .A3(n8835), .A4(n8216), .ZN(n8218)
         );
  NOR4_X1 U9458 ( .A1(n8228), .A2(n8219), .A3(n8805), .A4(n8218), .ZN(n8220)
         );
  XNOR2_X1 U9459 ( .A(n8220), .B(n10815), .ZN(n8221) );
  AOI211_X1 U9460 ( .C1(n8222), .C2(n5028), .A(n8227), .B(n8221), .ZN(n8238)
         );
  INV_X1 U9461 ( .A(n8223), .ZN(n8224) );
  OAI211_X1 U9462 ( .C1(n8230), .C2(n9038), .A(n8652), .B(n8227), .ZN(n8234)
         );
  AOI21_X1 U9463 ( .B1(n8230), .B2(n8229), .A(n8228), .ZN(n8233) );
  INV_X1 U9464 ( .A(n8231), .ZN(n8232) );
  INV_X1 U9465 ( .A(n8235), .ZN(n8236) );
  NOR4_X1 U9466 ( .A1(n8240), .A2(n10792), .A3(n8239), .A4(n9140), .ZN(n8243)
         );
  OAI21_X1 U9467 ( .B1(n8244), .B2(n8241), .A(P2_B_REG_SCAN_IN), .ZN(n8242) );
  NAND2_X1 U9468 ( .A1(n10333), .A2(n7802), .ZN(n8252) );
  NAND2_X1 U9469 ( .A1(n8412), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U9470 ( .A1(n7753), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8249) );
  INV_X1 U9471 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8245) );
  OR2_X1 U9472 ( .A1(n5034), .A2(n8245), .ZN(n8248) );
  INV_X1 U9473 ( .A(n8410), .ZN(n8246) );
  NAND2_X1 U9474 ( .A1(n8246), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8428) );
  INV_X1 U9475 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8437) );
  XNOR2_X1 U9476 ( .A(n8428), .B(n8437), .ZN(n10093) );
  OR2_X1 U9477 ( .A1(n8432), .A2(n10093), .ZN(n8247) );
  NAND2_X1 U9478 ( .A1(n9610), .A2(n9181), .ZN(n8251) );
  NAND2_X1 U9479 ( .A1(n8252), .A2(n8251), .ZN(n8253) );
  XNOR2_X1 U9480 ( .A(n8253), .B(n9185), .ZN(n8255) );
  NOR2_X1 U9481 ( .A1(n10111), .A2(n8396), .ZN(n8254) );
  AOI21_X1 U9482 ( .B1(n10333), .B2(n9181), .A(n8254), .ZN(n8256) );
  NAND2_X1 U9483 ( .A1(n8255), .A2(n8256), .ZN(n9196) );
  INV_X1 U9484 ( .A(n8255), .ZN(n8258) );
  INV_X1 U9485 ( .A(n8256), .ZN(n8257) );
  NAND2_X1 U9486 ( .A1(n8258), .A2(n8257), .ZN(n9180) );
  NAND2_X1 U9487 ( .A1(n9196), .A2(n9180), .ZN(n8425) );
  NAND2_X1 U9488 ( .A1(n7753), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8264) );
  NAND2_X1 U9489 ( .A1(n8412), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8263) );
  INV_X1 U9490 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8259) );
  OR2_X1 U9491 ( .A1(n5034), .A2(n8259), .ZN(n8262) );
  NOR2_X1 U9492 ( .A1(n8281), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8260) );
  OR2_X1 U9493 ( .A1(n8301), .A2(n8260), .ZN(n10270) );
  OR2_X1 U9494 ( .A1(n8432), .A2(n10270), .ZN(n8261) );
  AOI22_X1 U9495 ( .A1(n10389), .A2(n7802), .B1(n9181), .B2(n10294), .ZN(n8265) );
  XNOR2_X1 U9496 ( .A(n8265), .B(n8418), .ZN(n8299) );
  AOI22_X1 U9497 ( .A1(n10389), .A2(n9181), .B1(n9182), .B2(n10294), .ZN(n8298) );
  NAND2_X1 U9498 ( .A1(n10398), .A2(n7802), .ZN(n8269) );
  NAND2_X1 U9499 ( .A1(n10007), .A2(n9181), .ZN(n8268) );
  NAND2_X1 U9500 ( .A1(n8269), .A2(n8268), .ZN(n8270) );
  XNOR2_X1 U9501 ( .A(n8270), .B(n8418), .ZN(n9260) );
  NAND2_X1 U9502 ( .A1(n10398), .A2(n9181), .ZN(n8272) );
  NAND2_X1 U9503 ( .A1(n10007), .A2(n9182), .ZN(n8271) );
  NAND2_X1 U9504 ( .A1(n8272), .A2(n8271), .ZN(n9261) );
  AND2_X1 U9505 ( .A1(n10293), .A2(n9182), .ZN(n8273) );
  AOI21_X1 U9506 ( .B1(n10316), .B2(n9181), .A(n8273), .ZN(n9152) );
  INV_X1 U9507 ( .A(n9152), .ZN(n8274) );
  NOR2_X1 U9508 ( .A1(n9151), .A2(n8274), .ZN(n8293) );
  NAND2_X1 U9509 ( .A1(n10316), .A2(n7802), .ZN(n8276) );
  NAND2_X1 U9510 ( .A1(n10293), .A2(n9181), .ZN(n8275) );
  NAND2_X1 U9511 ( .A1(n8276), .A2(n8275), .ZN(n8277) );
  XNOR2_X1 U9512 ( .A(n8277), .B(n9185), .ZN(n9153) );
  NAND2_X1 U9513 ( .A1(n10393), .A2(n7802), .ZN(n8287) );
  NAND2_X1 U9514 ( .A1(n7239), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8285) );
  NAND2_X1 U9515 ( .A1(n8412), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8284) );
  INV_X1 U9516 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n8278) );
  OR2_X1 U9517 ( .A1(n5034), .A2(n8278), .ZN(n8283) );
  NOR2_X1 U9518 ( .A1(n8279), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8280) );
  OR2_X1 U9519 ( .A1(n8281), .A2(n8280), .ZN(n10287) );
  OR2_X1 U9520 ( .A1(n5032), .A2(n10287), .ZN(n8282) );
  NAND2_X1 U9521 ( .A1(n10276), .A2(n9181), .ZN(n8286) );
  NAND2_X1 U9522 ( .A1(n8287), .A2(n8286), .ZN(n8288) );
  XNOR2_X1 U9523 ( .A(n8288), .B(n9185), .ZN(n8294) );
  OAI21_X1 U9524 ( .B1(n8293), .B2(n9153), .A(n8289), .ZN(n9308) );
  NAND2_X1 U9525 ( .A1(n10393), .A2(n9181), .ZN(n8291) );
  NAND2_X1 U9526 ( .A1(n10276), .A2(n9182), .ZN(n8290) );
  NAND2_X1 U9527 ( .A1(n8291), .A2(n8290), .ZN(n9306) );
  NAND2_X1 U9528 ( .A1(n8292), .A2(n9153), .ZN(n8297) );
  INV_X1 U9529 ( .A(n8293), .ZN(n8296) );
  INV_X1 U9530 ( .A(n8294), .ZN(n8295) );
  XNOR2_X1 U9531 ( .A(n8299), .B(n8298), .ZN(n9225) );
  NAND2_X1 U9532 ( .A1(n10383), .A2(n7802), .ZN(n8308) );
  INV_X1 U9533 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8300) );
  OR2_X1 U9534 ( .A1(n5034), .A2(n8300), .ZN(n8306) );
  NOR2_X1 U9535 ( .A1(n8301), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8302) );
  OR2_X1 U9536 ( .A1(n8313), .A2(n8302), .ZN(n10260) );
  OR2_X1 U9537 ( .A1(n8432), .A2(n10260), .ZN(n8305) );
  NAND2_X1 U9538 ( .A1(n8412), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8304) );
  NAND2_X1 U9539 ( .A1(n7753), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8303) );
  NAND4_X1 U9540 ( .A1(n8306), .A2(n8305), .A3(n8304), .A4(n8303), .ZN(n10277)
         );
  NAND2_X1 U9541 ( .A1(n10277), .A2(n9181), .ZN(n8307) );
  NAND2_X1 U9542 ( .A1(n8308), .A2(n8307), .ZN(n8309) );
  XNOR2_X1 U9543 ( .A(n8309), .B(n9185), .ZN(n8312) );
  AND2_X1 U9544 ( .A1(n10277), .A2(n9182), .ZN(n8310) );
  AOI21_X1 U9545 ( .B1(n10383), .B2(n9181), .A(n8310), .ZN(n8311) );
  NOR2_X1 U9546 ( .A1(n8312), .A2(n8311), .ZN(n9233) );
  NAND2_X1 U9547 ( .A1(n8312), .A2(n8311), .ZN(n9231) );
  INV_X1 U9548 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10074) );
  OR2_X1 U9549 ( .A1(n5034), .A2(n10074), .ZN(n8320) );
  INV_X1 U9550 ( .A(n8313), .ZN(n8315) );
  INV_X1 U9551 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U9552 ( .A1(n8315), .A2(n8314), .ZN(n8316) );
  NAND2_X1 U9553 ( .A1(n8326), .A2(n8316), .ZN(n10237) );
  OR2_X1 U9554 ( .A1(n8432), .A2(n10237), .ZN(n8319) );
  NAND2_X1 U9555 ( .A1(n8412), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U9556 ( .A1(n7239), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8317) );
  NAND4_X1 U9557 ( .A1(n8320), .A2(n8319), .A3(n8318), .A4(n8317), .ZN(n10223)
         );
  AOI22_X1 U9558 ( .A1(n10378), .A2(n7802), .B1(n9181), .B2(n10223), .ZN(n8321) );
  XNOR2_X1 U9559 ( .A(n8321), .B(n8418), .ZN(n8322) );
  INV_X1 U9560 ( .A(n10378), .ZN(n10240) );
  OAI22_X1 U9561 ( .A1(n10240), .A2(n9187), .B1(n10251), .B2(n8396), .ZN(n9285) );
  NAND2_X1 U9562 ( .A1(n8323), .A2(n8322), .ZN(n9282) );
  INV_X1 U9563 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n8324) );
  OR2_X1 U9564 ( .A1(n5034), .A2(n8324), .ZN(n8331) );
  NAND2_X1 U9565 ( .A1(n8326), .A2(n8325), .ZN(n8327) );
  NAND2_X1 U9566 ( .A1(n8340), .A2(n8327), .ZN(n10231) );
  OR2_X1 U9567 ( .A1(n8432), .A2(n10231), .ZN(n8330) );
  NAND2_X1 U9568 ( .A1(n7753), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n8329) );
  NAND2_X1 U9569 ( .A1(n8412), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8328) );
  NAND4_X1 U9570 ( .A1(n8331), .A2(n8330), .A3(n8329), .A4(n8328), .ZN(n10243)
         );
  INV_X1 U9571 ( .A(n10243), .ZN(n10204) );
  OAI22_X1 U9572 ( .A1(n8332), .A2(n9187), .B1(n10204), .B2(n8396), .ZN(n8337)
         );
  NAND2_X1 U9573 ( .A1(n10374), .A2(n7802), .ZN(n8334) );
  NAND2_X1 U9574 ( .A1(n10243), .A2(n9181), .ZN(n8333) );
  NAND2_X1 U9575 ( .A1(n8334), .A2(n8333), .ZN(n8335) );
  XNOR2_X1 U9576 ( .A(n8335), .B(n8418), .ZN(n8336) );
  XOR2_X1 U9577 ( .A(n8337), .B(n8336), .Z(n9173) );
  INV_X1 U9578 ( .A(n8336), .ZN(n8339) );
  INV_X1 U9579 ( .A(n8337), .ZN(n8338) );
  NAND2_X1 U9580 ( .A1(n10368), .A2(n7802), .ZN(n8348) );
  AND2_X1 U9581 ( .A1(n8340), .A2(n9254), .ZN(n8341) );
  OR2_X1 U9582 ( .A1(n8341), .A2(n8353), .ZN(n10212) );
  INV_X1 U9583 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8342) );
  OR2_X1 U9584 ( .A1(n5034), .A2(n8342), .ZN(n8344) );
  NAND2_X1 U9585 ( .A1(n8412), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8343) );
  AND2_X1 U9586 ( .A1(n8344), .A2(n8343), .ZN(n8346) );
  NAND2_X1 U9587 ( .A1(n7239), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8345) );
  OAI211_X1 U9588 ( .C1(n10212), .C2(n8432), .A(n8346), .B(n8345), .ZN(n10224)
         );
  NAND2_X1 U9589 ( .A1(n10224), .A2(n9181), .ZN(n8347) );
  NAND2_X1 U9590 ( .A1(n8348), .A2(n8347), .ZN(n8349) );
  XNOR2_X1 U9591 ( .A(n8349), .B(n9185), .ZN(n9251) );
  AND2_X1 U9592 ( .A1(n10224), .A2(n9182), .ZN(n8350) );
  AOI21_X1 U9593 ( .B1(n10368), .B2(n9181), .A(n8350), .ZN(n8351) );
  INV_X1 U9594 ( .A(n9251), .ZN(n8352) );
  INV_X1 U9595 ( .A(n8351), .ZN(n9250) );
  NAND2_X1 U9596 ( .A1(n10364), .A2(n7802), .ZN(n8361) );
  OR2_X1 U9597 ( .A1(n8353), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8355) );
  AND2_X1 U9598 ( .A1(n8355), .A2(n8354), .ZN(n10197) );
  NAND2_X1 U9599 ( .A1(n10197), .A2(n5033), .ZN(n8359) );
  AOI22_X1 U9600 ( .A1(n8356), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n7753), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U9601 ( .A1(n8412), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8357) );
  OR2_X1 U9602 ( .A1(n10205), .A2(n9187), .ZN(n8360) );
  NAND2_X1 U9603 ( .A1(n8361), .A2(n8360), .ZN(n8362) );
  XNOR2_X1 U9604 ( .A(n8362), .B(n9185), .ZN(n8365) );
  NOR2_X1 U9605 ( .A1(n10205), .A2(n8396), .ZN(n8363) );
  AOI21_X1 U9606 ( .B1(n10364), .B2(n9181), .A(n8363), .ZN(n8364) );
  OR2_X1 U9607 ( .A1(n8365), .A2(n8364), .ZN(n9203) );
  INV_X1 U9608 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8366) );
  OR2_X1 U9609 ( .A1(n5034), .A2(n8366), .ZN(n8372) );
  OAI21_X1 U9610 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n8368), .A(n8367), .ZN(
        n10172) );
  OR2_X1 U9611 ( .A1(n5032), .A2(n10172), .ZN(n8371) );
  NAND2_X1 U9612 ( .A1(n5035), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U9613 ( .A1(n7239), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8369) );
  NAND4_X1 U9614 ( .A1(n8372), .A2(n8371), .A3(n8370), .A4(n8369), .ZN(n10192)
         );
  AOI22_X1 U9615 ( .A1(n10358), .A2(n7802), .B1(n9181), .B2(n10192), .ZN(n8373) );
  XNOR2_X1 U9616 ( .A(n8373), .B(n8418), .ZN(n8375) );
  AOI22_X1 U9617 ( .A1(n10358), .A2(n9181), .B1(n9182), .B2(n10192), .ZN(n8374) );
  NOR2_X1 U9618 ( .A1(n8375), .A2(n8374), .ZN(n9274) );
  NAND2_X1 U9619 ( .A1(n8375), .A2(n8374), .ZN(n9272) );
  NAND2_X1 U9620 ( .A1(n5035), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8381) );
  NAND2_X1 U9621 ( .A1(n7753), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8380) );
  INV_X1 U9622 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8376) );
  OR2_X1 U9623 ( .A1(n5034), .A2(n8376), .ZN(n8379) );
  OAI21_X1 U9624 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n8377), .A(n8388), .ZN(
        n10157) );
  OR2_X1 U9625 ( .A1(n5032), .A2(n10157), .ZN(n8378) );
  OAI22_X1 U9626 ( .A1(n10160), .A2(n8382), .B1(n8457), .B2(n9187), .ZN(n8383)
         );
  XOR2_X1 U9627 ( .A(n8418), .B(n8383), .Z(n8384) );
  OAI22_X1 U9628 ( .A1(n10160), .A2(n9187), .B1(n8457), .B2(n8396), .ZN(n9165)
         );
  NAND2_X1 U9629 ( .A1(n8385), .A2(n8384), .ZN(n9162) );
  OAI21_X1 U9630 ( .B1(n9164), .B2(n9165), .A(n9162), .ZN(n9242) );
  INV_X1 U9631 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8386) );
  OR2_X1 U9632 ( .A1(n5034), .A2(n8386), .ZN(n8394) );
  INV_X1 U9633 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U9634 ( .A1(n8388), .A2(n8387), .ZN(n8389) );
  NAND2_X1 U9635 ( .A1(n8390), .A2(n8389), .ZN(n9245) );
  OR2_X1 U9636 ( .A1(n8432), .A2(n9245), .ZN(n8393) );
  NAND2_X1 U9637 ( .A1(n8412), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8392) );
  NAND2_X1 U9638 ( .A1(n7239), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8391) );
  NAND4_X1 U9639 ( .A1(n8394), .A2(n8393), .A3(n8392), .A4(n8391), .ZN(n10164)
         );
  AOI22_X1 U9640 ( .A1(n10349), .A2(n7802), .B1(n9181), .B2(n10164), .ZN(n8395) );
  XOR2_X1 U9641 ( .A(n8418), .B(n8395), .Z(n8398) );
  INV_X1 U9642 ( .A(n10164), .ZN(n8482) );
  OAI22_X1 U9643 ( .A1(n5316), .A2(n9187), .B1(n8482), .B2(n8396), .ZN(n8397)
         );
  NOR2_X1 U9644 ( .A1(n8398), .A2(n8397), .ZN(n8399) );
  AOI21_X1 U9645 ( .B1(n8398), .B2(n8397), .A(n8399), .ZN(n9243) );
  NAND2_X1 U9646 ( .A1(n9242), .A2(n9243), .ZN(n9241) );
  INV_X1 U9647 ( .A(n8399), .ZN(n8400) );
  NAND2_X1 U9648 ( .A1(n9241), .A2(n8400), .ZN(n9216) );
  NAND2_X1 U9649 ( .A1(n10343), .A2(n7802), .ZN(n8402) );
  NAND2_X1 U9650 ( .A1(n10144), .A2(n9181), .ZN(n8401) );
  NAND2_X1 U9651 ( .A1(n8402), .A2(n8401), .ZN(n8403) );
  XNOR2_X1 U9652 ( .A(n8403), .B(n8418), .ZN(n8407) );
  NAND2_X1 U9653 ( .A1(n10343), .A2(n9181), .ZN(n8405) );
  NAND2_X1 U9654 ( .A1(n10144), .A2(n9182), .ZN(n8404) );
  NAND2_X1 U9655 ( .A1(n8405), .A2(n8404), .ZN(n8406) );
  NOR2_X1 U9656 ( .A1(n8407), .A2(n8406), .ZN(n9212) );
  NAND2_X1 U9657 ( .A1(n8407), .A2(n8406), .ZN(n9213) );
  INV_X1 U9658 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8408) );
  OR2_X1 U9659 ( .A1(n5034), .A2(n8408), .ZN(n8416) );
  INV_X1 U9660 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U9661 ( .A1(n8410), .A2(n8409), .ZN(n8411) );
  NAND2_X1 U9662 ( .A1(n8428), .A2(n8411), .ZN(n9299) );
  OR2_X1 U9663 ( .A1(n5032), .A2(n9299), .ZN(n8415) );
  NAND2_X1 U9664 ( .A1(n8412), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U9665 ( .A1(n7239), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8413) );
  NAND4_X1 U9666 ( .A1(n8416), .A2(n8415), .A3(n8414), .A4(n8413), .ZN(n10135)
         );
  AND2_X1 U9667 ( .A1(n10135), .A2(n9182), .ZN(n8417) );
  AOI21_X1 U9668 ( .B1(n10338), .B2(n9181), .A(n8417), .ZN(n8421) );
  AOI22_X1 U9669 ( .A1(n10338), .A2(n7802), .B1(n9181), .B2(n10135), .ZN(n8419) );
  XNOR2_X1 U9670 ( .A(n8419), .B(n8418), .ZN(n8420) );
  XOR2_X1 U9671 ( .A(n8421), .B(n8420), .Z(n9297) );
  INV_X1 U9672 ( .A(n8420), .ZN(n8423) );
  XOR2_X1 U9673 ( .A(n8425), .B(n9179), .Z(n8442) );
  NAND2_X1 U9674 ( .A1(n5035), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8436) );
  NAND2_X1 U9675 ( .A1(n7753), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8435) );
  INV_X1 U9676 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8426) );
  OR2_X1 U9677 ( .A1(n5034), .A2(n8426), .ZN(n8434) );
  INV_X1 U9678 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8427) );
  OAI21_X1 U9679 ( .B1(n8428), .B2(n8437), .A(n8427), .ZN(n8431) );
  INV_X1 U9680 ( .A(n8428), .ZN(n8430) );
  AND2_X1 U9681 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n8429) );
  NAND2_X1 U9682 ( .A1(n8430), .A2(n8429), .ZN(n8474) );
  NAND2_X1 U9683 ( .A1(n8431), .A2(n8474), .ZN(n8510) );
  OR2_X1 U9684 ( .A1(n5032), .A2(n8510), .ZN(n8433) );
  INV_X1 U9685 ( .A(n10135), .ZN(n8484) );
  OAI22_X1 U9686 ( .A1(n9314), .A2(n8484), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8437), .ZN(n8438) );
  AOI21_X1 U9687 ( .B1(n9318), .B2(n10102), .A(n8438), .ZN(n8439) );
  OAI21_X1 U9688 ( .B1(n9315), .B2(n10093), .A(n8439), .ZN(n8440) );
  AOI21_X1 U9689 ( .B1(n10333), .B2(n9292), .A(n8440), .ZN(n8441) );
  OAI21_X1 U9690 ( .B1(n8442), .B2(n9309), .A(n8441), .ZN(P1_U3212) );
  INV_X1 U9691 ( .A(n10328), .ZN(n8512) );
  OR2_X1 U9692 ( .A1(n10398), .A2(n10007), .ZN(n8444) );
  NOR2_X1 U9693 ( .A1(n10316), .A2(n10293), .ZN(n8446) );
  INV_X1 U9694 ( .A(n10316), .ZN(n11022) );
  NAND2_X1 U9695 ( .A1(n10393), .A2(n10304), .ZN(n9547) );
  NAND2_X1 U9696 ( .A1(n9546), .A2(n9547), .ZN(n10292) );
  NAND2_X1 U9697 ( .A1(n10393), .A2(n10276), .ZN(n8447) );
  NAND2_X1 U9698 ( .A1(n10389), .A2(n10250), .ZN(n9552) );
  NAND2_X1 U9699 ( .A1(n9551), .A2(n9552), .ZN(n10274) );
  OR2_X1 U9700 ( .A1(n10383), .A2(n10277), .ZN(n8448) );
  NAND2_X1 U9701 ( .A1(n10383), .A2(n10277), .ZN(n8449) );
  NAND2_X1 U9702 ( .A1(n10378), .A2(n10251), .ZN(n9560) );
  NAND2_X1 U9703 ( .A1(n9561), .A2(n9560), .ZN(n10241) );
  NAND2_X1 U9704 ( .A1(n10378), .A2(n10223), .ZN(n8450) );
  AND2_X1 U9705 ( .A1(n10374), .A2(n10243), .ZN(n8451) );
  OR2_X1 U9706 ( .A1(n10374), .A2(n10243), .ZN(n8452) );
  INV_X1 U9707 ( .A(n10224), .ZN(n9208) );
  OR2_X1 U9708 ( .A1(n10368), .A2(n9208), .ZN(n9368) );
  NAND2_X1 U9709 ( .A1(n10368), .A2(n9208), .ZN(n9359) );
  NAND2_X1 U9710 ( .A1(n9368), .A2(n9359), .ZN(n9444) );
  NAND2_X1 U9711 ( .A1(n10207), .A2(n9444), .ZN(n8454) );
  OR2_X1 U9712 ( .A1(n10368), .A2(n10224), .ZN(n8453) );
  OR2_X1 U9713 ( .A1(n10364), .A2(n10205), .ZN(n9369) );
  NAND2_X1 U9714 ( .A1(n10364), .A2(n10205), .ZN(n9484) );
  INV_X1 U9715 ( .A(n10205), .ZN(n10179) );
  NAND2_X1 U9716 ( .A1(n10364), .A2(n10179), .ZN(n8455) );
  OR2_X1 U9717 ( .A1(n10358), .A2(n10192), .ZN(n8456) );
  OR2_X1 U9718 ( .A1(n10353), .A2(n8457), .ZN(n9480) );
  NAND2_X1 U9719 ( .A1(n10353), .A2(n8457), .ZN(n9481) );
  OR2_X1 U9720 ( .A1(n10353), .A2(n10180), .ZN(n8458) );
  NAND2_X1 U9721 ( .A1(n10349), .A2(n10164), .ZN(n8459) );
  OR2_X1 U9722 ( .A1(n10349), .A2(n10164), .ZN(n8460) );
  OR2_X1 U9723 ( .A1(n10343), .A2(n10110), .ZN(n9476) );
  NAND2_X1 U9724 ( .A1(n10343), .A2(n10110), .ZN(n9477) );
  NAND2_X1 U9725 ( .A1(n9476), .A2(n9477), .ZN(n8483) );
  OR2_X1 U9726 ( .A1(n10343), .A2(n10144), .ZN(n8461) );
  NOR2_X1 U9727 ( .A1(n10338), .A2(n10135), .ZN(n8463) );
  NAND2_X1 U9728 ( .A1(n10338), .A2(n10135), .ZN(n8464) );
  NAND2_X1 U9729 ( .A1(n10333), .A2(n10111), .ZN(n9474) );
  OR2_X1 U9730 ( .A1(n10333), .A2(n9610), .ZN(n8465) );
  NAND2_X1 U9731 ( .A1(n10328), .A2(n9188), .ZN(n9466) );
  NAND2_X1 U9732 ( .A1(n8466), .A2(n9447), .ZN(n8502) );
  NAND2_X1 U9733 ( .A1(n7712), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8471) );
  NAND2_X1 U9734 ( .A1(n7753), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8470) );
  INV_X1 U9735 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n8467) );
  OR2_X1 U9736 ( .A1(n5034), .A2(n8467), .ZN(n8469) );
  OR2_X1 U9737 ( .A1(n8432), .A2(n8474), .ZN(n8468) );
  NAND2_X1 U9738 ( .A1(n10323), .A2(n9467), .ZN(n9422) );
  AOI21_X1 U9739 ( .B1(n10323), .B2(n8473), .A(n8472), .ZN(n10324) );
  INV_X1 U9740 ( .A(n10323), .ZN(n9464) );
  INV_X1 U9741 ( .A(n8474), .ZN(n8475) );
  AOI22_X1 U9742 ( .A1(n10296), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8475), .B2(
        n10724), .ZN(n8476) );
  OAI21_X1 U9743 ( .B1(n9464), .B2(n10935), .A(n8476), .ZN(n8494) );
  INV_X1 U9744 ( .A(n9523), .ZN(n8477) );
  NAND2_X1 U9745 ( .A1(n10316), .A2(n9533), .ZN(n9524) );
  INV_X1 U9746 ( .A(n10274), .ZN(n9549) );
  INV_X1 U9747 ( .A(n9551), .ZN(n9335) );
  INV_X1 U9748 ( .A(n10277), .ZN(n8479) );
  NAND2_X1 U9749 ( .A1(n10383), .A2(n8479), .ZN(n9556) );
  NAND2_X1 U9750 ( .A1(n9555), .A2(n9556), .ZN(n10252) );
  OAI21_X1 U9751 ( .B1(n10249), .B2(n10252), .A(n9555), .ZN(n10242) );
  INV_X1 U9752 ( .A(n10241), .ZN(n9558) );
  INV_X1 U9753 ( .A(n9561), .ZN(n8480) );
  AOI21_X1 U9754 ( .B1(n10242), .B2(n9558), .A(n8480), .ZN(n10221) );
  OR2_X1 U9755 ( .A1(n10374), .A2(n10204), .ZN(n9565) );
  NAND2_X1 U9756 ( .A1(n10374), .A2(n10204), .ZN(n9566) );
  NAND2_X1 U9757 ( .A1(n10221), .A2(n10222), .ZN(n10220) );
  NAND2_X1 U9758 ( .A1(n10220), .A2(n9566), .ZN(n10203) );
  INV_X1 U9759 ( .A(n10192), .ZN(n8481) );
  OR2_X1 U9760 ( .A1(n10358), .A2(n8481), .ZN(n9482) );
  NAND2_X1 U9761 ( .A1(n10358), .A2(n8481), .ZN(n9483) );
  NAND2_X1 U9762 ( .A1(n10177), .A2(n10178), .ZN(n10176) );
  NAND2_X1 U9763 ( .A1(n10176), .A2(n9483), .ZN(n10162) );
  OR2_X1 U9764 ( .A1(n10349), .A2(n8482), .ZN(n9479) );
  NAND2_X1 U9765 ( .A1(n10349), .A2(n8482), .ZN(n9478) );
  NAND2_X1 U9766 ( .A1(n10133), .A2(n10134), .ZN(n10132) );
  NAND2_X1 U9767 ( .A1(n10132), .A2(n9477), .ZN(n10109) );
  OR2_X1 U9768 ( .A1(n10338), .A2(n8484), .ZN(n9475) );
  NAND2_X1 U9769 ( .A1(n10338), .A2(n8484), .ZN(n10097) );
  INV_X1 U9770 ( .A(n10097), .ZN(n9385) );
  XOR2_X1 U9771 ( .A(n9582), .B(n8485), .Z(n8486) );
  INV_X1 U9772 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U9773 ( .A1(n7239), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U9774 ( .A1(n5035), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8487) );
  OAI211_X1 U9775 ( .C1(n5034), .C2(n8489), .A(n8488), .B(n8487), .ZN(n9608)
         );
  AND2_X1 U9776 ( .A1(n9608), .A2(n8490), .ZN(n8491) );
  AOI21_X1 U9777 ( .B1(n10102), .B2(n10843), .A(n8491), .ZN(n8492) );
  INV_X1 U9778 ( .A(n8495), .ZN(n10449) );
  OAI222_X1 U9779 ( .A1(n9147), .A2(n10449), .B1(n6253), .B2(P2_U3152), .C1(
        n8496), .C2(n9146), .ZN(P2_U3330) );
  INV_X1 U9780 ( .A(n8497), .ZN(n8517) );
  OAI222_X1 U9781 ( .A1(n9147), .A2(n8517), .B1(n8499), .B2(P2_U3152), .C1(
        n8498), .C2(n9146), .ZN(P2_U3328) );
  NAND2_X1 U9782 ( .A1(n8500), .A2(n9581), .ZN(n8501) );
  NAND2_X1 U9783 ( .A1(n8502), .A2(n8501), .ZN(n10332) );
  OAI21_X1 U9784 ( .B1(n9581), .B2(n8504), .A(n8503), .ZN(n8506) );
  OAI22_X1 U9785 ( .A1(n10111), .A2(n10915), .B1(n9467), .B2(n10917), .ZN(
        n8505) );
  AOI21_X1 U9786 ( .B1(n10328), .B2(n10090), .A(n8509), .ZN(n10329) );
  INV_X1 U9787 ( .A(n8510), .ZN(n9193) );
  AOI22_X1 U9788 ( .A1(n10296), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9193), .B2(
        n10724), .ZN(n8511) );
  OAI21_X1 U9789 ( .B1(n8512), .B2(n10935), .A(n8511), .ZN(n8514) );
  NOR2_X1 U9790 ( .A1(n10332), .A2(n10264), .ZN(n8513) );
  AOI211_X1 U9791 ( .C1(n10932), .C2(n10329), .A(n8514), .B(n8513), .ZN(n8515)
         );
  OAI21_X1 U9792 ( .B1(n10331), .B2(n10296), .A(n8515), .ZN(P1_U3263) );
  OAI222_X1 U9793 ( .A1(P1_U3084), .A2(n8518), .B1(n10461), .B2(n8517), .C1(
        n8516), .C2(n10454), .ZN(P1_U3323) );
  XNOR2_X1 U9794 ( .A(n8519), .B(n8520), .ZN(n8526) );
  NOR2_X1 U9795 ( .A1(n10968), .A2(n8521), .ZN(n8524) );
  AOI22_X1 U9796 ( .A1(n10884), .A2(n8654), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8522) );
  OAI21_X1 U9797 ( .B1(n8824), .B2(n10886), .A(n8522), .ZN(n8523) );
  AOI211_X1 U9798 ( .C1(n9046), .C2(n10963), .A(n8524), .B(n8523), .ZN(n8525)
         );
  OAI21_X1 U9799 ( .B1(n8526), .B2(n10890), .A(n8525), .ZN(P2_U3216) );
  NAND2_X1 U9800 ( .A1(n8612), .A2(n8527), .ZN(n8531) );
  XNOR2_X1 U9801 ( .A(n8529), .B(n8528), .ZN(n8530) );
  XNOR2_X1 U9802 ( .A(n8531), .B(n8530), .ZN(n8537) );
  NAND2_X1 U9803 ( .A1(n6450), .A2(n8886), .ZN(n8533) );
  AOI22_X1 U9804 ( .A1(n10884), .A2(n8880), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8532) );
  OAI211_X1 U9805 ( .C1(n8534), .C2(n10886), .A(n8533), .B(n8532), .ZN(n8535)
         );
  AOI21_X1 U9806 ( .B1(n9068), .B2(n10963), .A(n8535), .ZN(n8536) );
  OAI21_X1 U9807 ( .B1(n8537), .B2(n10890), .A(n8536), .ZN(P2_U3218) );
  AOI21_X1 U9808 ( .B1(n8539), .B2(n8538), .A(n10890), .ZN(n8541) );
  NAND2_X1 U9809 ( .A1(n8541), .A2(n8540), .ZN(n8547) );
  INV_X1 U9810 ( .A(n10886), .ZN(n8543) );
  AOI22_X1 U9811 ( .A1(n8543), .A2(n5815), .B1(n10884), .B2(n8542), .ZN(n8546)
         );
  MUX2_X1 U9812 ( .A(n10968), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n8545) );
  NAND2_X1 U9813 ( .A1(n10963), .A2(n10766), .ZN(n8544) );
  NAND4_X1 U9814 ( .A1(n8547), .A2(n8546), .A3(n8545), .A4(n8544), .ZN(
        P2_U3220) );
  XNOR2_X1 U9815 ( .A(n8549), .B(n8548), .ZN(n8556) );
  NOR2_X1 U9816 ( .A1(n10968), .A2(n8951), .ZN(n8554) );
  NAND2_X1 U9817 ( .A1(n8919), .A2(n9016), .ZN(n8551) );
  OR2_X1 U9818 ( .A1(n8591), .A2(n10792), .ZN(n8550) );
  AND2_X1 U9819 ( .A1(n8551), .A2(n8550), .ZN(n8948) );
  NAND2_X1 U9820 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8772) );
  OAI21_X1 U9821 ( .B1(n8948), .B2(n8552), .A(n8772), .ZN(n8553) );
  AOI211_X1 U9822 ( .C1(n9091), .C2(n10963), .A(n8554), .B(n8553), .ZN(n8555)
         );
  OAI21_X1 U9823 ( .B1(n8556), .B2(n10890), .A(n8555), .ZN(P2_U3221) );
  XNOR2_X1 U9824 ( .A(n8558), .B(n8557), .ZN(n8564) );
  NAND2_X1 U9825 ( .A1(n6450), .A2(n8912), .ZN(n8560) );
  AOI22_X1 U9826 ( .A1(n10884), .A2(n8918), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8559) );
  OAI211_X1 U9827 ( .C1(n8561), .C2(n10886), .A(n8560), .B(n8559), .ZN(n8562)
         );
  AOI21_X1 U9828 ( .B1(n9079), .B2(n10963), .A(n8562), .ZN(n8563) );
  OAI21_X1 U9829 ( .B1(n8564), .B2(n10890), .A(n8563), .ZN(P2_U3225) );
  XNOR2_X1 U9830 ( .A(n8566), .B(n8565), .ZN(n8573) );
  INV_X1 U9831 ( .A(n8849), .ZN(n8570) );
  OR2_X1 U9832 ( .A1(n8824), .A2(n10794), .ZN(n8567) );
  OAI21_X1 U9833 ( .B1(n8568), .B2(n10792), .A(n8567), .ZN(n8853) );
  AOI22_X1 U9834 ( .A1(n8853), .A2(n10955), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8569) );
  OAI21_X1 U9835 ( .B1(n10968), .B2(n8570), .A(n8569), .ZN(n8571) );
  AOI21_X1 U9836 ( .B1(n9057), .B2(n10963), .A(n8571), .ZN(n8572) );
  OAI21_X1 U9837 ( .B1(n8573), .B2(n10890), .A(n8572), .ZN(P2_U3227) );
  INV_X1 U9838 ( .A(n9105), .ZN(n8584) );
  OAI21_X1 U9839 ( .B1(n8576), .B2(n8575), .A(n8574), .ZN(n8577) );
  NAND2_X1 U9840 ( .A1(n8577), .A2(n10964), .ZN(n8583) );
  OAI22_X1 U9841 ( .A1(n8627), .A2(n10794), .B1(n8578), .B2(n10792), .ZN(n8997) );
  NOR2_X1 U9842 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8579), .ZN(n8720) );
  INV_X1 U9843 ( .A(n9002), .ZN(n8580) );
  NOR2_X1 U9844 ( .A1(n10968), .A2(n8580), .ZN(n8581) );
  AOI211_X1 U9845 ( .C1(n10955), .C2(n8997), .A(n8720), .B(n8581), .ZN(n8582)
         );
  OAI211_X1 U9846 ( .C1(n8584), .C2(n6439), .A(n8583), .B(n8582), .ZN(P2_U3228) );
  NAND2_X1 U9847 ( .A1(n6376), .A2(n8586), .ZN(n8587) );
  XNOR2_X1 U9848 ( .A(n8588), .B(n8587), .ZN(n8595) );
  INV_X1 U9849 ( .A(n8589), .ZN(n8988) );
  OAI22_X1 U9850 ( .A1(n8591), .A2(n10794), .B1(n8590), .B2(n10792), .ZN(n8980) );
  AOI22_X1 U9851 ( .A1(n8980), .A2(n10955), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8592) );
  OAI21_X1 U9852 ( .B1(n8988), .B2(n10968), .A(n8592), .ZN(n8593) );
  AOI21_X1 U9853 ( .B1(n9100), .B2(n10963), .A(n8593), .ZN(n8594) );
  OAI21_X1 U9854 ( .B1(n8595), .B2(n10890), .A(n8594), .ZN(P2_U3230) );
  XNOR2_X1 U9855 ( .A(n8597), .B(n8596), .ZN(n8602) );
  NOR2_X1 U9856 ( .A1(n10886), .A2(n8860), .ZN(n8599) );
  OAI22_X1 U9857 ( .A1(n8606), .A2(n8861), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9711), .ZN(n8598) );
  AOI211_X1 U9858 ( .C1(n6450), .C2(n8868), .A(n8599), .B(n8598), .ZN(n8601)
         );
  NAND2_X1 U9859 ( .A1(n9062), .A2(n10963), .ZN(n8600) );
  OAI211_X1 U9860 ( .C1(n8602), .C2(n10890), .A(n8601), .B(n8600), .ZN(
        P2_U3231) );
  XNOR2_X1 U9861 ( .A(n8604), .B(n8603), .ZN(n8611) );
  INV_X1 U9862 ( .A(n8605), .ZN(n8929) );
  NOR2_X1 U9863 ( .A1(n10886), .A2(n8935), .ZN(n8608) );
  INV_X1 U9864 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9715) );
  OAI22_X1 U9865 ( .A1(n8606), .A2(n8934), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9715), .ZN(n8607) );
  AOI211_X1 U9866 ( .C1(n6450), .C2(n8929), .A(n8608), .B(n8607), .ZN(n8610)
         );
  NAND2_X1 U9867 ( .A1(n9084), .A2(n10963), .ZN(n8609) );
  OAI211_X1 U9868 ( .C1(n8611), .C2(n10890), .A(n8610), .B(n8609), .ZN(
        P2_U3235) );
  INV_X1 U9869 ( .A(n8612), .ZN(n8613) );
  AOI21_X1 U9870 ( .B1(n8615), .B2(n8614), .A(n8613), .ZN(n8621) );
  INV_X1 U9871 ( .A(n8904), .ZN(n8618) );
  OR2_X1 U9872 ( .A1(n8860), .A2(n10794), .ZN(n8616) );
  OAI21_X1 U9873 ( .B1(n8934), .B2(n10792), .A(n8616), .ZN(n8902) );
  AOI22_X1 U9874 ( .A1(n8902), .A2(n10955), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8617) );
  OAI21_X1 U9875 ( .B1(n10968), .B2(n8618), .A(n8617), .ZN(n8619) );
  AOI21_X1 U9876 ( .B1(n9074), .B2(n10963), .A(n8619), .ZN(n8620) );
  OAI21_X1 U9877 ( .B1(n8621), .B2(n10890), .A(n8620), .ZN(P2_U3237) );
  NAND2_X1 U9878 ( .A1(n8623), .A2(n8622), .ZN(n8625) );
  XOR2_X1 U9879 ( .A(n8625), .B(n8624), .Z(n8631) );
  NOR2_X1 U9880 ( .A1(n10968), .A2(n8960), .ZN(n8629) );
  NAND2_X1 U9881 ( .A1(n10884), .A2(n8968), .ZN(n8626) );
  NAND2_X1 U9882 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8742) );
  OAI211_X1 U9883 ( .C1(n8627), .C2(n10886), .A(n8626), .B(n8742), .ZN(n8628)
         );
  AOI211_X1 U9884 ( .C1(n9094), .C2(n10963), .A(n8629), .B(n8628), .ZN(n8630)
         );
  OAI21_X1 U9885 ( .B1(n8631), .B2(n10890), .A(n8630), .ZN(P2_U3240) );
  XNOR2_X1 U9886 ( .A(n8632), .B(n8633), .ZN(n8640) );
  INV_X1 U9887 ( .A(n8840), .ZN(n8637) );
  NAND2_X1 U9888 ( .A1(n8634), .A2(n9016), .ZN(n8635) );
  OAI21_X1 U9889 ( .B1(n8861), .B2(n10792), .A(n8635), .ZN(n8836) );
  AOI22_X1 U9890 ( .A1(n8836), .A2(n10955), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8636) );
  OAI21_X1 U9891 ( .B1(n10968), .B2(n8637), .A(n8636), .ZN(n8638) );
  AOI21_X1 U9892 ( .B1(n9052), .B2(n10963), .A(n8638), .ZN(n8639) );
  OAI21_X1 U9893 ( .B1(n8640), .B2(n10890), .A(n8639), .ZN(P2_U3242) );
  OAI21_X1 U9894 ( .B1(n8643), .B2(n8642), .A(n8641), .ZN(n8644) );
  NAND2_X1 U9895 ( .A1(n8644), .A2(n10964), .ZN(n8650) );
  NAND2_X1 U9896 ( .A1(n10884), .A2(n8657), .ZN(n8645) );
  NAND2_X1 U9897 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8697) );
  OAI211_X1 U9898 ( .C1(n8646), .C2(n10886), .A(n8645), .B(n8697), .ZN(n8647)
         );
  AOI21_X1 U9899 ( .B1(n8648), .B2(n6450), .A(n8647), .ZN(n8649) );
  OAI211_X1 U9900 ( .C1(n8651), .C2(n6439), .A(n8650), .B(n8649), .ZN(P2_U3243) );
  INV_X1 U9901 ( .A(n8652), .ZN(n8778) );
  MUX2_X1 U9902 ( .A(n8778), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8665), .Z(
        P2_U3583) );
  MUX2_X1 U9903 ( .A(n8653), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8665), .Z(
        P2_U3582) );
  MUX2_X1 U9904 ( .A(n8654), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8665), .Z(
        P2_U3580) );
  MUX2_X1 U9905 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8655), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9906 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8880), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9907 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n5536), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9908 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8918), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9909 ( .A(n8919), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8665), .Z(
        P2_U3572) );
  MUX2_X1 U9910 ( .A(n8968), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8665), .Z(
        P2_U3571) );
  MUX2_X1 U9911 ( .A(n8656), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8665), .Z(
        P2_U3570) );
  MUX2_X1 U9912 ( .A(n8657), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8665), .Z(
        P2_U3568) );
  MUX2_X1 U9913 ( .A(n8658), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8665), .Z(
        P2_U3567) );
  MUX2_X1 U9914 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8659), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9915 ( .A(n8660), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8665), .Z(
        P2_U3565) );
  MUX2_X1 U9916 ( .A(n8661), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8665), .Z(
        P2_U3564) );
  MUX2_X1 U9917 ( .A(n8662), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8665), .Z(
        P2_U3563) );
  MUX2_X1 U9918 ( .A(n8663), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8665), .Z(
        P2_U3562) );
  MUX2_X1 U9919 ( .A(n10883), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8665), .Z(
        P2_U3560) );
  MUX2_X1 U9920 ( .A(n9017), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8665), .Z(
        P2_U3559) );
  MUX2_X1 U9921 ( .A(n8664), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8665), .Z(
        P2_U3558) );
  MUX2_X1 U9922 ( .A(n9015), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8665), .Z(
        P2_U3557) );
  MUX2_X1 U9923 ( .A(n6230), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8665), .Z(
        P2_U3552) );
  NOR2_X1 U9924 ( .A1(n10638), .A2(n8666), .ZN(n8667) );
  AOI211_X1 U9925 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n10647), .A(n8668), .B(
        n8667), .ZN(n8678) );
  NAND2_X1 U9926 ( .A1(n8670), .A2(n8669), .ZN(n8671) );
  NAND3_X1 U9927 ( .A1(n10622), .A2(n8672), .A3(n8671), .ZN(n8677) );
  OAI211_X1 U9928 ( .C1(n8675), .C2(n8674), .A(n10656), .B(n8673), .ZN(n8676)
         );
  NAND3_X1 U9929 ( .A1(n8678), .A2(n8677), .A3(n8676), .ZN(P2_U3253) );
  OAI211_X1 U9930 ( .C1(n8681), .C2(n8680), .A(n10656), .B(n8679), .ZN(n8691)
         );
  NOR2_X1 U9931 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8682), .ZN(n8683) );
  AOI21_X1 U9932 ( .B1(n10647), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8683), .ZN(
        n8690) );
  OAI211_X1 U9933 ( .C1(n8686), .C2(n8685), .A(n10622), .B(n8684), .ZN(n8689)
         );
  NAND2_X1 U9934 ( .A1(n10654), .A2(n8687), .ZN(n8688) );
  NAND4_X1 U9935 ( .A1(n8691), .A2(n8690), .A3(n8689), .A4(n8688), .ZN(
        P2_U3254) );
  OAI21_X1 U9936 ( .B1(n8693), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8692), .ZN(
        n8705) );
  XNOR2_X1 U9937 ( .A(n8714), .B(n8705), .ZN(n8695) );
  INV_X1 U9938 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U9939 ( .A1(n8695), .A2(n8694), .ZN(n8707) );
  OAI21_X1 U9940 ( .B1(n8695), .B2(n8694), .A(n8707), .ZN(n8696) );
  AOI22_X1 U9941 ( .A1(n8714), .A2(n10654), .B1(n10622), .B2(n8696), .ZN(n8704) );
  INV_X1 U9942 ( .A(n8697), .ZN(n8698) );
  AOI21_X1 U9943 ( .B1(n10647), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8698), .ZN(
        n8703) );
  AOI21_X1 U9944 ( .B1(n8700), .B2(n7305), .A(n8699), .ZN(n8713) );
  XNOR2_X1 U9945 ( .A(n8706), .B(n8713), .ZN(n8701) );
  NAND2_X1 U9946 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n8701), .ZN(n8715) );
  OAI211_X1 U9947 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n8701), .A(n10656), .B(
        n8715), .ZN(n8702) );
  NAND3_X1 U9948 ( .A1(n8704), .A2(n8703), .A3(n8702), .ZN(P2_U3260) );
  NAND2_X1 U9949 ( .A1(n8706), .A2(n8705), .ZN(n8708) );
  NAND2_X1 U9950 ( .A1(n8708), .A2(n8707), .ZN(n8712) );
  INV_X1 U9951 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8709) );
  MUX2_X1 U9952 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n8709), .S(n8726), .Z(n8710)
         );
  INV_X1 U9953 ( .A(n8710), .ZN(n8711) );
  NOR2_X1 U9954 ( .A1(n8712), .A2(n8711), .ZN(n8725) );
  AOI211_X1 U9955 ( .C1(n8712), .C2(n8711), .A(n8725), .B(n10648), .ZN(n8724)
         );
  NAND2_X1 U9956 ( .A1(n8714), .A2(n8713), .ZN(n8716) );
  NAND2_X1 U9957 ( .A1(n8716), .A2(n8715), .ZN(n8718) );
  XNOR2_X1 U9958 ( .A(n8726), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8717) );
  NOR2_X1 U9959 ( .A1(n8718), .A2(n8717), .ZN(n8731) );
  AOI21_X1 U9960 ( .B1(n8718), .B2(n8717), .A(n8731), .ZN(n8719) );
  NOR2_X1 U9961 ( .A1(n8719), .A2(n10624), .ZN(n8723) );
  AOI21_X1 U9962 ( .B1(n10647), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8720), .ZN(
        n8721) );
  OAI21_X1 U9963 ( .B1(n10638), .B2(n8733), .A(n8721), .ZN(n8722) );
  OR3_X1 U9964 ( .A1(n8724), .A2(n8723), .A3(n8722), .ZN(P2_U3261) );
  AOI21_X1 U9965 ( .B1(n8726), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8725), .ZN(
        n8730) );
  INV_X1 U9966 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8727) );
  MUX2_X1 U9967 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n8727), .S(n8753), .Z(n8728)
         );
  INV_X1 U9968 ( .A(n8728), .ZN(n8729) );
  NOR2_X1 U9969 ( .A1(n8730), .A2(n8729), .ZN(n8752) );
  AOI211_X1 U9970 ( .C1(n8730), .C2(n8729), .A(n8752), .B(n10648), .ZN(n8741)
         );
  INV_X1 U9971 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8732) );
  AOI21_X1 U9972 ( .B1(n8733), .B2(n8732), .A(n8731), .ZN(n8735) );
  XNOR2_X1 U9973 ( .A(n8744), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U9974 ( .A1(n8734), .A2(n8735), .ZN(n8743) );
  OAI211_X1 U9975 ( .C1(n8735), .C2(n8734), .A(n10656), .B(n8743), .ZN(n8739)
         );
  NOR2_X1 U9976 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8736), .ZN(n8737) );
  AOI21_X1 U9977 ( .B1(n10647), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8737), .ZN(
        n8738) );
  OAI211_X1 U9978 ( .C1(n10638), .C2(n8744), .A(n8739), .B(n8738), .ZN(n8740)
         );
  OR2_X1 U9979 ( .A1(n8741), .A2(n8740), .ZN(P2_U3262) );
  INV_X1 U9980 ( .A(n8742), .ZN(n8751) );
  INV_X1 U9981 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8745) );
  OAI21_X1 U9982 ( .B1(n8745), .B2(n8744), .A(n8743), .ZN(n8748) );
  INV_X1 U9983 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U9984 ( .A1(n8760), .A2(n8746), .ZN(n8766) );
  OAI21_X1 U9985 ( .B1(n8760), .B2(n8746), .A(n8766), .ZN(n8747) );
  NOR2_X1 U9986 ( .A1(n8747), .A2(n8748), .ZN(n8768) );
  AOI21_X1 U9987 ( .B1(n8748), .B2(n8747), .A(n8768), .ZN(n8749) );
  NOR2_X1 U9988 ( .A1(n8749), .A2(n10624), .ZN(n8750) );
  AOI211_X1 U9989 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n10647), .A(n8751), .B(
        n8750), .ZN(n8759) );
  AOI21_X1 U9990 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n8753), .A(n8752), .ZN(
        n8756) );
  INV_X1 U9991 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8754) );
  MUX2_X1 U9992 ( .A(P2_REG2_REG_18__SCAN_IN), .B(n8754), .S(n8762), .Z(n8755)
         );
  NAND2_X1 U9993 ( .A1(n8755), .A2(n8756), .ZN(n8761) );
  OAI21_X1 U9994 ( .B1(n8756), .B2(n8755), .A(n8761), .ZN(n8757) );
  NAND2_X1 U9995 ( .A1(n10622), .A2(n8757), .ZN(n8758) );
  OAI211_X1 U9996 ( .C1(n10638), .C2(n8760), .A(n8759), .B(n8758), .ZN(
        P2_U3263) );
  OAI21_X1 U9997 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8762), .A(n8761), .ZN(
        n8765) );
  INV_X1 U9998 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8763) );
  MUX2_X1 U9999 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8763), .S(n6223), .Z(n8764)
         );
  XNOR2_X1 U10000 ( .A(n8765), .B(n8764), .ZN(n8776) );
  INV_X1 U10001 ( .A(n8766), .ZN(n8767) );
  NOR2_X1 U10002 ( .A1(n8768), .A2(n8767), .ZN(n8770) );
  XNOR2_X1 U10003 ( .A(n6223), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8769) );
  XNOR2_X1 U10004 ( .A(n8770), .B(n8769), .ZN(n8773) );
  NAND2_X1 U10005 ( .A1(n10647), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8771) );
  OAI211_X1 U10006 ( .C1(n8773), .C2(n10624), .A(n8772), .B(n8771), .ZN(n8774)
         );
  AOI21_X1 U10007 ( .B1(n10815), .B2(n10654), .A(n8774), .ZN(n8775) );
  OAI21_X1 U10008 ( .B1(n8776), .B2(n10648), .A(n8775), .ZN(P2_U3264) );
  NAND2_X1 U10009 ( .A1(n8778), .A2(n8777), .ZN(n9036) );
  NOR2_X1 U10010 ( .A1(n10821), .A2(n9036), .ZN(n8786) );
  AOI21_X1 U10011 ( .B1(n10821), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8786), .ZN(
        n8780) );
  NAND2_X1 U10012 ( .A1(n9032), .A2(n10767), .ZN(n8779) );
  OAI211_X1 U10013 ( .C1(n9034), .C2(n8788), .A(n8780), .B(n8779), .ZN(
        P2_U3265) );
  OR2_X1 U10014 ( .A1(n8784), .A2(n8781), .ZN(n8782) );
  NAND2_X1 U10015 ( .A1(n8783), .A2(n8782), .ZN(n9035) );
  NOR2_X1 U10016 ( .A1(n8784), .A2(n8963), .ZN(n8785) );
  AOI211_X1 U10017 ( .C1(n10821), .C2(P2_REG2_REG_30__SCAN_IN), .A(n8786), .B(
        n8785), .ZN(n8787) );
  OAI21_X1 U10018 ( .B1(n8788), .B2(n9035), .A(n8787), .ZN(P2_U3266) );
  NAND2_X1 U10019 ( .A1(n8789), .A2(n10764), .ZN(n8792) );
  AOI22_X1 U10020 ( .A1(n10821), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8790), 
        .B2(n10813), .ZN(n8791) );
  OAI211_X1 U10021 ( .C1(n8793), .C2(n8963), .A(n8792), .B(n8791), .ZN(n8794)
         );
  AOI21_X1 U10022 ( .B1(n8795), .B2(n9024), .A(n8794), .ZN(n8796) );
  OAI21_X1 U10023 ( .B1(n8797), .B2(n10821), .A(n8796), .ZN(P2_U3267) );
  XNOR2_X1 U10024 ( .A(n8799), .B(n8798), .ZN(n9045) );
  AOI21_X1 U10025 ( .B1(n9041), .B2(n8815), .A(n8800), .ZN(n9042) );
  AOI22_X1 U10026 ( .A1(n10821), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8801), 
        .B2(n10813), .ZN(n8802) );
  OAI21_X1 U10027 ( .B1(n8803), .B2(n8963), .A(n8802), .ZN(n8811) );
  INV_X1 U10028 ( .A(n8804), .ZN(n8806) );
  AOI21_X1 U10029 ( .B1(n8806), .B2(n8805), .A(n8932), .ZN(n8809) );
  AOI21_X1 U10030 ( .B1(n8809), .B2(n8808), .A(n8807), .ZN(n9044) );
  NOR2_X1 U10031 ( .A1(n9044), .A2(n10821), .ZN(n8810) );
  AOI211_X1 U10032 ( .C1(n10764), .C2(n9042), .A(n8811), .B(n8810), .ZN(n8812)
         );
  OAI21_X1 U10033 ( .B1(n9045), .B2(n9008), .A(n8812), .ZN(P2_U3268) );
  XNOR2_X1 U10034 ( .A(n8814), .B(n8813), .ZN(n9050) );
  INV_X1 U10035 ( .A(n8815), .ZN(n8816) );
  AOI21_X1 U10036 ( .B1(n9046), .B2(n8838), .A(n8816), .ZN(n9047) );
  AOI22_X1 U10037 ( .A1(n10821), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8817), 
        .B2(n10813), .ZN(n8818) );
  OAI21_X1 U10038 ( .B1(n8819), .B2(n8963), .A(n8818), .ZN(n8829) );
  INV_X1 U10039 ( .A(n8820), .ZN(n8822) );
  AOI21_X1 U10040 ( .B1(n8822), .B2(n8821), .A(n8932), .ZN(n8827) );
  OAI22_X1 U10041 ( .A1(n8824), .A2(n10792), .B1(n8823), .B2(n10794), .ZN(
        n8825) );
  AOI21_X1 U10042 ( .B1(n8827), .B2(n8826), .A(n8825), .ZN(n9049) );
  NOR2_X1 U10043 ( .A1(n9049), .A2(n10821), .ZN(n8828) );
  AOI211_X1 U10044 ( .C1(n9047), .C2(n10764), .A(n8829), .B(n8828), .ZN(n8830)
         );
  OAI21_X1 U10045 ( .B1(n9050), .B2(n9008), .A(n8830), .ZN(P2_U3269) );
  XOR2_X1 U10046 ( .A(n8835), .B(n8831), .Z(n9055) );
  NOR2_X1 U10047 ( .A1(n8832), .A2(n8963), .ZN(n8843) );
  NAND2_X1 U10048 ( .A1(n8854), .A2(n8833), .ZN(n8834) );
  XOR2_X1 U10049 ( .A(n8835), .B(n8834), .Z(n8837) );
  AOI21_X1 U10050 ( .B1(n8837), .B2(n10808), .A(n8836), .ZN(n9054) );
  INV_X1 U10051 ( .A(n8838), .ZN(n8839) );
  AOI211_X1 U10052 ( .C1(n9052), .C2(n5273), .A(n11030), .B(n8839), .ZN(n9051)
         );
  AOI22_X1 U10053 ( .A1(n9051), .A2(n6223), .B1(n10813), .B2(n8840), .ZN(n8841) );
  AOI21_X1 U10054 ( .B1(n9054), .B2(n8841), .A(n10821), .ZN(n8842) );
  AOI211_X1 U10055 ( .C1(n10821), .C2(P2_REG2_REG_26__SCAN_IN), .A(n8843), .B(
        n8842), .ZN(n8844) );
  OAI21_X1 U10056 ( .B1(n9055), .B2(n9008), .A(n8844), .ZN(P2_U3270) );
  XNOR2_X1 U10057 ( .A(n8846), .B(n8845), .ZN(n9060) );
  AOI211_X1 U10058 ( .C1(n9057), .C2(n8848), .A(n11030), .B(n8847), .ZN(n9056)
         );
  AOI22_X1 U10059 ( .A1(n10821), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8849), 
        .B2(n10813), .ZN(n8850) );
  OAI21_X1 U10060 ( .B1(n8851), .B2(n8963), .A(n8850), .ZN(n8857) );
  AOI21_X1 U10061 ( .B1(n5065), .B2(n8852), .A(n8932), .ZN(n8855) );
  AOI21_X1 U10062 ( .B1(n8855), .B2(n8854), .A(n8853), .ZN(n9059) );
  NOR2_X1 U10063 ( .A1(n9059), .A2(n10821), .ZN(n8856) );
  AOI211_X1 U10064 ( .C1(n9056), .C2(n9011), .A(n8857), .B(n8856), .ZN(n8858)
         );
  OAI21_X1 U10065 ( .B1(n9060), .B2(n9008), .A(n8858), .ZN(P2_U3271) );
  AOI21_X1 U10066 ( .B1(n8859), .B2(n8866), .A(n8932), .ZN(n8864) );
  OAI22_X1 U10067 ( .A1(n8861), .A2(n10794), .B1(n8860), .B2(n10792), .ZN(
        n8862) );
  AOI21_X1 U10068 ( .B1(n8864), .B2(n8863), .A(n8862), .ZN(n9065) );
  OAI21_X1 U10069 ( .B1(n8867), .B2(n8866), .A(n8865), .ZN(n9061) );
  NAND2_X1 U10070 ( .A1(n9061), .A2(n9024), .ZN(n8874) );
  XNOR2_X1 U10071 ( .A(n8885), .B(n9062), .ZN(n9063) );
  INV_X1 U10072 ( .A(n8868), .ZN(n8871) );
  NAND2_X1 U10073 ( .A1(n9062), .A2(n10767), .ZN(n8870) );
  NAND2_X1 U10074 ( .A1(n10821), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8869) );
  OAI211_X1 U10075 ( .C1(n8987), .C2(n8871), .A(n8870), .B(n8869), .ZN(n8872)
         );
  AOI21_X1 U10076 ( .B1(n9063), .B2(n10764), .A(n8872), .ZN(n8873) );
  OAI211_X1 U10077 ( .C1(n10821), .C2(n9065), .A(n8874), .B(n8873), .ZN(
        P2_U3272) );
  INV_X1 U10078 ( .A(n8875), .ZN(n8900) );
  OAI21_X1 U10079 ( .B1(n8900), .B2(n8877), .A(n8876), .ZN(n8879) );
  NAND2_X1 U10080 ( .A1(n8879), .A2(n8878), .ZN(n8881) );
  AOI222_X1 U10081 ( .A1(n10808), .A2(n8881), .B1(n8880), .B2(n9016), .C1(
        n8918), .C2(n9014), .ZN(n9071) );
  NAND2_X1 U10082 ( .A1(n8883), .A2(n8882), .ZN(n9067) );
  NAND3_X1 U10083 ( .A1(n5477), .A2(n9024), .A3(n9067), .ZN(n8891) );
  AND2_X1 U10084 ( .A1(n9068), .A2(n8894), .ZN(n8884) );
  NOR2_X1 U10085 ( .A1(n8885), .A2(n8884), .ZN(n9069) );
  INV_X1 U10086 ( .A(n9068), .ZN(n8888) );
  AOI22_X1 U10087 ( .A1(n10821), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8886), 
        .B2(n10813), .ZN(n8887) );
  OAI21_X1 U10088 ( .B1(n8888), .B2(n8963), .A(n8887), .ZN(n8889) );
  AOI21_X1 U10089 ( .B1(n9069), .B2(n10764), .A(n8889), .ZN(n8890) );
  OAI211_X1 U10090 ( .C1(n10821), .C2(n9071), .A(n8891), .B(n8890), .ZN(
        P2_U3273) );
  XOR2_X1 U10091 ( .A(n8899), .B(n8892), .Z(n9078) );
  INV_X1 U10092 ( .A(n8894), .ZN(n8895) );
  AOI21_X1 U10093 ( .B1(n9074), .B2(n8911), .A(n8895), .ZN(n9075) );
  INV_X1 U10094 ( .A(n9074), .ZN(n8897) );
  INV_X1 U10095 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8896) );
  OAI22_X1 U10096 ( .A1(n8897), .A2(n8963), .B1(n10818), .B2(n8896), .ZN(n8907) );
  INV_X1 U10097 ( .A(n8898), .ZN(n8901) );
  AOI211_X1 U10098 ( .C1(n8901), .C2(n5585), .A(n8932), .B(n8900), .ZN(n8903)
         );
  NOR2_X1 U10099 ( .A1(n8903), .A2(n8902), .ZN(n9077) );
  NAND2_X1 U10100 ( .A1(n10813), .A2(n8904), .ZN(n8905) );
  AOI21_X1 U10101 ( .B1(n9077), .B2(n8905), .A(n10821), .ZN(n8906) );
  AOI211_X1 U10102 ( .C1(n9075), .C2(n10764), .A(n8907), .B(n8906), .ZN(n8908)
         );
  OAI21_X1 U10103 ( .B1(n9078), .B2(n9008), .A(n8908), .ZN(P2_U3274) );
  AOI21_X1 U10104 ( .B1(n8916), .B2(n8910), .A(n8909), .ZN(n9083) );
  AOI21_X1 U10105 ( .B1(n9079), .B2(n8927), .A(n8893), .ZN(n9080) );
  AOI22_X1 U10106 ( .A1(n10821), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8912), 
        .B2(n10813), .ZN(n8913) );
  OAI21_X1 U10107 ( .B1(n8914), .B2(n8963), .A(n8913), .ZN(n8923) );
  OAI211_X1 U10108 ( .C1(n8917), .C2(n8916), .A(n8915), .B(n10808), .ZN(n8921)
         );
  AOI22_X1 U10109 ( .A1(n8919), .A2(n9014), .B1(n8918), .B2(n9016), .ZN(n8920)
         );
  AND2_X1 U10110 ( .A1(n8921), .A2(n8920), .ZN(n9082) );
  NOR2_X1 U10111 ( .A1(n9082), .A2(n10821), .ZN(n8922) );
  AOI211_X1 U10112 ( .C1(n9080), .C2(n10764), .A(n8923), .B(n8922), .ZN(n8924)
         );
  OAI21_X1 U10113 ( .B1(n9083), .B2(n9008), .A(n8924), .ZN(P2_U3275) );
  OAI21_X1 U10114 ( .B1(n8926), .B2(n8933), .A(n8925), .ZN(n9088) );
  INV_X1 U10115 ( .A(n8927), .ZN(n8928) );
  AOI21_X1 U10116 ( .B1(n9084), .B2(n5275), .A(n8928), .ZN(n9085) );
  AOI22_X1 U10117 ( .A1(n10821), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8929), 
        .B2(n10813), .ZN(n8930) );
  OAI21_X1 U10118 ( .B1(n8931), .B2(n8963), .A(n8930), .ZN(n8940) );
  AOI21_X1 U10119 ( .B1(n5093), .B2(n8933), .A(n8932), .ZN(n8938) );
  OAI22_X1 U10120 ( .A1(n8935), .A2(n10792), .B1(n8934), .B2(n10794), .ZN(
        n8936) );
  AOI21_X1 U10121 ( .B1(n8938), .B2(n8937), .A(n8936), .ZN(n9087) );
  NOR2_X1 U10122 ( .A1(n9087), .A2(n10821), .ZN(n8939) );
  AOI211_X1 U10123 ( .C1(n9085), .C2(n10764), .A(n8940), .B(n8939), .ZN(n8941)
         );
  OAI21_X1 U10124 ( .B1(n9008), .B2(n9088), .A(n8941), .ZN(P2_U3276) );
  OAI21_X1 U10125 ( .B1(n8944), .B2(n8943), .A(n8942), .ZN(n9093) );
  AOI22_X1 U10126 ( .A1(n9091), .A2(n10767), .B1(P2_REG2_REG_19__SCAN_IN), 
        .B2(n10821), .ZN(n8955) );
  OAI211_X1 U10127 ( .C1(n8947), .C2(n8946), .A(n8945), .B(n10808), .ZN(n8949)
         );
  NAND2_X1 U10128 ( .A1(n8949), .A2(n8948), .ZN(n9089) );
  AOI211_X1 U10129 ( .C1(n9091), .C2(n8957), .A(n11030), .B(n8950), .ZN(n9090)
         );
  INV_X1 U10130 ( .A(n9090), .ZN(n8952) );
  OAI22_X1 U10131 ( .A1(n8952), .A2(n10815), .B1(n8987), .B2(n8951), .ZN(n8953) );
  OAI21_X1 U10132 ( .B1(n9089), .B2(n8953), .A(n10818), .ZN(n8954) );
  OAI211_X1 U10133 ( .C1(n9093), .C2(n9008), .A(n8955), .B(n8954), .ZN(
        P2_U3277) );
  XNOR2_X1 U10134 ( .A(n8956), .B(n8966), .ZN(n9098) );
  INV_X1 U10135 ( .A(n8957), .ZN(n8958) );
  AOI21_X1 U10136 ( .B1(n9094), .B2(n8959), .A(n8958), .ZN(n9095) );
  INV_X1 U10137 ( .A(n8960), .ZN(n8961) );
  AOI22_X1 U10138 ( .A1(n10821), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8961), 
        .B2(n10813), .ZN(n8962) );
  OAI21_X1 U10139 ( .B1(n8964), .B2(n8963), .A(n8962), .ZN(n8973) );
  OAI211_X1 U10140 ( .C1(n8967), .C2(n8966), .A(n8965), .B(n10808), .ZN(n8971)
         );
  AOI22_X1 U10141 ( .A1(n9014), .A2(n8969), .B1(n8968), .B2(n9016), .ZN(n8970)
         );
  AND2_X1 U10142 ( .A1(n8971), .A2(n8970), .ZN(n9097) );
  NOR2_X1 U10143 ( .A1(n9097), .A2(n10821), .ZN(n8972) );
  AOI211_X1 U10144 ( .C1(n9095), .C2(n10764), .A(n8973), .B(n8972), .ZN(n8974)
         );
  OAI21_X1 U10145 ( .B1(n9098), .B2(n9008), .A(n8974), .ZN(P2_U3278) );
  NAND2_X1 U10146 ( .A1(n8976), .A2(n8978), .ZN(n8977) );
  XOR2_X1 U10147 ( .A(n8979), .B(n8978), .Z(n8981) );
  AOI21_X1 U10148 ( .B1(n8981), .B2(n10808), .A(n8980), .ZN(n9102) );
  INV_X1 U10149 ( .A(n8982), .ZN(n9000) );
  XNOR2_X1 U10150 ( .A(n9000), .B(n9100), .ZN(n8983) );
  NOR2_X1 U10151 ( .A1(n8983), .A2(n11030), .ZN(n9099) );
  NAND2_X1 U10152 ( .A1(n9099), .A2(n6223), .ZN(n8984) );
  OAI211_X1 U10153 ( .C1(n9103), .C2(n8985), .A(n9102), .B(n8984), .ZN(n8986)
         );
  NAND2_X1 U10154 ( .A1(n8986), .A2(n10818), .ZN(n8991) );
  OAI22_X1 U10155 ( .A1(n10818), .A2(n8727), .B1(n8988), .B2(n8987), .ZN(n8989) );
  AOI21_X1 U10156 ( .B1(n9100), .B2(n10767), .A(n8989), .ZN(n8990) );
  OAI211_X1 U10157 ( .C1(n9103), .C2(n8992), .A(n8991), .B(n8990), .ZN(
        P2_U3279) );
  AOI21_X1 U10158 ( .B1(n7939), .B2(n8994), .A(n8993), .ZN(n8996) );
  XNOR2_X1 U10159 ( .A(n8996), .B(n8995), .ZN(n8998) );
  AOI21_X1 U10160 ( .B1(n8998), .B2(n10808), .A(n8997), .ZN(n9107) );
  AOI21_X1 U10161 ( .B1(n9105), .B2(n8999), .A(n11030), .ZN(n9001) );
  AND2_X1 U10162 ( .A1(n9001), .A2(n9000), .ZN(n9104) );
  NAND2_X1 U10163 ( .A1(n9105), .A2(n10767), .ZN(n9004) );
  NAND2_X1 U10164 ( .A1(n10813), .A2(n9002), .ZN(n9003) );
  OAI211_X1 U10165 ( .C1(n10818), .C2(n8709), .A(n9004), .B(n9003), .ZN(n9010)
         );
  OAI21_X1 U10166 ( .B1(n9007), .B2(n9006), .A(n9005), .ZN(n9108) );
  NOR2_X1 U10167 ( .A1(n9108), .A2(n9008), .ZN(n9009) );
  AOI211_X1 U10168 ( .C1(n9104), .C2(n9011), .A(n9010), .B(n9009), .ZN(n9012)
         );
  OAI21_X1 U10169 ( .B1(n10821), .B2(n9107), .A(n9012), .ZN(P2_U3280) );
  XNOR2_X1 U10170 ( .A(n9022), .B(n9013), .ZN(n9018) );
  AOI222_X1 U10171 ( .A1(n10808), .A2(n9018), .B1(n9017), .B2(n9016), .C1(
        n9015), .C2(n9014), .ZN(n10871) );
  MUX2_X1 U10172 ( .A(n6735), .B(n10871), .S(n10818), .Z(n9031) );
  AOI22_X1 U10173 ( .A1(n10767), .A2(n10863), .B1(n9019), .B2(n10813), .ZN(
        n9030) );
  NAND2_X1 U10174 ( .A1(n9021), .A2(n9020), .ZN(n9023) );
  NAND2_X1 U10175 ( .A1(n9023), .A2(n9022), .ZN(n10867) );
  NAND3_X1 U10176 ( .A1(n10868), .A2(n10867), .A3(n9024), .ZN(n9029) );
  AND2_X1 U10177 ( .A1(n10863), .A2(n9025), .ZN(n9026) );
  NOR2_X1 U10178 ( .A1(n9027), .A2(n9026), .ZN(n10866) );
  NAND2_X1 U10179 ( .A1(n10866), .A2(n10764), .ZN(n9028) );
  NAND4_X1 U10180 ( .A1(n9031), .A2(n9030), .A3(n9029), .A4(n9028), .ZN(
        P2_U3290) );
  NAND2_X1 U10181 ( .A1(n9032), .A2(n10864), .ZN(n9033) );
  MUX2_X1 U10182 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9114), .S(n11037), .Z(
        P2_U3551) );
  INV_X1 U10183 ( .A(n9036), .ZN(n9037) );
  AOI21_X1 U10184 ( .B1(n9038), .B2(n10864), .A(n9037), .ZN(n9039) );
  NAND2_X1 U10185 ( .A1(n9040), .A2(n9039), .ZN(n9115) );
  MUX2_X1 U10186 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9115), .S(n11037), .Z(
        P2_U3550) );
  AOI22_X1 U10187 ( .A1(n9042), .A2(n10865), .B1(n10864), .B2(n9041), .ZN(
        n9043) );
  OAI211_X1 U10188 ( .C1(n9045), .C2(n11008), .A(n9044), .B(n9043), .ZN(n9116)
         );
  MUX2_X1 U10189 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9116), .S(n11037), .Z(
        P2_U3548) );
  AOI22_X1 U10190 ( .A1(n9047), .A2(n10865), .B1(n10864), .B2(n9046), .ZN(
        n9048) );
  OAI211_X1 U10191 ( .C1(n9050), .C2(n11008), .A(n9049), .B(n9048), .ZN(n9117)
         );
  MUX2_X1 U10192 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9117), .S(n11037), .Z(
        P2_U3547) );
  AOI21_X1 U10193 ( .B1(n10864), .B2(n9052), .A(n9051), .ZN(n9053) );
  OAI211_X1 U10194 ( .C1(n9055), .C2(n11008), .A(n9054), .B(n9053), .ZN(n9118)
         );
  MUX2_X1 U10195 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9118), .S(n11037), .Z(
        P2_U3546) );
  AOI21_X1 U10196 ( .B1(n10864), .B2(n9057), .A(n9056), .ZN(n9058) );
  OAI211_X1 U10197 ( .C1(n9060), .C2(n11008), .A(n9059), .B(n9058), .ZN(n9119)
         );
  MUX2_X1 U10198 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9119), .S(n11037), .Z(
        P2_U3545) );
  INV_X1 U10199 ( .A(n9061), .ZN(n9066) );
  AOI22_X1 U10200 ( .A1(n9063), .A2(n10865), .B1(n10864), .B2(n9062), .ZN(
        n9064) );
  OAI211_X1 U10201 ( .C1(n9066), .C2(n11008), .A(n9065), .B(n9064), .ZN(n9120)
         );
  MUX2_X1 U10202 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9120), .S(n11037), .Z(
        P2_U3544) );
  NAND2_X1 U10203 ( .A1(n9067), .A2(n11034), .ZN(n9072) );
  AOI22_X1 U10204 ( .A1(n9069), .A2(n10865), .B1(n10864), .B2(n9068), .ZN(
        n9070) );
  OAI211_X1 U10205 ( .C1(n9073), .C2(n9072), .A(n9071), .B(n9070), .ZN(n9121)
         );
  MUX2_X1 U10206 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9121), .S(n11037), .Z(
        P2_U3543) );
  AOI22_X1 U10207 ( .A1(n9075), .A2(n10865), .B1(n10864), .B2(n9074), .ZN(
        n9076) );
  OAI211_X1 U10208 ( .C1(n9078), .C2(n11008), .A(n9077), .B(n9076), .ZN(n9122)
         );
  MUX2_X1 U10209 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9122), .S(n11037), .Z(
        P2_U3542) );
  AOI22_X1 U10210 ( .A1(n9080), .A2(n10865), .B1(n10864), .B2(n9079), .ZN(
        n9081) );
  OAI211_X1 U10211 ( .C1(n9083), .C2(n11008), .A(n9082), .B(n9081), .ZN(n9123)
         );
  MUX2_X1 U10212 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9123), .S(n11037), .Z(
        P2_U3541) );
  AOI22_X1 U10213 ( .A1(n9085), .A2(n10865), .B1(n10864), .B2(n9084), .ZN(
        n9086) );
  OAI211_X1 U10214 ( .C1(n9088), .C2(n11008), .A(n9087), .B(n9086), .ZN(n9124)
         );
  MUX2_X1 U10215 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9124), .S(n11037), .Z(
        P2_U3540) );
  AOI211_X1 U10216 ( .C1(n10864), .C2(n9091), .A(n9090), .B(n9089), .ZN(n9092)
         );
  OAI21_X1 U10217 ( .B1(n9093), .B2(n11008), .A(n9092), .ZN(n9125) );
  MUX2_X1 U10218 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9125), .S(n11037), .Z(
        P2_U3539) );
  AOI22_X1 U10219 ( .A1(n9095), .A2(n10865), .B1(n10864), .B2(n9094), .ZN(
        n9096) );
  OAI211_X1 U10220 ( .C1(n9098), .C2(n11008), .A(n9097), .B(n9096), .ZN(n9126)
         );
  MUX2_X1 U10221 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9126), .S(n11037), .Z(
        P2_U3538) );
  AOI21_X1 U10222 ( .B1(n10864), .B2(n9100), .A(n9099), .ZN(n9101) );
  OAI211_X1 U10223 ( .C1(n9103), .C2(n11008), .A(n9102), .B(n9101), .ZN(n9127)
         );
  MUX2_X1 U10224 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9127), .S(n11037), .Z(
        P2_U3537) );
  AOI21_X1 U10225 ( .B1(n10864), .B2(n9105), .A(n9104), .ZN(n9106) );
  OAI211_X1 U10226 ( .C1(n9108), .C2(n11008), .A(n9107), .B(n9106), .ZN(n9128)
         );
  MUX2_X1 U10227 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9128), .S(n11037), .Z(
        P2_U3536) );
  AOI22_X1 U10228 ( .A1(n9110), .A2(n10865), .B1(n10864), .B2(n9109), .ZN(
        n9111) );
  OAI211_X1 U10229 ( .C1(n9113), .C2(n11008), .A(n9112), .B(n9111), .ZN(n9129)
         );
  MUX2_X1 U10230 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9129), .S(n11037), .Z(
        P2_U3535) );
  MUX2_X1 U10231 ( .A(n9115), .B(P2_REG0_REG_30__SCAN_IN), .S(n11038), .Z(
        P2_U3518) );
  MUX2_X1 U10232 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9116), .S(n11041), .Z(
        P2_U3516) );
  MUX2_X1 U10233 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9117), .S(n11041), .Z(
        P2_U3515) );
  MUX2_X1 U10234 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9118), .S(n11041), .Z(
        P2_U3514) );
  MUX2_X1 U10235 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9119), .S(n11041), .Z(
        P2_U3513) );
  MUX2_X1 U10236 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9120), .S(n11041), .Z(
        P2_U3512) );
  MUX2_X1 U10237 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9121), .S(n11041), .Z(
        P2_U3511) );
  MUX2_X1 U10238 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9122), .S(n11041), .Z(
        P2_U3510) );
  MUX2_X1 U10239 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9123), .S(n11041), .Z(
        P2_U3509) );
  MUX2_X1 U10240 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9124), .S(n11041), .Z(
        P2_U3508) );
  MUX2_X1 U10241 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9125), .S(n11041), .Z(
        P2_U3507) );
  MUX2_X1 U10242 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9126), .S(n11041), .Z(
        P2_U3505) );
  MUX2_X1 U10243 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9127), .S(n11041), .Z(
        P2_U3502) );
  MUX2_X1 U10244 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9128), .S(n11041), .Z(
        P2_U3499) );
  MUX2_X1 U10245 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9129), .S(n11041), .Z(
        P2_U3496) );
  INV_X1 U10246 ( .A(n9391), .ZN(n10444) );
  INV_X1 U10247 ( .A(n9130), .ZN(n9132) );
  NOR4_X1 U10248 ( .A1(n9132), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n9131), .ZN(n9133) );
  AOI21_X1 U10249 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9134), .A(n9133), .ZN(
        n9135) );
  OAI21_X1 U10250 ( .B1(n10444), .B2(n9147), .A(n9135), .ZN(P2_U3327) );
  INV_X1 U10251 ( .A(n9136), .ZN(n10446) );
  OAI222_X1 U10252 ( .A1(n9147), .A2(n10446), .B1(n9138), .B2(P2_U3152), .C1(
        n9137), .C2(n9146), .ZN(P2_U3329) );
  INV_X1 U10253 ( .A(n10451), .ZN(n9141) );
  OAI222_X1 U10254 ( .A1(n9147), .A2(n9141), .B1(n9140), .B2(P2_U3152), .C1(
        n9139), .C2(n9146), .ZN(P2_U3331) );
  INV_X1 U10255 ( .A(n9142), .ZN(n10456) );
  OAI222_X1 U10256 ( .A1(n9147), .A2(n10456), .B1(P2_U3152), .B2(n9144), .C1(
        n9143), .C2(n9146), .ZN(P2_U3332) );
  INV_X1 U10257 ( .A(n10469), .ZN(n9148) );
  INV_X1 U10258 ( .A(n9145), .ZN(n10460) );
  OAI222_X1 U10259 ( .A1(P2_U3152), .A2(n9148), .B1(n9147), .B2(n10460), .C1(
        n9146), .C2(n6142), .ZN(P2_U3333) );
  MUX2_X1 U10260 ( .A(n9150), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10261 ( .A(n9151), .ZN(n9155) );
  XNOR2_X1 U10262 ( .A(n9153), .B(n9152), .ZN(n9154) );
  XNOR2_X1 U10263 ( .A(n9155), .B(n9154), .ZN(n9161) );
  NOR2_X1 U10264 ( .A1(n9314), .A2(n10303), .ZN(n9156) );
  AOI211_X1 U10265 ( .C1(n9300), .C2(n10276), .A(n9157), .B(n9156), .ZN(n9158)
         );
  OAI21_X1 U10266 ( .B1(n9315), .B2(n10310), .A(n9158), .ZN(n9159) );
  AOI21_X1 U10267 ( .B1(n10316), .B2(n9292), .A(n9159), .ZN(n9160) );
  OAI21_X1 U10268 ( .B1(n9161), .B2(n9309), .A(n9160), .ZN(P1_U3213) );
  INV_X1 U10269 ( .A(n9162), .ZN(n9163) );
  NOR2_X1 U10270 ( .A1(n9164), .A2(n9163), .ZN(n9166) );
  XNOR2_X1 U10271 ( .A(n9166), .B(n9165), .ZN(n9171) );
  AOI22_X1 U10272 ( .A1(n9318), .A2(n10164), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9168) );
  NAND2_X1 U10273 ( .A1(n9289), .A2(n10192), .ZN(n9167) );
  OAI211_X1 U10274 ( .C1(n9315), .C2(n10157), .A(n9168), .B(n9167), .ZN(n9169)
         );
  AOI21_X1 U10275 ( .B1(n10353), .B2(n9220), .A(n9169), .ZN(n9170) );
  OAI21_X1 U10276 ( .B1(n9171), .B2(n9309), .A(n9170), .ZN(P1_U3214) );
  XOR2_X1 U10277 ( .A(n9173), .B(n9172), .Z(n9178) );
  NAND2_X1 U10278 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10081)
         );
  OAI21_X1 U10279 ( .B1(n9287), .B2(n9208), .A(n10081), .ZN(n9174) );
  AOI21_X1 U10280 ( .B1(n9289), .B2(n10223), .A(n9174), .ZN(n9175) );
  OAI21_X1 U10281 ( .B1(n9315), .B2(n10231), .A(n9175), .ZN(n9176) );
  AOI21_X1 U10282 ( .B1(n10374), .B2(n9292), .A(n9176), .ZN(n9177) );
  OAI21_X1 U10283 ( .B1(n9178), .B2(n9309), .A(n9177), .ZN(P1_U3217) );
  NAND2_X1 U10284 ( .A1(n10328), .A2(n9181), .ZN(n9184) );
  NAND2_X1 U10285 ( .A1(n10102), .A2(n9182), .ZN(n9183) );
  NAND2_X1 U10286 ( .A1(n9184), .A2(n9183), .ZN(n9186) );
  XNOR2_X1 U10287 ( .A(n9186), .B(n9185), .ZN(n9191) );
  NOR2_X1 U10288 ( .A1(n9188), .A2(n9187), .ZN(n9189) );
  AOI21_X1 U10289 ( .B1(n10328), .B2(n7802), .A(n9189), .ZN(n9190) );
  XNOR2_X1 U10290 ( .A(n9191), .B(n9190), .ZN(n9197) );
  NAND4_X1 U10291 ( .A1(n9192), .A2(n9295), .A3(n9196), .A4(n9197), .ZN(n9202)
         );
  AOI22_X1 U10292 ( .A1(n9289), .A2(n9610), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n9195) );
  NAND2_X1 U10293 ( .A1(n9303), .A2(n9193), .ZN(n9194) );
  OAI211_X1 U10294 ( .C1(n9467), .C2(n9287), .A(n9195), .B(n9194), .ZN(n9199)
         );
  NOR3_X1 U10295 ( .A1(n9197), .A2(n9309), .A3(n9196), .ZN(n9198) );
  AOI211_X1 U10296 ( .C1(n10328), .C2(n9220), .A(n9199), .B(n9198), .ZN(n9200)
         );
  NAND3_X1 U10297 ( .A1(n9202), .A2(n9201), .A3(n9200), .ZN(P1_U3218) );
  NAND2_X1 U10298 ( .A1(n5104), .A2(n9203), .ZN(n9204) );
  XNOR2_X1 U10299 ( .A(n9205), .B(n9204), .ZN(n9211) );
  NAND2_X1 U10300 ( .A1(n9303), .A2(n10197), .ZN(n9207) );
  AOI22_X1 U10301 ( .A1(n9318), .A2(n10192), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9206) );
  OAI211_X1 U10302 ( .C1(n9208), .C2(n9314), .A(n9207), .B(n9206), .ZN(n9209)
         );
  AOI21_X1 U10303 ( .B1(n10364), .B2(n9292), .A(n9209), .ZN(n9210) );
  OAI21_X1 U10304 ( .B1(n9211), .B2(n9309), .A(n9210), .ZN(P1_U3221) );
  INV_X1 U10305 ( .A(n9212), .ZN(n9214) );
  NAND2_X1 U10306 ( .A1(n9214), .A2(n9213), .ZN(n9215) );
  XNOR2_X1 U10307 ( .A(n9216), .B(n9215), .ZN(n9222) );
  AOI22_X1 U10308 ( .A1(n9318), .A2(n10135), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9218) );
  NAND2_X1 U10309 ( .A1(n9289), .A2(n10164), .ZN(n9217) );
  OAI211_X1 U10310 ( .C1(n9315), .C2(n10128), .A(n9218), .B(n9217), .ZN(n9219)
         );
  AOI21_X1 U10311 ( .B1(n10343), .B2(n9220), .A(n9219), .ZN(n9221) );
  OAI21_X1 U10312 ( .B1(n9222), .B2(n9309), .A(n9221), .ZN(P1_U3223) );
  AOI21_X1 U10313 ( .B1(n9225), .B2(n9224), .A(n9223), .ZN(n9230) );
  NAND2_X1 U10314 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10052)
         );
  OAI21_X1 U10315 ( .B1(n9314), .B2(n10304), .A(n10052), .ZN(n9226) );
  AOI21_X1 U10316 ( .B1(n9300), .B2(n10277), .A(n9226), .ZN(n9227) );
  OAI21_X1 U10317 ( .B1(n9315), .B2(n10270), .A(n9227), .ZN(n9228) );
  AOI21_X1 U10318 ( .B1(n10389), .B2(n9292), .A(n9228), .ZN(n9229) );
  OAI21_X1 U10319 ( .B1(n9230), .B2(n9309), .A(n9229), .ZN(P1_U3224) );
  INV_X1 U10320 ( .A(n9231), .ZN(n9232) );
  NOR2_X1 U10321 ( .A1(n9233), .A2(n9232), .ZN(n9234) );
  XNOR2_X1 U10322 ( .A(n9235), .B(n9234), .ZN(n9240) );
  NAND2_X1 U10323 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10058)
         );
  OAI21_X1 U10324 ( .B1(n9287), .B2(n10251), .A(n10058), .ZN(n9236) );
  AOI21_X1 U10325 ( .B1(n9289), .B2(n10294), .A(n9236), .ZN(n9237) );
  OAI21_X1 U10326 ( .B1(n9315), .B2(n10260), .A(n9237), .ZN(n9238) );
  AOI21_X1 U10327 ( .B1(n10383), .B2(n9292), .A(n9238), .ZN(n9239) );
  OAI21_X1 U10328 ( .B1(n9240), .B2(n9309), .A(n9239), .ZN(P1_U3226) );
  OAI21_X1 U10329 ( .B1(n9243), .B2(n9242), .A(n9241), .ZN(n9244) );
  NAND2_X1 U10330 ( .A1(n9244), .A2(n9295), .ZN(n9249) );
  INV_X1 U10331 ( .A(n9245), .ZN(n10147) );
  AOI22_X1 U10332 ( .A1(n9289), .A2(n10180), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9246) );
  OAI21_X1 U10333 ( .B1(n10110), .B2(n9287), .A(n9246), .ZN(n9247) );
  AOI21_X1 U10334 ( .B1(n10147), .B2(n9303), .A(n9247), .ZN(n9248) );
  OAI211_X1 U10335 ( .C1(n5316), .C2(n9321), .A(n9249), .B(n9248), .ZN(
        P1_U3227) );
  XNOR2_X1 U10336 ( .A(n9251), .B(n9250), .ZN(n9252) );
  XNOR2_X1 U10337 ( .A(n9253), .B(n9252), .ZN(n9259) );
  OAI22_X1 U10338 ( .A1(n10205), .A2(n9287), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9254), .ZN(n9255) );
  AOI21_X1 U10339 ( .B1(n9289), .B2(n10243), .A(n9255), .ZN(n9256) );
  OAI21_X1 U10340 ( .B1(n9315), .B2(n10212), .A(n9256), .ZN(n9257) );
  AOI21_X1 U10341 ( .B1(n10368), .B2(n9292), .A(n9257), .ZN(n9258) );
  OAI21_X1 U10342 ( .B1(n9259), .B2(n9309), .A(n9258), .ZN(P1_U3231) );
  XOR2_X1 U10343 ( .A(n9261), .B(n9260), .Z(n9262) );
  XNOR2_X1 U10344 ( .A(n9263), .B(n9262), .ZN(n9271) );
  NOR2_X1 U10345 ( .A1(n9314), .A2(n9264), .ZN(n9265) );
  AOI211_X1 U10346 ( .C1(n9318), .C2(n10293), .A(n9266), .B(n9265), .ZN(n9267)
         );
  OAI21_X1 U10347 ( .B1(n9315), .B2(n9268), .A(n9267), .ZN(n9269) );
  AOI21_X1 U10348 ( .B1(n10398), .B2(n9292), .A(n9269), .ZN(n9270) );
  OAI21_X1 U10349 ( .B1(n9271), .B2(n9309), .A(n9270), .ZN(P1_U3232) );
  INV_X1 U10350 ( .A(n9272), .ZN(n9273) );
  NOR2_X1 U10351 ( .A1(n9274), .A2(n9273), .ZN(n9275) );
  XNOR2_X1 U10352 ( .A(n9276), .B(n9275), .ZN(n9281) );
  NAND2_X1 U10353 ( .A1(n10179), .A2(n9289), .ZN(n9278) );
  AOI22_X1 U10354 ( .A1(n10180), .A2(n9300), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3084), .ZN(n9277) );
  OAI211_X1 U10355 ( .C1(n9315), .C2(n10172), .A(n9278), .B(n9277), .ZN(n9279)
         );
  AOI21_X1 U10356 ( .B1(n10358), .B2(n9292), .A(n9279), .ZN(n9280) );
  OAI21_X1 U10357 ( .B1(n9281), .B2(n9309), .A(n9280), .ZN(P1_U3233) );
  INV_X1 U10358 ( .A(n9282), .ZN(n9283) );
  NOR2_X1 U10359 ( .A1(n9284), .A2(n9283), .ZN(n9286) );
  XNOR2_X1 U10360 ( .A(n9286), .B(n9285), .ZN(n9294) );
  NAND2_X1 U10361 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10580)
         );
  OAI21_X1 U10362 ( .B1(n9287), .B2(n10204), .A(n10580), .ZN(n9288) );
  AOI21_X1 U10363 ( .B1(n9289), .B2(n10277), .A(n9288), .ZN(n9290) );
  OAI21_X1 U10364 ( .B1(n9315), .B2(n10237), .A(n9290), .ZN(n9291) );
  AOI21_X1 U10365 ( .B1(n10378), .B2(n9292), .A(n9291), .ZN(n9293) );
  OAI21_X1 U10366 ( .B1(n9294), .B2(n9309), .A(n9293), .ZN(P1_U3236) );
  INV_X1 U10367 ( .A(n10338), .ZN(n10120) );
  OAI211_X1 U10368 ( .C1(n9298), .C2(n9297), .A(n9296), .B(n9295), .ZN(n9305)
         );
  INV_X1 U10369 ( .A(n9299), .ZN(n10118) );
  AOI22_X1 U10370 ( .A1(n9610), .A2(n9300), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9301) );
  OAI21_X1 U10371 ( .B1(n10110), .B2(n9314), .A(n9301), .ZN(n9302) );
  AOI21_X1 U10372 ( .B1(n10118), .B2(n9303), .A(n9302), .ZN(n9304) );
  OAI211_X1 U10373 ( .C1(n10120), .C2(n9321), .A(n9305), .B(n9304), .ZN(
        P1_U3238) );
  INV_X1 U10374 ( .A(n9307), .ZN(n9313) );
  AOI21_X1 U10375 ( .B1(n9308), .B2(n9307), .A(n9306), .ZN(n9310) );
  NOR2_X1 U10376 ( .A1(n9310), .A2(n9309), .ZN(n9311) );
  OAI21_X1 U10377 ( .B1(n9313), .B2(n9312), .A(n9311), .ZN(n9320) );
  NAND2_X1 U10378 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10029)
         );
  OAI21_X1 U10379 ( .B1(n9314), .B2(n9533), .A(n10029), .ZN(n9317) );
  NOR2_X1 U10380 ( .A1(n9315), .A2(n10287), .ZN(n9316) );
  AOI211_X1 U10381 ( .C1(n9318), .C2(n10294), .A(n9317), .B(n9316), .ZN(n9319)
         );
  OAI211_X1 U10382 ( .C1(n10290), .C2(n9321), .A(n9320), .B(n9319), .ZN(
        P1_U3239) );
  NAND2_X1 U10383 ( .A1(n9511), .A2(n9506), .ZN(n9322) );
  NAND2_X1 U10384 ( .A1(n9322), .A2(n9510), .ZN(n9323) );
  AND3_X1 U10385 ( .A1(n9530), .A2(n9518), .A3(n9323), .ZN(n9324) );
  NAND2_X1 U10386 ( .A1(n9523), .A2(n9324), .ZN(n9351) );
  NAND2_X1 U10387 ( .A1(n9510), .A2(n9325), .ZN(n9508) );
  NOR2_X1 U10388 ( .A1(n9508), .A2(n9326), .ZN(n9327) );
  OR2_X1 U10389 ( .A1(n9351), .A2(n9327), .ZN(n9331) );
  NAND2_X1 U10390 ( .A1(n9530), .A2(n5456), .ZN(n9328) );
  NAND2_X1 U10391 ( .A1(n9328), .A2(n9526), .ZN(n9329) );
  NAND2_X1 U10392 ( .A1(n9523), .A2(n9329), .ZN(n9330) );
  NAND4_X1 U10393 ( .A1(n9331), .A2(n9528), .A3(n9527), .A4(n9330), .ZN(n9332)
         );
  NAND3_X1 U10394 ( .A1(n9547), .A2(n9524), .A3(n9332), .ZN(n9333) );
  NAND2_X1 U10395 ( .A1(n9333), .A2(n9546), .ZN(n9334) );
  AND2_X1 U10396 ( .A1(n9556), .A2(n9552), .ZN(n9350) );
  OAI211_X1 U10397 ( .C1(n9335), .C2(n9334), .A(n9560), .B(n9350), .ZN(n9412)
         );
  INV_X1 U10398 ( .A(n9336), .ZN(n9337) );
  OAI211_X1 U10399 ( .C1(n9338), .C2(n10726), .A(n9595), .B(n9337), .ZN(n9340)
         );
  NAND2_X1 U10400 ( .A1(n9340), .A2(n9339), .ZN(n9343) );
  OAI22_X1 U10401 ( .A1(n9344), .A2(n9343), .B1(n9342), .B2(n9341), .ZN(n9347)
         );
  AND2_X1 U10402 ( .A1(n9404), .A2(n9345), .ZN(n9431) );
  INV_X1 U10403 ( .A(n9431), .ZN(n9346) );
  AOI21_X1 U10404 ( .B1(n9347), .B2(n9403), .A(n9346), .ZN(n9348) );
  NOR3_X1 U10405 ( .A1(n9348), .A2(n5457), .A3(n9401), .ZN(n9358) );
  NAND2_X1 U10406 ( .A1(n9496), .A2(n9349), .ZN(n9491) );
  INV_X1 U10407 ( .A(n9491), .ZN(n9409) );
  NAND2_X1 U10408 ( .A1(n9409), .A2(n9399), .ZN(n9357) );
  INV_X1 U10409 ( .A(n9350), .ZN(n9354) );
  INV_X1 U10410 ( .A(n9351), .ZN(n9352) );
  NAND4_X1 U10411 ( .A1(n9547), .A2(n9352), .A3(n9524), .A4(n10911), .ZN(n9353) );
  NOR2_X1 U10412 ( .A1(n9354), .A2(n9353), .ZN(n9355) );
  NAND2_X1 U10413 ( .A1(n9355), .A2(n9560), .ZN(n9414) );
  INV_X1 U10414 ( .A(n9414), .ZN(n9356) );
  OAI211_X1 U10415 ( .C1(n9358), .C2(n9357), .A(n9356), .B(n9500), .ZN(n9367)
         );
  INV_X1 U10416 ( .A(n9359), .ZN(n9360) );
  NAND2_X1 U10417 ( .A1(n9369), .A2(n9360), .ZN(n9361) );
  AND2_X1 U10418 ( .A1(n9361), .A2(n9484), .ZN(n9486) );
  INV_X1 U10419 ( .A(n9486), .ZN(n9363) );
  INV_X1 U10420 ( .A(n9566), .ZN(n9362) );
  NOR2_X1 U10421 ( .A1(n9363), .A2(n9362), .ZN(n9364) );
  AND4_X1 U10422 ( .A1(n9478), .A2(n9364), .A3(n9481), .A4(n9483), .ZN(n9365)
         );
  AND2_X1 U10423 ( .A1(n9477), .A2(n9365), .ZN(n9416) );
  INV_X1 U10424 ( .A(n9416), .ZN(n9366) );
  AOI21_X1 U10425 ( .B1(n9412), .B2(n9367), .A(n9366), .ZN(n9382) );
  NAND2_X1 U10426 ( .A1(n9369), .A2(n9368), .ZN(n9485) );
  INV_X1 U10427 ( .A(n9555), .ZN(n9370) );
  NAND2_X1 U10428 ( .A1(n9560), .A2(n9370), .ZN(n9371) );
  NAND2_X1 U10429 ( .A1(n9371), .A2(n9561), .ZN(n9372) );
  NAND2_X1 U10430 ( .A1(n9566), .A2(n9372), .ZN(n9373) );
  NAND2_X1 U10431 ( .A1(n9373), .A2(n9565), .ZN(n9374) );
  OAI211_X1 U10432 ( .C1(n9485), .C2(n9374), .A(n9486), .B(n9483), .ZN(n9375)
         );
  NAND2_X1 U10433 ( .A1(n9375), .A2(n9482), .ZN(n9376) );
  NAND2_X1 U10434 ( .A1(n9376), .A2(n9481), .ZN(n9377) );
  NAND3_X1 U10435 ( .A1(n9479), .A2(n9377), .A3(n9480), .ZN(n9378) );
  NAND3_X1 U10436 ( .A1(n9477), .A2(n9478), .A3(n9378), .ZN(n9379) );
  AND2_X1 U10437 ( .A1(n9379), .A2(n9476), .ZN(n9380) );
  AND2_X1 U10438 ( .A1(n9380), .A2(n9475), .ZN(n9418) );
  INV_X1 U10439 ( .A(n9418), .ZN(n9381) );
  NOR3_X1 U10440 ( .A1(n5184), .A2(n9382), .A3(n9381), .ZN(n9387) );
  INV_X1 U10441 ( .A(n9474), .ZN(n9384) );
  INV_X1 U10442 ( .A(n9466), .ZN(n9383) );
  AOI211_X1 U10443 ( .C1(n9385), .C2(n9473), .A(n9384), .B(n9383), .ZN(n9421)
         );
  INV_X1 U10444 ( .A(n9421), .ZN(n9386) );
  NOR2_X1 U10445 ( .A1(n9387), .A2(n9386), .ZN(n9389) );
  NAND2_X1 U10446 ( .A1(n9388), .A2(n9468), .ZN(n9419) );
  INV_X1 U10447 ( .A(n9608), .ZN(n9395) );
  NAND2_X1 U10448 ( .A1(n11047), .A2(n9395), .ZN(n9448) );
  OAI211_X1 U10449 ( .C1(n9389), .C2(n9419), .A(n9448), .B(n9422), .ZN(n9396)
         );
  NAND2_X1 U10450 ( .A1(n9391), .A2(n9390), .ZN(n9394) );
  INV_X1 U10451 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9392) );
  OR2_X1 U10452 ( .A1(n7060), .A2(n9392), .ZN(n9393) );
  INV_X1 U10453 ( .A(n10322), .ZN(n9460) );
  INV_X1 U10454 ( .A(n9607), .ZN(n9426) );
  OR2_X1 U10455 ( .A1(n11047), .A2(n9395), .ZN(n9459) );
  NAND3_X1 U10456 ( .A1(n9396), .A2(n9456), .A3(n9459), .ZN(n9397) );
  NAND2_X1 U10457 ( .A1(n9397), .A2(n9594), .ZN(n9398) );
  XNOR2_X1 U10458 ( .A(n9398), .B(n10730), .ZN(n9599) );
  NAND3_X1 U10459 ( .A1(n9400), .A2(n9431), .A3(n9399), .ZN(n9408) );
  INV_X1 U10460 ( .A(n9401), .ZN(n9407) );
  AND2_X1 U10461 ( .A1(n9403), .A2(n9402), .ZN(n9430) );
  INV_X1 U10462 ( .A(n9430), .ZN(n9405) );
  NAND3_X1 U10463 ( .A1(n9405), .A2(n9404), .A3(n10837), .ZN(n9406) );
  NAND3_X1 U10464 ( .A1(n9408), .A2(n9407), .A3(n9406), .ZN(n9410) );
  NAND2_X1 U10465 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  NAND2_X1 U10466 ( .A1(n9411), .A2(n9500), .ZN(n9413) );
  OAI21_X1 U10467 ( .B1(n9414), .B2(n9413), .A(n9412), .ZN(n9415) );
  NAND2_X1 U10468 ( .A1(n9416), .A2(n9415), .ZN(n9417) );
  NAND3_X1 U10469 ( .A1(n9473), .A2(n9418), .A3(n9417), .ZN(n9420) );
  AOI21_X1 U10470 ( .B1(n9421), .B2(n9420), .A(n9419), .ZN(n9425) );
  INV_X1 U10471 ( .A(n9422), .ZN(n9424) );
  NAND2_X1 U10472 ( .A1(n11047), .A2(n9426), .ZN(n9423) );
  NAND2_X1 U10473 ( .A1(n9448), .A2(n9423), .ZN(n9462) );
  NOR3_X1 U10474 ( .A1(n9425), .A2(n9424), .A3(n9462), .ZN(n9428) );
  OR2_X1 U10475 ( .A1(n9459), .A2(n9426), .ZN(n9427) );
  NAND2_X1 U10476 ( .A1(n9456), .A2(n9427), .ZN(n9458) );
  OAI211_X1 U10477 ( .C1(n9428), .C2(n9458), .A(n9595), .B(n9594), .ZN(n9454)
         );
  INV_X1 U10478 ( .A(n10143), .ZN(n9445) );
  INV_X1 U10479 ( .A(n10178), .ZN(n10169) );
  INV_X1 U10480 ( .A(n10709), .ZN(n10715) );
  NAND4_X1 U10481 ( .A1(n9432), .A2(n9431), .A3(n9488), .A4(n9430), .ZN(n9433)
         );
  INV_X1 U10482 ( .A(n10838), .ZN(n10832) );
  NOR4_X1 U10483 ( .A1(n10715), .A2(n9434), .A3(n9433), .A4(n10832), .ZN(n9436) );
  NAND4_X1 U10484 ( .A1(n9436), .A2(n10913), .A3(n9503), .A4(n9435), .ZN(n9437) );
  NOR4_X1 U10485 ( .A1(n9438), .A2(n9514), .A3(n5452), .A4(n9437), .ZN(n9439)
         );
  NAND3_X1 U10486 ( .A1(n10307), .A2(n9440), .A3(n9439), .ZN(n9441) );
  NOR4_X1 U10487 ( .A1(n10252), .A2(n10274), .A3(n10292), .A4(n9441), .ZN(
        n9442) );
  NAND4_X1 U10488 ( .A1(n10191), .A2(n10222), .A3(n9558), .A4(n9442), .ZN(
        n9443) );
  NOR4_X1 U10489 ( .A1(n9445), .A2(n10169), .A3(n9444), .A4(n9443), .ZN(n9446)
         );
  NOR3_X1 U10490 ( .A1(n9451), .A2(n9450), .A3(n9449), .ZN(n9452) );
  NOR2_X1 U10491 ( .A1(n9452), .A2(n9595), .ZN(n9590) );
  INV_X1 U10492 ( .A(n9590), .ZN(n9453) );
  NAND2_X1 U10493 ( .A1(n9462), .A2(n9559), .ZN(n9455) );
  NAND2_X1 U10494 ( .A1(n9455), .A2(n9594), .ZN(n9457) );
  NAND2_X1 U10495 ( .A1(n9457), .A2(n9456), .ZN(n9589) );
  INV_X1 U10496 ( .A(n9559), .ZN(n9564) );
  NAND2_X1 U10497 ( .A1(n9458), .A2(n9564), .ZN(n9588) );
  NAND2_X1 U10498 ( .A1(n9459), .A2(n9607), .ZN(n9461) );
  NAND2_X1 U10499 ( .A1(n9461), .A2(n9460), .ZN(n9587) );
  INV_X1 U10500 ( .A(n9462), .ZN(n9586) );
  NAND2_X1 U10501 ( .A1(n9468), .A2(n9467), .ZN(n9463) );
  NAND3_X1 U10502 ( .A1(n9464), .A2(n9559), .A3(n9463), .ZN(n9472) );
  INV_X1 U10503 ( .A(n9467), .ZN(n9609) );
  NAND2_X1 U10504 ( .A1(n9466), .A2(n9609), .ZN(n9465) );
  NAND3_X1 U10505 ( .A1(n9465), .A2(n10323), .A3(n9564), .ZN(n9471) );
  OR3_X1 U10506 ( .A1(n9466), .A2(n9609), .A3(n9559), .ZN(n9470) );
  OR3_X1 U10507 ( .A1(n9468), .A2(n9467), .A3(n9564), .ZN(n9469) );
  AND4_X1 U10508 ( .A1(n9472), .A2(n9471), .A3(n9470), .A4(n9469), .ZN(n9585)
         );
  MUX2_X1 U10509 ( .A(n9474), .B(n9473), .S(n9564), .Z(n9580) );
  MUX2_X1 U10510 ( .A(n10097), .B(n9475), .S(n9559), .Z(n9578) );
  MUX2_X1 U10511 ( .A(n9477), .B(n9476), .S(n9564), .Z(n9576) );
  MUX2_X1 U10512 ( .A(n9479), .B(n9478), .S(n9564), .Z(n9574) );
  MUX2_X1 U10513 ( .A(n9481), .B(n9480), .S(n9564), .Z(n9572) );
  MUX2_X1 U10514 ( .A(n9483), .B(n9482), .S(n9559), .Z(n9571) );
  NAND2_X1 U10515 ( .A1(n9485), .A2(n9484), .ZN(n9487) );
  MUX2_X1 U10516 ( .A(n9487), .B(n9486), .S(n9559), .Z(n9570) );
  NAND2_X1 U10517 ( .A1(n9489), .A2(n9488), .ZN(n9490) );
  OAI211_X1 U10518 ( .C1(n9559), .C2(n10835), .A(n9490), .B(n10838), .ZN(n9495) );
  INV_X1 U10519 ( .A(n9495), .ZN(n9492) );
  OAI21_X1 U10520 ( .B1(n9492), .B2(n9491), .A(n10911), .ZN(n9499) );
  OAI211_X1 U10521 ( .C1(n9495), .C2(n9494), .A(n10911), .B(n9493), .ZN(n9497)
         );
  NAND2_X1 U10522 ( .A1(n9497), .A2(n9496), .ZN(n9498) );
  MUX2_X1 U10523 ( .A(n9499), .B(n9498), .S(n9559), .Z(n9505) );
  MUX2_X1 U10524 ( .A(n9501), .B(n9500), .S(n9559), .Z(n9502) );
  OAI21_X1 U10525 ( .B1(n9506), .B2(n9559), .A(n9511), .ZN(n9507) );
  AOI21_X1 U10526 ( .B1(n9508), .B2(n9559), .A(n9507), .ZN(n9509) );
  MUX2_X1 U10527 ( .A(n9511), .B(n9510), .S(n9564), .Z(n9512) );
  NAND2_X1 U10528 ( .A1(n9513), .A2(n9512), .ZN(n9516) );
  INV_X1 U10529 ( .A(n9514), .ZN(n9515) );
  NAND2_X1 U10530 ( .A1(n9516), .A2(n9515), .ZN(n9520) );
  MUX2_X1 U10531 ( .A(n9518), .B(n9517), .S(n9564), .Z(n9519) );
  NAND2_X1 U10532 ( .A1(n9520), .A2(n9519), .ZN(n9522) );
  NAND3_X1 U10533 ( .A1(n9524), .A2(n9564), .A3(n9523), .ZN(n9525) );
  AOI21_X1 U10534 ( .B1(n9531), .B2(n9526), .A(n9525), .ZN(n9545) );
  NAND3_X1 U10535 ( .A1(n9528), .A2(n9527), .A3(n9559), .ZN(n9529) );
  AOI21_X1 U10536 ( .B1(n9531), .B2(n9530), .A(n9529), .ZN(n9544) );
  NAND2_X1 U10537 ( .A1(n10303), .A2(n9559), .ZN(n9537) );
  INV_X1 U10538 ( .A(n9537), .ZN(n9532) );
  AOI22_X1 U10539 ( .A1(n10398), .A2(n9532), .B1(n9533), .B2(n9559), .ZN(n9542) );
  NAND2_X1 U10540 ( .A1(n10007), .A2(n9564), .ZN(n9535) );
  OAI22_X1 U10541 ( .A1(n10398), .A2(n9535), .B1(n9533), .B2(n9559), .ZN(n9534) );
  NAND2_X1 U10542 ( .A1(n11022), .A2(n9534), .ZN(n9541) );
  INV_X1 U10543 ( .A(n9535), .ZN(n9536) );
  AND2_X1 U10544 ( .A1(n9536), .A2(n10293), .ZN(n9539) );
  OAI21_X1 U10545 ( .B1(n10293), .B2(n9537), .A(n10398), .ZN(n9538) );
  OAI21_X1 U10546 ( .B1(n9539), .B2(n10398), .A(n9538), .ZN(n9540) );
  OAI211_X1 U10547 ( .C1(n11022), .C2(n9542), .A(n9541), .B(n9540), .ZN(n9543)
         );
  MUX2_X1 U10548 ( .A(n9547), .B(n9546), .S(n9559), .Z(n9548) );
  NAND3_X1 U10549 ( .A1(n9550), .A2(n9549), .A3(n9548), .ZN(n9554) );
  INV_X1 U10550 ( .A(n10252), .ZN(n10248) );
  MUX2_X1 U10551 ( .A(n9552), .B(n9551), .S(n9564), .Z(n9553) );
  MUX2_X1 U10552 ( .A(n9556), .B(n9555), .S(n9559), .Z(n9557) );
  MUX2_X1 U10553 ( .A(n9561), .B(n9560), .S(n9559), .Z(n9562) );
  NAND2_X1 U10554 ( .A1(n9563), .A2(n10222), .ZN(n9568) );
  MUX2_X1 U10555 ( .A(n9566), .B(n9565), .S(n9564), .Z(n9567) );
  NAND3_X1 U10556 ( .A1(n10134), .A2(n9574), .A3(n9573), .ZN(n9575) );
  NAND3_X1 U10557 ( .A1(n10112), .A2(n9576), .A3(n9575), .ZN(n9577) );
  NAND3_X1 U10558 ( .A1(n10098), .A2(n9578), .A3(n9577), .ZN(n9579) );
  NAND3_X1 U10559 ( .A1(n9581), .A2(n9580), .A3(n9579), .ZN(n9583) );
  OR2_X1 U10560 ( .A1(n9583), .A2(n9582), .ZN(n9584) );
  AOI21_X1 U10561 ( .B1(n9593), .B2(n9591), .A(n9590), .ZN(n9592) );
  INV_X1 U10562 ( .A(n9593), .ZN(n9596) );
  NAND4_X1 U10563 ( .A1(n9596), .A2(n9595), .A3(n6889), .A4(n9594), .ZN(n9597)
         );
  NAND3_X1 U10564 ( .A1(n9601), .A2(n10669), .A3(n9600), .ZN(n9602) );
  OAI211_X1 U10565 ( .C1(n9603), .C2(n9605), .A(n9602), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9604) );
  OAI21_X1 U10566 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(P1_U3240) );
  MUX2_X1 U10567 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9607), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10568 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9608), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10569 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9609), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10570 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n10102), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10571 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9610), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10572 ( .A(n10135), .B(P1_DATAO_REG_26__SCAN_IN), .S(n10671), .Z(
        P1_U3581) );
  MUX2_X1 U10573 ( .A(n10164), .B(P1_DATAO_REG_24__SCAN_IN), .S(n10671), .Z(
        P1_U3579) );
  MUX2_X1 U10574 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n10180), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10575 ( .A(n10192), .B(P1_DATAO_REG_22__SCAN_IN), .S(n10671), .Z(
        P1_U3577) );
  MUX2_X1 U10576 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10179), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10577 ( .A(n10224), .B(P1_DATAO_REG_20__SCAN_IN), .S(n10671), .Z(
        P1_U3575) );
  MUX2_X1 U10578 ( .A(n10243), .B(P1_DATAO_REG_19__SCAN_IN), .S(n10671), .Z(
        P1_U3574) );
  INV_X1 U10579 ( .A(keyinput_233), .ZN(n9784) );
  XNOR2_X1 U10580 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .ZN(n9757)
         );
  AOI22_X1 U10581 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput_203), .B1(
        n9612), .B2(keyinput_204), .ZN(n9611) );
  OAI221_X1 U10582 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_203), .C1(
        n9612), .C2(keyinput_204), .A(n9611), .ZN(n9742) );
  INV_X1 U10583 ( .A(keyinput_199), .ZN(n9737) );
  INV_X1 U10584 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9614) );
  OAI22_X1 U10585 ( .A1(n9614), .A2(keyinput_191), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_194), .ZN(n9613) );
  AOI221_X1 U10586 ( .B1(n9614), .B2(keyinput_191), .C1(keyinput_194), .C2(
        P2_DATAO_REG_30__SCAN_IN), .A(n9613), .ZN(n9618) );
  OAI22_X1 U10587 ( .A1(n10445), .A2(keyinput_195), .B1(n9616), .B2(
        keyinput_192), .ZN(n9615) );
  AOI221_X1 U10588 ( .B1(n10445), .B2(keyinput_195), .C1(keyinput_192), .C2(
        n9616), .A(n9615), .ZN(n9617) );
  OAI211_X1 U10589 ( .C1(P2_DATAO_REG_31__SCAN_IN), .C2(keyinput_193), .A(
        n9618), .B(n9617), .ZN(n9619) );
  AOI21_X1 U10590 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_193), .A(n9619), .ZN(n9735) );
  INV_X1 U10591 ( .A(keyinput_190), .ZN(n9729) );
  INV_X1 U10592 ( .A(keyinput_189), .ZN(n9727) );
  OAI22_X1 U10593 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_181), .B1(
        keyinput_182), .B2(P2_REG3_REG_0__SCAN_IN), .ZN(n9620) );
  AOI221_X1 U10594 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_181), .C1(
        P2_REG3_REG_0__SCAN_IN), .C2(keyinput_182), .A(n9620), .ZN(n9716) );
  OAI22_X1 U10595 ( .A1(n9622), .A2(keyinput_177), .B1(keyinput_176), .B2(
        P2_REG3_REG_16__SCAN_IN), .ZN(n9621) );
  AOI221_X1 U10596 ( .B1(n9622), .B2(keyinput_177), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_176), .A(n9621), .ZN(n9707) );
  AOI22_X1 U10597 ( .A1(SI_3_), .A2(keyinput_157), .B1(SI_4_), .B2(
        keyinput_156), .ZN(n9623) );
  OAI221_X1 U10598 ( .B1(SI_3_), .B2(keyinput_157), .C1(SI_4_), .C2(
        keyinput_156), .A(n9623), .ZN(n9676) );
  INV_X1 U10599 ( .A(keyinput_151), .ZN(n9669) );
  AOI22_X1 U10600 ( .A1(SI_15_), .A2(keyinput_145), .B1(n9625), .B2(
        keyinput_144), .ZN(n9624) );
  OAI221_X1 U10601 ( .B1(SI_15_), .B2(keyinput_145), .C1(n9625), .C2(
        keyinput_144), .A(n9624), .ZN(n9660) );
  INV_X1 U10602 ( .A(keyinput_143), .ZN(n9659) );
  INV_X1 U10603 ( .A(SI_17_), .ZN(n9658) );
  AOI22_X1 U10604 ( .A1(SI_20_), .A2(keyinput_140), .B1(n9627), .B2(
        keyinput_141), .ZN(n9626) );
  OAI221_X1 U10605 ( .B1(SI_20_), .B2(keyinput_140), .C1(n9627), .C2(
        keyinput_141), .A(n9626), .ZN(n9655) );
  OAI22_X1 U10606 ( .A1(SI_31_), .A2(keyinput_129), .B1(P2_WR_REG_SCAN_IN), 
        .B2(keyinput_128), .ZN(n9628) );
  INV_X1 U10607 ( .A(keyinput_130), .ZN(n9629) );
  MUX2_X1 U10608 ( .A(n9629), .B(keyinput_130), .S(SI_30_), .Z(n9630) );
  OAI22_X1 U10609 ( .A1(n9632), .A2(keyinput_132), .B1(n9631), .B2(
        keyinput_131), .ZN(n9636) );
  INV_X1 U10610 ( .A(SI_24_), .ZN(n9644) );
  AOI22_X1 U10611 ( .A1(n9644), .A2(keyinput_136), .B1(n9643), .B2(
        keyinput_135), .ZN(n9642) );
  OAI221_X1 U10612 ( .B1(n9644), .B2(keyinput_136), .C1(n9643), .C2(
        keyinput_135), .A(n9642), .ZN(n9645) );
  OAI22_X1 U10613 ( .A1(SI_26_), .A2(keyinput_134), .B1(SI_23_), .B2(
        keyinput_137), .ZN(n9646) );
  AOI221_X1 U10614 ( .B1(SI_26_), .B2(keyinput_134), .C1(keyinput_137), .C2(
        SI_23_), .A(n9646), .ZN(n9647) );
  AOI22_X1 U10615 ( .A1(SI_21_), .A2(keyinput_139), .B1(n9650), .B2(
        keyinput_138), .ZN(n9649) );
  OAI221_X1 U10616 ( .B1(SI_21_), .B2(keyinput_139), .C1(n9650), .C2(
        keyinput_138), .A(n9649), .ZN(n9651) );
  OAI22_X1 U10617 ( .A1(keyinput_142), .A2(n9657), .B1(n9655), .B2(n9654), 
        .ZN(n9656) );
  AOI22_X1 U10618 ( .A1(SI_13_), .A2(keyinput_147), .B1(n9662), .B2(
        keyinput_150), .ZN(n9661) );
  OAI221_X1 U10619 ( .B1(SI_13_), .B2(keyinput_147), .C1(n9662), .C2(
        keyinput_150), .A(n9661), .ZN(n9665) );
  AOI22_X1 U10620 ( .A1(SI_12_), .A2(keyinput_148), .B1(SI_11_), .B2(
        keyinput_149), .ZN(n9663) );
  OAI221_X1 U10621 ( .B1(SI_12_), .B2(keyinput_148), .C1(SI_11_), .C2(
        keyinput_149), .A(n9663), .ZN(n9664) );
  AOI22_X1 U10622 ( .A1(n9672), .A2(keyinput_152), .B1(keyinput_154), .B2(
        n9671), .ZN(n9670) );
  OAI221_X1 U10623 ( .B1(n9672), .B2(keyinput_152), .C1(n9671), .C2(
        keyinput_154), .A(n9670), .ZN(n9675) );
  AOI22_X1 U10624 ( .A1(SI_5_), .A2(keyinput_155), .B1(SI_7_), .B2(
        keyinput_153), .ZN(n9673) );
  OAI221_X1 U10625 ( .B1(SI_5_), .B2(keyinput_155), .C1(SI_7_), .C2(
        keyinput_153), .A(n9673), .ZN(n9674) );
  OAI22_X1 U10626 ( .A1(SI_2_), .A2(keyinput_158), .B1(keyinput_159), .B2(
        SI_1_), .ZN(n9677) );
  AOI221_X1 U10627 ( .B1(SI_2_), .B2(keyinput_158), .C1(SI_1_), .C2(
        keyinput_159), .A(n9677), .ZN(n9684) );
  AOI22_X1 U10628 ( .A1(P2_U3152), .A2(keyinput_162), .B1(n9679), .B2(
        keyinput_164), .ZN(n9678) );
  OAI221_X1 U10629 ( .B1(P2_U3152), .B2(keyinput_162), .C1(n9679), .C2(
        keyinput_164), .A(n9678), .ZN(n9683) );
  AOI22_X1 U10630 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_161), .B1(n9681), 
        .B2(keyinput_163), .ZN(n9680) );
  OAI221_X1 U10631 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_161), .C1(n9681), 
        .C2(keyinput_163), .A(n9680), .ZN(n9682) );
  AOI22_X1 U10632 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_166), .B1(n5991), .B2(keyinput_165), .ZN(n9686) );
  OAI221_X1 U10633 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_166), .C1(
        n5991), .C2(keyinput_165), .A(n9686), .ZN(n9691) );
  XNOR2_X1 U10634 ( .A(keyinput_167), .B(n9687), .ZN(n9690) );
  OAI22_X1 U10635 ( .A1(n10763), .A2(keyinput_168), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_169), .ZN(n9688) );
  AOI221_X1 U10636 ( .B1(n10763), .B2(keyinput_168), .C1(keyinput_169), .C2(
        P2_REG3_REG_19__SCAN_IN), .A(n9688), .ZN(n9689) );
  OAI211_X1 U10637 ( .C1(n9692), .C2(n9691), .A(n9690), .B(n9689), .ZN(n9698)
         );
  OAI22_X1 U10638 ( .A1(n9694), .A2(keyinput_170), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(keyinput_171), .ZN(n9693) );
  AOI221_X1 U10639 ( .B1(n9694), .B2(keyinput_170), .C1(keyinput_171), .C2(
        P2_REG3_REG_8__SCAN_IN), .A(n9693), .ZN(n9697) );
  INV_X1 U10640 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9696) );
  NOR2_X1 U10641 ( .A1(n9696), .A2(keyinput_172), .ZN(n9695) );
  AOI221_X1 U10642 ( .B1(n9698), .B2(n9697), .C1(keyinput_172), .C2(n9696), 
        .A(n9695), .ZN(n9705) );
  AOI22_X1 U10643 ( .A1(n9701), .A2(keyinput_173), .B1(n9700), .B2(
        keyinput_174), .ZN(n9699) );
  OAI221_X1 U10644 ( .B1(n9701), .B2(keyinput_173), .C1(n9700), .C2(
        keyinput_174), .A(n9699), .ZN(n9704) );
  INV_X1 U10645 ( .A(keyinput_178), .ZN(n9714) );
  AOI22_X1 U10646 ( .A1(n9711), .A2(keyinput_179), .B1(n9710), .B2(
        keyinput_180), .ZN(n9709) );
  OAI221_X1 U10647 ( .B1(n9711), .B2(keyinput_179), .C1(n9710), .C2(
        keyinput_180), .A(n9709), .ZN(n9712) );
  INV_X1 U10648 ( .A(n9712), .ZN(n9713) );
  XNOR2_X1 U10649 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_184), .ZN(n9723)
         );
  INV_X1 U10650 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9718) );
  OAI22_X1 U10651 ( .A1(n9719), .A2(keyinput_186), .B1(n9718), .B2(
        keyinput_188), .ZN(n9717) );
  AOI221_X1 U10652 ( .B1(n9719), .B2(keyinput_186), .C1(keyinput_188), .C2(
        n9718), .A(n9717), .ZN(n9722) );
  OAI22_X1 U10653 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_185), .B1(
        keyinput_187), .B2(P2_REG3_REG_2__SCAN_IN), .ZN(n9720) );
  AOI221_X1 U10654 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_185), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_187), .A(n9720), .ZN(n9721) );
  OAI211_X1 U10655 ( .C1(n9724), .C2(n9723), .A(n9722), .B(n9721), .ZN(n9725)
         );
  OAI221_X1 U10656 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(n9727), .C1(n9726), .C2(
        keyinput_189), .A(n9725), .ZN(n9728) );
  OAI221_X1 U10657 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_190), .C1(
        n9730), .C2(n9729), .A(n9728), .ZN(n9734) );
  XOR2_X1 U10658 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .Z(n9733)
         );
  AOI22_X1 U10659 ( .A1(n10448), .A2(keyinput_196), .B1(keyinput_198), .B2(
        n10455), .ZN(n9731) );
  OAI221_X1 U10660 ( .B1(n10448), .B2(keyinput_196), .C1(n10455), .C2(
        keyinput_198), .A(n9731), .ZN(n9732) );
  AOI221_X1 U10661 ( .B1(P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_199), .C1(
        n10459), .C2(n9737), .A(n9736), .ZN(n9741) );
  OAI22_X1 U10662 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_200), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(keyinput_202), .ZN(n9738) );
  AOI221_X1 U10663 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_200), .C1(
        keyinput_202), .C2(P2_DATAO_REG_22__SCAN_IN), .A(n9738), .ZN(n9739) );
  OAI21_X1 U10664 ( .B1(keyinput_201), .B2(P2_DATAO_REG_23__SCAN_IN), .A(n9739), .ZN(n9740) );
  AOI22_X1 U10665 ( .A1(n9746), .A2(keyinput_206), .B1(keyinput_208), .B2(
        n9745), .ZN(n9744) );
  OAI221_X1 U10666 ( .B1(n9746), .B2(keyinput_206), .C1(n9745), .C2(
        keyinput_208), .A(n9744), .ZN(n9747) );
  OAI21_X1 U10667 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_207), .A(n9748), .ZN(n9756) );
  AOI22_X1 U10668 ( .A1(n9751), .A2(keyinput_213), .B1(n9750), .B2(
        keyinput_210), .ZN(n9749) );
  OAI221_X1 U10669 ( .B1(n9751), .B2(keyinput_213), .C1(n9750), .C2(
        keyinput_210), .A(n9749), .ZN(n9755) );
  AOI22_X1 U10670 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(keyinput_212), .B1(
        n9753), .B2(keyinput_211), .ZN(n9752) );
  OAI221_X1 U10671 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_212), .C1(
        n9753), .C2(keyinput_211), .A(n9752), .ZN(n9754) );
  XNOR2_X1 U10672 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n9763)
         );
  OAI22_X1 U10673 ( .A1(n9759), .A2(keyinput_216), .B1(keyinput_215), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n9758) );
  AOI221_X1 U10674 ( .B1(n9759), .B2(keyinput_216), .C1(
        P2_DATAO_REG_9__SCAN_IN), .C2(keyinput_215), .A(n9758), .ZN(n9762) );
  OAI22_X1 U10675 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_217), .B1(
        keyinput_218), .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n9760) );
  AOI221_X1 U10676 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_217), .C1(
        P2_DATAO_REG_6__SCAN_IN), .C2(keyinput_218), .A(n9760), .ZN(n9761) );
  OAI211_X1 U10677 ( .C1(n9764), .C2(n9763), .A(n9762), .B(n9761), .ZN(n9769)
         );
  OAI22_X1 U10678 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_220), .B1(
        keyinput_219), .B2(P1_IR_REG_0__SCAN_IN), .ZN(n9765) );
  AOI221_X1 U10679 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_220), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput_219), .A(n9765), .ZN(n9768) );
  XOR2_X1 U10680 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_222), .Z(n9767) );
  XNOR2_X1 U10681 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_221), .ZN(n9766) );
  AOI211_X1 U10682 ( .C1(n9769), .C2(n9768), .A(n9767), .B(n9766), .ZN(n9774)
         );
  XOR2_X1 U10683 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_223), .Z(n9773) );
  OAI22_X1 U10684 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(keyinput_224), .B1(
        keyinput_225), .B2(P1_IR_REG_6__SCAN_IN), .ZN(n9770) );
  AOI221_X1 U10685 ( .B1(P1_IR_REG_5__SCAN_IN), .B2(keyinput_224), .C1(
        P1_IR_REG_6__SCAN_IN), .C2(keyinput_225), .A(n9770), .ZN(n9771) );
  INV_X1 U10686 ( .A(n9771), .ZN(n9772) );
  OAI22_X1 U10687 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_228), .B1(
        keyinput_229), .B2(P1_IR_REG_10__SCAN_IN), .ZN(n9775) );
  AOI221_X1 U10688 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_228), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_229), .A(n9775), .ZN(n9778) );
  XNOR2_X1 U10689 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_227), .ZN(n9777) );
  XNOR2_X1 U10690 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_226), .ZN(n9776) );
  XNOR2_X1 U10691 ( .A(n9779), .B(keyinput_230), .ZN(n9781) );
  XNOR2_X1 U10692 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_231), .ZN(n9780) );
  NOR2_X1 U10693 ( .A1(n9781), .A2(n9780), .ZN(n9782) );
  OAI221_X1 U10694 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_233), .C1(n9968), 
        .C2(n9784), .A(n9783), .ZN(n9788) );
  OAI22_X1 U10695 ( .A1(n7187), .A2(keyinput_236), .B1(P1_IR_REG_16__SCAN_IN), 
        .B2(keyinput_235), .ZN(n9785) );
  AOI221_X1 U10696 ( .B1(n7187), .B2(keyinput_236), .C1(keyinput_235), .C2(
        P1_IR_REG_16__SCAN_IN), .A(n9785), .ZN(n9787) );
  XNOR2_X1 U10697 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_234), .ZN(n9786) );
  INV_X1 U10698 ( .A(keyinput_237), .ZN(n9789) );
  MUX2_X1 U10699 ( .A(keyinput_237), .B(n9789), .S(P1_IR_REG_18__SCAN_IN), .Z(
        n9790) );
  AOI22_X1 U10700 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_243), .B1(
        P1_IR_REG_21__SCAN_IN), .B2(keyinput_240), .ZN(n9791) );
  OAI221_X1 U10701 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_243), .C1(
        P1_IR_REG_21__SCAN_IN), .C2(keyinput_240), .A(n9791), .ZN(n9795) );
  XOR2_X1 U10702 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_244), .Z(n9794) );
  XNOR2_X1 U10703 ( .A(n5471), .B(keyinput_242), .ZN(n9793) );
  XNOR2_X1 U10704 ( .A(keyinput_241), .B(n6493), .ZN(n9792) );
  NOR4_X1 U10705 ( .A1(n9795), .A2(n9794), .A3(n9793), .A4(n9792), .ZN(n9798)
         );
  OAI22_X1 U10706 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput_238), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput_239), .ZN(n9796) );
  AOI221_X1 U10707 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput_238), .C1(
        keyinput_239), .C2(P1_IR_REG_20__SCAN_IN), .A(n9796), .ZN(n9797) );
  AND2_X1 U10708 ( .A1(n9798), .A2(n9797), .ZN(n9799) );
  INV_X1 U10709 ( .A(keyinput_246), .ZN(n9800) );
  MUX2_X1 U10710 ( .A(n9800), .B(keyinput_246), .S(P1_IR_REG_27__SCAN_IN), .Z(
        n9801) );
  NAND2_X1 U10711 ( .A1(n9802), .A2(n9801), .ZN(n9805) );
  INV_X1 U10712 ( .A(keyinput_247), .ZN(n9803) );
  MUX2_X1 U10713 ( .A(keyinput_247), .B(n9803), .S(P1_IR_REG_28__SCAN_IN), .Z(
        n9804) );
  NAND2_X1 U10714 ( .A1(n9805), .A2(n9804), .ZN(n9808) );
  INV_X1 U10715 ( .A(keyinput_248), .ZN(n9806) );
  MUX2_X1 U10716 ( .A(keyinput_248), .B(n9806), .S(P1_IR_REG_29__SCAN_IN), .Z(
        n9807) );
  NAND2_X1 U10717 ( .A1(n9808), .A2(n9807), .ZN(n9813) );
  INV_X1 U10718 ( .A(keyinput_249), .ZN(n9809) );
  MUX2_X1 U10719 ( .A(n9809), .B(keyinput_249), .S(P1_IR_REG_30__SCAN_IN), .Z(
        n9812) );
  XOR2_X1 U10720 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_250), .Z(n9811) );
  XNOR2_X1 U10721 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_251), .ZN(n9810) );
  XNOR2_X1 U10722 ( .A(keyinput_252), .B(P1_D_REG_1__SCAN_IN), .ZN(n9815) );
  XNOR2_X1 U10723 ( .A(keyinput_253), .B(P1_D_REG_2__SCAN_IN), .ZN(n9814) );
  OAI21_X1 U10724 ( .B1(n9816), .B2(n9815), .A(n9814), .ZN(n9819) );
  XOR2_X1 U10725 ( .A(keyinput_255), .B(P1_D_REG_4__SCAN_IN), .Z(n9818) );
  INV_X1 U10726 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10465) );
  XNOR2_X1 U10727 ( .A(n10465), .B(keyinput_254), .ZN(n9817) );
  NAND3_X1 U10728 ( .A1(n9819), .A2(n9818), .A3(n9817), .ZN(n10004) );
  XOR2_X1 U10729 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_127), .Z(n10003) );
  XOR2_X1 U10730 ( .A(SI_30_), .B(keyinput_2), .Z(n9822) );
  XNOR2_X1 U10731 ( .A(SI_31_), .B(keyinput_1), .ZN(n9821) );
  XNOR2_X1 U10732 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n9820) );
  NOR3_X1 U10733 ( .A1(n9822), .A2(n9821), .A3(n9820), .ZN(n9825) );
  XNOR2_X1 U10734 ( .A(SI_28_), .B(keyinput_4), .ZN(n9824) );
  XNOR2_X1 U10735 ( .A(SI_29_), .B(keyinput_3), .ZN(n9823) );
  NOR3_X1 U10736 ( .A1(n9825), .A2(n9824), .A3(n9823), .ZN(n9832) );
  XNOR2_X1 U10737 ( .A(SI_27_), .B(keyinput_5), .ZN(n9831) );
  XOR2_X1 U10738 ( .A(SI_23_), .B(keyinput_9), .Z(n9829) );
  XOR2_X1 U10739 ( .A(SI_26_), .B(keyinput_6), .Z(n9828) );
  XOR2_X1 U10740 ( .A(SI_25_), .B(keyinput_7), .Z(n9827) );
  XNOR2_X1 U10741 ( .A(SI_24_), .B(keyinput_8), .ZN(n9826) );
  NOR4_X1 U10742 ( .A1(n9829), .A2(n9828), .A3(n9827), .A4(n9826), .ZN(n9830)
         );
  OAI21_X1 U10743 ( .B1(n9832), .B2(n9831), .A(n9830), .ZN(n9835) );
  XNOR2_X1 U10744 ( .A(SI_22_), .B(keyinput_10), .ZN(n9834) );
  XNOR2_X1 U10745 ( .A(SI_21_), .B(keyinput_11), .ZN(n9833) );
  NAND3_X1 U10746 ( .A1(n9835), .A2(n9834), .A3(n9833), .ZN(n9838) );
  XOR2_X1 U10747 ( .A(SI_19_), .B(keyinput_13), .Z(n9837) );
  XNOR2_X1 U10748 ( .A(SI_20_), .B(keyinput_12), .ZN(n9836) );
  NAND3_X1 U10749 ( .A1(n9838), .A2(n9837), .A3(n9836), .ZN(n9841) );
  XNOR2_X1 U10750 ( .A(SI_18_), .B(keyinput_14), .ZN(n9840) );
  XOR2_X1 U10751 ( .A(SI_17_), .B(keyinput_15), .Z(n9839) );
  AOI21_X1 U10752 ( .B1(n9841), .B2(n9840), .A(n9839), .ZN(n9844) );
  XOR2_X1 U10753 ( .A(SI_15_), .B(keyinput_17), .Z(n9843) );
  XNOR2_X1 U10754 ( .A(SI_16_), .B(keyinput_16), .ZN(n9842) );
  NOR3_X1 U10755 ( .A1(n9844), .A2(n9843), .A3(n9842), .ZN(n9851) );
  XNOR2_X1 U10756 ( .A(SI_14_), .B(keyinput_18), .ZN(n9850) );
  XOR2_X1 U10757 ( .A(SI_12_), .B(keyinput_20), .Z(n9848) );
  XOR2_X1 U10758 ( .A(SI_11_), .B(keyinput_21), .Z(n9847) );
  XNOR2_X1 U10759 ( .A(SI_10_), .B(keyinput_22), .ZN(n9846) );
  XNOR2_X1 U10760 ( .A(SI_13_), .B(keyinput_19), .ZN(n9845) );
  NOR4_X1 U10761 ( .A1(n9848), .A2(n9847), .A3(n9846), .A4(n9845), .ZN(n9849)
         );
  OAI21_X1 U10762 ( .B1(n9851), .B2(n9850), .A(n9849), .ZN(n9858) );
  XNOR2_X1 U10763 ( .A(SI_9_), .B(keyinput_23), .ZN(n9857) );
  XOR2_X1 U10764 ( .A(SI_5_), .B(keyinput_27), .Z(n9855) );
  XOR2_X1 U10765 ( .A(SI_8_), .B(keyinput_24), .Z(n9854) );
  XOR2_X1 U10766 ( .A(SI_6_), .B(keyinput_26), .Z(n9853) );
  XNOR2_X1 U10767 ( .A(SI_7_), .B(keyinput_25), .ZN(n9852) );
  NAND4_X1 U10768 ( .A1(n9855), .A2(n9854), .A3(n9853), .A4(n9852), .ZN(n9856)
         );
  AOI21_X1 U10769 ( .B1(n9858), .B2(n9857), .A(n9856), .ZN(n9861) );
  XNOR2_X1 U10770 ( .A(SI_3_), .B(keyinput_29), .ZN(n9860) );
  XNOR2_X1 U10771 ( .A(SI_4_), .B(keyinput_28), .ZN(n9859) );
  NOR3_X1 U10772 ( .A1(n9861), .A2(n9860), .A3(n9859), .ZN(n9865) );
  XOR2_X1 U10773 ( .A(SI_0_), .B(keyinput_32), .Z(n9864) );
  XOR2_X1 U10774 ( .A(SI_1_), .B(keyinput_31), .Z(n9863) );
  XOR2_X1 U10775 ( .A(SI_2_), .B(keyinput_30), .Z(n9862) );
  NOR4_X1 U10776 ( .A1(n9865), .A2(n9864), .A3(n9863), .A4(n9862), .ZN(n9873)
         );
  XOR2_X1 U10777 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .Z(n9869) );
  XOR2_X1 U10778 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_34), .Z(n9868) );
  XOR2_X1 U10779 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .Z(n9867) );
  XNOR2_X1 U10780 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n9866) );
  NAND4_X1 U10781 ( .A1(n9869), .A2(n9868), .A3(n9867), .A4(n9866), .ZN(n9872)
         );
  XOR2_X1 U10782 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_37), .Z(n9871) );
  XNOR2_X1 U10783 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n9870)
         );
  OAI211_X1 U10784 ( .C1(n9873), .C2(n9872), .A(n9871), .B(n9870), .ZN(n9877)
         );
  XOR2_X1 U10785 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .Z(n9876) );
  XOR2_X1 U10786 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_41), .Z(n9875) );
  XOR2_X1 U10787 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .Z(n9874) );
  NAND4_X1 U10788 ( .A1(n9877), .A2(n9876), .A3(n9875), .A4(n9874), .ZN(n9880)
         );
  XOR2_X1 U10789 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_43), .Z(n9879) );
  XNOR2_X1 U10790 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n9878)
         );
  NAND3_X1 U10791 ( .A1(n9880), .A2(n9879), .A3(n9878), .ZN(n9886) );
  XOR2_X1 U10792 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n9885) );
  XNOR2_X1 U10793 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n9883)
         );
  XNOR2_X1 U10794 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_47), .ZN(n9882)
         );
  XNOR2_X1 U10795 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput_45), .ZN(n9881)
         );
  NAND3_X1 U10796 ( .A1(n9883), .A2(n9882), .A3(n9881), .ZN(n9884) );
  AOI21_X1 U10797 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9889) );
  XOR2_X1 U10798 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_48), .Z(n9888) );
  XOR2_X1 U10799 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_49), .Z(n9887) );
  NOR3_X1 U10800 ( .A1(n9889), .A2(n9888), .A3(n9887), .ZN(n9896) );
  XOR2_X1 U10801 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_50), .Z(n9895) );
  XOR2_X1 U10802 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_53), .Z(n9893) );
  XNOR2_X1 U10803 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n9892) );
  XNOR2_X1 U10804 ( .A(P2_REG3_REG_24__SCAN_IN), .B(keyinput_51), .ZN(n9891)
         );
  XNOR2_X1 U10805 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n9890) );
  NOR4_X1 U10806 ( .A1(n9893), .A2(n9892), .A3(n9891), .A4(n9890), .ZN(n9894)
         );
  OAI21_X1 U10807 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(n9899) );
  XNOR2_X1 U10808 ( .A(P2_REG3_REG_20__SCAN_IN), .B(keyinput_55), .ZN(n9898)
         );
  XOR2_X1 U10809 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput_56), .Z(n9897) );
  AOI21_X1 U10810 ( .B1(n9899), .B2(n9898), .A(n9897), .ZN(n9906) );
  XOR2_X1 U10811 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .Z(n9903) );
  XOR2_X1 U10812 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .Z(n9902) );
  XNOR2_X1 U10813 ( .A(P2_REG3_REG_11__SCAN_IN), .B(keyinput_58), .ZN(n9901)
         );
  XNOR2_X1 U10814 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_57), .ZN(n9900)
         );
  NAND4_X1 U10815 ( .A1(n9903), .A2(n9902), .A3(n9901), .A4(n9900), .ZN(n9905)
         );
  XNOR2_X1 U10816 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n9904) );
  OAI21_X1 U10817 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9915) );
  XNOR2_X1 U10818 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n9914)
         );
  XOR2_X1 U10819 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_66), .Z(n9909) );
  XOR2_X1 U10820 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_65), .Z(n9908) );
  XOR2_X1 U10821 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .Z(n9907) );
  NOR3_X1 U10822 ( .A1(n9909), .A2(n9908), .A3(n9907), .ZN(n9912) );
  XNOR2_X1 U10823 ( .A(P2_REG3_REG_15__SCAN_IN), .B(keyinput_63), .ZN(n9911)
         );
  XNOR2_X1 U10824 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_64), .ZN(n9910) );
  NAND3_X1 U10825 ( .A1(n9912), .A2(n9911), .A3(n9910), .ZN(n9913) );
  AOI21_X1 U10826 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9922) );
  INV_X1 U10827 ( .A(keyinput_69), .ZN(n9919) );
  XOR2_X1 U10828 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_70), .Z(n9918) );
  OAI22_X1 U10829 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(keyinput_68), .B1(
        keyinput_69), .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9916) );
  AOI21_X1 U10830 ( .B1(P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_68), .A(n9916), 
        .ZN(n9917) );
  OAI211_X1 U10831 ( .C1(n7034), .C2(n9919), .A(n9918), .B(n9917), .ZN(n9921)
         );
  XNOR2_X1 U10832 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n9920)
         );
  OAI21_X1 U10833 ( .B1(n9922), .B2(n9921), .A(n9920), .ZN(n9929) );
  XOR2_X1 U10834 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_72), .Z(n9925) );
  XNOR2_X1 U10835 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_74), .ZN(n9924)
         );
  XNOR2_X1 U10836 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n9923)
         );
  NOR3_X1 U10837 ( .A1(n9925), .A2(n9924), .A3(n9923), .ZN(n9928) );
  XNOR2_X1 U10838 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_76), .ZN(n9927)
         );
  XNOR2_X1 U10839 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .ZN(n9926)
         );
  AOI211_X1 U10840 ( .C1(n9929), .C2(n9928), .A(n9927), .B(n9926), .ZN(n9935)
         );
  XNOR2_X1 U10841 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n9934)
         );
  XOR2_X1 U10842 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n9932) );
  XOR2_X1 U10843 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(keyinput_80), .Z(n9931) );
  XNOR2_X1 U10844 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .ZN(n9930)
         );
  NOR3_X1 U10845 ( .A1(n9932), .A2(n9931), .A3(n9930), .ZN(n9933) );
  OAI21_X1 U10846 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(n9942) );
  XOR2_X1 U10847 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .Z(n9941) );
  XOR2_X1 U10848 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .Z(n9939) );
  XOR2_X1 U10849 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .Z(n9938) );
  XNOR2_X1 U10850 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n9937)
         );
  XNOR2_X1 U10851 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput_82), .ZN(n9936)
         );
  NAND4_X1 U10852 ( .A1(n9939), .A2(n9938), .A3(n9937), .A4(n9936), .ZN(n9940)
         );
  AOI21_X1 U10853 ( .B1(n9942), .B2(n9941), .A(n9940), .ZN(n9949) );
  XNOR2_X1 U10854 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .ZN(n9948)
         );
  XOR2_X1 U10855 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput_90), .Z(n9946) );
  XNOR2_X1 U10856 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .ZN(n9945)
         );
  XNOR2_X1 U10857 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n9944)
         );
  XNOR2_X1 U10858 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .ZN(n9943)
         );
  NOR4_X1 U10859 ( .A1(n9946), .A2(n9945), .A3(n9944), .A4(n9943), .ZN(n9947)
         );
  OAI21_X1 U10860 ( .B1(n9949), .B2(n9948), .A(n9947), .ZN(n9952) );
  XOR2_X1 U10861 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_91), .Z(n9951) );
  XNOR2_X1 U10862 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_92), .ZN(n9950) );
  NAND3_X1 U10863 ( .A1(n9952), .A2(n9951), .A3(n9950), .ZN(n9955) );
  XOR2_X1 U10864 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_94), .Z(n9954) );
  XOR2_X1 U10865 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_93), .Z(n9953) );
  NAND3_X1 U10866 ( .A1(n9955), .A2(n9954), .A3(n9953), .ZN(n9959) );
  XOR2_X1 U10867 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_96), .Z(n9958) );
  XNOR2_X1 U10868 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_97), .ZN(n9957) );
  XNOR2_X1 U10869 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_95), .ZN(n9956) );
  NAND4_X1 U10870 ( .A1(n9959), .A2(n9958), .A3(n9957), .A4(n9956), .ZN(n9967)
         );
  XOR2_X1 U10871 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_98), .Z(n9963) );
  XOR2_X1 U10872 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_99), .Z(n9962) );
  XNOR2_X1 U10873 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_101), .ZN(n9961) );
  XNOR2_X1 U10874 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_100), .ZN(n9960) );
  NOR4_X1 U10875 ( .A1(n9963), .A2(n9962), .A3(n9961), .A4(n9960), .ZN(n9966)
         );
  XOR2_X1 U10876 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_103), .Z(n9965) );
  XNOR2_X1 U10877 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_102), .ZN(n9964) );
  AOI211_X1 U10878 ( .C1(n9967), .C2(n9966), .A(n9965), .B(n9964), .ZN(n9971)
         );
  XNOR2_X1 U10879 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_104), .ZN(n9970) );
  XNOR2_X1 U10880 ( .A(n9968), .B(keyinput_105), .ZN(n9969) );
  OAI21_X1 U10881 ( .B1(n9971), .B2(n9970), .A(n9969), .ZN(n9975) );
  XOR2_X1 U10882 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_106), .Z(n9974) );
  XOR2_X1 U10883 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_107), .Z(n9973) );
  XOR2_X1 U10884 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_108), .Z(n9972) );
  NAND4_X1 U10885 ( .A1(n9975), .A2(n9974), .A3(n9973), .A4(n9972), .ZN(n9977)
         );
  XNOR2_X1 U10886 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_109), .ZN(n9976) );
  NAND2_X1 U10887 ( .A1(n9977), .A2(n9976), .ZN(n9987) );
  XOR2_X1 U10888 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput_116), .Z(n9986) );
  XOR2_X1 U10889 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_110), .Z(n9983) );
  XOR2_X1 U10890 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_112), .Z(n9982) );
  XOR2_X1 U10891 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_114), .Z(n9981) );
  OR2_X1 U10892 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_113), .ZN(n9979) );
  AOI22_X1 U10893 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_115), .B1(
        P1_IR_REG_22__SCAN_IN), .B2(keyinput_113), .ZN(n9978) );
  OAI211_X1 U10894 ( .C1(P1_IR_REG_24__SCAN_IN), .C2(keyinput_115), .A(n9979), 
        .B(n9978), .ZN(n9980) );
  NOR4_X1 U10895 ( .A1(n9983), .A2(n9982), .A3(n9981), .A4(n9980), .ZN(n9985)
         );
  XNOR2_X1 U10896 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_111), .ZN(n9984) );
  NAND4_X1 U10897 ( .A1(n9987), .A2(n9986), .A3(n9985), .A4(n9984), .ZN(n9990)
         );
  XOR2_X1 U10898 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_117), .Z(n9989) );
  XOR2_X1 U10899 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_118), .Z(n9988) );
  AOI21_X1 U10900 ( .B1(n9990), .B2(n9989), .A(n9988), .ZN(n9993) );
  XOR2_X1 U10901 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput_119), .Z(n9992) );
  XOR2_X1 U10902 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_120), .Z(n9991) );
  OAI21_X1 U10903 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(n9997) );
  XOR2_X1 U10904 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_121), .Z(n9996) );
  XOR2_X1 U10905 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_122), .Z(n9995) );
  XOR2_X1 U10906 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_123), .Z(n9994) );
  AOI211_X1 U10907 ( .C1(n9997), .C2(n9996), .A(n9995), .B(n9994), .ZN(n10000)
         );
  XNOR2_X1 U10908 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_124), .ZN(n9999) );
  INV_X1 U10909 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10464) );
  XNOR2_X1 U10910 ( .A(n10464), .B(keyinput_125), .ZN(n9998) );
  OAI21_X1 U10911 ( .B1(n10000), .B2(n9999), .A(n9998), .ZN(n10002) );
  XNOR2_X1 U10912 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_126), .ZN(n10001) );
  NAND4_X1 U10913 ( .A1(n10004), .A2(n10003), .A3(n10002), .A4(n10001), .ZN(
        n10006) );
  MUX2_X1 U10914 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10223), .S(P1_U4006), .Z(
        n10005) );
  XNOR2_X1 U10915 ( .A(n10006), .B(n10005), .ZN(P1_U3573) );
  MUX2_X1 U10916 ( .A(n10277), .B(P1_DATAO_REG_17__SCAN_IN), .S(n10671), .Z(
        P1_U3572) );
  MUX2_X1 U10917 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n10294), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10918 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10276), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10919 ( .A(n10007), .B(P1_DATAO_REG_13__SCAN_IN), .S(n10671), .Z(
        P1_U3568) );
  MUX2_X1 U10920 ( .A(n10008), .B(P1_DATAO_REG_12__SCAN_IN), .S(n10671), .Z(
        P1_U3567) );
  MUX2_X1 U10921 ( .A(n10009), .B(P1_DATAO_REG_11__SCAN_IN), .S(n10671), .Z(
        P1_U3566) );
  MUX2_X1 U10922 ( .A(n10010), .B(P1_DATAO_REG_10__SCAN_IN), .S(n10671), .Z(
        P1_U3565) );
  MUX2_X1 U10923 ( .A(n10011), .B(P1_DATAO_REG_9__SCAN_IN), .S(n10671), .Z(
        P1_U3564) );
  MUX2_X1 U10924 ( .A(n10012), .B(P1_DATAO_REG_8__SCAN_IN), .S(n10671), .Z(
        P1_U3563) );
  MUX2_X1 U10925 ( .A(n10841), .B(P1_DATAO_REG_7__SCAN_IN), .S(n10671), .Z(
        P1_U3562) );
  MUX2_X1 U10926 ( .A(n10013), .B(P1_DATAO_REG_6__SCAN_IN), .S(n10671), .Z(
        P1_U3561) );
  MUX2_X1 U10927 ( .A(n10844), .B(P1_DATAO_REG_5__SCAN_IN), .S(n10671), .Z(
        P1_U3560) );
  MUX2_X1 U10928 ( .A(n10014), .B(P1_DATAO_REG_4__SCAN_IN), .S(n10671), .Z(
        P1_U3559) );
  MUX2_X1 U10929 ( .A(n10015), .B(P1_DATAO_REG_3__SCAN_IN), .S(n10671), .Z(
        P1_U3558) );
  MUX2_X1 U10930 ( .A(n6949), .B(P1_DATAO_REG_2__SCAN_IN), .S(n10671), .Z(
        P1_U3557) );
  MUX2_X1 U10931 ( .A(n7107), .B(P1_DATAO_REG_1__SCAN_IN), .S(n10671), .Z(
        P1_U3556) );
  MUX2_X1 U10932 ( .A(n6910), .B(P1_DATAO_REG_0__SCAN_IN), .S(n10671), .Z(
        P1_U3555) );
  NOR2_X1 U10933 ( .A1(n10691), .A2(n10016), .ZN(n10017) );
  AOI211_X1 U10934 ( .C1(n10664), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n10018), .B(
        n10017), .ZN(n10028) );
  AOI211_X1 U10935 ( .C1(n10021), .C2(n10020), .A(n10019), .B(n10665), .ZN(
        n10022) );
  INV_X1 U10936 ( .A(n10022), .ZN(n10027) );
  OAI211_X1 U10937 ( .C1(n10025), .C2(n10024), .A(n10677), .B(n10023), .ZN(
        n10026) );
  NAND3_X1 U10938 ( .A1(n10028), .A2(n10027), .A3(n10026), .ZN(P1_U3244) );
  NAND2_X1 U10939 ( .A1(n10664), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n10030) );
  OAI211_X1 U10940 ( .C1(n10047), .C2(n10691), .A(n10030), .B(n10029), .ZN(
        n10039) );
  INV_X1 U10941 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10032) );
  AOI211_X1 U10942 ( .C1(n10033), .C2(n10032), .A(n10041), .B(n10665), .ZN(
        n10038) );
  OAI21_X1 U10943 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n10035), .A(n10034), 
        .ZN(n10046) );
  XNOR2_X1 U10944 ( .A(n10047), .B(n10046), .ZN(n10036) );
  NOR2_X1 U10945 ( .A1(n8278), .A2(n10036), .ZN(n10048) );
  AOI211_X1 U10946 ( .C1(n8278), .C2(n10036), .A(n10048), .B(n10694), .ZN(
        n10037) );
  OR3_X1 U10947 ( .A1(n10039), .A2(n10038), .A3(n10037), .ZN(P1_U3256) );
  NOR2_X1 U10948 ( .A1(n10040), .A2(n10047), .ZN(n10042) );
  NAND2_X1 U10949 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n10066), .ZN(n10043) );
  OAI21_X1 U10950 ( .B1(n10066), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10043), 
        .ZN(n10044) );
  NOR2_X1 U10951 ( .A1(n10045), .A2(n10044), .ZN(n10059) );
  AOI211_X1 U10952 ( .C1(n10045), .C2(n10044), .A(n10059), .B(n10665), .ZN(
        n10057) );
  NOR2_X1 U10953 ( .A1(n10047), .A2(n10046), .ZN(n10049) );
  NOR2_X1 U10954 ( .A1(n10049), .A2(n10048), .ZN(n10051) );
  XNOR2_X1 U10955 ( .A(n10066), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10050) );
  NOR2_X1 U10956 ( .A1(n10051), .A2(n10050), .ZN(n10065) );
  AOI211_X1 U10957 ( .C1(n10051), .C2(n10050), .A(n10065), .B(n10694), .ZN(
        n10056) );
  NAND2_X1 U10958 ( .A1(n10664), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n10053) );
  OAI211_X1 U10959 ( .C1(n10054), .C2(n10691), .A(n10053), .B(n10052), .ZN(
        n10055) );
  OR3_X1 U10960 ( .A1(n10057), .A2(n10056), .A3(n10055), .ZN(P1_U3257) );
  INV_X1 U10961 ( .A(n10058), .ZN(n10064) );
  AOI21_X1 U10962 ( .B1(n10066), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10059), 
        .ZN(n10062) );
  NAND2_X1 U10963 ( .A1(n10078), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n10060) );
  OAI21_X1 U10964 ( .B1(n10078), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10060), 
        .ZN(n10061) );
  NOR2_X1 U10965 ( .A1(n10062), .A2(n10061), .ZN(n10077) );
  AOI211_X1 U10966 ( .C1(n10062), .C2(n10061), .A(n10077), .B(n10665), .ZN(
        n10063) );
  AOI211_X1 U10967 ( .C1(n10078), .C2(n10662), .A(n10064), .B(n10063), .ZN(
        n10071) );
  AOI21_X1 U10968 ( .B1(n10066), .B2(P1_REG1_REG_16__SCAN_IN), .A(n10065), 
        .ZN(n10068) );
  XNOR2_X1 U10969 ( .A(n10078), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n10067) );
  NOR2_X1 U10970 ( .A1(n10068), .A2(n10067), .ZN(n10072) );
  AOI211_X1 U10971 ( .C1(n10068), .C2(n10067), .A(n10072), .B(n10694), .ZN(
        n10069) );
  AOI21_X1 U10972 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n10664), .A(n10069), 
        .ZN(n10070) );
  NAND2_X1 U10973 ( .A1(n10071), .A2(n10070), .ZN(P1_U3258) );
  AOI21_X1 U10974 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n10078), .A(n10072), 
        .ZN(n10578) );
  AOI22_X1 U10975 ( .A1(n10586), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n10074), 
        .B2(n10073), .ZN(n10577) );
  NAND2_X1 U10976 ( .A1(n10578), .A2(n10577), .ZN(n10576) );
  OAI21_X1 U10977 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n10586), .A(n10576), 
        .ZN(n10076) );
  XNOR2_X1 U10978 ( .A(n10730), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n10075) );
  XNOR2_X1 U10979 ( .A(n10076), .B(n10075), .ZN(n10084) );
  AOI21_X1 U10980 ( .B1(n10078), .B2(P1_REG2_REG_17__SCAN_IN), .A(n10077), 
        .ZN(n10583) );
  INV_X1 U10981 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10080) );
  NOR2_X1 U10982 ( .A1(n10586), .A2(n10080), .ZN(n10079) );
  AOI21_X1 U10983 ( .B1(n10586), .B2(n10080), .A(n10079), .ZN(n10582) );
  NOR2_X1 U10984 ( .A1(n10583), .A2(n10582), .ZN(n10581) );
  OAI21_X1 U10985 ( .B1(n10691), .B2(n10229), .A(n10081), .ZN(n10082) );
  OAI21_X1 U10986 ( .B1(n10084), .B2(n10694), .A(n10083), .ZN(P1_U3260) );
  XNOR2_X1 U10987 ( .A(n10085), .B(n10322), .ZN(n10320) );
  NAND2_X1 U10988 ( .A1(n10320), .A2(n10932), .ZN(n10088) );
  AOI21_X1 U10989 ( .B1(n10296), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10086), 
        .ZN(n10087) );
  OAI211_X1 U10990 ( .C1(n10322), .C2(n10935), .A(n10088), .B(n10087), .ZN(
        P1_U3261) );
  XNOR2_X1 U10991 ( .A(n10089), .B(n5184), .ZN(n10337) );
  INV_X1 U10992 ( .A(n10117), .ZN(n10092) );
  INV_X1 U10993 ( .A(n10090), .ZN(n10091) );
  AOI21_X1 U10994 ( .B1(n10333), .B2(n10092), .A(n10091), .ZN(n10334) );
  INV_X1 U10995 ( .A(n10093), .ZN(n10094) );
  AOI22_X1 U10996 ( .A1(n10296), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10094), 
        .B2(n10724), .ZN(n10095) );
  OAI21_X1 U10997 ( .B1(n10096), .B2(n10935), .A(n10095), .ZN(n10106) );
  NAND2_X1 U10998 ( .A1(n10108), .A2(n10097), .ZN(n10099) );
  XNOR2_X1 U10999 ( .A(n10099), .B(n10098), .ZN(n10100) );
  AND2_X1 U11000 ( .A1(n10135), .A2(n10843), .ZN(n10101) );
  AOI21_X1 U11001 ( .B1(n10102), .B2(n10842), .A(n10101), .ZN(n10103) );
  AOI211_X1 U11002 ( .C1(n10932), .C2(n10334), .A(n10106), .B(n10105), .ZN(
        n10107) );
  OAI21_X1 U11003 ( .B1(n10337), .B2(n10300), .A(n10107), .ZN(P1_U3264) );
  OAI21_X1 U11004 ( .B1(n10112), .B2(n10109), .A(n10108), .ZN(n10116) );
  OAI22_X1 U11005 ( .A1(n10111), .A2(n10917), .B1(n10110), .B2(n10915), .ZN(
        n10115) );
  XNOR2_X1 U11006 ( .A(n10113), .B(n10112), .ZN(n10342) );
  NOR2_X1 U11007 ( .A1(n10342), .A2(n10923), .ZN(n10114) );
  AOI211_X1 U11008 ( .C1(n10920), .C2(n10116), .A(n10115), .B(n10114), .ZN(
        n10341) );
  AOI21_X1 U11009 ( .B1(n10338), .B2(n10125), .A(n10117), .ZN(n10339) );
  AOI22_X1 U11010 ( .A1(n10296), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n10118), 
        .B2(n10724), .ZN(n10119) );
  OAI21_X1 U11011 ( .B1(n10120), .B2(n10935), .A(n10119), .ZN(n10122) );
  NOR2_X1 U11012 ( .A1(n10342), .A2(n10264), .ZN(n10121) );
  AOI211_X1 U11013 ( .C1(n10339), .C2(n10932), .A(n10122), .B(n10121), .ZN(
        n10123) );
  OAI21_X1 U11014 ( .B1(n10341), .B2(n10296), .A(n10123), .ZN(P1_U3265) );
  XNOR2_X1 U11015 ( .A(n10124), .B(n10134), .ZN(n10347) );
  INV_X1 U11016 ( .A(n10146), .ZN(n10127) );
  INV_X1 U11017 ( .A(n10125), .ZN(n10126) );
  AOI21_X1 U11018 ( .B1(n10343), .B2(n10127), .A(n10126), .ZN(n10344) );
  INV_X1 U11019 ( .A(n10128), .ZN(n10129) );
  AOI22_X1 U11020 ( .A1(n10296), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10129), 
        .B2(n10724), .ZN(n10130) );
  OAI21_X1 U11021 ( .B1(n10131), .B2(n10935), .A(n10130), .ZN(n10138) );
  OAI21_X1 U11022 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(n10136) );
  AOI222_X1 U11023 ( .A1(n10920), .A2(n10136), .B1(n10135), .B2(n10842), .C1(
        n10164), .C2(n10843), .ZN(n10346) );
  NOR2_X1 U11024 ( .A1(n10346), .A2(n10296), .ZN(n10137) );
  AOI211_X1 U11025 ( .C1(n10344), .C2(n10932), .A(n10138), .B(n10137), .ZN(
        n10139) );
  OAI21_X1 U11026 ( .B1(n10347), .B2(n10300), .A(n10139), .ZN(P1_U3266) );
  XNOR2_X1 U11027 ( .A(n10140), .B(n10143), .ZN(n10352) );
  NOR2_X1 U11028 ( .A1(n5316), .A2(n10935), .ZN(n10150) );
  OAI21_X1 U11029 ( .B1(n10143), .B2(n10142), .A(n10141), .ZN(n10145) );
  AOI222_X1 U11030 ( .A1(n10920), .A2(n10145), .B1(n10144), .B2(n10842), .C1(
        n10180), .C2(n10843), .ZN(n10351) );
  AOI211_X1 U11031 ( .C1(n10349), .C2(n10155), .A(n11043), .B(n10146), .ZN(
        n10348) );
  AOI22_X1 U11032 ( .A1(n10348), .A2(n10229), .B1(n10724), .B2(n10147), .ZN(
        n10148) );
  AOI21_X1 U11033 ( .B1(n10351), .B2(n10148), .A(n10296), .ZN(n10149) );
  AOI211_X1 U11034 ( .C1(n10296), .C2(P1_REG2_REG_24__SCAN_IN), .A(n10150), 
        .B(n10149), .ZN(n10151) );
  OAI21_X1 U11035 ( .B1(n10352), .B2(n10300), .A(n10151), .ZN(P1_U3267) );
  INV_X1 U11036 ( .A(n10152), .ZN(n10153) );
  AOI21_X1 U11037 ( .B1(n10163), .B2(n10154), .A(n10153), .ZN(n10357) );
  INV_X1 U11038 ( .A(n10155), .ZN(n10156) );
  AOI21_X1 U11039 ( .B1(n10353), .B2(n5320), .A(n10156), .ZN(n10354) );
  INV_X1 U11040 ( .A(n10157), .ZN(n10158) );
  AOI22_X1 U11041 ( .A1(n10296), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n10158), 
        .B2(n10724), .ZN(n10159) );
  OAI21_X1 U11042 ( .B1(n10160), .B2(n10935), .A(n10159), .ZN(n10167) );
  OAI21_X1 U11043 ( .B1(n10163), .B2(n10162), .A(n10161), .ZN(n10165) );
  AOI222_X1 U11044 ( .A1(n10920), .A2(n10165), .B1(n10164), .B2(n10842), .C1(
        n10192), .C2(n10843), .ZN(n10356) );
  NOR2_X1 U11045 ( .A1(n10356), .A2(n10296), .ZN(n10166) );
  AOI211_X1 U11046 ( .C1(n10354), .C2(n10932), .A(n10167), .B(n10166), .ZN(
        n10168) );
  OAI21_X1 U11047 ( .B1(n10357), .B2(n10300), .A(n10168), .ZN(P1_U3268) );
  XNOR2_X1 U11048 ( .A(n10170), .B(n10169), .ZN(n10362) );
  AOI21_X1 U11049 ( .B1(n10358), .B2(n10194), .A(n10171), .ZN(n10359) );
  INV_X1 U11050 ( .A(n10358), .ZN(n10175) );
  INV_X1 U11051 ( .A(n10172), .ZN(n10173) );
  AOI22_X1 U11052 ( .A1(n10296), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n10173), 
        .B2(n10724), .ZN(n10174) );
  OAI21_X1 U11053 ( .B1(n10175), .B2(n10935), .A(n10174), .ZN(n10183) );
  OAI21_X1 U11054 ( .B1(n10178), .B2(n10177), .A(n10176), .ZN(n10181) );
  AOI222_X1 U11055 ( .A1(n10920), .A2(n10181), .B1(n10180), .B2(n10842), .C1(
        n10179), .C2(n10843), .ZN(n10361) );
  NOR2_X1 U11056 ( .A1(n10361), .A2(n10296), .ZN(n10182) );
  AOI211_X1 U11057 ( .C1(n10359), .C2(n10932), .A(n10183), .B(n10182), .ZN(
        n10184) );
  OAI21_X1 U11058 ( .B1(n10300), .B2(n10362), .A(n10184), .ZN(P1_U3269) );
  INV_X1 U11059 ( .A(n10185), .ZN(n10187) );
  OAI21_X1 U11060 ( .B1(n10187), .B2(n5444), .A(n10186), .ZN(n10367) );
  NOR2_X1 U11061 ( .A1(n10188), .A2(n10935), .ZN(n10200) );
  OAI21_X1 U11062 ( .B1(n10191), .B2(n10190), .A(n10189), .ZN(n10193) );
  AOI222_X1 U11063 ( .A1(n10920), .A2(n10193), .B1(n10192), .B2(n10842), .C1(
        n10224), .C2(n10843), .ZN(n10366) );
  INV_X1 U11064 ( .A(n10211), .ZN(n10196) );
  INV_X1 U11065 ( .A(n10194), .ZN(n10195) );
  AOI211_X1 U11066 ( .C1(n10364), .C2(n10196), .A(n11043), .B(n10195), .ZN(
        n10363) );
  AOI22_X1 U11067 ( .A1(n10363), .A2(n10229), .B1(n10724), .B2(n10197), .ZN(
        n10198) );
  AOI21_X1 U11068 ( .B1(n10366), .B2(n10198), .A(n10296), .ZN(n10199) );
  AOI211_X1 U11069 ( .C1(n10296), .C2(P1_REG2_REG_21__SCAN_IN), .A(n10200), 
        .B(n10199), .ZN(n10201) );
  OAI21_X1 U11070 ( .B1(n10300), .B2(n10367), .A(n10201), .ZN(P1_U3270) );
  OAI21_X1 U11071 ( .B1(n10206), .B2(n10203), .A(n10202), .ZN(n10210) );
  OAI22_X1 U11072 ( .A1(n10205), .A2(n10917), .B1(n10204), .B2(n10915), .ZN(
        n10209) );
  XNOR2_X1 U11073 ( .A(n10207), .B(n10206), .ZN(n10372) );
  NOR2_X1 U11074 ( .A1(n10372), .A2(n10923), .ZN(n10208) );
  AOI211_X1 U11075 ( .C1(n10920), .C2(n10210), .A(n10209), .B(n10208), .ZN(
        n10371) );
  AOI21_X1 U11076 ( .B1(n10368), .B2(n10226), .A(n10211), .ZN(n10369) );
  INV_X1 U11077 ( .A(n10368), .ZN(n10215) );
  INV_X1 U11078 ( .A(n10212), .ZN(n10213) );
  AOI22_X1 U11079 ( .A1(n10296), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10213), 
        .B2(n10724), .ZN(n10214) );
  OAI21_X1 U11080 ( .B1(n10215), .B2(n10935), .A(n10214), .ZN(n10217) );
  NOR2_X1 U11081 ( .A1(n10372), .A2(n10264), .ZN(n10216) );
  AOI211_X1 U11082 ( .C1(n10369), .C2(n10932), .A(n10217), .B(n10216), .ZN(
        n10218) );
  OAI21_X1 U11083 ( .B1(n10371), .B2(n10296), .A(n10218), .ZN(P1_U3271) );
  XOR2_X1 U11084 ( .A(n10222), .B(n10219), .Z(n10377) );
  OAI21_X1 U11085 ( .B1(n10222), .B2(n10221), .A(n10220), .ZN(n10225) );
  AOI222_X1 U11086 ( .A1(n10920), .A2(n10225), .B1(n10224), .B2(n10842), .C1(
        n10223), .C2(n10843), .ZN(n10376) );
  INV_X1 U11087 ( .A(n10236), .ZN(n10228) );
  INV_X1 U11088 ( .A(n10226), .ZN(n10227) );
  AOI211_X1 U11089 ( .C1(n10374), .C2(n10228), .A(n11043), .B(n10227), .ZN(
        n10373) );
  NAND2_X1 U11090 ( .A1(n10373), .A2(n10229), .ZN(n10230) );
  OAI211_X1 U11091 ( .C1(n10937), .C2(n10231), .A(n10376), .B(n10230), .ZN(
        n10232) );
  NAND2_X1 U11092 ( .A1(n10232), .A2(n10942), .ZN(n10234) );
  AOI22_X1 U11093 ( .A1(n10374), .A2(n10317), .B1(P1_REG2_REG_19__SCAN_IN), 
        .B2(n10296), .ZN(n10233) );
  OAI211_X1 U11094 ( .C1(n10377), .C2(n10300), .A(n10234), .B(n10233), .ZN(
        P1_U3272) );
  XNOR2_X1 U11095 ( .A(n10235), .B(n10241), .ZN(n10382) );
  AOI21_X1 U11096 ( .B1(n10378), .B2(n10257), .A(n10236), .ZN(n10379) );
  INV_X1 U11097 ( .A(n10237), .ZN(n10238) );
  AOI22_X1 U11098 ( .A1(n10296), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10238), 
        .B2(n10724), .ZN(n10239) );
  OAI21_X1 U11099 ( .B1(n10240), .B2(n10935), .A(n10239), .ZN(n10246) );
  XNOR2_X1 U11100 ( .A(n10242), .B(n10241), .ZN(n10244) );
  AOI222_X1 U11101 ( .A1(n10920), .A2(n10244), .B1(n10243), .B2(n10842), .C1(
        n10277), .C2(n10843), .ZN(n10381) );
  NOR2_X1 U11102 ( .A1(n10381), .A2(n10296), .ZN(n10245) );
  AOI211_X1 U11103 ( .C1(n10379), .C2(n10932), .A(n10246), .B(n10245), .ZN(
        n10247) );
  OAI21_X1 U11104 ( .B1(n10300), .B2(n10382), .A(n10247), .ZN(P1_U3273) );
  XNOR2_X1 U11105 ( .A(n10249), .B(n10248), .ZN(n10256) );
  OAI22_X1 U11106 ( .A1(n10251), .A2(n10917), .B1(n10250), .B2(n10915), .ZN(
        n10255) );
  XNOR2_X1 U11107 ( .A(n10253), .B(n10252), .ZN(n10387) );
  NOR2_X1 U11108 ( .A1(n10387), .A2(n10923), .ZN(n10254) );
  AOI211_X1 U11109 ( .C1(n10920), .C2(n10256), .A(n10255), .B(n10254), .ZN(
        n10386) );
  INV_X1 U11110 ( .A(n10269), .ZN(n10259) );
  INV_X1 U11111 ( .A(n10257), .ZN(n10258) );
  AOI21_X1 U11112 ( .B1(n10383), .B2(n10259), .A(n10258), .ZN(n10384) );
  INV_X1 U11113 ( .A(n10260), .ZN(n10261) );
  AOI22_X1 U11114 ( .A1(n10296), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n10261), 
        .B2(n10724), .ZN(n10262) );
  OAI21_X1 U11115 ( .B1(n10263), .B2(n10935), .A(n10262), .ZN(n10266) );
  NOR2_X1 U11116 ( .A1(n10387), .A2(n10264), .ZN(n10265) );
  AOI211_X1 U11117 ( .C1(n10384), .C2(n10932), .A(n10266), .B(n10265), .ZN(
        n10267) );
  OAI21_X1 U11118 ( .B1(n10386), .B2(n10296), .A(n10267), .ZN(P1_U3274) );
  XNOR2_X1 U11119 ( .A(n10268), .B(n10274), .ZN(n10392) );
  AOI211_X1 U11120 ( .C1(n10389), .C2(n10285), .A(n11043), .B(n10269), .ZN(
        n10388) );
  INV_X1 U11121 ( .A(n10389), .ZN(n10273) );
  INV_X1 U11122 ( .A(n10270), .ZN(n10271) );
  AOI22_X1 U11123 ( .A1(n10296), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10271), 
        .B2(n10724), .ZN(n10272) );
  OAI21_X1 U11124 ( .B1(n10273), .B2(n10935), .A(n10272), .ZN(n10280) );
  XNOR2_X1 U11125 ( .A(n10275), .B(n10274), .ZN(n10278) );
  AOI222_X1 U11126 ( .A1(n10920), .A2(n10278), .B1(n10277), .B2(n10842), .C1(
        n10276), .C2(n10843), .ZN(n10391) );
  NOR2_X1 U11127 ( .A1(n10391), .A2(n10296), .ZN(n10279) );
  AOI211_X1 U11128 ( .C1(n10388), .C2(n10281), .A(n10280), .B(n10279), .ZN(
        n10282) );
  OAI21_X1 U11129 ( .B1(n10300), .B2(n10392), .A(n10282), .ZN(P1_U3275) );
  XNOR2_X1 U11130 ( .A(n10283), .B(n10292), .ZN(n10397) );
  INV_X1 U11131 ( .A(n10284), .ZN(n10312) );
  INV_X1 U11132 ( .A(n10285), .ZN(n10286) );
  AOI21_X1 U11133 ( .B1(n10393), .B2(n10312), .A(n10286), .ZN(n10394) );
  INV_X1 U11134 ( .A(n10287), .ZN(n10288) );
  AOI22_X1 U11135 ( .A1(n10296), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10288), 
        .B2(n10724), .ZN(n10289) );
  OAI21_X1 U11136 ( .B1(n10290), .B2(n10935), .A(n10289), .ZN(n10298) );
  XOR2_X1 U11137 ( .A(n10292), .B(n10291), .Z(n10295) );
  AOI222_X1 U11138 ( .A1(n10920), .A2(n10295), .B1(n10294), .B2(n10842), .C1(
        n10293), .C2(n10843), .ZN(n10396) );
  NOR2_X1 U11139 ( .A1(n10396), .A2(n10296), .ZN(n10297) );
  AOI211_X1 U11140 ( .C1(n10394), .C2(n10932), .A(n10298), .B(n10297), .ZN(
        n10299) );
  OAI21_X1 U11141 ( .B1(n10300), .B2(n10397), .A(n10299), .ZN(P1_U3276) );
  INV_X1 U11142 ( .A(n10307), .ZN(n10301) );
  XNOR2_X1 U11143 ( .A(n10302), .B(n10301), .ZN(n10306) );
  OAI22_X1 U11144 ( .A1(n10304), .A2(n10917), .B1(n10303), .B2(n10915), .ZN(
        n10305) );
  AOI21_X1 U11145 ( .B1(n10306), .B2(n10920), .A(n10305), .ZN(n11020) );
  XOR2_X1 U11146 ( .A(n10308), .B(n10307), .Z(n11025) );
  NAND2_X1 U11147 ( .A1(n11025), .A2(n10309), .ZN(n10319) );
  OAI22_X1 U11148 ( .A1(n10942), .A2(n7273), .B1(n10310), .B2(n10937), .ZN(
        n10315) );
  OAI211_X1 U11149 ( .C1(n11022), .C2(n5324), .A(n10312), .B(n10711), .ZN(
        n11019) );
  NOR2_X1 U11150 ( .A1(n11019), .A2(n10313), .ZN(n10314) );
  AOI211_X1 U11151 ( .C1(n10317), .C2(n10316), .A(n10315), .B(n10314), .ZN(
        n10318) );
  OAI211_X1 U11152 ( .C1(n10296), .C2(n11020), .A(n10319), .B(n10318), .ZN(
        P1_U3277) );
  NAND2_X1 U11153 ( .A1(n10320), .A2(n10711), .ZN(n10321) );
  OAI211_X1 U11154 ( .C1(n10322), .C2(n11021), .A(n10321), .B(n11042), .ZN(
        n10418) );
  MUX2_X1 U11155 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10418), .S(n11050), .Z(
        P1_U3554) );
  AOI22_X1 U11156 ( .A1(n10329), .A2(n10711), .B1(n11048), .B2(n10328), .ZN(
        n10330) );
  OAI211_X1 U11157 ( .C1(n10707), .C2(n10332), .A(n10331), .B(n10330), .ZN(
        n10419) );
  MUX2_X1 U11158 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10419), .S(n11050), .Z(
        P1_U3551) );
  AOI22_X1 U11159 ( .A1(n10334), .A2(n10711), .B1(n11048), .B2(n10333), .ZN(
        n10335) );
  OAI211_X1 U11160 ( .C1(n10415), .C2(n10337), .A(n10336), .B(n10335), .ZN(
        n10420) );
  MUX2_X1 U11161 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10420), .S(n11050), .Z(
        P1_U3550) );
  AOI22_X1 U11162 ( .A1(n10339), .A2(n10711), .B1(n11048), .B2(n10338), .ZN(
        n10340) );
  OAI211_X1 U11163 ( .C1(n10342), .C2(n10707), .A(n10341), .B(n10340), .ZN(
        n10421) );
  MUX2_X1 U11164 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10421), .S(n11050), .Z(
        P1_U3549) );
  AOI22_X1 U11165 ( .A1(n10344), .A2(n10711), .B1(n11048), .B2(n10343), .ZN(
        n10345) );
  OAI211_X1 U11166 ( .C1(n10415), .C2(n10347), .A(n10346), .B(n10345), .ZN(
        n10422) );
  MUX2_X1 U11167 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10422), .S(n11050), .Z(
        P1_U3548) );
  AOI21_X1 U11168 ( .B1(n11048), .B2(n10349), .A(n10348), .ZN(n10350) );
  OAI211_X1 U11169 ( .C1(n10415), .C2(n10352), .A(n10351), .B(n10350), .ZN(
        n10423) );
  MUX2_X1 U11170 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10423), .S(n11050), .Z(
        P1_U3547) );
  AOI22_X1 U11171 ( .A1(n10354), .A2(n10711), .B1(n11048), .B2(n10353), .ZN(
        n10355) );
  OAI211_X1 U11172 ( .C1(n10357), .C2(n10415), .A(n10356), .B(n10355), .ZN(
        n10424) );
  MUX2_X1 U11173 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10424), .S(n11050), .Z(
        P1_U3546) );
  AOI22_X1 U11174 ( .A1(n10359), .A2(n10711), .B1(n11048), .B2(n10358), .ZN(
        n10360) );
  OAI211_X1 U11175 ( .C1(n10415), .C2(n10362), .A(n10361), .B(n10360), .ZN(
        n10425) );
  MUX2_X1 U11176 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10425), .S(n11050), .Z(
        P1_U3545) );
  AOI21_X1 U11177 ( .B1(n11048), .B2(n10364), .A(n10363), .ZN(n10365) );
  OAI211_X1 U11178 ( .C1(n10415), .C2(n10367), .A(n10366), .B(n10365), .ZN(
        n10426) );
  MUX2_X1 U11179 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10426), .S(n11050), .Z(
        P1_U3544) );
  AOI22_X1 U11180 ( .A1(n10369), .A2(n10711), .B1(n11048), .B2(n10368), .ZN(
        n10370) );
  OAI211_X1 U11181 ( .C1(n10372), .C2(n10707), .A(n10371), .B(n10370), .ZN(
        n10427) );
  MUX2_X1 U11182 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10427), .S(n11050), .Z(
        P1_U3543) );
  AOI21_X1 U11183 ( .B1(n11048), .B2(n10374), .A(n10373), .ZN(n10375) );
  OAI211_X1 U11184 ( .C1(n10377), .C2(n10415), .A(n10376), .B(n10375), .ZN(
        n10428) );
  MUX2_X1 U11185 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10428), .S(n11050), .Z(
        P1_U3542) );
  AOI22_X1 U11186 ( .A1(n10379), .A2(n10711), .B1(n11048), .B2(n10378), .ZN(
        n10380) );
  OAI211_X1 U11187 ( .C1(n10415), .C2(n10382), .A(n10381), .B(n10380), .ZN(
        n10429) );
  MUX2_X1 U11188 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10429), .S(n11050), .Z(
        P1_U3541) );
  AOI22_X1 U11189 ( .A1(n10384), .A2(n10711), .B1(n11048), .B2(n10383), .ZN(
        n10385) );
  OAI211_X1 U11190 ( .C1(n10707), .C2(n10387), .A(n10386), .B(n10385), .ZN(
        n10430) );
  MUX2_X1 U11191 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10430), .S(n11050), .Z(
        P1_U3540) );
  AOI21_X1 U11192 ( .B1(n11048), .B2(n10389), .A(n10388), .ZN(n10390) );
  OAI211_X1 U11193 ( .C1(n10392), .C2(n10415), .A(n10391), .B(n10390), .ZN(
        n10431) );
  MUX2_X1 U11194 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10431), .S(n11050), .Z(
        P1_U3539) );
  AOI22_X1 U11195 ( .A1(n10394), .A2(n10711), .B1(n11048), .B2(n10393), .ZN(
        n10395) );
  OAI211_X1 U11196 ( .C1(n10397), .C2(n10415), .A(n10396), .B(n10395), .ZN(
        n10432) );
  MUX2_X1 U11197 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10432), .S(n11050), .Z(
        P1_U3538) );
  INV_X1 U11198 ( .A(n10415), .ZN(n11024) );
  INV_X1 U11199 ( .A(n10398), .ZN(n10400) );
  OAI21_X1 U11200 ( .B1(n10400), .B2(n11021), .A(n10399), .ZN(n10401) );
  OR2_X1 U11201 ( .A1(n10402), .A2(n10401), .ZN(n10403) );
  AOI21_X1 U11202 ( .B1(n10404), .B2(n11024), .A(n10403), .ZN(n10434) );
  MUX2_X1 U11203 ( .A(n10434), .B(n7761), .S(n11049), .Z(n10405) );
  INV_X1 U11204 ( .A(n10405), .ZN(P1_U3536) );
  AOI22_X1 U11205 ( .A1(n10407), .A2(n10711), .B1(n11048), .B2(n10406), .ZN(
        n10408) );
  OAI211_X1 U11206 ( .C1(n10410), .C2(n10707), .A(n10409), .B(n10408), .ZN(
        n10436) );
  MUX2_X1 U11207 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10436), .S(n11050), .Z(
        P1_U3534) );
  AOI21_X1 U11208 ( .B1(n11048), .B2(n10412), .A(n10411), .ZN(n10413) );
  OAI211_X1 U11209 ( .C1(n10416), .C2(n10415), .A(n10414), .B(n10413), .ZN(
        n10437) );
  MUX2_X1 U11210 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10437), .S(n11050), .Z(
        P1_U3533) );
  MUX2_X1 U11211 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10417), .S(n11050), .Z(
        P1_U3523) );
  MUX2_X1 U11212 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10418), .S(n11054), .Z(
        P1_U3522) );
  MUX2_X1 U11213 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10419), .S(n11054), .Z(
        P1_U3519) );
  MUX2_X1 U11214 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10420), .S(n11054), .Z(
        P1_U3518) );
  MUX2_X1 U11215 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10421), .S(n11054), .Z(
        P1_U3517) );
  MUX2_X1 U11216 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10422), .S(n11054), .Z(
        P1_U3516) );
  MUX2_X1 U11217 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10423), .S(n11054), .Z(
        P1_U3515) );
  MUX2_X1 U11218 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10424), .S(n11054), .Z(
        P1_U3514) );
  MUX2_X1 U11219 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10425), .S(n11054), .Z(
        P1_U3513) );
  MUX2_X1 U11220 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10426), .S(n11054), .Z(
        P1_U3512) );
  MUX2_X1 U11221 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10427), .S(n11054), .Z(
        P1_U3511) );
  MUX2_X1 U11222 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10428), .S(n11054), .Z(
        P1_U3510) );
  MUX2_X1 U11223 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10429), .S(n11054), .Z(
        P1_U3508) );
  MUX2_X1 U11224 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10430), .S(n11054), .Z(
        P1_U3505) );
  MUX2_X1 U11225 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10431), .S(n11054), .Z(
        P1_U3502) );
  MUX2_X1 U11226 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10432), .S(n11054), .Z(
        P1_U3499) );
  INV_X1 U11227 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10433) );
  MUX2_X1 U11228 ( .A(n10434), .B(n10433), .S(n11051), .Z(n10435) );
  INV_X1 U11229 ( .A(n10435), .ZN(P1_U3493) );
  MUX2_X1 U11230 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10436), .S(n11054), .Z(
        P1_U3487) );
  MUX2_X1 U11231 ( .A(P1_REG0_REG_10__SCAN_IN), .B(n10437), .S(n11054), .Z(
        P1_U3484) );
  INV_X1 U11232 ( .A(n10438), .ZN(n10440) );
  NOR4_X1 U11233 ( .A1(n10440), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), 
        .A4(n10439), .ZN(n10441) );
  AOI21_X1 U11234 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n10442), .A(n10441), 
        .ZN(n10443) );
  OAI21_X1 U11235 ( .B1(n10444), .B2(n10461), .A(n10443), .ZN(P1_U3322) );
  OAI222_X1 U11236 ( .A1(P1_U3084), .A2(n10447), .B1(n10461), .B2(n10446), 
        .C1(n10445), .C2(n10454), .ZN(P1_U3324) );
  OAI222_X1 U11237 ( .A1(n10512), .A2(P1_U3084), .B1(n10461), .B2(n10449), 
        .C1(n10448), .C2(n10454), .ZN(P1_U3325) );
  NAND2_X1 U11238 ( .A1(n10451), .A2(n10450), .ZN(n10453) );
  OAI211_X1 U11239 ( .C1(n10454), .C2(n7034), .A(n10453), .B(n10452), .ZN(
        P1_U3326) );
  OAI222_X1 U11240 ( .A1(n10457), .A2(P1_U3084), .B1(n10461), .B2(n10456), 
        .C1(n10455), .C2(n10454), .ZN(P1_U3327) );
  INV_X1 U11241 ( .A(n10458), .ZN(n10462) );
  OAI222_X1 U11242 ( .A1(P1_U3084), .A2(n10462), .B1(n10461), .B2(n10460), 
        .C1(n10459), .C2(n10454), .ZN(P1_U3328) );
  MUX2_X1 U11243 ( .A(n10463), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U11244 ( .A(n10467), .ZN(n10466) );
  NOR2_X1 U11245 ( .A1(n10466), .A2(n10464), .ZN(P1_U3321) );
  NOR2_X1 U11246 ( .A1(n10466), .A2(n10465), .ZN(P1_U3320) );
  AND2_X1 U11247 ( .A1(n10467), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3319) );
  AND2_X1 U11248 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10467), .ZN(P1_U3318) );
  AND2_X1 U11249 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10467), .ZN(P1_U3317) );
  AND2_X1 U11250 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10467), .ZN(P1_U3316) );
  AND2_X1 U11251 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10467), .ZN(P1_U3315) );
  AND2_X1 U11252 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10467), .ZN(P1_U3314) );
  AND2_X1 U11253 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10467), .ZN(P1_U3313) );
  AND2_X1 U11254 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10467), .ZN(P1_U3312) );
  AND2_X1 U11255 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10467), .ZN(P1_U3311) );
  AND2_X1 U11256 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10467), .ZN(P1_U3310) );
  AND2_X1 U11257 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10467), .ZN(P1_U3309) );
  AND2_X1 U11258 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10467), .ZN(P1_U3308) );
  AND2_X1 U11259 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10467), .ZN(P1_U3307) );
  AND2_X1 U11260 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10467), .ZN(P1_U3306) );
  AND2_X1 U11261 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10467), .ZN(P1_U3305) );
  AND2_X1 U11262 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10467), .ZN(P1_U3304) );
  AND2_X1 U11263 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10467), .ZN(P1_U3303) );
  AND2_X1 U11264 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10467), .ZN(P1_U3302) );
  AND2_X1 U11265 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10467), .ZN(P1_U3301) );
  AND2_X1 U11266 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10467), .ZN(P1_U3300) );
  AND2_X1 U11267 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10467), .ZN(P1_U3299) );
  AND2_X1 U11268 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10467), .ZN(P1_U3298) );
  AND2_X1 U11269 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10467), .ZN(P1_U3297) );
  AND2_X1 U11270 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10467), .ZN(P1_U3296) );
  AND2_X1 U11271 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10467), .ZN(P1_U3295) );
  AND2_X1 U11272 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10467), .ZN(P1_U3294) );
  AND2_X1 U11273 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10467), .ZN(P1_U3293) );
  AND2_X1 U11274 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10467), .ZN(P1_U3292) );
  NOR2_X1 U11275 ( .A1(n10469), .A2(n10468), .ZN(n10473) );
  INV_X1 U11276 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U11277 ( .A1(n10621), .A2(n10473), .B1(n10472), .B2(n10618), .ZN(
        P2_U3438) );
  AND2_X1 U11278 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10618), .ZN(P2_U3326) );
  AND2_X1 U11279 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10618), .ZN(P2_U3325) );
  AND2_X1 U11280 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10618), .ZN(P2_U3324) );
  AND2_X1 U11281 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10618), .ZN(P2_U3323) );
  AND2_X1 U11282 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10618), .ZN(P2_U3322) );
  AND2_X1 U11283 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10618), .ZN(P2_U3321) );
  AND2_X1 U11284 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10618), .ZN(P2_U3320) );
  AND2_X1 U11285 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10618), .ZN(P2_U3319) );
  AND2_X1 U11286 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10618), .ZN(P2_U3318) );
  AND2_X1 U11287 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10618), .ZN(P2_U3317) );
  AND2_X1 U11288 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10618), .ZN(P2_U3316) );
  AND2_X1 U11289 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10618), .ZN(P2_U3315) );
  AND2_X1 U11290 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10618), .ZN(P2_U3314) );
  AND2_X1 U11291 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10618), .ZN(P2_U3313) );
  AND2_X1 U11292 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10618), .ZN(P2_U3312) );
  AND2_X1 U11293 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10618), .ZN(P2_U3311) );
  AND2_X1 U11294 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10618), .ZN(P2_U3310) );
  AND2_X1 U11295 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10618), .ZN(P2_U3309) );
  AND2_X1 U11296 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10618), .ZN(P2_U3308) );
  AND2_X1 U11297 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10618), .ZN(P2_U3307) );
  AND2_X1 U11298 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10618), .ZN(P2_U3306) );
  AND2_X1 U11299 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10618), .ZN(P2_U3305) );
  AND2_X1 U11300 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10618), .ZN(P2_U3304) );
  AND2_X1 U11301 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10618), .ZN(P2_U3303) );
  AND2_X1 U11302 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10618), .ZN(P2_U3302) );
  AND2_X1 U11303 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10618), .ZN(P2_U3301) );
  AND2_X1 U11304 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10618), .ZN(P2_U3300) );
  AND2_X1 U11305 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10618), .ZN(P2_U3299) );
  AND2_X1 U11306 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10618), .ZN(P2_U3298) );
  AND2_X1 U11307 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10618), .ZN(P2_U3297) );
  XOR2_X1 U11308 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  INV_X1 U11309 ( .A(n10474), .ZN(n10475) );
  NAND2_X1 U11310 ( .A1(n10476), .A2(n10475), .ZN(n10477) );
  XNOR2_X1 U11311 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10477), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11312 ( .A(n10479), .B(n10478), .Z(ADD_1071_U54) );
  XOR2_X1 U11313 ( .A(n10481), .B(n10480), .Z(ADD_1071_U53) );
  XNOR2_X1 U11314 ( .A(n10483), .B(n10482), .ZN(ADD_1071_U52) );
  NOR2_X1 U11315 ( .A1(n10485), .A2(n10484), .ZN(n10486) );
  XOR2_X1 U11316 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10486), .Z(ADD_1071_U51) );
  XOR2_X1 U11317 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10487), .Z(ADD_1071_U50) );
  XOR2_X1 U11318 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10488), .Z(ADD_1071_U49) );
  XOR2_X1 U11319 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10489), .Z(ADD_1071_U48) );
  XOR2_X1 U11320 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10490), .Z(ADD_1071_U47) );
  XOR2_X1 U11321 ( .A(n10492), .B(n10491), .Z(ADD_1071_U63) );
  XOR2_X1 U11322 ( .A(n10494), .B(n10493), .Z(ADD_1071_U62) );
  XNOR2_X1 U11323 ( .A(n10496), .B(n10495), .ZN(ADD_1071_U61) );
  XNOR2_X1 U11324 ( .A(n10498), .B(n10497), .ZN(ADD_1071_U60) );
  XNOR2_X1 U11325 ( .A(n10500), .B(n10499), .ZN(ADD_1071_U59) );
  XNOR2_X1 U11326 ( .A(n10502), .B(n10501), .ZN(ADD_1071_U58) );
  XNOR2_X1 U11327 ( .A(n10504), .B(n10503), .ZN(ADD_1071_U57) );
  XNOR2_X1 U11328 ( .A(n10506), .B(n10505), .ZN(ADD_1071_U56) );
  NOR2_X1 U11329 ( .A1(n10508), .A2(n10507), .ZN(n10509) );
  XOR2_X1 U11330 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10509), .Z(ADD_1071_U55)
         );
  NOR2_X1 U11331 ( .A1(n10669), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10515) );
  NOR2_X1 U11332 ( .A1(n10510), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10511) );
  NOR2_X1 U11333 ( .A1(n10512), .A2(n10511), .ZN(n10673) );
  INV_X1 U11334 ( .A(n10673), .ZN(n10513) );
  NOR2_X1 U11335 ( .A1(n10513), .A2(n10515), .ZN(n10514) );
  MUX2_X1 U11336 ( .A(n10515), .B(n10514), .S(P1_IR_REG_0__SCAN_IN), .Z(n10516) );
  NOR2_X1 U11337 ( .A1(n10673), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10672) );
  OR2_X1 U11338 ( .A1(n10516), .A2(n10672), .ZN(n10518) );
  AOI22_X1 U11339 ( .A1(n10664), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10517) );
  OAI21_X1 U11340 ( .B1(n10519), .B2(n10518), .A(n10517), .ZN(P1_U3241) );
  INV_X1 U11341 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n10531) );
  AOI211_X1 U11342 ( .C1(n10522), .C2(n10521), .A(n10520), .B(n10665), .ZN(
        n10523) );
  AOI211_X1 U11343 ( .C1(n10662), .C2(n10525), .A(n10524), .B(n10523), .ZN(
        n10530) );
  OAI211_X1 U11344 ( .C1(n10528), .C2(n10527), .A(n10677), .B(n10526), .ZN(
        n10529) );
  OAI211_X1 U11345 ( .C1(n10700), .C2(n10531), .A(n10530), .B(n10529), .ZN(
        P1_U3247) );
  INV_X1 U11346 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10544) );
  AOI211_X1 U11347 ( .C1(n10534), .C2(n10533), .A(n10532), .B(n10665), .ZN(
        n10535) );
  AOI211_X1 U11348 ( .C1(n10662), .C2(n10537), .A(n10536), .B(n10535), .ZN(
        n10543) );
  AOI21_X1 U11349 ( .B1(n10540), .B2(n10539), .A(n10538), .ZN(n10541) );
  OR2_X1 U11350 ( .A1(n10541), .A2(n10694), .ZN(n10542) );
  OAI211_X1 U11351 ( .C1(n10700), .C2(n10544), .A(n10543), .B(n10542), .ZN(
        P1_U3250) );
  INV_X1 U11352 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10557) );
  AOI211_X1 U11353 ( .C1(n10547), .C2(n10546), .A(n10545), .B(n10665), .ZN(
        n10548) );
  AOI211_X1 U11354 ( .C1(n10662), .C2(n10550), .A(n10549), .B(n10548), .ZN(
        n10556) );
  AOI21_X1 U11355 ( .B1(n10553), .B2(n10552), .A(n10551), .ZN(n10554) );
  OR2_X1 U11356 ( .A1(n10694), .A2(n10554), .ZN(n10555) );
  OAI211_X1 U11357 ( .C1(n10700), .C2(n10557), .A(n10556), .B(n10555), .ZN(
        P1_U3251) );
  INV_X1 U11358 ( .A(n10563), .ZN(n10558) );
  NOR3_X1 U11359 ( .A1(n10559), .A2(n10565), .A3(n10558), .ZN(n10560) );
  AOI211_X1 U11360 ( .C1(P1_ADDR_REG_11__SCAN_IN), .C2(n10664), .A(n10561), 
        .B(n10560), .ZN(n10575) );
  AOI211_X1 U11361 ( .C1(n10565), .C2(n10564), .A(n10563), .B(n10562), .ZN(
        n10569) );
  NAND3_X1 U11362 ( .A1(n10677), .A2(P1_REG1_REG_11__SCAN_IN), .A3(n10572), 
        .ZN(n10566) );
  NAND2_X1 U11363 ( .A1(n10566), .A2(n10691), .ZN(n10567) );
  AOI22_X1 U11364 ( .A1(n10569), .A2(n10687), .B1(n10568), .B2(n10567), .ZN(
        n10574) );
  OAI211_X1 U11365 ( .C1(n10572), .C2(n10571), .A(n10677), .B(n10570), .ZN(
        n10573) );
  NAND3_X1 U11366 ( .A1(n10575), .A2(n10574), .A3(n10573), .ZN(P1_U3252) );
  OAI21_X1 U11367 ( .B1(n10578), .B2(n10577), .A(n10576), .ZN(n10579) );
  AOI22_X1 U11368 ( .A1(n10579), .A2(n10677), .B1(n10664), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n10588) );
  INV_X1 U11369 ( .A(n10580), .ZN(n10585) );
  AOI211_X1 U11370 ( .C1(n10583), .C2(n10582), .A(n10581), .B(n10665), .ZN(
        n10584) );
  AOI211_X1 U11371 ( .C1(n10586), .C2(n10662), .A(n10585), .B(n10584), .ZN(
        n10587) );
  NAND2_X1 U11372 ( .A1(n10588), .A2(n10587), .ZN(P1_U3259) );
  INV_X1 U11373 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10601) );
  OAI21_X1 U11374 ( .B1(n10591), .B2(n10590), .A(n10589), .ZN(n10595) );
  NOR2_X1 U11375 ( .A1(n10691), .A2(n10592), .ZN(n10593) );
  AOI211_X1 U11376 ( .C1(n10687), .C2(n10595), .A(n10594), .B(n10593), .ZN(
        n10600) );
  OAI211_X1 U11377 ( .C1(n10598), .C2(n10597), .A(n10677), .B(n10596), .ZN(
        n10599) );
  OAI211_X1 U11378 ( .C1(n10700), .C2(n10601), .A(n10600), .B(n10599), .ZN(
        P1_U3246) );
  OAI211_X1 U11379 ( .C1(n10604), .C2(n10603), .A(n10687), .B(n10602), .ZN(
        n10606) );
  NAND2_X1 U11380 ( .A1(P1_U3084), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n10605) );
  OAI211_X1 U11381 ( .C1(n10691), .C2(n10607), .A(n10606), .B(n10605), .ZN(
        n10610) );
  INV_X1 U11382 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10608) );
  NOR2_X1 U11383 ( .A1(n10700), .A2(n10608), .ZN(n10609) );
  NOR2_X1 U11384 ( .A1(n10610), .A2(n10609), .ZN(n10616) );
  NOR2_X1 U11385 ( .A1(n5214), .A2(n10611), .ZN(n10613) );
  OAI211_X1 U11386 ( .C1(n10614), .C2(n10613), .A(n10677), .B(n10612), .ZN(
        n10615) );
  NAND2_X1 U11387 ( .A1(n10616), .A2(n10615), .ZN(P1_U3242) );
  INV_X1 U11388 ( .A(n10617), .ZN(n10620) );
  INV_X1 U11389 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U11390 ( .A1(n10621), .A2(n10620), .B1(n10619), .B2(n10618), .ZN(
        P2_U3437) );
  AOI22_X1 U11391 ( .A1(n10622), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n10656), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10628) );
  OR2_X1 U11392 ( .A1(n10648), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10623) );
  OAI211_X1 U11393 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10624), .A(n10623), .B(
        n10638), .ZN(n10625) );
  INV_X1 U11394 ( .A(n10625), .ZN(n10627) );
  AOI22_X1 U11395 ( .A1(n10647), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10626) );
  OAI221_X1 U11396 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10628), .C1(n10641), .C2(
        n10627), .A(n10626), .ZN(P2_U3245) );
  NAND2_X1 U11397 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n10629) );
  NAND2_X1 U11398 ( .A1(n10630), .A2(n10629), .ZN(n10633) );
  INV_X1 U11399 ( .A(n10631), .ZN(n10632) );
  NAND2_X1 U11400 ( .A1(n10633), .A2(n10632), .ZN(n10634) );
  OR2_X1 U11401 ( .A1(n10648), .A2(n10634), .ZN(n10636) );
  AOI22_X1 U11402 ( .A1(n10647), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n10635) );
  OAI211_X1 U11403 ( .C1(n10638), .C2(n10637), .A(n10636), .B(n10635), .ZN(
        n10639) );
  INV_X1 U11404 ( .A(n10639), .ZN(n10646) );
  NOR2_X1 U11405 ( .A1(n10641), .A2(n10640), .ZN(n10644) );
  OAI211_X1 U11406 ( .C1(n10644), .C2(n10643), .A(n10656), .B(n10642), .ZN(
        n10645) );
  NAND2_X1 U11407 ( .A1(n10646), .A2(n10645), .ZN(P2_U3246) );
  AOI22_X1 U11408 ( .A1(n10647), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10661) );
  AOI211_X1 U11409 ( .C1(n10651), .C2(n10650), .A(n10649), .B(n10648), .ZN(
        n10652) );
  AOI21_X1 U11410 ( .B1(n10654), .B2(n10653), .A(n10652), .ZN(n10660) );
  OAI211_X1 U11411 ( .C1(n10658), .C2(n10657), .A(n10656), .B(n10655), .ZN(
        n10659) );
  NAND3_X1 U11412 ( .A1(n10661), .A2(n10660), .A3(n10659), .ZN(P2_U3247) );
  XNOR2_X1 U11413 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI22_X1 U11414 ( .A1(n10664), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(n10663), 
        .B2(n10662), .ZN(n10682) );
  AOI211_X1 U11415 ( .C1(n10668), .C2(n10667), .A(n10666), .B(n10665), .ZN(
        n10675) );
  MUX2_X1 U11416 ( .A(n10670), .B(P1_IR_REG_0__SCAN_IN), .S(n10669), .Z(n10674) );
  AOI211_X1 U11417 ( .C1(n10674), .C2(n10673), .A(n10672), .B(n10671), .ZN(
        n10697) );
  AOI211_X1 U11418 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(P1_U3084), .A(n10675), 
        .B(n10697), .ZN(n10681) );
  OAI211_X1 U11419 ( .C1(n10679), .C2(n10678), .A(n10677), .B(n10676), .ZN(
        n10680) );
  NAND3_X1 U11420 ( .A1(n10682), .A2(n10681), .A3(n10680), .ZN(P1_U3243) );
  INV_X1 U11421 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10701) );
  OAI21_X1 U11422 ( .B1(n10685), .B2(n10684), .A(n10683), .ZN(n10686) );
  AND2_X1 U11423 ( .A1(n10687), .A2(n10686), .ZN(n10696) );
  AOI21_X1 U11424 ( .B1(n10690), .B2(n10689), .A(n10688), .ZN(n10693) );
  OAI22_X1 U11425 ( .A1(n10694), .A2(n10693), .B1(n10692), .B2(n10691), .ZN(
        n10695) );
  NOR4_X1 U11426 ( .A1(n10698), .A2(n10697), .A3(n10696), .A4(n10695), .ZN(
        n10699) );
  OAI21_X1 U11427 ( .B1(n10701), .B2(n10700), .A(n10699), .ZN(P1_U3245) );
  AOI21_X1 U11428 ( .B1(n10702), .B2(n10935), .A(n10712), .ZN(n10705) );
  NOR2_X1 U11429 ( .A1(n10703), .A2(n10296), .ZN(n10704) );
  AOI211_X1 U11430 ( .C1(n10296), .C2(P1_REG2_REG_0__SCAN_IN), .A(n10705), .B(
        n10704), .ZN(n10706) );
  OAI21_X1 U11431 ( .B1(n10937), .B2(n6866), .A(n10706), .ZN(P1_U3291) );
  INV_X1 U11432 ( .A(n10707), .ZN(n10926) );
  XNOR2_X1 U11433 ( .A(n10709), .B(n10708), .ZN(n10731) );
  OAI211_X1 U11434 ( .C1(n10713), .C2(n10712), .A(n10711), .B(n10710), .ZN(
        n10729) );
  OAI21_X1 U11435 ( .B1(n10713), .B2(n11021), .A(n10729), .ZN(n10720) );
  XNOR2_X1 U11436 ( .A(n10715), .B(n10714), .ZN(n10717) );
  AOI22_X1 U11437 ( .A1(n10843), .A2(n6910), .B1(n6949), .B2(n10842), .ZN(
        n10716) );
  OAI21_X1 U11438 ( .B1(n10717), .B2(n10848), .A(n10716), .ZN(n10718) );
  AOI21_X1 U11439 ( .B1(n10840), .B2(n10731), .A(n10718), .ZN(n10728) );
  INV_X1 U11440 ( .A(n10728), .ZN(n10719) );
  AOI211_X1 U11441 ( .C1(n10926), .C2(n10731), .A(n10720), .B(n10719), .ZN(
        n10723) );
  AOI22_X1 U11442 ( .A1(n11050), .A2(n10723), .B1(n10721), .B2(n11049), .ZN(
        P1_U3524) );
  INV_X1 U11443 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10722) );
  AOI22_X1 U11444 ( .A1(n11054), .A2(n10723), .B1(n10722), .B2(n11051), .ZN(
        P1_U3457) );
  INV_X1 U11445 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10734) );
  AOI22_X1 U11446 ( .A1(n10726), .A2(n10725), .B1(n10724), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10727) );
  OAI211_X1 U11447 ( .C1(n10730), .C2(n10729), .A(n10728), .B(n10727), .ZN(
        n10732) );
  AOI22_X1 U11448 ( .A1(n10732), .A2(n10942), .B1(n10731), .B2(n10933), .ZN(
        n10733) );
  OAI21_X1 U11449 ( .B1(n10734), .B2(n10942), .A(n10733), .ZN(P1_U3290) );
  INV_X1 U11450 ( .A(n10735), .ZN(n10740) );
  OAI22_X1 U11451 ( .A1(n10737), .A2(n11043), .B1(n10736), .B2(n11021), .ZN(
        n10739) );
  AOI211_X1 U11452 ( .C1(n10926), .C2(n10740), .A(n10739), .B(n10738), .ZN(
        n10742) );
  AOI22_X1 U11453 ( .A1(n11050), .A2(n10742), .B1(n6876), .B2(n11049), .ZN(
        P1_U3525) );
  INV_X1 U11454 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10741) );
  AOI22_X1 U11455 ( .A1(n11054), .A2(n10742), .B1(n10741), .B2(n11051), .ZN(
        P1_U3460) );
  INV_X1 U11456 ( .A(n10743), .ZN(n10984) );
  OAI22_X1 U11457 ( .A1(n10745), .A2(n11030), .B1(n10744), .B2(n11028), .ZN(
        n10747) );
  AOI211_X1 U11458 ( .C1(n10984), .C2(n10748), .A(n10747), .B(n10746), .ZN(
        n10751) );
  AOI22_X1 U11459 ( .A1(n11037), .A2(n10751), .B1(n10749), .B2(n11036), .ZN(
        P2_U3522) );
  INV_X1 U11460 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10750) );
  AOI22_X1 U11461 ( .A1(n11041), .A2(n10751), .B1(n10750), .B2(n11038), .ZN(
        P2_U3457) );
  OAI22_X1 U11462 ( .A1(n10753), .A2(n11043), .B1(n10752), .B2(n11021), .ZN(
        n10754) );
  AOI21_X1 U11463 ( .B1(n10755), .B2(n10926), .A(n10754), .ZN(n10756) );
  AND2_X1 U11464 ( .A1(n10757), .A2(n10756), .ZN(n10759) );
  AOI22_X1 U11465 ( .A1(n11050), .A2(n10759), .B1(n6551), .B2(n11049), .ZN(
        P1_U3526) );
  INV_X1 U11466 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U11467 ( .A1(n11054), .A2(n10759), .B1(n10758), .B2(n11051), .ZN(
        P1_U3463) );
  INV_X1 U11468 ( .A(n10760), .ZN(n10761) );
  AOI21_X1 U11469 ( .B1(n10762), .B2(n10772), .A(n10761), .ZN(n10774) );
  AOI22_X1 U11470 ( .A1(n10765), .A2(n10764), .B1(n10813), .B2(n10763), .ZN(
        n10769) );
  NAND2_X1 U11471 ( .A1(n10767), .A2(n10766), .ZN(n10768) );
  OAI211_X1 U11472 ( .C1(n6650), .C2(n10818), .A(n10769), .B(n10768), .ZN(
        n10770) );
  AOI21_X1 U11473 ( .B1(n10772), .B2(n10771), .A(n10770), .ZN(n10773) );
  OAI21_X1 U11474 ( .B1(n10821), .B2(n10774), .A(n10773), .ZN(P2_U3293) );
  NAND2_X1 U11475 ( .A1(n10780), .A2(n10926), .ZN(n10776) );
  OAI211_X1 U11476 ( .C1(n10777), .C2(n11021), .A(n10776), .B(n10775), .ZN(
        n10779) );
  AOI211_X1 U11477 ( .C1(n10840), .C2(n10780), .A(n10779), .B(n10778), .ZN(
        n10783) );
  AOI22_X1 U11478 ( .A1(n11050), .A2(n10783), .B1(n10781), .B2(n11049), .ZN(
        P1_U3527) );
  INV_X1 U11479 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10782) );
  AOI22_X1 U11480 ( .A1(n11054), .A2(n10783), .B1(n10782), .B2(n11051), .ZN(
        P1_U3466) );
  OAI22_X1 U11481 ( .A1(n10785), .A2(n11030), .B1(n10784), .B2(n11028), .ZN(
        n10787) );
  AOI211_X1 U11482 ( .C1(n11034), .C2(n10788), .A(n10787), .B(n10786), .ZN(
        n10791) );
  AOI22_X1 U11483 ( .A1(n11037), .A2(n10791), .B1(n10789), .B2(n11036), .ZN(
        P2_U3524) );
  INV_X1 U11484 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10790) );
  AOI22_X1 U11485 ( .A1(n11041), .A2(n10791), .B1(n10790), .B2(n11038), .ZN(
        P2_U3463) );
  OAI22_X1 U11486 ( .A1(n10887), .A2(n10794), .B1(n10793), .B2(n10792), .ZN(
        n10807) );
  AOI22_X1 U11487 ( .A1(n10807), .A2(n10955), .B1(P2_REG3_REG_5__SCAN_IN), 
        .B2(P2_U3152), .ZN(n10800) );
  OAI21_X1 U11488 ( .B1(n10797), .B2(n10796), .A(n10795), .ZN(n10798) );
  AOI22_X1 U11489 ( .A1(n10798), .A2(n10964), .B1(n10963), .B2(n10810), .ZN(
        n10799) );
  OAI211_X1 U11490 ( .C1(n10801), .C2(n10968), .A(n10800), .B(n10799), .ZN(
        P2_U3229) );
  INV_X1 U11491 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10820) );
  XNOR2_X1 U11492 ( .A(n10802), .B(n10805), .ZN(n10826) );
  XNOR2_X1 U11493 ( .A(n10803), .B(n10824), .ZN(n10804) );
  NAND2_X1 U11494 ( .A1(n10804), .A2(n10865), .ZN(n10822) );
  XNOR2_X1 U11495 ( .A(n10806), .B(n10805), .ZN(n10809) );
  AOI21_X1 U11496 ( .B1(n10809), .B2(n10808), .A(n10807), .ZN(n10823) );
  AOI22_X1 U11497 ( .A1(n10813), .A2(n10812), .B1(n10811), .B2(n10810), .ZN(
        n10814) );
  OAI211_X1 U11498 ( .C1(n10815), .C2(n10822), .A(n10823), .B(n10814), .ZN(
        n10816) );
  AOI21_X1 U11499 ( .B1(n10817), .B2(n10826), .A(n10816), .ZN(n10819) );
  AOI22_X1 U11500 ( .A1(n10821), .A2(n10820), .B1(n10819), .B2(n10818), .ZN(
        P2_U3291) );
  OAI211_X1 U11501 ( .C1(n10824), .C2(n11028), .A(n10823), .B(n10822), .ZN(
        n10825) );
  AOI21_X1 U11502 ( .B1(n11034), .B2(n10826), .A(n10825), .ZN(n10829) );
  AOI22_X1 U11503 ( .A1(n11037), .A2(n10829), .B1(n10827), .B2(n11036), .ZN(
        P2_U3525) );
  INV_X1 U11504 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10828) );
  AOI22_X1 U11505 ( .A1(n11041), .A2(n10829), .B1(n10828), .B2(n11038), .ZN(
        P2_U3466) );
  OAI21_X1 U11506 ( .B1(n7521), .B2(n10832), .A(n10831), .ZN(n10854) );
  OAI21_X1 U11507 ( .B1(n5314), .B2(n10855), .A(n10834), .ZN(n10852) );
  OAI22_X1 U11508 ( .A1(n10852), .A2(n11043), .B1(n10855), .B2(n11021), .ZN(
        n10849) );
  INV_X1 U11509 ( .A(n10835), .ZN(n10836) );
  XNOR2_X1 U11510 ( .A(n10839), .B(n10838), .ZN(n10847) );
  NAND2_X1 U11511 ( .A1(n10854), .A2(n10840), .ZN(n10846) );
  AOI22_X1 U11512 ( .A1(n10844), .A2(n10843), .B1(n10842), .B2(n10841), .ZN(
        n10845) );
  OAI211_X1 U11513 ( .C1(n10848), .C2(n10847), .A(n10846), .B(n10845), .ZN(
        n10860) );
  AOI211_X1 U11514 ( .C1(n10926), .C2(n10854), .A(n10849), .B(n10860), .ZN(
        n10851) );
  AOI22_X1 U11515 ( .A1(n11050), .A2(n10851), .B1(n7240), .B2(n11049), .ZN(
        P1_U3529) );
  INV_X1 U11516 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U11517 ( .A1(n11054), .A2(n10851), .B1(n10850), .B2(n11051), .ZN(
        P1_U3472) );
  INV_X1 U11518 ( .A(n10852), .ZN(n10853) );
  AOI22_X1 U11519 ( .A1(n10854), .A2(n10933), .B1(n10932), .B2(n10853), .ZN(
        n10862) );
  NOR2_X1 U11520 ( .A1(n10935), .A2(n10855), .ZN(n10859) );
  INV_X1 U11521 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10857) );
  OAI22_X1 U11522 ( .A1(n10942), .A2(n10857), .B1(n10856), .B2(n10937), .ZN(
        n10858) );
  AOI211_X1 U11523 ( .C1(n10860), .C2(n10942), .A(n10859), .B(n10858), .ZN(
        n10861) );
  NAND2_X1 U11524 ( .A1(n10862), .A2(n10861), .ZN(P1_U3285) );
  AOI22_X1 U11525 ( .A1(n10866), .A2(n10865), .B1(n10864), .B2(n10863), .ZN(
        n10870) );
  NAND3_X1 U11526 ( .A1(n10868), .A2(n10867), .A3(n11034), .ZN(n10869) );
  AND3_X1 U11527 ( .A1(n10871), .A2(n10870), .A3(n10869), .ZN(n10874) );
  AOI22_X1 U11528 ( .A1(n11037), .A2(n10874), .B1(n10872), .B2(n11036), .ZN(
        P2_U3526) );
  INV_X1 U11529 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U11530 ( .A1(n11041), .A2(n10874), .B1(n10873), .B2(n11038), .ZN(
        P2_U3469) );
  OAI21_X1 U11531 ( .B1(n10876), .B2(n11021), .A(n10875), .ZN(n10877) );
  AOI21_X1 U11532 ( .B1(n10878), .B2(n10926), .A(n10877), .ZN(n10879) );
  AOI22_X1 U11533 ( .A1(n11050), .A2(n10882), .B1(n7347), .B2(n11049), .ZN(
        P1_U3530) );
  INV_X1 U11534 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U11535 ( .A1(n11054), .A2(n10882), .B1(n10881), .B2(n11051), .ZN(
        P1_U3475) );
  AOI22_X1 U11536 ( .A1(n10884), .A2(n10883), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(P2_U3152), .ZN(n10885) );
  OAI21_X1 U11537 ( .B1(n10887), .B2(n10886), .A(n10885), .ZN(n10894) );
  INV_X1 U11538 ( .A(n10888), .ZN(n10889) );
  AOI211_X1 U11539 ( .C1(n10892), .C2(n10891), .A(n10890), .B(n10889), .ZN(
        n10893) );
  AOI211_X1 U11540 ( .C1(n10963), .C2(n10895), .A(n10894), .B(n10893), .ZN(
        n10896) );
  OAI21_X1 U11541 ( .B1(n10897), .B2(n10968), .A(n10896), .ZN(P2_U3215) );
  OAI22_X1 U11542 ( .A1(n10898), .A2(n11030), .B1(n5151), .B2(n11028), .ZN(
        n10900) );
  AOI211_X1 U11543 ( .C1(n11034), .C2(n10901), .A(n10900), .B(n10899), .ZN(
        n10903) );
  AOI22_X1 U11544 ( .A1(n11037), .A2(n10903), .B1(n6746), .B2(n11036), .ZN(
        P2_U3527) );
  INV_X1 U11545 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U11546 ( .A1(n11041), .A2(n10903), .B1(n10902), .B2(n11038), .ZN(
        P2_U3472) );
  NAND2_X1 U11547 ( .A1(n10905), .A2(n10904), .ZN(n10906) );
  NAND2_X1 U11548 ( .A1(n10906), .A2(n10913), .ZN(n10907) );
  NAND2_X1 U11549 ( .A1(n10908), .A2(n10907), .ZN(n10924) );
  INV_X1 U11550 ( .A(n10924), .ZN(n10934) );
  OAI21_X1 U11551 ( .B1(n10910), .B2(n10936), .A(n10909), .ZN(n10930) );
  OAI22_X1 U11552 ( .A1(n10930), .A2(n11043), .B1(n10936), .B2(n11021), .ZN(
        n10925) );
  NAND2_X1 U11553 ( .A1(n10912), .A2(n10911), .ZN(n10914) );
  XNOR2_X1 U11554 ( .A(n10914), .B(n10913), .ZN(n10921) );
  OAI22_X1 U11555 ( .A1(n10918), .A2(n10917), .B1(n10916), .B2(n10915), .ZN(
        n10919) );
  AOI21_X1 U11556 ( .B1(n10921), .B2(n10920), .A(n10919), .ZN(n10922) );
  OAI21_X1 U11557 ( .B1(n10924), .B2(n10923), .A(n10922), .ZN(n10943) );
  AOI211_X1 U11558 ( .C1(n10926), .C2(n10934), .A(n10925), .B(n10943), .ZN(
        n10929) );
  AOI22_X1 U11559 ( .A1(n11050), .A2(n10929), .B1(n10927), .B2(n11049), .ZN(
        P1_U3531) );
  INV_X1 U11560 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U11561 ( .A1(n11054), .A2(n10929), .B1(n10928), .B2(n11051), .ZN(
        P1_U3478) );
  INV_X1 U11562 ( .A(n10930), .ZN(n10931) );
  AOI22_X1 U11563 ( .A1(n10934), .A2(n10933), .B1(n10932), .B2(n10931), .ZN(
        n10945) );
  NOR2_X1 U11564 ( .A1(n10936), .A2(n10935), .ZN(n10941) );
  INV_X1 U11565 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10939) );
  OAI22_X1 U11566 ( .A1(n10942), .A2(n10939), .B1(n10938), .B2(n10937), .ZN(
        n10940) );
  AOI211_X1 U11567 ( .C1(n10943), .C2(n10942), .A(n10941), .B(n10940), .ZN(
        n10944) );
  NAND2_X1 U11568 ( .A1(n10945), .A2(n10944), .ZN(P1_U3283) );
  NOR2_X1 U11569 ( .A1(n10946), .A2(n11008), .ZN(n10951) );
  OAI21_X1 U11570 ( .B1(n10948), .B2(n11028), .A(n10947), .ZN(n10950) );
  AOI211_X1 U11571 ( .C1(n10951), .C2(n7375), .A(n10950), .B(n10949), .ZN(
        n10953) );
  AOI22_X1 U11572 ( .A1(n11037), .A2(n10953), .B1(n6789), .B2(n11036), .ZN(
        P2_U3528) );
  INV_X1 U11573 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U11574 ( .A1(n11041), .A2(n10953), .B1(n10952), .B2(n11038), .ZN(
        P2_U3475) );
  AOI22_X1 U11575 ( .A1(n10956), .A2(n10955), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(P2_U3152), .ZN(n10967) );
  INV_X1 U11576 ( .A(n10957), .ZN(n10959) );
  NAND2_X1 U11577 ( .A1(n10959), .A2(n10958), .ZN(n10960) );
  XNOR2_X1 U11578 ( .A(n10961), .B(n10960), .ZN(n10965) );
  AOI22_X1 U11579 ( .A1(n10965), .A2(n10964), .B1(n10963), .B2(n10962), .ZN(
        n10966) );
  OAI211_X1 U11580 ( .C1(n10969), .C2(n10968), .A(n10967), .B(n10966), .ZN(
        P2_U3233) );
  OAI22_X1 U11581 ( .A1(n10971), .A2(n11030), .B1(n10970), .B2(n11028), .ZN(
        n10973) );
  AOI211_X1 U11582 ( .C1(n10974), .C2(n11034), .A(n10973), .B(n10972), .ZN(
        n10977) );
  AOI22_X1 U11583 ( .A1(n11037), .A2(n10977), .B1(n10975), .B2(n11036), .ZN(
        P2_U3529) );
  INV_X1 U11584 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10976) );
  AOI22_X1 U11585 ( .A1(n11041), .A2(n10977), .B1(n10976), .B2(n11038), .ZN(
        P2_U3478) );
  INV_X1 U11586 ( .A(n10978), .ZN(n10983) );
  OAI22_X1 U11587 ( .A1(n10980), .A2(n11030), .B1(n10979), .B2(n11028), .ZN(
        n10982) );
  AOI211_X1 U11588 ( .C1(n10984), .C2(n10983), .A(n10982), .B(n10981), .ZN(
        n10986) );
  AOI22_X1 U11589 ( .A1(n11037), .A2(n10986), .B1(n6791), .B2(n11036), .ZN(
        P2_U3530) );
  INV_X1 U11590 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U11591 ( .A1(n11041), .A2(n10986), .B1(n10985), .B2(n11038), .ZN(
        P2_U3481) );
  OAI21_X1 U11592 ( .B1(n10988), .B2(n11028), .A(n10987), .ZN(n10990) );
  AOI211_X1 U11593 ( .C1(n10991), .C2(n11034), .A(n10990), .B(n10989), .ZN(
        n10993) );
  AOI22_X1 U11594 ( .A1(n11037), .A2(n10993), .B1(n6812), .B2(n11036), .ZN(
        P2_U3531) );
  INV_X1 U11595 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10992) );
  AOI22_X1 U11596 ( .A1(n11041), .A2(n10993), .B1(n10992), .B2(n11038), .ZN(
        P2_U3484) );
  OAI211_X1 U11597 ( .C1(n10996), .C2(n11021), .A(n10995), .B(n10994), .ZN(
        n10997) );
  AOI21_X1 U11598 ( .B1(n10998), .B2(n11024), .A(n10997), .ZN(n11000) );
  AOI22_X1 U11599 ( .A1(n11050), .A2(n11000), .B1(n7754), .B2(n11049), .ZN(
        P1_U3535) );
  INV_X1 U11600 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U11601 ( .A1(n11054), .A2(n11000), .B1(n10999), .B2(n11051), .ZN(
        P1_U3490) );
  OAI22_X1 U11602 ( .A1(n11001), .A2(n11030), .B1(n5276), .B2(n11028), .ZN(
        n11003) );
  AOI211_X1 U11603 ( .C1(n11004), .C2(n11034), .A(n11003), .B(n11002), .ZN(
        n11007) );
  AOI22_X1 U11604 ( .A1(n11037), .A2(n11007), .B1(n11005), .B2(n11036), .ZN(
        P2_U3532) );
  INV_X1 U11605 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U11606 ( .A1(n11041), .A2(n11007), .B1(n11006), .B2(n11038), .ZN(
        P2_U3487) );
  NOR2_X1 U11607 ( .A1(n11009), .A2(n11008), .ZN(n11015) );
  OAI22_X1 U11608 ( .A1(n11011), .A2(n11030), .B1(n11010), .B2(n11028), .ZN(
        n11013) );
  AOI211_X1 U11609 ( .C1(n11015), .C2(n11014), .A(n11013), .B(n11012), .ZN(
        n11018) );
  AOI22_X1 U11610 ( .A1(n11037), .A2(n11018), .B1(n11016), .B2(n11036), .ZN(
        P2_U3533) );
  INV_X1 U11611 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U11612 ( .A1(n11041), .A2(n11018), .B1(n11017), .B2(n11038), .ZN(
        P2_U3490) );
  OAI211_X1 U11613 ( .C1(n11022), .C2(n11021), .A(n11020), .B(n11019), .ZN(
        n11023) );
  AOI21_X1 U11614 ( .B1(n11025), .B2(n11024), .A(n11023), .ZN(n11027) );
  AOI22_X1 U11615 ( .A1(n11050), .A2(n11027), .B1(n7267), .B2(n11049), .ZN(
        P1_U3537) );
  INV_X1 U11616 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U11617 ( .A1(n11054), .A2(n11027), .B1(n11026), .B2(n11051), .ZN(
        P1_U3496) );
  OAI22_X1 U11618 ( .A1(n11031), .A2(n11030), .B1(n11029), .B2(n11028), .ZN(
        n11032) );
  AOI211_X1 U11619 ( .C1(n11035), .C2(n11034), .A(n11033), .B(n11032), .ZN(
        n11040) );
  AOI22_X1 U11620 ( .A1(n11037), .A2(n11040), .B1(n7305), .B2(n11036), .ZN(
        P2_U3534) );
  INV_X1 U11621 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n11039) );
  AOI22_X1 U11622 ( .A1(n11041), .A2(n11040), .B1(n11039), .B2(n11038), .ZN(
        P2_U3493) );
  INV_X1 U11623 ( .A(n11042), .ZN(n11046) );
  NOR2_X1 U11624 ( .A1(n11044), .A2(n11043), .ZN(n11045) );
  AOI211_X2 U11625 ( .C1(n11048), .C2(n11047), .A(n11046), .B(n11045), .ZN(
        n11053) );
  AOI22_X1 U11626 ( .A1(n11050), .A2(n11053), .B1(n8489), .B2(n11049), .ZN(
        P1_U3553) );
  INV_X1 U11627 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n11052) );
  AOI22_X1 U11628 ( .A1(n11054), .A2(n11053), .B1(n11052), .B2(n11051), .ZN(
        P1_U3521) );
  XNOR2_X1 U11629 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  CLKBUF_X1 U5296 ( .A(n6303), .Z(n6427) );
  CLKBUF_X1 U5369 ( .A(n5830), .Z(n6128) );
endmodule

