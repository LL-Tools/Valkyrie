

module b14_C_gen_AntiSAT_k_128_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, 
        U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, 
        U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, 
        U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, 
        U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, 
        U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, 
        U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, 
        U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, 
        U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, 
        U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, 
        U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, 
        U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, 
        U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, 
        U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, 
        U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, 
        U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, 
        U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, 
        U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, 
        U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, 
        U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, 
        U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, 
        U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, 
        U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, 
        U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, 
        U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704;

  NAND2_X1 U2287 ( .A1(n2394), .A2(n2393), .ZN(n3875) );
  INV_X1 U2288 ( .A(n2355), .ZN(n2609) );
  BUF_X1 U2289 ( .A(n4359), .Z(n2048) );
  XNOR2_X1 U2290 ( .A(n2371), .B(IR_REG_2__SCAN_IN), .ZN(n4359) );
  CLKBUF_X1 U2291 ( .A(n3839), .Z(n2045) );
  NOR2_X1 U2292 ( .A1(n2892), .A2(n4181), .ZN(n3839) );
  INV_X1 U2293 ( .A(n3697), .ZN(n3702) );
  INV_X2 U2294 ( .A(n3428), .ZN(n2771) );
  OAI21_X1 U2295 ( .B1(n2354), .B2(n2152), .A(n2151), .ZN(n3029) );
  INV_X1 U2296 ( .A(IR_REG_31__SCAN_IN), .ZN(n2642) );
  NAND2_X1 U2298 ( .A1(n2677), .A2(n2068), .ZN(n2309) );
  XNOR2_X2 U2299 ( .A(n2685), .B(IR_REG_24__SCAN_IN), .ZN(n2688) );
  XNOR2_X2 U2300 ( .A(n2634), .B(n2633), .ZN(n2640) );
  BUF_X1 U2301 ( .A(n2320), .Z(n2046) );
  XNOR2_X2 U2302 ( .A(n2308), .B(IR_REG_30__SCAN_IN), .ZN(n4349) );
  NAND2_X2 U2303 ( .A1(n2309), .A2(IR_REG_31__SCAN_IN), .ZN(n2308) );
  CLKBUF_X1 U2304 ( .A(n4359), .Z(n2047) );
  NAND2_X1 U2305 ( .A1(n3757), .A2(n2288), .ZN(n3797) );
  NAND2_X1 U2306 ( .A1(n3587), .A2(n3586), .ZN(n3585) );
  NAND2_X1 U2307 ( .A1(n3259), .A2(n3258), .ZN(n2178) );
  NAND2_X1 U2308 ( .A1(n2413), .A2(n2412), .ZN(n3060) );
  NAND2_X1 U2309 ( .A1(n2993), .A2(n2397), .ZN(n3049) );
  AND3_X1 U2310 ( .A1(n2096), .A2(n2930), .A3(n2931), .ZN(n2958) );
  AND2_X1 U2311 ( .A1(n2940), .A2(n2361), .ZN(n2372) );
  NOR2_X1 U2312 ( .A1(n2825), .A2(n2124), .ZN(n2840) );
  NAND2_X2 U2313 ( .A1(n3515), .A2(n3519), .ZN(n2650) );
  INV_X1 U2314 ( .A(n3876), .ZN(n3041) );
  CLKBUF_X2 U2315 ( .A(n2904), .Z(n3877) );
  NAND4_X2 U2316 ( .A1(n2377), .A2(n2376), .A3(n2375), .A4(n2374), .ZN(n3876)
         );
  INV_X1 U2317 ( .A(n3708), .ZN(n2903) );
  OR2_X1 U2318 ( .A1(n3470), .A2(n2764), .ZN(n2908) );
  NAND2_X1 U2319 ( .A1(n2119), .A2(n4350), .ZN(n2365) );
  NAND2_X1 U2320 ( .A1(n2684), .A2(IR_REG_31__SCAN_IN), .ZN(n2685) );
  AOI21_X1 U2321 ( .B1(n2683), .B2(IR_REG_31__SCAN_IN), .A(n2094), .ZN(n2093)
         );
  MUX2_X1 U2322 ( .A(IR_REG_31__SCAN_IN), .B(n2312), .S(IR_REG_29__SCAN_IN), 
        .Z(n2313) );
  NAND2_X1 U2323 ( .A1(n2560), .A2(IR_REG_31__SCAN_IN), .ZN(n2631) );
  NOR3_X1 U2324 ( .A1(n2679), .A2(IR_REG_25__SCAN_IN), .A3(n2114), .ZN(n2320)
         );
  AND2_X1 U2325 ( .A1(n2551), .A2(n2065), .ZN(n2627) );
  AND4_X1 U2326 ( .A1(n2335), .A2(n2299), .A3(n2298), .A4(n2297), .ZN(n2300)
         );
  NOR2_X1 U2327 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2107)
         );
  NOR2_X1 U2328 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2106)
         );
  INV_X1 U2329 ( .A(IR_REG_3__SCAN_IN), .ZN(n2379) );
  NOR2_X1 U2330 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2297)
         );
  NOR2_X1 U2331 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2299)
         );
  NOR2_X1 U2332 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2298)
         );
  OAI22_X2 U2333 ( .A1(n3060), .A2(n2425), .B1(n3084), .B2(n3873), .ZN(n3106)
         );
  NOR2_X1 U2334 ( .A1(n2583), .A2(n2073), .ZN(n2252) );
  NAND2_X1 U2335 ( .A1(n2627), .A2(n2626), .ZN(n2635) );
  NOR2_X1 U2336 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2626)
         );
  INV_X1 U2337 ( .A(IR_REG_21__SCAN_IN), .ZN(n2628) );
  INV_X1 U2338 ( .A(n2296), .ZN(n2232) );
  NAND2_X1 U2339 ( .A1(n2183), .A2(n2076), .ZN(n3614) );
  OR2_X1 U2340 ( .A1(n3399), .A2(n2184), .ZN(n2183) );
  NAND2_X1 U2341 ( .A1(n2181), .A2(n3599), .ZN(n2180) );
  OR2_X1 U2342 ( .A1(n4350), .A2(n4349), .ZN(n2364) );
  NAND2_X1 U2343 ( .A1(n3898), .A2(n2138), .ZN(n2137) );
  NAND2_X1 U2344 ( .A1(n2048), .A2(REG2_REG_2__SCAN_IN), .ZN(n2138) );
  NAND2_X1 U2345 ( .A1(n2274), .A2(n2502), .ZN(n2273) );
  OR2_X1 U2346 ( .A1(n3605), .A2(n3400), .ZN(n2502) );
  NAND2_X1 U2347 ( .A1(n3490), .A2(n2492), .ZN(n2274) );
  NAND2_X1 U2348 ( .A1(n3523), .A2(n3520), .ZN(n2651) );
  INV_X1 U2349 ( .A(n2908), .ZN(n2856) );
  NOR2_X1 U2350 ( .A1(n2706), .A2(n2762), .ZN(n2689) );
  OR2_X1 U2351 ( .A1(n2617), .A2(n3715), .ZN(n2644) );
  NAND2_X1 U2352 ( .A1(n2575), .A2(n2574), .ZN(n2585) );
  OAI22_X1 U2353 ( .A1(n3602), .A2(n2964), .B1(n3702), .B2(n3606), .ZN(n3612)
         );
  NAND2_X1 U2354 ( .A1(n3354), .A2(n3353), .ZN(n3399) );
  OR2_X1 U2355 ( .A1(n2889), .A2(n4352), .ZN(n2909) );
  OR2_X1 U2356 ( .A1(n2871), .A2(n2062), .ZN(n2142) );
  NAND2_X1 U2357 ( .A1(n2794), .A2(n2141), .ZN(n2144) );
  NOR2_X1 U2358 ( .A1(n2796), .A2(n2876), .ZN(n2141) );
  AND2_X1 U2359 ( .A1(n2262), .A2(n3501), .ZN(n2258) );
  NOR2_X1 U2360 ( .A1(n4005), .A2(n3994), .ZN(n2263) );
  AOI21_X1 U2361 ( .B1(n2080), .B2(n2249), .A(n2248), .ZN(n2247) );
  NOR2_X1 U2362 ( .A1(n4225), .A2(n4027), .ZN(n2248) );
  AND2_X1 U2363 ( .A1(n3291), .A2(n3293), .ZN(n3490) );
  INV_X1 U2364 ( .A(n2651), .ZN(n3480) );
  MUX2_X1 U2365 ( .A(n2726), .B(n2725), .S(IR_REG_28__SCAN_IN), .Z(n2354) );
  NAND2_X1 U2366 ( .A1(n2165), .A2(n2169), .ZN(n2723) );
  NAND2_X1 U2367 ( .A1(n4017), .A2(n2171), .ZN(n2165) );
  OR2_X1 U2368 ( .A1(n4009), .A2(n4199), .ZN(n3988) );
  AND4_X1 U2369 ( .A1(n2486), .A2(n2485), .A3(n2484), .A4(n2483), .ZN(n3356)
         );
  INV_X1 U2370 ( .A(n4169), .ZN(n4070) );
  INV_X1 U2371 ( .A(n2277), .ZN(n2114) );
  INV_X1 U2372 ( .A(n2635), .ZN(n2636) );
  INV_X1 U2373 ( .A(n4216), .ZN(n4200) );
  INV_X1 U2374 ( .A(n4199), .ZN(n3994) );
  NOR2_X1 U2375 ( .A1(n3434), .A2(n3437), .ZN(n2175) );
  INV_X1 U2376 ( .A(n3401), .ZN(n3173) );
  INV_X1 U2377 ( .A(n3817), .ZN(n2214) );
  NOR2_X1 U2378 ( .A1(n3638), .A2(n2227), .ZN(n2226) );
  INV_X1 U2379 ( .A(n3635), .ZN(n2227) );
  NAND2_X1 U2380 ( .A1(n2123), .A2(n2122), .ZN(n3937) );
  NAND2_X1 U2381 ( .A1(n4354), .A2(REG1_REG_7__SCAN_IN), .ZN(n2122) );
  OR2_X1 U2382 ( .A1(n2840), .A2(n2839), .ZN(n2123) );
  AND2_X1 U2383 ( .A1(n3436), .A2(n2175), .ZN(n2174) );
  NAND2_X1 U2384 ( .A1(n4155), .A2(n4137), .ZN(n2561) );
  NOR2_X1 U2385 ( .A1(n2241), .A2(n2238), .ZN(n2237) );
  INV_X1 U2386 ( .A(n2244), .ZN(n2238) );
  INV_X1 U2387 ( .A(n4261), .ZN(n2245) );
  AND2_X1 U2388 ( .A1(n2052), .A2(n2541), .ZN(n2244) );
  INV_X1 U2389 ( .A(n3525), .ZN(n2104) );
  AND2_X1 U2390 ( .A1(n2171), .A2(n3422), .ZN(n2168) );
  OAI21_X1 U2391 ( .B1(n2169), .B2(n2167), .A(n3425), .ZN(n2166) );
  INV_X1 U2392 ( .A(n3422), .ZN(n2167) );
  INV_X1 U2393 ( .A(n3859), .ZN(n2163) );
  INV_X1 U2394 ( .A(n4058), .ZN(n2709) );
  NAND2_X1 U2395 ( .A1(n4115), .A2(n4072), .ZN(n2130) );
  NOR2_X1 U2396 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2301)
         );
  NOR2_X1 U2397 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2302)
         );
  INV_X1 U2398 ( .A(IR_REG_23__SCAN_IN), .ZN(n2691) );
  INV_X1 U2399 ( .A(IR_REG_19__SCAN_IN), .ZN(n2630) );
  INV_X1 U2400 ( .A(IR_REG_18__SCAN_IN), .ZN(n2092) );
  NOR2_X1 U2401 ( .A1(n2511), .A2(IR_REG_13__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U2402 ( .A1(n2107), .A2(n2106), .ZN(n2296) );
  INV_X1 U2403 ( .A(IR_REG_2__SCAN_IN), .ZN(n2293) );
  AND2_X1 U2404 ( .A1(n3172), .A2(n3170), .ZN(n2195) );
  NAND2_X1 U2405 ( .A1(n3169), .A2(n3168), .ZN(n2194) );
  NAND2_X1 U2406 ( .A1(n2089), .A2(n3847), .ZN(n3630) );
  NOR2_X1 U2407 ( .A1(n2222), .A2(n2218), .ZN(n2217) );
  INV_X1 U2408 ( .A(n3780), .ZN(n2218) );
  INV_X1 U2409 ( .A(n2223), .ZN(n2222) );
  NOR2_X1 U2410 ( .A1(n3825), .A2(n2224), .ZN(n2223) );
  INV_X1 U2411 ( .A(n3637), .ZN(n2224) );
  INV_X1 U2412 ( .A(n2226), .ZN(n2221) );
  OR2_X1 U2413 ( .A1(n2365), .A2(n2801), .ZN(n2366) );
  OR2_X1 U2414 ( .A1(n3397), .A2(n3398), .ZN(n2182) );
  AND2_X1 U2415 ( .A1(n3397), .A2(n3398), .ZN(n2186) );
  OR2_X1 U2416 ( .A1(n3647), .A2(n3646), .ZN(n3648) );
  OAI22_X1 U2417 ( .A1(n2925), .A2(n3708), .B1(n3707), .B2(n2927), .ZN(n2926)
         );
  NAND2_X1 U2418 ( .A1(n2928), .A2(n2913), .ZN(n2930) );
  AOI21_X1 U2419 ( .B1(n3910), .B2(REG2_REG_3__SCAN_IN), .A(n2061), .ZN(n2793)
         );
  AND2_X1 U2420 ( .A1(n2142), .A2(n2063), .ZN(n2829) );
  XNOR2_X1 U2421 ( .A(n3937), .B(n2121), .ZN(n3940) );
  NAND2_X1 U2422 ( .A1(n4396), .A2(REG2_REG_12__SCAN_IN), .ZN(n4395) );
  NAND2_X1 U2423 ( .A1(n2140), .A2(n2139), .ZN(n3926) );
  OR2_X1 U2424 ( .A1(n4488), .A2(REG2_REG_13__SCAN_IN), .ZN(n2139) );
  OR2_X1 U2425 ( .A1(n4408), .A2(n4404), .ZN(n2140) );
  XNOR2_X1 U2426 ( .A(n3929), .B(n3954), .ZN(n4439) );
  NAND2_X1 U2427 ( .A1(n4431), .A2(n3953), .ZN(n3955) );
  NOR2_X1 U2428 ( .A1(n4426), .A2(n2147), .ZN(n3929) );
  AND2_X1 U2429 ( .A1(n4485), .A2(REG2_REG_15__SCAN_IN), .ZN(n2147) );
  NAND2_X1 U2430 ( .A1(n4439), .A2(n2530), .ZN(n4438) );
  NAND2_X1 U2431 ( .A1(n4447), .A2(n2158), .ZN(n2157) );
  NAND2_X1 U2432 ( .A1(n4483), .A2(n2547), .ZN(n2158) );
  NOR2_X1 U2433 ( .A1(n2157), .A2(n4458), .ZN(n4457) );
  NAND2_X1 U2434 ( .A1(n2260), .A2(n2266), .ZN(n2259) );
  INV_X1 U2435 ( .A(n2264), .ZN(n2260) );
  AOI21_X1 U2436 ( .B1(n2721), .B2(n2263), .A(n2072), .ZN(n2262) );
  NAND2_X1 U2437 ( .A1(n2262), .A2(n2257), .ZN(n2256) );
  NAND2_X1 U2438 ( .A1(n2264), .A2(n3501), .ZN(n2257) );
  INV_X1 U2439 ( .A(n2252), .ZN(n2251) );
  AOI21_X1 U2440 ( .B1(n2252), .B2(n2250), .A(n2079), .ZN(n2249) );
  INV_X1 U2441 ( .A(n2584), .ZN(n2250) );
  NAND2_X1 U2442 ( .A1(n3585), .A2(n2244), .ZN(n2243) );
  NAND2_X1 U2443 ( .A1(n2052), .A2(n2071), .ZN(n2242) );
  NAND2_X1 U2444 ( .A1(n3366), .A2(n3508), .ZN(n3595) );
  NAND2_X1 U2445 ( .A1(n3595), .A2(n3594), .ZN(n3593) );
  INV_X1 U2446 ( .A(n2272), .ZN(n2271) );
  OAI21_X1 U2447 ( .B1(n2273), .B2(n2492), .A(n2284), .ZN(n2272) );
  OAI21_X1 U2448 ( .B1(n3094), .B2(n2655), .A(n3536), .ZN(n3204) );
  OAI21_X1 U2449 ( .B1(n3050), .B2(n3048), .A(n3503), .ZN(n3061) );
  AND2_X1 U2450 ( .A1(n3526), .A2(n3530), .ZN(n3482) );
  NAND4_X1 U2451 ( .A1(n2352), .A2(n2351), .A3(n2350), .A4(n2349), .ZN(n2904)
         );
  OR2_X1 U2452 ( .A1(n2364), .A2(n2346), .ZN(n2352) );
  NAND2_X1 U2453 ( .A1(n2355), .A2(REG3_REG_1__SCAN_IN), .ZN(n2351) );
  OR2_X1 U2454 ( .A1(n2365), .A2(n2348), .ZN(n2349) );
  NAND2_X1 U2455 ( .A1(n2108), .A2(n3480), .ZN(n2743) );
  NAND2_X1 U2456 ( .A1(n2109), .A2(n3519), .ZN(n2108) );
  INV_X1 U2457 ( .A(n2944), .ZN(n2109) );
  AND2_X1 U2458 ( .A1(n2624), .A2(n2623), .ZN(n4202) );
  NOR2_X1 U2459 ( .A1(n2050), .A2(n4221), .ZN(n4036) );
  AND4_X1 U2460 ( .A1(n2510), .A2(n2509), .A3(n2508), .A4(n2507), .ZN(n3602)
         );
  NAND2_X1 U2461 ( .A1(n2674), .A2(n3456), .ZN(n4169) );
  NAND2_X1 U2462 ( .A1(n2100), .A2(n3480), .ZN(n2741) );
  INV_X1 U2463 ( .A(n2372), .ZN(n2100) );
  AND2_X1 U2464 ( .A1(n2848), .A2(n2640), .ZN(n4276) );
  NAND2_X1 U2465 ( .A1(n3721), .A2(n2687), .ZN(n2776) );
  NAND2_X1 U2466 ( .A1(n2858), .A2(n2778), .ZN(n2895) );
  INV_X1 U2467 ( .A(IR_REG_29__SCAN_IN), .ZN(n2307) );
  AND2_X1 U2468 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2324)
         );
  NAND2_X1 U2469 ( .A1(n2323), .A2(n2322), .ZN(n2726) );
  INV_X1 U2470 ( .A(n2046), .ZN(n2323) );
  XNOR2_X1 U2471 ( .A(n2638), .B(n2637), .ZN(n2889) );
  INV_X1 U2472 ( .A(IR_REG_22__SCAN_IN), .ZN(n2637) );
  NAND2_X1 U2473 ( .A1(n2551), .A2(n2325), .ZN(n2559) );
  NOR2_X1 U2474 ( .A1(n2404), .A2(n2296), .ZN(n2333) );
  INV_X1 U2475 ( .A(IR_REG_7__SCAN_IN), .ZN(n2434) );
  AND2_X1 U2476 ( .A1(n2605), .A2(n2604), .ZN(n4216) );
  NAND2_X1 U2477 ( .A1(n2099), .A2(n3835), .ZN(n2098) );
  NAND2_X1 U2478 ( .A1(n2207), .A2(n2204), .ZN(n2099) );
  XNOR2_X1 U2479 ( .A(n3705), .B(n3706), .ZN(n3736) );
  NAND2_X1 U2480 ( .A1(n2178), .A2(n2058), .ZN(n3354) );
  NAND2_X1 U2481 ( .A1(n2196), .A2(n2199), .ZN(n3714) );
  INV_X1 U2482 ( .A(n2200), .ZN(n2199) );
  NAND2_X1 U2483 ( .A1(n3691), .A2(n2197), .ZN(n2196) );
  OAI22_X1 U2484 ( .A1(n3736), .A2(n2201), .B1(n3705), .B2(n3706), .ZN(n2200)
         );
  AND2_X1 U2485 ( .A1(n2591), .A2(n2590), .ZN(n4054) );
  INV_X1 U2486 ( .A(n3875), .ZN(n3120) );
  AND2_X1 U2487 ( .A1(n2582), .A2(n2581), .ZN(n3819) );
  INV_X1 U2488 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4635) );
  OR2_X1 U2489 ( .A1(n2921), .A2(n2898), .ZN(n3840) );
  AND4_X1 U2490 ( .A1(n2403), .A2(n2402), .A3(n2401), .A4(n2400), .ZN(n3133)
         );
  INV_X1 U2491 ( .A(n4038), .ZN(n4225) );
  OR2_X1 U2492 ( .A1(n2921), .A2(n2920), .ZN(n3851) );
  INV_X1 U2493 ( .A(n3819), .ZN(n4222) );
  OAI21_X1 U2494 ( .B1(n2148), .B2(n2789), .A(n2125), .ZN(n3883) );
  NAND2_X1 U2495 ( .A1(n2148), .A2(n2789), .ZN(n2125) );
  NAND2_X1 U2496 ( .A1(n3883), .A2(n2790), .ZN(n3895) );
  XNOR2_X1 U2497 ( .A(n3955), .B(n3954), .ZN(n4442) );
  NOR2_X1 U2498 ( .A1(n4442), .A2(REG1_REG_16__SCAN_IN), .ZN(n4443) );
  AOI21_X1 U2499 ( .B1(n4460), .B2(ADDR_REG_18__SCAN_IN), .A(n4459), .ZN(n2154) );
  NOR2_X1 U2500 ( .A1(n4453), .A2(n3958), .ZN(n4463) );
  NAND2_X1 U2501 ( .A1(n4463), .A2(n4464), .ZN(n4461) );
  INV_X1 U2502 ( .A(n4457), .ZN(n2156) );
  AOI21_X1 U2503 ( .B1(n2157), .B2(n4458), .A(n4456), .ZN(n2155) );
  AND2_X1 U2504 ( .A1(n2797), .A2(n2795), .ZN(n4462) );
  OAI21_X1 U2505 ( .B1(n2710), .B2(n3729), .A(n2054), .ZN(n3725) );
  INV_X1 U2506 ( .A(n2263), .ZN(n2261) );
  NAND2_X1 U2507 ( .A1(n2173), .A2(n2171), .ZN(n3987) );
  NAND2_X1 U2508 ( .A1(n2111), .A2(n3985), .ZN(n3986) );
  NAND2_X1 U2509 ( .A1(n2173), .A2(n3563), .ZN(n2111) );
  NAND2_X1 U2510 ( .A1(n3232), .A2(n2492), .ZN(n3308) );
  OR2_X1 U2511 ( .A1(n2365), .A2(n2357), .ZN(n2358) );
  OR2_X1 U2512 ( .A1(n2364), .A2(n2356), .ZN(n2360) );
  INV_X1 U2513 ( .A(n4468), .ZN(n4181) );
  NAND2_X1 U2514 ( .A1(n2731), .A2(n2161), .ZN(n2160) );
  NAND2_X1 U2515 ( .A1(n3427), .A2(n4282), .ZN(n2161) );
  OR2_X1 U2516 ( .A1(n3725), .A2(n4294), .ZN(n2716) );
  NAND2_X1 U2517 ( .A1(n2056), .A2(n4512), .ZN(n2159) );
  OR2_X1 U2518 ( .A1(n3725), .A2(n4347), .ZN(n2712) );
  INV_X1 U2519 ( .A(n3933), .ZN(n4482) );
  INV_X1 U2520 ( .A(n2182), .ZN(n2181) );
  OR2_X1 U2521 ( .A1(n2185), .A2(n2186), .ZN(n2184) );
  INV_X1 U2522 ( .A(n3599), .ZN(n2185) );
  INV_X1 U2523 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U2524 ( .A1(n2721), .A2(n2265), .ZN(n2264) );
  INV_X1 U2525 ( .A(n2616), .ZN(n2265) );
  NOR2_X1 U2526 ( .A1(n2544), .A2(n4626), .ZN(n2328) );
  AND2_X1 U2527 ( .A1(n2328), .A2(REG3_REG_18__SCAN_IN), .ZN(n2327) );
  INV_X1 U2528 ( .A(n2470), .ZN(n2290) );
  INV_X1 U2529 ( .A(n2373), .ZN(n2270) );
  OR2_X1 U2530 ( .A1(n2720), .A2(n3427), .ZN(n2136) );
  AOI21_X1 U2531 ( .B1(n2171), .B2(n3557), .A(n2170), .ZN(n2169) );
  INV_X1 U2532 ( .A(n3424), .ZN(n2170) );
  NAND2_X1 U2533 ( .A1(n3593), .A2(n2175), .ZN(n4125) );
  NOR2_X1 U2534 ( .A1(n3369), .A2(n4283), .ZN(n2127) );
  NAND2_X1 U2535 ( .A1(n3152), .A2(n2075), .ZN(n2126) );
  NAND2_X1 U2536 ( .A1(n3121), .A2(n3042), .ZN(n2133) );
  OR2_X1 U2537 ( .A1(n2776), .A2(n2703), .ZN(n2747) );
  AND2_X1 U2538 ( .A1(n2321), .A2(n2306), .ZN(n2277) );
  AND2_X1 U2539 ( .A1(n2277), .A2(n2310), .ZN(n2276) );
  INV_X1 U2540 ( .A(IR_REG_27__SCAN_IN), .ZN(n2321) );
  INV_X1 U2541 ( .A(IR_REG_17__SCAN_IN), .ZN(n2325) );
  OR2_X1 U2542 ( .A1(n3622), .A2(n3621), .ZN(n3743) );
  AOI21_X1 U2543 ( .B1(n2209), .B2(n2213), .A(n2077), .ZN(n2208) );
  NAND2_X1 U2544 ( .A1(n2205), .A2(n3835), .ZN(n2201) );
  NOR2_X1 U2545 ( .A1(n2202), .A2(n2198), .ZN(n2197) );
  OR2_X1 U2546 ( .A1(n3736), .A2(n2203), .ZN(n2202) );
  INV_X1 U2547 ( .A(n3835), .ZN(n2203) );
  INV_X1 U2548 ( .A(n3186), .ZN(n2191) );
  NAND2_X1 U2549 ( .A1(n2193), .A2(n3186), .ZN(n2192) );
  INV_X1 U2550 ( .A(n2195), .ZN(n2193) );
  NAND2_X1 U2551 ( .A1(n3698), .A2(n2948), .ZN(n2091) );
  INV_X1 U2552 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4665) );
  OR2_X1 U2553 ( .A1(n2532), .A2(n2531), .ZN(n2544) );
  NAND2_X1 U2554 ( .A1(n3634), .A2(n3633), .ZN(n3635) );
  INV_X1 U2555 ( .A(n3632), .ZN(n3633) );
  INV_X1 U2556 ( .A(n3631), .ZN(n3634) );
  XOR2_X1 U2557 ( .A(n3261), .B(n3260), .Z(n3258) );
  NAND2_X1 U2558 ( .A1(n3771), .A2(n3770), .ZN(n2215) );
  NAND2_X1 U2559 ( .A1(n3804), .A2(n2212), .ZN(n2211) );
  OR2_X1 U2560 ( .A1(n2564), .A2(n4630), .ZN(n2576) );
  NAND2_X1 U2561 ( .A1(n2228), .A2(n2226), .ZN(n2225) );
  NAND2_X1 U2562 ( .A1(n2339), .A2(REG3_REG_15__SCAN_IN), .ZN(n2532) );
  NAND3_X1 U2563 ( .A1(n2886), .A2(n2885), .A3(n2884), .ZN(n2921) );
  AND4_X1 U2564 ( .A1(n2432), .A2(n2431), .A3(n2430), .A4(n2429), .ZN(n3206)
         );
  XNOR2_X1 U2565 ( .A(n2137), .B(n2804), .ZN(n3910) );
  OR2_X1 U2566 ( .A1(n2871), .A2(n2146), .ZN(n2143) );
  AOI22_X1 U2567 ( .A1(n2831), .A2(REG2_REG_6__SCAN_IN), .B1(n4355), .B2(n2830), .ZN(n2833) );
  AND2_X1 U2568 ( .A1(n3563), .A2(n2172), .ZN(n2171) );
  NAND2_X1 U2569 ( .A1(n2112), .A2(n2673), .ZN(n2173) );
  NAND2_X1 U2570 ( .A1(n4067), .A2(n4094), .ZN(n2234) );
  NOR2_X1 U2571 ( .A1(n4067), .A2(n4094), .ZN(n2235) );
  NAND2_X1 U2572 ( .A1(n2113), .A2(n3554), .ZN(n4084) );
  NAND2_X1 U2573 ( .A1(n3593), .A2(n2074), .ZN(n2113) );
  NAND2_X1 U2574 ( .A1(n3593), .A2(n2174), .ZN(n4102) );
  AOI21_X1 U2575 ( .B1(n4151), .B2(n2240), .A(n2081), .ZN(n2239) );
  NAND2_X1 U2576 ( .A1(n3585), .A2(n2237), .ZN(n2236) );
  INV_X1 U2577 ( .A(n2242), .ZN(n2240) );
  OR2_X1 U2578 ( .A1(n3365), .A2(n3493), .ZN(n3366) );
  NAND2_X1 U2579 ( .A1(n3323), .A2(n2231), .ZN(n3368) );
  NAND2_X1 U2580 ( .A1(n4289), .A2(n3617), .ZN(n2231) );
  OAI21_X1 U2581 ( .B1(n3141), .B2(n3140), .A(n3539), .ZN(n3150) );
  NAND2_X1 U2582 ( .A1(n2118), .A2(n3535), .ZN(n3141) );
  NAND2_X1 U2583 ( .A1(n3204), .A2(n3538), .ZN(n2118) );
  NAND2_X1 U2584 ( .A1(n3061), .A2(n3528), .ZN(n2653) );
  AND2_X1 U2585 ( .A1(n2654), .A2(n3536), .ZN(n3533) );
  NAND2_X1 U2586 ( .A1(n2105), .A2(n3530), .ZN(n3050) );
  NAND2_X1 U2587 ( .A1(n2977), .A2(n2103), .ZN(n2105) );
  NOR2_X1 U2588 ( .A1(n2652), .A2(n2104), .ZN(n2103) );
  NAND2_X1 U2589 ( .A1(n2372), .A2(n2651), .ZN(n2742) );
  INV_X1 U2590 ( .A(n4276), .ZN(n3098) );
  NOR2_X1 U2591 ( .A1(n2650), .A2(n3514), .ZN(n2944) );
  OR2_X1 U2592 ( .A1(n2882), .A2(n2880), .ZN(n2887) );
  OR2_X1 U2593 ( .A1(n2776), .A2(D_REG_1__SCAN_IN), .ZN(n2884) );
  AND2_X1 U2594 ( .A1(n2747), .A2(n2777), .ZN(n2885) );
  AOI21_X1 U2595 ( .B1(n2730), .B2(n4169), .A(n2162), .ZN(n3976) );
  NOR2_X1 U2596 ( .A1(n2164), .A2(n2163), .ZN(n2162) );
  INV_X1 U2597 ( .A(n3968), .ZN(n2164) );
  NOR2_X1 U2598 ( .A1(n3988), .A2(n2135), .ZN(n4194) );
  OR2_X1 U2599 ( .A1(n2136), .A2(n4197), .ZN(n2135) );
  NAND2_X1 U2600 ( .A1(n4023), .A2(n4010), .ZN(n4009) );
  AND2_X1 U2601 ( .A1(n4036), .A2(n4027), .ZN(n4023) );
  INV_X1 U2602 ( .A(n4042), .ZN(n4221) );
  OR3_X1 U2603 ( .A1(n2130), .A2(n4239), .A3(n2709), .ZN(n2129) );
  NAND2_X1 U2604 ( .A1(n3428), .A2(DATAI_23_), .ZN(n4058) );
  NOR3_X1 U2605 ( .A1(n4136), .A2(n4239), .A3(n4105), .ZN(n4088) );
  NOR2_X1 U2606 ( .A1(n4136), .A2(n4105), .ZN(n4113) );
  NAND2_X1 U2607 ( .A1(n4175), .A2(n4159), .ZN(n4158) );
  OR2_X1 U2608 ( .A1(n4158), .A2(n4132), .ZN(n4136) );
  NAND2_X1 U2609 ( .A1(n2127), .A2(n3628), .ZN(n4174) );
  NOR2_X1 U2610 ( .A1(n4174), .A2(n4260), .ZN(n4175) );
  INV_X1 U2611 ( .A(n4186), .ZN(n4260) );
  INV_X1 U2612 ( .A(n2127), .ZN(n3588) );
  NAND2_X1 U2613 ( .A1(n3326), .A2(n3617), .ZN(n3369) );
  NOR2_X1 U2614 ( .A1(n2126), .A2(n3296), .ZN(n3326) );
  NAND2_X1 U2615 ( .A1(n3152), .A2(n2049), .ZN(n3311) );
  INV_X1 U2616 ( .A(n3266), .ZN(n3275) );
  AND2_X1 U2617 ( .A1(n3213), .A2(n3253), .ZN(n3152) );
  INV_X1 U2618 ( .A(n3205), .ZN(n3215) );
  OR2_X1 U2619 ( .A1(n3100), .A2(n3099), .ZN(n3214) );
  NOR2_X1 U2620 ( .A1(n3214), .A2(n3215), .ZN(n3213) );
  NAND2_X1 U2621 ( .A1(n2132), .A2(n2131), .ZN(n3100) );
  INV_X1 U2622 ( .A(n2133), .ZN(n2132) );
  AND3_X1 U2623 ( .A1(n3011), .A2(n2974), .A3(n3134), .ZN(n2131) );
  NOR2_X1 U2624 ( .A1(n2133), .A2(n3002), .ZN(n3065) );
  NAND2_X1 U2625 ( .A1(n2134), .A2(n3042), .ZN(n3054) );
  INV_X1 U2626 ( .A(n2980), .ZN(n3011) );
  INV_X1 U2627 ( .A(n4273), .ZN(n4284) );
  INV_X1 U2628 ( .A(n2749), .ZN(n2886) );
  INV_X1 U2629 ( .A(IR_REG_28__SCAN_IN), .ZN(n2310) );
  NAND2_X1 U2630 ( .A1(n2678), .A2(n2229), .ZN(n2706) );
  AOI21_X1 U2631 ( .B1(n2681), .B2(n2057), .A(n2230), .ZN(n2229) );
  NOR2_X1 U2632 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2230)
         );
  AND4_X1 U2633 ( .A1(n2304), .A2(n2303), .A3(n2302), .A4(n2301), .ZN(n2305)
         );
  NOR2_X1 U2634 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2304)
         );
  NOR2_X1 U2635 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2303)
         );
  NAND2_X1 U2636 ( .A1(n2095), .A2(n2691), .ZN(n2094) );
  NAND2_X1 U2637 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2095) );
  OAI21_X1 U2638 ( .B1(n2683), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2690) );
  XNOR2_X1 U2639 ( .A(n2629), .B(n2628), .ZN(n3470) );
  INV_X1 U2640 ( .A(IR_REG_20__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U2641 ( .A1(n2632), .A2(IR_REG_31__SCAN_IN), .ZN(n2634) );
  OR3_X1 U2642 ( .A1(n2487), .A2(IR_REG_12__SCAN_IN), .A3(n2336), .ZN(n2511)
         );
  CLKBUF_X1 U2643 ( .A(n2404), .Z(n2405) );
  INV_X1 U2644 ( .A(IR_REG_5__SCAN_IN), .ZN(n2407) );
  NOR2_X2 U2645 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2370)
         );
  INV_X1 U2646 ( .A(IR_REG_6__SCAN_IN), .ZN(n4519) );
  OAI21_X1 U2647 ( .B1(n3171), .B2(n2195), .A(n2194), .ZN(n3187) );
  AND4_X1 U2648 ( .A1(n2522), .A2(n2521), .A3(n2520), .A4(n2519), .ZN(n4269)
         );
  NAND2_X1 U2649 ( .A1(n3613), .A2(n3612), .ZN(n2177) );
  NAND2_X1 U2650 ( .A1(n3616), .A2(n3615), .ZN(n2176) );
  CLKBUF_X1 U2651 ( .A(n3757), .Z(n3758) );
  AOI21_X1 U2652 ( .B1(n2221), .B2(n2223), .A(n2220), .ZN(n2219) );
  INV_X1 U2653 ( .A(n3826), .ZN(n2220) );
  XOR2_X1 U2654 ( .A(n3646), .B(n3647), .Z(n3765) );
  AND2_X1 U2655 ( .A1(n2644), .A2(n2618), .ZN(n3726) );
  NOR2_X2 U2656 ( .A1(n2369), .A2(n2283), .ZN(n2925) );
  AND2_X1 U2657 ( .A1(n2355), .A2(REG3_REG_2__SCAN_IN), .ZN(n2283) );
  OR2_X1 U2658 ( .A1(n2364), .A2(n2363), .ZN(n2367) );
  INV_X1 U2659 ( .A(n4090), .ZN(n4244) );
  INV_X1 U2660 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4630) );
  NAND2_X1 U2661 ( .A1(n3804), .A2(n3808), .ZN(n3773) );
  OR2_X1 U2662 ( .A1(n3399), .A2(n2186), .ZN(n2179) );
  INV_X1 U2663 ( .A(n2090), .ZN(n3129) );
  AND2_X1 U2664 ( .A1(n2597), .A2(n2586), .ZN(n4039) );
  AND4_X1 U2665 ( .A1(n2442), .A2(n2441), .A3(n2440), .A4(n2439), .ZN(n3252)
         );
  INV_X1 U2666 ( .A(n3247), .ZN(n3253) );
  AND4_X1 U2667 ( .A1(n2498), .A2(n2497), .A3(n2496), .A4(n2495), .ZN(n3605)
         );
  NAND2_X1 U2668 ( .A1(n2211), .A2(n2215), .ZN(n3816) );
  NAND2_X1 U2669 ( .A1(n2931), .A2(n2930), .ZN(n2097) );
  INV_X1 U2670 ( .A(n2045), .ZN(n3782) );
  INV_X1 U2671 ( .A(n2932), .ZN(n2096) );
  AND3_X1 U2672 ( .A1(n2550), .A2(n2549), .A3(n2548), .ZN(n4274) );
  INV_X1 U2673 ( .A(n3084), .ZN(n3134) );
  INV_X1 U2674 ( .A(n3845), .ZN(n3849) );
  NOR2_X1 U2675 ( .A1(n3702), .A2(n2890), .ZN(n3579) );
  INV_X1 U2676 ( .A(n4352), .ZN(n3963) );
  NAND2_X1 U2677 ( .A1(n2614), .A2(n2613), .ZN(n3861) );
  NAND2_X1 U2678 ( .A1(n2596), .A2(n2595), .ZN(n4038) );
  INV_X1 U2679 ( .A(n4054), .ZN(n4213) );
  OAI211_X1 U2680 ( .C1(n3419), .C2(n4251), .A(n2567), .B(n2566), .ZN(n4241)
         );
  OAI211_X1 U2681 ( .C1(n4161), .C2(n2609), .A(n2332), .B(n2331), .ZN(n4261)
         );
  INV_X1 U2682 ( .A(n4274), .ZN(n4153) );
  INV_X1 U2683 ( .A(n3602), .ZN(n3865) );
  INV_X1 U2684 ( .A(n3605), .ZN(n3866) );
  INV_X1 U2685 ( .A(n3356), .ZN(n3867) );
  INV_X1 U2686 ( .A(n3252), .ZN(n3870) );
  INV_X1 U2687 ( .A(n3206), .ZN(n3871) );
  INV_X1 U2688 ( .A(n3133), .ZN(n3874) );
  AND3_X1 U2689 ( .A1(n2389), .A2(n2388), .A3(n2387), .ZN(n2394) );
  OR2_X1 U2690 ( .A1(n2609), .A2(REG3_REG_3__SCAN_IN), .ZN(n2376) );
  OR2_X1 U2691 ( .A1(n2314), .A2(n3909), .ZN(n2374) );
  NAND2_X1 U2692 ( .A1(n2791), .A2(n2792), .ZN(n3898) );
  NAND2_X1 U2693 ( .A1(n2142), .A2(n2144), .ZN(n2813) );
  NAND2_X1 U2694 ( .A1(n2794), .A2(n4357), .ZN(n2145) );
  AND2_X1 U2695 ( .A1(n2826), .A2(n4355), .ZN(n2124) );
  INV_X1 U2696 ( .A(IR_REG_8__SCAN_IN), .ZN(n2444) );
  INV_X1 U2697 ( .A(n3940), .ZN(n3936) );
  AND2_X1 U2698 ( .A1(n2797), .A2(n3578), .ZN(n4406) );
  NAND2_X1 U2699 ( .A1(n4395), .A2(n3925), .ZN(n4408) );
  XNOR2_X1 U2700 ( .A(n3926), .B(n4487), .ZN(n4419) );
  NOR2_X1 U2701 ( .A1(n4443), .A2(n3956), .ZN(n4452) );
  NAND2_X1 U2702 ( .A1(n4438), .A2(n3930), .ZN(n4446) );
  INV_X1 U2703 ( .A(n4406), .ZN(n4456) );
  XNOR2_X1 U2704 ( .A(n2120), .B(n3960), .ZN(n3965) );
  NAND2_X1 U2705 ( .A1(n4461), .A2(n2088), .ZN(n2120) );
  AOI21_X1 U2706 ( .B1(n2051), .B2(n4197), .A(n4194), .ZN(n4361) );
  OAI21_X1 U2707 ( .B1(n2262), .B2(n2266), .A(n2256), .ZN(n2255) );
  INV_X1 U2708 ( .A(n4212), .ZN(n4027) );
  OAI21_X1 U2709 ( .B1(n4047), .B2(n2251), .A(n2249), .ZN(n4021) );
  NAND2_X1 U2710 ( .A1(n4047), .A2(n2584), .ZN(n2253) );
  NAND2_X1 U2711 ( .A1(n4148), .A2(n4151), .ZN(n4147) );
  NAND2_X1 U2712 ( .A1(n2243), .A2(n2242), .ZN(n4148) );
  NAND2_X1 U2713 ( .A1(n3593), .A2(n3510), .ZN(n4168) );
  NAND2_X1 U2714 ( .A1(n3585), .A2(n2541), .ZN(n4171) );
  INV_X1 U2715 ( .A(n4283), .ZN(n3852) );
  INV_X1 U2716 ( .A(n3869), .ZN(n3274) );
  NAND2_X1 U2717 ( .A1(n2977), .A2(n3525), .ZN(n2996) );
  OAI21_X1 U2718 ( .B1(n3480), .B2(n2108), .A(n2743), .ZN(n2744) );
  OR2_X1 U2719 ( .A1(n4160), .A2(n3098), .ZN(n4139) );
  INV_X1 U2720 ( .A(DATAI_1_), .ZN(n2152) );
  AND2_X1 U2721 ( .A1(n4164), .A2(n4240), .ZN(n4179) );
  INV_X2 U2722 ( .A(n4515), .ZN(n4517) );
  AND3_X1 U2723 ( .A1(n3343), .A2(n3342), .A3(n3341), .ZN(n3346) );
  INV_X2 U2724 ( .A(n4510), .ZN(n4512) );
  INV_X1 U2725 ( .A(n2688), .ZN(n3722) );
  NAND2_X1 U2726 ( .A1(n2776), .A2(n2775), .ZN(n4479) );
  INV_X1 U2727 ( .A(n2706), .ZN(n3721) );
  NAND2_X1 U2728 ( .A1(n2772), .A2(STATE_REG_SCAN_IN), .ZN(n4480) );
  INV_X1 U2729 ( .A(n2889), .ZN(n3581) );
  XNOR2_X1 U2730 ( .A(n2631), .B(IR_REG_19__SCAN_IN), .ZN(n4352) );
  AND2_X1 U2731 ( .A1(n2539), .A2(n2528), .ZN(n4485) );
  OR2_X1 U2732 ( .A1(n2464), .A2(n2463), .ZN(n4493) );
  AND2_X1 U2733 ( .A1(n2395), .A2(n2381), .ZN(n4358) );
  XNOR2_X1 U2734 ( .A(n2098), .B(n3736), .ZN(n3741) );
  AOI21_X1 U2735 ( .B1(n2156), .B2(n2155), .A(n2153), .ZN(n4466) );
  INV_X1 U2736 ( .A(n2154), .ZN(n2153) );
  AND2_X1 U2737 ( .A1(n2716), .A2(n2278), .ZN(n2719) );
  OR2_X1 U2738 ( .A1(n4305), .A2(n4294), .ZN(n2101) );
  NAND2_X1 U2739 ( .A1(n2159), .A2(n2053), .ZN(n2740) );
  AOI21_X1 U2740 ( .B1(n2717), .B2(n4512), .A(n2713), .ZN(n2714) );
  NAND2_X1 U2741 ( .A1(n2712), .A2(n2280), .ZN(n2713) );
  OR2_X1 U2742 ( .A1(n4305), .A2(n4347), .ZN(n2102) );
  NAND2_X1 U2743 ( .A1(n2150), .A2(n2149), .ZN(U3351) );
  NAND2_X1 U2744 ( .A1(U3149), .A2(DATAI_1_), .ZN(n2149) );
  AND2_X1 U2745 ( .A1(n3275), .A2(n3360), .ZN(n2049) );
  OR2_X1 U2746 ( .A1(n4136), .A2(n2129), .ZN(n2050) );
  OR2_X1 U2747 ( .A1(n3988), .A2(n2136), .ZN(n2051) );
  AND2_X1 U2748 ( .A1(n2253), .A2(n2254), .ZN(n4034) );
  AND2_X1 U2749 ( .A1(n4222), .A2(n2709), .ZN(n2583) );
  NOR2_X1 U2750 ( .A1(n2188), .A2(n2190), .ZN(n3244) );
  INV_X1 U2751 ( .A(n3747), .ZN(n3617) );
  NAND2_X1 U2752 ( .A1(n4153), .A2(n4260), .ZN(n2052) );
  INV_X1 U2753 ( .A(n3233), .ZN(n3360) );
  NAND2_X1 U2754 ( .A1(n2319), .A2(n2318), .ZN(n4106) );
  INV_X1 U2755 ( .A(n2213), .ZN(n2212) );
  NAND2_X1 U2756 ( .A1(n3808), .A2(n2070), .ZN(n2213) );
  AND2_X1 U2757 ( .A1(n2443), .A2(n2436), .ZN(n4354) );
  OR2_X1 U2758 ( .A1(n4512), .A2(REG0_REG_29__SCAN_IN), .ZN(n2053) );
  OR2_X1 U2759 ( .A1(n3988), .A2(n2720), .ZN(n2054) );
  AND2_X1 U2760 ( .A1(n2211), .A2(n2209), .ZN(n2055) );
  NAND2_X1 U2761 ( .A1(n2228), .A2(n3635), .ZN(n3788) );
  AND2_X1 U2762 ( .A1(n2207), .A2(n2206), .ZN(n3833) );
  INV_X1 U2763 ( .A(n4349), .ZN(n2119) );
  AND2_X1 U2764 ( .A1(n2115), .A2(n3976), .ZN(n2056) );
  NAND2_X1 U2765 ( .A1(n3649), .A2(n3648), .ZN(n3805) );
  INV_X1 U2766 ( .A(n2112), .ZN(n4017) );
  NOR2_X1 U2767 ( .A1(n4032), .A2(n3461), .ZN(n2112) );
  AND2_X1 U2768 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2057)
         );
  AND2_X1 U2769 ( .A1(n3272), .A2(n3264), .ZN(n2058) );
  INV_X1 U2770 ( .A(n3121), .ZN(n3114) );
  OR2_X1 U2771 ( .A1(n2818), .A2(n2399), .ZN(n2059) );
  NAND2_X1 U2772 ( .A1(n3185), .A2(n3184), .ZN(n2060) );
  AND2_X1 U2773 ( .A1(n2137), .A2(n4358), .ZN(n2061) );
  NAND2_X1 U2774 ( .A1(n2225), .A2(n3637), .ZN(n3824) );
  OR2_X1 U2775 ( .A1(n2796), .A2(n2146), .ZN(n2062) );
  AND2_X1 U2776 ( .A1(n2144), .A2(n2059), .ZN(n2063) );
  AND2_X1 U2777 ( .A1(n2859), .A2(n2860), .ZN(n2064) );
  AND2_X1 U2778 ( .A1(n2325), .A2(n2092), .ZN(n2065) );
  AND2_X1 U2779 ( .A1(n2189), .A2(n3243), .ZN(n2066) );
  NAND2_X1 U2780 ( .A1(n3128), .A2(n3127), .ZN(n2067) );
  AND2_X1 U2781 ( .A1(n2276), .A2(n2307), .ZN(n2068) );
  INV_X1 U2782 ( .A(n3985), .ZN(n2172) );
  OR2_X1 U2783 ( .A1(n4038), .A2(n4212), .ZN(n2069) );
  INV_X1 U2784 ( .A(n4151), .ZN(n2241) );
  INV_X1 U2785 ( .A(n3501), .ZN(n2266) );
  NAND2_X1 U2786 ( .A1(n2177), .A2(n2176), .ZN(n3742) );
  NAND2_X1 U2787 ( .A1(n3246), .A2(n3245), .ZN(n3259) );
  NAND2_X1 U2788 ( .A1(n2179), .A2(n2182), .ZN(n3600) );
  INV_X1 U2789 ( .A(n3690), .ZN(n2198) );
  OR2_X1 U2790 ( .A1(n3771), .A2(n3770), .ZN(n2070) );
  NAND2_X1 U2791 ( .A1(n2178), .A2(n3264), .ZN(n3270) );
  AND2_X1 U2792 ( .A1(n4274), .A2(n4186), .ZN(n2071) );
  AND2_X1 U2793 ( .A1(n3990), .A2(n2720), .ZN(n2072) );
  INV_X1 U2794 ( .A(n2128), .ZN(n4074) );
  NOR3_X1 U2795 ( .A1(n4136), .A2(n2130), .A3(n4239), .ZN(n2128) );
  NOR2_X1 U2796 ( .A1(n4054), .A2(n4042), .ZN(n2073) );
  AND2_X1 U2797 ( .A1(n2174), .A2(n3435), .ZN(n2074) );
  AND2_X1 U2798 ( .A1(n2049), .A2(n3400), .ZN(n2075) );
  AND2_X1 U2799 ( .A1(n2084), .A2(n2180), .ZN(n2076) );
  INV_X1 U2800 ( .A(n2275), .ZN(n3232) );
  NOR2_X1 U2801 ( .A1(n3231), .A2(n3490), .ZN(n2275) );
  OR2_X1 U2802 ( .A1(n3755), .A2(n3756), .ZN(n2077) );
  AND2_X1 U2803 ( .A1(n4269), .A2(n3852), .ZN(n2078) );
  INV_X1 U2804 ( .A(n2210), .ZN(n2209) );
  NAND2_X1 U2805 ( .A1(n2214), .A2(n2215), .ZN(n2210) );
  NOR2_X1 U2806 ( .A1(n4213), .A2(n4221), .ZN(n2079) );
  INV_X1 U2807 ( .A(n4289), .ZN(n3864) );
  AND4_X1 U2808 ( .A1(n2345), .A2(n2344), .A3(n2343), .A4(n2342), .ZN(n4289)
         );
  AND2_X1 U2809 ( .A1(n2251), .A2(n2069), .ZN(n2080) );
  AND2_X1 U2810 ( .A1(n2245), .A2(n4159), .ZN(n2081) );
  INV_X1 U2811 ( .A(n2205), .ZN(n2204) );
  NAND2_X1 U2812 ( .A1(n2206), .A2(n3834), .ZN(n2205) );
  AND2_X1 U2813 ( .A1(n2249), .A2(n2069), .ZN(n2082) );
  INV_X1 U2814 ( .A(n2583), .ZN(n2254) );
  NOR2_X1 U2815 ( .A1(n2771), .A2(n2568), .ZN(n4105) );
  AND2_X1 U2816 ( .A1(n3152), .A2(n3275), .ZN(n2083) );
  INV_X1 U2817 ( .A(n2190), .ZN(n2189) );
  OAI21_X1 U2818 ( .B1(n2194), .B2(n2191), .A(n2060), .ZN(n2190) );
  OR2_X1 U2819 ( .A1(n2994), .A2(n3482), .ZN(n2993) );
  NAND2_X1 U2820 ( .A1(n2742), .A2(n2373), .ZN(n2976) );
  OR2_X1 U2821 ( .A1(n2881), .A2(n2640), .ZN(n4066) );
  NAND2_X1 U2822 ( .A1(n3011), .A2(n2974), .ZN(n3002) );
  INV_X1 U2823 ( .A(n3002), .ZN(n2134) );
  NAND2_X1 U2824 ( .A1(n3406), .A2(n3405), .ZN(n2084) );
  AND2_X1 U2825 ( .A1(n2097), .A2(n2932), .ZN(n2085) );
  AND2_X1 U2826 ( .A1(n2677), .A2(n2276), .ZN(n2086) );
  AND2_X1 U2827 ( .A1(n2143), .A2(n2145), .ZN(n2087) );
  INV_X1 U2828 ( .A(n3957), .ZN(n4483) );
  INV_X1 U2829 ( .A(n4353), .ZN(n2121) );
  OR2_X1 U2830 ( .A1(n4482), .A2(n3959), .ZN(n2088) );
  NAND2_X1 U2831 ( .A1(n2286), .A2(n2089), .ZN(n3848) );
  OAI21_X1 U2832 ( .B1(n3778), .B2(n3847), .A(n2089), .ZN(n3779) );
  NAND2_X1 U2833 ( .A1(n3627), .A2(n3626), .ZN(n2089) );
  NAND2_X1 U2834 ( .A1(n2370), .A2(n2293), .ZN(n2378) );
  AND2_X2 U2835 ( .A1(n2090), .A2(n2067), .ZN(n3171) );
  OR2_X2 U2836 ( .A1(n3118), .A2(n3117), .ZN(n2090) );
  NOR2_X1 U2837 ( .A1(n3112), .A2(n3111), .ZN(n3118) );
  NOR2_X2 U2838 ( .A1(n3038), .A2(n3039), .ZN(n3112) );
  NAND2_X1 U2839 ( .A1(n2091), .A2(n2859), .ZN(n2914) );
  NAND2_X1 U2840 ( .A1(n2064), .A2(n2091), .ZN(n2866) );
  INV_X1 U2841 ( .A(n2093), .ZN(n2684) );
  NOR2_X1 U2842 ( .A1(n2958), .A2(n2085), .ZN(n2937) );
  NAND2_X1 U2843 ( .A1(n3757), .A2(n3672), .ZN(n3675) );
  OAI21_X2 U2844 ( .B1(n3804), .B2(n2210), .A(n2208), .ZN(n3757) );
  NAND2_X2 U2845 ( .A1(n3805), .A2(n3806), .ZN(n3804) );
  NAND2_X1 U2846 ( .A1(n4207), .A2(n2101), .ZN(U3545) );
  NAND2_X1 U2847 ( .A1(n4304), .A2(n2102), .ZN(U3513) );
  INV_X1 U2848 ( .A(n2110), .ZN(n4078) );
  OAI21_X2 U2849 ( .B1(n4087), .B2(n2235), .A(n2234), .ZN(n2110) );
  AOI21_X2 U2850 ( .B1(n4099), .B2(n3465), .A(n3466), .ZN(n4087) );
  NAND2_X2 U2851 ( .A1(n2562), .A2(n2561), .ZN(n4099) );
  NAND2_X1 U2852 ( .A1(n2269), .A2(n2267), .ZN(n2994) );
  AOI21_X2 U2853 ( .B1(n3368), .B2(n2529), .A(n2078), .ZN(n3587) );
  NOR2_X2 U2854 ( .A1(n2679), .A2(IR_REG_25__SCAN_IN), .ZN(n2677) );
  NAND2_X1 U2855 ( .A1(n2677), .A2(n2306), .ZN(n2678) );
  AOI21_X1 U2856 ( .B1(n3973), .B2(n4504), .A(n2160), .ZN(n2115) );
  NAND3_X1 U2857 ( .A1(n2117), .A2(n2116), .A3(n2255), .ZN(n3973) );
  NAND2_X1 U2858 ( .A1(n3984), .A2(n2258), .ZN(n2116) );
  OR2_X1 U2859 ( .A1(n3984), .A2(n2259), .ZN(n2117) );
  INV_X2 U2860 ( .A(n2362), .ZN(n2347) );
  OR2_X2 U2861 ( .A1(n4350), .A2(n2119), .ZN(n2362) );
  AND2_X2 U2862 ( .A1(n2313), .A2(n2309), .ZN(n4350) );
  XNOR2_X2 U2863 ( .A(n2353), .B(IR_REG_1__SCAN_IN), .ZN(n2148) );
  INV_X1 U2864 ( .A(n2126), .ZN(n3312) );
  INV_X1 U2865 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2146) );
  NAND2_X1 U2866 ( .A1(n2148), .A2(REG2_REG_1__SCAN_IN), .ZN(n3894) );
  NAND2_X1 U2867 ( .A1(n2148), .A2(REG1_REG_1__SCAN_IN), .ZN(n2802) );
  NAND2_X1 U2868 ( .A1(n2148), .A2(STATE_REG_SCAN_IN), .ZN(n2150) );
  XNOR2_X1 U2869 ( .A(n2148), .B(n2348), .ZN(n3881) );
  NAND2_X1 U2870 ( .A1(n2354), .A2(n2148), .ZN(n2151) );
  NAND2_X1 U2871 ( .A1(n3906), .A2(n2148), .ZN(n3887) );
  NOR2_X1 U2872 ( .A1(n3927), .A2(n4418), .ZN(n4428) );
  NAND2_X1 U2873 ( .A1(n4448), .A2(n4446), .ZN(n4447) );
  NAND2_X1 U2874 ( .A1(n3920), .A2(n4367), .ZN(n3921) );
  NAND2_X1 U2875 ( .A1(n3923), .A2(n4387), .ZN(n3924) );
  INV_X2 U2876 ( .A(n2354), .ZN(n3428) );
  AOI21_X1 U2877 ( .B1(n4017), .B2(n2168), .A(n2166), .ZN(n2724) );
  OAI21_X2 U2878 ( .B1(n3742), .B2(n3744), .A(n3743), .ZN(n3627) );
  NAND2_X1 U2879 ( .A1(n2187), .A2(n2066), .ZN(n3246) );
  OR2_X2 U2880 ( .A1(n3171), .A2(n2192), .ZN(n2187) );
  INV_X1 U2881 ( .A(n2187), .ZN(n2188) );
  NAND2_X1 U2882 ( .A1(n3691), .A2(n3690), .ZN(n2207) );
  INV_X1 U2883 ( .A(n3689), .ZN(n2206) );
  NAND2_X1 U2884 ( .A1(n2216), .A2(n2219), .ZN(n3764) );
  NAND3_X1 U2885 ( .A1(n2286), .A2(n3630), .A3(n2217), .ZN(n2216) );
  NAND3_X1 U2886 ( .A1(n3630), .A2(n2286), .A3(n3780), .ZN(n2228) );
  NAND2_X2 U2887 ( .A1(n3325), .A2(n3324), .ZN(n3323) );
  AOI21_X2 U2888 ( .B1(n2514), .B2(n2285), .A(n2279), .ZN(n3325) );
  NAND2_X1 U2889 ( .A1(n2300), .A2(n2232), .ZN(n2233) );
  NOR2_X2 U2890 ( .A1(n2233), .A2(n2404), .ZN(n2551) );
  NAND2_X1 U2891 ( .A1(n2236), .A2(n2239), .ZN(n4123) );
  NAND2_X1 U2892 ( .A1(n4047), .A2(n2082), .ZN(n2246) );
  NAND2_X1 U2893 ( .A1(n2246), .A2(n2247), .ZN(n3999) );
  OAI21_X1 U2894 ( .B1(n3984), .B2(n2616), .A(n2261), .ZN(n2722) );
  AND2_X1 U2895 ( .A1(n2383), .A2(n2268), .ZN(n2267) );
  NAND2_X1 U2896 ( .A1(n2382), .A2(n2270), .ZN(n2268) );
  NAND3_X1 U2897 ( .A1(n2372), .A2(n2651), .A3(n2382), .ZN(n2269) );
  OAI21_X1 U2898 ( .B1(n3231), .B2(n2273), .A(n2271), .ZN(n3301) );
  OR2_X1 U2899 ( .A1(n2914), .A2(n3401), .ZN(n2915) );
  NAND2_X2 U2900 ( .A1(n2856), .A2(n2858), .ZN(n3708) );
  NAND2_X1 U2901 ( .A1(n3029), .A2(n2861), .ZN(n2906) );
  INV_X1 U2902 ( .A(n2904), .ZN(n2912) );
  AOI21_X2 U2903 ( .B1(n2960), .B2(n2959), .A(n2958), .ZN(n3037) );
  OAI21_X2 U2904 ( .B1(n3151), .B2(n2479), .A(n2478), .ZN(n3231) );
  OAI21_X2 U2905 ( .B1(n3147), .B2(n2466), .A(n2465), .ZN(n3151) );
  AND2_X2 U2906 ( .A1(n4349), .A2(n4350), .ZN(n2355) );
  OR2_X1 U2907 ( .A1(n4517), .A2(n2621), .ZN(n2278) );
  AND2_X1 U2908 ( .A1(n3865), .A2(n3296), .ZN(n2279) );
  OR2_X1 U2909 ( .A1(n4512), .A2(n2711), .ZN(n2280) );
  AND4_X1 U2910 ( .A1(n2538), .A2(n2537), .A3(n2536), .A4(n2535), .ZN(n4264)
         );
  INV_X1 U2911 ( .A(n4264), .ZN(n4285) );
  NAND2_X1 U2912 ( .A1(n2355), .A2(REG3_REG_0__SCAN_IN), .ZN(n2281) );
  AND2_X1 U2913 ( .A1(n2294), .A2(n2379), .ZN(n2282) );
  OR2_X1 U2914 ( .A1(n3866), .A2(n3411), .ZN(n2284) );
  INV_X1 U2915 ( .A(n4294), .ZN(n2734) );
  NAND2_X1 U2916 ( .A1(n3602), .A2(n3606), .ZN(n2285) );
  XNOR2_X1 U2917 ( .A(n2926), .B(n3401), .ZN(n2957) );
  NAND2_X1 U2918 ( .A1(n4512), .A2(n4276), .ZN(n4347) );
  INV_X1 U2919 ( .A(n4347), .ZN(n2738) );
  INV_X1 U2920 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2503) );
  OAI22_X1 U2921 ( .A1(n3176), .A2(n2964), .B1(n3702), .B2(n3134), .ZN(n3168)
         );
  INV_X1 U2922 ( .A(n4137), .ZN(n4132) );
  OR2_X1 U2923 ( .A1(n3627), .A2(n3626), .ZN(n2286) );
  OR2_X1 U2924 ( .A1(n4244), .A2(n4072), .ZN(n2287) );
  AND2_X1 U2925 ( .A1(n3672), .A2(n3673), .ZN(n2288) );
  OR2_X1 U2926 ( .A1(n4155), .A2(n4137), .ZN(n2289) );
  INV_X1 U2927 ( .A(n4155), .ZN(n3862) );
  AND2_X1 U2928 ( .A1(n2558), .A2(n2557), .ZN(n4155) );
  NAND2_X2 U2929 ( .A1(n2752), .A2(n4468), .ZN(n4164) );
  INV_X1 U2930 ( .A(IR_REG_4__SCAN_IN), .ZN(n2294) );
  INV_X1 U2931 ( .A(n3615), .ZN(n3611) );
  INV_X1 U2932 ( .A(n3261), .ZN(n3262) );
  INV_X1 U2933 ( .A(IR_REG_26__SCAN_IN), .ZN(n2306) );
  NAND2_X1 U2934 ( .A1(n3263), .A2(n3262), .ZN(n3264) );
  OR2_X1 U2935 ( .A1(n4090), .A2(n4072), .ZN(n4051) );
  NAND2_X1 U2936 ( .A1(n3120), .A2(n2997), .ZN(n3526) );
  INV_X1 U2937 ( .A(n3169), .ZN(n3172) );
  INV_X1 U2938 ( .A(n2964), .ZN(n3704) );
  AND2_X1 U2939 ( .A1(n3110), .A2(n3109), .ZN(n3111) );
  OR2_X1 U2940 ( .A1(n2607), .A2(n4554), .ZN(n2617) );
  NAND2_X1 U2941 ( .A1(n2327), .A2(n2291), .ZN(n2564) );
  NOR2_X1 U2942 ( .A1(n2771), .A2(n2625), .ZN(n2720) );
  OR2_X1 U2943 ( .A1(n4222), .A2(n4058), .ZN(n3463) );
  NAND2_X1 U2944 ( .A1(n4270), .A2(n4285), .ZN(n2541) );
  OR2_X1 U2945 ( .A1(n3359), .A2(n3275), .ZN(n2478) );
  NAND2_X1 U2946 ( .A1(n3581), .A2(n4351), .ZN(n2882) );
  NOR2_X1 U2947 ( .A1(n2771), .A2(n4604), .ZN(n4212) );
  INV_X1 U2948 ( .A(n4493), .ZN(n3935) );
  INV_X1 U2949 ( .A(IR_REG_9__SCAN_IN), .ZN(n2334) );
  OR2_X1 U2950 ( .A1(n2585), .A2(n4635), .ZN(n2597) );
  AND2_X1 U2951 ( .A1(n2437), .A2(REG3_REG_8__SCAN_IN), .ZN(n2452) );
  OR2_X1 U2952 ( .A1(n2493), .A2(n4665), .ZN(n2504) );
  AND2_X1 U2953 ( .A1(n2290), .A2(REG3_REG_10__SCAN_IN), .ZN(n2468) );
  INV_X1 U2954 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2814) );
  NOR2_X1 U2955 ( .A1(n2506), .A2(n3748), .ZN(n2339) );
  OR2_X1 U2956 ( .A1(n3837), .A2(n2609), .ZN(n2605) );
  INV_X1 U2957 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3748) );
  INV_X1 U2958 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4626) );
  INV_X1 U2959 ( .A(n3861), .ZN(n4005) );
  NAND2_X1 U2960 ( .A1(n3428), .A2(DATAI_24_), .ZN(n4042) );
  NAND2_X1 U2961 ( .A1(n2897), .A2(n2773), .ZN(n4273) );
  INV_X1 U2962 ( .A(n4270), .ZN(n3628) );
  OR2_X1 U2963 ( .A1(n2776), .A2(D_REG_0__SCAN_IN), .ZN(n2708) );
  NOR2_X1 U2964 ( .A1(n2771), .A2(n2615), .ZN(n4199) );
  NAND2_X1 U2965 ( .A1(n3428), .A2(DATAI_22_), .ZN(n4072) );
  INV_X1 U2966 ( .A(n3400), .ZN(n3411) );
  INV_X1 U2967 ( .A(n4240), .ZN(n4288) );
  AND2_X1 U2968 ( .A1(n2678), .A2(n2324), .ZN(n2725) );
  AND2_X1 U2969 ( .A1(n2426), .A2(REG3_REG_7__SCAN_IN), .ZN(n2437) );
  AND2_X1 U2970 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2398) );
  NAND2_X1 U2971 ( .A1(n2452), .A2(REG3_REG_9__SCAN_IN), .ZN(n2470) );
  OR2_X1 U2972 ( .A1(n2504), .A2(n2503), .ZN(n2506) );
  NAND2_X1 U2973 ( .A1(n2468), .A2(REG3_REG_11__SCAN_IN), .ZN(n2493) );
  NOR2_X1 U2974 ( .A1(n2414), .A2(n2814), .ZN(n2426) );
  NAND3_X1 U2975 ( .A1(n2968), .A2(n2967), .A3(n3583), .ZN(n3843) );
  OR2_X1 U2976 ( .A1(n3737), .A2(n2609), .ZN(n2614) );
  INV_X1 U2977 ( .A(n2925), .ZN(n2941) );
  AND2_X1 U2978 ( .A1(n2782), .A2(n2781), .ZN(n2797) );
  INV_X1 U2979 ( .A(n4066), .ZN(n4282) );
  INV_X1 U2980 ( .A(n4167), .ZN(n4173) );
  INV_X1 U2981 ( .A(n4139), .ZN(n4473) );
  AND2_X1 U2982 ( .A1(n4164), .A2(n4284), .ZN(n4178) );
  OR2_X1 U2983 ( .A1(n2895), .A2(n2751), .ZN(n4468) );
  NAND2_X1 U2984 ( .A1(n2708), .A2(n2707), .ZN(n2749) );
  INV_X1 U2985 ( .A(n4504), .ZN(n4280) );
  NAND2_X1 U2986 ( .A1(n4111), .A2(n3281), .ZN(n4504) );
  AND2_X1 U2987 ( .A1(n2851), .A2(n2889), .ZN(n4502) );
  AND2_X1 U2988 ( .A1(n2491), .A2(n2499), .ZN(n3934) );
  AND2_X1 U2989 ( .A1(n2782), .A2(n2774), .ZN(n4460) );
  OR2_X1 U2990 ( .A1(n2921), .A2(n2896), .ZN(n3845) );
  INV_X1 U2991 ( .A(n4202), .ZN(n3990) );
  NAND2_X1 U2992 ( .A1(n2573), .A2(n2572), .ZN(n4090) );
  INV_X1 U2993 ( .A(n4269), .ZN(n3863) );
  INV_X1 U2995 ( .A(n4488), .ZN(n4417) );
  NAND2_X1 U2996 ( .A1(n2797), .A2(n2897), .ZN(n4467) );
  INV_X1 U2997 ( .A(n4164), .ZN(n4360) );
  INV_X1 U2998 ( .A(n4164), .ZN(n4118) );
  NAND2_X1 U2999 ( .A1(n4164), .A2(n3008), .ZN(n4167) );
  NAND2_X1 U3000 ( .A1(n4517), .A2(n4276), .ZN(n4294) );
  OR2_X1 U3001 ( .A1(n2715), .A2(n2749), .ZN(n4515) );
  NAND2_X1 U3002 ( .A1(n2735), .A2(n2738), .ZN(n2739) );
  AND3_X1 U3003 ( .A1(n4509), .A2(n4508), .A3(n4507), .ZN(n4516) );
  OR2_X1 U3004 ( .A1(n2715), .A2(n2886), .ZN(n4510) );
  INV_X1 U3005 ( .A(n4480), .ZN(n2778) );
  INV_X1 U3006 ( .A(n3946), .ZN(n4490) );
  AND2_X1 U3007 ( .A1(n2424), .A2(n2433), .ZN(n4355) );
  INV_X1 U3008 ( .A(n2714), .ZN(U3514) );
  NAND2_X1 U3009 ( .A1(n2398), .A2(REG3_REG_5__SCAN_IN), .ZN(n2414) );
  AND2_X1 U3010 ( .A1(REG3_REG_19__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .ZN(
        n2291) );
  NAND2_X1 U3011 ( .A1(n2564), .A2(n4630), .ZN(n2292) );
  AND2_X1 U3012 ( .A1(n2576), .A2(n2292), .ZN(n4091) );
  INV_X1 U3013 ( .A(n2378), .ZN(n2295) );
  NAND2_X1 U3014 ( .A1(n2295), .A2(n2282), .ZN(n2404) );
  NOR2_X2 U3015 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2335)
         );
  NAND2_X1 U3016 ( .A1(n2551), .A2(n2305), .ZN(n2679) );
  NAND2_X1 U3017 ( .A1(n2046), .A2(n2310), .ZN(n2311) );
  NAND2_X1 U3018 ( .A1(n2311), .A2(IR_REG_31__SCAN_IN), .ZN(n2312) );
  NAND2_X1 U3019 ( .A1(n4091), .A2(n2355), .ZN(n2319) );
  INV_X1 U3020 ( .A(n2365), .ZN(n2338) );
  INV_X2 U3021 ( .A(n2338), .ZN(n3419) );
  INV_X1 U3022 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4247) );
  INV_X2 U3023 ( .A(n2364), .ZN(n2645) );
  NAND2_X1 U3024 ( .A1(n2645), .A2(REG0_REG_21__SCAN_IN), .ZN(n2316) );
  NAND2_X1 U3026 ( .A1(n2384), .A2(REG2_REG_21__SCAN_IN), .ZN(n2315) );
  OAI211_X1 U3027 ( .C1(n3419), .C2(n4247), .A(n2316), .B(n2315), .ZN(n2317)
         );
  INV_X1 U3028 ( .A(n2317), .ZN(n2318) );
  INV_X1 U3029 ( .A(n4106), .ZN(n4067) );
  NAND2_X1 U3030 ( .A1(n2321), .A2(n2642), .ZN(n2322) );
  NAND2_X1 U3031 ( .A1(n3428), .A2(DATAI_21_), .ZN(n4094) );
  INV_X1 U3032 ( .A(n4094), .ZN(n4239) );
  INV_X1 U3033 ( .A(DATAI_18_), .ZN(n4632) );
  NAND2_X1 U3034 ( .A1(n2559), .A2(IR_REG_31__SCAN_IN), .ZN(n2326) );
  XNOR2_X1 U3035 ( .A(n2326), .B(IR_REG_18__SCAN_IN), .ZN(n3933) );
  MUX2_X1 U3036 ( .A(n4632), .B(n4482), .S(n2771), .Z(n4159) );
  INV_X1 U3037 ( .A(n4159), .ZN(n4152) );
  INV_X1 U3038 ( .A(n2327), .ZN(n2563) );
  INV_X1 U3039 ( .A(n2328), .ZN(n2546) );
  INV_X1 U3040 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2329) );
  NAND2_X1 U3041 ( .A1(n2546), .A2(n2329), .ZN(n2330) );
  NAND2_X1 U3042 ( .A1(n2563), .A2(n2330), .ZN(n4161) );
  AOI22_X1 U3043 ( .A1(n2338), .A2(REG1_REG_18__SCAN_IN), .B1(n2645), .B2(
        REG0_REG_18__SCAN_IN), .ZN(n2332) );
  NAND2_X1 U3044 ( .A1(n2347), .A2(REG2_REG_18__SCAN_IN), .ZN(n2331) );
  NAND2_X1 U3045 ( .A1(n2333), .A2(n2334), .ZN(n2487) );
  INV_X1 U3046 ( .A(n2335), .ZN(n2336) );
  OR2_X1 U3047 ( .A1(n2524), .A2(n2642), .ZN(n2337) );
  XNOR2_X1 U3048 ( .A(n2337), .B(IR_REG_14__SCAN_IN), .ZN(n3950) );
  MUX2_X1 U3049 ( .A(DATAI_14_), .B(n3950), .S(n2771), .Z(n3747) );
  NAND2_X1 U3050 ( .A1(n2645), .A2(REG0_REG_14__SCAN_IN), .ZN(n2345) );
  INV_X1 U3051 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3394) );
  OR2_X1 U3052 ( .A1(n2365), .A2(n3394), .ZN(n2344) );
  INV_X1 U3053 ( .A(n2339), .ZN(n2517) );
  NAND2_X1 U3054 ( .A1(n2506), .A2(n3748), .ZN(n2340) );
  NAND2_X1 U3055 ( .A1(n2517), .A2(n2340), .ZN(n3328) );
  OR2_X1 U3056 ( .A1(n2609), .A2(n3328), .ZN(n2343) );
  INV_X1 U3057 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2341) );
  OR2_X1 U3058 ( .A1(n2314), .A2(n2341), .ZN(n2342) );
  INV_X1 U3059 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2346) );
  NAND2_X1 U3060 ( .A1(n2347), .A2(REG2_REG_1__SCAN_IN), .ZN(n2350) );
  INV_X1 U3061 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U3062 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2353)
         );
  INV_X1 U3063 ( .A(n3029), .ZN(n2905) );
  NAND2_X1 U3064 ( .A1(n3877), .A2(n2905), .ZN(n3515) );
  NAND2_X1 U3065 ( .A1(n2912), .A2(n3029), .ZN(n3519) );
  INV_X1 U3066 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2356) );
  INV_X1 U3067 ( .A(n2362), .ZN(n2384) );
  NAND2_X1 U3068 ( .A1(n2384), .A2(REG2_REG_0__SCAN_IN), .ZN(n2359) );
  INV_X1 U3069 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2357) );
  NAND4_X1 U3070 ( .A1(n2281), .A2(n2360), .A3(n2359), .A4(n2358), .ZN(n2857)
         );
  MUX2_X1 U3071 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(n2354), .Z(n2948) );
  AND2_X1 U3072 ( .A1(n2857), .A2(n2948), .ZN(n2938) );
  NAND2_X1 U3073 ( .A1(n2650), .A2(n2938), .ZN(n2940) );
  NAND2_X1 U3074 ( .A1(n3877), .A2(n3029), .ZN(n2361) );
  OR2_X1 U3075 ( .A1(n2362), .A2(n3893), .ZN(n2368) );
  INV_X1 U3076 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2363) );
  INV_X1 U3077 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2801) );
  NAND3_X1 U3078 ( .A1(n2368), .A2(n2367), .A3(n2366), .ZN(n2369) );
  OR2_X1 U3079 ( .A1(n2370), .A2(n2642), .ZN(n2371) );
  MUX2_X1 U3080 ( .A(DATAI_2_), .B(n2048), .S(n2354), .Z(n2984) );
  INV_X1 U3081 ( .A(n2984), .ZN(n2927) );
  NAND2_X1 U3082 ( .A1(n2941), .A2(n2927), .ZN(n3523) );
  NAND2_X1 U3083 ( .A1(n2925), .A2(n2984), .ZN(n3520) );
  NAND2_X1 U3084 ( .A1(n2925), .A2(n2927), .ZN(n2373) );
  NAND2_X1 U3085 ( .A1(n2645), .A2(REG0_REG_3__SCAN_IN), .ZN(n2377) );
  INV_X1 U3086 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3018) );
  OR2_X1 U3087 ( .A1(n3419), .A2(n3018), .ZN(n2375) );
  INV_X1 U3088 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3909) );
  NAND2_X1 U3089 ( .A1(n2378), .A2(IR_REG_31__SCAN_IN), .ZN(n2380) );
  NAND2_X1 U3090 ( .A1(n2380), .A2(n2379), .ZN(n2395) );
  OR2_X1 U3091 ( .A1(n2380), .A2(n2379), .ZN(n2381) );
  MUX2_X1 U3092 ( .A(DATAI_3_), .B(n4358), .S(n2771), .Z(n2980) );
  NAND2_X1 U3093 ( .A1(n3876), .A2(n2980), .ZN(n2382) );
  NAND2_X1 U3094 ( .A1(n3041), .A2(n3011), .ZN(n2383) );
  NAND2_X1 U3095 ( .A1(n2384), .A2(REG2_REG_4__SCAN_IN), .ZN(n2389) );
  INV_X1 U3096 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2385) );
  OR2_X1 U3097 ( .A1(n2365), .A2(n2385), .ZN(n2388) );
  INV_X1 U3098 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2386) );
  OR2_X1 U3099 ( .A1(n2364), .A2(n2386), .ZN(n2387) );
  INV_X1 U3100 ( .A(n2398), .ZN(n2392) );
  INV_X1 U3101 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2969) );
  INV_X1 U3102 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3103 ( .A1(n2969), .A2(n2390), .ZN(n2391) );
  NAND2_X1 U3104 ( .A1(n2392), .A2(n2391), .ZN(n3047) );
  OR2_X1 U3105 ( .A1(n2609), .A2(n3047), .ZN(n2393) );
  NAND2_X1 U3106 ( .A1(n2395), .A2(IR_REG_31__SCAN_IN), .ZN(n2396) );
  XNOR2_X1 U3107 ( .A(n2396), .B(IR_REG_4__SCAN_IN), .ZN(n4357) );
  MUX2_X1 U3108 ( .A(DATAI_4_), .B(n4357), .S(n2354), .Z(n2997) );
  INV_X1 U3109 ( .A(n2997), .ZN(n3042) );
  NAND2_X1 U3110 ( .A1(n3875), .A2(n3042), .ZN(n3530) );
  NAND2_X1 U3111 ( .A1(n3875), .A2(n2997), .ZN(n2397) );
  NAND2_X1 U3112 ( .A1(n2645), .A2(REG0_REG_5__SCAN_IN), .ZN(n2403) );
  INV_X1 U3113 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2817) );
  OR2_X1 U3114 ( .A1(n3419), .A2(n2817), .ZN(n2402) );
  OAI21_X1 U3115 ( .B1(n2398), .B2(REG3_REG_5__SCAN_IN), .A(n2414), .ZN(n3126)
         );
  OR2_X1 U3116 ( .A1(n2609), .A2(n3126), .ZN(n2401) );
  INV_X1 U3117 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2399) );
  OR2_X1 U3118 ( .A1(n2314), .A2(n2399), .ZN(n2400) );
  INV_X1 U3119 ( .A(DATAI_5_), .ZN(n2410) );
  NAND2_X1 U3120 ( .A1(n2405), .A2(IR_REG_31__SCAN_IN), .ZN(n2406) );
  MUX2_X1 U3121 ( .A(n2406), .B(IR_REG_31__SCAN_IN), .S(n2407), .Z(n2409) );
  INV_X1 U3122 ( .A(n2405), .ZN(n2408) );
  NAND2_X1 U3123 ( .A1(n2408), .A2(n2407), .ZN(n2422) );
  NAND2_X1 U3124 ( .A1(n2409), .A2(n2422), .ZN(n2818) );
  MUX2_X1 U3125 ( .A(n2410), .B(n2818), .S(n2771), .Z(n3121) );
  NAND2_X1 U3126 ( .A1(n3133), .A2(n3121), .ZN(n2411) );
  NAND2_X1 U3127 ( .A1(n3049), .A2(n2411), .ZN(n2413) );
  NAND2_X1 U3128 ( .A1(n3874), .A2(n3114), .ZN(n2412) );
  NAND2_X1 U3129 ( .A1(n2645), .A2(REG0_REG_6__SCAN_IN), .ZN(n2420) );
  INV_X1 U3130 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3085) );
  OR2_X1 U3131 ( .A1(n2314), .A2(n3085), .ZN(n2419) );
  AND2_X1 U3132 ( .A1(n2414), .A2(n2814), .ZN(n2415) );
  OR2_X1 U3133 ( .A1(n2415), .A2(n2426), .ZN(n3139) );
  OR2_X1 U3134 ( .A1(n2609), .A2(n3139), .ZN(n2418) );
  INV_X1 U3135 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2416) );
  OR2_X1 U3136 ( .A1(n3419), .A2(n2416), .ZN(n2417) );
  NAND4_X1 U3137 ( .A1(n2420), .A2(n2419), .A3(n2418), .A4(n2417), .ZN(n3873)
         );
  NAND2_X1 U3138 ( .A1(n2422), .A2(IR_REG_31__SCAN_IN), .ZN(n2421) );
  MUX2_X1 U3139 ( .A(n2421), .B(IR_REG_31__SCAN_IN), .S(n4519), .Z(n2424) );
  INV_X1 U3140 ( .A(n2422), .ZN(n2423) );
  NAND2_X1 U3141 ( .A1(n2423), .A2(n4519), .ZN(n2433) );
  MUX2_X1 U3142 ( .A(DATAI_6_), .B(n4355), .S(n2771), .Z(n3084) );
  AND2_X1 U3143 ( .A1(n3873), .A2(n3084), .ZN(n2425) );
  NAND2_X1 U3144 ( .A1(n2645), .A2(REG0_REG_7__SCAN_IN), .ZN(n2432) );
  OR2_X1 U3145 ( .A1(n2314), .A2(n3102), .ZN(n2431) );
  NOR2_X1 U3146 ( .A1(n2426), .A2(REG3_REG_7__SCAN_IN), .ZN(n2427) );
  OR2_X1 U3147 ( .A1(n2437), .A2(n2427), .ZN(n3182) );
  OR2_X1 U31480 ( .A1(n2609), .A2(n3182), .ZN(n2430) );
  INV_X1 U31490 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2428) );
  OR2_X1 U3150 ( .A1(n3419), .A2(n2428), .ZN(n2429) );
  NAND2_X1 U3151 ( .A1(n2433), .A2(IR_REG_31__SCAN_IN), .ZN(n2435) );
  NAND2_X1 U3152 ( .A1(n2435), .A2(n2434), .ZN(n2443) );
  OR2_X1 U3153 ( .A1(n2435), .A2(n2434), .ZN(n2436) );
  MUX2_X1 U3154 ( .A(DATAI_7_), .B(n4354), .S(n2771), .Z(n3099) );
  NAND2_X1 U3155 ( .A1(n3206), .A2(n3099), .ZN(n2654) );
  INV_X1 U3156 ( .A(n3099), .ZN(n3177) );
  NAND2_X1 U3157 ( .A1(n3871), .A2(n3177), .ZN(n3536) );
  NAND2_X1 U3158 ( .A1(n2645), .A2(REG0_REG_8__SCAN_IN), .ZN(n2442) );
  INV_X1 U3159 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3939) );
  OR2_X1 U3160 ( .A1(n3419), .A2(n3939), .ZN(n2441) );
  NOR2_X1 U3161 ( .A1(n2437), .A2(REG3_REG_8__SCAN_IN), .ZN(n2438) );
  OR2_X1 U3162 ( .A1(n2452), .A2(n2438), .ZN(n4469) );
  OR2_X1 U3163 ( .A1(n2609), .A2(n4469), .ZN(n2440) );
  INV_X1 U3164 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4470) );
  OR2_X1 U3165 ( .A1(n2314), .A2(n4470), .ZN(n2439) );
  INV_X1 U3166 ( .A(DATAI_8_), .ZN(n2446) );
  NAND2_X1 U3167 ( .A1(n2443), .A2(IR_REG_31__SCAN_IN), .ZN(n2445) );
  XNOR2_X1 U3168 ( .A(n2445), .B(n2444), .ZN(n4353) );
  MUX2_X1 U3169 ( .A(n2446), .B(n4353), .S(n2771), .Z(n3205) );
  AND2_X1 U3170 ( .A1(n3252), .A2(n3205), .ZN(n2449) );
  OR2_X1 U3171 ( .A1(n3533), .A2(n2449), .ZN(n2451) );
  NAND2_X1 U3172 ( .A1(n3871), .A2(n3099), .ZN(n3202) );
  NAND2_X1 U3173 ( .A1(n3870), .A2(n3215), .ZN(n2447) );
  AND2_X1 U3174 ( .A1(n3202), .A2(n2447), .ZN(n2448) );
  OR2_X1 U3175 ( .A1(n2449), .A2(n2448), .ZN(n2450) );
  OAI21_X2 U3176 ( .B1(n3106), .B2(n2451), .A(n2450), .ZN(n3147) );
  NAND2_X1 U3177 ( .A1(n2645), .A2(REG0_REG_9__SCAN_IN), .ZN(n2461) );
  INV_X1 U3178 ( .A(n2452), .ZN(n2454) );
  INV_X1 U3179 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2453) );
  NAND2_X1 U3180 ( .A1(n2454), .A2(n2453), .ZN(n2455) );
  NAND2_X1 U3181 ( .A1(n2470), .A2(n2455), .ZN(n3257) );
  OR2_X1 U3182 ( .A1(n2609), .A2(n3257), .ZN(n2460) );
  INV_X1 U3183 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2456) );
  OR2_X1 U3184 ( .A1(n3419), .A2(n2456), .ZN(n2459) );
  INV_X1 U3185 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2457) );
  OR2_X1 U3186 ( .A1(n2314), .A2(n2457), .ZN(n2458) );
  NAND4_X1 U3187 ( .A1(n2461), .A2(n2460), .A3(n2459), .A4(n2458), .ZN(n3869)
         );
  NOR2_X1 U3188 ( .A1(n2333), .A2(n2642), .ZN(n2462) );
  MUX2_X1 U3189 ( .A(n2642), .B(n2462), .S(IR_REG_9__SCAN_IN), .Z(n2464) );
  INV_X1 U3190 ( .A(n2487), .ZN(n2463) );
  MUX2_X1 U3191 ( .A(DATAI_9_), .B(n3935), .S(n2771), .Z(n3247) );
  AND2_X1 U3192 ( .A1(n3869), .A2(n3247), .ZN(n2466) );
  NAND2_X1 U3193 ( .A1(n3274), .A2(n3253), .ZN(n2465) );
  NAND2_X1 U3194 ( .A1(n2645), .A2(REG0_REG_10__SCAN_IN), .ZN(n2476) );
  INV_X1 U3195 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2467) );
  OR2_X1 U3196 ( .A1(n3419), .A2(n2467), .ZN(n2475) );
  INV_X1 U3197 ( .A(n2468), .ZN(n2481) );
  INV_X1 U3198 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3199 ( .A1(n2470), .A2(n2469), .ZN(n2471) );
  NAND2_X1 U3200 ( .A1(n2481), .A2(n2471), .ZN(n3280) );
  OR2_X1 U3201 ( .A1(n2609), .A2(n3280), .ZN(n2474) );
  INV_X1 U3202 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2472) );
  OR2_X1 U3203 ( .A1(n2314), .A2(n2472), .ZN(n2473) );
  NAND4_X1 U3204 ( .A1(n2476), .A2(n2475), .A3(n2474), .A4(n2473), .ZN(n3868)
         );
  NAND2_X1 U3205 ( .A1(n2487), .A2(IR_REG_31__SCAN_IN), .ZN(n2477) );
  XNOR2_X1 U3206 ( .A(n2477), .B(IR_REG_10__SCAN_IN), .ZN(n3942) );
  MUX2_X1 U3207 ( .A(DATAI_10_), .B(n3942), .S(n2771), .Z(n3266) );
  NOR2_X1 U3208 ( .A1(n3868), .A2(n3266), .ZN(n2479) );
  INV_X1 U3209 ( .A(n3868), .ZN(n3359) );
  NAND2_X1 U32100 ( .A1(n2645), .A2(REG0_REG_11__SCAN_IN), .ZN(n2486) );
  INV_X1 U32110 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3288) );
  OR2_X1 U32120 ( .A1(n3419), .A2(n3288), .ZN(n2485) );
  INV_X1 U32130 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2480) );
  NAND2_X1 U32140 ( .A1(n2481), .A2(n2480), .ZN(n2482) );
  NAND2_X1 U32150 ( .A1(n2493), .A2(n2482), .ZN(n3364) );
  OR2_X1 U32160 ( .A1(n2609), .A2(n3364), .ZN(n2484) );
  INV_X1 U32170 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3237) );
  OR2_X1 U32180 ( .A1(n2314), .A2(n3237), .ZN(n2483) );
  OR2_X1 U32190 ( .A1(n2487), .A2(IR_REG_10__SCAN_IN), .ZN(n2488) );
  NAND2_X1 U32200 ( .A1(n2488), .A2(IR_REG_31__SCAN_IN), .ZN(n2490) );
  INV_X1 U32210 ( .A(IR_REG_11__SCAN_IN), .ZN(n2489) );
  OR2_X1 U32220 ( .A1(n2490), .A2(n2489), .ZN(n2491) );
  NAND2_X1 U32230 ( .A1(n2490), .A2(n2489), .ZN(n2499) );
  MUX2_X1 U32240 ( .A(DATAI_11_), .B(n3934), .S(n2771), .Z(n3233) );
  NAND2_X1 U32250 ( .A1(n3356), .A2(n3233), .ZN(n3291) );
  NAND2_X1 U32260 ( .A1(n3867), .A2(n3360), .ZN(n3293) );
  NAND2_X1 U32270 ( .A1(n3356), .A2(n3360), .ZN(n2492) );
  NAND2_X1 U32280 ( .A1(n2645), .A2(REG0_REG_12__SCAN_IN), .ZN(n2498) );
  INV_X1 U32290 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3314) );
  OR2_X1 U32300 ( .A1(n2314), .A2(n3314), .ZN(n2497) );
  NAND2_X1 U32310 ( .A1(n2493), .A2(n4665), .ZN(n2494) );
  NAND2_X1 U32320 ( .A1(n2504), .A2(n2494), .ZN(n3410) );
  OR2_X1 U32330 ( .A1(n2609), .A2(n3410), .ZN(n2496) );
  INV_X1 U32340 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3344) );
  OR2_X1 U32350 ( .A1(n3419), .A2(n3344), .ZN(n2495) );
  INV_X1 U32360 ( .A(DATAI_12_), .ZN(n2501) );
  NAND2_X1 U32370 ( .A1(n2499), .A2(IR_REG_31__SCAN_IN), .ZN(n2500) );
  XNOR2_X1 U32380 ( .A(n2500), .B(IR_REG_12__SCAN_IN), .ZN(n3946) );
  MUX2_X1 U32390 ( .A(n2501), .B(n4490), .S(n2771), .Z(n3400) );
  INV_X1 U32400 ( .A(n3301), .ZN(n2514) );
  NAND2_X1 U32410 ( .A1(n2645), .A2(REG0_REG_13__SCAN_IN), .ZN(n2510) );
  INV_X1 U32420 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4405) );
  OR2_X1 U32430 ( .A1(n2314), .A2(n4405), .ZN(n2509) );
  NAND2_X1 U32440 ( .A1(n2504), .A2(n2503), .ZN(n2505) );
  NAND2_X1 U32450 ( .A1(n2506), .A2(n2505), .ZN(n3610) );
  OR2_X1 U32460 ( .A1(n2609), .A2(n3610), .ZN(n2508) );
  INV_X1 U32470 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3380) );
  OR2_X1 U32480 ( .A1(n2365), .A2(n3380), .ZN(n2507) );
  INV_X1 U32490 ( .A(DATAI_13_), .ZN(n2513) );
  NAND2_X1 U32500 ( .A1(n2511), .A2(IR_REG_31__SCAN_IN), .ZN(n2512) );
  XNOR2_X1 U32510 ( .A(n2512), .B(IR_REG_13__SCAN_IN), .ZN(n4488) );
  MUX2_X1 U32520 ( .A(n2513), .B(n4417), .S(n2771), .Z(n3606) );
  INV_X1 U32530 ( .A(n3606), .ZN(n3296) );
  NAND2_X1 U32540 ( .A1(n4289), .A2(n3747), .ZN(n3432) );
  NAND2_X1 U32550 ( .A1(n3864), .A2(n3617), .ZN(n3509) );
  NAND2_X1 U32560 ( .A1(n3432), .A2(n3509), .ZN(n3324) );
  NAND2_X1 U32570 ( .A1(n2645), .A2(REG0_REG_15__SCAN_IN), .ZN(n2522) );
  INV_X1 U32580 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2515) );
  OR2_X1 U32590 ( .A1(n2314), .A2(n2515), .ZN(n2521) );
  INV_X1 U32600 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2516) );
  NAND2_X1 U32610 ( .A1(n2517), .A2(n2516), .ZN(n2518) );
  NAND2_X1 U32620 ( .A1(n2532), .A2(n2518), .ZN(n3857) );
  OR2_X1 U32630 ( .A1(n2609), .A2(n3857), .ZN(n2520) );
  INV_X1 U32640 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4292) );
  OR2_X1 U32650 ( .A1(n2365), .A2(n4292), .ZN(n2519) );
  INV_X1 U32660 ( .A(IR_REG_14__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U32670 ( .A1(n2524), .A2(n2523), .ZN(n2525) );
  NAND2_X1 U32680 ( .A1(n2525), .A2(IR_REG_31__SCAN_IN), .ZN(n2527) );
  INV_X1 U32690 ( .A(IR_REG_15__SCAN_IN), .ZN(n2526) );
  NAND2_X1 U32700 ( .A1(n2527), .A2(n2526), .ZN(n2539) );
  OR2_X1 U32710 ( .A1(n2527), .A2(n2526), .ZN(n2528) );
  MUX2_X1 U32720 ( .A(DATAI_15_), .B(n4485), .S(n2771), .Z(n4283) );
  NAND2_X1 U32730 ( .A1(n3863), .A2(n4283), .ZN(n2529) );
  NAND2_X1 U32740 ( .A1(n2645), .A2(REG0_REG_16__SCAN_IN), .ZN(n2538) );
  INV_X1 U32750 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2530) );
  OR2_X1 U32760 ( .A1(n2314), .A2(n2530), .ZN(n2537) );
  NAND2_X1 U32770 ( .A1(n2532), .A2(n2531), .ZN(n2533) );
  NAND2_X1 U32780 ( .A1(n2544), .A2(n2533), .ZN(n3590) );
  OR2_X1 U32790 ( .A1(n3590), .A2(n2609), .ZN(n2536) );
  INV_X1 U32800 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2534) );
  OR2_X1 U32810 ( .A1(n3419), .A2(n2534), .ZN(n2535) );
  NAND2_X1 U32820 ( .A1(n2539), .A2(IR_REG_31__SCAN_IN), .ZN(n2540) );
  XNOR2_X1 U32830 ( .A(n2540), .B(IR_REG_16__SCAN_IN), .ZN(n3954) );
  MUX2_X1 U32840 ( .A(DATAI_16_), .B(n3954), .S(n2771), .Z(n4270) );
  NAND2_X1 U32850 ( .A1(n4264), .A2(n4270), .ZN(n3441) );
  NAND2_X1 U32860 ( .A1(n4285), .A2(n3628), .ZN(n3510) );
  NAND2_X1 U32870 ( .A1(n3441), .A2(n3510), .ZN(n3586) );
  INV_X1 U32880 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4340) );
  OR2_X1 U32890 ( .A1(n2364), .A2(n4340), .ZN(n2543) );
  INV_X1 U32900 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4267) );
  OR2_X1 U32910 ( .A1(n3419), .A2(n4267), .ZN(n2542) );
  AND2_X1 U32920 ( .A1(n2543), .A2(n2542), .ZN(n2550) );
  NAND2_X1 U32930 ( .A1(n2544), .A2(n4626), .ZN(n2545) );
  NAND2_X1 U32940 ( .A1(n2546), .A2(n2545), .ZN(n4180) );
  OR2_X1 U32950 ( .A1(n4180), .A2(n2609), .ZN(n2549) );
  INV_X1 U32960 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2547) );
  OR2_X1 U32970 ( .A1(n2314), .A2(n2547), .ZN(n2548) );
  INV_X1 U32980 ( .A(DATAI_17_), .ZN(n2553) );
  OR2_X1 U32990 ( .A1(n2551), .A2(n2642), .ZN(n2552) );
  XNOR2_X1 U33000 ( .A(n2552), .B(IR_REG_17__SCAN_IN), .ZN(n3957) );
  MUX2_X1 U33010 ( .A(n2553), .B(n4483), .S(n2771), .Z(n4186) );
  OR2_X1 U33020 ( .A1(n4261), .A2(n4159), .ZN(n4126) );
  NAND2_X1 U33030 ( .A1(n4261), .A2(n4159), .ZN(n4127) );
  NAND2_X1 U33040 ( .A1(n4126), .A2(n4127), .ZN(n4151) );
  XNOR2_X1 U33050 ( .A(n2563), .B(REG3_REG_19__SCAN_IN), .ZN(n4140) );
  NAND2_X1 U33060 ( .A1(n4140), .A2(n2355), .ZN(n2558) );
  INV_X1 U33070 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4255) );
  NAND2_X1 U33080 ( .A1(n2645), .A2(REG0_REG_19__SCAN_IN), .ZN(n2555) );
  INV_X1 U33090 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4142) );
  OR2_X1 U33100 ( .A1(n2314), .A2(n4142), .ZN(n2554) );
  OAI211_X1 U33110 ( .C1(n4255), .C2(n3419), .A(n2555), .B(n2554), .ZN(n2556)
         );
  INV_X1 U33120 ( .A(n2556), .ZN(n2557) );
  INV_X1 U33130 ( .A(DATAI_19_), .ZN(n4544) );
  INV_X1 U33140 ( .A(n2627), .ZN(n2560) );
  MUX2_X1 U33150 ( .A(n4544), .B(n3963), .S(n2771), .Z(n4137) );
  NAND2_X1 U33160 ( .A1(n4123), .A2(n2289), .ZN(n2562) );
  INV_X1 U33170 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4251) );
  INV_X1 U33180 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4616) );
  INV_X1 U33190 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3811) );
  OAI21_X1 U33200 ( .B1(n2563), .B2(n4616), .A(n3811), .ZN(n2565) );
  NAND2_X1 U33210 ( .A1(n2565), .A2(n2564), .ZN(n3810) );
  OR2_X1 U33220 ( .A1(n3810), .A2(n2609), .ZN(n2567) );
  AOI22_X1 U33230 ( .A1(n2347), .A2(REG2_REG_20__SCAN_IN), .B1(n2645), .B2(
        REG0_REG_20__SCAN_IN), .ZN(n2566) );
  INV_X1 U33240 ( .A(DATAI_20_), .ZN(n2568) );
  NAND2_X1 U33250 ( .A1(n4241), .A2(n4105), .ZN(n3465) );
  NOR2_X1 U33260 ( .A1(n4241), .A2(n4105), .ZN(n3466) );
  XNOR2_X1 U33270 ( .A(n2576), .B(REG3_REG_22__SCAN_IN), .ZN(n4075) );
  NAND2_X1 U33280 ( .A1(n4075), .A2(n2355), .ZN(n2573) );
  INV_X1 U33290 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4237) );
  NAND2_X1 U33300 ( .A1(n2645), .A2(REG0_REG_22__SCAN_IN), .ZN(n2570) );
  NAND2_X1 U33310 ( .A1(n2384), .A2(REG2_REG_22__SCAN_IN), .ZN(n2569) );
  OAI211_X1 U33320 ( .C1(n2365), .C2(n4237), .A(n2570), .B(n2569), .ZN(n2571)
         );
  INV_X1 U33330 ( .A(n2571), .ZN(n2572) );
  NAND2_X1 U33340 ( .A1(n4090), .A2(n4072), .ZN(n2667) );
  NAND2_X1 U33350 ( .A1(n4051), .A2(n2667), .ZN(n4077) );
  NAND2_X2 U33360 ( .A1(n4078), .A2(n4077), .ZN(n4079) );
  NAND2_X2 U33370 ( .A1(n4079), .A2(n2287), .ZN(n4047) );
  INV_X1 U33380 ( .A(n2576), .ZN(n2575) );
  AND2_X1 U33390 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2574) );
  INV_X1 U33400 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3818) );
  INV_X1 U33410 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4627) );
  OAI21_X1 U33420 ( .B1(n2576), .B2(n3818), .A(n4627), .ZN(n2577) );
  NAND2_X1 U33430 ( .A1(n2585), .A2(n2577), .ZN(n4059) );
  OR2_X1 U33440 ( .A1(n4059), .A2(n2609), .ZN(n2582) );
  INV_X1 U33450 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4232) );
  NAND2_X1 U33460 ( .A1(n2347), .A2(REG2_REG_23__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U33470 ( .A1(n2645), .A2(REG0_REG_23__SCAN_IN), .ZN(n2578) );
  OAI211_X1 U33480 ( .C1(n4232), .C2(n3419), .A(n2579), .B(n2578), .ZN(n2580)
         );
  INV_X1 U33490 ( .A(n2580), .ZN(n2581) );
  NAND2_X1 U33500 ( .A1(n3819), .A2(n4058), .ZN(n2584) );
  NAND2_X1 U33510 ( .A1(n2585), .A2(n4635), .ZN(n2586) );
  NAND2_X1 U33520 ( .A1(n4039), .A2(n2355), .ZN(n2591) );
  INV_X1 U3353 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4228) );
  NAND2_X1 U33540 ( .A1(n2347), .A2(REG2_REG_24__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U3355 ( .A1(n2645), .A2(REG0_REG_24__SCAN_IN), .ZN(n2587) );
  OAI211_X1 U3356 ( .C1(n4228), .C2(n3419), .A(n2588), .B(n2587), .ZN(n2589)
         );
  INV_X1 U3357 ( .A(n2589), .ZN(n2590) );
  XNOR2_X1 U3358 ( .A(n2597), .B(REG3_REG_25__SCAN_IN), .ZN(n4024) );
  NAND2_X1 U3359 ( .A1(n4024), .A2(n2355), .ZN(n2596) );
  INV_X1 U3360 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4219) );
  NAND2_X1 U3361 ( .A1(n2347), .A2(REG2_REG_25__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U3362 ( .A1(n2645), .A2(REG0_REG_25__SCAN_IN), .ZN(n2592) );
  OAI211_X1 U3363 ( .C1(n4219), .C2(n3419), .A(n2593), .B(n2592), .ZN(n2594)
         );
  INV_X1 U3364 ( .A(n2594), .ZN(n2595) );
  INV_X1 U3365 ( .A(DATAI_25_), .ZN(n4604) );
  INV_X1 U3366 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4541) );
  INV_X1 U3367 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3838) );
  OAI21_X1 U3368 ( .B1(n2597), .B2(n4541), .A(n3838), .ZN(n2600) );
  INV_X1 U3369 ( .A(n2597), .ZN(n2599) );
  AND2_X1 U3370 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2598) );
  NAND2_X1 U3371 ( .A1(n2599), .A2(n2598), .ZN(n2607) );
  NAND2_X1 U3372 ( .A1(n2600), .A2(n2607), .ZN(n3837) );
  INV_X1 U3373 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4210) );
  NAND2_X1 U3374 ( .A1(n2384), .A2(REG2_REG_26__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U3375 ( .A1(n2645), .A2(REG0_REG_26__SCAN_IN), .ZN(n2601) );
  OAI211_X1 U3376 ( .C1(n4210), .C2(n3419), .A(n2602), .B(n2601), .ZN(n2603)
         );
  INV_X1 U3377 ( .A(n2603), .ZN(n2604) );
  NAND2_X1 U3378 ( .A1(n3428), .A2(DATAI_26_), .ZN(n4010) );
  NOR2_X1 U3379 ( .A1(n4216), .A2(n4010), .ZN(n2606) );
  INV_X1 U3380 ( .A(n4010), .ZN(n2671) );
  OAI22_X2 U3381 ( .A1(n3999), .A2(n2606), .B1(n2671), .B2(n4200), .ZN(n3984)
         );
  INV_X1 U3382 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4554) );
  NAND2_X1 U3383 ( .A1(n2607), .A2(n4554), .ZN(n2608) );
  NAND2_X1 U3384 ( .A1(n2617), .A2(n2608), .ZN(n3737) );
  INV_X1 U3385 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4206) );
  NAND2_X1 U3386 ( .A1(n2347), .A2(REG2_REG_27__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U3387 ( .A1(n2645), .A2(REG0_REG_27__SCAN_IN), .ZN(n2610) );
  OAI211_X1 U3388 ( .C1(n4206), .C2(n3419), .A(n2611), .B(n2610), .ZN(n2612)
         );
  INV_X1 U3389 ( .A(n2612), .ZN(n2613) );
  INV_X1 U3390 ( .A(DATAI_27_), .ZN(n2615) );
  NOR2_X1 U3391 ( .A1(n3861), .A2(n4199), .ZN(n2616) );
  INV_X1 U3392 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U3393 ( .A1(n2617), .A2(n3715), .ZN(n2618) );
  NAND2_X1 U3394 ( .A1(n3726), .A2(n2355), .ZN(n2624) );
  INV_X1 U3395 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2621) );
  NAND2_X1 U3396 ( .A1(n2347), .A2(REG2_REG_28__SCAN_IN), .ZN(n2620) );
  NAND2_X1 U3397 ( .A1(n2645), .A2(REG0_REG_28__SCAN_IN), .ZN(n2619) );
  OAI211_X1 U3398 ( .C1(n2621), .C2(n3419), .A(n2620), .B(n2619), .ZN(n2622)
         );
  INV_X1 U3399 ( .A(n2622), .ZN(n2623) );
  INV_X1 U3400 ( .A(DATAI_28_), .ZN(n2625) );
  NAND2_X1 U3401 ( .A1(n4202), .A2(n2720), .ZN(n3425) );
  INV_X1 U3402 ( .A(n2720), .ZN(n3729) );
  NAND2_X1 U3403 ( .A1(n3990), .A2(n3729), .ZN(n3422) );
  NAND2_X1 U3404 ( .A1(n3425), .A2(n3422), .ZN(n2721) );
  XNOR2_X1 U3405 ( .A(n2722), .B(n2721), .ZN(n3735) );
  NAND2_X1 U3406 ( .A1(n2635), .A2(IR_REG_31__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U3407 ( .A1(n2631), .A2(n2630), .ZN(n2632) );
  INV_X1 U3408 ( .A(n2640), .ZN(n2764) );
  NAND2_X1 U3409 ( .A1(n2636), .A2(n2628), .ZN(n2683) );
  NAND2_X1 U3410 ( .A1(n2683), .A2(IR_REG_31__SCAN_IN), .ZN(n2638) );
  XNOR2_X1 U3411 ( .A(n2908), .B(n3581), .ZN(n2639) );
  NAND2_X1 U3412 ( .A1(n2639), .A2(n3963), .ZN(n4111) );
  AND2_X1 U3413 ( .A1(n2640), .A2(n4352), .ZN(n2851) );
  INV_X1 U3414 ( .A(n4502), .ZN(n3281) );
  NOR2_X1 U3415 ( .A1(n2046), .A2(n2642), .ZN(n2641) );
  MUX2_X1 U3416 ( .A(n2642), .B(n2641), .S(IR_REG_28__SCAN_IN), .Z(n2643) );
  OR2_X1 U3417 ( .A1(n2643), .A2(n2086), .ZN(n2897) );
  INV_X1 U3418 ( .A(n3470), .ZN(n4351) );
  INV_X1 U3419 ( .A(n2882), .ZN(n2773) );
  INV_X1 U3420 ( .A(n2644), .ZN(n3974) );
  INV_X1 U3421 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2732) );
  NAND2_X1 U3422 ( .A1(n2347), .A2(REG2_REG_29__SCAN_IN), .ZN(n2647) );
  NAND2_X1 U3423 ( .A1(n2645), .A2(REG0_REG_29__SCAN_IN), .ZN(n2646) );
  OAI211_X1 U3424 ( .C1(n2732), .C2(n3419), .A(n2647), .B(n2646), .ZN(n2648)
         );
  AOI21_X1 U3425 ( .B1(n3974), .B2(n2355), .A(n2648), .ZN(n3716) );
  INV_X1 U3426 ( .A(n3716), .ZN(n3860) );
  NOR2_X2 U3427 ( .A1(n2897), .A2(n2882), .ZN(n4240) );
  NAND2_X1 U3428 ( .A1(n2889), .A2(n3470), .ZN(n2881) );
  OAI22_X1 U3429 ( .A1(n4005), .A2(n4288), .B1(n4066), .B2(n3729), .ZN(n2649)
         );
  AOI21_X1 U3430 ( .B1(n4284), .B2(n3860), .A(n2649), .ZN(n2676) );
  INV_X1 U3431 ( .A(n2857), .ZN(n2943) );
  NAND2_X1 U3432 ( .A1(n2943), .A2(n2948), .ZN(n3514) );
  NAND2_X1 U3433 ( .A1(n2743), .A2(n3520), .ZN(n2978) );
  NAND2_X1 U3434 ( .A1(n3041), .A2(n2980), .ZN(n3525) );
  NAND2_X1 U3435 ( .A1(n3876), .A2(n3011), .ZN(n3522) );
  AND2_X1 U3436 ( .A1(n3525), .A2(n3522), .ZN(n3483) );
  NAND2_X1 U3437 ( .A1(n2978), .A2(n3483), .ZN(n2977) );
  INV_X1 U3438 ( .A(n3526), .ZN(n2652) );
  AND2_X1 U3439 ( .A1(n3874), .A2(n3121), .ZN(n3048) );
  NAND2_X1 U3440 ( .A1(n3133), .A2(n3114), .ZN(n3503) );
  NAND2_X1 U3441 ( .A1(n3873), .A2(n3134), .ZN(n3528) );
  INV_X1 U3442 ( .A(n3873), .ZN(n3176) );
  NAND2_X1 U3443 ( .A1(n3176), .A2(n3084), .ZN(n3532) );
  NAND2_X1 U3444 ( .A1(n2653), .A2(n3532), .ZN(n3094) );
  INV_X1 U3445 ( .A(n2654), .ZN(n2655) );
  NAND2_X1 U3446 ( .A1(n3252), .A2(n3215), .ZN(n3538) );
  NAND2_X1 U3447 ( .A1(n3870), .A2(n3205), .ZN(n3535) );
  AND2_X1 U3448 ( .A1(n3869), .A2(n3253), .ZN(n3140) );
  NAND2_X1 U3449 ( .A1(n3274), .A2(n3247), .ZN(n3539) );
  NAND2_X1 U3450 ( .A1(n3868), .A2(n3275), .ZN(n3502) );
  NAND2_X1 U3451 ( .A1(n3150), .A2(n3502), .ZN(n2656) );
  NAND2_X1 U3452 ( .A1(n3359), .A2(n3266), .ZN(n3507) );
  NAND2_X1 U3453 ( .A1(n2656), .A2(n3507), .ZN(n3294) );
  NAND2_X1 U3454 ( .A1(n3866), .A2(n3400), .ZN(n3309) );
  NAND2_X1 U3455 ( .A1(n3865), .A2(n3606), .ZN(n2657) );
  NAND2_X1 U3456 ( .A1(n3309), .A2(n2657), .ZN(n3543) );
  INV_X1 U3457 ( .A(n3293), .ZN(n3546) );
  NOR2_X1 U34580 ( .A1(n3543), .A2(n3546), .ZN(n2658) );
  NAND2_X1 U34590 ( .A1(n3294), .A2(n2658), .ZN(n2662) );
  NAND2_X1 U3460 ( .A1(n3605), .A2(n3411), .ZN(n3310) );
  NAND2_X1 U3461 ( .A1(n3291), .A2(n3310), .ZN(n2661) );
  INV_X1 U3462 ( .A(n3543), .ZN(n2660) );
  NOR2_X1 U3463 ( .A1(n3865), .A2(n3606), .ZN(n2659) );
  AOI21_X1 U3464 ( .B1(n2661), .B2(n2660), .A(n2659), .ZN(n3547) );
  NAND2_X1 U3465 ( .A1(n2662), .A2(n3547), .ZN(n3440) );
  INV_X1 U3466 ( .A(n3324), .ZN(n3481) );
  NAND2_X1 U34670 ( .A1(n3440), .A2(n3481), .ZN(n2663) );
  NAND2_X1 U3468 ( .A1(n2663), .A2(n3432), .ZN(n3365) );
  NAND2_X1 U34690 ( .A1(n4269), .A2(n4283), .ZN(n3439) );
  NAND2_X1 U3470 ( .A1(n3863), .A2(n3852), .ZN(n3508) );
  NAND2_X1 U34710 ( .A1(n3439), .A2(n3508), .ZN(n3493) );
  INV_X1 U3472 ( .A(n3586), .ZN(n3594) );
  AND2_X1 U34730 ( .A1(n4153), .A2(n4186), .ZN(n3434) );
  NAND2_X1 U3474 ( .A1(n3862), .A2(n4137), .ZN(n3471) );
  NAND2_X1 U34750 ( .A1(n3471), .A2(n4127), .ZN(n3433) );
  INV_X1 U3476 ( .A(n4105), .ZN(n4115) );
  NAND2_X1 U34770 ( .A1(n4241), .A2(n4115), .ZN(n3435) );
  NAND2_X1 U3478 ( .A1(n4274), .A2(n4260), .ZN(n4124) );
  AND2_X1 U34790 ( .A1(n4126), .A2(n4124), .ZN(n2664) );
  OR2_X1 U3480 ( .A1(n3862), .A2(n4137), .ZN(n3472) );
  OAI21_X1 U34810 ( .B1(n3433), .B2(n2664), .A(n3472), .ZN(n4100) );
  NOR2_X1 U3482 ( .A1(n4241), .A2(n4115), .ZN(n2665) );
  OR2_X1 U34830 ( .A1(n4100), .A2(n2665), .ZN(n2666) );
  NAND2_X1 U3484 ( .A1(n2666), .A2(n3435), .ZN(n3554) );
  OR2_X1 U34850 ( .A1(n4106), .A2(n4094), .ZN(n3489) );
  AND2_X1 U3486 ( .A1(n4051), .A2(n3489), .ZN(n3555) );
  INV_X1 U34870 ( .A(n3555), .ZN(n2669) );
  NAND2_X1 U3488 ( .A1(n4222), .A2(n4058), .ZN(n3462) );
  AND2_X1 U34890 ( .A1(n3462), .A2(n2667), .ZN(n3560) );
  AND2_X1 U3490 ( .A1(n4106), .A2(n4094), .ZN(n4048) );
  NAND2_X1 U34910 ( .A1(n4051), .A2(n4048), .ZN(n2668) );
  AND2_X1 U3492 ( .A1(n3560), .A2(n2668), .ZN(n3446) );
  OAI21_X1 U34930 ( .B1(n4084), .B2(n2669), .A(n3446), .ZN(n2670) );
  NAND2_X1 U3494 ( .A1(n2670), .A2(n3463), .ZN(n4032) );
  NOR2_X1 U34950 ( .A1(n4213), .A2(n4042), .ZN(n3461) );
  NAND2_X1 U3496 ( .A1(n4216), .A2(n2671), .ZN(n2672) );
  OR2_X1 U34970 ( .A1(n4038), .A2(n4027), .ZN(n4000) );
  AND2_X1 U3498 ( .A1(n2672), .A2(n4000), .ZN(n2673) );
  INV_X1 U34990 ( .A(n2673), .ZN(n3557) );
  NAND2_X1 U3500 ( .A1(n4038), .A2(n4027), .ZN(n3459) );
  NAND2_X1 U35010 ( .A1(n4213), .A2(n4042), .ZN(n4016) );
  NAND2_X1 U3502 ( .A1(n3459), .A2(n4016), .ZN(n4001) );
  AND2_X1 U35030 ( .A1(n4200), .A2(n4010), .ZN(n3423) );
  AOI21_X1 U3504 ( .B1(n2673), .B2(n4001), .A(n3423), .ZN(n3563) );
  XNOR2_X1 U35050 ( .A(n3861), .B(n3994), .ZN(n3985) );
  NAND2_X1 U35060 ( .A1(n4005), .A2(n4199), .ZN(n3424) );
  INV_X1 U35070 ( .A(n2721), .ZN(n3458) );
  XNOR2_X1 U35080 ( .A(n2723), .B(n3458), .ZN(n2675) );
  NAND2_X1 U35090 ( .A1(n3581), .A2(n4352), .ZN(n2674) );
  NAND2_X1 U35100 ( .A1(n4351), .A2(n2764), .ZN(n3456) );
  NAND2_X1 U35110 ( .A1(n2675), .A2(n4169), .ZN(n3730) );
  OAI211_X1 U35120 ( .C1(n3735), .C2(n4280), .A(n2676), .B(n3730), .ZN(n2717)
         );
  INV_X1 U35130 ( .A(n2677), .ZN(n2681) );
  NAND2_X1 U35140 ( .A1(n2679), .A2(IR_REG_31__SCAN_IN), .ZN(n2680) );
  MUX2_X1 U35150 ( .A(IR_REG_31__SCAN_IN), .B(n2680), .S(IR_REG_25__SCAN_IN), 
        .Z(n2682) );
  NAND2_X1 U35160 ( .A1(n2682), .A2(n2681), .ZN(n2762) );
  NAND2_X1 U35170 ( .A1(n2762), .A2(B_REG_SCAN_IN), .ZN(n2686) );
  MUX2_X1 U35180 ( .A(n2686), .B(B_REG_SCAN_IN), .S(n2688), .Z(n2687) );
  NAND2_X1 U35190 ( .A1(n2706), .A2(n2762), .ZN(n2777) );
  NAND2_X1 U35200 ( .A1(n2884), .A2(n2777), .ZN(n2705) );
  XNOR2_X1 U35210 ( .A(n2690), .B(n2691), .ZN(n2772) );
  NAND2_X1 U35220 ( .A1(n4502), .A2(n3470), .ZN(n2751) );
  AND2_X1 U35230 ( .A1(n2640), .A2(n3963), .ZN(n2880) );
  NAND2_X1 U35240 ( .A1(n2751), .A2(n2887), .ZN(n2692) );
  NOR2_X1 U35250 ( .A1(n2895), .A2(n2692), .ZN(n2704) );
  NOR4_X1 U35260 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2696) );
  NOR4_X1 U35270 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2695) );
  NOR4_X1 U35280 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2694) );
  NOR4_X1 U35290 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2693) );
  NAND4_X1 U35300 ( .A1(n2696), .A2(n2695), .A3(n2694), .A4(n2693), .ZN(n2702)
         );
  NOR2_X1 U35310 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .ZN(n2700) );
  NOR4_X1 U35320 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2699) );
  NOR4_X1 U35330 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2698) );
  NOR4_X1 U35340 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2697) );
  NAND4_X1 U35350 ( .A1(n2700), .A2(n2699), .A3(n2698), .A4(n2697), .ZN(n2701)
         );
  NOR2_X1 U35360 ( .A1(n2702), .A2(n2701), .ZN(n2703) );
  NAND3_X1 U35370 ( .A1(n2705), .A2(n2704), .A3(n2747), .ZN(n2715) );
  NAND2_X1 U35380 ( .A1(n3722), .A2(n2706), .ZN(n2707) );
  INV_X1 U35390 ( .A(n2948), .ZN(n2849) );
  NAND2_X1 U35400 ( .A1(n2905), .A2(n2849), .ZN(n2950) );
  NOR2_X1 U35410 ( .A1(n2950), .A2(n2984), .ZN(n2974) );
  INV_X1 U35420 ( .A(n3988), .ZN(n2710) );
  INV_X1 U35430 ( .A(n2881), .ZN(n2848) );
  INV_X1 U35440 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2711) );
  NAND2_X1 U35450 ( .A1(n2717), .A2(n4517), .ZN(n2718) );
  NAND2_X1 U35460 ( .A1(n2719), .A2(n2718), .ZN(U3546) );
  NAND2_X1 U35470 ( .A1(n3428), .A2(DATAI_29_), .ZN(n3979) );
  XOR2_X1 U35480 ( .A(n3979), .B(n3716), .Z(n3501) );
  XNOR2_X1 U35490 ( .A(n2724), .B(n3501), .ZN(n2730) );
  NOR2_X1 U35500 ( .A1(n2726), .A2(n2725), .ZN(n2868) );
  AOI21_X1 U35510 ( .B1(B_REG_SCAN_IN), .B2(n2868), .A(n4273), .ZN(n3968) );
  INV_X1 U35520 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2729) );
  NAND2_X1 U35530 ( .A1(n2384), .A2(REG2_REG_30__SCAN_IN), .ZN(n2728) );
  NAND2_X1 U35540 ( .A1(n2645), .A2(REG0_REG_30__SCAN_IN), .ZN(n2727) );
  OAI211_X1 U35550 ( .C1(n3419), .C2(n2729), .A(n2728), .B(n2727), .ZN(n3859)
         );
  NAND2_X1 U35560 ( .A1(n3990), .A2(n4240), .ZN(n2731) );
  MUX2_X1 U35570 ( .A(n2732), .B(n2056), .S(n4517), .Z(n2737) );
  INV_X1 U35580 ( .A(n3979), .ZN(n3427) );
  NAND2_X1 U35590 ( .A1(n2054), .A2(n3427), .ZN(n2733) );
  NAND2_X1 U35600 ( .A1(n2051), .A2(n2733), .ZN(n3977) );
  INV_X1 U35610 ( .A(n3977), .ZN(n2735) );
  NAND2_X1 U35620 ( .A1(n2735), .A2(n2734), .ZN(n2736) );
  NAND2_X1 U35630 ( .A1(n2737), .A2(n2736), .ZN(U3547) );
  NAND2_X1 U35640 ( .A1(n2740), .A2(n2739), .ZN(U3515) );
  INV_X2 U35650 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U35660 ( .A1(n2742), .A2(n2741), .ZN(n2988) );
  INV_X1 U35670 ( .A(n4111), .ZN(n3211) );
  NAND2_X1 U35680 ( .A1(n2988), .A2(n3211), .ZN(n2746) );
  NAND2_X1 U35690 ( .A1(n2744), .A2(n4169), .ZN(n2745) );
  NAND2_X1 U35700 ( .A1(n2746), .A2(n2745), .ZN(n2986) );
  INV_X1 U35710 ( .A(n2887), .ZN(n2748) );
  NOR2_X1 U35720 ( .A1(n2895), .A2(n2748), .ZN(n2750) );
  NAND4_X1 U35730 ( .A1(n2885), .A2(n2750), .A3(n2749), .A4(n2884), .ZN(n2752)
         );
  MUX2_X1 U35740 ( .A(REG2_REG_2__SCAN_IN), .B(n2986), .S(n4164), .Z(n2760) );
  NAND2_X1 U35750 ( .A1(n2856), .A2(n4352), .ZN(n3007) );
  INV_X1 U35760 ( .A(n3007), .ZN(n2753) );
  AND2_X1 U35770 ( .A1(n4164), .A2(n2753), .ZN(n4474) );
  INV_X1 U35780 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3888) );
  NOR2_X1 U35790 ( .A1(n4468), .A2(n3888), .ZN(n2754) );
  AOI21_X1 U35800 ( .B1(n2988), .B2(n4474), .A(n2754), .ZN(n2758) );
  NAND2_X1 U35810 ( .A1(n4164), .A2(n4282), .ZN(n4185) );
  INV_X1 U3582 ( .A(n4185), .ZN(n3327) );
  AOI22_X1 U3583 ( .A1(n3327), .A2(n2984), .B1(n4178), .B2(n3876), .ZN(n2757)
         );
  NAND2_X1 U3584 ( .A1(n4164), .A2(n3963), .ZN(n4160) );
  XNOR2_X1 U3585 ( .A(n2950), .B(n2927), .ZN(n2990) );
  NAND2_X1 U3586 ( .A1(n4473), .A2(n2990), .ZN(n2756) );
  NAND2_X1 U3587 ( .A1(n4179), .A2(n3877), .ZN(n2755) );
  NAND4_X1 U3588 ( .A1(n2758), .A2(n2757), .A3(n2756), .A4(n2755), .ZN(n2759)
         );
  OR2_X1 U3589 ( .A1(n2760), .A2(n2759), .ZN(U3288) );
  NAND2_X1 U3590 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2761) );
  OAI21_X1 U3591 ( .B1(n2762), .B2(U3149), .A(n2761), .ZN(U3327) );
  INV_X1 U3592 ( .A(DATAI_26_), .ZN(n4552) );
  NAND2_X1 U3593 ( .A1(n3721), .A2(STATE_REG_SCAN_IN), .ZN(n2763) );
  OAI21_X1 U3594 ( .B1(STATE_REG_SCAN_IN), .B2(n4552), .A(n2763), .ZN(U3326)
         );
  NAND2_X1 U3595 ( .A1(n2764), .A2(STATE_REG_SCAN_IN), .ZN(n2765) );
  OAI21_X1 U3596 ( .B1(STATE_REG_SCAN_IN), .B2(n2568), .A(n2765), .ZN(U3332)
         );
  INV_X1 U3597 ( .A(DATAI_22_), .ZN(n4644) );
  NAND2_X1 U3598 ( .A1(n3581), .A2(STATE_REG_SCAN_IN), .ZN(n2766) );
  OAI21_X1 U3599 ( .B1(STATE_REG_SCAN_IN), .B2(n4644), .A(n2766), .ZN(U3330)
         );
  INV_X1 U3600 ( .A(DATAI_24_), .ZN(n4542) );
  NAND2_X1 U3601 ( .A1(n2688), .A2(STATE_REG_SCAN_IN), .ZN(n2767) );
  OAI21_X1 U3602 ( .B1(STATE_REG_SCAN_IN), .B2(n4542), .A(n2767), .ZN(U3328)
         );
  NAND2_X1 U3603 ( .A1(n2868), .A2(STATE_REG_SCAN_IN), .ZN(n2768) );
  OAI21_X1 U3604 ( .B1(STATE_REG_SCAN_IN), .B2(n2615), .A(n2768), .ZN(U3325)
         );
  INV_X1 U3605 ( .A(DATAI_31_), .ZN(n4677) );
  OR4_X1 U3606 ( .A1(n2309), .A2(IR_REG_30__SCAN_IN), .A3(n2642), .A4(U3149), 
        .ZN(n2769) );
  OAI21_X1 U3607 ( .B1(STATE_REG_SCAN_IN), .B2(n4677), .A(n2769), .ZN(U3321)
         );
  INV_X1 U3608 ( .A(n2897), .ZN(n2919) );
  NAND2_X1 U3609 ( .A1(n2919), .A2(STATE_REG_SCAN_IN), .ZN(n2770) );
  OAI21_X1 U3610 ( .B1(STATE_REG_SCAN_IN), .B2(n2625), .A(n2770), .ZN(U3324)
         );
  OR2_X1 U3611 ( .A1(n2772), .A2(U3149), .ZN(n3583) );
  NAND2_X1 U3612 ( .A1(n2895), .A2(n3583), .ZN(n2782) );
  AOI21_X1 U3613 ( .B1(n2773), .B2(n2772), .A(n2771), .ZN(n2781) );
  INV_X1 U3614 ( .A(n2781), .ZN(n2774) );
  NOR2_X1 U3615 ( .A1(n4460), .A2(U4043), .ZN(U3148) );
  INV_X1 U3616 ( .A(n2895), .ZN(n2775) );
  INV_X1 U3617 ( .A(D_REG_1__SCAN_IN), .ZN(n2780) );
  INV_X1 U3618 ( .A(n2777), .ZN(n2779) );
  AOI22_X1 U3619 ( .A1(n4479), .A2(n2780), .B1(n2779), .B2(n2778), .ZN(U3459)
         );
  INV_X1 U3620 ( .A(n2797), .ZN(n2785) );
  INV_X1 U3621 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2855) );
  AOI21_X1 U3622 ( .B1(n2868), .B2(n2855), .A(n2897), .ZN(n2870) );
  OAI21_X1 U3623 ( .B1(REG1_REG_0__SCAN_IN), .B2(n2868), .A(n2870), .ZN(n2783)
         );
  MUX2_X1 U3624 ( .A(n2783), .B(n2870), .S(IR_REG_0__SCAN_IN), .Z(n2784) );
  INV_X1 U3625 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2902) );
  OAI22_X1 U3626 ( .A1(n2785), .A2(n2784), .B1(STATE_REG_SCAN_IN), .B2(n2902), 
        .ZN(n2786) );
  AOI21_X1 U3627 ( .B1(n4460), .B2(ADDR_REG_0__SCAN_IN), .A(n2786), .ZN(n2788)
         );
  INV_X1 U3628 ( .A(n2868), .ZN(n2795) );
  NAND3_X1 U3629 ( .A1(n4462), .A2(IR_REG_0__SCAN_IN), .A3(n2357), .ZN(n2787)
         );
  NAND2_X1 U3630 ( .A1(n2788), .A2(n2787), .ZN(U3240) );
  INV_X1 U3631 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3893) );
  INV_X1 U3632 ( .A(n2048), .ZN(n3891) );
  MUX2_X1 U3633 ( .A(REG2_REG_2__SCAN_IN), .B(n3893), .S(n2047), .Z(n2792) );
  INV_X1 U3634 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2789) );
  AND2_X1 U3635 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2790)
         );
  NAND2_X1 U3636 ( .A1(n3895), .A2(n3894), .ZN(n2791) );
  INV_X1 U3637 ( .A(n4358), .ZN(n2804) );
  INV_X1 U3638 ( .A(n4357), .ZN(n2876) );
  XNOR2_X1 U3639 ( .A(n2793), .B(n2876), .ZN(n2871) );
  INV_X1 U3640 ( .A(n2793), .ZN(n2794) );
  MUX2_X1 U3641 ( .A(REG2_REG_5__SCAN_IN), .B(n2399), .S(n2818), .Z(n2796) );
  NOR2_X1 U3642 ( .A1(n2897), .A2(n2795), .ZN(n3578) );
  AOI211_X1 U3643 ( .C1(n2087), .C2(n2796), .A(n2813), .B(n4456), .ZN(n2800)
         );
  INV_X1 U3644 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4645) );
  NOR2_X1 U3645 ( .A1(STATE_REG_SCAN_IN), .A2(n4645), .ZN(n3123) );
  AOI21_X1 U3646 ( .B1(n4460), .B2(ADDR_REG_5__SCAN_IN), .A(n3123), .ZN(n2798)
         );
  OAI21_X1 U3647 ( .B1(n4467), .B2(n2818), .A(n2798), .ZN(n2799) );
  NOR2_X1 U3648 ( .A1(n2800), .A2(n2799), .ZN(n2812) );
  XNOR2_X1 U3649 ( .A(n2818), .B(REG1_REG_5__SCAN_IN), .ZN(n2810) );
  XNOR2_X1 U3650 ( .A(n2048), .B(n2801), .ZN(n3901) );
  AND2_X1 U3651 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3880)
         );
  NAND2_X1 U3652 ( .A1(n3881), .A2(n3880), .ZN(n3879) );
  NAND2_X1 U3653 ( .A1(n3879), .A2(n2802), .ZN(n3900) );
  NAND2_X1 U3654 ( .A1(n3901), .A2(n3900), .ZN(n3899) );
  NAND2_X1 U3655 ( .A1(n2048), .A2(REG1_REG_2__SCAN_IN), .ZN(n2803) );
  NAND2_X1 U3656 ( .A1(n3899), .A2(n2803), .ZN(n2805) );
  XNOR2_X1 U3657 ( .A(n2805), .B(n2804), .ZN(n3908) );
  NAND2_X1 U3658 ( .A1(n3908), .A2(REG1_REG_3__SCAN_IN), .ZN(n3907) );
  NAND2_X1 U3659 ( .A1(n2805), .A2(n4358), .ZN(n2806) );
  NAND2_X1 U3660 ( .A1(n3907), .A2(n2806), .ZN(n2807) );
  INV_X1 U3661 ( .A(n2807), .ZN(n2808) );
  XNOR2_X1 U3662 ( .A(n2807), .B(n2876), .ZN(n2873) );
  NAND2_X1 U3663 ( .A1(n2873), .A2(REG1_REG_4__SCAN_IN), .ZN(n2872) );
  OAI21_X1 U3664 ( .B1(n2808), .B2(n2876), .A(n2872), .ZN(n2809) );
  NAND2_X1 U3665 ( .A1(n2809), .A2(n2810), .ZN(n2816) );
  OAI211_X1 U3666 ( .C1(n2810), .C2(n2809), .A(n4462), .B(n2816), .ZN(n2811)
         );
  NAND2_X1 U3667 ( .A1(n2812), .A2(n2811), .ZN(U3245) );
  INV_X1 U3668 ( .A(n2818), .ZN(n4356) );
  XNOR2_X1 U3669 ( .A(n2829), .B(n4355), .ZN(n2831) );
  XNOR2_X1 U3670 ( .A(n2831), .B(REG2_REG_6__SCAN_IN), .ZN(n2824) );
  INV_X1 U3671 ( .A(n4467), .ZN(n3906) );
  NOR2_X1 U3672 ( .A1(STATE_REG_SCAN_IN), .A2(n2814), .ZN(n3136) );
  AOI21_X1 U3673 ( .B1(n4460), .B2(ADDR_REG_6__SCAN_IN), .A(n3136), .ZN(n2815)
         );
  INV_X1 U3674 ( .A(n2815), .ZN(n2822) );
  OAI21_X1 U3675 ( .B1(n2818), .B2(n2817), .A(n2816), .ZN(n2826) );
  XNOR2_X1 U3676 ( .A(n2826), .B(n4355), .ZN(n2820) );
  NOR2_X1 U3677 ( .A1(n2820), .A2(n2416), .ZN(n2825) );
  INV_X1 U3678 ( .A(n4462), .ZN(n2819) );
  AOI211_X1 U3679 ( .C1(n2820), .C2(n2416), .A(n2825), .B(n2819), .ZN(n2821)
         );
  AOI211_X1 U3680 ( .C1(n3906), .C2(n4355), .A(n2822), .B(n2821), .ZN(n2823)
         );
  OAI21_X1 U3681 ( .B1(n2824), .B2(n4456), .A(n2823), .ZN(U3246) );
  MUX2_X1 U3682 ( .A(REG1_REG_7__SCAN_IN), .B(n2428), .S(n4354), .Z(n2827) );
  XNOR2_X1 U3683 ( .A(n2840), .B(n2827), .ZN(n2836) );
  INV_X1 U3684 ( .A(n4354), .ZN(n2838) );
  INV_X1 U3685 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4606) );
  NOR2_X1 U3686 ( .A1(STATE_REG_SCAN_IN), .A2(n4606), .ZN(n3179) );
  AOI21_X1 U3687 ( .B1(n4460), .B2(ADDR_REG_7__SCAN_IN), .A(n3179), .ZN(n2828)
         );
  OAI21_X1 U3688 ( .B1(n4467), .B2(n2838), .A(n2828), .ZN(n2835) );
  INV_X1 U3689 ( .A(n2829), .ZN(n2830) );
  INV_X1 U3690 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3102) );
  MUX2_X1 U3691 ( .A(n3102), .B(REG2_REG_7__SCAN_IN), .S(n4354), .Z(n2832) );
  NOR2_X1 U3692 ( .A1(n2833), .A2(n2832), .ZN(n2842) );
  AOI211_X1 U3693 ( .C1(n2833), .C2(n2832), .A(n4456), .B(n2842), .ZN(n2834)
         );
  AOI211_X1 U3694 ( .C1(n4462), .C2(n2836), .A(n2835), .B(n2834), .ZN(n2837)
         );
  INV_X1 U3695 ( .A(n2837), .ZN(U3247) );
  NOR2_X1 U3696 ( .A1(n4354), .A2(REG1_REG_7__SCAN_IN), .ZN(n2839) );
  XOR2_X1 U3697 ( .A(REG1_REG_8__SCAN_IN), .B(n3936), .Z(n2841) );
  NAND2_X1 U3698 ( .A1(n2841), .A2(n4462), .ZN(n2847) );
  AOI21_X1 U3699 ( .B1(n4354), .B2(REG2_REG_7__SCAN_IN), .A(n2842), .ZN(n3918)
         );
  XNOR2_X1 U3700 ( .A(n3918), .B(n4353), .ZN(n3919) );
  XNOR2_X1 U3701 ( .A(REG2_REG_8__SCAN_IN), .B(n3919), .ZN(n2843) );
  NAND2_X1 U3702 ( .A1(n4406), .A2(n2843), .ZN(n2844) );
  NAND2_X1 U3703 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3196) );
  NAND2_X1 U3704 ( .A1(n2844), .A2(n3196), .ZN(n2845) );
  AOI21_X1 U3705 ( .B1(n4460), .B2(ADDR_REG_8__SCAN_IN), .A(n2845), .ZN(n2846)
         );
  OAI211_X1 U3706 ( .C1(n4467), .C2(n4353), .A(n2847), .B(n2846), .ZN(U3248)
         );
  NAND2_X1 U3707 ( .A1(n2948), .A2(n2848), .ZN(n4494) );
  NAND2_X1 U3708 ( .A1(n2857), .A2(n2849), .ZN(n3516) );
  NAND2_X1 U3709 ( .A1(n3514), .A2(n3516), .ZN(n4498) );
  NAND2_X1 U3710 ( .A1(n4111), .A2(n4070), .ZN(n2850) );
  AOI22_X1 U3711 ( .A1(n4498), .A2(n2850), .B1(n4284), .B2(n3877), .ZN(n4495)
         );
  OAI21_X1 U3712 ( .B1(n2851), .B2(n4494), .A(n4495), .ZN(n2852) );
  AOI22_X1 U3713 ( .A1(n2852), .A2(n4164), .B1(REG3_REG_0__SCAN_IN), .B2(n4181), .ZN(n2854) );
  NAND2_X1 U3714 ( .A1(n4474), .A2(n4498), .ZN(n2853) );
  OAI211_X1 U3715 ( .C1(n4164), .C2(n2855), .A(n2854), .B(n2853), .ZN(U3290)
         );
  NAND2_X1 U3716 ( .A1(n2857), .A2(n2903), .ZN(n2859) );
  NAND2_X4 U3717 ( .A1(n2858), .A2(n2908), .ZN(n3707) );
  INV_X1 U3718 ( .A(n3707), .ZN(n3698) );
  INV_X1 U3719 ( .A(n2858), .ZN(n2965) );
  NAND2_X1 U3720 ( .A1(n2965), .A2(REG1_REG_0__SCAN_IN), .ZN(n2860) );
  INV_X1 U3721 ( .A(n3707), .ZN(n2861) );
  NAND2_X4 U3722 ( .A1(n2861), .A2(n3098), .ZN(n2964) );
  INV_X1 U3723 ( .A(n2964), .ZN(n2862) );
  NAND2_X1 U3724 ( .A1(n2862), .A2(n2857), .ZN(n2864) );
  AOI22_X1 U3725 ( .A1(n3697), .A2(n2948), .B1(n2965), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2863) );
  NAND2_X1 U3726 ( .A1(n2864), .A2(n2863), .ZN(n2865) );
  NAND2_X1 U3727 ( .A1(n2866), .A2(n2865), .ZN(n2916) );
  OAI21_X1 U3728 ( .B1(n2866), .B2(n2865), .A(n2916), .ZN(n2899) );
  NAND2_X1 U3729 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3882) );
  AOI21_X1 U3730 ( .B1(n2868), .B2(n3882), .A(n2897), .ZN(n2867) );
  OAI21_X1 U3731 ( .B1(n2899), .B2(n2868), .A(n2867), .ZN(n2869) );
  CLKBUF_X2 U3732 ( .A(U4043), .Z(n3872) );
  OAI211_X1 U3733 ( .C1(IR_REG_0__SCAN_IN), .C2(n2870), .A(n2869), .B(n3872), 
        .ZN(n3905) );
  XNOR2_X1 U3734 ( .A(n2871), .B(REG2_REG_4__SCAN_IN), .ZN(n2878) );
  OAI211_X1 U3735 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2873), .A(n4462), .B(n2872), 
        .ZN(n2875) );
  AND2_X1 U3736 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3044) );
  AOI21_X1 U3737 ( .B1(n4460), .B2(ADDR_REG_4__SCAN_IN), .A(n3044), .ZN(n2874)
         );
  OAI211_X1 U3738 ( .C1(n4467), .C2(n2876), .A(n2875), .B(n2874), .ZN(n2877)
         );
  AOI21_X1 U3739 ( .B1(n4406), .B2(n2878), .A(n2877), .ZN(n2879) );
  NAND2_X1 U3740 ( .A1(n3905), .A2(n2879), .ZN(U3244) );
  OR2_X1 U3741 ( .A1(n2881), .A2(n2880), .ZN(n2883) );
  AND2_X1 U3742 ( .A1(n2883), .A2(n2882), .ZN(n2893) );
  OAI21_X1 U3743 ( .B1(n2893), .B2(n4282), .A(n2921), .ZN(n2888) );
  NAND2_X1 U3744 ( .A1(n2888), .A2(n2887), .ZN(n2966) );
  OR2_X1 U3745 ( .A1(n2909), .A2(n4480), .ZN(n2890) );
  NAND2_X1 U3746 ( .A1(n2921), .A2(n3579), .ZN(n2967) );
  INV_X1 U3747 ( .A(n2967), .ZN(n2891) );
  NOR3_X1 U3748 ( .A1(n2966), .A2(n2891), .A3(n2895), .ZN(n2933) );
  NOR3_X1 U3749 ( .A1(n2921), .A2(n2895), .A3(n4066), .ZN(n2892) );
  INV_X1 U3750 ( .A(n2893), .ZN(n2894) );
  OR2_X1 U3751 ( .A1(n2895), .A2(n2894), .ZN(n2896) );
  NAND2_X1 U3752 ( .A1(n3579), .A2(n2897), .ZN(n2898) );
  OAI22_X1 U3753 ( .A1(n2899), .A2(n3845), .B1(n3840), .B2(n2912), .ZN(n2900)
         );
  AOI21_X1 U3754 ( .B1(n3782), .B2(n2948), .A(n2900), .ZN(n2901) );
  OAI21_X1 U3755 ( .B1(n2933), .B2(n2902), .A(n2901), .ZN(U3229) );
  INV_X1 U3756 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3025) );
  NAND2_X1 U3757 ( .A1(n2904), .A2(n2903), .ZN(n2907) );
  NAND2_X1 U3758 ( .A1(n2907), .A2(n2906), .ZN(n2910) );
  NAND2_X1 U3759 ( .A1(n2909), .A2(n2908), .ZN(n3401) );
  XNOR2_X1 U3760 ( .A(n2910), .B(n3401), .ZN(n2928) );
  NAND2_X1 U3761 ( .A1(n2903), .A2(n3029), .ZN(n2911) );
  OAI21_X1 U3762 ( .B1(n2964), .B2(n2912), .A(n2911), .ZN(n2913) );
  INV_X1 U3763 ( .A(n2913), .ZN(n2929) );
  XNOR2_X1 U3764 ( .A(n2928), .B(n2929), .ZN(n2917) );
  NAND2_X1 U3765 ( .A1(n2916), .A2(n2915), .ZN(n2918) );
  NAND2_X1 U3766 ( .A1(n2917), .A2(n2918), .ZN(n2931) );
  OAI211_X1 U3767 ( .C1(n2917), .C2(n2918), .A(n2931), .B(n3849), .ZN(n2924)
         );
  NAND2_X1 U3768 ( .A1(n3579), .A2(n2919), .ZN(n2920) );
  OAI22_X1 U3769 ( .A1(n2943), .A2(n3851), .B1(n3840), .B2(n2925), .ZN(n2922)
         );
  AOI21_X1 U3770 ( .B1(n3782), .B2(n3029), .A(n2922), .ZN(n2923) );
  OAI211_X1 U3771 ( .C1(n2933), .C2(n3025), .A(n2924), .B(n2923), .ZN(U3219)
         );
  OAI22_X1 U3772 ( .A1(n2925), .A2(n2964), .B1(n3708), .B2(n2927), .ZN(n2956)
         );
  XNOR2_X1 U3773 ( .A(n2957), .B(n2956), .ZN(n2932) );
  OAI22_X1 U3774 ( .A1(n3041), .A2(n3840), .B1(n3851), .B2(n2912), .ZN(n2935)
         );
  NOR2_X1 U3775 ( .A1(n2933), .A2(n3888), .ZN(n2934) );
  AOI211_X1 U3776 ( .C1(n2984), .C2(n3782), .A(n2935), .B(n2934), .ZN(n2936)
         );
  OAI21_X1 U3777 ( .B1(n2937), .B2(n3845), .A(n2936), .ZN(U3234) );
  OR2_X1 U3778 ( .A1(n2938), .A2(n2650), .ZN(n2939) );
  NAND2_X1 U3779 ( .A1(n2940), .A2(n2939), .ZN(n2945) );
  INV_X1 U3780 ( .A(n2945), .ZN(n3023) );
  AOI22_X1 U3781 ( .A1(n2941), .A2(n4284), .B1(n4282), .B2(n3029), .ZN(n2942)
         );
  OAI21_X1 U3782 ( .B1(n2943), .B2(n4288), .A(n2942), .ZN(n2947) );
  AOI21_X1 U3783 ( .B1(n2650), .B2(n3514), .A(n2944), .ZN(n2946) );
  OAI22_X1 U3784 ( .A1(n2946), .A2(n4070), .B1(n4111), .B2(n2945), .ZN(n3026)
         );
  AOI211_X1 U3785 ( .C1(n4502), .C2(n3023), .A(n2947), .B(n3026), .ZN(n2955)
         );
  NAND2_X1 U3786 ( .A1(n3029), .A2(n2948), .ZN(n2949) );
  NAND2_X1 U3787 ( .A1(n2950), .A2(n2949), .ZN(n3032) );
  OAI22_X1 U3788 ( .A1(n4294), .A2(n3032), .B1(n4517), .B2(n2348), .ZN(n2951)
         );
  INV_X1 U3789 ( .A(n2951), .ZN(n2952) );
  OAI21_X1 U3790 ( .B1(n2955), .B2(n4515), .A(n2952), .ZN(U3519) );
  OAI22_X1 U3791 ( .A1(n4347), .A2(n3032), .B1(n4512), .B2(n2346), .ZN(n2953)
         );
  INV_X1 U3792 ( .A(n2953), .ZN(n2954) );
  OAI21_X1 U3793 ( .B1(n2955), .B2(n4510), .A(n2954), .ZN(U3469) );
  INV_X1 U3794 ( .A(n2956), .ZN(n2960) );
  INV_X1 U3795 ( .A(n2957), .ZN(n2959) );
  NAND2_X1 U3796 ( .A1(n3876), .A2(n3697), .ZN(n2962) );
  NAND2_X1 U3797 ( .A1(n3698), .A2(n2980), .ZN(n2961) );
  NAND2_X1 U3798 ( .A1(n2962), .A2(n2961), .ZN(n2963) );
  XNOR2_X1 U3799 ( .A(n2963), .B(n3401), .ZN(n3035) );
  OAI22_X1 U3800 ( .A1(n3041), .A2(n2964), .B1(n3708), .B2(n3011), .ZN(n3034)
         );
  XNOR2_X1 U3801 ( .A(n3035), .B(n3034), .ZN(n3036) );
  XOR2_X1 U3802 ( .A(n3037), .B(n3036), .Z(n2973) );
  OAI22_X1 U3803 ( .A1(n2925), .A2(n3851), .B1(n3840), .B2(n3120), .ZN(n2971)
         );
  OAI21_X1 U3804 ( .B1(n2966), .B2(n2965), .A(STATE_REG_SCAN_IN), .ZN(n2968)
         );
  MUX2_X1 U3805 ( .A(U3149), .B(n3843), .S(n2969), .Z(n2970) );
  AOI211_X1 U3806 ( .C1(n2980), .C2(n3782), .A(n2971), .B(n2970), .ZN(n2972)
         );
  OAI21_X1 U3807 ( .B1(n2973), .B2(n3845), .A(n2972), .ZN(U3215) );
  OR2_X1 U3808 ( .A1(n2974), .A2(n3011), .ZN(n2975) );
  NAND2_X1 U3809 ( .A1(n2975), .A2(n3002), .ZN(n3019) );
  XNOR2_X1 U3810 ( .A(n2976), .B(n3483), .ZN(n3017) );
  OAI21_X1 U3811 ( .B1(n3483), .B2(n2978), .A(n2977), .ZN(n2979) );
  AOI22_X1 U3812 ( .A1(n2979), .A2(n4169), .B1(n4240), .B2(n2941), .ZN(n3012)
         );
  AOI22_X1 U3813 ( .A1(n3875), .A2(n4284), .B1(n4282), .B2(n2980), .ZN(n2981)
         );
  OAI211_X1 U3814 ( .C1(n4280), .C2(n3017), .A(n3012), .B(n2981), .ZN(n3021)
         );
  NAND2_X1 U3815 ( .A1(n3021), .A2(n4512), .ZN(n2983) );
  NAND2_X1 U3816 ( .A1(n4510), .A2(REG0_REG_3__SCAN_IN), .ZN(n2982) );
  OAI211_X1 U3817 ( .C1(n3019), .C2(n4347), .A(n2983), .B(n2982), .ZN(U3473)
         );
  AOI22_X1 U3818 ( .A1(n3876), .A2(n4284), .B1(n2984), .B2(n4282), .ZN(n2985)
         );
  OAI21_X1 U3819 ( .B1(n2912), .B2(n4288), .A(n2985), .ZN(n2987) );
  AOI211_X1 U3820 ( .C1(n4502), .C2(n2988), .A(n2987), .B(n2986), .ZN(n2992)
         );
  AOI22_X1 U3821 ( .A1(n2738), .A2(n2990), .B1(REG0_REG_2__SCAN_IN), .B2(n4510), .ZN(n2989) );
  OAI21_X1 U3822 ( .B1(n2992), .B2(n4510), .A(n2989), .ZN(U3471) );
  AOI22_X1 U3823 ( .A1(n2734), .A2(n2990), .B1(REG1_REG_2__SCAN_IN), .B2(n4515), .ZN(n2991) );
  OAI21_X1 U3824 ( .B1(n2992), .B2(n4515), .A(n2991), .ZN(U3520) );
  NAND2_X1 U3825 ( .A1(n2994), .A2(n3482), .ZN(n2995) );
  AND2_X1 U3826 ( .A1(n2993), .A2(n2995), .ZN(n4503) );
  INV_X1 U3827 ( .A(n4503), .ZN(n3006) );
  INV_X1 U3828 ( .A(n4474), .ZN(n3242) );
  XOR2_X1 U3829 ( .A(n3482), .B(n2996), .Z(n3001) );
  AOI22_X1 U3830 ( .A1(n3876), .A2(n4240), .B1(n2997), .B2(n4282), .ZN(n2998)
         );
  OAI21_X1 U3831 ( .B1(n3133), .B2(n4273), .A(n2998), .ZN(n2999) );
  AOI21_X1 U3832 ( .B1(n4503), .B2(n3211), .A(n2999), .ZN(n3000) );
  OAI21_X1 U3833 ( .B1(n3001), .B2(n4070), .A(n3000), .ZN(n4500) );
  OAI211_X1 U3834 ( .C1(n2134), .C2(n3042), .A(n4276), .B(n3054), .ZN(n4499)
         );
  OAI22_X1 U3835 ( .A1(n4499), .A2(n4352), .B1(n4468), .B2(n3047), .ZN(n3003)
         );
  OAI21_X1 U3836 ( .B1(n4500), .B2(n3003), .A(n4164), .ZN(n3005) );
  NAND2_X1 U3837 ( .A1(n4118), .A2(REG2_REG_4__SCAN_IN), .ZN(n3004) );
  OAI211_X1 U3838 ( .C1(n3006), .C2(n3242), .A(n3005), .B(n3004), .ZN(U3286)
         );
  NAND2_X1 U3839 ( .A1(n4111), .A2(n3007), .ZN(n3008) );
  INV_X1 U3840 ( .A(n3019), .ZN(n3015) );
  OAI22_X1 U3841 ( .A1(n4164), .A2(n3909), .B1(REG3_REG_3__SCAN_IN), .B2(n4468), .ZN(n3009) );
  AOI21_X1 U3842 ( .B1(n4178), .B2(n3875), .A(n3009), .ZN(n3010) );
  OAI21_X1 U3843 ( .B1(n3011), .B2(n4185), .A(n3010), .ZN(n3014) );
  NOR2_X1 U3844 ( .A1(n3012), .A2(n4360), .ZN(n3013) );
  AOI211_X1 U3845 ( .C1(n3015), .C2(n4473), .A(n3014), .B(n3013), .ZN(n3016)
         );
  OAI21_X1 U3846 ( .B1(n4167), .B2(n3017), .A(n3016), .ZN(U3287) );
  OAI22_X1 U3847 ( .A1(n4294), .A2(n3019), .B1(n4517), .B2(n3018), .ZN(n3020)
         );
  AOI21_X1 U3848 ( .B1(n3021), .B2(n4517), .A(n3020), .ZN(n3022) );
  INV_X1 U3849 ( .A(n3022), .ZN(U3521) );
  NAND2_X1 U3850 ( .A1(n4474), .A2(n3023), .ZN(n3024) );
  OAI21_X1 U3851 ( .B1(n4468), .B2(n3025), .A(n3024), .ZN(n3028) );
  MUX2_X1 U3852 ( .A(REG2_REG_1__SCAN_IN), .B(n3026), .S(n4164), .Z(n3027) );
  AOI211_X1 U3853 ( .C1(n4179), .C2(n2857), .A(n3028), .B(n3027), .ZN(n3031)
         );
  AOI22_X1 U3854 ( .A1(n3327), .A2(n3029), .B1(n4178), .B2(n2941), .ZN(n3030)
         );
  OAI211_X1 U3855 ( .C1(n4139), .C2(n3032), .A(n3031), .B(n3030), .ZN(U3289)
         );
  INV_X1 U3856 ( .A(n3843), .ZN(n3858) );
  OAI22_X1 U3857 ( .A1(n3120), .A2(n3708), .B1(n3707), .B2(n3042), .ZN(n3033)
         );
  XNOR2_X1 U3858 ( .A(n3033), .B(n3709), .ZN(n3110) );
  OAI22_X1 U3859 ( .A1(n3120), .A2(n2964), .B1(n3702), .B2(n3042), .ZN(n3109)
         );
  XNOR2_X1 U3860 ( .A(n3110), .B(n3109), .ZN(n3039) );
  OAI22_X1 U3861 ( .A1(n3037), .A2(n3036), .B1(n3035), .B2(n3034), .ZN(n3038)
         );
  AOI211_X1 U3862 ( .C1(n3039), .C2(n3038), .A(n3845), .B(n3112), .ZN(n3040)
         );
  INV_X1 U3863 ( .A(n3040), .ZN(n3046) );
  INV_X1 U3864 ( .A(n3840), .ZN(n3854) );
  OAI22_X1 U3865 ( .A1(n2045), .A2(n3042), .B1(n3041), .B2(n3851), .ZN(n3043)
         );
  AOI211_X1 U3866 ( .C1(n3854), .C2(n3874), .A(n3044), .B(n3043), .ZN(n3045)
         );
  OAI211_X1 U3867 ( .C1(n3858), .C2(n3047), .A(n3046), .B(n3045), .ZN(U3227)
         );
  INV_X1 U3868 ( .A(n3048), .ZN(n3529) );
  NAND2_X1 U3869 ( .A1(n3529), .A2(n3503), .ZN(n3476) );
  XOR2_X1 U3870 ( .A(n3049), .B(n3476), .Z(n3079) );
  XNOR2_X1 U3871 ( .A(n3050), .B(n3476), .ZN(n3051) );
  NAND2_X1 U3872 ( .A1(n3051), .A2(n4169), .ZN(n3081) );
  AOI22_X1 U3873 ( .A1(n3873), .A2(n4284), .B1(n4282), .B2(n3114), .ZN(n3052)
         );
  OAI211_X1 U3874 ( .C1(n3120), .C2(n4288), .A(n3081), .B(n3052), .ZN(n3053)
         );
  AOI21_X1 U3875 ( .B1(n3079), .B2(n4504), .A(n3053), .ZN(n3059) );
  AND2_X1 U3876 ( .A1(n3054), .A2(n3114), .ZN(n3055) );
  NOR2_X1 U3877 ( .A1(n3065), .A2(n3055), .ZN(n3073) );
  AOI22_X1 U3878 ( .A1(n2738), .A2(n3073), .B1(REG0_REG_5__SCAN_IN), .B2(n4510), .ZN(n3056) );
  OAI21_X1 U3879 ( .B1(n3059), .B2(n4510), .A(n3056), .ZN(U3477) );
  NAND2_X1 U3880 ( .A1(n4515), .A2(REG1_REG_5__SCAN_IN), .ZN(n3058) );
  NAND2_X1 U3881 ( .A1(n2734), .A2(n3073), .ZN(n3057) );
  OAI211_X1 U3882 ( .C1(n3059), .C2(n4515), .A(n3058), .B(n3057), .ZN(U3523)
         );
  NAND2_X1 U3883 ( .A1(n3532), .A2(n3528), .ZN(n3485) );
  XNOR2_X1 U3884 ( .A(n3060), .B(n3485), .ZN(n3083) );
  XOR2_X1 U3885 ( .A(n3485), .B(n3061), .Z(n3082) );
  AOI22_X1 U3886 ( .A1(n3871), .A2(n4284), .B1(n3084), .B2(n4282), .ZN(n3062)
         );
  OAI21_X1 U3887 ( .B1(n3133), .B2(n4288), .A(n3062), .ZN(n3063) );
  AOI21_X1 U3888 ( .B1(n3082), .B2(n4169), .A(n3063), .ZN(n3064) );
  OAI21_X1 U3889 ( .B1(n4280), .B2(n3083), .A(n3064), .ZN(n3071) );
  OR2_X1 U3890 ( .A1(n3065), .A2(n3134), .ZN(n3066) );
  NAND2_X1 U3891 ( .A1(n3100), .A2(n3066), .ZN(n3089) );
  OAI22_X1 U3892 ( .A1(n4294), .A2(n3089), .B1(n4517), .B2(n2416), .ZN(n3067)
         );
  AOI21_X1 U3893 ( .B1(n3071), .B2(n4517), .A(n3067), .ZN(n3068) );
  INV_X1 U3894 ( .A(n3068), .ZN(U3524) );
  INV_X1 U3895 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3069) );
  OAI22_X1 U3896 ( .A1(n4347), .A2(n3089), .B1(n4512), .B2(n3069), .ZN(n3070)
         );
  AOI21_X1 U3897 ( .B1(n3071), .B2(n4512), .A(n3070), .ZN(n3072) );
  INV_X1 U3898 ( .A(n3072), .ZN(U3479) );
  INV_X1 U3899 ( .A(n3073), .ZN(n3077) );
  AOI22_X1 U3900 ( .A1(n4179), .A2(n3875), .B1(n4178), .B2(n3873), .ZN(n3076)
         );
  OAI22_X1 U3901 ( .A1(n4164), .A2(n2399), .B1(n3126), .B2(n4468), .ZN(n3074)
         );
  AOI21_X1 U3902 ( .B1(n3114), .B2(n3327), .A(n3074), .ZN(n3075) );
  OAI211_X1 U3903 ( .C1(n4139), .C2(n3077), .A(n3076), .B(n3075), .ZN(n3078)
         );
  AOI21_X1 U3904 ( .B1(n3079), .B2(n4173), .A(n3078), .ZN(n3080) );
  OAI21_X1 U3905 ( .B1(n4118), .B2(n3081), .A(n3080), .ZN(U3285) );
  INV_X1 U3906 ( .A(n3082), .ZN(n3093) );
  NAND2_X1 U3907 ( .A1(n4164), .A2(n4169), .ZN(n3336) );
  INV_X1 U3908 ( .A(n3083), .ZN(n3091) );
  AOI22_X1 U3909 ( .A1(n3327), .A2(n3084), .B1(n4178), .B2(n3871), .ZN(n3088)
         );
  OAI22_X1 U3910 ( .A1(n4164), .A2(n3085), .B1(n3139), .B2(n4468), .ZN(n3086)
         );
  AOI21_X1 U3911 ( .B1(n4179), .B2(n3874), .A(n3086), .ZN(n3087) );
  OAI211_X1 U3912 ( .C1(n4139), .C2(n3089), .A(n3088), .B(n3087), .ZN(n3090)
         );
  AOI21_X1 U3913 ( .B1(n3091), .B2(n4173), .A(n3090), .ZN(n3092) );
  OAI21_X1 U3914 ( .B1(n3093), .B2(n3336), .A(n3092), .ZN(U3284) );
  XNOR2_X1 U3915 ( .A(n3094), .B(n3533), .ZN(n3097) );
  AOI22_X1 U3916 ( .A1(n3870), .A2(n4284), .B1(n4282), .B2(n3099), .ZN(n3095)
         );
  OAI21_X1 U3917 ( .B1(n3176), .B2(n4288), .A(n3095), .ZN(n3096) );
  AOI21_X1 U3918 ( .B1(n3097), .B2(n4169), .A(n3096), .ZN(n4509) );
  AOI21_X1 U3919 ( .B1(n3100), .B2(n3099), .A(n3098), .ZN(n3101) );
  NAND2_X1 U3920 ( .A1(n3101), .A2(n3214), .ZN(n4508) );
  INV_X1 U3921 ( .A(n4508), .ZN(n3105) );
  INV_X1 U3922 ( .A(n4160), .ZN(n3104) );
  OAI22_X1 U3923 ( .A1(n4164), .A2(n3102), .B1(n3182), .B2(n4468), .ZN(n3103)
         );
  AOI21_X1 U3924 ( .B1(n3105), .B2(n3104), .A(n3103), .ZN(n3108) );
  OR2_X1 U3925 ( .A1(n3106), .A2(n3533), .ZN(n4506) );
  NAND2_X1 U3926 ( .A1(n3106), .A2(n3533), .ZN(n4505) );
  NAND3_X1 U3927 ( .A1(n4506), .A2(n4505), .A3(n4173), .ZN(n3107) );
  OAI211_X1 U3928 ( .C1(n4509), .C2(n4118), .A(n3108), .B(n3107), .ZN(U3283)
         );
  OAI22_X1 U3929 ( .A1(n3133), .A2(n3708), .B1(n3707), .B2(n3121), .ZN(n3113)
         );
  INV_X2 U3930 ( .A(n3173), .ZN(n3709) );
  XNOR2_X1 U3931 ( .A(n3113), .B(n3709), .ZN(n3128) );
  OR2_X1 U3932 ( .A1(n3133), .A2(n2964), .ZN(n3116) );
  NAND2_X1 U3933 ( .A1(n3677), .A2(n3114), .ZN(n3115) );
  NAND2_X1 U3934 ( .A1(n3116), .A2(n3115), .ZN(n3127) );
  XNOR2_X1 U3935 ( .A(n3128), .B(n3127), .ZN(n3117) );
  AOI211_X1 U3936 ( .C1(n3118), .C2(n3117), .A(n3845), .B(n3129), .ZN(n3119)
         );
  INV_X1 U3937 ( .A(n3119), .ZN(n3125) );
  OAI22_X1 U3938 ( .A1(n2045), .A2(n3121), .B1(n3120), .B2(n3851), .ZN(n3122)
         );
  AOI211_X1 U3939 ( .C1(n3854), .C2(n3873), .A(n3123), .B(n3122), .ZN(n3124)
         );
  OAI211_X1 U3940 ( .C1(n3858), .C2(n3126), .A(n3125), .B(n3124), .ZN(U3224)
         );
  OAI22_X1 U3941 ( .A1(n3176), .A2(n3708), .B1(n3707), .B2(n3134), .ZN(n3130)
         );
  XNOR2_X1 U3942 ( .A(n3130), .B(n3709), .ZN(n3169) );
  INV_X1 U3943 ( .A(n3168), .ZN(n3170) );
  XNOR2_X1 U3944 ( .A(n3169), .B(n3170), .ZN(n3131) );
  XNOR2_X1 U3945 ( .A(n3171), .B(n3131), .ZN(n3132) );
  NAND2_X1 U3946 ( .A1(n3132), .A2(n3849), .ZN(n3138) );
  OAI22_X1 U3947 ( .A1(n2045), .A2(n3134), .B1(n3133), .B2(n3851), .ZN(n3135)
         );
  AOI211_X1 U3948 ( .C1(n3854), .C2(n3871), .A(n3136), .B(n3135), .ZN(n3137)
         );
  OAI211_X1 U3949 ( .C1(n3858), .C2(n3139), .A(n3138), .B(n3137), .ZN(U3236)
         );
  INV_X1 U3950 ( .A(n3140), .ZN(n3511) );
  AND2_X1 U3951 ( .A1(n3511), .A2(n3539), .ZN(n3491) );
  XOR2_X1 U3952 ( .A(n3491), .B(n3141), .Z(n3142) );
  NAND2_X1 U3953 ( .A1(n3142), .A2(n4169), .ZN(n3161) );
  INV_X1 U3954 ( .A(n3213), .ZN(n3143) );
  AOI21_X1 U3955 ( .B1(n3247), .B2(n3143), .A(n3152), .ZN(n3165) );
  INV_X1 U3956 ( .A(n4179), .ZN(n3331) );
  AOI22_X1 U3957 ( .A1(n3327), .A2(n3247), .B1(n4178), .B2(n3868), .ZN(n3144)
         );
  OAI21_X1 U3958 ( .B1(n3252), .B2(n3331), .A(n3144), .ZN(n3146) );
  OAI22_X1 U3959 ( .A1(n3257), .A2(n4468), .B1(n2457), .B2(n4164), .ZN(n3145)
         );
  AOI211_X1 U3960 ( .C1(n3165), .C2(n4473), .A(n3146), .B(n3145), .ZN(n3149)
         );
  XNOR2_X1 U3961 ( .A(n3147), .B(n3491), .ZN(n3163) );
  NAND2_X1 U3962 ( .A1(n3163), .A2(n4173), .ZN(n3148) );
  OAI211_X1 U3963 ( .C1(n3161), .C2(n4118), .A(n3149), .B(n3148), .ZN(U3281)
         );
  NAND2_X1 U3964 ( .A1(n3507), .A2(n3502), .ZN(n3474) );
  XNOR2_X1 U3965 ( .A(n3150), .B(n3474), .ZN(n3224) );
  XNOR2_X1 U3966 ( .A(n3151), .B(n3474), .ZN(n3226) );
  NAND2_X1 U3967 ( .A1(n3226), .A2(n4173), .ZN(n3159) );
  INV_X1 U3968 ( .A(n3152), .ZN(n3153) );
  AOI21_X1 U3969 ( .B1(n3266), .B2(n3153), .A(n2083), .ZN(n3228) );
  AOI22_X1 U3970 ( .A1(n3327), .A2(n3266), .B1(n4178), .B2(n3867), .ZN(n3156)
         );
  INV_X1 U3971 ( .A(n3280), .ZN(n3154) );
  AOI22_X1 U3972 ( .A1(n4118), .A2(REG2_REG_10__SCAN_IN), .B1(n3154), .B2(
        n4181), .ZN(n3155) );
  OAI211_X1 U3973 ( .C1(n3274), .C2(n3331), .A(n3156), .B(n3155), .ZN(n3157)
         );
  AOI21_X1 U3974 ( .B1(n3228), .B2(n4473), .A(n3157), .ZN(n3158) );
  OAI211_X1 U3975 ( .C1(n3224), .C2(n3336), .A(n3159), .B(n3158), .ZN(U3280)
         );
  AOI22_X1 U3976 ( .A1(n3868), .A2(n4284), .B1(n4282), .B2(n3247), .ZN(n3160)
         );
  OAI211_X1 U3977 ( .C1(n3252), .C2(n4288), .A(n3161), .B(n3160), .ZN(n3162)
         );
  AOI21_X1 U3978 ( .B1(n3163), .B2(n4504), .A(n3162), .ZN(n3167) );
  AOI22_X1 U3979 ( .A1(n3165), .A2(n2734), .B1(REG1_REG_9__SCAN_IN), .B2(n4515), .ZN(n3164) );
  OAI21_X1 U3980 ( .B1(n3167), .B2(n4515), .A(n3164), .ZN(U3527) );
  AOI22_X1 U3981 ( .A1(n3165), .A2(n2738), .B1(REG0_REG_9__SCAN_IN), .B2(n4510), .ZN(n3166) );
  OAI21_X1 U3982 ( .B1(n3167), .B2(n4510), .A(n3166), .ZN(U3485) );
  OAI22_X1 U3983 ( .A1(n3206), .A2(n3708), .B1(n3707), .B2(n3177), .ZN(n3174)
         );
  XNOR2_X1 U3984 ( .A(n3174), .B(n3173), .ZN(n3183) );
  OAI22_X1 U3985 ( .A1(n3206), .A2(n2964), .B1(n3702), .B2(n3177), .ZN(n3184)
         );
  XNOR2_X1 U3986 ( .A(n3183), .B(n3184), .ZN(n3186) );
  XOR2_X1 U3987 ( .A(n3187), .B(n3186), .Z(n3175) );
  NAND2_X1 U3988 ( .A1(n3175), .A2(n3849), .ZN(n3181) );
  OAI22_X1 U3989 ( .A1(n2045), .A2(n3177), .B1(n3176), .B2(n3851), .ZN(n3178)
         );
  AOI211_X1 U3990 ( .C1(n3854), .C2(n3870), .A(n3179), .B(n3178), .ZN(n3180)
         );
  OAI211_X1 U3991 ( .C1(n3858), .C2(n3182), .A(n3181), .B(n3180), .ZN(U3210)
         );
  INV_X1 U3992 ( .A(n3183), .ZN(n3185) );
  OAI22_X1 U3993 ( .A1(n3252), .A2(n3702), .B1(n3707), .B2(n3205), .ZN(n3188)
         );
  XNOR2_X1 U3994 ( .A(n3188), .B(n3709), .ZN(n3191) );
  OR2_X1 U3995 ( .A1(n3252), .A2(n2964), .ZN(n3190) );
  NAND2_X1 U3996 ( .A1(n3677), .A2(n3215), .ZN(n3189) );
  NAND2_X1 U3997 ( .A1(n3190), .A2(n3189), .ZN(n3192) );
  NAND2_X1 U3998 ( .A1(n3191), .A2(n3192), .ZN(n3243) );
  INV_X1 U3999 ( .A(n3191), .ZN(n3194) );
  INV_X1 U4000 ( .A(n3192), .ZN(n3193) );
  NAND2_X1 U4001 ( .A1(n3194), .A2(n3193), .ZN(n3245) );
  NAND2_X1 U4002 ( .A1(n3243), .A2(n3245), .ZN(n3195) );
  XNOR2_X1 U4003 ( .A(n3244), .B(n3195), .ZN(n3201) );
  INV_X1 U4004 ( .A(n4469), .ZN(n3199) );
  INV_X1 U4005 ( .A(n3851), .ZN(n3781) );
  AOI22_X1 U4006 ( .A1(n3782), .A2(n3215), .B1(n3781), .B2(n3871), .ZN(n3197)
         );
  OAI211_X1 U4007 ( .C1(n3274), .C2(n3840), .A(n3197), .B(n3196), .ZN(n3198)
         );
  AOI21_X1 U4008 ( .B1(n3199), .B2(n3843), .A(n3198), .ZN(n3200) );
  OAI21_X1 U4009 ( .B1(n3201), .B2(n3845), .A(n3200), .ZN(U3218) );
  NAND2_X1 U4010 ( .A1(n3538), .A2(n3535), .ZN(n3486) );
  NAND2_X1 U4011 ( .A1(n4506), .A2(n3202), .ZN(n3203) );
  XOR2_X1 U4012 ( .A(n3486), .B(n3203), .Z(n4475) );
  INV_X1 U4013 ( .A(n4475), .ZN(n3212) );
  XOR2_X1 U4014 ( .A(n3486), .B(n3204), .Z(n3209) );
  OAI22_X1 U4015 ( .A1(n3206), .A2(n4288), .B1(n3205), .B2(n4066), .ZN(n3207)
         );
  AOI21_X1 U4016 ( .B1(n4284), .B2(n3869), .A(n3207), .ZN(n3208) );
  OAI21_X1 U4017 ( .B1(n3209), .B2(n4070), .A(n3208), .ZN(n3210) );
  AOI21_X1 U4018 ( .B1(n3211), .B2(n4475), .A(n3210), .ZN(n4478) );
  OAI21_X1 U4019 ( .B1(n3281), .B2(n3212), .A(n4478), .ZN(n3218) );
  NAND2_X1 U4020 ( .A1(n3218), .A2(n4517), .ZN(n3217) );
  AOI21_X1 U4021 ( .B1(n3215), .B2(n3214), .A(n3213), .ZN(n4472) );
  NAND2_X1 U4022 ( .A1(n4472), .A2(n2734), .ZN(n3216) );
  OAI211_X1 U4023 ( .C1(n4517), .C2(n3939), .A(n3217), .B(n3216), .ZN(U3526)
         );
  INV_X1 U4024 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4025 ( .A1(n3218), .A2(n4512), .ZN(n3220) );
  NAND2_X1 U4026 ( .A1(n4472), .A2(n2738), .ZN(n3219) );
  OAI211_X1 U4027 ( .C1(n4512), .C2(n3221), .A(n3220), .B(n3219), .ZN(U3483)
         );
  OAI22_X1 U4028 ( .A1(n3356), .A2(n4273), .B1(n4066), .B2(n3275), .ZN(n3222)
         );
  AOI21_X1 U4029 ( .B1(n4240), .B2(n3869), .A(n3222), .ZN(n3223) );
  OAI21_X1 U4030 ( .B1(n3224), .B2(n4070), .A(n3223), .ZN(n3225) );
  AOI21_X1 U4031 ( .B1(n4504), .B2(n3226), .A(n3225), .ZN(n3230) );
  AOI22_X1 U4032 ( .A1(n3228), .A2(n2734), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4515), .ZN(n3227) );
  OAI21_X1 U4033 ( .B1(n3230), .B2(n4515), .A(n3227), .ZN(U3528) );
  AOI22_X1 U4034 ( .A1(n3228), .A2(n2738), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4510), .ZN(n3229) );
  OAI21_X1 U4035 ( .B1(n3230), .B2(n4510), .A(n3229), .ZN(U3487) );
  AOI21_X1 U4036 ( .B1(n3490), .B2(n3231), .A(n2275), .ZN(n3282) );
  AOI22_X1 U4037 ( .A1(n3866), .A2(n4284), .B1(n4282), .B2(n3233), .ZN(n3236)
         );
  XNOR2_X1 U4038 ( .A(n3294), .B(n3490), .ZN(n3234) );
  NAND2_X1 U4039 ( .A1(n3234), .A2(n4169), .ZN(n3235) );
  OAI211_X1 U4040 ( .C1(n3282), .C2(n4111), .A(n3236), .B(n3235), .ZN(n3284)
         );
  NAND2_X1 U4041 ( .A1(n3284), .A2(n4164), .ZN(n3241) );
  OAI22_X1 U4042 ( .A1(n4164), .A2(n3237), .B1(n3364), .B2(n4468), .ZN(n3239)
         );
  OAI21_X1 U40430 ( .B1(n2083), .B2(n3360), .A(n3311), .ZN(n3290) );
  NOR2_X1 U4044 ( .A1(n3290), .A2(n4139), .ZN(n3238) );
  AOI211_X1 U4045 ( .C1(n4179), .C2(n3868), .A(n3239), .B(n3238), .ZN(n3240)
         );
  OAI211_X1 U4046 ( .C1(n3282), .C2(n3242), .A(n3241), .B(n3240), .ZN(U3279)
         );
  OAI22_X1 U4047 ( .A1(n3274), .A2(n2964), .B1(n3702), .B2(n3253), .ZN(n3261)
         );
  NAND2_X1 U4048 ( .A1(n3869), .A2(n3677), .ZN(n3249) );
  NAND2_X1 U4049 ( .A1(n3698), .A2(n3247), .ZN(n3248) );
  NAND2_X1 U4050 ( .A1(n3249), .A2(n3248), .ZN(n3250) );
  XNOR2_X1 U4051 ( .A(n3250), .B(n3709), .ZN(n3260) );
  XNOR2_X1 U4052 ( .A(n3259), .B(n3258), .ZN(n3251) );
  NAND2_X1 U4053 ( .A1(n3251), .A2(n3849), .ZN(n3256) );
  NOR2_X1 U4054 ( .A1(STATE_REG_SCAN_IN), .A2(n2453), .ZN(n4373) );
  OAI22_X1 U4055 ( .A1(n2045), .A2(n3253), .B1(n3252), .B2(n3851), .ZN(n3254)
         );
  AOI211_X1 U4056 ( .C1(n3854), .C2(n3868), .A(n4373), .B(n3254), .ZN(n3255)
         );
  OAI211_X1 U4057 ( .C1(n3858), .C2(n3257), .A(n3256), .B(n3255), .ZN(U3228)
         );
  INV_X1 U4058 ( .A(n3260), .ZN(n3263) );
  NOR2_X1 U4059 ( .A1(n3702), .A2(n3275), .ZN(n3265) );
  AOI21_X1 U4060 ( .B1(n3704), .B2(n3868), .A(n3265), .ZN(n3350) );
  NAND2_X1 U4061 ( .A1(n3868), .A2(n3677), .ZN(n3268) );
  NAND2_X1 U4062 ( .A1(n3698), .A2(n3266), .ZN(n3267) );
  NAND2_X1 U4063 ( .A1(n3268), .A2(n3267), .ZN(n3269) );
  XNOR2_X1 U4064 ( .A(n3269), .B(n3709), .ZN(n3352) );
  XOR2_X1 U4065 ( .A(n3350), .B(n3352), .Z(n3271) );
  AOI21_X1 U4066 ( .B1(n3270), .B2(n3271), .A(n3845), .ZN(n3273) );
  INV_X1 U4067 ( .A(n3271), .ZN(n3272) );
  NAND2_X1 U4068 ( .A1(n3273), .A2(n3354), .ZN(n3279) );
  NAND2_X1 U4069 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4377) );
  INV_X1 U4070 ( .A(n4377), .ZN(n3277) );
  OAI22_X1 U4071 ( .A1(n2045), .A2(n3275), .B1(n3274), .B2(n3851), .ZN(n3276)
         );
  AOI211_X1 U4072 ( .C1(n3854), .C2(n3867), .A(n3277), .B(n3276), .ZN(n3278)
         );
  OAI211_X1 U4073 ( .C1(n3858), .C2(n3280), .A(n3279), .B(n3278), .ZN(U3214)
         );
  INV_X1 U4074 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3285) );
  OAI22_X1 U4075 ( .A1(n3282), .A2(n3281), .B1(n3359), .B2(n4288), .ZN(n3283)
         );
  NOR2_X1 U4076 ( .A1(n3284), .A2(n3283), .ZN(n3287) );
  MUX2_X1 U4077 ( .A(n3285), .B(n3287), .S(n4512), .Z(n3286) );
  OAI21_X1 U4078 ( .B1(n3290), .B2(n4347), .A(n3286), .ZN(U3489) );
  MUX2_X1 U4079 ( .A(n3288), .B(n3287), .S(n4517), .Z(n3289) );
  OAI21_X1 U4080 ( .B1(n4294), .B2(n3290), .A(n3289), .ZN(U3529) );
  INV_X1 U4081 ( .A(n3291), .ZN(n3292) );
  AOI21_X1 U4082 ( .B1(n3294), .B2(n3293), .A(n3292), .ZN(n3318) );
  INV_X1 U4083 ( .A(n3309), .ZN(n3295) );
  AOI21_X1 U4084 ( .B1(n3318), .B2(n3310), .A(n3295), .ZN(n3297) );
  XNOR2_X1 U4085 ( .A(n3602), .B(n3296), .ZN(n3464) );
  XNOR2_X1 U4086 ( .A(n3297), .B(n3464), .ZN(n3300) );
  OAI22_X1 U4087 ( .A1(n4289), .A2(n4273), .B1(n4066), .B2(n3606), .ZN(n3298)
         );
  AOI21_X1 U4088 ( .B1(n4240), .B2(n3866), .A(n3298), .ZN(n3299) );
  OAI21_X1 U4089 ( .B1(n3300), .B2(n4070), .A(n3299), .ZN(n3378) );
  INV_X1 U4090 ( .A(n3378), .ZN(n3307) );
  XNOR2_X1 U4091 ( .A(n3301), .B(n3464), .ZN(n3379) );
  NOR2_X1 U4092 ( .A1(n3312), .A2(n3606), .ZN(n3302) );
  OR2_X1 U4093 ( .A1(n3326), .A2(n3302), .ZN(n3385) );
  INV_X1 U4094 ( .A(n3610), .ZN(n3303) );
  AOI22_X1 U4095 ( .A1(n4118), .A2(REG2_REG_13__SCAN_IN), .B1(n3303), .B2(
        n4181), .ZN(n3304) );
  OAI21_X1 U4096 ( .B1(n3385), .B2(n4139), .A(n3304), .ZN(n3305) );
  AOI21_X1 U4097 ( .B1(n3379), .B2(n4173), .A(n3305), .ZN(n3306) );
  OAI21_X1 U4098 ( .B1(n3307), .B2(n4360), .A(n3306), .ZN(U3277) );
  NAND2_X1 U4099 ( .A1(n3310), .A2(n3309), .ZN(n3475) );
  XNOR2_X1 U4100 ( .A(n3308), .B(n3475), .ZN(n3337) );
  AND2_X1 U4101 ( .A1(n3311), .A2(n3411), .ZN(n3313) );
  OR2_X1 U4102 ( .A1(n3313), .A2(n3312), .ZN(n3349) );
  OAI22_X1 U4103 ( .A1(n4164), .A2(n3314), .B1(n3410), .B2(n4468), .ZN(n3315)
         );
  AOI21_X1 U4104 ( .B1(n3411), .B2(n3327), .A(n3315), .ZN(n3317) );
  AOI22_X1 U4105 ( .A1(n4179), .A2(n3867), .B1(n4178), .B2(n3865), .ZN(n3316)
         );
  OAI211_X1 U4106 ( .C1(n3349), .C2(n4139), .A(n3317), .B(n3316), .ZN(n3321)
         );
  XNOR2_X1 U4107 ( .A(n3318), .B(n3475), .ZN(n3319) );
  NAND2_X1 U4108 ( .A1(n3319), .A2(n4169), .ZN(n3341) );
  NOR2_X1 U4109 ( .A1(n3341), .A2(n4360), .ZN(n3320) );
  AOI211_X1 U4110 ( .C1(n4173), .C2(n3337), .A(n3321), .B(n3320), .ZN(n3322)
         );
  INV_X1 U4111 ( .A(n3322), .ZN(U3278) );
  XNOR2_X1 U4112 ( .A(n3440), .B(n3324), .ZN(n3388) );
  OAI21_X1 U4113 ( .B1(n3325), .B2(n3324), .A(n3323), .ZN(n3390) );
  NAND2_X1 U4114 ( .A1(n3390), .A2(n4173), .ZN(n3335) );
  OAI21_X1 U4115 ( .B1(n3326), .B2(n3617), .A(n3369), .ZN(n3396) );
  INV_X1 U4116 ( .A(n3396), .ZN(n3333) );
  AOI22_X1 U4117 ( .A1(n3327), .A2(n3747), .B1(n4178), .B2(n3863), .ZN(n3330)
         );
  INV_X1 U4118 ( .A(n3328), .ZN(n3752) );
  AOI22_X1 U4119 ( .A1(n4118), .A2(REG2_REG_14__SCAN_IN), .B1(n3752), .B2(
        n4181), .ZN(n3329) );
  OAI211_X1 U4120 ( .C1(n3602), .C2(n3331), .A(n3330), .B(n3329), .ZN(n3332)
         );
  AOI21_X1 U4121 ( .B1(n3333), .B2(n4473), .A(n3332), .ZN(n3334) );
  OAI211_X1 U4122 ( .C1(n3388), .C2(n3336), .A(n3335), .B(n3334), .ZN(U3276)
         );
  NAND2_X1 U4123 ( .A1(n3337), .A2(n4504), .ZN(n3343) );
  OR2_X1 U4124 ( .A1(n3356), .A2(n4288), .ZN(n3339) );
  NAND2_X1 U4125 ( .A1(n3411), .A2(n4282), .ZN(n3338) );
  OAI211_X1 U4126 ( .C1(n3602), .C2(n4273), .A(n3339), .B(n3338), .ZN(n3340)
         );
  INV_X1 U4127 ( .A(n3340), .ZN(n3342) );
  MUX2_X1 U4128 ( .A(n3344), .B(n3346), .S(n4517), .Z(n3345) );
  OAI21_X1 U4129 ( .B1(n4294), .B2(n3349), .A(n3345), .ZN(U3530) );
  INV_X1 U4130 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3347) );
  MUX2_X1 U4131 ( .A(n3347), .B(n3346), .S(n4512), .Z(n3348) );
  OAI21_X1 U4132 ( .B1(n3349), .B2(n4347), .A(n3348), .ZN(U3491) );
  INV_X1 U4133 ( .A(n3350), .ZN(n3351) );
  NAND2_X1 U4134 ( .A1(n3352), .A2(n3351), .ZN(n3353) );
  OAI22_X1 U4135 ( .A1(n3356), .A2(n3708), .B1(n3707), .B2(n3360), .ZN(n3355)
         );
  XNOR2_X1 U4136 ( .A(n3355), .B(n3709), .ZN(n3397) );
  OAI22_X1 U4137 ( .A1(n3356), .A2(n2964), .B1(n3702), .B2(n3360), .ZN(n3398)
         );
  XNOR2_X1 U4138 ( .A(n3397), .B(n3398), .ZN(n3357) );
  XNOR2_X1 U4139 ( .A(n3399), .B(n3357), .ZN(n3358) );
  NAND2_X1 U4140 ( .A1(n3358), .A2(n3849), .ZN(n3363) );
  AND2_X1 U4141 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4393) );
  OAI22_X1 U4142 ( .A1(n2045), .A2(n3360), .B1(n3359), .B2(n3851), .ZN(n3361)
         );
  AOI211_X1 U4143 ( .C1(n3854), .C2(n3866), .A(n4393), .B(n3361), .ZN(n3362)
         );
  OAI211_X1 U4144 ( .C1(n3858), .C2(n3364), .A(n3363), .B(n3362), .ZN(U3233)
         );
  AOI21_X1 U4145 ( .B1(n3365), .B2(n3493), .A(n4070), .ZN(n3367) );
  NAND2_X1 U4146 ( .A1(n3367), .A2(n3366), .ZN(n4287) );
  XNOR2_X1 U4147 ( .A(n3368), .B(n3493), .ZN(n4291) );
  NAND2_X1 U4148 ( .A1(n4291), .A2(n4173), .ZN(n3377) );
  INV_X1 U4149 ( .A(n3369), .ZN(n3370) );
  OAI21_X1 U4150 ( .B1(n3370), .B2(n3852), .A(n3588), .ZN(n4348) );
  INV_X1 U4151 ( .A(n4348), .ZN(n3375) );
  AOI22_X1 U4152 ( .A1(n4178), .A2(n4285), .B1(n4179), .B2(n3864), .ZN(n3373)
         );
  INV_X1 U4153 ( .A(n3857), .ZN(n3371) );
  AOI22_X1 U4154 ( .A1(n4118), .A2(REG2_REG_15__SCAN_IN), .B1(n3371), .B2(
        n4181), .ZN(n3372) );
  OAI211_X1 U4155 ( .C1(n3852), .C2(n4185), .A(n3373), .B(n3372), .ZN(n3374)
         );
  AOI21_X1 U4156 ( .B1(n3375), .B2(n4473), .A(n3374), .ZN(n3376) );
  OAI211_X1 U4157 ( .C1(n4118), .C2(n4287), .A(n3377), .B(n3376), .ZN(U3275)
         );
  AOI21_X1 U4158 ( .B1(n4504), .B2(n3379), .A(n3378), .ZN(n3382) );
  MUX2_X1 U4159 ( .A(n3380), .B(n3382), .S(n4517), .Z(n3381) );
  OAI21_X1 U4160 ( .B1(n4294), .B2(n3385), .A(n3381), .ZN(U3531) );
  INV_X1 U4161 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3383) );
  MUX2_X1 U4162 ( .A(n3383), .B(n3382), .S(n4512), .Z(n3384) );
  OAI21_X1 U4163 ( .B1(n3385), .B2(n4347), .A(n3384), .ZN(U3493) );
  INV_X1 U4164 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3391) );
  OAI22_X1 U4165 ( .A1(n4269), .A2(n4273), .B1(n4066), .B2(n3617), .ZN(n3386)
         );
  AOI21_X1 U4166 ( .B1(n4240), .B2(n3865), .A(n3386), .ZN(n3387) );
  OAI21_X1 U4167 ( .B1(n3388), .B2(n4070), .A(n3387), .ZN(n3389) );
  AOI21_X1 U4168 ( .B1(n3390), .B2(n4504), .A(n3389), .ZN(n3393) );
  MUX2_X1 U4169 ( .A(n3391), .B(n3393), .S(n4512), .Z(n3392) );
  OAI21_X1 U4170 ( .B1(n3396), .B2(n4347), .A(n3392), .ZN(U3495) );
  MUX2_X1 U4171 ( .A(n3394), .B(n3393), .S(n4517), .Z(n3395) );
  OAI21_X1 U4172 ( .B1(n4294), .B2(n3396), .A(n3395), .ZN(U3532) );
  OAI22_X1 U4173 ( .A1(n3605), .A2(n3702), .B1(n3707), .B2(n3400), .ZN(n3402)
         );
  XNOR2_X1 U4174 ( .A(n3402), .B(n3173), .ZN(n3406) );
  OR2_X1 U4175 ( .A1(n3605), .A2(n2964), .ZN(n3404) );
  NAND2_X1 U4176 ( .A1(n3677), .A2(n3411), .ZN(n3403) );
  NAND2_X1 U4177 ( .A1(n3404), .A2(n3403), .ZN(n3407) );
  INV_X1 U4178 ( .A(n3407), .ZN(n3405) );
  INV_X1 U4179 ( .A(n3406), .ZN(n3408) );
  NAND2_X1 U4180 ( .A1(n3408), .A2(n3407), .ZN(n3599) );
  NAND2_X1 U4181 ( .A1(n2084), .A2(n3599), .ZN(n3409) );
  XNOR2_X1 U4182 ( .A(n3600), .B(n3409), .ZN(n3416) );
  INV_X1 U4183 ( .A(n3410), .ZN(n3414) );
  AOI22_X1 U4184 ( .A1(n3782), .A2(n3411), .B1(n3781), .B2(n3867), .ZN(n3412)
         );
  NAND2_X1 U4185 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4397) );
  OAI211_X1 U4186 ( .C1(n3602), .C2(n3840), .A(n3412), .B(n4397), .ZN(n3413)
         );
  AOI21_X1 U4187 ( .B1(n3414), .B2(n3843), .A(n3413), .ZN(n3415) );
  OAI21_X1 U4188 ( .B1(n3416), .B2(n3845), .A(n3415), .ZN(U3221) );
  INV_X1 U4189 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4191) );
  NAND2_X1 U4190 ( .A1(n2347), .A2(REG2_REG_31__SCAN_IN), .ZN(n3418) );
  NAND2_X1 U4191 ( .A1(n2645), .A2(REG0_REG_31__SCAN_IN), .ZN(n3417) );
  OAI211_X1 U4192 ( .C1(n3419), .C2(n4191), .A(n3418), .B(n3417), .ZN(n3969)
         );
  INV_X1 U4193 ( .A(DATAI_30_), .ZN(n3420) );
  NOR2_X1 U4194 ( .A1(n2771), .A2(n3420), .ZN(n4197) );
  INV_X1 U4195 ( .A(n4197), .ZN(n3455) );
  OR2_X1 U4196 ( .A1(n3716), .A2(n3427), .ZN(n3421) );
  AND2_X1 U4197 ( .A1(n3422), .A2(n3421), .ZN(n3426) );
  INV_X1 U4198 ( .A(n3426), .ZN(n3562) );
  NOR3_X1 U4199 ( .A1(n3562), .A2(n3985), .A3(n3423), .ZN(n3453) );
  NAND2_X1 U4200 ( .A1(n3425), .A2(n3424), .ZN(n3449) );
  NAND2_X1 U4201 ( .A1(n3426), .A2(n3449), .ZN(n3431) );
  NAND2_X1 U4202 ( .A1(n3716), .A2(n3427), .ZN(n3429) );
  NAND2_X1 U4203 ( .A1(n3428), .A2(DATAI_31_), .ZN(n3970) );
  NAND2_X1 U4204 ( .A1(n3969), .A2(n3970), .ZN(n3569) );
  OAI211_X1 U4205 ( .C1(n3455), .C2(n3859), .A(n3429), .B(n3569), .ZN(n3448)
         );
  INV_X1 U4206 ( .A(n3448), .ZN(n3430) );
  NAND2_X1 U4207 ( .A1(n3431), .A2(n3430), .ZN(n3565) );
  NAND2_X1 U4208 ( .A1(n3432), .A2(n3439), .ZN(n3549) );
  NAND2_X1 U4209 ( .A1(n3508), .A2(n3509), .ZN(n3438) );
  INV_X1 U4210 ( .A(n3510), .ZN(n3437) );
  INV_X1 U4211 ( .A(n3433), .ZN(n3436) );
  INV_X1 U4212 ( .A(n3434), .ZN(n3473) );
  NAND3_X1 U4213 ( .A1(n3436), .A2(n3435), .A3(n3473), .ZN(n3513) );
  AOI211_X1 U4214 ( .C1(n3439), .C2(n3438), .A(n3437), .B(n3513), .ZN(n3548)
         );
  OAI21_X1 U4215 ( .B1(n3440), .B2(n3549), .A(n3548), .ZN(n3444) );
  INV_X1 U4216 ( .A(n3513), .ZN(n3443) );
  INV_X1 U4217 ( .A(n3441), .ZN(n3442) );
  NAND2_X1 U4218 ( .A1(n3443), .A2(n3442), .ZN(n3553) );
  NAND4_X1 U4219 ( .A1(n3444), .A2(n3555), .A3(n3554), .A4(n3553), .ZN(n3447)
         );
  INV_X1 U4220 ( .A(n3461), .ZN(n3445) );
  NAND2_X1 U4221 ( .A1(n3445), .A2(n3463), .ZN(n3558) );
  AOI21_X1 U4222 ( .B1(n3447), .B2(n3446), .A(n3558), .ZN(n3451) );
  NOR3_X1 U4223 ( .A1(n3449), .A2(n3448), .A3(n3557), .ZN(n3450) );
  OAI21_X1 U4224 ( .B1(n3451), .B2(n4001), .A(n3450), .ZN(n3452) );
  OAI21_X1 U4225 ( .B1(n3453), .B2(n3565), .A(n3452), .ZN(n3454) );
  OAI21_X1 U4226 ( .B1(n3969), .B2(n3455), .A(n3454), .ZN(n3576) );
  NAND2_X1 U4227 ( .A1(n3859), .A2(n3455), .ZN(n3566) );
  AOI21_X1 U4228 ( .B1(n3566), .B2(n3969), .A(n3970), .ZN(n3457) );
  NOR2_X1 U4229 ( .A1(n3457), .A2(n3456), .ZN(n3575) );
  XNOR2_X1 U4230 ( .A(n4216), .B(n4010), .ZN(n4002) );
  NAND3_X1 U4231 ( .A1(n3458), .A2(n2172), .A3(n4002), .ZN(n3500) );
  NAND2_X1 U4232 ( .A1(n4000), .A2(n3459), .ZN(n4020) );
  INV_X1 U4233 ( .A(n4016), .ZN(n3460) );
  OR2_X1 U4234 ( .A1(n3461), .A2(n3460), .ZN(n4035) );
  NAND2_X1 U4235 ( .A1(n3463), .A2(n3462), .ZN(n4052) );
  NOR4_X1 U4236 ( .A1(n4035), .A2(n4077), .A3(n4052), .A4(n3464), .ZN(n3498)
         );
  INV_X1 U4237 ( .A(n3465), .ZN(n3467) );
  OR2_X1 U4238 ( .A1(n3467), .A2(n3466), .ZN(n4103) );
  INV_X1 U4239 ( .A(n3969), .ZN(n3469) );
  INV_X1 U4240 ( .A(n3970), .ZN(n3468) );
  NAND2_X1 U4241 ( .A1(n3469), .A2(n3468), .ZN(n3567) );
  NAND4_X1 U4242 ( .A1(n4103), .A2(n3470), .A3(n3569), .A4(n3567), .ZN(n3479)
         );
  NAND2_X1 U4243 ( .A1(n3472), .A2(n3471), .ZN(n4129) );
  XOR2_X1 U4244 ( .A(n4197), .B(n3859), .Z(n3478) );
  NAND2_X1 U4245 ( .A1(n3473), .A2(n4124), .ZN(n4172) );
  OR4_X1 U4246 ( .A1(n4172), .A2(n3476), .A3(n3475), .A4(n3474), .ZN(n3477) );
  NOR4_X1 U4247 ( .A1(n3479), .A2(n4129), .A3(n3478), .A4(n3477), .ZN(n3497)
         );
  NAND4_X1 U4248 ( .A1(n3482), .A2(n3481), .A3(n2241), .A4(n3480), .ZN(n3488)
         );
  INV_X1 U4249 ( .A(n2650), .ZN(n3484) );
  NAND2_X1 U4250 ( .A1(n3484), .A2(n3483), .ZN(n3487) );
  NOR4_X1 U4251 ( .A1(n3488), .A2(n3487), .A3(n3486), .A4(n3485), .ZN(n3496)
         );
  INV_X1 U4252 ( .A(n3489), .ZN(n4049) );
  NOR2_X1 U4253 ( .A1(n4049), .A2(n4048), .ZN(n4086) );
  INV_X1 U4254 ( .A(n4086), .ZN(n3494) );
  NAND4_X1 U4255 ( .A1(n3491), .A2(n3594), .A3(n3490), .A4(n3533), .ZN(n3492)
         );
  NOR4_X1 U4256 ( .A1(n3494), .A2(n3493), .A3(n3492), .A4(n4498), .ZN(n3495)
         );
  NAND4_X1 U4257 ( .A1(n3498), .A2(n3497), .A3(n3496), .A4(n3495), .ZN(n3499)
         );
  NOR4_X1 U4258 ( .A1(n3501), .A2(n3500), .A3(n4020), .A4(n3499), .ZN(n3573)
         );
  INV_X1 U4259 ( .A(n3502), .ZN(n3545) );
  INV_X1 U4260 ( .A(n3536), .ZN(n3504) );
  NOR2_X1 U4261 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  NAND4_X1 U4262 ( .A1(n3505), .A2(n3511), .A3(n3535), .A4(n3528), .ZN(n3506)
         );
  NAND2_X1 U4263 ( .A1(n3507), .A2(n3506), .ZN(n3542) );
  NAND4_X1 U4264 ( .A1(n3511), .A2(n3510), .A3(n3509), .A4(n3508), .ZN(n3512)
         );
  NOR2_X1 U4265 ( .A1(n3513), .A2(n3512), .ZN(n3541) );
  INV_X1 U4266 ( .A(n3514), .ZN(n3517) );
  OAI211_X1 U4267 ( .C1(n4351), .C2(n3517), .A(n3516), .B(n3515), .ZN(n3518)
         );
  NAND3_X1 U4268 ( .A1(n3520), .A2(n3519), .A3(n3518), .ZN(n3521) );
  NAND3_X1 U4269 ( .A1(n3523), .A2(n3522), .A3(n3521), .ZN(n3524) );
  NAND3_X1 U4270 ( .A1(n3526), .A2(n3525), .A3(n3524), .ZN(n3527) );
  NAND4_X1 U4271 ( .A1(n3530), .A2(n3529), .A3(n3528), .A4(n3527), .ZN(n3531)
         );
  NAND3_X1 U4272 ( .A1(n3533), .A2(n3532), .A3(n3531), .ZN(n3534) );
  NAND3_X1 U4273 ( .A1(n3536), .A2(n3535), .A3(n3534), .ZN(n3537) );
  NAND3_X1 U4274 ( .A1(n3539), .A2(n3538), .A3(n3537), .ZN(n3540) );
  AOI22_X1 U4275 ( .A1(n3548), .A2(n3542), .B1(n3541), .B2(n3540), .ZN(n3544)
         );
  OR4_X1 U4276 ( .A1(n3546), .A2(n3545), .A3(n3544), .A4(n3543), .ZN(n3552) );
  INV_X1 U4277 ( .A(n3547), .ZN(n3550) );
  OAI21_X1 U4278 ( .B1(n3550), .B2(n3549), .A(n3548), .ZN(n3551) );
  AND4_X1 U4279 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n3556)
         );
  OAI21_X1 U4280 ( .B1(n4048), .B2(n3556), .A(n3555), .ZN(n3559) );
  AOI211_X1 U4281 ( .C1(n3560), .C2(n3559), .A(n3558), .B(n3557), .ZN(n3561)
         );
  AOI211_X1 U4282 ( .C1(n3861), .C2(n3994), .A(n3562), .B(n3561), .ZN(n3564)
         );
  NAND2_X1 U4283 ( .A1(n3564), .A2(n3563), .ZN(n3571) );
  INV_X1 U4284 ( .A(n3565), .ZN(n3570) );
  NAND2_X1 U4285 ( .A1(n3567), .A2(n3566), .ZN(n3568) );
  AOI22_X1 U4286 ( .A1(n3571), .A2(n3570), .B1(n3569), .B2(n3568), .ZN(n3572)
         );
  MUX2_X1 U4287 ( .A(n3573), .B(n3572), .S(n2640), .Z(n3574) );
  AOI21_X1 U4288 ( .B1(n3576), .B2(n3575), .A(n3574), .ZN(n3577) );
  XNOR2_X1 U4289 ( .A(n3577), .B(n3963), .ZN(n3584) );
  NAND2_X1 U4290 ( .A1(n3579), .A2(n3578), .ZN(n3580) );
  OAI211_X1 U4291 ( .C1(n3581), .C2(n3583), .A(n3580), .B(B_REG_SCAN_IN), .ZN(
        n3582) );
  OAI21_X1 U4292 ( .B1(n3584), .B2(n3583), .A(n3582), .ZN(U3239) );
  OAI21_X1 U4293 ( .B1(n3587), .B2(n3586), .A(n3585), .ZN(n4281) );
  NAND2_X1 U4294 ( .A1(n3588), .A2(n4270), .ZN(n3589) );
  AND2_X1 U4295 ( .A1(n4174), .A2(n3589), .ZN(n4277) );
  AOI22_X1 U4296 ( .A1(n4179), .A2(n3863), .B1(n4178), .B2(n4153), .ZN(n3592)
         );
  INV_X1 U4297 ( .A(n3590), .ZN(n3785) );
  AOI22_X1 U4298 ( .A1(n4360), .A2(REG2_REG_16__SCAN_IN), .B1(n3785), .B2(
        n4181), .ZN(n3591) );
  OAI211_X1 U4299 ( .C1(n3628), .C2(n4185), .A(n3592), .B(n3591), .ZN(n3597)
         );
  OAI211_X1 U4300 ( .C1(n3595), .C2(n3594), .A(n3593), .B(n4169), .ZN(n4278)
         );
  NOR2_X1 U4301 ( .A1(n4278), .A2(n4360), .ZN(n3596) );
  AOI211_X1 U4302 ( .C1(n4277), .C2(n4473), .A(n3597), .B(n3596), .ZN(n3598)
         );
  OAI21_X1 U4303 ( .B1(n4281), .B2(n4167), .A(n3598), .ZN(U3274) );
  OAI22_X1 U4304 ( .A1(n3602), .A2(n3708), .B1(n3707), .B2(n3606), .ZN(n3601)
         );
  XNOR2_X1 U4305 ( .A(n3601), .B(n3709), .ZN(n3615) );
  XNOR2_X1 U4306 ( .A(n3615), .B(n3612), .ZN(n3603) );
  XNOR2_X1 U4307 ( .A(n3616), .B(n3603), .ZN(n3604) );
  NAND2_X1 U4308 ( .A1(n3604), .A2(n3849), .ZN(n3609) );
  NOR2_X1 U4309 ( .A1(STATE_REG_SCAN_IN), .A2(n2503), .ZN(n4410) );
  OAI22_X1 U4310 ( .A1(n2045), .A2(n3606), .B1(n3605), .B2(n3851), .ZN(n3607)
         );
  AOI211_X1 U4311 ( .C1(n3854), .C2(n3864), .A(n4410), .B(n3607), .ZN(n3608)
         );
  OAI211_X1 U4312 ( .C1(n3858), .C2(n3610), .A(n3609), .B(n3608), .ZN(U3231)
         );
  NAND2_X1 U4313 ( .A1(n3614), .A2(n3611), .ZN(n3613) );
  INV_X1 U4314 ( .A(n3614), .ZN(n3616) );
  OAI22_X1 U4315 ( .A1(n4289), .A2(n3708), .B1(n3707), .B2(n3617), .ZN(n3618)
         );
  XNOR2_X1 U4316 ( .A(n3618), .B(n3709), .ZN(n3622) );
  OR2_X1 U4317 ( .A1(n4289), .A2(n2964), .ZN(n3620) );
  NAND2_X1 U4318 ( .A1(n3677), .A2(n3747), .ZN(n3619) );
  NAND2_X1 U4319 ( .A1(n3620), .A2(n3619), .ZN(n3621) );
  AND2_X1 U4320 ( .A1(n3622), .A2(n3621), .ZN(n3744) );
  OAI22_X1 U4321 ( .A1(n4269), .A2(n3708), .B1(n3707), .B2(n3852), .ZN(n3623)
         );
  XOR2_X1 U4322 ( .A(n3709), .B(n3623), .Z(n3626) );
  OR2_X1 U4323 ( .A1(n4269), .A2(n2964), .ZN(n3625) );
  INV_X1 U4324 ( .A(n3708), .ZN(n3697) );
  NAND2_X1 U4325 ( .A1(n3697), .A2(n4283), .ZN(n3624) );
  NAND2_X1 U4326 ( .A1(n3625), .A2(n3624), .ZN(n3847) );
  OAI22_X1 U4327 ( .A1(n4264), .A2(n2964), .B1(n3702), .B2(n3628), .ZN(n3632)
         );
  OAI22_X1 U4328 ( .A1(n4264), .A2(n3708), .B1(n3707), .B2(n3628), .ZN(n3629)
         );
  XNOR2_X1 U4329 ( .A(n3629), .B(n3709), .ZN(n3631) );
  XOR2_X1 U4330 ( .A(n3632), .B(n3631), .Z(n3780) );
  OAI22_X1 U4331 ( .A1(n4274), .A2(n3702), .B1(n3707), .B2(n4186), .ZN(n3636)
         );
  XNOR2_X1 U4332 ( .A(n3636), .B(n3709), .ZN(n3789) );
  OAI22_X1 U4333 ( .A1(n4274), .A2(n2964), .B1(n3702), .B2(n4186), .ZN(n3790)
         );
  NOR2_X1 U4334 ( .A1(n3789), .A2(n3790), .ZN(n3638) );
  NAND2_X1 U4335 ( .A1(n3789), .A2(n3790), .ZN(n3637) );
  INV_X1 U4336 ( .A(n3708), .ZN(n3677) );
  NAND2_X1 U4337 ( .A1(n4261), .A2(n3677), .ZN(n3640) );
  NAND2_X1 U4338 ( .A1(n3698), .A2(n4152), .ZN(n3639) );
  NAND2_X1 U4339 ( .A1(n3640), .A2(n3639), .ZN(n3641) );
  XNOR2_X1 U4340 ( .A(n3641), .B(n3173), .ZN(n3644) );
  NOR2_X1 U4341 ( .A1(n3702), .A2(n4159), .ZN(n3642) );
  AOI21_X1 U4342 ( .B1(n4261), .B2(n3704), .A(n3642), .ZN(n3643) );
  NOR2_X1 U4343 ( .A1(n3644), .A2(n3643), .ZN(n3825) );
  NAND2_X1 U4344 ( .A1(n3644), .A2(n3643), .ZN(n3826) );
  OAI22_X1 U4345 ( .A1(n4155), .A2(n2964), .B1(n3702), .B2(n4137), .ZN(n3646)
         );
  OAI22_X1 U4346 ( .A1(n4155), .A2(n3708), .B1(n3707), .B2(n4137), .ZN(n3645)
         );
  XNOR2_X1 U4347 ( .A(n3645), .B(n3709), .ZN(n3647) );
  NAND2_X1 U4348 ( .A1(n3764), .A2(n3765), .ZN(n3649) );
  NAND2_X1 U4349 ( .A1(n4241), .A2(n3677), .ZN(n3651) );
  NAND2_X1 U4350 ( .A1(n3698), .A2(n4105), .ZN(n3650) );
  NAND2_X1 U4351 ( .A1(n3651), .A2(n3650), .ZN(n3652) );
  XNOR2_X1 U4352 ( .A(n3652), .B(n3709), .ZN(n3655) );
  NAND2_X1 U4353 ( .A1(n4241), .A2(n3704), .ZN(n3654) );
  NAND2_X1 U4354 ( .A1(n3697), .A2(n4105), .ZN(n3653) );
  NAND2_X1 U4355 ( .A1(n3654), .A2(n3653), .ZN(n3656) );
  NAND2_X1 U4356 ( .A1(n3655), .A2(n3656), .ZN(n3806) );
  INV_X1 U4357 ( .A(n3655), .ZN(n3658) );
  INV_X1 U4358 ( .A(n3656), .ZN(n3657) );
  NAND2_X1 U4359 ( .A1(n3658), .A2(n3657), .ZN(n3808) );
  NAND2_X1 U4360 ( .A1(n4106), .A2(n3677), .ZN(n3660) );
  NAND2_X1 U4361 ( .A1(n3698), .A2(n4239), .ZN(n3659) );
  NAND2_X1 U4362 ( .A1(n3660), .A2(n3659), .ZN(n3661) );
  XNOR2_X1 U4363 ( .A(n3661), .B(n3709), .ZN(n3771) );
  NAND2_X1 U4364 ( .A1(n4106), .A2(n3704), .ZN(n3663) );
  NAND2_X1 U4365 ( .A1(n3677), .A2(n4239), .ZN(n3662) );
  NAND2_X1 U4366 ( .A1(n3663), .A2(n3662), .ZN(n3770) );
  OAI22_X1 U4367 ( .A1(n4244), .A2(n3708), .B1(n3707), .B2(n4072), .ZN(n3664)
         );
  XNOR2_X1 U4368 ( .A(n3664), .B(n3709), .ZN(n3667) );
  OAI22_X1 U4369 ( .A1(n4244), .A2(n2964), .B1(n3702), .B2(n4072), .ZN(n3666)
         );
  XNOR2_X1 U4370 ( .A(n3667), .B(n3666), .ZN(n3817) );
  OAI22_X1 U4371 ( .A1(n3819), .A2(n3708), .B1(n3707), .B2(n4058), .ZN(n3665)
         );
  XNOR2_X1 U4372 ( .A(n3665), .B(n3709), .ZN(n3669) );
  OAI22_X1 U4373 ( .A1(n3819), .A2(n2964), .B1(n3702), .B2(n4058), .ZN(n3668)
         );
  XNOR2_X1 U4374 ( .A(n3669), .B(n3668), .ZN(n3755) );
  NOR2_X1 U4375 ( .A1(n3667), .A2(n3666), .ZN(n3756) );
  NAND2_X1 U4376 ( .A1(n3669), .A2(n3668), .ZN(n3672) );
  NOR2_X1 U4377 ( .A1(n3702), .A2(n4042), .ZN(n3670) );
  AOI21_X1 U4378 ( .B1(n4213), .B2(n3704), .A(n3670), .ZN(n3673) );
  OAI22_X1 U4379 ( .A1(n4054), .A2(n3708), .B1(n3707), .B2(n4042), .ZN(n3671)
         );
  XNOR2_X1 U4380 ( .A(n3671), .B(n3709), .ZN(n3799) );
  NAND2_X1 U4381 ( .A1(n3797), .A2(n3799), .ZN(n3676) );
  INV_X1 U4382 ( .A(n3673), .ZN(n3674) );
  NAND2_X1 U4383 ( .A1(n3675), .A2(n3674), .ZN(n3796) );
  NAND2_X1 U4384 ( .A1(n3676), .A2(n3796), .ZN(n3691) );
  NAND2_X1 U4385 ( .A1(n4038), .A2(n3677), .ZN(n3679) );
  NAND2_X1 U4386 ( .A1(n3698), .A2(n4212), .ZN(n3678) );
  NAND2_X1 U4387 ( .A1(n3679), .A2(n3678), .ZN(n3680) );
  XNOR2_X1 U4388 ( .A(n3680), .B(n3173), .ZN(n3683) );
  NOR2_X1 U4389 ( .A1(n3702), .A2(n4027), .ZN(n3681) );
  AOI21_X1 U4390 ( .B1(n4038), .B2(n3704), .A(n3681), .ZN(n3682) );
  NOR2_X1 U4391 ( .A1(n3683), .A2(n3682), .ZN(n3689) );
  NAND2_X1 U4392 ( .A1(n3683), .A2(n3682), .ZN(n3690) );
  NOR2_X1 U4393 ( .A1(n3689), .A2(n2198), .ZN(n3684) );
  XNOR2_X1 U4394 ( .A(n3691), .B(n3684), .ZN(n3688) );
  OAI22_X1 U4395 ( .A1(n2045), .A2(n4027), .B1(n4054), .B2(n3851), .ZN(n3686)
         );
  OAI22_X1 U4396 ( .A1(n4216), .A2(n3840), .B1(STATE_REG_SCAN_IN), .B2(n4541), 
        .ZN(n3685) );
  AOI211_X1 U4397 ( .C1(n4024), .C2(n3843), .A(n3686), .B(n3685), .ZN(n3687)
         );
  OAI21_X1 U4398 ( .B1(n3688), .B2(n3845), .A(n3687), .ZN(U3222) );
  OAI22_X1 U4399 ( .A1(n4216), .A2(n3708), .B1(n3707), .B2(n4010), .ZN(n3692)
         );
  XNOR2_X1 U4400 ( .A(n3692), .B(n3709), .ZN(n3693) );
  OAI22_X1 U4401 ( .A1(n4216), .A2(n2964), .B1(n3702), .B2(n4010), .ZN(n3694)
         );
  NAND2_X1 U4402 ( .A1(n3693), .A2(n3694), .ZN(n3834) );
  INV_X1 U4403 ( .A(n3693), .ZN(n3696) );
  INV_X1 U4404 ( .A(n3694), .ZN(n3695) );
  NAND2_X1 U4405 ( .A1(n3696), .A2(n3695), .ZN(n3835) );
  NAND2_X1 U4406 ( .A1(n3861), .A2(n3697), .ZN(n3700) );
  NAND2_X1 U4407 ( .A1(n3698), .A2(n4199), .ZN(n3699) );
  NAND2_X1 U4408 ( .A1(n3700), .A2(n3699), .ZN(n3701) );
  XNOR2_X1 U4409 ( .A(n3701), .B(n3173), .ZN(n3705) );
  NOR2_X1 U4410 ( .A1(n3702), .A2(n3994), .ZN(n3703) );
  AOI21_X1 U4411 ( .B1(n3861), .B2(n3704), .A(n3703), .ZN(n3706) );
  OAI22_X1 U4412 ( .A1(n4202), .A2(n3708), .B1(n3707), .B2(n3729), .ZN(n3712)
         );
  OAI22_X1 U4413 ( .A1(n4202), .A2(n2964), .B1(n3702), .B2(n3729), .ZN(n3710)
         );
  XNOR2_X1 U4414 ( .A(n3710), .B(n3709), .ZN(n3711) );
  XOR2_X1 U4415 ( .A(n3712), .B(n3711), .Z(n3713) );
  XNOR2_X1 U4416 ( .A(n3714), .B(n3713), .ZN(n3720) );
  OAI22_X1 U4417 ( .A1(n4005), .A2(n3851), .B1(STATE_REG_SCAN_IN), .B2(n3715), 
        .ZN(n3718) );
  OAI22_X1 U4418 ( .A1(n3716), .A2(n3840), .B1(n2045), .B2(n3729), .ZN(n3717)
         );
  AOI211_X1 U4419 ( .C1(n3726), .C2(n3843), .A(n3718), .B(n3717), .ZN(n3719)
         );
  OAI21_X1 U4420 ( .B1(n3720), .B2(n3845), .A(n3719), .ZN(U3217) );
  INV_X1 U4421 ( .A(D_REG_0__SCAN_IN), .ZN(n3724) );
  NOR2_X1 U4422 ( .A1(n4480), .A2(n3721), .ZN(n3723) );
  AOI22_X1 U4423 ( .A1(n4479), .A2(n3724), .B1(n3723), .B2(n3722), .ZN(U3458)
         );
  INV_X1 U4424 ( .A(n3725), .ZN(n3733) );
  AOI22_X1 U4425 ( .A1(n3860), .A2(n4178), .B1(n4179), .B2(n3861), .ZN(n3728)
         );
  AOI22_X1 U4426 ( .A1(n3726), .A2(n4181), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4360), .ZN(n3727) );
  OAI211_X1 U4427 ( .C1(n3729), .C2(n4185), .A(n3728), .B(n3727), .ZN(n3732)
         );
  NOR2_X1 U4428 ( .A1(n3730), .A2(n4360), .ZN(n3731) );
  AOI211_X1 U4429 ( .C1(n4473), .C2(n3733), .A(n3732), .B(n3731), .ZN(n3734)
         );
  OAI21_X1 U4430 ( .B1(n3735), .B2(n4167), .A(n3734), .ZN(U3262) );
  INV_X1 U4431 ( .A(n3737), .ZN(n3991) );
  OAI22_X1 U4432 ( .A1(n4216), .A2(n3851), .B1(n2045), .B2(n3994), .ZN(n3739)
         );
  OAI22_X1 U4433 ( .A1(n4202), .A2(n3840), .B1(STATE_REG_SCAN_IN), .B2(n4554), 
        .ZN(n3738) );
  AOI211_X1 U4434 ( .C1(n3991), .C2(n3843), .A(n3739), .B(n3738), .ZN(n3740)
         );
  OAI21_X1 U4435 ( .B1(n3741), .B2(n3845), .A(n3740), .ZN(U3211) );
  INV_X1 U4436 ( .A(n3743), .ZN(n3745) );
  NOR2_X1 U4437 ( .A1(n3745), .A2(n3744), .ZN(n3746) );
  XNOR2_X1 U4438 ( .A(n3742), .B(n3746), .ZN(n3754) );
  AOI22_X1 U4439 ( .A1(n3782), .A2(n3747), .B1(n3781), .B2(n3865), .ZN(n3750)
         );
  NOR2_X1 U4440 ( .A1(n3748), .A2(STATE_REG_SCAN_IN), .ZN(n4421) );
  INV_X1 U4441 ( .A(n4421), .ZN(n3749) );
  OAI211_X1 U4442 ( .C1(n4269), .C2(n3840), .A(n3750), .B(n3749), .ZN(n3751)
         );
  AOI21_X1 U4443 ( .B1(n3752), .B2(n3843), .A(n3751), .ZN(n3753) );
  OAI21_X1 U4444 ( .B1(n3754), .B2(n3845), .A(n3753), .ZN(U3212) );
  OAI21_X1 U4445 ( .B1(n2055), .B2(n3756), .A(n3755), .ZN(n3759) );
  NAND3_X1 U4446 ( .A1(n3759), .A2(n3849), .A3(n3758), .ZN(n3763) );
  OAI22_X1 U4447 ( .A1(n2045), .A2(n4058), .B1(n4054), .B2(n3840), .ZN(n3761)
         );
  OAI22_X1 U4448 ( .A1(n4244), .A2(n3851), .B1(STATE_REG_SCAN_IN), .B2(n4627), 
        .ZN(n3760) );
  NOR2_X1 U4449 ( .A1(n3761), .A2(n3760), .ZN(n3762) );
  OAI211_X1 U4450 ( .C1(n3858), .C2(n4059), .A(n3763), .B(n3762), .ZN(U3213)
         );
  XOR2_X1 U4451 ( .A(n3765), .B(n3764), .Z(n3769) );
  INV_X1 U4452 ( .A(n4241), .ZN(n4135) );
  AOI22_X1 U4453 ( .A1(n3782), .A2(n4132), .B1(n3781), .B2(n4261), .ZN(n3766)
         );
  NAND2_X1 U4454 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3962) );
  OAI211_X1 U4455 ( .C1(n4135), .C2(n3840), .A(n3766), .B(n3962), .ZN(n3767)
         );
  AOI21_X1 U4456 ( .B1(n4140), .B2(n3843), .A(n3767), .ZN(n3768) );
  OAI21_X1 U4457 ( .B1(n3769), .B2(n3845), .A(n3768), .ZN(U3216) );
  XNOR2_X1 U4458 ( .A(n3771), .B(n3770), .ZN(n3772) );
  XNOR2_X1 U4459 ( .A(n3773), .B(n3772), .ZN(n3777) );
  OAI22_X1 U4460 ( .A1(n4244), .A2(n3840), .B1(STATE_REG_SCAN_IN), .B2(n4630), 
        .ZN(n3775) );
  OAI22_X1 U4461 ( .A1(n2045), .A2(n4094), .B1(n4135), .B2(n3851), .ZN(n3774)
         );
  AOI211_X1 U4462 ( .C1(n4091), .C2(n3843), .A(n3775), .B(n3774), .ZN(n3776)
         );
  OAI21_X1 U4463 ( .B1(n3777), .B2(n3845), .A(n3776), .ZN(U3220) );
  INV_X1 U4464 ( .A(n2286), .ZN(n3778) );
  XOR2_X1 U4465 ( .A(n3780), .B(n3779), .Z(n3787) );
  AOI22_X1 U4466 ( .A1(n3782), .A2(n4270), .B1(n3781), .B2(n3863), .ZN(n3783)
         );
  NAND2_X1 U4467 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4437) );
  OAI211_X1 U4468 ( .C1(n4274), .C2(n3840), .A(n3783), .B(n4437), .ZN(n3784)
         );
  AOI21_X1 U4469 ( .B1(n3785), .B2(n3843), .A(n3784), .ZN(n3786) );
  OAI21_X1 U4470 ( .B1(n3787), .B2(n3845), .A(n3786), .ZN(U3223) );
  XOR2_X1 U4471 ( .A(n3790), .B(n3789), .Z(n3791) );
  XNOR2_X1 U4472 ( .A(n3788), .B(n3791), .ZN(n3792) );
  NAND2_X1 U4473 ( .A1(n3792), .A2(n3849), .ZN(n3795) );
  NOR2_X1 U4474 ( .A1(n4626), .A2(STATE_REG_SCAN_IN), .ZN(n4450) );
  OAI22_X1 U4475 ( .A1(n2045), .A2(n4186), .B1(n4264), .B2(n3851), .ZN(n3793)
         );
  AOI211_X1 U4476 ( .C1(n3854), .C2(n4261), .A(n4450), .B(n3793), .ZN(n3794)
         );
  OAI211_X1 U4477 ( .C1(n3858), .C2(n4180), .A(n3795), .B(n3794), .ZN(U3225)
         );
  NAND2_X1 U4478 ( .A1(n3796), .A2(n3797), .ZN(n3798) );
  XOR2_X1 U4479 ( .A(n3799), .B(n3798), .Z(n3803) );
  OAI22_X1 U4480 ( .A1(n3819), .A2(n3851), .B1(STATE_REG_SCAN_IN), .B2(n4635), 
        .ZN(n3801) );
  OAI22_X1 U4481 ( .A1(n4225), .A2(n3840), .B1(n2045), .B2(n4042), .ZN(n3800)
         );
  AOI211_X1 U4482 ( .C1(n4039), .C2(n3843), .A(n3801), .B(n3800), .ZN(n3802)
         );
  OAI21_X1 U4483 ( .B1(n3803), .B2(n3845), .A(n3802), .ZN(U3226) );
  INV_X1 U4484 ( .A(n3804), .ZN(n3809) );
  AOI21_X1 U4485 ( .B1(n3808), .B2(n3806), .A(n3805), .ZN(n3807) );
  AOI21_X1 U4486 ( .B1(n3809), .B2(n3808), .A(n3807), .ZN(n3815) );
  INV_X1 U4487 ( .A(n3810), .ZN(n4117) );
  OAI22_X1 U4488 ( .A1(n3840), .A2(n4067), .B1(STATE_REG_SCAN_IN), .B2(n3811), 
        .ZN(n3813) );
  OAI22_X1 U4489 ( .A1(n2045), .A2(n4115), .B1(n4155), .B2(n3851), .ZN(n3812)
         );
  AOI211_X1 U4490 ( .C1(n4117), .C2(n3843), .A(n3813), .B(n3812), .ZN(n3814)
         );
  OAI21_X1 U4491 ( .B1(n3815), .B2(n3845), .A(n3814), .ZN(U3230) );
  AOI21_X1 U4492 ( .B1(n3817), .B2(n3816), .A(n2055), .ZN(n3823) );
  OAI22_X1 U4493 ( .A1(n3851), .A2(n4067), .B1(STATE_REG_SCAN_IN), .B2(n3818), 
        .ZN(n3821) );
  OAI22_X1 U4494 ( .A1(n2045), .A2(n4072), .B1(n3819), .B2(n3840), .ZN(n3820)
         );
  AOI211_X1 U4495 ( .C1(n4075), .C2(n3843), .A(n3821), .B(n3820), .ZN(n3822)
         );
  OAI21_X1 U4496 ( .B1(n3823), .B2(n3845), .A(n3822), .ZN(U3232) );
  INV_X1 U4497 ( .A(n3825), .ZN(n3827) );
  NAND2_X1 U4498 ( .A1(n3827), .A2(n3826), .ZN(n3828) );
  XNOR2_X1 U4499 ( .A(n3824), .B(n3828), .ZN(n3829) );
  NAND2_X1 U4500 ( .A1(n3829), .A2(n3849), .ZN(n3832) );
  AND2_X1 U4501 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4459) );
  OAI22_X1 U4502 ( .A1(n2045), .A2(n4159), .B1(n4274), .B2(n3851), .ZN(n3830)
         );
  AOI211_X1 U4503 ( .C1(n3854), .C2(n3862), .A(n4459), .B(n3830), .ZN(n3831)
         );
  OAI211_X1 U4504 ( .C1(n3858), .C2(n4161), .A(n3832), .B(n3831), .ZN(U3235)
         );
  NAND2_X1 U4505 ( .A1(n3835), .A2(n3834), .ZN(n3836) );
  XNOR2_X1 U4506 ( .A(n3833), .B(n3836), .ZN(n3846) );
  INV_X1 U4507 ( .A(n3837), .ZN(n4011) );
  OAI22_X1 U4508 ( .A1(n4225), .A2(n3851), .B1(STATE_REG_SCAN_IN), .B2(n3838), 
        .ZN(n3842) );
  OAI22_X1 U4509 ( .A1(n4005), .A2(n3840), .B1(n2045), .B2(n4010), .ZN(n3841)
         );
  AOI211_X1 U4510 ( .C1(n4011), .C2(n3843), .A(n3842), .B(n3841), .ZN(n3844)
         );
  OAI21_X1 U4511 ( .B1(n3846), .B2(n3845), .A(n3844), .ZN(U3237) );
  XNOR2_X1 U4512 ( .A(n3848), .B(n3847), .ZN(n3850) );
  NAND2_X1 U4513 ( .A1(n3850), .A2(n3849), .ZN(n3856) );
  AND2_X1 U4514 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4430) );
  OAI22_X1 U4515 ( .A1(n2045), .A2(n3852), .B1(n4289), .B2(n3851), .ZN(n3853)
         );
  AOI211_X1 U4516 ( .C1(n3854), .C2(n4285), .A(n4430), .B(n3853), .ZN(n3855)
         );
  OAI211_X1 U4517 ( .C1(n3858), .C2(n3857), .A(n3856), .B(n3855), .ZN(U3238)
         );
  MUX2_X1 U4518 ( .A(DATAO_REG_31__SCAN_IN), .B(n3969), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4519 ( .A(DATAO_REG_30__SCAN_IN), .B(n3859), .S(n3872), .Z(U3580)
         );
  MUX2_X1 U4520 ( .A(DATAO_REG_29__SCAN_IN), .B(n3860), .S(n3872), .Z(U3579)
         );
  MUX2_X1 U4521 ( .A(DATAO_REG_28__SCAN_IN), .B(n3990), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4522 ( .A(DATAO_REG_27__SCAN_IN), .B(n3861), .S(n3872), .Z(U3577)
         );
  MUX2_X1 U4523 ( .A(DATAO_REG_26__SCAN_IN), .B(n4200), .S(n3872), .Z(U3576)
         );
  MUX2_X1 U4524 ( .A(DATAO_REG_25__SCAN_IN), .B(n4038), .S(n3872), .Z(U3575)
         );
  MUX2_X1 U4525 ( .A(DATAO_REG_24__SCAN_IN), .B(n4213), .S(n3872), .Z(U3574)
         );
  MUX2_X1 U4526 ( .A(DATAO_REG_23__SCAN_IN), .B(n4222), .S(n3872), .Z(U3573)
         );
  MUX2_X1 U4527 ( .A(DATAO_REG_22__SCAN_IN), .B(n4090), .S(n3872), .Z(U3572)
         );
  MUX2_X1 U4528 ( .A(DATAO_REG_21__SCAN_IN), .B(n4106), .S(n3872), .Z(U3571)
         );
  MUX2_X1 U4529 ( .A(DATAO_REG_20__SCAN_IN), .B(n4241), .S(n3872), .Z(U3570)
         );
  MUX2_X1 U4530 ( .A(DATAO_REG_19__SCAN_IN), .B(n3862), .S(n3872), .Z(U3569)
         );
  MUX2_X1 U4531 ( .A(DATAO_REG_18__SCAN_IN), .B(n4261), .S(n3872), .Z(U3568)
         );
  MUX2_X1 U4532 ( .A(DATAO_REG_17__SCAN_IN), .B(n4153), .S(n3872), .Z(U3567)
         );
  MUX2_X1 U4533 ( .A(DATAO_REG_16__SCAN_IN), .B(n4285), .S(n3872), .Z(U3566)
         );
  MUX2_X1 U4534 ( .A(DATAO_REG_15__SCAN_IN), .B(n3863), .S(n3872), .Z(U3565)
         );
  MUX2_X1 U4535 ( .A(DATAO_REG_14__SCAN_IN), .B(n3864), .S(n3872), .Z(U3564)
         );
  MUX2_X1 U4536 ( .A(DATAO_REG_13__SCAN_IN), .B(n3865), .S(n3872), .Z(U3563)
         );
  MUX2_X1 U4537 ( .A(DATAO_REG_12__SCAN_IN), .B(n3866), .S(n3872), .Z(U3562)
         );
  MUX2_X1 U4538 ( .A(DATAO_REG_11__SCAN_IN), .B(n3867), .S(n3872), .Z(U3561)
         );
  MUX2_X1 U4539 ( .A(DATAO_REG_10__SCAN_IN), .B(n3868), .S(n3872), .Z(U3560)
         );
  MUX2_X1 U4540 ( .A(DATAO_REG_9__SCAN_IN), .B(n3869), .S(n3872), .Z(U3559) );
  MUX2_X1 U4541 ( .A(DATAO_REG_8__SCAN_IN), .B(n3870), .S(n3872), .Z(U3558) );
  MUX2_X1 U4542 ( .A(DATAO_REG_7__SCAN_IN), .B(n3871), .S(n3872), .Z(U3557) );
  MUX2_X1 U4543 ( .A(DATAO_REG_6__SCAN_IN), .B(n3873), .S(n3872), .Z(U3556) );
  MUX2_X1 U4544 ( .A(DATAO_REG_5__SCAN_IN), .B(n3874), .S(U4043), .Z(U3555) );
  MUX2_X1 U4545 ( .A(DATAO_REG_4__SCAN_IN), .B(n3875), .S(U4043), .Z(U3554) );
  MUX2_X1 U4546 ( .A(DATAO_REG_3__SCAN_IN), .B(n3876), .S(U4043), .Z(U3553) );
  MUX2_X1 U4547 ( .A(DATAO_REG_2__SCAN_IN), .B(n2941), .S(U4043), .Z(U3552) );
  MUX2_X1 U4548 ( .A(DATAO_REG_1__SCAN_IN), .B(n3877), .S(U4043), .Z(U3551) );
  MUX2_X1 U4549 ( .A(DATAO_REG_0__SCAN_IN), .B(n2857), .S(U4043), .Z(U3550) );
  OAI211_X1 U4550 ( .C1(n3881), .C2(n3880), .A(n4462), .B(n3879), .ZN(n3886)
         );
  OAI211_X1 U4551 ( .C1(n2790), .C2(n3883), .A(n4406), .B(n3895), .ZN(n3885)
         );
  AOI22_X1 U4552 ( .A1(n4460), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3884) );
  NAND4_X1 U4553 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(U3241)
         );
  NOR2_X1 U4554 ( .A1(n3888), .A2(STATE_REG_SCAN_IN), .ZN(n3889) );
  AOI21_X1 U4555 ( .B1(n4460), .B2(ADDR_REG_2__SCAN_IN), .A(n3889), .ZN(n3890)
         );
  OAI21_X1 U4556 ( .B1(n4467), .B2(n3891), .A(n3890), .ZN(n3892) );
  INV_X1 U4557 ( .A(n3892), .ZN(n3904) );
  MUX2_X1 U4558 ( .A(n3893), .B(REG2_REG_2__SCAN_IN), .S(n2048), .Z(n3896) );
  NAND3_X1 U4559 ( .A1(n3896), .A2(n3895), .A3(n3894), .ZN(n3897) );
  NAND3_X1 U4560 ( .A1(n4406), .A2(n3898), .A3(n3897), .ZN(n3903) );
  OAI211_X1 U4561 ( .C1(n3901), .C2(n3900), .A(n4462), .B(n3899), .ZN(n3902)
         );
  NAND4_X1 U4562 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(U3242)
         );
  NAND2_X1 U4563 ( .A1(n3906), .A2(n4358), .ZN(n3915) );
  OAI211_X1 U4564 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3908), .A(n4462), .B(n3907), 
        .ZN(n3914) );
  AOI22_X1 U4565 ( .A1(n4460), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3913) );
  XNOR2_X1 U4566 ( .A(n3910), .B(n3909), .ZN(n3911) );
  NAND2_X1 U4567 ( .A1(n4406), .A2(n3911), .ZN(n3912) );
  NAND4_X1 U4568 ( .A1(n3915), .A2(n3914), .A3(n3913), .A4(n3912), .ZN(U3243)
         );
  MUX2_X1 U4569 ( .A(REG2_REG_19__SCAN_IN), .B(n4142), .S(n4352), .Z(n3932) );
  INV_X1 U4570 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4571 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4482), .B1(n3933), .B2(
        n3916), .ZN(n4458) );
  NOR2_X1 U4572 ( .A1(n3957), .A2(REG2_REG_17__SCAN_IN), .ZN(n3917) );
  AOI21_X1 U4573 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3957), .A(n3917), .ZN(n4448) );
  INV_X1 U4574 ( .A(n3950), .ZN(n4487) );
  NOR2_X1 U4575 ( .A1(n4405), .A2(n4417), .ZN(n4404) );
  NAND2_X1 U4576 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3934), .ZN(n3923) );
  INV_X1 U4577 ( .A(n3934), .ZN(n4491) );
  AOI22_X1 U4578 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3934), .B1(n4491), .B2(
        n3237), .ZN(n4389) );
  NAND2_X1 U4579 ( .A1(n3935), .A2(REG2_REG_9__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4580 ( .A1(n3935), .A2(REG2_REG_9__SCAN_IN), .B1(n2457), .B2(n4493), .ZN(n4369) );
  OAI22_X1 U4581 ( .A1(n3919), .A2(n4470), .B1(n3918), .B2(n4353), .ZN(n4368)
         );
  NAND2_X1 U4582 ( .A1(n4369), .A2(n4368), .ZN(n4367) );
  NAND2_X1 U4583 ( .A1(n3942), .A2(n3921), .ZN(n3922) );
  INV_X1 U4584 ( .A(n3942), .ZN(n4492) );
  XNOR2_X1 U4585 ( .A(n3921), .B(n4492), .ZN(n4376) );
  NAND2_X1 U4586 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4376), .ZN(n4375) );
  NAND2_X1 U4587 ( .A1(n3922), .A2(n4375), .ZN(n4388) );
  NAND2_X1 U4588 ( .A1(n4389), .A2(n4388), .ZN(n4387) );
  NAND2_X1 U4589 ( .A1(n3946), .A2(n3924), .ZN(n3925) );
  XNOR2_X1 U4590 ( .A(n3924), .B(n4490), .ZN(n4396) );
  NOR2_X1 U4591 ( .A1(n4487), .A2(n3926), .ZN(n3927) );
  NOR2_X1 U4592 ( .A1(n2341), .A2(n4419), .ZN(n4418) );
  NAND2_X1 U4593 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4485), .ZN(n3928) );
  OAI21_X1 U4594 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4485), .A(n3928), .ZN(n4427) );
  NOR2_X1 U4595 ( .A1(n4428), .A2(n4427), .ZN(n4426) );
  INV_X1 U4596 ( .A(n3954), .ZN(n4484) );
  NAND2_X1 U4597 ( .A1(n3929), .A2(n4484), .ZN(n3930) );
  AOI21_X1 U4598 ( .B1(n3933), .B2(REG2_REG_18__SCAN_IN), .A(n4457), .ZN(n3931) );
  XOR2_X1 U4599 ( .A(n3932), .B(n3931), .Z(n3967) );
  INV_X1 U4600 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4601 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3933), .B1(n4482), .B2(
        n3959), .ZN(n4464) );
  NOR2_X1 U4602 ( .A1(n3957), .A2(REG1_REG_17__SCAN_IN), .ZN(n3958) );
  NAND2_X1 U4603 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4485), .ZN(n3953) );
  INV_X1 U4604 ( .A(n4485), .ZN(n4436) );
  AOI22_X1 U4605 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4485), .B1(n4436), .B2(
        n4292), .ZN(n4433) );
  NAND2_X1 U4606 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4488), .ZN(n3949) );
  AOI22_X1 U4607 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4488), .B1(n4417), .B2(
        n3380), .ZN(n4414) );
  NAND2_X1 U4608 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3934), .ZN(n3945) );
  AOI22_X1 U4609 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3934), .B1(n4491), .B2(
        n3288), .ZN(n4386) );
  NAND2_X1 U4610 ( .A1(n3935), .A2(REG1_REG_9__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4611 ( .A1(n3935), .A2(REG1_REG_9__SCAN_IN), .B1(n2456), .B2(n4493), .ZN(n4366) );
  INV_X1 U4612 ( .A(n3937), .ZN(n3938) );
  OAI22_X1 U4613 ( .A1(n3940), .A2(n3939), .B1(n3938), .B2(n4353), .ZN(n4365)
         );
  NAND2_X1 U4614 ( .A1(n4366), .A2(n4365), .ZN(n4364) );
  NAND2_X1 U4615 ( .A1(n3941), .A2(n4364), .ZN(n3943) );
  NAND2_X1 U4616 ( .A1(n3942), .A2(n3943), .ZN(n3944) );
  XNOR2_X1 U4617 ( .A(n3943), .B(n4492), .ZN(n4381) );
  NAND2_X1 U4618 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4381), .ZN(n4380) );
  NAND2_X1 U4619 ( .A1(n3944), .A2(n4380), .ZN(n4385) );
  NAND2_X1 U4620 ( .A1(n4386), .A2(n4385), .ZN(n4384) );
  NAND2_X1 U4621 ( .A1(n3945), .A2(n4384), .ZN(n3947) );
  NAND2_X1 U4622 ( .A1(n3946), .A2(n3947), .ZN(n3948) );
  XNOR2_X1 U4623 ( .A(n3947), .B(n4490), .ZN(n4401) );
  NAND2_X1 U4624 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4401), .ZN(n4400) );
  NAND2_X1 U4625 ( .A1(n3948), .A2(n4400), .ZN(n4413) );
  NAND2_X1 U4626 ( .A1(n4414), .A2(n4413), .ZN(n4412) );
  NAND2_X1 U4627 ( .A1(n3949), .A2(n4412), .ZN(n3951) );
  NAND2_X1 U4628 ( .A1(n3950), .A2(n3951), .ZN(n3952) );
  XNOR2_X1 U4629 ( .A(n3951), .B(n4487), .ZN(n4423) );
  NAND2_X1 U4630 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4423), .ZN(n4422) );
  NAND2_X1 U4631 ( .A1(n3952), .A2(n4422), .ZN(n4432) );
  NAND2_X1 U4632 ( .A1(n4433), .A2(n4432), .ZN(n4431) );
  NOR2_X1 U4633 ( .A1(n3954), .A2(n3955), .ZN(n3956) );
  AOI22_X1 U4634 ( .A1(n3957), .A2(n4267), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4483), .ZN(n4451) );
  NOR2_X1 U4635 ( .A1(n4452), .A2(n4451), .ZN(n4453) );
  MUX2_X1 U4636 ( .A(n4255), .B(REG1_REG_19__SCAN_IN), .S(n4352), .Z(n3960) );
  NAND2_X1 U4637 ( .A1(n4460), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3961) );
  OAI211_X1 U4638 ( .C1(n4467), .C2(n3963), .A(n3962), .B(n3961), .ZN(n3964)
         );
  AOI21_X1 U4639 ( .B1(n3965), .B2(n4462), .A(n3964), .ZN(n3966) );
  OAI21_X1 U4640 ( .B1(n3967), .B2(n4456), .A(n3966), .ZN(U3259) );
  XNOR2_X1 U4641 ( .A(n4194), .B(n3970), .ZN(n4298) );
  NAND2_X1 U4642 ( .A1(n3969), .A2(n3968), .ZN(n4195) );
  OAI21_X1 U4643 ( .B1(n3970), .B2(n4066), .A(n4195), .ZN(n4295) );
  NAND2_X1 U4644 ( .A1(n4164), .A2(n4295), .ZN(n3972) );
  NAND2_X1 U4645 ( .A1(n4118), .A2(REG2_REG_31__SCAN_IN), .ZN(n3971) );
  OAI211_X1 U4646 ( .C1(n4298), .C2(n4139), .A(n3972), .B(n3971), .ZN(U3260)
         );
  INV_X1 U4647 ( .A(n3973), .ZN(n3983) );
  NAND2_X1 U4648 ( .A1(n3974), .A2(n4181), .ZN(n3975) );
  OAI211_X1 U4649 ( .C1(n3977), .C2(n4139), .A(n3976), .B(n3975), .ZN(n3981)
         );
  AOI22_X1 U4650 ( .A1(n3990), .A2(n4179), .B1(n4118), .B2(
        REG2_REG_29__SCAN_IN), .ZN(n3978) );
  OAI21_X1 U4651 ( .B1(n3979), .B2(n4185), .A(n3978), .ZN(n3980) );
  AOI21_X1 U4652 ( .B1(n3981), .B2(n4164), .A(n3980), .ZN(n3982) );
  OAI21_X1 U4653 ( .B1(n3983), .B2(n4167), .A(n3982), .ZN(U3354) );
  XNOR2_X1 U4654 ( .A(n3984), .B(n3985), .ZN(n4205) );
  INV_X1 U4655 ( .A(n4205), .ZN(n3998) );
  AOI21_X1 U4656 ( .B1(n3987), .B2(n3986), .A(n4070), .ZN(n4204) );
  INV_X1 U4657 ( .A(n4009), .ZN(n3989) );
  OAI21_X1 U4658 ( .B1(n3989), .B2(n3994), .A(n3988), .ZN(n4305) );
  NOR2_X1 U4659 ( .A1(n4305), .A2(n4139), .ZN(n3996) );
  AOI22_X1 U4660 ( .A1(n3990), .A2(n4178), .B1(n4179), .B2(n4200), .ZN(n3993)
         );
  AOI22_X1 U4661 ( .A1(n3991), .A2(n4181), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4360), .ZN(n3992) );
  OAI211_X1 U4662 ( .C1(n3994), .C2(n4185), .A(n3993), .B(n3992), .ZN(n3995)
         );
  AOI211_X1 U4663 ( .C1(n4204), .C2(n4164), .A(n3996), .B(n3995), .ZN(n3997)
         );
  OAI21_X1 U4664 ( .B1(n3998), .B2(n4167), .A(n3997), .ZN(U3263) );
  XNOR2_X1 U4665 ( .A(n3999), .B(n4002), .ZN(n4209) );
  INV_X1 U4666 ( .A(n4209), .ZN(n4015) );
  OAI21_X1 U4667 ( .B1(n2112), .B2(n4001), .A(n4000), .ZN(n4004) );
  INV_X1 U4668 ( .A(n4002), .ZN(n4003) );
  XNOR2_X1 U4669 ( .A(n4004), .B(n4003), .ZN(n4008) );
  OAI22_X1 U4670 ( .A1(n4005), .A2(n4273), .B1(n4066), .B2(n4010), .ZN(n4006)
         );
  AOI21_X1 U4671 ( .B1(n4240), .B2(n4038), .A(n4006), .ZN(n4007) );
  OAI21_X1 U4672 ( .B1(n4008), .B2(n4070), .A(n4007), .ZN(n4208) );
  OAI21_X1 U4673 ( .B1(n4023), .B2(n4010), .A(n4009), .ZN(n4309) );
  AOI22_X1 U4674 ( .A1(n4011), .A2(n4181), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4360), .ZN(n4012) );
  OAI21_X1 U4675 ( .B1(n4309), .B2(n4139), .A(n4012), .ZN(n4013) );
  AOI21_X1 U4676 ( .B1(n4208), .B2(n4164), .A(n4013), .ZN(n4014) );
  OAI21_X1 U4677 ( .B1(n4015), .B2(n4167), .A(n4014), .ZN(U3264) );
  NAND2_X1 U4678 ( .A1(n4017), .A2(n4016), .ZN(n4018) );
  XNOR2_X1 U4679 ( .A(n4018), .B(n4020), .ZN(n4019) );
  NAND2_X1 U4680 ( .A1(n4019), .A2(n4169), .ZN(n4215) );
  XNOR2_X1 U4681 ( .A(n4021), .B(n4020), .ZN(n4218) );
  NAND2_X1 U4682 ( .A1(n4218), .A2(n4173), .ZN(n4031) );
  NOR2_X1 U4683 ( .A1(n4036), .A2(n4027), .ZN(n4022) );
  OR2_X1 U4684 ( .A1(n4023), .A2(n4022), .ZN(n4313) );
  INV_X1 U4685 ( .A(n4313), .ZN(n4029) );
  AOI22_X1 U4686 ( .A1(n4200), .A2(n4178), .B1(n4179), .B2(n4213), .ZN(n4026)
         );
  AOI22_X1 U4687 ( .A1(n4024), .A2(n4181), .B1(n4118), .B2(
        REG2_REG_25__SCAN_IN), .ZN(n4025) );
  OAI211_X1 U4688 ( .C1(n4027), .C2(n4185), .A(n4026), .B(n4025), .ZN(n4028)
         );
  AOI21_X1 U4689 ( .B1(n4029), .B2(n4473), .A(n4028), .ZN(n4030) );
  OAI211_X1 U4690 ( .C1(n4118), .C2(n4215), .A(n4031), .B(n4030), .ZN(U3265)
         );
  XOR2_X1 U4691 ( .A(n4035), .B(n4032), .Z(n4033) );
  NAND2_X1 U4692 ( .A1(n4033), .A2(n4169), .ZN(n4224) );
  XNOR2_X1 U4693 ( .A(n4034), .B(n4035), .ZN(n4227) );
  NAND2_X1 U4694 ( .A1(n4227), .A2(n4173), .ZN(n4046) );
  AND2_X1 U4695 ( .A1(n2050), .A2(n4221), .ZN(n4037) );
  OR2_X1 U4696 ( .A1(n4037), .A2(n4036), .ZN(n4317) );
  INV_X1 U4697 ( .A(n4317), .ZN(n4044) );
  AOI22_X1 U4698 ( .A1(n4038), .A2(n4178), .B1(n4179), .B2(n4222), .ZN(n4041)
         );
  AOI22_X1 U4699 ( .A1(REG2_REG_24__SCAN_IN), .A2(n4118), .B1(n4039), .B2(
        n4181), .ZN(n4040) );
  OAI211_X1 U4700 ( .C1(n4042), .C2(n4185), .A(n4041), .B(n4040), .ZN(n4043)
         );
  AOI21_X1 U4701 ( .B1(n4044), .B2(n4473), .A(n4043), .ZN(n4045) );
  OAI211_X1 U4702 ( .C1(n4118), .C2(n4224), .A(n4046), .B(n4045), .ZN(U3266)
         );
  XOR2_X1 U4703 ( .A(n4052), .B(n4047), .Z(n4231) );
  INV_X1 U4704 ( .A(n4231), .ZN(n4064) );
  INV_X1 U4705 ( .A(n4048), .ZN(n4050) );
  AOI21_X1 U4706 ( .B1(n4084), .B2(n4050), .A(n4049), .ZN(n4065) );
  OAI21_X1 U4707 ( .B1(n4065), .B2(n4077), .A(n4051), .ZN(n4053) );
  XNOR2_X1 U4708 ( .A(n4053), .B(n4052), .ZN(n4057) );
  OAI22_X1 U4709 ( .A1(n4054), .A2(n4273), .B1(n4058), .B2(n4066), .ZN(n4055)
         );
  AOI21_X1 U4710 ( .B1(n4240), .B2(n4090), .A(n4055), .ZN(n4056) );
  OAI21_X1 U4711 ( .B1(n4057), .B2(n4070), .A(n4056), .ZN(n4230) );
  OAI21_X1 U4712 ( .B1(n2128), .B2(n4058), .A(n2050), .ZN(n4321) );
  INV_X1 U4713 ( .A(n4059), .ZN(n4060) );
  AOI22_X1 U4714 ( .A1(n4118), .A2(REG2_REG_23__SCAN_IN), .B1(n4060), .B2(
        n4181), .ZN(n4061) );
  OAI21_X1 U4715 ( .B1(n4321), .B2(n4139), .A(n4061), .ZN(n4062) );
  AOI21_X1 U4716 ( .B1(n4230), .B2(n4164), .A(n4062), .ZN(n4063) );
  OAI21_X1 U4717 ( .B1(n4064), .B2(n4167), .A(n4063), .ZN(U3267) );
  XOR2_X1 U4718 ( .A(n4077), .B(n4065), .Z(n4071) );
  OAI22_X1 U4719 ( .A1(n4067), .A2(n4288), .B1(n4072), .B2(n4066), .ZN(n4068)
         );
  AOI21_X1 U4720 ( .B1(n4284), .B2(n4222), .A(n4068), .ZN(n4069) );
  OAI21_X1 U4721 ( .B1(n4071), .B2(n4070), .A(n4069), .ZN(n4235) );
  OR2_X1 U4722 ( .A1(n4088), .A2(n4072), .ZN(n4073) );
  NAND2_X1 U4723 ( .A1(n4074), .A2(n4073), .ZN(n4325) );
  AOI22_X1 U4724 ( .A1(n4118), .A2(REG2_REG_22__SCAN_IN), .B1(n4075), .B2(
        n4181), .ZN(n4076) );
  OAI21_X1 U4725 ( .B1(n4325), .B2(n4139), .A(n4076), .ZN(n4082) );
  NOR2_X1 U4726 ( .A1(n4078), .A2(n4077), .ZN(n4234) );
  INV_X1 U4727 ( .A(n4079), .ZN(n4080) );
  NOR3_X1 U4728 ( .A1(n4234), .A2(n4080), .A3(n4167), .ZN(n4081) );
  AOI211_X1 U4729 ( .C1(n4164), .C2(n4235), .A(n4082), .B(n4081), .ZN(n4083)
         );
  INV_X1 U4730 ( .A(n4083), .ZN(U3268) );
  XNOR2_X1 U4731 ( .A(n4084), .B(n4086), .ZN(n4085) );
  NAND2_X1 U4732 ( .A1(n4085), .A2(n4169), .ZN(n4243) );
  XNOR2_X1 U4733 ( .A(n4087), .B(n4086), .ZN(n4246) );
  NAND2_X1 U4734 ( .A1(n4246), .A2(n4173), .ZN(n4098) );
  INV_X1 U4735 ( .A(n4088), .ZN(n4089) );
  OAI21_X1 U4736 ( .B1(n4113), .B2(n4094), .A(n4089), .ZN(n4329) );
  INV_X1 U4737 ( .A(n4329), .ZN(n4096) );
  AOI22_X1 U4738 ( .A1(n4179), .A2(n4241), .B1(n4178), .B2(n4090), .ZN(n4093)
         );
  AOI22_X1 U4739 ( .A1(n4118), .A2(REG2_REG_21__SCAN_IN), .B1(n4091), .B2(
        n4181), .ZN(n4092) );
  OAI211_X1 U4740 ( .C1(n4094), .C2(n4185), .A(n4093), .B(n4092), .ZN(n4095)
         );
  AOI21_X1 U4741 ( .B1(n4096), .B2(n4473), .A(n4095), .ZN(n4097) );
  OAI211_X1 U4742 ( .C1(n4118), .C2(n4243), .A(n4098), .B(n4097), .ZN(U3269)
         );
  XNOR2_X1 U4743 ( .A(n4099), .B(n4103), .ZN(n4112) );
  INV_X1 U4744 ( .A(n4100), .ZN(n4101) );
  NAND2_X1 U4745 ( .A1(n4102), .A2(n4101), .ZN(n4104) );
  XNOR2_X1 U4746 ( .A(n4104), .B(n4103), .ZN(n4109) );
  AOI22_X1 U4747 ( .A1(n4106), .A2(n4284), .B1(n4282), .B2(n4105), .ZN(n4107)
         );
  OAI21_X1 U4748 ( .B1(n4155), .B2(n4288), .A(n4107), .ZN(n4108) );
  AOI21_X1 U4749 ( .B1(n4109), .B2(n4169), .A(n4108), .ZN(n4110) );
  OAI21_X1 U4750 ( .B1(n4112), .B2(n4111), .A(n4110), .ZN(n4249) );
  INV_X1 U4751 ( .A(n4249), .ZN(n4122) );
  INV_X1 U4752 ( .A(n4112), .ZN(n4250) );
  INV_X1 U4753 ( .A(n4136), .ZN(n4116) );
  INV_X1 U4754 ( .A(n4113), .ZN(n4114) );
  OAI21_X1 U4755 ( .B1(n4116), .B2(n4115), .A(n4114), .ZN(n4333) );
  AOI22_X1 U4756 ( .A1(n4118), .A2(REG2_REG_20__SCAN_IN), .B1(n4117), .B2(
        n4181), .ZN(n4119) );
  OAI21_X1 U4757 ( .B1(n4333), .B2(n4139), .A(n4119), .ZN(n4120) );
  AOI21_X1 U4758 ( .B1(n4250), .B2(n4474), .A(n4120), .ZN(n4121) );
  OAI21_X1 U4759 ( .B1(n4122), .B2(n4360), .A(n4121), .ZN(U3270) );
  XNOR2_X1 U4760 ( .A(n4123), .B(n4129), .ZN(n4254) );
  INV_X1 U4761 ( .A(n4254), .ZN(n4146) );
  NAND2_X1 U4762 ( .A1(n4125), .A2(n4124), .ZN(n4150) );
  INV_X1 U4763 ( .A(n4126), .ZN(n4128) );
  OAI21_X1 U4764 ( .B1(n4150), .B2(n4128), .A(n4127), .ZN(n4130) );
  XNOR2_X1 U4765 ( .A(n4130), .B(n4129), .ZN(n4131) );
  NAND2_X1 U4766 ( .A1(n4131), .A2(n4169), .ZN(n4134) );
  AOI22_X1 U4767 ( .A1(n4261), .A2(n4240), .B1(n4282), .B2(n4132), .ZN(n4133)
         );
  OAI211_X1 U4768 ( .C1(n4135), .C2(n4273), .A(n4134), .B(n4133), .ZN(n4253)
         );
  INV_X1 U4769 ( .A(n4158), .ZN(n4138) );
  OAI21_X1 U4770 ( .B1(n4138), .B2(n4137), .A(n4136), .ZN(n4337) );
  NOR2_X1 U4771 ( .A1(n4337), .A2(n4139), .ZN(n4144) );
  INV_X1 U4772 ( .A(n4140), .ZN(n4141) );
  OAI22_X1 U4773 ( .A1(n4164), .A2(n4142), .B1(n4141), .B2(n4468), .ZN(n4143)
         );
  AOI211_X1 U4774 ( .C1(n4253), .C2(n4164), .A(n4144), .B(n4143), .ZN(n4145)
         );
  OAI21_X1 U4775 ( .B1(n4146), .B2(n4167), .A(n4145), .ZN(U3271) );
  OAI21_X1 U4776 ( .B1(n4148), .B2(n4151), .A(n4147), .ZN(n4149) );
  INV_X1 U4777 ( .A(n4149), .ZN(n4259) );
  XOR2_X1 U4778 ( .A(n4151), .B(n4150), .Z(n4157) );
  AOI22_X1 U4779 ( .A1(n4153), .A2(n4240), .B1(n4152), .B2(n4282), .ZN(n4154)
         );
  OAI21_X1 U4780 ( .B1(n4155), .B2(n4273), .A(n4154), .ZN(n4156) );
  AOI21_X1 U4781 ( .B1(n4157), .B2(n4169), .A(n4156), .ZN(n4258) );
  INV_X1 U4782 ( .A(n4258), .ZN(n4165) );
  OAI211_X1 U4783 ( .C1(n4175), .C2(n4159), .A(n4158), .B(n4276), .ZN(n4257)
         );
  NOR2_X1 U4784 ( .A1(n4257), .A2(n4160), .ZN(n4163) );
  OAI22_X1 U4785 ( .A1(n4164), .A2(n3916), .B1(n4161), .B2(n4468), .ZN(n4162)
         );
  AOI211_X1 U4786 ( .C1(n4165), .C2(n4164), .A(n4163), .B(n4162), .ZN(n4166)
         );
  OAI21_X1 U4787 ( .B1(n4259), .B2(n4167), .A(n4166), .ZN(U3272) );
  XNOR2_X1 U4788 ( .A(n4168), .B(n4172), .ZN(n4170) );
  NAND2_X1 U4789 ( .A1(n4170), .A2(n4169), .ZN(n4263) );
  XOR2_X1 U4790 ( .A(n4172), .B(n4171), .Z(n4266) );
  NAND2_X1 U4791 ( .A1(n4266), .A2(n4173), .ZN(n4190) );
  INV_X1 U4792 ( .A(n4174), .ZN(n4177) );
  INV_X1 U4793 ( .A(n4175), .ZN(n4176) );
  OAI21_X1 U4794 ( .B1(n4177), .B2(n4186), .A(n4176), .ZN(n4342) );
  INV_X1 U4795 ( .A(n4342), .ZN(n4188) );
  AOI22_X1 U4796 ( .A1(n4179), .A2(n4285), .B1(n4178), .B2(n4261), .ZN(n4184)
         );
  INV_X1 U4797 ( .A(n4180), .ZN(n4182) );
  AOI22_X1 U4798 ( .A1(n4118), .A2(REG2_REG_17__SCAN_IN), .B1(n4182), .B2(
        n4181), .ZN(n4183) );
  OAI211_X1 U4799 ( .C1(n4186), .C2(n4185), .A(n4184), .B(n4183), .ZN(n4187)
         );
  AOI21_X1 U4800 ( .B1(n4188), .B2(n4473), .A(n4187), .ZN(n4189) );
  OAI211_X1 U4801 ( .C1(n4118), .C2(n4263), .A(n4190), .B(n4189), .ZN(U3273)
         );
  NOR2_X1 U4802 ( .A1(n4517), .A2(n4191), .ZN(n4192) );
  AOI21_X1 U4803 ( .B1(n4517), .B2(n4295), .A(n4192), .ZN(n4193) );
  OAI21_X1 U4804 ( .B1(n4298), .B2(n4294), .A(n4193), .ZN(U3549) );
  INV_X1 U4805 ( .A(n4361), .ZN(n4301) );
  INV_X1 U4806 ( .A(n4195), .ZN(n4196) );
  AOI21_X1 U4807 ( .B1(n4197), .B2(n4282), .A(n4196), .ZN(n4363) );
  MUX2_X1 U4808 ( .A(n4363), .B(n2729), .S(n4515), .Z(n4198) );
  OAI21_X1 U4809 ( .B1(n4301), .B2(n4294), .A(n4198), .ZN(U3548) );
  AOI22_X1 U4810 ( .A1(n4200), .A2(n4240), .B1(n4199), .B2(n4282), .ZN(n4201)
         );
  OAI21_X1 U4811 ( .B1(n4202), .B2(n4273), .A(n4201), .ZN(n4203) );
  AOI211_X1 U4812 ( .C1(n4205), .C2(n4504), .A(n4204), .B(n4203), .ZN(n4302)
         );
  MUX2_X1 U4813 ( .A(n4206), .B(n4302), .S(n4517), .Z(n4207) );
  AOI21_X1 U4814 ( .B1(n4209), .B2(n4504), .A(n4208), .ZN(n4306) );
  MUX2_X1 U4815 ( .A(n4210), .B(n4306), .S(n4517), .Z(n4211) );
  OAI21_X1 U4816 ( .B1(n4294), .B2(n4309), .A(n4211), .ZN(U3544) );
  AOI22_X1 U4817 ( .A1(n4213), .A2(n4240), .B1(n4212), .B2(n4282), .ZN(n4214)
         );
  OAI211_X1 U4818 ( .C1(n4216), .C2(n4273), .A(n4215), .B(n4214), .ZN(n4217)
         );
  AOI21_X1 U4819 ( .B1(n4218), .B2(n4504), .A(n4217), .ZN(n4310) );
  MUX2_X1 U4820 ( .A(n4219), .B(n4310), .S(n4517), .Z(n4220) );
  OAI21_X1 U4821 ( .B1(n4294), .B2(n4313), .A(n4220), .ZN(U3543) );
  AOI22_X1 U4822 ( .A1(n4222), .A2(n4240), .B1(n4282), .B2(n4221), .ZN(n4223)
         );
  OAI211_X1 U4823 ( .C1(n4225), .C2(n4273), .A(n4224), .B(n4223), .ZN(n4226)
         );
  AOI21_X1 U4824 ( .B1(n4227), .B2(n4504), .A(n4226), .ZN(n4314) );
  MUX2_X1 U4825 ( .A(n4228), .B(n4314), .S(n4517), .Z(n4229) );
  OAI21_X1 U4826 ( .B1(n4294), .B2(n4317), .A(n4229), .ZN(U3542) );
  AOI21_X1 U4827 ( .B1(n4231), .B2(n4504), .A(n4230), .ZN(n4318) );
  MUX2_X1 U4828 ( .A(n4232), .B(n4318), .S(n4517), .Z(n4233) );
  OAI21_X1 U4829 ( .B1(n4294), .B2(n4321), .A(n4233), .ZN(U3541) );
  NOR2_X1 U4830 ( .A1(n4234), .A2(n4280), .ZN(n4236) );
  AOI21_X1 U4831 ( .B1(n4236), .B2(n4079), .A(n4235), .ZN(n4322) );
  MUX2_X1 U4832 ( .A(n4237), .B(n4322), .S(n4517), .Z(n4238) );
  OAI21_X1 U4833 ( .B1(n4294), .B2(n4325), .A(n4238), .ZN(U3540) );
  AOI22_X1 U4834 ( .A1(n4241), .A2(n4240), .B1(n4239), .B2(n4282), .ZN(n4242)
         );
  OAI211_X1 U4835 ( .C1(n4244), .C2(n4273), .A(n4243), .B(n4242), .ZN(n4245)
         );
  AOI21_X1 U4836 ( .B1(n4246), .B2(n4504), .A(n4245), .ZN(n4326) );
  MUX2_X1 U4837 ( .A(n4247), .B(n4326), .S(n4517), .Z(n4248) );
  OAI21_X1 U4838 ( .B1(n4294), .B2(n4329), .A(n4248), .ZN(U3539) );
  AOI21_X1 U4839 ( .B1(n4502), .B2(n4250), .A(n4249), .ZN(n4330) );
  MUX2_X1 U4840 ( .A(n4251), .B(n4330), .S(n4517), .Z(n4252) );
  OAI21_X1 U4841 ( .B1(n4294), .B2(n4333), .A(n4252), .ZN(U3538) );
  AOI21_X1 U4842 ( .B1(n4254), .B2(n4504), .A(n4253), .ZN(n4334) );
  MUX2_X1 U4843 ( .A(n4255), .B(n4334), .S(n4517), .Z(n4256) );
  OAI21_X1 U4844 ( .B1(n4294), .B2(n4337), .A(n4256), .ZN(U3537) );
  OAI211_X1 U4845 ( .C1(n4259), .C2(n4280), .A(n4258), .B(n4257), .ZN(n4338)
         );
  MUX2_X1 U4846 ( .A(REG1_REG_18__SCAN_IN), .B(n4338), .S(n4517), .Z(U3536) );
  AOI22_X1 U4847 ( .A1(n4261), .A2(n4284), .B1(n4282), .B2(n4260), .ZN(n4262)
         );
  OAI211_X1 U4848 ( .C1(n4264), .C2(n4288), .A(n4263), .B(n4262), .ZN(n4265)
         );
  AOI21_X1 U4849 ( .B1(n4266), .B2(n4504), .A(n4265), .ZN(n4339) );
  MUX2_X1 U4850 ( .A(n4267), .B(n4339), .S(n4517), .Z(n4268) );
  OAI21_X1 U4851 ( .B1(n4294), .B2(n4342), .A(n4268), .ZN(U3535) );
  OR2_X1 U4852 ( .A1(n4269), .A2(n4288), .ZN(n4272) );
  NAND2_X1 U4853 ( .A1(n4270), .A2(n4282), .ZN(n4271) );
  OAI211_X1 U4854 ( .C1(n4274), .C2(n4273), .A(n4272), .B(n4271), .ZN(n4275)
         );
  AOI21_X1 U4855 ( .B1(n4277), .B2(n4276), .A(n4275), .ZN(n4279) );
  OAI211_X1 U4856 ( .C1(n4281), .C2(n4280), .A(n4279), .B(n4278), .ZN(n4343)
         );
  MUX2_X1 U4857 ( .A(REG1_REG_16__SCAN_IN), .B(n4343), .S(n4517), .Z(U3534) );
  AOI22_X1 U4858 ( .A1(n4285), .A2(n4284), .B1(n4283), .B2(n4282), .ZN(n4286)
         );
  OAI211_X1 U4859 ( .C1(n4289), .C2(n4288), .A(n4287), .B(n4286), .ZN(n4290)
         );
  AOI21_X1 U4860 ( .B1(n4291), .B2(n4504), .A(n4290), .ZN(n4344) );
  MUX2_X1 U4861 ( .A(n4292), .B(n4344), .S(n4517), .Z(n4293) );
  OAI21_X1 U4862 ( .B1(n4294), .B2(n4348), .A(n4293), .ZN(U3533) );
  NAND2_X1 U4863 ( .A1(n4512), .A2(n4295), .ZN(n4297) );
  NAND2_X1 U4864 ( .A1(n4510), .A2(REG0_REG_31__SCAN_IN), .ZN(n4296) );
  OAI211_X1 U4865 ( .C1(n4298), .C2(n4347), .A(n4297), .B(n4296), .ZN(U3517)
         );
  INV_X1 U4866 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4299) );
  MUX2_X1 U4867 ( .A(n4363), .B(n4299), .S(n4510), .Z(n4300) );
  OAI21_X1 U4868 ( .B1(n4301), .B2(n4347), .A(n4300), .ZN(U3516) );
  INV_X1 U4869 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4303) );
  MUX2_X1 U4870 ( .A(n4303), .B(n4302), .S(n4512), .Z(n4304) );
  INV_X1 U4871 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4307) );
  MUX2_X1 U4872 ( .A(n4307), .B(n4306), .S(n4512), .Z(n4308) );
  OAI21_X1 U4873 ( .B1(n4309), .B2(n4347), .A(n4308), .ZN(U3512) );
  INV_X1 U4874 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4311) );
  MUX2_X1 U4875 ( .A(n4311), .B(n4310), .S(n4512), .Z(n4312) );
  OAI21_X1 U4876 ( .B1(n4313), .B2(n4347), .A(n4312), .ZN(U3511) );
  INV_X1 U4877 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4315) );
  MUX2_X1 U4878 ( .A(n4315), .B(n4314), .S(n4512), .Z(n4316) );
  OAI21_X1 U4879 ( .B1(n4317), .B2(n4347), .A(n4316), .ZN(U3510) );
  INV_X1 U4880 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4319) );
  MUX2_X1 U4881 ( .A(n4319), .B(n4318), .S(n4512), .Z(n4320) );
  OAI21_X1 U4882 ( .B1(n4321), .B2(n4347), .A(n4320), .ZN(U3509) );
  INV_X1 U4883 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4323) );
  MUX2_X1 U4884 ( .A(n4323), .B(n4322), .S(n4512), .Z(n4324) );
  OAI21_X1 U4885 ( .B1(n4325), .B2(n4347), .A(n4324), .ZN(U3508) );
  INV_X1 U4886 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4327) );
  MUX2_X1 U4887 ( .A(n4327), .B(n4326), .S(n4512), .Z(n4328) );
  OAI21_X1 U4888 ( .B1(n4329), .B2(n4347), .A(n4328), .ZN(U3507) );
  INV_X1 U4889 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4331) );
  MUX2_X1 U4890 ( .A(n4331), .B(n4330), .S(n4512), .Z(n4332) );
  OAI21_X1 U4891 ( .B1(n4333), .B2(n4347), .A(n4332), .ZN(U3506) );
  INV_X1 U4892 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4335) );
  MUX2_X1 U4893 ( .A(n4335), .B(n4334), .S(n4512), .Z(n4336) );
  OAI21_X1 U4894 ( .B1(n4337), .B2(n4347), .A(n4336), .ZN(U3505) );
  MUX2_X1 U4895 ( .A(REG0_REG_18__SCAN_IN), .B(n4338), .S(n4512), .Z(U3503) );
  MUX2_X1 U4896 ( .A(n4340), .B(n4339), .S(n4512), .Z(n4341) );
  OAI21_X1 U4897 ( .B1(n4342), .B2(n4347), .A(n4341), .ZN(U3501) );
  MUX2_X1 U4898 ( .A(REG0_REG_16__SCAN_IN), .B(n4343), .S(n4512), .Z(U3499) );
  INV_X1 U4899 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4345) );
  MUX2_X1 U4900 ( .A(n4345), .B(n4344), .S(n4512), .Z(n4346) );
  OAI21_X1 U4901 ( .B1(n4348), .B2(n4347), .A(n4346), .ZN(U3497) );
  MUX2_X1 U4902 ( .A(DATAI_30_), .B(n4349), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4903 ( .A(DATAI_29_), .B(n4350), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U4904 ( .A(DATAI_21_), .B(n4351), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U4905 ( .A(n4352), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4906 ( .A(DATAI_8_), .B(n2121), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4907 ( .A(n4354), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4908 ( .A(n4355), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4909 ( .A(n4356), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4910 ( .A(DATAI_4_), .B(n4357), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4911 ( .A(n4358), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4912 ( .A(n2048), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  AOI22_X1 U4913 ( .A1(n4361), .A2(n4473), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4360), .ZN(n4362) );
  OAI21_X1 U4914 ( .B1(n4118), .B2(n4363), .A(n4362), .ZN(U3261) );
  OAI211_X1 U4915 ( .C1(n4366), .C2(n4365), .A(n4462), .B(n4364), .ZN(n4371)
         );
  OAI211_X1 U4916 ( .C1(n4369), .C2(n4368), .A(n4406), .B(n4367), .ZN(n4370)
         );
  OAI211_X1 U4917 ( .C1(n4467), .C2(n4493), .A(n4371), .B(n4370), .ZN(n4372)
         );
  AOI211_X1 U4918 ( .C1(n4460), .C2(ADDR_REG_9__SCAN_IN), .A(n4373), .B(n4372), 
        .ZN(n4374) );
  INV_X1 U4919 ( .A(n4374), .ZN(U3249) );
  OAI211_X1 U4920 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4376), .A(n4406), .B(n4375), .ZN(n4378) );
  NAND2_X1 U4921 ( .A1(n4378), .A2(n4377), .ZN(n4379) );
  AOI21_X1 U4922 ( .B1(n4460), .B2(ADDR_REG_10__SCAN_IN), .A(n4379), .ZN(n4383) );
  OAI211_X1 U4923 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4381), .A(n4462), .B(n4380), .ZN(n4382) );
  OAI211_X1 U4924 ( .C1(n4467), .C2(n4492), .A(n4383), .B(n4382), .ZN(U3250)
         );
  OAI211_X1 U4925 ( .C1(n4386), .C2(n4385), .A(n4462), .B(n4384), .ZN(n4391)
         );
  OAI211_X1 U4926 ( .C1(n4389), .C2(n4388), .A(n4406), .B(n4387), .ZN(n4390)
         );
  OAI211_X1 U4927 ( .C1(n4467), .C2(n4491), .A(n4391), .B(n4390), .ZN(n4392)
         );
  AOI211_X1 U4928 ( .C1(n4460), .C2(ADDR_REG_11__SCAN_IN), .A(n4393), .B(n4392), .ZN(n4394) );
  INV_X1 U4929 ( .A(n4394), .ZN(U3251) );
  OAI211_X1 U4930 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4396), .A(n4406), .B(n4395), .ZN(n4398) );
  NAND2_X1 U4931 ( .A1(n4398), .A2(n4397), .ZN(n4399) );
  AOI21_X1 U4932 ( .B1(n4460), .B2(ADDR_REG_12__SCAN_IN), .A(n4399), .ZN(n4403) );
  OAI211_X1 U4933 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4401), .A(n4462), .B(n4400), .ZN(n4402) );
  OAI211_X1 U4934 ( .C1(n4467), .C2(n4490), .A(n4403), .B(n4402), .ZN(U3252)
         );
  AOI21_X1 U4935 ( .B1(n4405), .B2(n4417), .A(n4404), .ZN(n4409) );
  OAI21_X1 U4936 ( .B1(n4409), .B2(n4408), .A(n4406), .ZN(n4407) );
  AOI21_X1 U4937 ( .B1(n4409), .B2(n4408), .A(n4407), .ZN(n4411) );
  AOI211_X1 U4938 ( .C1(n4460), .C2(ADDR_REG_13__SCAN_IN), .A(n4411), .B(n4410), .ZN(n4416) );
  OAI211_X1 U4939 ( .C1(n4414), .C2(n4413), .A(n4462), .B(n4412), .ZN(n4415)
         );
  OAI211_X1 U4940 ( .C1(n4467), .C2(n4417), .A(n4416), .B(n4415), .ZN(U3253)
         );
  AOI211_X1 U4941 ( .C1(n2341), .C2(n4419), .A(n4418), .B(n4456), .ZN(n4420)
         );
  AOI211_X1 U4942 ( .C1(n4460), .C2(ADDR_REG_14__SCAN_IN), .A(n4421), .B(n4420), .ZN(n4425) );
  OAI211_X1 U4943 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4423), .A(n4462), .B(n4422), .ZN(n4424) );
  OAI211_X1 U4944 ( .C1(n4467), .C2(n4487), .A(n4425), .B(n4424), .ZN(U3254)
         );
  AOI211_X1 U4945 ( .C1(n4428), .C2(n4427), .A(n4426), .B(n4456), .ZN(n4429)
         );
  AOI211_X1 U4946 ( .C1(n4460), .C2(ADDR_REG_15__SCAN_IN), .A(n4430), .B(n4429), .ZN(n4435) );
  OAI211_X1 U4947 ( .C1(n4433), .C2(n4432), .A(n4462), .B(n4431), .ZN(n4434)
         );
  OAI211_X1 U4948 ( .C1(n4467), .C2(n4436), .A(n4435), .B(n4434), .ZN(U3255)
         );
  INV_X1 U4949 ( .A(n4437), .ZN(n4441) );
  AOI221_X1 U4950 ( .B1(n4439), .B2(n4438), .C1(n2530), .C2(n4438), .A(n4456), 
        .ZN(n4440) );
  AOI211_X1 U4951 ( .C1(n4460), .C2(ADDR_REG_16__SCAN_IN), .A(n4441), .B(n4440), .ZN(n4445) );
  OAI221_X1 U4952 ( .B1(n4443), .B2(REG1_REG_16__SCAN_IN), .C1(n4443), .C2(
        n4442), .A(n4462), .ZN(n4444) );
  OAI211_X1 U4953 ( .C1(n4467), .C2(n4484), .A(n4445), .B(n4444), .ZN(U3256)
         );
  AOI221_X1 U4954 ( .B1(n4448), .B2(n4447), .C1(n4446), .C2(n4447), .A(n4456), 
        .ZN(n4449) );
  AOI211_X1 U4955 ( .C1(n4460), .C2(ADDR_REG_17__SCAN_IN), .A(n4450), .B(n4449), .ZN(n4455) );
  OAI221_X1 U4956 ( .B1(n4453), .B2(n4452), .C1(n4453), .C2(n4451), .A(n4462), 
        .ZN(n4454) );
  OAI211_X1 U4957 ( .C1(n4467), .C2(n4483), .A(n4455), .B(n4454), .ZN(U3257)
         );
  OAI211_X1 U4958 ( .C1(n4464), .C2(n4463), .A(n4462), .B(n4461), .ZN(n4465)
         );
  OAI211_X1 U4959 ( .C1(n4467), .C2(n4482), .A(n4466), .B(n4465), .ZN(U3258)
         );
  OAI22_X1 U4960 ( .A1(n4164), .A2(n4470), .B1(n4469), .B2(n4468), .ZN(n4471)
         );
  INV_X1 U4961 ( .A(n4471), .ZN(n4477) );
  AOI22_X1 U4962 ( .A1(n4475), .A2(n4474), .B1(n4473), .B2(n4472), .ZN(n4476)
         );
  OAI211_X1 U4963 ( .C1(n4118), .C2(n4478), .A(n4477), .B(n4476), .ZN(U3282)
         );
  AND2_X1 U4964 ( .A1(D_REG_31__SCAN_IN), .A2(n4479), .ZN(U3291) );
  AND2_X1 U4965 ( .A1(D_REG_30__SCAN_IN), .A2(n4479), .ZN(U3292) );
  AND2_X1 U4966 ( .A1(D_REG_29__SCAN_IN), .A2(n4479), .ZN(U3293) );
  AND2_X1 U4967 ( .A1(D_REG_28__SCAN_IN), .A2(n4479), .ZN(U3294) );
  AND2_X1 U4968 ( .A1(D_REG_27__SCAN_IN), .A2(n4479), .ZN(U3295) );
  AND2_X1 U4969 ( .A1(D_REG_26__SCAN_IN), .A2(n4479), .ZN(U3296) );
  AND2_X1 U4970 ( .A1(D_REG_25__SCAN_IN), .A2(n4479), .ZN(U3297) );
  AND2_X1 U4971 ( .A1(D_REG_24__SCAN_IN), .A2(n4479), .ZN(U3298) );
  AND2_X1 U4972 ( .A1(D_REG_23__SCAN_IN), .A2(n4479), .ZN(U3299) );
  AND2_X1 U4973 ( .A1(D_REG_22__SCAN_IN), .A2(n4479), .ZN(U3300) );
  AND2_X1 U4974 ( .A1(D_REG_21__SCAN_IN), .A2(n4479), .ZN(U3301) );
  AND2_X1 U4975 ( .A1(D_REG_20__SCAN_IN), .A2(n4479), .ZN(U3302) );
  AND2_X1 U4976 ( .A1(D_REG_19__SCAN_IN), .A2(n4479), .ZN(U3303) );
  AND2_X1 U4977 ( .A1(D_REG_18__SCAN_IN), .A2(n4479), .ZN(U3304) );
  AND2_X1 U4978 ( .A1(D_REG_17__SCAN_IN), .A2(n4479), .ZN(U3305) );
  AND2_X1 U4979 ( .A1(D_REG_16__SCAN_IN), .A2(n4479), .ZN(U3306) );
  AND2_X1 U4980 ( .A1(D_REG_15__SCAN_IN), .A2(n4479), .ZN(U3307) );
  AND2_X1 U4981 ( .A1(D_REG_14__SCAN_IN), .A2(n4479), .ZN(U3308) );
  AND2_X1 U4982 ( .A1(D_REG_13__SCAN_IN), .A2(n4479), .ZN(U3309) );
  AND2_X1 U4983 ( .A1(D_REG_12__SCAN_IN), .A2(n4479), .ZN(U3310) );
  AND2_X1 U4984 ( .A1(D_REG_11__SCAN_IN), .A2(n4479), .ZN(U3311) );
  AND2_X1 U4985 ( .A1(D_REG_10__SCAN_IN), .A2(n4479), .ZN(U3312) );
  AND2_X1 U4986 ( .A1(D_REG_9__SCAN_IN), .A2(n4479), .ZN(U3313) );
  AND2_X1 U4987 ( .A1(D_REG_8__SCAN_IN), .A2(n4479), .ZN(U3314) );
  AND2_X1 U4988 ( .A1(D_REG_7__SCAN_IN), .A2(n4479), .ZN(U3315) );
  AND2_X1 U4989 ( .A1(D_REG_6__SCAN_IN), .A2(n4479), .ZN(U3316) );
  AND2_X1 U4990 ( .A1(D_REG_5__SCAN_IN), .A2(n4479), .ZN(U3317) );
  AND2_X1 U4991 ( .A1(D_REG_4__SCAN_IN), .A2(n4479), .ZN(U3318) );
  AND2_X1 U4992 ( .A1(D_REG_3__SCAN_IN), .A2(n4479), .ZN(U3319) );
  AND2_X1 U4993 ( .A1(D_REG_2__SCAN_IN), .A2(n4479), .ZN(U3320) );
  OAI21_X1 U4994 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4480), .ZN(
        n4481) );
  INV_X1 U4995 ( .A(n4481), .ZN(U3329) );
  AOI22_X1 U4996 ( .A1(STATE_REG_SCAN_IN), .A2(n4482), .B1(n4632), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U4997 ( .A1(STATE_REG_SCAN_IN), .A2(n4483), .B1(n2553), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U4998 ( .A(DATAI_16_), .ZN(n4642) );
  AOI22_X1 U4999 ( .A1(STATE_REG_SCAN_IN), .A2(n4484), .B1(n4642), .B2(U3149), 
        .ZN(U3336) );
  OAI22_X1 U5000 ( .A1(U3149), .A2(n4485), .B1(DATAI_15_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4486) );
  INV_X1 U5001 ( .A(n4486), .ZN(U3337) );
  INV_X1 U5002 ( .A(DATAI_14_), .ZN(n4615) );
  AOI22_X1 U5003 ( .A1(STATE_REG_SCAN_IN), .A2(n4487), .B1(n4615), .B2(U3149), 
        .ZN(U3338) );
  OAI22_X1 U5004 ( .A1(U3149), .A2(n4488), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4489) );
  INV_X1 U5005 ( .A(n4489), .ZN(U3339) );
  AOI22_X1 U5006 ( .A1(STATE_REG_SCAN_IN), .A2(n4490), .B1(n2501), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5007 ( .A(DATAI_11_), .ZN(n4539) );
  AOI22_X1 U5008 ( .A1(STATE_REG_SCAN_IN), .A2(n4491), .B1(n4539), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5009 ( .A(DATAI_10_), .ZN(n4529) );
  AOI22_X1 U5010 ( .A1(STATE_REG_SCAN_IN), .A2(n4492), .B1(n4529), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5011 ( .A(DATAI_9_), .ZN(n4605) );
  AOI22_X1 U5012 ( .A1(STATE_REG_SCAN_IN), .A2(n4493), .B1(n4605), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5013 ( .A(n4494), .ZN(n4497) );
  INV_X1 U5014 ( .A(n4495), .ZN(n4496) );
  AOI211_X1 U5015 ( .C1(n4502), .C2(n4498), .A(n4497), .B(n4496), .ZN(n4513)
         );
  AOI22_X1 U5016 ( .A1(n4512), .A2(n4513), .B1(n2356), .B2(n4510), .ZN(U3467)
         );
  INV_X1 U5017 ( .A(n4499), .ZN(n4501) );
  AOI211_X1 U5018 ( .C1(n4503), .C2(n4502), .A(n4501), .B(n4500), .ZN(n4514)
         );
  AOI22_X1 U5019 ( .A1(n4512), .A2(n4514), .B1(n2386), .B2(n4510), .ZN(U3475)
         );
  NAND3_X1 U5020 ( .A1(n4506), .A2(n4505), .A3(n4504), .ZN(n4507) );
  INV_X1 U5021 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4511) );
  AOI22_X1 U5022 ( .A1(n4512), .A2(n4516), .B1(n4511), .B2(n4510), .ZN(U3481)
         );
  AOI22_X1 U5023 ( .A1(n4517), .A2(n4513), .B1(n2357), .B2(n4515), .ZN(U3518)
         );
  AOI22_X1 U5024 ( .A1(n4517), .A2(n4514), .B1(n2385), .B2(n4515), .ZN(U3522)
         );
  AOI22_X1 U5025 ( .A1(n4517), .A2(n4516), .B1(n2428), .B2(n4515), .ZN(U3525)
         );
  AOI22_X1 U5026 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n4704) );
  AOI22_X1 U5027 ( .A1(n2453), .A2(keyinput_g51), .B1(keyinput_g23), .B2(n2446), .ZN(n4518) );
  OAI221_X1 U5028 ( .B1(n2453), .B2(keyinput_g51), .C1(n2446), .C2(
        keyinput_g23), .A(n4518), .ZN(n4527) );
  XNOR2_X1 U5029 ( .A(n4519), .B(keyinput_g61), .ZN(n4526) );
  XNOR2_X1 U5030 ( .A(keyinput_g19), .B(n2501), .ZN(n4525) );
  XNOR2_X1 U5031 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_g57), .ZN(n4523) );
  XNOR2_X1 U5032 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_g52), .ZN(n4522) );
  XNOR2_X1 U5033 ( .A(DATAI_0_), .B(keyinput_g31), .ZN(n4521) );
  XNOR2_X1 U5034 ( .A(DATAI_9_), .B(keyinput_g22), .ZN(n4520) );
  NAND4_X1 U5035 ( .A1(n4523), .A2(n4522), .A3(n4521), .A4(n4520), .ZN(n4524)
         );
  NOR4_X1 U5036 ( .A1(n4527), .A2(n4526), .A3(n4525), .A4(n4524), .ZN(n4565)
         );
  AOI22_X1 U5037 ( .A1(n2568), .A2(keyinput_g11), .B1(n4606), .B2(keyinput_g33), .ZN(n4528) );
  OAI221_X1 U5038 ( .B1(n2568), .B2(keyinput_g11), .C1(n4606), .C2(
        keyinput_g33), .A(n4528), .ZN(n4537) );
  XNOR2_X1 U5039 ( .A(keyinput_g21), .B(n4529), .ZN(n4536) );
  XNOR2_X1 U5040 ( .A(keyinput_g4), .B(n2615), .ZN(n4535) );
  XNOR2_X1 U5041 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_g56), .ZN(n4533) );
  XNOR2_X1 U5042 ( .A(DATAI_30_), .B(keyinput_g1), .ZN(n4532) );
  XNOR2_X1 U5043 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_g50), .ZN(n4531) );
  XNOR2_X1 U5044 ( .A(DATAI_3_), .B(keyinput_g28), .ZN(n4530) );
  NAND4_X1 U5045 ( .A1(n4533), .A2(n4532), .A3(n4531), .A4(n4530), .ZN(n4534)
         );
  NOR4_X1 U5046 ( .A1(n4537), .A2(n4536), .A3(n4535), .A4(n4534), .ZN(n4564)
         );
  INV_X1 U5047 ( .A(DATAI_4_), .ZN(n4633) );
  AOI22_X1 U5048 ( .A1(n4539), .A2(keyinput_g20), .B1(keyinput_g27), .B2(n4633), .ZN(n4538) );
  OAI221_X1 U5049 ( .B1(n4539), .B2(keyinput_g20), .C1(n4633), .C2(
        keyinput_g27), .A(n4538), .ZN(n4550) );
  AOI22_X1 U5050 ( .A1(n4542), .A2(keyinput_g7), .B1(n4541), .B2(keyinput_g45), 
        .ZN(n4540) );
  OAI221_X1 U5051 ( .B1(n4542), .B2(keyinput_g7), .C1(n4541), .C2(keyinput_g45), .A(n4540), .ZN(n4549) );
  AOI22_X1 U5052 ( .A1(n4544), .A2(keyinput_g12), .B1(n4635), .B2(keyinput_g49), .ZN(n4543) );
  OAI221_X1 U5053 ( .B1(n4544), .B2(keyinput_g12), .C1(n4635), .C2(
        keyinput_g49), .A(n4543), .ZN(n4548) );
  XNOR2_X1 U5054 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_g44), .ZN(n4546) );
  XNOR2_X1 U5055 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_g38), .ZN(n4545) );
  NAND2_X1 U5056 ( .A1(n4546), .A2(n4545), .ZN(n4547) );
  NOR4_X1 U5057 ( .A1(n4550), .A2(n4549), .A3(n4548), .A4(n4547), .ZN(n4563)
         );
  AOI22_X1 U5058 ( .A1(n4645), .A2(keyinput_g47), .B1(keyinput_g5), .B2(n4552), 
        .ZN(n4551) );
  OAI221_X1 U5059 ( .B1(n4645), .B2(keyinput_g47), .C1(n4552), .C2(keyinput_g5), .A(n4551), .ZN(n4561) );
  AOI22_X1 U5060 ( .A1(n4554), .A2(keyinput_g34), .B1(n3715), .B2(keyinput_g40), .ZN(n4553) );
  OAI221_X1 U5061 ( .B1(n4554), .B2(keyinput_g34), .C1(n3715), .C2(
        keyinput_g40), .A(n4553), .ZN(n4560) );
  XNOR2_X1 U5062 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_g43), .ZN(n4558) );
  XNOR2_X1 U5063 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_g58), .ZN(n4557) );
  XNOR2_X1 U5064 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_g55), .ZN(n4556) );
  XNOR2_X1 U5065 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_g35), .ZN(n4555) );
  NAND4_X1 U5066 ( .A1(n4558), .A2(n4557), .A3(n4556), .A4(n4555), .ZN(n4559)
         );
  NOR3_X1 U5067 ( .A1(n4561), .A2(n4560), .A3(n4559), .ZN(n4562) );
  NAND4_X1 U5068 ( .A1(n4565), .A2(n4564), .A3(n4563), .A4(n4562), .ZN(n4702)
         );
  AOI22_X1 U5069 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(DATAI_22_), .B2(
        keyinput_g9), .ZN(n4566) );
  OAI221_X1 U5070 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(DATAI_22_), .C2(
        keyinput_g9), .A(n4566), .ZN(n4573) );
  AOI22_X1 U5071 ( .A1(DATAI_23_), .A2(keyinput_g8), .B1(DATAI_25_), .B2(
        keyinput_g6), .ZN(n4567) );
  OAI221_X1 U5072 ( .B1(DATAI_23_), .B2(keyinput_g8), .C1(DATAI_25_), .C2(
        keyinput_g6), .A(n4567), .ZN(n4572) );
  AOI22_X1 U5073 ( .A1(DATAI_6_), .A2(keyinput_g25), .B1(DATAI_15_), .B2(
        keyinput_g16), .ZN(n4568) );
  OAI221_X1 U5074 ( .B1(DATAI_6_), .B2(keyinput_g25), .C1(DATAI_15_), .C2(
        keyinput_g16), .A(n4568), .ZN(n4571) );
  AOI22_X1 U5075 ( .A1(DATAI_18_), .A2(keyinput_g13), .B1(REG3_REG_1__SCAN_IN), 
        .B2(keyinput_g42), .ZN(n4569) );
  OAI221_X1 U5076 ( .B1(DATAI_18_), .B2(keyinput_g13), .C1(REG3_REG_1__SCAN_IN), .C2(keyinput_g42), .A(n4569), .ZN(n4570) );
  NOR4_X1 U5077 ( .A1(n4573), .A2(n4572), .A3(n4571), .A4(n4570), .ZN(n4600)
         );
  XOR2_X1 U5078 ( .A(U3149), .B(keyinput_g32), .Z(n4580) );
  AOI22_X1 U5079 ( .A1(DATAI_1_), .A2(keyinput_g30), .B1(n2553), .B2(
        keyinput_g14), .ZN(n4574) );
  OAI221_X1 U5080 ( .B1(DATAI_1_), .B2(keyinput_g30), .C1(n2553), .C2(
        keyinput_g14), .A(n4574), .ZN(n4579) );
  AOI22_X1 U5081 ( .A1(DATAI_28_), .A2(keyinput_g3), .B1(DATAI_29_), .B2(
        keyinput_g2), .ZN(n4575) );
  OAI221_X1 U5082 ( .B1(DATAI_28_), .B2(keyinput_g3), .C1(DATAI_29_), .C2(
        keyinput_g2), .A(n4575), .ZN(n4578) );
  AOI22_X1 U5083 ( .A1(DATAI_31_), .A2(keyinput_g0), .B1(REG3_REG_20__SCAN_IN), 
        .B2(keyinput_g53), .ZN(n4576) );
  OAI221_X1 U5084 ( .B1(DATAI_31_), .B2(keyinput_g0), .C1(REG3_REG_20__SCAN_IN), .C2(keyinput_g53), .A(n4576), .ZN(n4577) );
  NOR4_X1 U5085 ( .A1(n4580), .A2(n4579), .A3(n4578), .A4(n4577), .ZN(n4599)
         );
  AOI22_X1 U5086 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_g37), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .ZN(n4581) );
  OAI221_X1 U5087 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_g37), .C1(
        REG3_REG_16__SCAN_IN), .C2(keyinput_g46), .A(n4581), .ZN(n4588) );
  AOI22_X1 U5088 ( .A1(REG3_REG_17__SCAN_IN), .A2(keyinput_g48), .B1(
        REG3_REG_23__SCAN_IN), .B2(keyinput_g36), .ZN(n4582) );
  OAI221_X1 U5089 ( .B1(REG3_REG_17__SCAN_IN), .B2(keyinput_g48), .C1(
        REG3_REG_23__SCAN_IN), .C2(keyinput_g36), .A(n4582), .ZN(n4587) );
  AOI22_X1 U5090 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_g39), .B1(n2503), 
        .B2(keyinput_g54), .ZN(n4583) );
  OAI221_X1 U5091 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_g39), .C1(n2503), 
        .C2(keyinput_g54), .A(n4583), .ZN(n4586) );
  AOI22_X1 U5092 ( .A1(DATAI_16_), .A2(keyinput_g15), .B1(REG3_REG_8__SCAN_IN), 
        .B2(keyinput_g41), .ZN(n4584) );
  OAI221_X1 U5093 ( .B1(DATAI_16_), .B2(keyinput_g15), .C1(REG3_REG_8__SCAN_IN), .C2(keyinput_g41), .A(n4584), .ZN(n4585) );
  NOR4_X1 U5094 ( .A1(n4588), .A2(n4587), .A3(n4586), .A4(n4585), .ZN(n4598)
         );
  AOI22_X1 U5095 ( .A1(DATAI_13_), .A2(keyinput_g18), .B1(IR_REG_7__SCAN_IN), 
        .B2(keyinput_g62), .ZN(n4589) );
  OAI221_X1 U5096 ( .B1(DATAI_13_), .B2(keyinput_g18), .C1(IR_REG_7__SCAN_IN), 
        .C2(keyinput_g62), .A(n4589), .ZN(n4596) );
  AOI22_X1 U5097 ( .A1(DATAI_5_), .A2(keyinput_g26), .B1(DATAI_14_), .B2(
        keyinput_g17), .ZN(n4590) );
  OAI221_X1 U5098 ( .B1(DATAI_5_), .B2(keyinput_g26), .C1(DATAI_14_), .C2(
        keyinput_g17), .A(n4590), .ZN(n4595) );
  AOI22_X1 U5099 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput_g60), .B1(
        IR_REG_8__SCAN_IN), .B2(keyinput_g63), .ZN(n4591) );
  OAI221_X1 U5100 ( .B1(IR_REG_5__SCAN_IN), .B2(keyinput_g60), .C1(
        IR_REG_8__SCAN_IN), .C2(keyinput_g63), .A(n4591), .ZN(n4594) );
  AOI22_X1 U5101 ( .A1(DATAI_2_), .A2(keyinput_g29), .B1(IR_REG_4__SCAN_IN), 
        .B2(keyinput_g59), .ZN(n4592) );
  OAI221_X1 U5102 ( .B1(DATAI_2_), .B2(keyinput_g29), .C1(IR_REG_4__SCAN_IN), 
        .C2(keyinput_g59), .A(n4592), .ZN(n4593) );
  NOR4_X1 U5103 ( .A1(n4596), .A2(n4595), .A3(n4594), .A4(n4593), .ZN(n4597)
         );
  NAND4_X1 U5104 ( .A1(n4600), .A2(n4599), .A3(n4598), .A4(n4597), .ZN(n4701)
         );
  INV_X1 U5105 ( .A(DATAI_7_), .ZN(n4696) );
  INV_X1 U5106 ( .A(DATAI_21_), .ZN(n4602) );
  AOI22_X1 U5107 ( .A1(n4602), .A2(keyinput_f10), .B1(n2453), .B2(keyinput_f51), .ZN(n4601) );
  OAI221_X1 U5108 ( .B1(n4602), .B2(keyinput_f10), .C1(n2453), .C2(
        keyinput_f51), .A(n4601), .ZN(n4613) );
  AOI22_X1 U5109 ( .A1(n4605), .A2(keyinput_f22), .B1(n4604), .B2(keyinput_f6), 
        .ZN(n4603) );
  OAI221_X1 U5110 ( .B1(n4605), .B2(keyinput_f22), .C1(n4604), .C2(keyinput_f6), .A(n4603), .ZN(n4612) );
  XOR2_X1 U5111 ( .A(n4606), .B(keyinput_f33), .Z(n4610) );
  XNOR2_X1 U5112 ( .A(DATAI_0_), .B(keyinput_f31), .ZN(n4609) );
  XNOR2_X1 U5113 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n4608) );
  XNOR2_X1 U5114 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_f56), .ZN(n4607) );
  NAND4_X1 U5115 ( .A1(n4610), .A2(n4609), .A3(n4608), .A4(n4607), .ZN(n4611)
         );
  NOR3_X1 U5116 ( .A1(n4613), .A2(n4612), .A3(n4611), .ZN(n4656) );
  AOI22_X1 U5117 ( .A1(n4616), .A2(keyinput_f39), .B1(keyinput_f17), .B2(n4615), .ZN(n4614) );
  OAI221_X1 U5118 ( .B1(n4616), .B2(keyinput_f39), .C1(n4615), .C2(
        keyinput_f17), .A(n4614), .ZN(n4624) );
  XNOR2_X1 U5119 ( .A(keyinput_f54), .B(n2503), .ZN(n4623) );
  XNOR2_X1 U5120 ( .A(keyinput_f4), .B(n2615), .ZN(n4622) );
  XNOR2_X1 U5121 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_f62), .ZN(n4620) );
  XNOR2_X1 U5122 ( .A(DATAI_3_), .B(keyinput_f28), .ZN(n4619) );
  XNOR2_X1 U5123 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_f50), .ZN(n4618) );
  XNOR2_X1 U5124 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_f57), .ZN(n4617) );
  NAND4_X1 U5125 ( .A1(n4620), .A2(n4619), .A3(n4618), .A4(n4617), .ZN(n4621)
         );
  NOR4_X1 U5126 ( .A1(n4624), .A2(n4623), .A3(n4622), .A4(n4621), .ZN(n4655)
         );
  AOI22_X1 U5127 ( .A1(n4627), .A2(keyinput_f36), .B1(keyinput_f48), .B2(n4626), .ZN(n4625) );
  OAI221_X1 U5128 ( .B1(n4627), .B2(keyinput_f36), .C1(n4626), .C2(
        keyinput_f48), .A(n4625), .ZN(n4640) );
  INV_X1 U5129 ( .A(DATAI_2_), .ZN(n4629) );
  AOI22_X1 U5130 ( .A1(n4630), .A2(keyinput_f43), .B1(keyinput_f29), .B2(n4629), .ZN(n4628) );
  OAI221_X1 U5131 ( .B1(n4630), .B2(keyinput_f43), .C1(n4629), .C2(
        keyinput_f29), .A(n4628), .ZN(n4639) );
  AOI22_X1 U5132 ( .A1(n4633), .A2(keyinput_f27), .B1(keyinput_f13), .B2(n4632), .ZN(n4631) );
  OAI221_X1 U5133 ( .B1(n4633), .B2(keyinput_f27), .C1(n4632), .C2(
        keyinput_f13), .A(n4631), .ZN(n4638) );
  INV_X1 U5134 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5135 ( .A1(n4636), .A2(keyinput_f41), .B1(n4635), .B2(keyinput_f49), .ZN(n4634) );
  OAI221_X1 U5136 ( .B1(n4636), .B2(keyinput_f41), .C1(n4635), .C2(
        keyinput_f49), .A(n4634), .ZN(n4637) );
  NOR4_X1 U5137 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n4654)
         );
  AOI22_X1 U5138 ( .A1(n4642), .A2(keyinput_f15), .B1(keyinput_f19), .B2(n2501), .ZN(n4641) );
  OAI221_X1 U5139 ( .B1(n4642), .B2(keyinput_f15), .C1(n2501), .C2(
        keyinput_f19), .A(n4641), .ZN(n4652) );
  AOI22_X1 U5140 ( .A1(n4645), .A2(keyinput_f47), .B1(keyinput_f9), .B2(n4644), 
        .ZN(n4643) );
  OAI221_X1 U5141 ( .B1(n4645), .B2(keyinput_f47), .C1(n4644), .C2(keyinput_f9), .A(n4643), .ZN(n4651) );
  XNOR2_X1 U5142 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_f55), .ZN(n4649) );
  XNOR2_X1 U5143 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_f63), .ZN(n4648) );
  XNOR2_X1 U5144 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_f58), .ZN(n4647) );
  XNOR2_X1 U5145 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_f35), .ZN(n4646) );
  NAND4_X1 U5146 ( .A1(n4649), .A2(n4648), .A3(n4647), .A4(n4646), .ZN(n4650)
         );
  NOR3_X1 U5147 ( .A1(n4652), .A2(n4651), .A3(n4650), .ZN(n4653) );
  NAND4_X1 U5148 ( .A1(n4656), .A2(n4655), .A3(n4654), .A4(n4653), .ZN(n4695)
         );
  AOI22_X1 U5149 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(DATAI_23_), .B2(
        keyinput_f8), .ZN(n4657) );
  OAI221_X1 U5150 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(DATAI_23_), .C2(
        keyinput_f8), .A(n4657), .ZN(n4664) );
  AOI22_X1 U5151 ( .A1(DATAI_26_), .A2(keyinput_f5), .B1(DATAI_29_), .B2(
        keyinput_f2), .ZN(n4658) );
  OAI221_X1 U5152 ( .B1(DATAI_26_), .B2(keyinput_f5), .C1(DATAI_29_), .C2(
        keyinput_f2), .A(n4658), .ZN(n4663) );
  AOI22_X1 U5153 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_f42), .B1(DATAI_15_), 
        .B2(keyinput_f16), .ZN(n4659) );
  OAI221_X1 U5154 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_f42), .C1(DATAI_15_), .C2(keyinput_f16), .A(n4659), .ZN(n4662) );
  AOI22_X1 U5155 ( .A1(DATAI_19_), .A2(keyinput_f12), .B1(REG3_REG_3__SCAN_IN), 
        .B2(keyinput_f38), .ZN(n4660) );
  OAI221_X1 U5156 ( .B1(DATAI_19_), .B2(keyinput_f12), .C1(REG3_REG_3__SCAN_IN), .C2(keyinput_f38), .A(n4660), .ZN(n4661) );
  NOR4_X1 U5157 ( .A1(n4664), .A2(n4663), .A3(n4662), .A4(n4661), .ZN(n4693)
         );
  XNOR2_X1 U5158 ( .A(n4665), .B(keyinput_f44), .ZN(n4672) );
  AOI22_X1 U5159 ( .A1(REG3_REG_25__SCAN_IN), .A2(keyinput_f45), .B1(
        STATE_REG_SCAN_IN), .B2(keyinput_f32), .ZN(n4666) );
  OAI221_X1 U5160 ( .B1(REG3_REG_25__SCAN_IN), .B2(keyinput_f45), .C1(
        STATE_REG_SCAN_IN), .C2(keyinput_f32), .A(n4666), .ZN(n4671) );
  AOI22_X1 U5161 ( .A1(REG3_REG_20__SCAN_IN), .A2(keyinput_f53), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput_f40), .ZN(n4667) );
  OAI221_X1 U5162 ( .B1(REG3_REG_20__SCAN_IN), .B2(keyinput_f53), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput_f40), .A(n4667), .ZN(n4670) );
  AOI22_X1 U5163 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_f52), .B1(DATAI_1_), 
        .B2(keyinput_f30), .ZN(n4668) );
  OAI221_X1 U5164 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_f52), .C1(DATAI_1_), 
        .C2(keyinput_f30), .A(n4668), .ZN(n4669) );
  NOR4_X1 U5165 ( .A1(n4672), .A2(n4671), .A3(n4670), .A4(n4669), .ZN(n4692)
         );
  AOI22_X1 U5166 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_f34), .ZN(n4673) );
  OAI221_X1 U5167 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_f34), .A(n4673), .ZN(n4681) );
  AOI22_X1 U5168 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_f37), .B1(
        REG3_REG_16__SCAN_IN), .B2(keyinput_f46), .ZN(n4674) );
  OAI221_X1 U5169 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_f37), .C1(
        REG3_REG_16__SCAN_IN), .C2(keyinput_f46), .A(n4674), .ZN(n4680) );
  AOI22_X1 U5170 ( .A1(n2625), .A2(keyinput_f3), .B1(keyinput_f14), .B2(n2553), 
        .ZN(n4675) );
  OAI221_X1 U5171 ( .B1(n2625), .B2(keyinput_f3), .C1(n2553), .C2(keyinput_f14), .A(n4675), .ZN(n4679) );
  AOI22_X1 U5172 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(n4677), .B2(
        keyinput_f0), .ZN(n4676) );
  OAI221_X1 U5173 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(n4677), .C2(
        keyinput_f0), .A(n4676), .ZN(n4678) );
  NOR4_X1 U5174 ( .A1(n4681), .A2(n4680), .A3(n4679), .A4(n4678), .ZN(n4691)
         );
  AOI22_X1 U5175 ( .A1(DATAI_10_), .A2(keyinput_f21), .B1(DATAI_13_), .B2(
        keyinput_f18), .ZN(n4682) );
  OAI221_X1 U5176 ( .B1(DATAI_10_), .B2(keyinput_f21), .C1(DATAI_13_), .C2(
        keyinput_f18), .A(n4682), .ZN(n4689) );
  AOI22_X1 U5177 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(DATAI_6_), .B2(
        keyinput_f25), .ZN(n4683) );
  OAI221_X1 U5178 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(DATAI_6_), .C2(
        keyinput_f25), .A(n4683), .ZN(n4688) );
  AOI22_X1 U5179 ( .A1(DATAI_8_), .A2(keyinput_f23), .B1(DATAI_11_), .B2(
        keyinput_f20), .ZN(n4684) );
  OAI221_X1 U5180 ( .B1(DATAI_8_), .B2(keyinput_f23), .C1(DATAI_11_), .C2(
        keyinput_f20), .A(n4684), .ZN(n4687) );
  AOI22_X1 U5181 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_f59), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_f60), .ZN(n4685) );
  OAI221_X1 U5182 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_f59), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_f60), .A(n4685), .ZN(n4686) );
  NOR4_X1 U5183 ( .A1(n4689), .A2(n4688), .A3(n4687), .A4(n4686), .ZN(n4690)
         );
  NAND4_X1 U5184 ( .A1(n4693), .A2(n4692), .A3(n4691), .A4(n4690), .ZN(n4694)
         );
  OAI22_X1 U5185 ( .A1(keyinput_f24), .A2(n4696), .B1(n4695), .B2(n4694), .ZN(
        n4697) );
  OAI21_X1 U5186 ( .B1(n4697), .B2(keyinput_f24), .A(n4696), .ZN(n4699) );
  NAND3_X1 U5187 ( .A1(n4697), .A2(keyinput_g24), .A3(DATAI_7_), .ZN(n4698) );
  OAI21_X1 U5188 ( .B1(keyinput_g24), .B2(n4699), .A(n4698), .ZN(n4700) );
  OAI21_X1 U5189 ( .B1(n4702), .B2(n4701), .A(n4700), .ZN(n4703) );
  XOR2_X1 U5190 ( .A(n4704), .B(n4703), .Z(U3352) );
  CLKBUF_X1 U2297 ( .A(n2362), .Z(n2314) );
  NOR2_X2 U2994 ( .A1(n2858), .A2(n4480), .ZN(U4043) );
  NAND2_X2 U3025 ( .A1(n2689), .A2(n2688), .ZN(n2858) );
endmodule

