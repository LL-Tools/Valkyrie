

module b20_C_gen_AntiSAT_k_256_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4502, n4503, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5349, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497,
         n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507,
         n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517,
         n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527,
         n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537,
         n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547,
         n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557,
         n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
         n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577,
         n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587,
         n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597,
         n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607,
         n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
         n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627,
         n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637,
         n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647,
         n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
         n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
         n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
         n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687,
         n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
         n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707,
         n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717,
         n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727,
         n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737,
         n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747,
         n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757,
         n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767,
         n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777,
         n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787,
         n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817,
         n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827,
         n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837,
         n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
         n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857,
         n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867,
         n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877,
         n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887,
         n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897,
         n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907,
         n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917,
         n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927,
         n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
         n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
         n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957,
         n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
         n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987,
         n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997,
         n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007,
         n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017,
         n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027,
         n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037,
         n8038, n8039, n8040, n8041, n8042, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10533;

  AND2_X1 U5008 ( .A1(n8209), .A2(n8208), .ZN(n4502) );
  AND2_X1 U5010 ( .A1(n9123), .A2(n9124), .ZN(n4508) );
  AND4_X1 U5011 ( .A1(n8913), .A2(n9122), .A3(n4510), .A4(n5995), .ZN(n8960)
         );
  INV_X1 U5012 ( .A(n8914), .ZN(n4510) );
  CLKBUF_X1 U5013 ( .A(n7191), .Z(n4503) );
  OR4_X1 U5014 ( .A1(n8908), .A2(n8907), .A3(n9401), .A4(n9410), .ZN(n8909) );
  INV_X1 U5015 ( .A(n5479), .ZN(n7210) );
  AND2_X1 U5016 ( .A1(n4980), .A2(n4979), .ZN(n8358) );
  OR2_X1 U5017 ( .A1(n8330), .A2(n5262), .ZN(n4980) );
  NAND2_X1 U5018 ( .A1(n8075), .A2(n8241), .ZN(n8123) );
  AND2_X1 U5019 ( .A1(n8011), .A2(n7816), .ZN(n8001) );
  OR2_X1 U5020 ( .A1(n9560), .A2(n8835), .ZN(n9104) );
  AND2_X1 U5021 ( .A1(n7814), .A2(n5852), .ZN(n8142) );
  AOI21_X1 U5022 ( .B1(n8842), .B2(n5535), .A(n7794), .ZN(n8580) );
  AOI22_X1 U5023 ( .A1(n8547), .A2(n8545), .B1(n8536), .B2(n8709), .ZN(n8534)
         );
  XNOR2_X1 U5024 ( .A(n5808), .B(n5822), .ZN(n7731) );
  AND3_X1 U5025 ( .A1(n4983), .A2(n4981), .A3(n4607), .ZN(n5259) );
  NAND2_X1 U5026 ( .A1(n7532), .A2(n5568), .ZN(n7670) );
  OR2_X1 U5027 ( .A1(n7453), .A2(n7834), .ZN(n7454) );
  NAND2_X1 U5028 ( .A1(n5773), .A2(n5772), .ZN(n5789) );
  OAI21_X1 U5029 ( .B1(n9927), .B2(n4992), .A(n4993), .ZN(n5253) );
  NOR2_X1 U5030 ( .A1(n9928), .A2(n9929), .ZN(n9927) );
  NAND2_X1 U5031 ( .A1(n5078), .A2(n5076), .ZN(n5479) );
  OAI21_X1 U5032 ( .B1(n7320), .B2(n4974), .A(n4972), .ZN(n7550) );
  AND2_X1 U5033 ( .A1(n4991), .A2(n4540), .ZN(n9907) );
  NAND2_X1 U5034 ( .A1(n6957), .A2(n6956), .ZN(n6995) );
  AOI21_X1 U5035 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6619), .A(n6700), .ZN(
        n5242) );
  CLKBUF_X1 U5036 ( .A(n6605), .Z(n4506) );
  AND2_X1 U5037 ( .A1(n8997), .A2(n8984), .ZN(n8889) );
  CLKBUF_X1 U5038 ( .A(n7059), .Z(n4509) );
  NOR2_X1 U5039 ( .A1(n5240), .A2(n6670), .ZN(n6697) );
  OR2_X1 U5040 ( .A1(n6814), .A2(n6815), .ZN(n6862) );
  CLKBUF_X2 U5041 ( .A(n5452), .Z(n6572) );
  NOR2_X1 U5042 ( .A1(n9876), .A2(n9877), .ZN(n9875) );
  CLKBUF_X3 U5043 ( .A(n8087), .Z(n4514) );
  OR2_X1 U5045 ( .A1(n8293), .A2(n6846), .ZN(n7857) );
  CLKBUF_X2 U5046 ( .A(n8087), .Z(n4511) );
  INV_X1 U5047 ( .A(n6934), .ZN(n10011) );
  BUF_X2 U5048 ( .A(n8845), .Z(n4521) );
  INV_X1 U5049 ( .A(n5382), .ZN(n4879) );
  NOR2_X1 U5050 ( .A1(n6682), .A2(n6683), .ZN(n6681) );
  XNOR2_X1 U5051 ( .A(n8087), .B(n6810), .ZN(n6811) );
  NAND2_X1 U5052 ( .A1(n6807), .A2(n4539), .ZN(n8087) );
  INV_X1 U5053 ( .A(n5402), .ZN(n5832) );
  AND4_X2 U5054 ( .A1(n6011), .A2(n6012), .A3(n6013), .A4(n6010), .ZN(n7059)
         );
  INV_X1 U5055 ( .A(n8041), .ZN(n5357) );
  NAND2_X1 U5056 ( .A1(n8042), .A2(n8041), .ZN(n5452) );
  NAND2_X1 U5057 ( .A1(n5180), .A2(n5181), .ZN(n6678) );
  OAI21_X1 U5058 ( .B1(n6625), .B2(P2_D_REG_0__SCAN_IN), .A(n6626), .ZN(n6802)
         );
  OR2_X1 U5059 ( .A1(n5354), .A2(n5195), .ZN(n5356) );
  NAND2_X1 U5060 ( .A1(n5859), .A2(n5858), .ZN(n6625) );
  NAND2_X1 U5061 ( .A1(n8726), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5353) );
  XNOR2_X1 U5062 ( .A(n5144), .B(n5352), .ZN(n5235) );
  NAND2_X1 U5063 ( .A1(n9627), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5985) );
  OAI21_X1 U5064 ( .B1(n5122), .B2(n5085), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5144) );
  XNOR2_X1 U5065 ( .A(n5117), .B(n5116), .ZN(n7686) );
  AND2_X1 U5066 ( .A1(n5120), .A2(n5083), .ZN(n5354) );
  OR2_X1 U5067 ( .A1(n5227), .A2(n5135), .ZN(n5840) );
  INV_X2 U5068 ( .A(n7798), .ZN(n6605) );
  NAND2_X1 U5069 ( .A1(n5368), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5369) );
  INV_X1 U5070 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5367) );
  INV_X1 U5071 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U5072 ( .A1(n6863), .A2(n6864), .ZN(n6925) );
  NOR2_X2 U5073 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4875) );
  NAND2_X2 U5074 ( .A1(n5235), .A2(n5236), .ZN(n5374) );
  NOR2_X2 U5075 ( .A1(n5111), .A2(n5110), .ZN(n5112) );
  NAND2_X2 U5076 ( .A1(n8083), .A2(n8149), .ZN(n8151) );
  NAND2_X1 U5077 ( .A1(n6996), .A2(n6997), .ZN(n7032) );
  NAND2_X1 U5078 ( .A1(n7619), .A2(n7618), .ZN(n7634) );
  NAND2_X1 U5079 ( .A1(n8159), .A2(n8158), .ZN(n8053) );
  NAND2_X1 U5080 ( .A1(n8110), .A2(n4604), .ZN(n8177) );
  XNOR2_X2 U5081 ( .A(n5138), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6805) );
  OAI21_X1 U5082 ( .B1(n8210), .B2(n8264), .A(n4502), .ZN(P2_U3169) );
  NAND2_X2 U5083 ( .A1(n8151), .A2(n8086), .ZN(n8233) );
  NOR2_X2 U5084 ( .A1(n6579), .A2(n4548), .ZN(n8032) );
  AND4_X2 U5085 ( .A1(n4875), .A2(n5104), .A3(n5173), .A4(n4873), .ZN(n5194)
         );
  OAI211_X1 U5086 ( .C1(n5351), .C2(n9953), .A(n4505), .B(n10533), .ZN(
        P2_U3201) );
  NAND2_X1 U5087 ( .A1(n5349), .A2(n5002), .ZN(n4505) );
  XNOR2_X1 U5088 ( .A(n5247), .B(n9930), .ZN(n9928) );
  NOR2_X1 U5089 ( .A1(n8331), .A2(n8332), .ZN(n8330) );
  XNOR2_X1 U5090 ( .A(n5261), .B(n5620), .ZN(n8331) );
  NAND2_X1 U5091 ( .A1(n5474), .A2(n5473), .ZN(n5491) );
  NAND2_X1 U5092 ( .A1(n5414), .A2(n5413), .ZN(n5430) );
  NAND2_X1 U5093 ( .A1(n4507), .A2(n5601), .ZN(n5615) );
  NAND2_X1 U5094 ( .A1(n5532), .A2(n5100), .ZN(n5534) );
  OAI21_X1 U5095 ( .B1(n5381), .B2(n5373), .A(n6022), .ZN(n5390) );
  OAI21_X1 U5096 ( .B1(n5618), .B2(n4826), .A(n4824), .ZN(n5665) );
  OAI21_X1 U5097 ( .B1(n5680), .B2(n5679), .A(n5678), .ZN(n5696) );
  NAND2_X1 U5098 ( .A1(n5599), .A2(n5598), .ZN(n4507) );
  OAI21_X2 U5099 ( .B1(n8880), .B2(n7179), .A(n7079), .ZN(n7097) );
  AOI21_X1 U5100 ( .B1(n9126), .B2(n9125), .A(n4508), .ZN(n9132) );
  INV_X1 U5101 ( .A(n8025), .ZN(n5324) );
  NAND2_X1 U5102 ( .A1(n4786), .A2(n4787), .ZN(n5199) );
  INV_X1 U5103 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5176) );
  CLKBUF_X2 U5104 ( .A(n6054), .Z(n4512) );
  INV_X1 U5105 ( .A(n6054), .ZN(n6081) );
  INV_X1 U5106 ( .A(n6154), .ZN(n8841) );
  INV_X1 U5107 ( .A(n7807), .ZN(n6569) );
  INV_X2 U5108 ( .A(n8009), .ZN(n8012) );
  BUF_X1 U5109 ( .A(n5374), .Z(n6576) );
  INV_X1 U5110 ( .A(n7215), .ZN(n10021) );
  INV_X2 U5111 ( .A(n6304), .ZN(n6419) );
  OR2_X1 U5112 ( .A1(n6074), .A2(n6009), .ZN(n6011) );
  AND2_X1 U5113 ( .A1(n6377), .A2(n6376), .ZN(n9515) );
  NOR2_X1 U5114 ( .A1(n7178), .A2(n7186), .ZN(n7179) );
  INV_X1 U5115 ( .A(n5409), .ZN(n5535) );
  INV_X1 U5116 ( .A(n5988), .ZN(n9635) );
  AND2_X2 U5117 ( .A1(n7058), .A2(n9522), .ZN(n9730) );
  NOR2_X2 U5118 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6090) );
  OAI222_X1 U5119 ( .A1(n7790), .A2(P1_U3086), .B1(n9634), .B2(n8044), .C1(
        n10253), .C2(n9632), .ZN(P1_U3325) );
  AND2_X1 U5120 ( .A1(n7790), .A2(n9635), .ZN(n6025) );
  NAND2_X1 U5121 ( .A1(n5980), .A2(n6019), .ZN(n6054) );
  OAI21_X2 U5122 ( .B1(n7433), .B2(n4784), .A(n4783), .ZN(n7658) );
  XNOR2_X2 U5123 ( .A(n5219), .B(n6657), .ZN(n7433) );
  NAND2_X4 U5124 ( .A1(n5358), .A2(n5357), .ZN(n5402) );
  XNOR2_X2 U5125 ( .A(n5353), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5358) );
  AOI22_X1 U5126 ( .A1(n9382), .A2(n9381), .B1(n9380), .B2(n9379), .ZN(n9384)
         );
  AOI21_X1 U5128 ( .B1(n9490), .B2(n5033), .A(n4589), .ZN(n5031) );
  NAND2_X1 U5129 ( .A1(n8057), .A2(n8108), .ZN(n8110) );
  OR2_X1 U5130 ( .A1(n8649), .A2(n8435), .ZN(n7982) );
  NAND2_X1 U5131 ( .A1(n4893), .A2(n4892), .ZN(n6309) );
  OR2_X1 U5132 ( .A1(n9952), .A2(n9951), .ZN(n9955) );
  INV_X1 U5133 ( .A(n6056), .ZN(n6449) );
  AND3_X1 U5134 ( .A1(n5451), .A2(n5450), .A3(n5449), .ZN(n7023) );
  INV_X1 U5135 ( .A(n6125), .ZN(n6304) );
  INV_X2 U5136 ( .A(n4515), .ZN(n4517) );
  INV_X1 U5137 ( .A(n6074), .ZN(n8845) );
  INV_X1 U5138 ( .A(n6025), .ZN(n4515) );
  INV_X2 U5139 ( .A(n5452), .ZN(n5401) );
  INV_X1 U5140 ( .A(n5995), .ZN(n6726) );
  INV_X1 U5141 ( .A(n6016), .ZN(n9738) );
  CLKBUF_X2 U5142 ( .A(n5423), .Z(n7811) );
  INV_X1 U5143 ( .A(n7807), .ZN(n5420) );
  INV_X4 U5144 ( .A(n7798), .ZN(n6600) );
  NAND2_X1 U5145 ( .A1(n5194), .A2(n5105), .ZN(n5154) );
  AOI21_X1 U5146 ( .B1(n8024), .B2(n6804), .A(n8023), .ZN(n8031) );
  AND2_X1 U5147 ( .A1(n6407), .A2(n6408), .ZN(n4914) );
  CLKBUF_X1 U5148 ( .A(n6406), .Z(n4910) );
  NAND2_X1 U5149 ( .A1(n5031), .A2(n5030), .ZN(n9439) );
  AOI21_X1 U5150 ( .B1(n8415), .B2(n9981), .A(n8414), .ZN(n8640) );
  AND2_X1 U5151 ( .A1(n5049), .A2(n5048), .ZN(n8424) );
  NAND2_X1 U5152 ( .A1(n5019), .A2(n5018), .ZN(n7764) );
  NOR2_X1 U5153 ( .A1(n8395), .A2(n8394), .ZN(n8393) );
  XNOR2_X1 U5154 ( .A(n7797), .B(n7796), .ZN(n8842) );
  AND2_X1 U5155 ( .A1(n4902), .A2(n4898), .ZN(n7756) );
  AOI21_X1 U5156 ( .B1(n6312), .B2(n4555), .A(n4899), .ZN(n4898) );
  NAND2_X1 U5157 ( .A1(n6312), .A2(n6311), .ZN(n7702) );
  NAND2_X1 U5158 ( .A1(n6309), .A2(n6310), .ZN(n7701) );
  INV_X1 U5159 ( .A(n6309), .ZN(n6312) );
  AND2_X1 U5160 ( .A1(n5838), .A2(n5837), .ZN(n8101) );
  OAI22_X1 U5161 ( .A1(n8534), .A2(n8535), .B1(n8187), .B2(n8550), .ZN(n8526)
         );
  NAND2_X1 U5162 ( .A1(n5827), .A2(n5826), .ZN(n6559) );
  NAND2_X1 U5163 ( .A1(n5056), .A2(n5054), .ZN(n8547) );
  NAND2_X1 U5164 ( .A1(n6442), .A2(n6441), .ZN(n9570) );
  NAND2_X1 U5165 ( .A1(n4989), .A2(n4988), .ZN(n4987) );
  NAND2_X1 U5166 ( .A1(n6390), .A2(n6389), .ZN(n9593) );
  OR2_X1 U5167 ( .A1(n8294), .A2(n5260), .ZN(n4989) );
  NAND2_X1 U5168 ( .A1(n5780), .A2(n5779), .ZN(n5811) );
  INV_X1 U5169 ( .A(n5781), .ZN(n5780) );
  NAND2_X1 U5170 ( .A1(n5761), .A2(n10473), .ZN(n5781) );
  NAND2_X1 U5171 ( .A1(n4777), .A2(n4776), .ZN(n5213) );
  NAND2_X1 U5172 ( .A1(n4530), .A2(n4613), .ZN(n4777) );
  NAND2_X1 U5173 ( .A1(n6236), .A2(n6235), .ZN(n7569) );
  INV_X1 U5174 ( .A(n10043), .ZN(n7620) );
  AND2_X1 U5175 ( .A1(n5538), .A2(n5537), .ZN(n10043) );
  OAI21_X2 U5176 ( .B1(n6623), .B2(n6154), .A(n6158), .ZN(n9779) );
  XNOR2_X1 U5177 ( .A(n5532), .B(n5100), .ZN(n6638) );
  AND4_X1 U5178 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n7085)
         );
  AND4_X1 U5179 ( .A1(n6139), .A2(n6138), .A3(n6137), .A4(n6136), .ZN(n7279)
         );
  XNOR2_X1 U5180 ( .A(n4707), .B(n5505), .ZN(n6623) );
  OAI21_X1 U5181 ( .B1(n5524), .B2(n5523), .A(n5522), .ZN(n5532) );
  INV_X2 U5183 ( .A(n6336), .ZN(n8868) );
  NAND4_X1 U5184 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(n9984)
         );
  OAI211_X1 U5185 ( .C1(n6154), .C2(n6612), .A(n6045), .B(n6044), .ZN(n9745)
         );
  AND2_X1 U5186 ( .A1(n5191), .A2(n9896), .ZN(n5192) );
  NAND4_X1 U5187 ( .A1(n5380), .A2(n5379), .A3(n5378), .A4(n5377), .ZN(n8293)
         );
  OR2_X1 U5188 ( .A1(n6525), .A2(n5995), .ZN(n6723) );
  INV_X1 U5189 ( .A(n7803), .ZN(n5685) );
  NAND2_X1 U5190 ( .A1(n7850), .A2(n7852), .ZN(n8021) );
  XNOR2_X1 U5191 ( .A(n4885), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U5192 ( .A1(n4883), .A2(n4882), .ZN(n6525) );
  NAND2_X1 U5193 ( .A1(n5843), .A2(n5842), .ZN(n7852) );
  NAND2_X1 U5194 ( .A1(n6650), .A2(n6600), .ZN(n6154) );
  INV_X2 U5195 ( .A(n6650), .ZN(n6360) );
  NAND2_X1 U5196 ( .A1(n5233), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4976) );
  AOI21_X1 U5197 ( .B1(n4799), .B2(n4801), .A(n4567), .ZN(n4797) );
  NAND2_X1 U5198 ( .A1(n5127), .A2(n5126), .ZN(n7585) );
  XNOR2_X1 U5199 ( .A(n5987), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U5200 ( .A1(n5126), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5117) );
  OAI21_X1 U5201 ( .B1(n5962), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U5202 ( .A1(n5986), .A2(n5948), .ZN(n7793) );
  XNOR2_X1 U5203 ( .A(n5950), .B(n5949), .ZN(n6764) );
  OR2_X1 U5204 ( .A1(n5125), .A2(n5124), .ZN(n5127) );
  NAND2_X1 U5205 ( .A1(n4545), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5950) );
  NOR2_X1 U5206 ( .A1(n5154), .A2(n5075), .ZN(n4977) );
  NAND2_X1 U5207 ( .A1(n5178), .A2(n5184), .ZN(n9871) );
  INV_X1 U5208 ( .A(n5154), .ZN(n5073) );
  AND2_X1 U5209 ( .A1(n5112), .A2(n4563), .ZN(n5074) );
  OAI21_X1 U5210 ( .B1(n5177), .B2(n5176), .A(n5175), .ZN(n5178) );
  NAND2_X1 U5211 ( .A1(n5366), .A2(n5365), .ZN(n5370) );
  INV_X1 U5212 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5364) );
  INV_X1 U5213 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5363) );
  INV_X4 U5214 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U5215 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5107) );
  INV_X1 U5216 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5116) );
  INV_X1 U5217 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5958) );
  INV_X1 U5218 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5984) );
  INV_X1 U5219 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5974) );
  INV_X1 U5220 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5210) );
  INV_X1 U5221 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5158) );
  INV_X1 U5222 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5156) );
  NOR2_X1 U5223 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5933) );
  NOR2_X1 U5224 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5934) );
  NOR2_X2 U5225 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5237) );
  OAI21_X1 U5226 ( .B1(n9560), .B2(n9420), .A(n9400), .ZN(n9382) );
  NAND2_X2 U5227 ( .A1(n7819), .A2(n7816), .ZN(n8005) );
  XNOR2_X2 U5228 ( .A(n9384), .B(n9383), .ZN(n9552) );
  AND2_X1 U5229 ( .A1(n7790), .A2(n5988), .ZN(n6047) );
  MUX2_X1 U5230 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9636), .S(n6650), .Z(n7233) );
  OAI22_X2 U5231 ( .A1(n8444), .A2(n5769), .B1(n8281), .B2(n8662), .ZN(n8433)
         );
  OAI22_X2 U5232 ( .A1(n8457), .A2(n5752), .B1(n8467), .B2(n8594), .ZN(n8444)
         );
  NAND2_X1 U5233 ( .A1(n9647), .A2(n5020), .ZN(n5019) );
  INV_X2 U5235 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10269) );
  INV_X2 U5237 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10223) );
  NAND2_X1 U5238 ( .A1(n5979), .A2(n6019), .ZN(n6056) );
  INV_X1 U5239 ( .A(n6336), .ZN(n4519) );
  INV_X2 U5240 ( .A(n6336), .ZN(n4520) );
  CLKBUF_X1 U5241 ( .A(n6764), .Z(n4522) );
  AND2_X1 U5242 ( .A1(n5989), .A2(n5988), .ZN(n4523) );
  OR2_X2 U5243 ( .A1(n6584), .A2(n8142), .ZN(n7819) );
  AOI21_X2 U5244 ( .B1(n9411), .B2(n9410), .A(n5003), .ZN(n9402) );
  OAI21_X2 U5245 ( .B1(n5005), .B2(n5004), .A(n4566), .ZN(n9411) );
  OAI22_X2 U5246 ( .A1(n9503), .A2(n7767), .B1(n9532), .B2(n9515), .ZN(n9490)
         );
  NAND2_X1 U5247 ( .A1(n5821), .A2(n8426), .ZN(n5050) );
  INV_X1 U5248 ( .A(n8493), .ZN(n5723) );
  OR2_X1 U5249 ( .A1(n8633), .A2(n8278), .ZN(n8016) );
  NAND2_X1 U5250 ( .A1(n4626), .A2(n4694), .ZN(n4691) );
  AOI21_X1 U5251 ( .B1(n4694), .B2(n4693), .A(n8013), .ZN(n4692) );
  INV_X1 U5252 ( .A(n8004), .ZN(n4626) );
  INV_X1 U5253 ( .A(n7811), .ZN(n6568) );
  AND4_X1 U5254 ( .A1(n5630), .A2(n5629), .A3(n5628), .A4(n5627), .ZN(n8564)
         );
  NAND2_X1 U5255 ( .A1(n5374), .A2(n7798), .ZN(n5409) );
  NAND2_X1 U5256 ( .A1(n4927), .A2(n8773), .ZN(n4921) );
  NAND2_X1 U5257 ( .A1(n4635), .A2(n4634), .ZN(n4633) );
  NOR2_X1 U5258 ( .A1(n7946), .A2(n8009), .ZN(n4634) );
  NAND2_X1 U5259 ( .A1(n7948), .A2(n7947), .ZN(n4635) );
  NAND2_X1 U5260 ( .A1(n4623), .A2(n7972), .ZN(n7994) );
  INV_X1 U5261 ( .A(n8006), .ZN(n4703) );
  NAND2_X1 U5262 ( .A1(n8637), .A2(n7815), .ZN(n8011) );
  NOR2_X1 U5263 ( .A1(n5725), .A2(n4811), .ZN(n4810) );
  INV_X1 U5264 ( .A(n4813), .ZN(n4811) );
  INV_X1 U5265 ( .A(n5631), .ZN(n5632) );
  INV_X1 U5266 ( .A(SI_15_), .ZN(n10429) );
  NAND2_X1 U5267 ( .A1(n4700), .A2(n4697), .ZN(n4696) );
  AND2_X1 U5268 ( .A1(n4699), .A2(n8006), .ZN(n4697) );
  INV_X1 U5269 ( .A(n8008), .ZN(n4699) );
  INV_X1 U5270 ( .A(n5119), .ZN(n4834) );
  NOR2_X1 U5271 ( .A1(n7039), .A2(n7023), .ZN(n5079) );
  NOR2_X1 U5272 ( .A1(n5082), .A2(n5081), .ZN(n5080) );
  AND2_X1 U5273 ( .A1(n7039), .A2(n7023), .ZN(n5081) );
  INV_X1 U5274 ( .A(n5436), .ZN(n5082) );
  OR2_X1 U5275 ( .A1(n9971), .A2(n10016), .ZN(n7890) );
  NAND2_X1 U5276 ( .A1(n5876), .A2(n7854), .ZN(n7825) );
  NAND2_X1 U5277 ( .A1(n4571), .A2(n5051), .ZN(n5046) );
  NAND2_X1 U5278 ( .A1(n5118), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5131) );
  INV_X1 U5279 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5132) );
  INV_X1 U5280 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5228) );
  OR2_X1 U5281 ( .A1(n5154), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5203) );
  INV_X1 U5282 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5105) );
  AOI21_X1 U5283 ( .B1(n4895), .B2(n4897), .A(n4559), .ZN(n4892) );
  NAND2_X1 U5284 ( .A1(n7487), .A2(n4895), .ZN(n4893) );
  AND2_X1 U5285 ( .A1(n4670), .A2(n4666), .ZN(n4665) );
  OR2_X1 U5286 ( .A1(n9359), .A2(n9116), .ZN(n4666) );
  AND2_X1 U5287 ( .A1(n9539), .A2(n9134), .ZN(n4670) );
  OR2_X1 U5288 ( .A1(n9549), .A2(n8872), .ZN(n9109) );
  OR2_X1 U5289 ( .A1(n9565), .A2(n8756), .ZN(n9099) );
  OR2_X1 U5290 ( .A1(n9474), .A2(n5035), .ZN(n5028) );
  NAND2_X1 U5291 ( .A1(n5756), .A2(n5755), .ZN(n5771) );
  NAND2_X1 U5292 ( .A1(n5754), .A2(n5753), .ZN(n5756) );
  NAND2_X1 U5293 ( .A1(n5701), .A2(n5700), .ZN(n5712) );
  INV_X1 U5294 ( .A(n8090), .ZN(n4966) );
  AND2_X1 U5295 ( .A1(n4963), .A2(n8094), .ZN(n4962) );
  OR2_X1 U5296 ( .A1(n8095), .A2(n4969), .ZN(n4963) );
  INV_X1 U5297 ( .A(n6929), .ZN(n6926) );
  AND2_X1 U5298 ( .A1(n7814), .A2(n7813), .ZN(n8278) );
  NAND2_X1 U5299 ( .A1(n8042), .A2(n5357), .ZN(n5423) );
  OAI211_X1 U5300 ( .C1(n5199), .C2(n4782), .A(n4780), .B(n4778), .ZN(n9940)
         );
  AOI21_X1 U5301 ( .B1(n9904), .B2(n4781), .A(n4565), .ZN(n4780) );
  OR2_X1 U5302 ( .A1(n7194), .A2(n10060), .ZN(n4613) );
  INV_X1 U5303 ( .A(n8359), .ZN(n4979) );
  XNOR2_X1 U5304 ( .A(n5264), .B(n8375), .ZN(n8366) );
  NAND2_X1 U5305 ( .A1(n4573), .A2(n4528), .ZN(n5070) );
  NAND2_X1 U5306 ( .A1(n8494), .A2(n5709), .ZN(n5072) );
  NAND2_X1 U5307 ( .A1(n4528), .A2(n5709), .ZN(n5071) );
  AOI21_X1 U5308 ( .B1(n5061), .B2(n5059), .A(n5058), .ZN(n5057) );
  INV_X1 U5309 ( .A(n5581), .ZN(n5059) );
  INV_X1 U5310 ( .A(n7713), .ZN(n5058) );
  INV_X1 U5311 ( .A(n5061), .ZN(n5060) );
  AND3_X1 U5312 ( .A1(n5736), .A2(n5735), .A3(n5734), .ZN(n8480) );
  AND2_X1 U5313 ( .A1(n7940), .A2(n7936), .ZN(n4858) );
  AND2_X1 U5314 ( .A1(n5853), .A2(n8012), .ZN(n9983) );
  AND2_X1 U5315 ( .A1(n6816), .A2(n8012), .ZN(n9986) );
  OR2_X1 U5316 ( .A1(n4945), .A2(n8823), .ZN(n4940) );
  NAND2_X1 U5317 ( .A1(n4924), .A2(n4928), .ZN(n4922) );
  NAND2_X1 U5318 ( .A1(n4906), .A2(n7702), .ZN(n6329) );
  NAND2_X1 U5319 ( .A1(n9184), .A2(n9185), .ZN(n9183) );
  OR2_X1 U5320 ( .A1(n9261), .A2(n9262), .ZN(n4713) );
  NAND2_X1 U5321 ( .A1(n9403), .A2(n4732), .ZN(n9367) );
  NOR2_X1 U5322 ( .A1(n9359), .A2(n4733), .ZN(n4732) );
  OR2_X1 U5323 ( .A1(n9549), .A2(n9554), .ZN(n4733) );
  AND2_X1 U5324 ( .A1(n9575), .A2(n9461), .ZN(n4615) );
  XNOR2_X1 U5325 ( .A(n5793), .B(n5792), .ZN(n7698) );
  INV_X1 U5326 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5365) );
  INV_X1 U5327 ( .A(n8282), .ZN(n8467) );
  MUX2_X1 U5328 ( .A(P2_REG2_REG_26__SCAN_IN), .B(n8646), .S(n9999), .Z(n8430)
         );
  NAND2_X1 U5329 ( .A1(n8640), .A2(n10064), .ZN(n8581) );
  NAND2_X1 U5330 ( .A1(n5810), .A2(n5809), .ZN(n8642) );
  AND2_X1 U5331 ( .A1(n8980), .A2(n8982), .ZN(n4656) );
  NOR2_X1 U5332 ( .A1(n8996), .A2(n4658), .ZN(n4657) );
  NAND2_X1 U5333 ( .A1(n8983), .A2(n8997), .ZN(n4659) );
  OAI211_X1 U5334 ( .C1(n9005), .C2(n4644), .A(n4641), .B(n9009), .ZN(n9022)
         );
  NAND2_X1 U5335 ( .A1(n8990), .A2(n4642), .ZN(n4641) );
  NAND2_X1 U5336 ( .A1(n4690), .A2(n4685), .ZN(n7906) );
  INV_X1 U5337 ( .A(n4631), .ZN(n7902) );
  NAND2_X1 U5338 ( .A1(n4621), .A2(n7921), .ZN(n7923) );
  NAND2_X1 U5339 ( .A1(n4633), .A2(n4632), .ZN(n7950) );
  NAND2_X1 U5340 ( .A1(n4653), .A2(n4652), .ZN(n4651) );
  NAND2_X1 U5341 ( .A1(n4650), .A2(n4554), .ZN(n4649) );
  NAND2_X1 U5342 ( .A1(n8580), .A2(n8279), .ZN(n4795) );
  AND2_X1 U5343 ( .A1(n9102), .A2(n9103), .ZN(n4676) );
  OAI21_X1 U5344 ( .B1(n9100), .B2(n9094), .A(n4675), .ZN(n4674) );
  OR2_X1 U5345 ( .A1(n5711), .A2(n10442), .ZN(n4814) );
  INV_X1 U5346 ( .A(n8125), .ZN(n4953) );
  AOI21_X1 U5347 ( .B1(n8125), .B2(n4952), .A(n4951), .ZN(n4950) );
  INV_X1 U5348 ( .A(n8003), .ZN(n4702) );
  NAND2_X1 U5349 ( .A1(n4538), .A2(n8008), .ZN(n4701) );
  OAI21_X1 U5350 ( .B1(n8001), .B2(n8012), .A(n4794), .ZN(n8003) );
  NOR2_X1 U5351 ( .A1(n7976), .A2(n7975), .ZN(n4627) );
  INV_X1 U5352 ( .A(n7995), .ZN(n4628) );
  INV_X1 U5353 ( .A(n4795), .ZN(n8010) );
  NAND2_X1 U5354 ( .A1(n4795), .A2(n7819), .ZN(n8002) );
  AOI21_X1 U5355 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n4513), .A(n9875), .ZN(
        n5240) );
  OR2_X1 U5356 ( .A1(n5192), .A2(n9888), .ZN(n4786) );
  OR2_X1 U5357 ( .A1(n5203), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5166) );
  INV_X1 U5358 ( .A(n7337), .ZN(n4997) );
  OAI21_X1 U5359 ( .B1(n4836), .B2(n4835), .A(n4837), .ZN(n7806) );
  INV_X1 U5360 ( .A(n4838), .ZN(n4837) );
  NAND2_X1 U5361 ( .A1(n4529), .A2(n5839), .ZN(n4835) );
  OAI22_X1 U5362 ( .A1(n4840), .A2(n7820), .B1(n8144), .B2(n8101), .ZN(n4838)
         );
  NOR2_X1 U5363 ( .A1(n4857), .A2(n4850), .ZN(n4849) );
  INV_X1 U5364 ( .A(n7822), .ZN(n4850) );
  INV_X1 U5365 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10248) );
  NOR2_X1 U5366 ( .A1(n7922), .A2(n5062), .ZN(n5061) );
  INV_X1 U5367 ( .A(n5582), .ZN(n5062) );
  OR2_X1 U5368 ( .A1(n7616), .A2(n10039), .ZN(n7903) );
  NOR2_X1 U5369 ( .A1(n7881), .A2(n4872), .ZN(n4871) );
  NOR2_X1 U5370 ( .A1(n7829), .A2(n4869), .ZN(n4868) );
  INV_X1 U5371 ( .A(n5880), .ZN(n4869) );
  NOR2_X1 U5372 ( .A1(n5079), .A2(n8290), .ZN(n5077) );
  AND2_X1 U5373 ( .A1(n5861), .A2(n5899), .ZN(n6740) );
  NAND2_X1 U5374 ( .A1(n5050), .A2(n4552), .ZN(n5045) );
  NOR2_X1 U5375 ( .A1(n8655), .A2(n5053), .ZN(n5052) );
  INV_X1 U5376 ( .A(n8446), .ZN(n5053) );
  OR2_X1 U5377 ( .A1(n8662), .A2(n8460), .ZN(n7980) );
  OR2_X1 U5378 ( .A1(n8470), .A2(n8480), .ZN(n7968) );
  INV_X1 U5379 ( .A(n8528), .ZN(n8071) );
  AND2_X1 U5380 ( .A1(n8513), .A2(n7823), .ZN(n4854) );
  OR2_X1 U5381 ( .A1(n8697), .A2(n8516), .ZN(n7822) );
  OR2_X1 U5382 ( .A1(n8703), .A2(n8550), .ZN(n7940) );
  NOR3_X1 U5383 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5119) );
  INV_X1 U5384 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U5385 ( .A1(n5842), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5138) );
  INV_X1 U5386 ( .A(n5152), .ZN(n5133) );
  INV_X1 U5387 ( .A(n7752), .ZN(n4901) );
  NAND2_X1 U5388 ( .A1(n9460), .A2(n4750), .ZN(n4749) );
  INV_X1 U5389 ( .A(n8851), .ZN(n4750) );
  INV_X1 U5390 ( .A(n9492), .ZN(n4755) );
  NOR2_X1 U5391 ( .A1(n4744), .A2(n9608), .ZN(n4743) );
  INV_X1 U5392 ( .A(n4745), .ZN(n4744) );
  NOR2_X1 U5393 ( .A1(n8778), .A2(n5024), .ZN(n5023) );
  NOR2_X1 U5394 ( .A1(n7691), .A2(n5025), .ZN(n5024) );
  INV_X1 U5395 ( .A(n5023), .ZN(n5022) );
  NAND2_X1 U5396 ( .A1(n7691), .A2(n5025), .ZN(n5021) );
  AOI21_X1 U5397 ( .B1(n5017), .B2(n7609), .A(n5016), .ZN(n5015) );
  INV_X1 U5398 ( .A(n5015), .ZN(n5014) );
  NOR2_X1 U5399 ( .A1(n7470), .A2(n9031), .ZN(n4729) );
  AND2_X1 U5400 ( .A1(n7396), .A2(n7378), .ZN(n5006) );
  INV_X1 U5401 ( .A(n7381), .ZN(n5009) );
  INV_X1 U5402 ( .A(n6644), .ZN(n6521) );
  OR2_X1 U5404 ( .A1(n9490), .A2(n7769), .ZN(n5036) );
  INV_X1 U5405 ( .A(n7604), .ZN(n7605) );
  OR2_X1 U5406 ( .A1(n9116), .A2(n4510), .ZN(n9736) );
  NAND2_X1 U5407 ( .A1(n6019), .A2(n6598), .ZN(n6533) );
  NAND2_X1 U5408 ( .A1(n5803), .A2(n5802), .ZN(n5825) );
  AND2_X1 U5409 ( .A1(n5801), .A2(n5800), .ZN(n5802) );
  NAND2_X1 U5410 ( .A1(n5789), .A2(n5788), .ZN(n5803) );
  AND2_X1 U5411 ( .A1(n5772), .A2(n5759), .ZN(n5770) );
  NAND2_X1 U5412 ( .A1(n5712), .A2(n4814), .ZN(n4812) );
  NAND2_X1 U5413 ( .A1(n5711), .A2(n10442), .ZN(n4813) );
  INV_X1 U5414 ( .A(n4825), .ZN(n4824) );
  OAI21_X1 U5415 ( .B1(n4827), .B2(n4826), .A(n5649), .ZN(n4825) );
  NAND2_X1 U5416 ( .A1(n4816), .A2(n4815), .ZN(n5599) );
  AOI21_X1 U5417 ( .B1(n4817), .B2(n4533), .A(n4568), .ZN(n4815) );
  NOR2_X1 U5418 ( .A1(n5553), .A2(n4822), .ZN(n4821) );
  INV_X1 U5419 ( .A(n5533), .ZN(n4822) );
  AND2_X1 U5420 ( .A1(n7325), .A2(n7319), .ZN(n4975) );
  INV_X1 U5421 ( .A(n8286), .ZN(n8050) );
  INV_X1 U5422 ( .A(n8548), .ZN(n8223) );
  NOR2_X1 U5423 ( .A1(n8221), .A2(n4971), .ZN(n4970) );
  INV_X1 U5424 ( .A(n8052), .ZN(n4971) );
  INV_X1 U5425 ( .A(n4514), .ZN(n8136) );
  NAND2_X1 U5426 ( .A1(n4957), .A2(n4968), .ZN(n4956) );
  INV_X1 U5427 ( .A(n4959), .ZN(n4957) );
  AOI21_X1 U5428 ( .B1(n4962), .B2(n4965), .A(n4960), .ZN(n4959) );
  INV_X1 U5429 ( .A(n4962), .ZN(n4961) );
  NAND2_X1 U5430 ( .A1(n5143), .A2(n5086), .ZN(n5085) );
  OAI21_X1 U5431 ( .B1(n6678), .B2(n4998), .A(n5238), .ZN(n6682) );
  NOR2_X1 U5432 ( .A1(n6844), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4998) );
  OAI21_X1 U5433 ( .B1(n6678), .B2(n4789), .A(n5182), .ZN(n6680) );
  NOR2_X1 U5434 ( .A1(n9865), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4789) );
  NOR2_X1 U5435 ( .A1(n6680), .A2(n10050), .ZN(n6679) );
  XNOR2_X1 U5436 ( .A(n9871), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9877) );
  NOR2_X1 U5437 ( .A1(n4786), .A2(n5193), .ZN(n9887) );
  NAND2_X1 U5438 ( .A1(n4788), .A2(n4787), .ZN(n9889) );
  INV_X1 U5439 ( .A(n4991), .ZN(n4990) );
  AND2_X1 U5440 ( .A1(n9906), .A2(n5200), .ZN(n5201) );
  NAND2_X1 U5441 ( .A1(n9946), .A2(n5252), .ZN(n4993) );
  OR2_X1 U5442 ( .A1(n5250), .A2(n4994), .ZN(n4992) );
  INV_X1 U5443 ( .A(n5252), .ZN(n4994) );
  XNOR2_X1 U5444 ( .A(n5208), .B(n7196), .ZN(n7194) );
  NAND2_X1 U5445 ( .A1(n4785), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4784) );
  NAND2_X1 U5446 ( .A1(n5220), .A2(n4785), .ZN(n4783) );
  INV_X1 U5447 ( .A(n7659), .ZN(n4785) );
  OR2_X1 U5448 ( .A1(n7432), .A2(n4984), .ZN(n4983) );
  OR2_X1 U5449 ( .A1(n7656), .A2(n7536), .ZN(n4984) );
  NAND2_X1 U5450 ( .A1(n5258), .A2(n4982), .ZN(n4981) );
  INV_X1 U5451 ( .A(n7656), .ZN(n4982) );
  OR2_X1 U5452 ( .A1(n7432), .A2(n7536), .ZN(n4985) );
  INV_X1 U5453 ( .A(n8322), .ZN(n4988) );
  NOR2_X1 U5454 ( .A1(n5265), .A2(n8365), .ZN(n8395) );
  OR2_X1 U5455 ( .A1(n5830), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8033) );
  AOI21_X1 U5456 ( .B1(n5047), .B2(n5044), .A(n5041), .ZN(n6566) );
  NAND2_X1 U5457 ( .A1(n4574), .A2(n5042), .ZN(n5041) );
  AND2_X1 U5458 ( .A1(n4547), .A2(n6556), .ZN(n5044) );
  AOI21_X1 U5459 ( .B1(n4841), .B2(n8406), .A(n7996), .ZN(n4840) );
  INV_X1 U5460 ( .A(n4843), .ZN(n4841) );
  NAND2_X1 U5461 ( .A1(n5813), .A2(n8099), .ZN(n5830) );
  INV_X1 U5462 ( .A(n5762), .ZN(n5761) );
  AND2_X1 U5463 ( .A1(n7968), .A2(n7969), .ZN(n8468) );
  AOI21_X1 U5464 ( .B1(n8495), .B2(n7953), .A(n5885), .ZN(n8482) );
  NAND2_X1 U5465 ( .A1(n8490), .A2(n8489), .ZN(n8488) );
  OR2_X1 U5466 ( .A1(n5498), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U5467 ( .A1(n5515), .A2(n5514), .ZN(n5540) );
  INV_X1 U5468 ( .A(n5516), .ZN(n5515) );
  NAND2_X1 U5469 ( .A1(n6973), .A2(n4871), .ZN(n4870) );
  NAND2_X1 U5470 ( .A1(n4870), .A2(n4868), .ZN(n7411) );
  INV_X1 U5471 ( .A(n5079), .ZN(n5076) );
  AND3_X1 U5472 ( .A1(n5397), .A2(n5396), .A3(n5395), .ZN(n9989) );
  OR2_X1 U5473 ( .A1(n6576), .A2(n4513), .ZN(n5395) );
  AND2_X1 U5474 ( .A1(n5066), .A2(n5065), .ZN(n5064) );
  OR2_X1 U5475 ( .A1(n8470), .A2(n8283), .ZN(n5065) );
  NOR2_X1 U5476 ( .A1(n10044), .A2(n6805), .ZN(n5920) );
  NAND2_X1 U5477 ( .A1(n5704), .A2(n5703), .ZN(n8211) );
  OR2_X1 U5478 ( .A1(n8614), .A2(n8071), .ZN(n8501) );
  AND2_X1 U5479 ( .A1(n8501), .A2(n7949), .ZN(n8513) );
  NAND2_X1 U5480 ( .A1(n4855), .A2(n4854), .ZN(n8512) );
  OR2_X1 U5481 ( .A1(n8709), .A2(n8564), .ZN(n7936) );
  AND2_X1 U5482 ( .A1(n7940), .A2(n7939), .ZN(n8535) );
  NAND2_X1 U5483 ( .A1(n5883), .A2(n7942), .ZN(n4859) );
  AND2_X1 U5484 ( .A1(n5055), .A2(n5612), .ZN(n5054) );
  AND2_X1 U5485 ( .A1(n5375), .A2(n4877), .ZN(n10002) );
  NAND2_X1 U5486 ( .A1(n6576), .A2(n4878), .ZN(n4877) );
  OAI22_X1 U5487 ( .A1(n6606), .A2(n6605), .B1(n6607), .B2(n7798), .ZN(n4878)
         );
  NOR2_X1 U5488 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5113) );
  INV_X1 U5489 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U5490 ( .A1(n5229), .A2(n5228), .ZN(n5233) );
  INV_X1 U5491 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5104) );
  INV_X1 U5492 ( .A(n4914), .ZN(n4911) );
  NAND2_X1 U5493 ( .A1(n6125), .A2(n7233), .ZN(n6034) );
  OR2_X1 U5494 ( .A1(n7178), .A2(n6083), .ZN(n6030) );
  INV_X1 U5495 ( .A(n7704), .ZN(n4904) );
  NOR2_X1 U5496 ( .A1(n4542), .A2(n4900), .ZN(n4899) );
  NAND2_X1 U5497 ( .A1(n6328), .A2(n4901), .ZN(n4900) );
  NAND2_X1 U5498 ( .A1(n7701), .A2(n7704), .ZN(n4906) );
  OR2_X1 U5499 ( .A1(n6525), .A2(n8881), .ZN(n7068) );
  NAND2_X1 U5500 ( .A1(n4662), .A2(n4660), .ZN(n9121) );
  NOR2_X1 U5501 ( .A1(n4667), .A2(n4661), .ZN(n4660) );
  AND2_X1 U5502 ( .A1(n4665), .A2(n9547), .ZN(n4661) );
  AND4_X1 U5503 ( .A1(n6448), .A2(n6447), .A3(n6446), .A4(n6445), .ZN(n8787)
         );
  NAND2_X1 U5504 ( .A1(n4717), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6092) );
  INV_X1 U5505 ( .A(n6043), .ZN(n4717) );
  NAND2_X1 U5506 ( .A1(n9183), .A2(n4557), .ZN(n9669) );
  NAND2_X1 U5507 ( .A1(n9669), .A2(n9668), .ZN(n4709) );
  NOR2_X1 U5508 ( .A1(n9214), .A2(n4593), .ZN(n9229) );
  OR2_X1 U5509 ( .A1(n9229), .A2(n9228), .ZN(n4711) );
  NOR2_X1 U5510 ( .A1(n9259), .A2(n4714), .ZN(n9261) );
  AND2_X1 U5511 ( .A1(n9260), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4714) );
  NOR2_X1 U5512 ( .A1(n9288), .A2(n9289), .ZN(n9291) );
  OR2_X1 U5513 ( .A1(n9291), .A2(n9290), .ZN(n4716) );
  AND2_X1 U5514 ( .A1(n4716), .A2(n4715), .ZN(n9320) );
  NAND2_X1 U5515 ( .A1(n9311), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U5516 ( .A1(n9403), .A2(n9380), .ZN(n9385) );
  NOR2_X1 U5517 ( .A1(n9560), .A2(n9413), .ZN(n9403) );
  AND2_X1 U5518 ( .A1(n9565), .A2(n9434), .ZN(n5003) );
  NAND2_X1 U5519 ( .A1(n5033), .A2(n5026), .ZN(n5030) );
  AOI21_X1 U5520 ( .B1(n5028), .B2(n4524), .A(n4569), .ZN(n5033) );
  NOR2_X1 U5521 ( .A1(n9580), .A2(n9479), .ZN(n9454) );
  INV_X1 U5522 ( .A(n5028), .ZN(n5029) );
  NAND2_X1 U5523 ( .A1(n8967), .A2(n4758), .ZN(n4757) );
  INV_X1 U5524 ( .A(n9504), .ZN(n4758) );
  NAND2_X1 U5525 ( .A1(n7775), .A2(n4759), .ZN(n4756) );
  AND2_X1 U5526 ( .A1(n8938), .A2(n8940), .ZN(n8900) );
  INV_X1 U5527 ( .A(n8898), .ZN(n7611) );
  NOR2_X1 U5528 ( .A1(n9687), .A2(n4766), .ZN(n4765) );
  NAND2_X1 U5529 ( .A1(n7476), .A2(n9041), .ZN(n9688) );
  AND4_X1 U5530 ( .A1(n6266), .A2(n6265), .A3(n6264), .A4(n6263), .ZN(n9027)
         );
  NAND2_X1 U5531 ( .A1(n7402), .A2(n7383), .ZN(n7476) );
  AND2_X1 U5532 ( .A1(n8933), .A2(n9018), .ZN(n8893) );
  AND2_X1 U5533 ( .A1(n7382), .A2(n9015), .ZN(n7403) );
  NAND2_X1 U5534 ( .A1(n7403), .A2(n8893), .ZN(n7402) );
  AND2_X1 U5535 ( .A1(n9015), .A2(n9017), .ZN(n8894) );
  CLKBUF_X1 U5536 ( .A(n7379), .Z(n7303) );
  AND4_X1 U5537 ( .A1(n6242), .A2(n6241), .A3(n6240), .A4(n6239), .ZN(n7380)
         );
  AND2_X1 U5538 ( .A1(n9014), .A2(n9012), .ZN(n8890) );
  OR2_X1 U5539 ( .A1(n6177), .A2(n6176), .ZN(n6195) );
  NOR2_X1 U5540 ( .A1(n9736), .A2(n8919), .ZN(n6717) );
  OR2_X1 U5541 ( .A1(n7068), .A2(n9173), .ZN(n9693) );
  OR2_X1 U5542 ( .A1(n7068), .A2(n7793), .ZN(n9691) );
  NOR2_X1 U5543 ( .A1(n6016), .A2(n7233), .ZN(n7184) );
  NAND2_X1 U5544 ( .A1(n7798), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4679) );
  NAND2_X1 U5545 ( .A1(n8866), .A2(n8865), .ZN(n9549) );
  AOI21_X1 U5546 ( .B1(n4804), .B2(n4807), .A(n4803), .ZN(n4802) );
  INV_X1 U5547 ( .A(n5737), .ZN(n4803) );
  AND2_X1 U5548 ( .A1(n5755), .A2(n5742), .ZN(n5753) );
  OAI21_X1 U5549 ( .B1(n5712), .B2(n4809), .A(n4807), .ZN(n5739) );
  XNOR2_X1 U5550 ( .A(n5975), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8919) );
  AND3_X1 U5551 ( .A1(n5039), .A2(n4930), .A3(n5038), .ZN(n5969) );
  AND2_X1 U5552 ( .A1(n4932), .A2(n5954), .ZN(n4930) );
  AND3_X1 U5553 ( .A1(n5967), .A2(n6356), .A3(n5953), .ZN(n5954) );
  INV_X1 U5554 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U5555 ( .A1(n4823), .A2(n5633), .ZN(n5647) );
  NOR2_X1 U5556 ( .A1(n6156), .A2(n5936), .ZN(n6293) );
  OAI21_X1 U5557 ( .B1(n5534), .B2(n4527), .A(n4817), .ZN(n5586) );
  CLKBUF_X1 U5558 ( .A(n6155), .Z(n6156) );
  XNOR2_X1 U5559 ( .A(n5392), .B(n5371), .ZN(n5391) );
  INV_X1 U5560 ( .A(n6576), .ZN(n5684) );
  INV_X1 U5561 ( .A(n8007), .ZN(n8144) );
  AND2_X1 U5562 ( .A1(n5708), .A2(n5707), .ZN(n8479) );
  AND2_X1 U5563 ( .A1(n6757), .A2(n6756), .ZN(n8264) );
  AOI21_X1 U5564 ( .B1(n4544), .B2(n8018), .A(n8017), .ZN(n8022) );
  INV_X1 U5565 ( .A(n7465), .ZN(n8027) );
  NAND2_X1 U5566 ( .A1(n5751), .A2(n5750), .ZN(n8282) );
  AND3_X1 U5567 ( .A1(n5722), .A2(n5721), .A3(n5720), .ZN(n8493) );
  INV_X1 U5568 ( .A(n8479), .ZN(n8505) );
  NAND4_X1 U5569 ( .A1(n5428), .A2(n5427), .A3(n5426), .A4(n5425), .ZN(n9971)
         );
  OR2_X1 U5570 ( .A1(n5452), .A2(n5385), .ZN(n5387) );
  XNOR2_X1 U5571 ( .A(n5190), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9896) );
  INV_X1 U5572 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4874) );
  INV_X1 U5573 ( .A(n4777), .ZN(n7341) );
  INV_X1 U5574 ( .A(n5213), .ZN(n7339) );
  NOR2_X1 U5575 ( .A1(n4503), .A2(n5254), .ZN(n7338) );
  NOR2_X1 U5576 ( .A1(n8373), .A2(n8372), .ZN(n8377) );
  AND2_X1 U5577 ( .A1(n4793), .A2(n4792), .ZN(n8382) );
  NOR2_X1 U5578 ( .A1(n8396), .A2(n5000), .ZN(n4999) );
  AND2_X1 U5579 ( .A1(n9933), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n5000) );
  NAND2_X1 U5580 ( .A1(n5336), .A2(n9964), .ZN(n5347) );
  NAND2_X1 U5581 ( .A1(n4791), .A2(n5231), .ZN(n4790) );
  NAND2_X1 U5582 ( .A1(n9868), .A2(n5315), .ZN(n9953) );
  OAI211_X1 U5583 ( .C1(n6623), .C2(n5409), .A(n5495), .B(n4562), .ZN(n7321)
         );
  INV_X1 U5584 ( .A(n8558), .ZN(n9977) );
  NAND2_X1 U5585 ( .A1(n5923), .A2(n8566), .ZN(n9975) );
  AOI21_X1 U5586 ( .B1(n7698), .B2(n5535), .A(n5794), .ZN(n8584) );
  INV_X1 U5587 ( .A(n8668), .ZN(n8594) );
  NAND2_X1 U5588 ( .A1(n5856), .A2(n5855), .ZN(n5921) );
  AOI21_X1 U5589 ( .B1(n8280), .B2(n9986), .A(n5854), .ZN(n5855) );
  NAND2_X1 U5590 ( .A1(n8413), .A2(n8412), .ZN(n8414) );
  NAND2_X1 U5591 ( .A1(n8411), .A2(n9986), .ZN(n8412) );
  NAND2_X1 U5592 ( .A1(n4839), .A2(n4843), .ZN(n8407) );
  OR2_X1 U5593 ( .A1(n4836), .A2(n4844), .ZN(n4839) );
  AOI21_X1 U5594 ( .B1(n8280), .B2(n9983), .A(n8427), .ZN(n8428) );
  NOR2_X1 U5595 ( .A1(n8446), .A2(n8563), .ZN(n8427) );
  OR2_X1 U5596 ( .A1(n8653), .A2(n10049), .ZN(n4611) );
  INV_X1 U5597 ( .A(n8683), .ZN(n8717) );
  NAND2_X1 U5598 ( .A1(n10048), .A2(n10040), .ZN(n8683) );
  XNOR2_X1 U5599 ( .A(n5211), .B(n5210), .ZN(n7343) );
  INV_X1 U5600 ( .A(n4940), .ZN(n4937) );
  NOR2_X1 U5601 ( .A1(n4941), .A2(n8823), .ZN(n4939) );
  INV_X1 U5602 ( .A(n4942), .ZN(n4941) );
  AOI21_X1 U5603 ( .B1(n6471), .B2(n4944), .A(n4943), .ZN(n4942) );
  OAI21_X1 U5604 ( .B1(n4940), .B2(n4936), .A(n4598), .ZN(n4935) );
  INV_X1 U5605 ( .A(n6471), .ZN(n4936) );
  AND4_X1 U5606 ( .A1(n6200), .A2(n6199), .A3(n6198), .A4(n6197), .ZN(n7524)
         );
  AND2_X1 U5607 ( .A1(n4922), .A2(n4588), .ZN(n4915) );
  NAND2_X1 U5608 ( .A1(n8764), .A2(n4918), .ZN(n4917) );
  OR2_X1 U5609 ( .A1(n8793), .A2(n6386), .ZN(n6385) );
  NAND2_X1 U5610 ( .A1(n6255), .A2(n5099), .ZN(n7487) );
  INV_X1 U5611 ( .A(n9338), .ZN(n9675) );
  INV_X1 U5612 ( .A(n9351), .ZN(n9679) );
  AND2_X1 U5613 ( .A1(n8876), .A2(n8875), .ZN(n9362) );
  AND2_X1 U5614 ( .A1(n4772), .A2(n4770), .ZN(n9556) );
  AOI21_X1 U5615 ( .B1(n9420), .B2(n9711), .A(n4771), .ZN(n4770) );
  NAND2_X1 U5616 ( .A1(n4773), .A2(n9491), .ZN(n4772) );
  AND2_X1 U5617 ( .A1(n9135), .A2(n9708), .ZN(n4771) );
  NAND2_X1 U5618 ( .A1(n7317), .A2(n7078), .ZN(n9486) );
  OR2_X1 U5619 ( .A1(n9730), .A2(n7071), .ZN(n9521) );
  INV_X1 U5620 ( .A(n9486), .ZN(n9537) );
  AND2_X1 U5621 ( .A1(n7712), .A2(n7596), .ZN(n6655) );
  NAND2_X1 U5622 ( .A1(n4655), .A2(n4654), .ZN(n8986) );
  AOI21_X1 U5623 ( .B1(n4657), .B2(n4659), .A(n7242), .ZN(n4654) );
  AND2_X1 U5624 ( .A1(n8988), .A2(n4643), .ZN(n4642) );
  AND2_X1 U5625 ( .A1(n8989), .A2(n4644), .ZN(n4643) );
  NAND2_X1 U5626 ( .A1(n7899), .A2(n7900), .ZN(n4631) );
  OAI21_X1 U5627 ( .B1(n7901), .B2(n4687), .A(n4686), .ZN(n4685) );
  NOR2_X1 U5628 ( .A1(n4689), .A2(n4688), .ZN(n4687) );
  AND2_X1 U5629 ( .A1(n7908), .A2(n4581), .ZN(n4686) );
  INV_X1 U5630 ( .A(n7898), .ZN(n4689) );
  NAND2_X1 U5631 ( .A1(n7905), .A2(n8009), .ZN(n4690) );
  INV_X1 U5632 ( .A(n4629), .ZN(n7905) );
  OAI211_X1 U5633 ( .C1(n7904), .C2(n4631), .A(n7903), .B(n4630), .ZN(n4629)
         );
  OAI21_X1 U5634 ( .B1(n9022), .B2(n9011), .A(n9010), .ZN(n9013) );
  OR2_X1 U5635 ( .A1(n7917), .A2(n8012), .ZN(n4622) );
  NAND2_X1 U5636 ( .A1(n7916), .A2(n4706), .ZN(n4705) );
  AND2_X1 U5637 ( .A1(n7915), .A2(n8012), .ZN(n4706) );
  OAI21_X1 U5638 ( .B1(n4646), .B2(n4645), .A(n9047), .ZN(n9051) );
  NAND2_X1 U5639 ( .A1(n9046), .A2(n9045), .ZN(n4645) );
  AOI21_X1 U5640 ( .B1(n9042), .B2(n9041), .A(n4647), .ZN(n4646) );
  NAND2_X1 U5641 ( .A1(n9044), .A2(n9043), .ZN(n4647) );
  NAND2_X1 U5642 ( .A1(n7949), .A2(n8009), .ZN(n4632) );
  NAND2_X1 U5643 ( .A1(n4636), .A2(n4684), .ZN(n7948) );
  AND2_X1 U5644 ( .A1(n8525), .A2(n4580), .ZN(n4684) );
  NAND2_X1 U5645 ( .A1(n7938), .A2(n4553), .ZN(n4636) );
  NAND2_X1 U5646 ( .A1(n9065), .A2(n9060), .ZN(n4650) );
  NAND2_X1 U5647 ( .A1(n9065), .A2(n9064), .ZN(n4653) );
  NOR2_X1 U5648 ( .A1(n9063), .A2(n4644), .ZN(n4652) );
  NAND2_X1 U5649 ( .A1(n9069), .A2(n9507), .ZN(n4648) );
  OR2_X1 U5650 ( .A1(n7966), .A2(n8012), .ZN(n4625) );
  OR2_X1 U5651 ( .A1(n7967), .A2(n8009), .ZN(n4624) );
  OAI21_X1 U5652 ( .B1(n4640), .B2(n9085), .A(n4644), .ZN(n4639) );
  AOI21_X1 U5653 ( .B1(n9083), .B2(n9474), .A(n9084), .ZN(n4640) );
  NOR2_X1 U5654 ( .A1(n9105), .A2(n9097), .ZN(n4675) );
  INV_X1 U5655 ( .A(SI_8_), .ZN(n10416) );
  NAND2_X1 U5656 ( .A1(n8002), .A2(n8012), .ZN(n4794) );
  AOI21_X1 U5657 ( .B1(n7994), .B2(n7993), .A(n4680), .ZN(n7995) );
  NAND2_X1 U5658 ( .A1(n4681), .A2(n8406), .ZN(n4680) );
  INV_X1 U5659 ( .A(n7992), .ZN(n4681) );
  AOI21_X1 U5660 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6619), .A(n6706), .ZN(
        n5191) );
  INV_X1 U5661 ( .A(n8468), .ZN(n5069) );
  NAND2_X1 U5662 ( .A1(n8649), .A2(n8411), .ZN(n5051) );
  CLKBUF_X1 U5663 ( .A(n5876), .Z(n7858) );
  INV_X1 U5664 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5106) );
  INV_X1 U5665 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5108) );
  AND2_X1 U5666 ( .A1(n7574), .A2(n4896), .ZN(n4895) );
  OR2_X1 U5667 ( .A1(n7488), .A2(n4897), .ZN(n4896) );
  INV_X1 U5668 ( .A(n6274), .ZN(n4897) );
  OR2_X1 U5669 ( .A1(n9554), .A2(n9379), .ZN(n9103) );
  INV_X1 U5670 ( .A(n5738), .ZN(n4806) );
  NAND2_X1 U5671 ( .A1(n4600), .A2(n5633), .ZN(n4826) );
  INV_X1 U5672 ( .A(SI_17_), .ZN(n5650) );
  INV_X1 U5673 ( .A(n5493), .ZN(n4801) );
  INV_X1 U5674 ( .A(n4800), .ZN(n4799) );
  OAI21_X1 U5675 ( .B1(n5490), .B2(n4801), .A(n5505), .ZN(n4800) );
  INV_X1 U5676 ( .A(SI_18_), .ZN(n10254) );
  INV_X1 U5677 ( .A(SI_9_), .ZN(n10228) );
  INV_X1 U5678 ( .A(n8170), .ZN(n4960) );
  INV_X1 U5679 ( .A(n4700), .ZN(n4693) );
  INV_X1 U5680 ( .A(n8014), .ZN(n4695) );
  AND2_X1 U5681 ( .A1(n5198), .A2(n9930), .ZN(n4779) );
  INV_X1 U5682 ( .A(n5247), .ZN(n5248) );
  NOR2_X1 U5683 ( .A1(n5637), .A2(n8539), .ZN(n4978) );
  NOR2_X1 U5684 ( .A1(n5637), .A2(n8620), .ZN(n4614) );
  NAND2_X1 U5685 ( .A1(n5043), .A2(n6556), .ZN(n5042) );
  INV_X1 U5686 ( .A(n5045), .ZN(n5043) );
  OR2_X1 U5687 ( .A1(n8082), .A2(n8493), .ZN(n7954) );
  OR2_X1 U5688 ( .A1(n8211), .A2(n8479), .ZN(n7953) );
  INV_X1 U5689 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7660) );
  AND2_X1 U5690 ( .A1(n7904), .A2(n4871), .ZN(n4866) );
  AND2_X1 U5691 ( .A1(n5070), .A2(n5069), .ZN(n5068) );
  AND2_X1 U5692 ( .A1(n8594), .A2(n8282), .ZN(n7973) );
  NAND2_X1 U5693 ( .A1(n7620), .A2(n7644), .ZN(n7908) );
  CLKBUF_X1 U5694 ( .A(n9980), .Z(n4612) );
  NAND2_X1 U5695 ( .A1(n7353), .A2(n6209), .ZN(n7516) );
  AOI21_X1 U5696 ( .B1(n8773), .B2(n4920), .A(n4526), .ZN(n4919) );
  NAND2_X1 U5697 ( .A1(n4673), .A2(n9107), .ZN(n9108) );
  NAND2_X1 U5698 ( .A1(n4572), .A2(n4664), .ZN(n4663) );
  INV_X1 U5699 ( .A(n4665), .ZN(n4664) );
  NAND2_X1 U5700 ( .A1(n4668), .A2(n9122), .ZN(n4667) );
  NAND2_X1 U5701 ( .A1(n4672), .A2(n4669), .ZN(n4668) );
  NOR2_X1 U5702 ( .A1(n9547), .A2(n9116), .ZN(n4669) );
  NOR2_X1 U5703 ( .A1(n8769), .A2(n8778), .ZN(n4745) );
  INV_X1 U5704 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6345) );
  INV_X1 U5705 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6333) );
  OR2_X1 U5706 ( .A1(n6334), .A2(n6333), .ZN(n6346) );
  INV_X1 U5707 ( .A(n9044), .ZN(n4762) );
  INV_X1 U5708 ( .A(n7383), .ZN(n4763) );
  NOR2_X1 U5709 ( .A1(n6195), .A2(n6791), .ZN(n6223) );
  OR2_X1 U5710 ( .A1(n7363), .A2(n7524), .ZN(n9010) );
  AND2_X1 U5711 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6117) );
  OAI21_X1 U5712 ( .B1(n7785), .B2(n10227), .A(n7784), .ZN(n7797) );
  XNOR2_X1 U5713 ( .A(n7783), .B(n7782), .ZN(n7785) );
  INV_X1 U5714 ( .A(SI_28_), .ZN(n10485) );
  NAND2_X1 U5715 ( .A1(n5771), .A2(n5770), .ZN(n5773) );
  AND2_X1 U5716 ( .A1(n5801), .A2(n5776), .ZN(n5788) );
  AND2_X1 U5717 ( .A1(n4809), .A2(n4806), .ZN(n4804) );
  INV_X1 U5718 ( .A(n4810), .ZN(n4809) );
  AOI21_X1 U5719 ( .B1(n4808), .B2(n4810), .A(n4599), .ZN(n4807) );
  INV_X1 U5720 ( .A(n4814), .ZN(n4808) );
  NOR2_X1 U5721 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4932) );
  INV_X1 U5722 ( .A(SI_20_), .ZN(n10442) );
  NOR2_X1 U5723 ( .A1(n4828), .A2(n5634), .ZN(n4827) );
  INV_X1 U5724 ( .A(n5617), .ZN(n4828) );
  INV_X1 U5725 ( .A(n5552), .ZN(n4819) );
  INV_X1 U5726 ( .A(n4818), .ZN(n4817) );
  OAI21_X1 U5727 ( .B1(n4821), .B2(n4527), .A(n5569), .ZN(n4818) );
  OAI21_X1 U5728 ( .B1(n7798), .B2(n4638), .A(n4637), .ZN(n5472) );
  NAND2_X1 U5729 ( .A1(n7798), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4637) );
  XNOR2_X1 U5730 ( .A(n5472), .B(SI_5_), .ZN(n5462) );
  INV_X1 U5731 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4683) );
  NAND2_X1 U5732 ( .A1(n7798), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4682) );
  INV_X1 U5733 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10467) );
  NAND2_X1 U5734 ( .A1(n8177), .A2(n8066), .ZN(n8176) );
  INV_X1 U5735 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10473) );
  NAND2_X1 U5736 ( .A1(n4950), .A2(n4953), .ZN(n4948) );
  OR2_X1 U5737 ( .A1(n5705), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U5738 ( .A1(n5717), .A2(n10467), .ZN(n5732) );
  INV_X1 U5739 ( .A(n5718), .ZN(n5717) );
  NAND2_X1 U5740 ( .A1(n4698), .A2(n4696), .ZN(n8015) );
  NAND2_X1 U5741 ( .A1(n8004), .A2(n4700), .ZN(n4698) );
  XNOR2_X1 U5742 ( .A(n5146), .B(n5143), .ZN(n5236) );
  OR2_X1 U5743 ( .A1(n5145), .A2(n5195), .ZN(n5146) );
  OR2_X1 U5744 ( .A1(n7811), .A2(n5424), .ZN(n5425) );
  OR2_X1 U5745 ( .A1(n5402), .A2(n6879), .ZN(n5359) );
  NAND2_X1 U5746 ( .A1(n5129), .A2(n5128), .ZN(n5899) );
  NOR2_X1 U5747 ( .A1(n6681), .A2(n5239), .ZN(n9876) );
  INV_X1 U5748 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4876) );
  INV_X1 U5749 ( .A(n5199), .ZN(n9903) );
  NOR2_X1 U5750 ( .A1(n9940), .A2(n10057), .ZN(n9939) );
  NOR2_X1 U5751 ( .A1(n9927), .A2(n5250), .ZN(n9947) );
  INV_X1 U5752 ( .A(n7340), .ZN(n4776) );
  NOR2_X1 U5753 ( .A1(n5166), .A2(n5155), .ZN(n5214) );
  AOI21_X1 U5754 ( .B1(n5254), .B2(n4997), .A(n4594), .ZN(n4996) );
  NOR2_X1 U5755 ( .A1(n7662), .A2(n7680), .ZN(n4616) );
  AND2_X1 U5756 ( .A1(n4987), .A2(n4986), .ZN(n5261) );
  NAND2_X1 U5757 ( .A1(n8320), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4986) );
  INV_X1 U5758 ( .A(n8383), .ZN(n4792) );
  AND2_X1 U5759 ( .A1(n5812), .A2(n10456), .ZN(n5813) );
  OR2_X1 U5760 ( .A1(n5732), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5745) );
  OR2_X1 U5761 ( .A1(n5745), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U5762 ( .A1(n4848), .A2(n4851), .ZN(n8495) );
  AOI21_X1 U5763 ( .B1(n4856), .B2(n4853), .A(n4852), .ZN(n4851) );
  INV_X1 U5764 ( .A(n4854), .ZN(n4853) );
  NAND2_X1 U5765 ( .A1(n5689), .A2(n5688), .ZN(n5705) );
  INV_X1 U5766 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5688) );
  INV_X1 U5767 ( .A(n5690), .ZN(n5689) );
  NAND2_X1 U5768 ( .A1(n5656), .A2(n10248), .ZN(n5669) );
  OR2_X1 U5769 ( .A1(n5669), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U5770 ( .A1(n5624), .A2(n5623), .ZN(n5640) );
  INV_X1 U5771 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5623) );
  INV_X1 U5772 ( .A(n5625), .ZN(n5624) );
  OR2_X1 U5773 ( .A1(n5640), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5657) );
  OR2_X1 U5774 ( .A1(n5606), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U5775 ( .A1(n5590), .A2(n5589), .ZN(n5606) );
  INV_X1 U5776 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5589) );
  INV_X1 U5777 ( .A(n5591), .ZN(n5590) );
  OR2_X1 U5778 ( .A1(n5562), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U5779 ( .A1(n5574), .A2(n7660), .ZN(n5591) );
  INV_X1 U5780 ( .A(n5575), .ZN(n5574) );
  OR2_X1 U5781 ( .A1(n5540), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5562) );
  NOR2_X1 U5782 ( .A1(n4865), .A2(n4864), .ZN(n7450) );
  OAI21_X1 U5783 ( .B1(n4868), .B2(n4867), .A(n7899), .ZN(n4865) );
  AND2_X1 U5784 ( .A1(n6973), .A2(n4866), .ZN(n4864) );
  INV_X1 U5785 ( .A(n7904), .ZN(n4867) );
  AND2_X1 U5786 ( .A1(n7903), .A2(n7900), .ZN(n7834) );
  NAND2_X1 U5787 ( .A1(n5483), .A2(n5482), .ZN(n5498) );
  INV_X1 U5788 ( .A(n5484), .ZN(n5483) );
  NAND2_X1 U5789 ( .A1(n6736), .A2(n5891), .ZN(n7502) );
  OR2_X1 U5790 ( .A1(n5454), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U5791 ( .A1(n7890), .A2(n7877), .ZN(n7824) );
  AND4_X1 U5792 ( .A1(n5444), .A2(n5443), .A3(n5442), .A4(n5441), .ZN(n7039)
         );
  XNOR2_X1 U5793 ( .A(n9984), .B(n6934), .ZN(n9974) );
  INV_X1 U5794 ( .A(n7857), .ZN(n6871) );
  INV_X1 U5795 ( .A(n7825), .ZN(n6874) );
  AND2_X1 U5796 ( .A1(n5860), .A2(n8009), .ZN(n5914) );
  NAND2_X1 U5797 ( .A1(n5873), .A2(n6629), .ZN(n5915) );
  AND3_X1 U5798 ( .A1(n6740), .A2(n5903), .A3(n6631), .ZN(n5919) );
  NAND2_X1 U5799 ( .A1(n5040), .A2(n5045), .ZN(n6557) );
  NAND2_X1 U5800 ( .A1(n5047), .A2(n4547), .ZN(n5040) );
  AND2_X1 U5801 ( .A1(n5829), .A2(n5828), .ZN(n8007) );
  NAND2_X1 U5802 ( .A1(n5047), .A2(n5046), .ZN(n8409) );
  NAND2_X1 U5803 ( .A1(n8410), .A2(n9983), .ZN(n8413) );
  NAND2_X1 U5804 ( .A1(n7982), .A2(n7987), .ZN(n4846) );
  OR2_X1 U5805 ( .A1(n7973), .A2(n8449), .ZN(n8458) );
  AND4_X1 U5806 ( .A1(n5645), .A2(n5644), .A3(n5643), .A4(n5642), .ZN(n8550)
         );
  NAND2_X1 U5807 ( .A1(n4863), .A2(n4861), .ZN(n8569) );
  AOI21_X1 U5808 ( .B1(n7838), .B2(n4531), .A(n4862), .ZN(n4861) );
  NOR2_X1 U5809 ( .A1(n7925), .A2(n8285), .ZN(n4862) );
  AOI21_X1 U5810 ( .B1(n7498), .B2(n5548), .A(n5547), .ZN(n7530) );
  AND3_X1 U5811 ( .A1(n5435), .A2(n5434), .A3(n5433), .ZN(n10016) );
  NOR2_X1 U5812 ( .A1(n6748), .A2(n5904), .ZN(n6755) );
  AND2_X1 U5813 ( .A1(n5899), .A2(n6631), .ZN(n6746) );
  NOR2_X1 U5814 ( .A1(n5084), .A2(n5085), .ZN(n5083) );
  NAND2_X1 U5815 ( .A1(n5119), .A2(n5352), .ZN(n5084) );
  INV_X1 U5816 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5355) );
  AND2_X1 U5817 ( .A1(n5123), .A2(n4832), .ZN(n5858) );
  NAND2_X1 U5818 ( .A1(n5115), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U5819 ( .A1(n5137), .A2(n5136), .ZN(n5842) );
  INV_X1 U5820 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5136) );
  INV_X1 U5821 ( .A(n5840), .ZN(n5137) );
  NAND2_X1 U5822 ( .A1(n4977), .A2(n5150), .ZN(n5152) );
  NAND2_X1 U5823 ( .A1(n5103), .A2(n5237), .ZN(n5186) );
  AND2_X1 U5824 ( .A1(n4876), .A2(n5176), .ZN(n5103) );
  OR2_X1 U5825 ( .A1(n6450), .A2(n7172), .ZN(n6126) );
  INV_X1 U5826 ( .A(n6592), .ZN(n4943) );
  INV_X1 U5827 ( .A(n6411), .ZN(n6412) );
  XNOR2_X1 U5828 ( .A(n6082), .B(n6081), .ZN(n6088) );
  OR2_X1 U5829 ( .A1(n4891), .A2(n6072), .ZN(n6080) );
  NOR2_X1 U5830 ( .A1(n4532), .A2(n4920), .ZN(n4918) );
  NAND2_X1 U5831 ( .A1(n8763), .A2(n4926), .ZN(n4916) );
  OR2_X1 U5832 ( .A1(n6592), .A2(n6591), .ZN(n4945) );
  NOR2_X1 U5833 ( .A1(n4890), .A2(n4889), .ZN(n4888) );
  INV_X1 U5834 ( .A(n7368), .ZN(n4889) );
  NAND2_X1 U5835 ( .A1(n4912), .A2(n8731), .ZN(n4909) );
  NAND2_X1 U5836 ( .A1(n8781), .A2(n6439), .ZN(n4912) );
  NAND2_X1 U5837 ( .A1(n4907), .A2(n4911), .ZN(n8783) );
  NAND2_X1 U5838 ( .A1(n6884), .A2(n6885), .ZN(n4886) );
  INV_X1 U5839 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6279) );
  AND2_X1 U5840 ( .A1(n6223), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U5841 ( .A1(n6237), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U5842 ( .A1(n6053), .A2(n5091), .ZN(n6055) );
  OR2_X1 U5843 ( .A1(n6083), .A2(n7063), .ZN(n5091) );
  NOR2_X1 U5844 ( .A1(n6346), .A2(n6345), .ZN(n6363) );
  AND2_X1 U5845 ( .A1(n6363), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6365) );
  INV_X1 U5846 ( .A(n6372), .ZN(n4925) );
  AND2_X1 U5847 ( .A1(n6535), .A2(n6534), .ZN(n8832) );
  AND4_X1 U5848 ( .A1(n6463), .A2(n6462), .A3(n6461), .A4(n6460), .ZN(n8756)
         );
  MUX2_X1 U5849 ( .A(n6009), .B(P1_REG2_REG_1__SCAN_IN), .S(n9158), .Z(n9154)
         );
  OR2_X1 U5850 ( .A1(n9165), .A2(n5101), .ZN(n9184) );
  AND2_X1 U5851 ( .A1(n4709), .A2(n4708), .ZN(n9203) );
  NAND2_X1 U5852 ( .A1(n9676), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4708) );
  NOR2_X1 U5853 ( .A1(n9203), .A2(n9202), .ZN(n9201) );
  AND2_X1 U5854 ( .A1(n4711), .A2(n4710), .ZN(n9242) );
  NAND2_X1 U5855 ( .A1(n6777), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4710) );
  NOR2_X1 U5856 ( .A1(n9242), .A2(n9241), .ZN(n9240) );
  AOI21_X1 U5857 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6776), .A(n9240), .ZN(
        n6772) );
  AOI21_X1 U5858 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6941), .A(n6940), .ZN(
        n6944) );
  OR2_X1 U5859 ( .A1(n6256), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6275) );
  AND2_X1 U5860 ( .A1(n4713), .A2(n9258), .ZN(n9287) );
  NAND2_X1 U5861 ( .A1(n9372), .A2(n4774), .ZN(n4773) );
  OR2_X1 U5862 ( .A1(n7778), .A2(n7779), .ZN(n4774) );
  NAND2_X1 U5863 ( .A1(n9412), .A2(n7770), .ZN(n9413) );
  NOR2_X1 U5864 ( .A1(n9570), .A2(n9449), .ZN(n5004) );
  OAI22_X1 U5865 ( .A1(n9467), .A2(n4747), .B1(n4748), .B2(n7776), .ZN(n9432)
         );
  NAND2_X1 U5866 ( .A1(n9460), .A2(n9091), .ZN(n4747) );
  AND2_X1 U5867 ( .A1(n7777), .A2(n4749), .ZN(n4748) );
  NAND2_X1 U5868 ( .A1(n9432), .A2(n9433), .ZN(n9431) );
  NOR2_X1 U5869 ( .A1(n9440), .A2(n9570), .ZN(n9412) );
  NAND2_X1 U5870 ( .A1(n9454), .A2(n9445), .ZN(n9440) );
  NAND2_X1 U5871 ( .A1(n9467), .A2(n8851), .ZN(n9459) );
  NAND2_X1 U5872 ( .A1(n9459), .A2(n9460), .ZN(n9458) );
  NAND2_X1 U5873 ( .A1(n7768), .A2(n7769), .ZN(n5027) );
  NAND2_X1 U5874 ( .A1(n9478), .A2(n9586), .ZN(n9479) );
  OAI21_X1 U5875 ( .B1(n7775), .B2(n4754), .A(n4751), .ZN(n9468) );
  AOI21_X1 U5876 ( .B1(n4753), .B2(n4760), .A(n4752), .ZN(n4751) );
  NAND2_X1 U5877 ( .A1(n7775), .A2(n9058), .ZN(n9505) );
  AND2_X1 U5878 ( .A1(n8967), .A2(n8969), .ZN(n9504) );
  AND2_X1 U5879 ( .A1(n7605), .A2(n4582), .ZN(n9519) );
  AND2_X1 U5880 ( .A1(n9066), .A2(n9058), .ZN(n9529) );
  NAND2_X1 U5881 ( .A1(n7605), .A2(n4743), .ZN(n9520) );
  OAI21_X1 U5882 ( .B1(n7742), .B2(n9054), .A(n8938), .ZN(n7743) );
  NAND2_X1 U5883 ( .A1(n7743), .A2(n7744), .ZN(n9528) );
  NAND2_X1 U5884 ( .A1(n5023), .A2(n5025), .ZN(n5018) );
  NAND2_X1 U5885 ( .A1(n5022), .A2(n5021), .ZN(n5020) );
  INV_X1 U5886 ( .A(n8902), .ZN(n7744) );
  NAND2_X1 U5887 ( .A1(n7687), .A2(n9048), .ZN(n7742) );
  NAND2_X1 U5888 ( .A1(n7605), .A2(n9645), .ZN(n7692) );
  AND2_X1 U5889 ( .A1(n9050), .A2(n9048), .ZN(n8898) );
  NAND2_X1 U5890 ( .A1(n5015), .A2(n7480), .ZN(n5011) );
  NAND2_X1 U5891 ( .A1(n4575), .A2(n5014), .ZN(n5013) );
  NOR2_X1 U5892 ( .A1(n7609), .A2(n4727), .ZN(n4725) );
  INV_X1 U5893 ( .A(n4767), .ZN(n7477) );
  OAI21_X1 U5894 ( .B1(n7402), .B2(n4764), .A(n4761), .ZN(n4767) );
  INV_X1 U5895 ( .A(n4765), .ZN(n4764) );
  AOI21_X1 U5896 ( .B1(n4765), .B2(n4763), .A(n4762), .ZN(n4761) );
  NAND2_X1 U5897 ( .A1(n7477), .A2(n8899), .ZN(n7600) );
  OR2_X1 U5898 ( .A1(n6280), .A2(n6279), .ZN(n6298) );
  NAND2_X1 U5899 ( .A1(n7397), .A2(n4729), .ZN(n9698) );
  AOI21_X1 U5900 ( .B1(n7396), .B2(n5009), .A(n4561), .ZN(n5007) );
  INV_X1 U5901 ( .A(n8895), .ZN(n7468) );
  AND2_X1 U5902 ( .A1(n7397), .A2(n9816), .ZN(n7398) );
  NOR2_X1 U5903 ( .A1(n7378), .A2(n7305), .ZN(n7306) );
  NOR2_X1 U5904 ( .A1(n4739), .A2(n9720), .ZN(n4737) );
  NAND2_X1 U5905 ( .A1(n9795), .A2(n4740), .ZN(n4739) );
  INV_X1 U5906 ( .A(n7286), .ZN(n4738) );
  NAND2_X1 U5907 ( .A1(n4738), .A2(n4735), .ZN(n7312) );
  NOR2_X1 U5908 ( .A1(n7526), .A2(n4736), .ZN(n4735) );
  INV_X1 U5909 ( .A(n4737), .ZN(n4736) );
  AND4_X1 U5910 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n7300)
         );
  NOR3_X1 U5911 ( .A1(n7286), .A2(n9720), .A3(n9779), .ZN(n9721) );
  NOR2_X1 U5912 ( .A1(n6134), .A2(n6133), .ZN(n6159) );
  NOR2_X1 U5913 ( .A1(n7286), .A2(n9779), .ZN(n9724) );
  AND4_X1 U5914 ( .A1(n6182), .A2(n6181), .A3(n6180), .A4(n6179), .ZN(n7361)
         );
  NOR2_X1 U5915 ( .A1(n7090), .A2(n9757), .ZN(n7270) );
  NAND2_X1 U5916 ( .A1(n4731), .A2(n6072), .ZN(n7090) );
  INV_X1 U5917 ( .A(n9693), .ZN(n9708) );
  INV_X1 U5918 ( .A(n9362), .ZN(n9539) );
  AND2_X1 U5919 ( .A1(n9387), .A2(n9386), .ZN(n9548) );
  NAND2_X1 U5920 ( .A1(n6455), .A2(n6454), .ZN(n9565) );
  NAND2_X1 U5921 ( .A1(n6410), .A2(n6409), .ZN(n9580) );
  AND2_X1 U5922 ( .A1(n5036), .A2(n5029), .ZN(n9476) );
  NAND2_X1 U5923 ( .A1(n5036), .A2(n7768), .ZN(n9475) );
  OR2_X1 U5924 ( .A1(n7072), .A2(n8955), .ZN(n9828) );
  NOR2_X1 U5925 ( .A1(n6721), .A2(n7054), .ZN(n9544) );
  NAND2_X1 U5926 ( .A1(n5825), .A2(n5824), .ZN(n5827) );
  INV_X1 U5927 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5949) );
  AND2_X1 U5928 ( .A1(n5825), .A2(n5823), .ZN(n5808) );
  NAND2_X1 U5929 ( .A1(n5961), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5957) );
  XNOR2_X1 U5930 ( .A(n6524), .B(n6523), .ZN(n7509) );
  NAND2_X1 U5931 ( .A1(n4881), .A2(n5977), .ZN(n6522) );
  AOI21_X1 U5932 ( .B1(n5976), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_22__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U5933 ( .A1(n4812), .A2(n4813), .ZN(n5726) );
  INV_X1 U5934 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U5935 ( .A1(n6357), .A2(n6356), .ZN(n6359) );
  NAND2_X1 U5936 ( .A1(n4820), .A2(n5552), .ZN(n5571) );
  INV_X1 U5937 ( .A(n5462), .ZN(n5467) );
  XNOR2_X1 U5938 ( .A(n5446), .B(n10266), .ZN(n5468) );
  XNOR2_X1 U5939 ( .A(n5412), .B(n5394), .ZN(n5410) );
  AND2_X1 U5940 ( .A1(n7320), .A2(n7319), .ZN(n7326) );
  OAI21_X1 U5941 ( .B1(n8435), .B2(n4967), .A(n8098), .ZN(n8135) );
  NAND2_X1 U5942 ( .A1(n4955), .A2(n4954), .ZN(n8098) );
  AOI21_X1 U5943 ( .B1(n4956), .B2(n4525), .A(n4536), .ZN(n4954) );
  AND2_X1 U5944 ( .A1(n5768), .A2(n5767), .ZN(n8460) );
  NAND2_X1 U5945 ( .A1(n8123), .A2(n8124), .ZN(n4949) );
  INV_X1 U5946 ( .A(n4973), .ZN(n4972) );
  OAI21_X1 U5947 ( .B1(n4975), .B2(n4974), .A(n7423), .ZN(n4973) );
  INV_X1 U5948 ( .A(n7424), .ZN(n4974) );
  NAND2_X1 U5949 ( .A1(n8049), .A2(n8048), .ZN(n8159) );
  NAND2_X1 U5950 ( .A1(n4958), .A2(n4962), .ZN(n8169) );
  NAND2_X1 U5951 ( .A1(n8233), .A2(n4964), .ZN(n4958) );
  INV_X1 U5952 ( .A(n8287), .ZN(n7644) );
  NAND2_X1 U5953 ( .A1(n8053), .A2(n8052), .ZN(n8222) );
  NAND2_X1 U5954 ( .A1(n5731), .A2(n5730), .ZN(n8470) );
  NAND2_X1 U5955 ( .A1(n6759), .A2(n9990), .ZN(n8236) );
  AND4_X1 U5956 ( .A1(n5695), .A2(n5694), .A3(n5693), .A4(n5692), .ZN(n8517)
         );
  AND2_X1 U5957 ( .A1(n6817), .A2(n6816), .ZN(n8269) );
  INV_X1 U5958 ( .A(n8264), .ZN(n8244) );
  NAND2_X1 U5959 ( .A1(n8110), .A2(n8060), .ZN(n8266) );
  OR2_X1 U5960 ( .A1(n6932), .A2(n6931), .ZN(n8273) );
  AOI21_X1 U5961 ( .B1(n7849), .B2(n6805), .A(n7848), .ZN(n7851) );
  NOR2_X1 U5962 ( .A1(n4550), .A2(n6805), .ZN(n7848) );
  INV_X1 U5963 ( .A(n8278), .ZN(n8400) );
  INV_X1 U5964 ( .A(n8101), .ZN(n8410) );
  NAND2_X1 U5965 ( .A1(n5820), .A2(n5819), .ZN(n8280) );
  AND2_X1 U5966 ( .A1(n5787), .A2(n5786), .ZN(n8446) );
  INV_X1 U5967 ( .A(n8460), .ZN(n8281) );
  INV_X1 U5968 ( .A(n8564), .ZN(n8536) );
  AND4_X1 U5969 ( .A1(n5521), .A2(n5520), .A3(n5519), .A4(n5518), .ZN(n7616)
         );
  NAND4_X1 U5970 ( .A1(n5504), .A2(n5503), .A3(n5502), .A4(n5501), .ZN(n8288)
         );
  INV_X1 U5971 ( .A(n7039), .ZN(n8291) );
  OR2_X1 U5972 ( .A1(n5899), .A2(n6751), .ZN(n8292) );
  INV_X1 U5973 ( .A(n6616), .ZN(n6670) );
  NAND2_X1 U5974 ( .A1(n4540), .A2(n5243), .ZN(n9891) );
  OR2_X1 U5975 ( .A1(n9947), .A2(n9946), .ZN(n9950) );
  INV_X1 U5976 ( .A(n4613), .ZN(n7193) );
  NOR2_X1 U5977 ( .A1(n7433), .A2(n5561), .ZN(n7436) );
  NAND2_X1 U5978 ( .A1(n4983), .A2(n4981), .ZN(n7655) );
  NOR2_X1 U5979 ( .A1(P2_U3150), .A2(n5343), .ZN(n9933) );
  INV_X1 U5980 ( .A(n4989), .ZN(n8323) );
  INV_X1 U5981 ( .A(n4987), .ZN(n8321) );
  INV_X1 U5982 ( .A(n4980), .ZN(n8360) );
  AND2_X1 U5983 ( .A1(n4842), .A2(n4840), .ZN(n6567) );
  OAI21_X1 U5984 ( .B1(n8490), .B2(n5071), .A(n5070), .ZN(n8465) );
  NAND2_X1 U5985 ( .A1(n8488), .A2(n5709), .ZN(n8477) );
  NAND2_X1 U5986 ( .A1(n5668), .A2(n5667), .ZN(n8614) );
  OAI21_X1 U5987 ( .B1(n7670), .B2(n5060), .A(n5057), .ZN(n8559) );
  INV_X1 U5988 ( .A(n7429), .ZN(n10031) );
  NAND2_X1 U5989 ( .A1(n4870), .A2(n5880), .ZN(n7256) );
  INV_X1 U5990 ( .A(n9975), .ZN(n8555) );
  AND2_X1 U5991 ( .A1(n5922), .A2(n9990), .ZN(n5088) );
  INV_X1 U5992 ( .A(n10042), .ZN(n10040) );
  INV_X2 U5993 ( .A(n5088), .ZN(n9999) );
  AOI21_X1 U5994 ( .B1(n7583), .B2(n5535), .A(n5760), .ZN(n8590) );
  NAND2_X1 U5995 ( .A1(n7805), .A2(n7804), .ZN(n8633) );
  INV_X1 U5996 ( .A(n8584), .ZN(n8649) );
  INV_X1 U5997 ( .A(n8590), .ZN(n8662) );
  NAND2_X1 U5998 ( .A1(n5744), .A2(n5743), .ZN(n8668) );
  INV_X1 U5999 ( .A(n8211), .ZN(n8684) );
  NAND2_X1 U6000 ( .A1(n5687), .A2(n5686), .ZN(n8687) );
  AND2_X1 U6001 ( .A1(n4855), .A2(n7823), .ZN(n8510) );
  NAND2_X1 U6002 ( .A1(n5655), .A2(n5654), .ZN(n8697) );
  NAND2_X1 U6003 ( .A1(n5639), .A2(n5638), .ZN(n8703) );
  NAND2_X1 U6004 ( .A1(n4859), .A2(n7936), .ZN(n8533) );
  NAND2_X1 U6005 ( .A1(n5622), .A2(n5621), .ZN(n8709) );
  NAND2_X1 U6006 ( .A1(n5605), .A2(n5604), .ZN(n8716) );
  NAND2_X1 U6007 ( .A1(n5588), .A2(n5587), .ZN(n8228) );
  NAND2_X1 U6008 ( .A1(n5063), .A2(n5582), .ZN(n7715) );
  NAND2_X1 U6009 ( .A1(n7670), .A2(n5581), .ZN(n5063) );
  NAND2_X1 U6010 ( .A1(n4860), .A2(n7920), .ZN(n7719) );
  OR2_X1 U6011 ( .A1(n7669), .A2(n7838), .ZN(n4860) );
  NAND2_X1 U6012 ( .A1(n5573), .A2(n5572), .ZN(n8166) );
  INV_X1 U6013 ( .A(n5858), .ZN(n7700) );
  INV_X1 U6014 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7584) );
  INV_X1 U6015 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7513) );
  INV_X1 U6016 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7466) );
  XNOR2_X1 U6017 ( .A(n5140), .B(n5139), .ZN(n7465) );
  INV_X1 U6018 ( .A(n6805), .ZN(n7856) );
  INV_X1 U6019 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7146) );
  INV_X1 U6020 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6968) );
  INV_X1 U6021 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6908) );
  INV_X1 U6022 ( .A(n5603), .ZN(n8320) );
  INV_X1 U6023 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6658) );
  INV_X1 U6024 ( .A(n7446), .ZN(n6657) );
  INV_X1 U6025 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6642) );
  INV_X1 U6026 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6639) );
  OR2_X1 U6027 ( .A1(n5197), .A2(n5073), .ZN(n9912) );
  NAND2_X1 U6028 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5176), .ZN(n5175) );
  MUX2_X1 U6029 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5179), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5181) );
  AND2_X1 U6030 ( .A1(n6528), .A2(n8830), .ZN(n6529) );
  AND4_X1 U6031 ( .A1(n6164), .A2(n6163), .A3(n6162), .A4(n6161), .ZN(n7371)
         );
  INV_X1 U6032 ( .A(n7271), .ZN(n9767) );
  OAI21_X1 U6033 ( .B1(n8764), .B2(n8763), .A(n4926), .ZN(n8772) );
  AOI21_X1 U6034 ( .B1(n8783), .B2(n8782), .A(n8781), .ZN(n8785) );
  NAND2_X1 U6035 ( .A1(n7354), .A2(n6205), .ZN(n7353) );
  NOR2_X1 U6036 ( .A1(n8738), .A2(n4597), .ZN(n8795) );
  AND4_X1 U6037 ( .A1(n6303), .A2(n6302), .A3(n6301), .A4(n6300), .ZN(n7577)
         );
  NAND2_X1 U6038 ( .A1(n7487), .A2(n7488), .ZN(n4894) );
  NAND2_X1 U6039 ( .A1(n5952), .A2(n5951), .ZN(n9584) );
  AND4_X1 U6040 ( .A1(n6480), .A2(n6479), .A3(n6478), .A4(n6477), .ZN(n8835)
         );
  NAND2_X1 U6041 ( .A1(n7701), .A2(n4903), .ZN(n4902) );
  NOR2_X1 U6042 ( .A1(n4542), .A2(n7752), .ZN(n4903) );
  AND2_X1 U6043 ( .A1(n4603), .A2(n4906), .ZN(n7753) );
  AND2_X1 U6044 ( .A1(n6828), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8837) );
  INV_X1 U6045 ( .A(n9121), .ZN(n9120) );
  INV_X1 U6046 ( .A(n8756), .ZN(n9434) );
  INV_X1 U6047 ( .A(n8787), .ZN(n9449) );
  INV_X1 U6048 ( .A(n7371), .ZN(n9710) );
  XNOR2_X1 U6049 ( .A(n6092), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9179) );
  INV_X1 U6050 ( .A(n4709), .ZN(n9671) );
  INV_X1 U6051 ( .A(n4711), .ZN(n9227) );
  INV_X1 U6052 ( .A(n4713), .ZN(n9267) );
  XNOR2_X1 U6053 ( .A(n9287), .B(n4712), .ZN(n9270) );
  INV_X1 U6054 ( .A(n4716), .ZN(n9310) );
  INV_X1 U6055 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4931) );
  AND2_X1 U6056 ( .A1(n9323), .A2(n9322), .ZN(n9329) );
  NOR2_X1 U6057 ( .A1(n9320), .A2(n9321), .ZN(n9319) );
  OR2_X1 U6058 ( .A1(n9353), .A2(n9351), .ZN(n4724) );
  OAI211_X1 U6059 ( .C1(n9356), .C2(n9672), .A(n9355), .B(n9354), .ZN(n4721)
         );
  CLKBUF_X1 U6060 ( .A(n5995), .Z(n9357) );
  INV_X1 U6061 ( .A(n4720), .ZN(n4719) );
  AOI21_X1 U6062 ( .B1(n9675), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n9358), .ZN(
        n4720) );
  INV_X1 U6063 ( .A(n9367), .ZN(n9366) );
  INV_X1 U6064 ( .A(n5005), .ZN(n9426) );
  INV_X1 U6065 ( .A(n9580), .ZN(n9457) );
  NAND2_X1 U6066 ( .A1(n4756), .A2(n4757), .ZN(n9493) );
  NAND2_X1 U6067 ( .A1(n9647), .A2(n7691), .ZN(n7737) );
  NAND2_X1 U6068 ( .A1(n7475), .A2(n7474), .ZN(n7608) );
  NAND2_X1 U6069 ( .A1(n7476), .A2(n4765), .ZN(n9690) );
  NAND2_X1 U6070 ( .A1(n7303), .A2(n7378), .ZN(n5010) );
  AND2_X1 U6071 ( .A1(n4775), .A2(n8928), .ZN(n7122) );
  NAND2_X1 U6072 ( .A1(n6650), .A2(n4677), .ZN(n4678) );
  INV_X1 U6073 ( .A(n9521), .ZN(n9719) );
  AND2_X2 U6074 ( .A1(n9544), .A2(n9543), .ZN(n9863) );
  INV_X1 U6075 ( .A(n9735), .ZN(n9731) );
  INV_X1 U6076 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5982) );
  XNOR2_X1 U6077 ( .A(n6559), .B(n6558), .ZN(n7791) );
  XNOR2_X1 U6078 ( .A(n5964), .B(n5963), .ZN(n7596) );
  INV_X1 U6079 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5963) );
  INV_X1 U6080 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10489) );
  INV_X1 U6081 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10415) );
  INV_X1 U6082 ( .A(n8919), .ZN(n8881) );
  XNOR2_X1 U6083 ( .A(n5972), .B(n5971), .ZN(n8914) );
  INV_X1 U6084 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10214) );
  INV_X1 U6085 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10403) );
  INV_X1 U6086 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6909) );
  INV_X1 U6087 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6659) );
  INV_X1 U6088 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10483) );
  NAND2_X1 U6089 ( .A1(n4798), .A2(n5493), .ZN(n4707) );
  NAND2_X1 U6090 ( .A1(n6925), .A2(n6924), .ZN(n6928) );
  NOR2_X1 U6091 ( .A1(n7338), .A2(n7337), .ZN(n7336) );
  OR2_X1 U6092 ( .A1(n8379), .A2(n4617), .ZN(P2_U3199) );
  OAI21_X1 U6093 ( .B1(n8381), .B2(n9948), .A(n4618), .ZN(n4617) );
  AOI21_X1 U6094 ( .B1(n8380), .B2(n9964), .A(n8378), .ZN(n4618) );
  AND2_X1 U6095 ( .A1(n5001), .A2(n4999), .ZN(n8397) );
  OAI21_X1 U6096 ( .B1(n8393), .B2(n4534), .A(n5002), .ZN(n5001) );
  NAND2_X1 U6098 ( .A1(n4620), .A2(n4619), .ZN(P2_U3207) );
  AOI21_X1 U6099 ( .B1(n8432), .B2(n9977), .A(n8431), .ZN(n4619) );
  INV_X1 U6100 ( .A(n8430), .ZN(n4620) );
  AOI21_X1 U6101 ( .B1(n6584), .B2(n8629), .A(n6589), .ZN(n6590) );
  AND2_X1 U6102 ( .A1(n5894), .A2(n5089), .ZN(n5895) );
  NAND2_X1 U6103 ( .A1(n8581), .A2(n5090), .ZN(n8583) );
  AND2_X1 U6104 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  NAND2_X1 U6105 ( .A1(n4611), .A2(n4610), .ZN(n8657) );
  NAND2_X1 U6106 ( .A1(n10049), .A2(n8654), .ZN(n4610) );
  AOI21_X1 U6107 ( .B1(n4939), .B2(n6591), .A(n4935), .ZN(n4934) );
  INV_X1 U6108 ( .A(n4939), .ZN(n4938) );
  NAND2_X1 U6109 ( .A1(n4722), .A2(n4718), .ZN(P1_U3262) );
  NAND2_X1 U6110 ( .A1(n4723), .A2(n6726), .ZN(n4722) );
  AOI21_X1 U6111 ( .B1(n4721), .B2(n9357), .A(n4719), .ZN(n4718) );
  OAI21_X1 U6112 ( .B1(n9352), .B2(n9672), .A(n4724), .ZN(n4723) );
  INV_X1 U6113 ( .A(n4768), .ZN(n7781) );
  OAI21_X1 U6114 ( .B1(n9556), .B2(n9730), .A(n4769), .ZN(n4768) );
  AOI21_X1 U6115 ( .B1(n9553), .B2(n9726), .A(n7780), .ZN(n4769) );
  NAND2_X1 U6116 ( .A1(n9584), .A2(n9462), .ZN(n4524) );
  OR2_X1 U6117 ( .A1(n4961), .A2(n5097), .ZN(n4525) );
  NAND2_X1 U6118 ( .A1(n6341), .A2(n6340), .ZN(n4926) );
  INV_X1 U6119 ( .A(n4926), .ZN(n4920) );
  NOR2_X1 U6120 ( .A1(n6530), .A2(n6527), .ZN(n8830) );
  AND2_X1 U6121 ( .A1(n6355), .A2(n6354), .ZN(n4526) );
  OR2_X1 U6122 ( .A1(n5570), .A2(n4819), .ZN(n4527) );
  OR2_X1 U6123 ( .A1(n9575), .A2(n8757), .ZN(n9091) );
  OR2_X1 U6124 ( .A1(n8082), .A2(n5723), .ZN(n4528) );
  AND2_X1 U6125 ( .A1(n4847), .A2(n8406), .ZN(n4529) );
  OR2_X1 U6126 ( .A1(n5528), .A2(n5207), .ZN(n4530) );
  AND2_X1 U6127 ( .A1(n4564), .A2(n7920), .ZN(n4531) );
  OR2_X1 U6128 ( .A1(n4526), .A2(n8814), .ZN(n4532) );
  NAND2_X1 U6129 ( .A1(n6810), .A2(n4879), .ZN(n5876) );
  INV_X1 U6130 ( .A(n7474), .ZN(n5017) );
  AND2_X1 U6131 ( .A1(n4527), .A2(n5583), .ZN(n4533) );
  NAND2_X1 U6132 ( .A1(n6425), .A2(n6424), .ZN(n9575) );
  INV_X1 U6133 ( .A(n4760), .ZN(n4759) );
  NAND2_X1 U6134 ( .A1(n8967), .A2(n9058), .ZN(n4760) );
  AND2_X1 U6135 ( .A1(n8395), .A2(n8394), .ZN(n4534) );
  OR2_X1 U6136 ( .A1(n9575), .A2(n9461), .ZN(n4535) );
  AND2_X1 U6137 ( .A1(n4967), .A2(n8435), .ZN(n4536) );
  AND2_X1 U6138 ( .A1(n9603), .A2(n9137), .ZN(n4537) );
  AND2_X1 U6139 ( .A1(n4704), .A2(n4703), .ZN(n4538) );
  NAND2_X1 U6140 ( .A1(n8844), .A2(n8843), .ZN(n9359) );
  INV_X1 U6141 ( .A(n9359), .ZN(n9547) );
  NAND2_X1 U6142 ( .A1(n7397), .A2(n4726), .ZN(n4730) );
  INV_X1 U6143 ( .A(n5026), .ZN(n5034) );
  INV_X1 U6144 ( .A(n9116), .ZN(n4644) );
  INV_X1 U6145 ( .A(n5236), .ZN(n8025) );
  NAND2_X1 U6146 ( .A1(n6316), .A2(n6315), .ZN(n7609) );
  INV_X1 U6147 ( .A(n7526), .ZN(n4741) );
  NAND2_X1 U6148 ( .A1(n7320), .A2(n4975), .ZN(n7422) );
  INV_X1 U6149 ( .A(n8124), .ZN(n4952) );
  NAND2_X1 U6150 ( .A1(n4886), .A2(n6089), .ZN(n7009) );
  NAND2_X1 U6151 ( .A1(n6153), .A2(n6152), .ZN(n7106) );
  AND2_X4 U6152 ( .A1(n6650), .A2(n7798), .ZN(n6066) );
  INV_X1 U6153 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5977) );
  CLKBUF_X1 U6154 ( .A(n5382), .Z(n9985) );
  AND2_X1 U6155 ( .A1(n6806), .A2(n8021), .ZN(n4539) );
  INV_X1 U6156 ( .A(n4891), .ZN(n6046) );
  NAND2_X1 U6157 ( .A1(n6019), .A2(n7076), .ZN(n6083) );
  OR2_X1 U6158 ( .A1(n5242), .A2(n9896), .ZN(n4540) );
  AND2_X1 U6159 ( .A1(n4949), .A2(n8125), .ZN(n4541) );
  AND2_X1 U6160 ( .A1(n4905), .A2(n4904), .ZN(n4542) );
  OAI21_X1 U6161 ( .B1(n9474), .B2(n5027), .A(n4524), .ZN(n5026) );
  AND2_X1 U6162 ( .A1(n8584), .A2(n8435), .ZN(n4543) );
  AND2_X1 U6163 ( .A1(n4692), .A2(n4691), .ZN(n4544) );
  OR2_X1 U6164 ( .A1(n9515), .A2(n9136), .ZN(n8967) );
  XNOR2_X1 U6165 ( .A(n8144), .B(n8101), .ZN(n7820) );
  INV_X1 U6166 ( .A(n7820), .ZN(n5839) );
  OR2_X1 U6167 ( .A1(n6313), .A2(n5092), .ZN(n4545) );
  OR2_X1 U6168 ( .A1(n8716), .A2(n8548), .ZN(n4546) );
  AND2_X1 U6169 ( .A1(n5046), .A2(n5050), .ZN(n4547) );
  INV_X1 U6170 ( .A(n8984), .ZN(n4658) );
  AND2_X1 U6171 ( .A1(n6580), .A2(n9981), .ZN(n4548) );
  AND2_X1 U6172 ( .A1(n5032), .A2(n5034), .ZN(n4549) );
  NOR4_X1 U6173 ( .A1(n7847), .A2(n8013), .A3(n8002), .A4(n7846), .ZN(n4550)
         );
  NAND2_X1 U6174 ( .A1(n5997), .A2(n5996), .ZN(n9603) );
  INV_X1 U6175 ( .A(n9603), .ZN(n4742) );
  XNOR2_X1 U6176 ( .A(n8642), .B(n8280), .ZN(n8406) );
  NAND2_X1 U6177 ( .A1(n5073), .A2(n5074), .ZN(n4551) );
  INV_X1 U6178 ( .A(n8814), .ZN(n4928) );
  AND2_X1 U6179 ( .A1(n8642), .A2(n8280), .ZN(n4552) );
  NAND2_X1 U6180 ( .A1(n6259), .A2(n6258), .ZN(n9031) );
  NAND2_X1 U6181 ( .A1(n6332), .A2(n6331), .ZN(n8769) );
  AND2_X1 U6182 ( .A1(n7939), .A2(n8012), .ZN(n4553) );
  INV_X1 U6183 ( .A(n4832), .ZN(n5145) );
  NAND2_X1 U6184 ( .A1(n6344), .A2(n6343), .ZN(n8778) );
  NOR2_X1 U6185 ( .A1(n9059), .A2(n9116), .ZN(n4554) );
  NAND2_X1 U6186 ( .A1(n5716), .A2(n5715), .ZN(n8082) );
  AND2_X1 U6187 ( .A1(n4901), .A2(n6311), .ZN(n4555) );
  AND2_X1 U6188 ( .A1(n8649), .A2(n8435), .ZN(n7988) );
  NAND2_X1 U6189 ( .A1(n5778), .A2(n5777), .ZN(n8655) );
  INV_X1 U6190 ( .A(n4630), .ZN(n7911) );
  NAND2_X1 U6191 ( .A1(n10043), .A2(n8287), .ZN(n4630) );
  NAND2_X1 U6192 ( .A1(n6362), .A2(n6361), .ZN(n9608) );
  AND4_X1 U6193 ( .A1(n5460), .A2(n5459), .A3(n5458), .A4(n5457), .ZN(n7331)
         );
  INV_X1 U6194 ( .A(n7331), .ZN(n8290) );
  AND2_X1 U6195 ( .A1(n4919), .A2(n6372), .ZN(n4556) );
  OR2_X1 U6196 ( .A1(n8655), .A2(n8446), .ZN(n7987) );
  INV_X1 U6197 ( .A(n4965), .ZN(n4964) );
  OR2_X1 U6198 ( .A1(n8095), .A2(n4966), .ZN(n4965) );
  OR2_X1 U6199 ( .A1(n6784), .A2(n6767), .ZN(n4557) );
  OR2_X1 U6200 ( .A1(n6440), .A2(n6423), .ZN(n4558) );
  NAND2_X1 U6201 ( .A1(n9955), .A2(n5206), .ZN(n5208) );
  INV_X1 U6202 ( .A(n6328), .ZN(n4905) );
  OR2_X1 U6203 ( .A1(n8211), .A2(n8505), .ZN(n5709) );
  AND2_X1 U6204 ( .A1(n6292), .A2(n6291), .ZN(n4559) );
  INV_X1 U6205 ( .A(n7899), .ZN(n4688) );
  AND2_X1 U6206 ( .A1(n4756), .A2(n4753), .ZN(n4560) );
  INV_X1 U6207 ( .A(n4857), .ZN(n4856) );
  NAND2_X1 U6208 ( .A1(n8503), .A2(n8501), .ZN(n4857) );
  NOR2_X1 U6209 ( .A1(n9031), .A2(n9143), .ZN(n4561) );
  OR2_X1 U6210 ( .A1(n6576), .A2(n9930), .ZN(n4562) );
  INV_X1 U6211 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5352) );
  AND4_X1 U6212 ( .A1(n5114), .A2(n5113), .A3(n5228), .A4(n5132), .ZN(n4563)
         );
  OR2_X1 U6213 ( .A1(n8228), .A2(n8562), .ZN(n4564) );
  NOR2_X1 U6214 ( .A1(n5200), .A2(n5249), .ZN(n4565) );
  OR2_X1 U6215 ( .A1(n9430), .A2(n8787), .ZN(n4566) );
  INV_X1 U6216 ( .A(n5097), .ZN(n4968) );
  INV_X1 U6217 ( .A(n4727), .ZN(n4726) );
  NAND2_X1 U6218 ( .A1(n4729), .A2(n4728), .ZN(n4727) );
  AND2_X1 U6219 ( .A1(n5506), .A2(SI_7_), .ZN(n4567) );
  INV_X1 U6220 ( .A(n4754), .ZN(n4753) );
  NAND2_X1 U6221 ( .A1(n4755), .A2(n4757), .ZN(n4754) );
  AND2_X1 U6222 ( .A1(n5585), .A2(SI_12_), .ZN(n4568) );
  NOR2_X1 U6223 ( .A1(n9580), .A2(n9470), .ZN(n4569) );
  AND2_X1 U6224 ( .A1(n4912), .A2(n4558), .ZN(n4570) );
  INV_X1 U6225 ( .A(n4924), .ZN(n4923) );
  OAI21_X1 U6226 ( .B1(n8773), .B2(n4526), .A(n4925), .ZN(n4924) );
  INV_X1 U6227 ( .A(n4734), .ZN(n9386) );
  NOR2_X1 U6228 ( .A1(n9385), .A2(n9549), .ZN(n4734) );
  AND2_X1 U6229 ( .A1(n9087), .A2(n9446), .ZN(n9460) );
  OR2_X1 U6230 ( .A1(n5052), .A2(n4543), .ZN(n4571) );
  INV_X1 U6231 ( .A(n7768), .ZN(n5035) );
  INV_X1 U6232 ( .A(n4847), .ZN(n4844) );
  NOR2_X1 U6233 ( .A1(n7988), .A2(n7979), .ZN(n4847) );
  NAND2_X1 U6234 ( .A1(n4672), .A2(n9547), .ZN(n4572) );
  NAND2_X1 U6235 ( .A1(n8481), .A2(n5072), .ZN(n4573) );
  INV_X1 U6236 ( .A(n8763), .ZN(n4927) );
  INV_X1 U6237 ( .A(n4782), .ZN(n4781) );
  NAND2_X1 U6238 ( .A1(n5200), .A2(n5249), .ZN(n4782) );
  NAND2_X1 U6239 ( .A1(n8144), .A2(n8410), .ZN(n4574) );
  INV_X1 U6240 ( .A(n6209), .ZN(n4890) );
  OR2_X1 U6241 ( .A1(n7609), .A2(n5017), .ZN(n4575) );
  INV_X1 U6242 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9626) );
  AND4_X1 U6243 ( .A1(n4875), .A2(n5173), .A3(n4874), .A4(n4876), .ZN(n4576)
         );
  AND2_X1 U6244 ( .A1(n9070), .A2(n4648), .ZN(n4577) );
  AND2_X1 U6245 ( .A1(n5057), .A2(n4546), .ZN(n4578) );
  INV_X1 U6246 ( .A(n7977), .ZN(n8423) );
  AND2_X1 U6247 ( .A1(n4845), .A2(n7982), .ZN(n7977) );
  AND2_X1 U6248 ( .A1(n8439), .A2(n5051), .ZN(n4579) );
  OR2_X1 U6249 ( .A1(n7939), .A2(n8012), .ZN(n4580) );
  INV_X1 U6250 ( .A(n9554), .ZN(n9380) );
  NAND2_X1 U6251 ( .A1(n6488), .A2(n6487), .ZN(n9554) );
  AND2_X1 U6252 ( .A1(n7900), .A2(n8012), .ZN(n4581) );
  AND2_X1 U6253 ( .A1(n4743), .A2(n4742), .ZN(n4582) );
  NOR2_X1 U6254 ( .A1(n4910), .A2(n4914), .ZN(n4583) );
  AND2_X1 U6255 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4584) );
  AND2_X1 U6256 ( .A1(n4817), .A2(n5583), .ZN(n4585) );
  AND2_X1 U6257 ( .A1(n6926), .A2(n6924), .ZN(n4586) );
  AND2_X1 U6258 ( .A1(n4917), .A2(n4915), .ZN(n4587) );
  OR2_X1 U6259 ( .A1(n4532), .A2(n4916), .ZN(n4588) );
  INV_X1 U6260 ( .A(n8089), .ZN(n4969) );
  NOR2_X1 U6261 ( .A1(n9457), .A2(n8809), .ZN(n4589) );
  INV_X1 U6262 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5086) );
  NAND2_X1 U6263 ( .A1(n8289), .A2(n7321), .ZN(n4590) );
  INV_X1 U6264 ( .A(n5226), .ZN(n4791) );
  AND2_X1 U6265 ( .A1(n5467), .A2(n5468), .ZN(n4591) );
  INV_X1 U6266 ( .A(n9730), .ZN(n9534) );
  NAND2_X1 U6267 ( .A1(n8524), .A2(n7822), .ZN(n4855) );
  INV_X1 U6268 ( .A(n9139), .ZN(n5025) );
  INV_X1 U6269 ( .A(n8253), .ZN(n4967) );
  NAND2_X1 U6270 ( .A1(n7605), .A2(n4745), .ZN(n4592) );
  INV_X1 U6271 ( .A(n7662), .ZN(n6716) );
  OR2_X1 U6272 ( .A1(n5966), .A2(n9626), .ZN(n6342) );
  NAND2_X1 U6273 ( .A1(n5010), .A2(n7381), .ZN(n7395) );
  NAND2_X1 U6274 ( .A1(n4894), .A2(n6274), .ZN(n7573) );
  INV_X1 U6275 ( .A(n5528), .ZN(n7196) );
  AND2_X1 U6276 ( .A1(n5170), .A2(n5209), .ZN(n5528) );
  AND2_X1 U6277 ( .A1(n6778), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4593) );
  AND2_X1 U6278 ( .A1(n7343), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4594) );
  INV_X1 U6279 ( .A(n9072), .ZN(n4752) );
  INV_X1 U6280 ( .A(n7958), .ZN(n4852) );
  INV_X1 U6281 ( .A(n6678), .ZN(n5288) );
  INV_X1 U6282 ( .A(n4977), .ZN(n5149) );
  AND2_X1 U6283 ( .A1(n8512), .A2(n4856), .ZN(n4595) );
  NOR2_X1 U6284 ( .A1(n7436), .A2(n5220), .ZN(n4596) );
  NOR2_X1 U6285 ( .A1(n9509), .A2(n9593), .ZN(n9478) );
  AND4_X1 U6286 ( .A1(n6431), .A2(n6430), .A3(n6429), .A4(n6428), .ZN(n8757)
         );
  INV_X1 U6287 ( .A(n6591), .ZN(n4944) );
  AND2_X1 U6288 ( .A1(n6374), .A2(n6375), .ZN(n4597) );
  NAND2_X1 U6289 ( .A1(n6476), .A2(n6475), .ZN(n9560) );
  AND2_X1 U6290 ( .A1(n6596), .A2(n6597), .ZN(n4598) );
  AND2_X1 U6291 ( .A1(n5724), .A2(SI_21_), .ZN(n4599) );
  OAI21_X1 U6292 ( .B1(n8772), .B2(n4526), .A(n4923), .ZN(n4929) );
  OR2_X1 U6293 ( .A1(n5648), .A2(SI_16_), .ZN(n4600) );
  AND2_X1 U6294 ( .A1(n4807), .A2(n4806), .ZN(n4601) );
  NAND3_X1 U6295 ( .A1(n5039), .A2(n5038), .A3(n4931), .ZN(n4602) );
  AND2_X1 U6296 ( .A1(n5172), .A2(n5203), .ZN(n5249) );
  INV_X1 U6297 ( .A(n5249), .ZN(n9930) );
  AND2_X1 U6298 ( .A1(n7702), .A2(n4905), .ZN(n4603) );
  AND2_X1 U6299 ( .A1(n8061), .A2(n8060), .ZN(n4604) );
  AND2_X1 U6300 ( .A1(n5256), .A2(n4985), .ZN(n4605) );
  AND2_X1 U6301 ( .A1(n4948), .A2(n8213), .ZN(n4606) );
  OR2_X1 U6302 ( .A1(n7662), .A2(n7675), .ZN(n4607) );
  INV_X1 U6303 ( .A(n8731), .ZN(n4913) );
  NAND2_X1 U6304 ( .A1(n6726), .A2(n8914), .ZN(n6526) );
  NAND2_X1 U6305 ( .A1(n6913), .A2(n7824), .ZN(n6912) );
  AND3_X1 U6306 ( .A1(n6323), .A2(n6322), .A3(n6321), .ZN(n9694) );
  INV_X1 U6307 ( .A(n9694), .ZN(n5016) );
  XNOR2_X1 U6308 ( .A(n5957), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U6309 ( .A1(n7367), .A2(n7368), .ZN(n7354) );
  NAND2_X1 U6310 ( .A1(n6296), .A2(n6295), .ZN(n9699) );
  INV_X1 U6311 ( .A(n9699), .ZN(n4728) );
  INV_X1 U6312 ( .A(n9041), .ZN(n4766) );
  NAND2_X1 U6313 ( .A1(n5480), .A2(n5481), .ZN(n7258) );
  NAND2_X1 U6314 ( .A1(n6912), .A2(n5436), .ZN(n6970) );
  INV_X2 U6315 ( .A(n10049), .ZN(n10048) );
  AND2_X1 U6316 ( .A1(n5907), .A2(n5906), .ZN(n10049) );
  INV_X1 U6317 ( .A(n8212), .ZN(n4951) );
  AND2_X1 U6318 ( .A1(n4738), .A2(n4737), .ZN(n4608) );
  INV_X1 U6319 ( .A(n9948), .ZN(n5002) );
  INV_X1 U6320 ( .A(n9281), .ZN(n4712) );
  AND4_X2 U6321 ( .A1(n5875), .A2(n5919), .A3(n5898), .A4(n5874), .ZN(n10064)
         );
  INV_X1 U6322 ( .A(n9981), .ZN(n8561) );
  INV_X1 U6323 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U6324 ( .A1(n6525), .A2(n9357), .ZN(n9116) );
  INV_X1 U6325 ( .A(n9779), .ZN(n4740) );
  NAND2_X1 U6326 ( .A1(n7184), .A2(n7101), .ZN(n7098) );
  INV_X1 U6327 ( .A(n7098), .ZN(n4731) );
  AND2_X1 U6328 ( .A1(n4990), .A2(n4540), .ZN(n4609) );
  INV_X1 U6329 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6523) );
  XNOR2_X1 U6330 ( .A(n4976), .B(n5134), .ZN(n7850) );
  INV_X1 U6331 ( .A(n7850), .ZN(n5901) );
  INV_X1 U6332 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5967) );
  INV_X1 U6333 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4638) );
  NAND2_X1 U6334 ( .A1(n5087), .A2(n5496), .ZN(n7408) );
  NAND2_X1 U6335 ( .A1(n4805), .A2(n4802), .ZN(n5754) );
  OAI21_X1 U6336 ( .B1(n5665), .B2(n5664), .A(n5663), .ZN(n5680) );
  NAND2_X1 U6337 ( .A1(n5391), .A2(n5390), .ZN(n4746) );
  NOR2_X2 U6338 ( .A1(n8739), .A2(n8740), .ZN(n8738) );
  OAI21_X2 U6339 ( .B1(n8764), .B2(n4921), .A(n4556), .ZN(n8813) );
  NAND2_X1 U6340 ( .A1(n7107), .A2(n6172), .ZN(n6189) );
  OAI21_X2 U6341 ( .B1(n9439), .B2(n4615), .A(n4535), .ZN(n5005) );
  OAI21_X2 U6342 ( .B1(n7764), .B2(n7763), .A(n7765), .ZN(n9518) );
  NAND2_X1 U6343 ( .A1(n7552), .A2(n7551), .ZN(n7619) );
  NAND2_X1 U6344 ( .A1(n6925), .A2(n4586), .ZN(n6952) );
  NAND3_X2 U6345 ( .A1(n5073), .A2(n5074), .A3(n5139), .ZN(n5118) );
  INV_X1 U6346 ( .A(n6811), .ZN(n4946) );
  AOI21_X2 U6347 ( .B1(n8233), .B2(n8090), .A(n8089), .ZN(n8201) );
  XNOR2_X1 U6348 ( .A(n5221), .B(n8305), .ZN(n8303) );
  NOR2_X2 U6349 ( .A1(n7658), .A2(n4616), .ZN(n5221) );
  NOR2_X2 U6350 ( .A1(n8347), .A2(n4614), .ZN(n5225) );
  NOR2_X1 U6351 ( .A1(n8371), .A2(n8617), .ZN(n8373) );
  NOR2_X1 U6352 ( .A1(n6679), .A2(n5183), .ZN(n9873) );
  AOI21_X1 U6353 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n4513), .A(n9872), .ZN(
        n5188) );
  OAI211_X1 U6354 ( .C1(n6205), .C2(n4890), .A(n6233), .B(n4887), .ZN(n6250)
         );
  NAND2_X1 U6355 ( .A1(n5012), .A2(n5011), .ZN(n7610) );
  NAND2_X1 U6356 ( .A1(n5067), .A2(n5064), .ZN(n8457) );
  NOR2_X1 U6357 ( .A1(n8337), .A2(n8623), .ZN(n8336) );
  XNOR2_X1 U6358 ( .A(n5223), .B(n5620), .ZN(n8337) );
  NOR2_X1 U6359 ( .A1(n5188), .A2(n6670), .ZN(n6703) );
  INV_X1 U6360 ( .A(n4833), .ZN(n5122) );
  NAND3_X1 U6361 ( .A1(n4705), .A2(n7918), .A3(n4622), .ZN(n4621) );
  NAND3_X1 U6362 ( .A1(n4625), .A2(n4624), .A3(n8468), .ZN(n4623) );
  OAI21_X2 U6363 ( .B1(n4628), .B2(n4627), .A(n8000), .ZN(n8004) );
  OAI211_X1 U6364 ( .C1(n9086), .C2(n4644), .A(n9089), .B(n4639), .ZN(n9093)
         );
  NOR2_X2 U6365 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6043) );
  NAND3_X1 U6366 ( .A1(n4651), .A2(n4649), .A3(n4577), .ZN(n9080) );
  NAND2_X1 U6367 ( .A1(n8981), .A2(n8980), .ZN(n8995) );
  NAND3_X1 U6368 ( .A1(n8981), .A2(n4656), .A3(n4657), .ZN(n4655) );
  NAND2_X1 U6369 ( .A1(n9115), .A2(n4663), .ZN(n4662) );
  AND2_X1 U6370 ( .A1(n9114), .A2(n9113), .ZN(n4672) );
  NAND3_X1 U6371 ( .A1(n9101), .A2(n4676), .A3(n4674), .ZN(n4673) );
  NAND2_X2 U6372 ( .A1(n6764), .A2(n7793), .ZN(n6650) );
  OAI21_X1 U6373 ( .B1(n6606), .B2(n7798), .A(n4679), .ZN(n4677) );
  OAI21_X2 U6374 ( .B1(n6650), .B2(n6008), .A(n4678), .ZN(n6016) );
  OAI21_X1 U6375 ( .B1(n7798), .B2(n4683), .A(n4682), .ZN(n5392) );
  NAND2_X4 U6376 ( .A1(n5369), .A2(n5370), .ZN(n7798) );
  AND2_X2 U6377 ( .A1(n4696), .A2(n4695), .ZN(n4694) );
  AND2_X2 U6378 ( .A1(n4702), .A2(n4701), .ZN(n4700) );
  INV_X1 U6379 ( .A(n8005), .ZN(n4704) );
  NAND2_X1 U6380 ( .A1(n7397), .A2(n4725), .ZN(n7604) );
  INV_X1 U6381 ( .A(n4730), .ZN(n7481) );
  NAND2_X1 U6382 ( .A1(n5411), .A2(n5410), .ZN(n5414) );
  MUX2_X1 U6383 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n7798), .Z(n5412) );
  NAND2_X1 U6384 ( .A1(n4746), .A2(n5393), .ZN(n5411) );
  NAND3_X1 U6385 ( .A1(n4775), .A2(n8890), .A3(n8928), .ZN(n7307) );
  NAND3_X1 U6386 ( .A1(n7121), .A2(n4657), .A3(n7119), .ZN(n4775) );
  NAND2_X1 U6387 ( .A1(n7119), .A2(n8984), .ZN(n7243) );
  OR2_X1 U6388 ( .A1(n7120), .A2(n8996), .ZN(n8918) );
  NAND2_X1 U6389 ( .A1(n5199), .A2(n4779), .ZN(n4778) );
  NAND2_X1 U6390 ( .A1(n5199), .A2(n5198), .ZN(n9906) );
  INV_X1 U6391 ( .A(n5193), .ZN(n4787) );
  INV_X1 U6392 ( .A(n5192), .ZN(n4788) );
  OR2_X1 U6393 ( .A1(n5226), .A2(n8373), .ZN(n4793) );
  OAI22_X1 U6394 ( .A1(n8373), .A2(n4790), .B1(n4792), .B2(n5232), .ZN(n5234)
         );
  INV_X1 U6395 ( .A(n4793), .ZN(n8384) );
  NAND2_X1 U6396 ( .A1(n5491), .A2(n4799), .ZN(n4796) );
  NAND2_X1 U6397 ( .A1(n4796), .A2(n4797), .ZN(n5524) );
  NAND2_X1 U6398 ( .A1(n5491), .A2(n5490), .ZN(n4798) );
  MUX2_X1 U6399 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7798), .Z(n5446) );
  NAND2_X1 U6400 ( .A1(n5712), .A2(n4601), .ZN(n4805) );
  NAND2_X1 U6401 ( .A1(n5534), .A2(n4585), .ZN(n4816) );
  NAND2_X1 U6402 ( .A1(n5534), .A2(n4821), .ZN(n4820) );
  NAND2_X1 U6403 ( .A1(n5534), .A2(n5533), .ZN(n5554) );
  NAND2_X1 U6404 ( .A1(n5618), .A2(n4827), .ZN(n4823) );
  NAND2_X1 U6405 ( .A1(n5618), .A2(n5617), .ZN(n5635) );
  NAND2_X1 U6406 ( .A1(n4831), .A2(n8032), .ZN(n6587) );
  OAI211_X1 U6407 ( .C1(n4831), .C2(n10062), .A(n4829), .B(n6590), .ZN(
        P2_U3488) );
  NAND2_X1 U6408 ( .A1(n4830), .A2(n10064), .ZN(n4829) );
  INV_X1 U6409 ( .A(n8032), .ZN(n4830) );
  NAND2_X1 U6410 ( .A1(n6583), .A2(n6582), .ZN(n4831) );
  INV_X1 U6411 ( .A(n5118), .ZN(n5120) );
  NAND2_X1 U6412 ( .A1(n4833), .A2(n5086), .ZN(n4832) );
  NOR2_X2 U6413 ( .A1(n5118), .A2(n4834), .ZN(n4833) );
  NAND2_X1 U6414 ( .A1(n8438), .A2(n4529), .ZN(n4842) );
  INV_X1 U6415 ( .A(n8438), .ZN(n4836) );
  NAND2_X1 U6416 ( .A1(n4846), .A2(n4845), .ZN(n4843) );
  AOI21_X1 U6417 ( .B1(n8438), .B2(n7984), .A(n5887), .ZN(n8420) );
  INV_X1 U6418 ( .A(n7988), .ZN(n4845) );
  NAND2_X1 U6419 ( .A1(n8524), .A2(n4849), .ZN(n4848) );
  NAND2_X1 U6420 ( .A1(n4859), .A2(n4858), .ZN(n5884) );
  NAND2_X1 U6421 ( .A1(n7669), .A2(n4531), .ZN(n4863) );
  NAND2_X1 U6422 ( .A1(n6973), .A2(n7879), .ZN(n7208) );
  INV_X1 U6423 ( .A(n7879), .ZN(n4872) );
  NOR2_X1 U6424 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4873) );
  NAND2_X2 U6425 ( .A1(n5374), .A2(n6605), .ZN(n7803) );
  NAND2_X1 U6426 ( .A1(n7863), .A2(n7864), .ZN(n9980) );
  AOI21_X2 U6427 ( .B1(n6662), .B2(n5189), .A(n6701), .ZN(n6706) );
  AOI21_X2 U6428 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8320), .A(n8312), .ZN(
        n5223) );
  NOR2_X1 U6429 ( .A1(n5222), .A2(n8301), .ZN(n8314) );
  NOR2_X1 U6430 ( .A1(n5224), .A2(n8336), .ZN(n8349) );
  NAND2_X1 U6431 ( .A1(n6153), .A2(n4880), .ZN(n7107) );
  AND2_X1 U6432 ( .A1(n6171), .A2(n6152), .ZN(n4880) );
  NAND2_X1 U6433 ( .A1(n6359), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U6434 ( .A1(n5976), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4881) );
  NAND2_X1 U6435 ( .A1(n5976), .A2(n4584), .ZN(n4882) );
  INV_X1 U6436 ( .A(n4884), .ZN(n4883) );
  NAND3_X1 U6437 ( .A1(n4886), .A2(n6089), .A3(n6109), .ZN(n7010) );
  NAND2_X1 U6438 ( .A1(n7367), .A2(n4888), .ZN(n4887) );
  OAI21_X1 U6439 ( .B1(n4891), .B2(n9738), .A(n6014), .ZN(n6015) );
  OAI21_X2 U6440 ( .B1(n5979), .B2(n5980), .A(n6019), .ZN(n4891) );
  NOR2_X1 U6441 ( .A1(n4910), .A2(n4913), .ZN(n4907) );
  AOI21_X2 U6442 ( .B1(n4911), .B2(n4908), .A(n4570), .ZN(n8754) );
  NOR2_X1 U6443 ( .A1(n6406), .A2(n4909), .ZN(n4908) );
  NAND2_X1 U6444 ( .A1(n8813), .A2(n4587), .ZN(n8739) );
  AND3_X1 U6445 ( .A1(n5039), .A2(n4932), .A3(n5038), .ZN(n5966) );
  NAND2_X1 U6446 ( .A1(n5039), .A2(n5038), .ZN(n6313) );
  NAND2_X1 U6447 ( .A1(n8828), .A2(n4937), .ZN(n4933) );
  NOR2_X1 U6448 ( .A1(n8828), .A2(n6471), .ZN(n8825) );
  OAI211_X1 U6449 ( .C1(n8828), .C2(n4938), .A(n4933), .B(n4934), .ZN(P1_U3214) );
  NOR2_X2 U6450 ( .A1(n8825), .A2(n4945), .ZN(n6593) );
  NAND2_X1 U6451 ( .A1(n4946), .A2(n9985), .ZN(n6812) );
  NAND2_X1 U6452 ( .A1(n4947), .A2(n4606), .ZN(n8147) );
  NAND2_X1 U6453 ( .A1(n8123), .A2(n4950), .ZN(n4947) );
  NAND2_X1 U6454 ( .A1(n8233), .A2(n4956), .ZN(n4955) );
  OAI21_X1 U6455 ( .B1(n8233), .B2(n4525), .A(n4956), .ZN(n8255) );
  NAND2_X1 U6456 ( .A1(n8053), .A2(n4970), .ZN(n8106) );
  NAND2_X1 U6457 ( .A1(n8106), .A2(n8107), .ZN(n8057) );
  NOR2_X2 U6459 ( .A1(n8358), .A2(n4978), .ZN(n5264) );
  INV_X1 U6460 ( .A(n4985), .ZN(n7431) );
  NAND2_X1 U6461 ( .A1(n5243), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4991) );
  NAND2_X1 U6462 ( .A1(n4995), .A2(n4996), .ZN(n5257) );
  NAND2_X1 U6463 ( .A1(n7191), .A2(n4997), .ZN(n4995) );
  OAI21_X2 U6464 ( .B1(n9518), .B2(n4537), .A(n7766), .ZN(n9503) );
  NAND2_X1 U6465 ( .A1(n7379), .A2(n5006), .ZN(n5008) );
  NAND2_X1 U6466 ( .A1(n5008), .A2(n5007), .ZN(n7469) );
  NAND2_X1 U6467 ( .A1(n7475), .A2(n5013), .ZN(n5012) );
  NAND2_X1 U6468 ( .A1(n9490), .A2(n5029), .ZN(n5032) );
  NOR2_X2 U6469 ( .A1(n5936), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5038) );
  INV_X2 U6470 ( .A(n6155), .ZN(n5039) );
  INV_X1 U6471 ( .A(n5092), .ZN(n5037) );
  NAND4_X1 U6472 ( .A1(n5037), .A2(n5949), .A3(n5038), .A4(n5039), .ZN(n5945)
         );
  NAND2_X1 U6473 ( .A1(n8433), .A2(n8439), .ZN(n5049) );
  NAND2_X1 U6474 ( .A1(n8433), .A2(n4579), .ZN(n5047) );
  INV_X1 U6475 ( .A(n5052), .ZN(n5048) );
  NAND2_X1 U6476 ( .A1(n7670), .A2(n4578), .ZN(n5056) );
  NAND3_X1 U6477 ( .A1(n5057), .A2(n5060), .A3(n4546), .ZN(n5055) );
  NAND2_X1 U6478 ( .A1(n8490), .A2(n5068), .ZN(n5067) );
  NAND3_X1 U6479 ( .A1(n5070), .A2(n5069), .A3(n5071), .ZN(n5066) );
  INV_X1 U6480 ( .A(n5112), .ZN(n5075) );
  NAND2_X1 U6481 ( .A1(n6912), .A2(n5080), .ZN(n5078) );
  NAND2_X1 U6482 ( .A1(n5078), .A2(n5077), .ZN(n5478) );
  NAND3_X1 U6483 ( .A1(n5481), .A2(n5480), .A3(n4590), .ZN(n5087) );
  NAND2_X1 U6484 ( .A1(n5125), .A2(n5124), .ZN(n5126) );
  NAND2_X2 U6485 ( .A1(n7036), .A2(n7035), .ZN(n7320) );
  NAND2_X1 U6486 ( .A1(n6250), .A2(n6249), .ZN(n6255) );
  NAND2_X1 U6487 ( .A1(n8429), .A2(n8428), .ZN(n8646) );
  NAND2_X1 U6488 ( .A1(n5921), .A2(n10048), .ZN(n5912) );
  NAND2_X1 U6489 ( .A1(n5921), .A2(n10064), .ZN(n5896) );
  NOR2_X1 U6490 ( .A1(n7700), .A2(n7585), .ZN(n5128) );
  NAND2_X1 U6491 ( .A1(n5947), .A2(n5946), .ZN(n5986) );
  NAND2_X1 U6492 ( .A1(n8425), .A2(n9981), .ZN(n8429) );
  NAND2_X2 U6493 ( .A1(n8991), .A2(n8982), .ZN(n8884) );
  NAND2_X1 U6494 ( .A1(n6746), .A2(n6625), .ZN(n6637) );
  OR2_X1 U6495 ( .A1(n6625), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5873) );
  OR2_X1 U6496 ( .A1(n6625), .A2(n5872), .ZN(n5903) );
  XNOR2_X1 U6497 ( .A(n7634), .B(n7644), .ZN(n7622) );
  OR2_X1 U6498 ( .A1(n6802), .A2(n5915), .ZN(n5898) );
  OR2_X1 U6499 ( .A1(n6083), .A2(n7059), .ZN(n6014) );
  INV_X1 U6500 ( .A(n5945), .ZN(n5947) );
  OR2_X2 U6501 ( .A1(n7063), .A2(n9745), .ZN(n8974) );
  NAND2_X2 U6502 ( .A1(n7612), .A2(n7611), .ZN(n9647) );
  INV_X1 U6503 ( .A(n5358), .ZN(n8042) );
  NAND2_X2 U6504 ( .A1(n5358), .A2(n8041), .ZN(n7807) );
  XNOR2_X1 U6505 ( .A(n8424), .B(n7977), .ZN(n8425) );
  INV_X1 U6506 ( .A(n6047), .ZN(n6336) );
  OR2_X1 U6507 ( .A1(n10064), .A2(n5893), .ZN(n5089) );
  OR2_X1 U6508 ( .A1(n10064), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5090) );
  OR2_X1 U6509 ( .A1(n5943), .A2(n5942), .ZN(n5092) );
  INV_X1 U6510 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5482) );
  AND2_X1 U6511 ( .A1(n5098), .A2(n6585), .ZN(n5093) );
  AND2_X1 U6512 ( .A1(n5977), .A2(n6523), .ZN(n5094) );
  OR2_X1 U6513 ( .A1(n9999), .A2(n5924), .ZN(n5095) );
  INV_X1 U6514 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8722) );
  AOI21_X1 U6515 ( .B1(n6532), .B2(n6531), .A(n9718), .ZN(n8840) );
  INV_X1 U6516 ( .A(n8840), .ZN(n8821) );
  AND2_X1 U6517 ( .A1(n5925), .A2(n5095), .ZN(n5096) );
  AND2_X1 U6518 ( .A1(n8097), .A2(n8446), .ZN(n5097) );
  OR2_X1 U6519 ( .A1(n8035), .A2(n8683), .ZN(n5098) );
  INV_X1 U6520 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6521 ( .A1(n6254), .A2(n6253), .ZN(n5099) );
  AND2_X1 U6522 ( .A1(n5533), .A2(n5527), .ZN(n5100) );
  INV_X1 U6523 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5514) );
  INV_X1 U6524 ( .A(n9983), .ZN(n8565) );
  INV_X1 U6525 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5946) );
  INV_X1 U6526 ( .A(n8280), .ZN(n8426) );
  INV_X1 U6527 ( .A(n9565), .ZN(n7770) );
  INV_X1 U6528 ( .A(n7609), .ZN(n7480) );
  AND2_X1 U6529 ( .A1(n9179), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6530 ( .A1(n8019), .A2(n7465), .ZN(n10044) );
  INV_X1 U6531 ( .A(n10044), .ZN(n6582) );
  AND2_X1 U6532 ( .A1(n5240), .A2(n6670), .ZN(n5102) );
  NAND2_X1 U6533 ( .A1(n6046), .A2(n7233), .ZN(n6035) );
  INV_X1 U6534 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5941) );
  INV_X1 U6535 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5109) );
  NAND2_X1 U6536 ( .A1(n7852), .A2(n6805), .ZN(n6806) );
  INV_X1 U6537 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5924) );
  INV_X1 U6538 ( .A(n5208), .ZN(n5207) );
  OR2_X1 U6539 ( .A1(n9985), .A2(n6810), .ZN(n5383) );
  INV_X1 U6540 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5134) );
  OR2_X1 U6541 ( .A1(n4518), .A2(n7059), .ZN(n6017) );
  AND2_X1 U6542 ( .A1(n6723), .A2(n5981), .ZN(n5980) );
  INV_X1 U6543 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6133) );
  INV_X1 U6544 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5931) );
  INV_X1 U6545 ( .A(n7555), .ZN(n7551) );
  NAND2_X1 U6546 ( .A1(n6803), .A2(n6804), .ZN(n6807) );
  NOR2_X1 U6547 ( .A1(n6697), .A2(n5102), .ZN(n6664) );
  INV_X1 U6548 ( .A(n5332), .ZN(n5269) );
  INV_X1 U6549 ( .A(n5657), .ZN(n5656) );
  NAND2_X1 U6550 ( .A1(n7454), .A2(n5531), .ZN(n7498) );
  XNOR2_X1 U6551 ( .A(n6015), .B(n6081), .ZN(n6038) );
  INV_X1 U6552 ( .A(n9478), .ZN(n9496) );
  INV_X1 U6553 ( .A(SI_26_), .ZN(n10427) );
  INV_X1 U6554 ( .A(SI_23_), .ZN(n10251) );
  INV_X1 U6555 ( .A(n5696), .ZN(n5699) );
  INV_X1 U6556 ( .A(n5646), .ZN(n5648) );
  INV_X1 U6557 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6211) );
  INV_X1 U6558 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6559 ( .A1(n8015), .A2(n8009), .ZN(n8018) );
  NAND2_X1 U6560 ( .A1(n5213), .A2(n5212), .ZN(n5219) );
  AND2_X1 U6561 ( .A1(n8371), .A2(n8617), .ZN(n8372) );
  NOR2_X1 U6562 ( .A1(n8142), .A2(n8565), .ZN(n5854) );
  AND2_X1 U6563 ( .A1(n7852), .A2(n5901), .ZN(n8019) );
  OR2_X1 U6564 ( .A1(n5216), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5157) );
  AND2_X1 U6565 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n6412), .ZN(n6413) );
  INV_X1 U6566 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6260) );
  INV_X1 U6567 ( .A(n8834), .ZN(n8796) );
  NAND2_X1 U6568 ( .A1(n6391), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6411) );
  AND2_X1 U6569 ( .A1(n6542), .A2(n6494), .ZN(n7773) );
  INV_X1 U6570 ( .A(n9608), .ZN(n7738) );
  INV_X1 U6571 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6297) );
  INV_X1 U6572 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6176) );
  AND2_X1 U6573 ( .A1(n9041), .A2(n9043), .ZN(n8895) );
  OR2_X1 U6574 ( .A1(n7783), .A2(n7782), .ZN(n7784) );
  AND2_X1 U6575 ( .A1(n5094), .A2(n5974), .ZN(n5955) );
  NAND2_X1 U6576 ( .A1(n5973), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5975) );
  OR2_X1 U6577 ( .A1(n5469), .A2(n4591), .ZN(n5470) );
  OR2_X1 U6578 ( .A1(n8087), .A2(n6808), .ZN(n6809) );
  INV_X1 U6579 ( .A(n8269), .ZN(n8256) );
  OR2_X1 U6580 ( .A1(n5423), .A2(n10050), .ZN(n5360) );
  INV_X1 U6581 ( .A(n9915), .ZN(n9957) );
  NAND2_X1 U6582 ( .A1(n5920), .A2(n6746), .ZN(n9990) );
  INV_X1 U6583 ( .A(n5914), .ZN(n5913) );
  OR2_X1 U6584 ( .A1(n10048), .A2(n5850), .ZN(n6585) );
  INV_X1 U6585 ( .A(n7842), .ZN(n8503) );
  INV_X1 U6586 ( .A(n7629), .ZN(n8162) );
  INV_X1 U6587 ( .A(n9986), .ZN(n8563) );
  NAND2_X1 U6588 ( .A1(n7856), .A2(n7465), .ZN(n10042) );
  INV_X1 U6589 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5124) );
  INV_X1 U6590 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5150) );
  AND2_X1 U6591 ( .A1(n6413), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6426) );
  OR2_X1 U6592 ( .A1(n8826), .A2(n8827), .ZN(n6471) );
  OR2_X1 U6593 ( .A1(n6261), .A2(n6260), .ZN(n6280) );
  AND2_X1 U6594 ( .A1(n6426), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6443) );
  AND2_X1 U6595 ( .A1(n6378), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6391) );
  AND2_X1 U6596 ( .A1(n6404), .A2(n6403), .ZN(n6405) );
  INV_X1 U6597 ( .A(n8832), .ZN(n8798) );
  OR2_X1 U6598 ( .A1(n6541), .A2(n6540), .ZN(n8834) );
  AND2_X1 U6599 ( .A1(n6365), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6378) );
  OR2_X1 U6600 ( .A1(n6074), .A2(n6024), .ZN(n6029) );
  INV_X1 U6601 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6791) );
  INV_X1 U6602 ( .A(n9412), .ZN(n9427) );
  INV_X1 U6603 ( .A(n9470), .ZN(n8809) );
  NOR2_X1 U6604 ( .A1(n6298), .A2(n6297), .ZN(n6319) );
  NOR2_X1 U6605 ( .A1(n7312), .A2(n7569), .ZN(n7397) );
  NAND2_X1 U6606 ( .A1(n8974), .A2(n8976), .ZN(n7096) );
  AOI21_X1 U6607 ( .B1(n6521), .B2(n10399), .A(n6646), .ZN(n7055) );
  INV_X1 U6608 ( .A(n9828), .ZN(n9758) );
  AND2_X1 U6609 ( .A1(n9046), .A2(n9047), .ZN(n8899) );
  INV_X1 U6610 ( .A(n8893), .ZN(n7396) );
  AND2_X1 U6611 ( .A1(n5826), .A2(n5807), .ZN(n5822) );
  INV_X1 U6612 ( .A(n8271), .ZN(n8258) );
  AND2_X1 U6613 ( .A1(n5799), .A2(n5798), .ZN(n8435) );
  AND4_X1 U6614 ( .A1(n5662), .A2(n5661), .A3(n5660), .A4(n5659), .ZN(n8516)
         );
  AND4_X1 U6615 ( .A1(n5567), .A2(n5566), .A3(n5565), .A4(n5564), .ZN(n7629)
         );
  NOR2_X1 U6616 ( .A1(n7192), .A2(n7460), .ZN(n7191) );
  INV_X1 U6617 ( .A(n7442), .ZN(n9964) );
  NOR2_X1 U6618 ( .A1(n5339), .A2(n7734), .ZN(n9868) );
  INV_X1 U6619 ( .A(n9990), .ZN(n8554) );
  NAND2_X1 U6620 ( .A1(n5845), .A2(n5844), .ZN(n9981) );
  INV_X1 U6621 ( .A(n8609), .ZN(n8629) );
  NAND2_X1 U6622 ( .A1(n7502), .A2(n10044), .ZN(n10035) );
  OR2_X1 U6623 ( .A1(n6758), .A2(n5902), .ZN(n5907) );
  AND2_X1 U6624 ( .A1(n6474), .A2(n6473), .ZN(n6591) );
  INV_X1 U6625 ( .A(n8825), .ZN(n8831) );
  AND4_X1 U6626 ( .A1(n6498), .A2(n6497), .A3(n6496), .A4(n6495), .ZN(n9379)
         );
  INV_X1 U6627 ( .A(n6073), .ZN(n6370) );
  AND4_X1 U6628 ( .A1(n6285), .A2(n6284), .A3(n6283), .A4(n6282), .ZN(n9692)
         );
  NAND2_X1 U6629 ( .A1(n6774), .A2(n9176), .ZN(n9672) );
  NOR2_X1 U6630 ( .A1(n9666), .A2(n9173), .ZN(n9677) );
  INV_X1 U6631 ( .A(n9541), .ZN(n9722) );
  AND2_X1 U6632 ( .A1(n6719), .A2(n6717), .ZN(n9718) );
  INV_X1 U6633 ( .A(n9691), .ZN(n9711) );
  INV_X1 U6634 ( .A(n9484), .ZN(n9726) );
  INV_X1 U6635 ( .A(n9718), .ZN(n9522) );
  AOI21_X1 U6636 ( .B1(n6521), .B2(n10424), .A(n6655), .ZN(n9543) );
  OR2_X1 U6637 ( .A1(n7072), .A2(n4510), .ZN(n9541) );
  AND2_X1 U6638 ( .A1(n7311), .A2(n9736), .ZN(n9762) );
  INV_X1 U6639 ( .A(n9762), .ZN(n9824) );
  INV_X1 U6640 ( .A(n6533), .ZN(n6719) );
  NOR2_X1 U6641 ( .A1(n6220), .A2(n6219), .ZN(n6941) );
  AND2_X1 U6642 ( .A1(n6113), .A2(n6096), .ZN(n9676) );
  OR2_X1 U6643 ( .A1(n6737), .A2(n6816), .ZN(n8271) );
  INV_X1 U6644 ( .A(n8273), .ZN(n8247) );
  INV_X1 U6645 ( .A(n8236), .ZN(n8276) );
  INV_X1 U6646 ( .A(n8435), .ZN(n8411) );
  INV_X1 U6647 ( .A(n8516), .ZN(n8537) );
  INV_X1 U6648 ( .A(n9933), .ZN(n9969) );
  NAND2_X1 U6649 ( .A1(n9868), .A2(n8025), .ZN(n9948) );
  NAND2_X1 U6650 ( .A1(n9999), .A2(n9995), .ZN(n8558) );
  INV_X1 U6651 ( .A(n6808), .ZN(n6846) );
  NAND2_X1 U6652 ( .A1(n10064), .A2(n10040), .ZN(n8609) );
  NAND2_X1 U6653 ( .A1(n10064), .A2(n10035), .ZN(n8626) );
  INV_X1 U6654 ( .A(n10064), .ZN(n10062) );
  INV_X1 U6655 ( .A(n8082), .ZN(n8679) );
  NAND2_X1 U6656 ( .A1(n10048), .A2(n10035), .ZN(n8712) );
  AND3_X1 U6657 ( .A1(n10019), .A2(n10018), .A3(n10017), .ZN(n10055) );
  AND2_X1 U6658 ( .A1(n6930), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6631) );
  INV_X1 U6659 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7732) );
  INV_X1 U6660 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6715) );
  AND2_X1 U6661 ( .A1(n7509), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6598) );
  INV_X1 U6662 ( .A(n9575), .ZN(n9445) );
  INV_X1 U6663 ( .A(n8830), .ZN(n8823) );
  INV_X1 U6664 ( .A(n8835), .ZN(n9420) );
  OAI21_X1 U6665 ( .B1(n8816), .B2(n6370), .A(n6369), .ZN(n9138) );
  INV_X1 U6666 ( .A(n7577), .ZN(n9141) );
  OR2_X1 U6667 ( .A1(n6763), .A2(n6762), .ZN(n9666) );
  INV_X1 U6668 ( .A(n9677), .ZN(n9354) );
  OR2_X1 U6669 ( .A1(n9730), .A2(n9357), .ZN(n9484) );
  OR2_X1 U6670 ( .A1(n9730), .A2(n7077), .ZN(n7317) );
  INV_X1 U6671 ( .A(n9863), .ZN(n9860) );
  INV_X1 U6672 ( .A(n9836), .ZN(n9834) );
  AND2_X2 U6673 ( .A1(n9544), .A2(n7056), .ZN(n9836) );
  AND2_X1 U6674 ( .A1(n6719), .A2(n6644), .ZN(n9735) );
  INV_X1 U6675 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10225) );
  INV_X1 U6676 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10237) );
  INV_X1 U6677 ( .A(n8292), .ZN(P2_U3893) );
  NAND2_X1 U6678 ( .A1(n5896), .A2(n5895), .ZN(P2_U3487) );
  NAND2_X1 U6679 ( .A1(n5912), .A2(n5911), .ZN(P2_U3455) );
  AND2_X2 U6680 ( .A1(n6599), .A2(n6598), .ZN(P1_U3973) );
  INV_X2 U6681 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NAND4_X1 U6682 ( .A1(n5107), .A2(n5156), .A3(n5210), .A4(n5106), .ZN(n5111)
         );
  NAND4_X1 U6683 ( .A1(n5168), .A2(n5109), .A3(n5158), .A4(n5108), .ZN(n5110)
         );
  NOR2_X1 U6684 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5114) );
  NAND2_X1 U6685 ( .A1(n5131), .A2(n5130), .ZN(n5115) );
  INV_X1 U6686 ( .A(n7686), .ZN(n5129) );
  NAND2_X1 U6687 ( .A1(n5122), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5121) );
  MUX2_X1 U6688 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5121), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5123) );
  XNOR2_X1 U6689 ( .A(n5131), .B(n5130), .ZN(n6930) );
  INV_X1 U6690 ( .A(n6930), .ZN(n5141) );
  OR2_X1 U6691 ( .A1(n5899), .A2(n5141), .ZN(n5342) );
  NAND2_X1 U6692 ( .A1(n5133), .A2(n5132), .ZN(n5227) );
  NAND2_X1 U6693 ( .A1(n5228), .A2(n5134), .ZN(n5135) );
  NAND2_X1 U6694 ( .A1(n4551), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5140) );
  OR2_X1 U6695 ( .A1(n8009), .A2(n5141), .ZN(n5142) );
  NAND2_X1 U6696 ( .A1(n5342), .A2(n5142), .ZN(n5339) );
  OR2_X1 U6697 ( .A1(n5339), .A2(n5684), .ZN(n5147) );
  NAND2_X1 U6698 ( .A1(n5147), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U6699 ( .A1(n5152), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5148) );
  XNOR2_X1 U6700 ( .A(n5148), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U6701 ( .A1(n5149), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5151) );
  MUX2_X1 U6702 ( .A(n5151), .B(P2_IR_REG_31__SCAN_IN), .S(n5150), .Z(n5153)
         );
  NAND2_X1 U6703 ( .A1(n5153), .A2(n5152), .ZN(n8354) );
  NAND2_X1 U6704 ( .A1(n5168), .A2(n5210), .ZN(n5155) );
  NAND2_X1 U6705 ( .A1(n5214), .A2(n5156), .ZN(n5216) );
  NAND2_X1 U6706 ( .A1(n5157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5164) );
  NAND2_X1 U6707 ( .A1(n5164), .A2(n5158), .ZN(n5159) );
  NAND2_X1 U6708 ( .A1(n5159), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5163) );
  INV_X1 U6709 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U6710 ( .A1(n5163), .A2(n5160), .ZN(n5161) );
  NAND2_X1 U6711 ( .A1(n5161), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5162) );
  XNOR2_X1 U6712 ( .A(n5162), .B(P2_IR_REG_15__SCAN_IN), .ZN(n5620) );
  XNOR2_X1 U6713 ( .A(n5163), .B(P2_IR_REG_14__SCAN_IN), .ZN(n5603) );
  XNOR2_X1 U6714 ( .A(n5164), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U6715 ( .A1(n5216), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5165) );
  XNOR2_X1 U6716 ( .A(n5165), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7662) );
  INV_X1 U6717 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U6718 ( .A1(n5166), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5169) );
  INV_X1 U6719 ( .A(n5169), .ZN(n5167) );
  NAND2_X1 U6720 ( .A1(n5167), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6721 ( .A1(n5169), .A2(n5168), .ZN(n5209) );
  NAND2_X1 U6722 ( .A1(n5154), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5171) );
  MUX2_X1 U6723 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5171), .S(
        P2_IR_REG_7__SCAN_IN), .Z(n5172) );
  NAND2_X1 U6724 ( .A1(n5186), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5174) );
  INV_X1 U6725 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5173) );
  XNOR2_X1 U6726 ( .A(n5174), .B(n5173), .ZN(n6619) );
  INV_X1 U6727 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5195) );
  NOR2_X1 U6728 ( .A1(n5237), .A2(n5195), .ZN(n5177) );
  NAND2_X1 U6729 ( .A1(n5237), .A2(n5176), .ZN(n5184) );
  INV_X1 U6730 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9865) );
  NAND2_X1 U6731 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5179) );
  INV_X1 U6732 ( .A(n5237), .ZN(n5180) );
  NAND2_X1 U6733 ( .A1(n5237), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5182) );
  INV_X1 U6734 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10050) );
  INV_X1 U6735 ( .A(n5182), .ZN(n5183) );
  XNOR2_X1 U6736 ( .A(n9871), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n9874) );
  NOR2_X1 U6737 ( .A1(n9873), .A2(n9874), .ZN(n9872) );
  NAND2_X1 U6738 ( .A1(n5184), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5185) );
  MUX2_X1 U6739 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5185), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5187) );
  NAND2_X1 U6740 ( .A1(n5187), .A2(n5186), .ZN(n6616) );
  AOI21_X1 U6741 ( .B1(n5188), .B2(n6670), .A(n6703), .ZN(n6661) );
  NAND2_X1 U6742 ( .A1(n6661), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6662) );
  INV_X1 U6743 ( .A(n6703), .ZN(n5189) );
  XNOR2_X1 U6744 ( .A(n6619), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n6701) );
  OR2_X1 U6745 ( .A1(n4576), .A2(n5195), .ZN(n5190) );
  NOR2_X1 U6746 ( .A1(n5191), .A2(n9896), .ZN(n5193) );
  INV_X1 U6747 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9888) );
  NOR2_X1 U6748 ( .A1(n5194), .A2(n5195), .ZN(n5196) );
  MUX2_X1 U6749 ( .A(n5195), .B(n5196), .S(P2_IR_REG_6__SCAN_IN), .Z(n5197) );
  NAND2_X1 U6750 ( .A1(n9912), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5200) );
  OAI21_X1 U6751 ( .B1(n9912), .B2(P2_REG1_REG_6__SCAN_IN), .A(n5200), .ZN(
        n9904) );
  INV_X1 U6752 ( .A(n9904), .ZN(n5198) );
  NOR2_X1 U6753 ( .A1(n5249), .A2(n5201), .ZN(n5202) );
  INV_X1 U6754 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10057) );
  NOR2_X1 U6755 ( .A1(n5202), .A2(n9939), .ZN(n9952) );
  NAND2_X1 U6756 ( .A1(n5203), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5204) );
  XNOR2_X1 U6757 ( .A(n5204), .B(P2_IR_REG_8__SCAN_IN), .ZN(n5510) );
  INV_X1 U6758 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5497) );
  OR2_X1 U6759 ( .A1(n5510), .A2(n5497), .ZN(n5206) );
  NAND2_X1 U6760 ( .A1(n5510), .A2(n5497), .ZN(n5205) );
  NAND2_X1 U6761 ( .A1(n5206), .A2(n5205), .ZN(n9951) );
  INV_X1 U6762 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U6763 ( .A1(n5209), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6764 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7343), .ZN(n5212) );
  OAI21_X1 U6765 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7343), .A(n5212), .ZN(
        n7340) );
  NOR2_X1 U6766 ( .A1(n5214), .A2(n5195), .ZN(n5215) );
  MUX2_X1 U6767 ( .A(n5195), .B(n5215), .S(P2_IR_REG_11__SCAN_IN), .Z(n5218)
         );
  INV_X1 U6768 ( .A(n5216), .ZN(n5217) );
  NOR2_X1 U6769 ( .A1(n5218), .A2(n5217), .ZN(n7446) );
  AND2_X1 U6770 ( .A1(n5219), .A2(n6657), .ZN(n5220) );
  INV_X1 U6771 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7680) );
  XNOR2_X1 U6772 ( .A(n7662), .B(n7680), .ZN(n7659) );
  NOR2_X1 U6773 ( .A1(n8305), .A2(n5221), .ZN(n5222) );
  INV_X1 U6774 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8302) );
  NOR2_X1 U6775 ( .A1(n8302), .A2(n8303), .ZN(n8301) );
  INV_X1 U6776 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8628) );
  XNOR2_X1 U6777 ( .A(n5603), .B(n8628), .ZN(n8313) );
  NOR2_X1 U6778 ( .A1(n8314), .A2(n8313), .ZN(n8312) );
  NOR2_X1 U6779 ( .A1(n5620), .A2(n5223), .ZN(n5224) );
  INV_X1 U6780 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8623) );
  XNOR2_X1 U6781 ( .A(n8354), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8348) );
  NOR2_X1 U6782 ( .A1(n8349), .A2(n8348), .ZN(n8347) );
  NOR2_X1 U6783 ( .A1(n8375), .A2(n5225), .ZN(n5226) );
  INV_X1 U6784 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8617) );
  XNOR2_X1 U6785 ( .A(n8375), .B(n5225), .ZN(n8371) );
  NAND2_X1 U6786 ( .A1(n5227), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5229) );
  OR2_X1 U6787 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  AND2_X1 U6788 ( .A1(n5233), .A2(n5230), .ZN(n5666) );
  INV_X1 U6789 ( .A(n5666), .ZN(n8391) );
  NAND2_X1 U6790 ( .A1(n8391), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5231) );
  OAI21_X1 U6791 ( .B1(n8391), .B2(P2_REG1_REG_18__SCAN_IN), .A(n5231), .ZN(
        n8383) );
  INV_X1 U6792 ( .A(n5231), .ZN(n5232) );
  XNOR2_X1 U6793 ( .A(n5901), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n5333) );
  XNOR2_X1 U6794 ( .A(n5234), .B(n5333), .ZN(n5351) );
  OR2_X1 U6795 ( .A1(n5235), .A2(P2_U3151), .ZN(n7734) );
  INV_X1 U6796 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9929) );
  INV_X1 U6797 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9890) );
  INV_X1 U6798 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U6799 ( .A1(n5237), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5238) );
  INV_X1 U6800 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6683) );
  INV_X1 U6801 ( .A(n5238), .ZN(n5239) );
  NAND2_X1 U6802 ( .A1(n6664), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6665) );
  INV_X1 U6803 ( .A(n6697), .ZN(n5241) );
  XNOR2_X1 U6804 ( .A(n6619), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6695) );
  AOI21_X1 U6805 ( .B1(n6665), .B2(n5241), .A(n6695), .ZN(n6700) );
  NAND2_X1 U6806 ( .A1(n5242), .A2(n9896), .ZN(n5243) );
  INV_X1 U6807 ( .A(n9907), .ZN(n5245) );
  NAND2_X1 U6808 ( .A1(n9912), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5246) );
  OAI21_X1 U6809 ( .B1(n9912), .B2(P2_REG2_REG_6__SCAN_IN), .A(n5246), .ZN(
        n9908) );
  INV_X1 U6810 ( .A(n9908), .ZN(n5244) );
  NAND2_X1 U6811 ( .A1(n5245), .A2(n5244), .ZN(n9910) );
  NAND2_X1 U6812 ( .A1(n9910), .A2(n5246), .ZN(n5247) );
  NOR2_X1 U6813 ( .A1(n5249), .A2(n5248), .ZN(n5250) );
  INV_X1 U6814 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5282) );
  OR2_X1 U6815 ( .A1(n5510), .A2(n5282), .ZN(n5252) );
  NAND2_X1 U6816 ( .A1(n5510), .A2(n5282), .ZN(n5251) );
  NAND2_X1 U6817 ( .A1(n5252), .A2(n5251), .ZN(n9946) );
  XNOR2_X1 U6818 ( .A(n5253), .B(n5528), .ZN(n7192) );
  INV_X1 U6819 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7460) );
  NOR2_X1 U6820 ( .A1(n5528), .A2(n5253), .ZN(n5254) );
  NAND2_X1 U6821 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7343), .ZN(n5255) );
  OAI21_X1 U6822 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7343), .A(n5255), .ZN(
        n7337) );
  NAND2_X1 U6823 ( .A1(n5257), .A2(n6657), .ZN(n5256) );
  INV_X1 U6824 ( .A(n5256), .ZN(n5258) );
  INV_X1 U6825 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7536) );
  OAI21_X1 U6826 ( .B1(n5257), .B2(n6657), .A(n5256), .ZN(n7432) );
  INV_X1 U6827 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7675) );
  AOI22_X1 U6828 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n7662), .B1(n6716), .B2(
        n7675), .ZN(n7656) );
  NOR2_X1 U6829 ( .A1(n8305), .A2(n5259), .ZN(n5260) );
  INV_X1 U6830 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8296) );
  XNOR2_X1 U6831 ( .A(n8305), .B(n5259), .ZN(n8295) );
  NOR2_X1 U6832 ( .A1(n8296), .A2(n8295), .ZN(n8294) );
  INV_X1 U6833 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8571) );
  AOI22_X1 U6834 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n5603), .B1(n8320), .B2(
        n8571), .ZN(n8322) );
  NOR2_X1 U6835 ( .A1(n5620), .A2(n5261), .ZN(n5262) );
  INV_X1 U6836 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8332) );
  INV_X1 U6837 ( .A(n5620), .ZN(n8341) );
  NAND2_X1 U6838 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8354), .ZN(n5263) );
  OAI21_X1 U6839 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8354), .A(n5263), .ZN(
        n8359) );
  NOR2_X1 U6840 ( .A1(n8375), .A2(n5264), .ZN(n5265) );
  INV_X1 U6841 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8367) );
  INV_X1 U6842 ( .A(n8375), .ZN(n6967) );
  NOR2_X1 U6843 ( .A1(n8367), .A2(n8366), .ZN(n8365) );
  NAND2_X1 U6844 ( .A1(n8391), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5266) );
  OAI21_X1 U6845 ( .B1(n8391), .B2(P2_REG2_REG_18__SCAN_IN), .A(n5266), .ZN(
        n8394) );
  INV_X1 U6846 ( .A(n5266), .ZN(n5267) );
  NOR2_X1 U6847 ( .A1(n8393), .A2(n5267), .ZN(n5270) );
  INV_X1 U6848 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5268) );
  MUX2_X1 U6849 ( .A(n5268), .B(P2_REG2_REG_19__SCAN_IN), .S(n5901), .Z(n5332)
         );
  XNOR2_X1 U6850 ( .A(n5270), .B(n5269), .ZN(n5349) );
  INV_X2 U6851 ( .A(n8025), .ZN(n5315) );
  NAND2_X1 U6852 ( .A1(n5324), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5271) );
  OAI21_X1 U6853 ( .B1(n5315), .B2(n8367), .A(n5271), .ZN(n5272) );
  OR2_X1 U6854 ( .A1(n5272), .A2(n6967), .ZN(n5323) );
  XNOR2_X1 U6855 ( .A(n5272), .B(n8375), .ZN(n8370) );
  INV_X1 U6856 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U6857 ( .A1(n5324), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5273) );
  OAI21_X1 U6858 ( .B1(n5315), .B2(n8539), .A(n5273), .ZN(n5274) );
  OR2_X1 U6859 ( .A1(n8354), .A2(n5274), .ZN(n5322) );
  INV_X1 U6860 ( .A(n8354), .ZN(n5637) );
  XNOR2_X1 U6861 ( .A(n5274), .B(n5637), .ZN(n8352) );
  NAND2_X1 U6862 ( .A1(n5315), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5275) );
  OAI21_X1 U6863 ( .B1(n5315), .B2(n8332), .A(n5275), .ZN(n5276) );
  OR2_X1 U6864 ( .A1(n8341), .A2(n5276), .ZN(n5321) );
  XNOR2_X1 U6865 ( .A(n5620), .B(n5276), .ZN(n8335) );
  OR2_X1 U6866 ( .A1(n5324), .A2(n8571), .ZN(n5278) );
  NAND2_X1 U6867 ( .A1(n5324), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5277) );
  NAND2_X1 U6868 ( .A1(n5278), .A2(n5277), .ZN(n5279) );
  OR2_X1 U6869 ( .A1(n8320), .A2(n5279), .ZN(n5320) );
  XNOR2_X1 U6870 ( .A(n5603), .B(n5279), .ZN(n8317) );
  NAND2_X1 U6871 ( .A1(n5315), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5280) );
  OAI21_X1 U6872 ( .B1(n5315), .B2(n8296), .A(n5280), .ZN(n5318) );
  INV_X1 U6873 ( .A(n5318), .ZN(n5281) );
  NAND2_X1 U6874 ( .A1(n8305), .A2(n5281), .ZN(n5319) );
  MUX2_X1 U6875 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n5315), .Z(n5311) );
  NOR2_X1 U6876 ( .A1(n5311), .A2(n6657), .ZN(n5313) );
  MUX2_X1 U6877 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n5315), .Z(n5308) );
  NOR2_X1 U6878 ( .A1(n5308), .A2(n7343), .ZN(n5310) );
  MUX2_X1 U6879 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n5315), .Z(n5305) );
  NOR2_X1 U6880 ( .A1(n5305), .A2(n7196), .ZN(n5307) );
  OR2_X1 U6881 ( .A1(n5324), .A2(n5282), .ZN(n5284) );
  NAND2_X1 U6882 ( .A1(n5315), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6883 ( .A1(n5284), .A2(n5283), .ZN(n5303) );
  INV_X1 U6884 ( .A(n5510), .ZN(n9956) );
  NOR2_X1 U6885 ( .A1(n5303), .A2(n9956), .ZN(n5304) );
  MUX2_X1 U6886 ( .A(n9929), .B(n10057), .S(n5315), .Z(n5301) );
  INV_X1 U6887 ( .A(n5301), .ZN(n5302) );
  MUX2_X1 U6888 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n5324), .Z(n5300) );
  INV_X1 U6889 ( .A(n6619), .ZN(n6710) );
  MUX2_X1 U6890 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n5315), .Z(n5295) );
  INV_X1 U6891 ( .A(n5295), .ZN(n5296) );
  OR2_X1 U6892 ( .A1(n5324), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6893 ( .A1(n5324), .A2(n10050), .ZN(n5285) );
  NAND2_X1 U6894 ( .A1(n5286), .A2(n5285), .ZN(n5289) );
  XOR2_X1 U6895 ( .A(n6678), .B(n5289), .Z(n6677) );
  MUX2_X1 U6896 ( .A(n6844), .B(n9865), .S(n5315), .Z(n5287) );
  AND2_X1 U6897 ( .A1(n5287), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9866) );
  OAI22_X1 U6898 ( .A1(n6677), .A2(n9866), .B1(n5288), .B2(n5289), .ZN(n9882)
         );
  INV_X1 U6899 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10001) );
  OR2_X1 U6900 ( .A1(n5324), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5291) );
  INV_X1 U6901 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10052) );
  NAND2_X1 U6902 ( .A1(n5315), .A2(n10052), .ZN(n5290) );
  NAND2_X1 U6903 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  XNOR2_X1 U6904 ( .A(n5292), .B(n4513), .ZN(n9883) );
  INV_X1 U6905 ( .A(n5292), .ZN(n5293) );
  AOI22_X1 U6906 ( .A1(n9882), .A2(n9883), .B1(n5293), .B2(n4513), .ZN(n6671)
         );
  INV_X1 U6907 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5403) );
  INV_X1 U6908 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5404) );
  MUX2_X1 U6909 ( .A(n5403), .B(n5404), .S(n5315), .Z(n5294) );
  XNOR2_X1 U6910 ( .A(n5294), .B(n6616), .ZN(n6672) );
  NAND2_X1 U6911 ( .A1(n6671), .A2(n6672), .ZN(n6691) );
  NAND2_X1 U6912 ( .A1(n5294), .A2(n6670), .ZN(n6690) );
  XNOR2_X1 U6913 ( .A(n5295), .B(n6710), .ZN(n6693) );
  NAND3_X1 U6914 ( .A1(n6691), .A2(n6690), .A3(n6693), .ZN(n6692) );
  OAI21_X1 U6915 ( .B1(n6710), .B2(n5296), .A(n6692), .ZN(n9897) );
  OR2_X1 U6916 ( .A1(n5324), .A2(n9890), .ZN(n5298) );
  NAND2_X1 U6917 ( .A1(n5315), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6918 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  XNOR2_X1 U6919 ( .A(n5299), .B(n9896), .ZN(n9898) );
  INV_X1 U6920 ( .A(n9896), .ZN(n6609) );
  AOI22_X1 U6921 ( .A1(n9897), .A2(n9898), .B1(n6609), .B2(n5299), .ZN(n9922)
         );
  XOR2_X1 U6922 ( .A(n9912), .B(n5300), .Z(n9921) );
  NAND2_X1 U6923 ( .A1(n9922), .A2(n9921), .ZN(n9920) );
  OAI21_X1 U6924 ( .B1(n5300), .B2(n9912), .A(n9920), .ZN(n9936) );
  XNOR2_X1 U6925 ( .A(n5301), .B(n9930), .ZN(n9937) );
  NAND2_X1 U6926 ( .A1(n9936), .A2(n9937), .ZN(n9935) );
  OAI21_X1 U6927 ( .B1(n5302), .B2(n9930), .A(n9935), .ZN(n9963) );
  AOI21_X1 U6928 ( .B1(n9956), .B2(n5303), .A(n5304), .ZN(n9962) );
  AND2_X1 U6929 ( .A1(n9963), .A2(n9962), .ZN(n9966) );
  NOR2_X1 U6930 ( .A1(n5304), .A2(n9966), .ZN(n7198) );
  AOI21_X1 U6931 ( .B1(n7196), .B2(n5305), .A(n5307), .ZN(n5306) );
  INV_X1 U6932 ( .A(n5306), .ZN(n7199) );
  NOR2_X1 U6933 ( .A1(n7198), .A2(n7199), .ZN(n7197) );
  NOR2_X1 U6934 ( .A1(n5307), .A2(n7197), .ZN(n7345) );
  AOI21_X1 U6935 ( .B1(n7343), .B2(n5308), .A(n5310), .ZN(n5309) );
  INV_X1 U6936 ( .A(n5309), .ZN(n7346) );
  NOR2_X1 U6937 ( .A1(n7345), .A2(n7346), .ZN(n7344) );
  NOR2_X1 U6938 ( .A1(n5310), .A2(n7344), .ZN(n7439) );
  AOI21_X1 U6939 ( .B1(n6657), .B2(n5311), .A(n5313), .ZN(n5312) );
  INV_X1 U6940 ( .A(n5312), .ZN(n7440) );
  NOR2_X1 U6941 ( .A1(n7439), .A2(n7440), .ZN(n7438) );
  NOR2_X1 U6942 ( .A1(n5313), .A2(n7438), .ZN(n7654) );
  AOI21_X1 U6943 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n5315), .A(n6716), .ZN(
        n5314) );
  OAI21_X1 U6944 ( .B1(n5315), .B2(n7675), .A(n5314), .ZN(n7651) );
  OR2_X1 U6945 ( .A1(n5324), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5317) );
  AOI21_X1 U6946 ( .B1(n5315), .B2(n7680), .A(n7662), .ZN(n5316) );
  AND2_X1 U6947 ( .A1(n5317), .A2(n5316), .ZN(n7650) );
  AOI21_X1 U6948 ( .B1(n7654), .B2(n7651), .A(n7650), .ZN(n8299) );
  XNOR2_X1 U6949 ( .A(n5318), .B(n8305), .ZN(n8298) );
  NAND2_X1 U6950 ( .A1(n8299), .A2(n8298), .ZN(n8297) );
  NAND2_X1 U6951 ( .A1(n5319), .A2(n8297), .ZN(n8316) );
  NAND2_X1 U6952 ( .A1(n8317), .A2(n8316), .ZN(n8315) );
  NAND2_X1 U6953 ( .A1(n5320), .A2(n8315), .ZN(n8334) );
  NAND2_X1 U6954 ( .A1(n8335), .A2(n8334), .ZN(n8333) );
  NAND2_X1 U6955 ( .A1(n5321), .A2(n8333), .ZN(n8351) );
  NAND2_X1 U6956 ( .A1(n8352), .A2(n8351), .ZN(n8350) );
  NAND2_X1 U6957 ( .A1(n5322), .A2(n8350), .ZN(n8369) );
  NAND2_X1 U6958 ( .A1(n8370), .A2(n8369), .ZN(n8368) );
  AND2_X1 U6959 ( .A1(n5323), .A2(n8368), .ZN(n5327) );
  INV_X1 U6960 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8519) );
  OR2_X1 U6961 ( .A1(n5324), .A2(n8519), .ZN(n5326) );
  NAND2_X1 U6962 ( .A1(n5324), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6963 ( .A1(n5326), .A2(n5325), .ZN(n5328) );
  NAND2_X1 U6964 ( .A1(n5327), .A2(n5328), .ZN(n8386) );
  NAND2_X1 U6965 ( .A1(n8386), .A2(n5666), .ZN(n5331) );
  INV_X1 U6966 ( .A(n5327), .ZN(n5330) );
  INV_X1 U6967 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U6968 ( .A1(n5330), .A2(n5329), .ZN(n8385) );
  NAND2_X1 U6969 ( .A1(n5331), .A2(n8385), .ZN(n5335) );
  MUX2_X1 U6970 ( .A(n5333), .B(n5332), .S(n8025), .Z(n5334) );
  XNOR2_X1 U6971 ( .A(n5335), .B(n5334), .ZN(n5336) );
  INV_X1 U6972 ( .A(n6631), .ZN(n6751) );
  INV_X1 U6973 ( .A(n5235), .ZN(n5847) );
  OR2_X1 U6974 ( .A1(n8292), .A2(n5847), .ZN(n7442) );
  NOR2_X1 U6975 ( .A1(n5315), .A2(P2_U3151), .ZN(n5337) );
  NAND2_X1 U6976 ( .A1(n5337), .A2(n5235), .ZN(n5338) );
  OR2_X1 U6977 ( .A1(n5339), .A2(n5338), .ZN(n5341) );
  OR2_X1 U6978 ( .A1(n5342), .A2(n7734), .ZN(n5340) );
  NAND2_X1 U6979 ( .A1(n5341), .A2(n5340), .ZN(n9915) );
  INV_X1 U6980 ( .A(n5342), .ZN(n5343) );
  NAND2_X1 U6981 ( .A1(n9933), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6982 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8127) );
  OAI211_X1 U6983 ( .C1(n9957), .C2(n7850), .A(n5344), .B(n8127), .ZN(n5345)
         );
  INV_X1 U6984 ( .A(n5345), .ZN(n5346) );
  NAND2_X1 U6985 ( .A1(n5354), .A2(n5355), .ZN(n8726) );
  NAND2_X1 U6987 ( .A1(n5401), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6988 ( .A1(n5420), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5361) );
  INV_X1 U6989 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6879) );
  NAND4_X1 U6990 ( .A1(n5362), .A2(n5361), .A3(n5360), .A4(n5359), .ZN(n5382)
         );
  NAND2_X1 U6991 ( .A1(n5364), .A2(n5363), .ZN(n5366) );
  NAND2_X1 U6992 ( .A1(n5367), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5368) );
  INV_X1 U6993 ( .A(SI_1_), .ZN(n5371) );
  NAND2_X1 U6994 ( .A1(n7798), .A2(SI_0_), .ZN(n5381) );
  INV_X1 U6995 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5373) );
  AND2_X1 U6996 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5372) );
  NAND2_X1 U6997 ( .A1(n6605), .A2(n5372), .ZN(n6022) );
  XNOR2_X1 U6998 ( .A(n5391), .B(n5390), .ZN(n6606) );
  INV_X1 U6999 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6607) );
  OR2_X1 U7000 ( .A1(n5374), .A2(n6678), .ZN(n5375) );
  NAND2_X1 U7001 ( .A1(n5382), .A2(n10002), .ZN(n7854) );
  NAND2_X1 U7002 ( .A1(n5832), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5380) );
  OR2_X1 U7003 ( .A1(n7807), .A2(n6844), .ZN(n5379) );
  INV_X1 U7004 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5376) );
  OR2_X1 U7005 ( .A1(n5452), .A2(n5376), .ZN(n5378) );
  OR2_X1 U7006 ( .A1(n5423), .A2(n9865), .ZN(n5377) );
  XNOR2_X1 U7007 ( .A(n5381), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8730) );
  MUX2_X1 U7008 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8730), .S(n6576), .Z(n6808) );
  NAND2_X1 U7009 ( .A1(n8293), .A2(n6808), .ZN(n6873) );
  NAND2_X1 U7010 ( .A1(n7825), .A2(n6873), .ZN(n5384) );
  INV_X1 U7011 ( .A(n10002), .ZN(n6810) );
  NAND2_X1 U7012 ( .A1(n5384), .A2(n5383), .ZN(n9979) );
  NAND2_X1 U7013 ( .A1(n5420), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5389) );
  INV_X1 U7014 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10468) );
  OR2_X1 U7015 ( .A1(n5402), .A2(n10468), .ZN(n5388) );
  INV_X1 U7016 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5385) );
  OR2_X1 U7017 ( .A1(n5423), .A2(n10052), .ZN(n5386) );
  NAND4_X1 U7018 ( .A1(n5389), .A2(n5388), .A3(n5387), .A4(n5386), .ZN(n5398)
         );
  NAND2_X1 U7019 ( .A1(n5392), .A2(SI_1_), .ZN(n5393) );
  INV_X1 U7020 ( .A(SI_2_), .ZN(n5394) );
  XNOR2_X1 U7021 ( .A(n5411), .B(n5410), .ZN(n6612) );
  OR2_X1 U7022 ( .A1(n5409), .A2(n6612), .ZN(n5397) );
  INV_X1 U7023 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6613) );
  OR2_X1 U7024 ( .A1(n7803), .A2(n6613), .ZN(n5396) );
  OR2_X1 U7025 ( .A1(n5398), .A2(n9989), .ZN(n7863) );
  NAND2_X1 U7026 ( .A1(n5398), .A2(n9989), .ZN(n7864) );
  NAND2_X1 U7027 ( .A1(n9979), .A2(n9980), .ZN(n5400) );
  INV_X1 U7028 ( .A(n9989), .ZN(n6860) );
  OR2_X1 U7029 ( .A1(n5398), .A2(n6860), .ZN(n5399) );
  NAND2_X1 U7030 ( .A1(n5400), .A2(n5399), .ZN(n9970) );
  NAND2_X1 U7031 ( .A1(n5401), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5408) );
  OR2_X1 U7032 ( .A1(n5402), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5407) );
  OR2_X1 U7033 ( .A1(n7807), .A2(n5403), .ZN(n5406) );
  OR2_X1 U7034 ( .A1(n5423), .A2(n5404), .ZN(n5405) );
  NAND2_X1 U7035 ( .A1(n5412), .A2(SI_2_), .ZN(n5413) );
  INV_X1 U7036 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6618) );
  INV_X1 U7037 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6603) );
  MUX2_X1 U7038 ( .A(n6618), .B(n6603), .S(n6600), .Z(n5431) );
  XNOR2_X1 U7039 ( .A(n5431), .B(SI_3_), .ZN(n5429) );
  XNOR2_X1 U7040 ( .A(n5429), .B(n5430), .ZN(n6617) );
  OR2_X1 U7041 ( .A1(n5409), .A2(n6617), .ZN(n5416) );
  OR2_X1 U7042 ( .A1(n7803), .A2(n6618), .ZN(n5415) );
  OAI211_X1 U7043 ( .C1(n6576), .C2(n6616), .A(n5416), .B(n5415), .ZN(n6934)
         );
  NOR2_X1 U7044 ( .A1(n9984), .A2(n6934), .ZN(n5417) );
  NAND2_X1 U7045 ( .A1(n9984), .A2(n6934), .ZN(n5418) );
  OAI21_X1 U7046 ( .B1(n9970), .B2(n5417), .A(n5418), .ZN(n5419) );
  INV_X1 U7047 ( .A(n5419), .ZN(n6913) );
  NAND2_X1 U7048 ( .A1(n5420), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5428) );
  INV_X1 U7049 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5421) );
  OR2_X1 U7050 ( .A1(n6572), .A2(n5421), .ZN(n5427) );
  NAND2_X1 U7051 ( .A1(n10269), .A2(n10223), .ZN(n5439) );
  NAND2_X1 U7052 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5422) );
  AND2_X1 U7053 ( .A1(n5439), .A2(n5422), .ZN(n6962) );
  OR2_X1 U7054 ( .A1(n5402), .A2(n6962), .ZN(n5426) );
  INV_X1 U7055 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U7056 ( .A1(n5430), .A2(n5429), .ZN(n5465) );
  INV_X1 U7057 ( .A(n5431), .ZN(n5432) );
  NAND2_X1 U7058 ( .A1(n5432), .A2(SI_3_), .ZN(n5463) );
  NAND2_X1 U7059 ( .A1(n5465), .A2(n5463), .ZN(n5445) );
  INV_X1 U7060 ( .A(SI_4_), .ZN(n10266) );
  XNOR2_X1 U7061 ( .A(n5445), .B(n5468), .ZN(n6620) );
  OR2_X1 U7062 ( .A1(n5409), .A2(n6620), .ZN(n5435) );
  INV_X1 U7063 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6621) );
  OR2_X1 U7064 ( .A1(n7803), .A2(n6621), .ZN(n5434) );
  OR2_X1 U7065 ( .A1(n6576), .A2(n6619), .ZN(n5433) );
  NAND2_X1 U7066 ( .A1(n9971), .A2(n10016), .ZN(n7877) );
  INV_X1 U7067 ( .A(n10016), .ZN(n6959) );
  OR2_X1 U7068 ( .A1(n9971), .A2(n6959), .ZN(n5436) );
  NAND2_X1 U7069 ( .A1(n5401), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5444) );
  OR2_X1 U7070 ( .A1(n7807), .A2(n9890), .ZN(n5443) );
  OR2_X1 U7071 ( .A1(n7811), .A2(n9888), .ZN(n5442) );
  INV_X1 U7072 ( .A(n5439), .ZN(n5438) );
  NAND2_X1 U7073 ( .A1(n5438), .A2(n5437), .ZN(n5454) );
  NAND2_X1 U7074 ( .A1(n5439), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5440) );
  AND2_X1 U7075 ( .A1(n5454), .A2(n5440), .ZN(n7003) );
  OR2_X1 U7076 ( .A1(n5402), .A2(n7003), .ZN(n5441) );
  NAND2_X1 U7077 ( .A1(n5445), .A2(n5468), .ZN(n5447) );
  NAND2_X1 U7078 ( .A1(n5446), .A2(SI_4_), .ZN(n5461) );
  NAND2_X1 U7079 ( .A1(n5447), .A2(n5461), .ZN(n5448) );
  INV_X1 U7080 ( .A(SI_5_), .ZN(n10474) );
  XNOR2_X1 U7081 ( .A(n5448), .B(n5467), .ZN(n6610) );
  OR2_X1 U7082 ( .A1(n5409), .A2(n6610), .ZN(n5451) );
  INV_X1 U7083 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6611) );
  OR2_X1 U7084 ( .A1(n7803), .A2(n6611), .ZN(n5450) );
  OR2_X1 U7085 ( .A1(n6576), .A2(n6609), .ZN(n5449) );
  NAND2_X1 U7086 ( .A1(n6569), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5460) );
  INV_X1 U7087 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5453) );
  OR2_X1 U7088 ( .A1(n6572), .A2(n5453), .ZN(n5459) );
  NAND2_X1 U7089 ( .A1(n5454), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5455) );
  AND2_X1 U7090 ( .A1(n5484), .A2(n5455), .ZN(n7213) );
  OR2_X1 U7091 ( .A1(n5402), .A2(n7213), .ZN(n5458) );
  INV_X1 U7092 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5456) );
  OR2_X1 U7093 ( .A1(n7811), .A2(n5456), .ZN(n5457) );
  OR2_X1 U7094 ( .A1(n5462), .A2(n5461), .ZN(n5466) );
  AND2_X1 U7095 ( .A1(n5463), .A2(n5466), .ZN(n5464) );
  NAND2_X1 U7096 ( .A1(n5465), .A2(n5464), .ZN(n5471) );
  INV_X1 U7097 ( .A(n5466), .ZN(n5469) );
  NAND2_X1 U7098 ( .A1(n5471), .A2(n5470), .ZN(n5474) );
  NAND2_X1 U7099 ( .A1(n5472), .A2(SI_5_), .ZN(n5473) );
  MUX2_X1 U7100 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6605), .Z(n5492) );
  INV_X1 U7101 ( .A(SI_6_), .ZN(n5475) );
  XNOR2_X1 U7102 ( .A(n5492), .B(n5475), .ZN(n5490) );
  XNOR2_X1 U7103 ( .A(n5491), .B(n5490), .ZN(n6614) );
  OR2_X1 U7104 ( .A1(n5409), .A2(n6614), .ZN(n5477) );
  INV_X1 U7105 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6615) );
  OR2_X1 U7106 ( .A1(n7803), .A2(n6615), .ZN(n5476) );
  OAI211_X1 U7107 ( .C1(n6576), .C2(n9912), .A(n5477), .B(n5476), .ZN(n7215)
         );
  NAND2_X1 U7108 ( .A1(n5478), .A2(n7215), .ZN(n5481) );
  NAND2_X1 U7109 ( .A1(n5479), .A2(n8290), .ZN(n5480) );
  NAND2_X1 U7110 ( .A1(n5401), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5489) );
  OR2_X1 U7111 ( .A1(n7811), .A2(n10057), .ZN(n5488) );
  OR2_X1 U7112 ( .A1(n7807), .A2(n9929), .ZN(n5487) );
  NAND2_X1 U7113 ( .A1(n5484), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5485) );
  AND2_X1 U7114 ( .A1(n5498), .A2(n5485), .ZN(n7327) );
  OR2_X1 U7115 ( .A1(n5402), .A2(n7327), .ZN(n5486) );
  NAND4_X1 U7116 ( .A1(n5489), .A2(n5488), .A3(n5487), .A4(n5486), .ZN(n8289)
         );
  NAND2_X1 U7117 ( .A1(n5492), .A2(SI_6_), .ZN(n5493) );
  MUX2_X1 U7118 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6605), .Z(n5506) );
  INV_X1 U7119 ( .A(SI_7_), .ZN(n5494) );
  XNOR2_X1 U7120 ( .A(n5506), .B(n5494), .ZN(n5505) );
  INV_X1 U7121 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6624) );
  OR2_X1 U7122 ( .A1(n7803), .A2(n6624), .ZN(n5495) );
  OR2_X1 U7123 ( .A1(n8289), .A2(n7321), .ZN(n5496) );
  NAND2_X1 U7124 ( .A1(n6569), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5504) );
  OR2_X1 U7125 ( .A1(n7811), .A2(n5497), .ZN(n5503) );
  NAND2_X1 U7126 ( .A1(n5498), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5499) );
  AND2_X1 U7127 ( .A1(n5516), .A2(n5499), .ZN(n7417) );
  OR2_X1 U7128 ( .A1(n5402), .A2(n7417), .ZN(n5502) );
  INV_X1 U7129 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5500) );
  OR2_X1 U7130 ( .A1(n6572), .A2(n5500), .ZN(n5501) );
  INV_X1 U7131 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6636) );
  INV_X1 U7132 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6634) );
  MUX2_X1 U7133 ( .A(n6636), .B(n6634), .S(n6605), .Z(n5507) );
  NAND2_X1 U7134 ( .A1(n5507), .A2(n10416), .ZN(n5522) );
  INV_X1 U7135 ( .A(n5507), .ZN(n5508) );
  NAND2_X1 U7136 ( .A1(n5508), .A2(SI_8_), .ZN(n5509) );
  NAND2_X1 U7137 ( .A1(n5522), .A2(n5509), .ZN(n5523) );
  XNOR2_X1 U7138 ( .A(n5524), .B(n5523), .ZN(n6633) );
  NAND2_X1 U7139 ( .A1(n6633), .A2(n5535), .ZN(n5512) );
  AOI22_X1 U7140 ( .A1(n5685), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5684), .B2(
        n5510), .ZN(n5511) );
  NAND2_X1 U7141 ( .A1(n5512), .A2(n5511), .ZN(n7429) );
  NOR2_X1 U7142 ( .A1(n8288), .A2(n7429), .ZN(n5513) );
  INV_X1 U7143 ( .A(n8288), .ZN(n7547) );
  OAI22_X1 U7144 ( .A1(n7408), .A2(n5513), .B1(n10031), .B2(n7547), .ZN(n7453)
         );
  NAND2_X1 U7145 ( .A1(n5401), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5521) );
  OR2_X1 U7146 ( .A1(n7807), .A2(n7460), .ZN(n5520) );
  NAND2_X1 U7147 ( .A1(n5516), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5517) );
  AND2_X1 U7148 ( .A1(n5540), .A2(n5517), .ZN(n7541) );
  OR2_X1 U7149 ( .A1(n5402), .A2(n7541), .ZN(n5519) );
  OR2_X1 U7150 ( .A1(n7811), .A2(n10060), .ZN(n5518) );
  MUX2_X1 U7151 ( .A(n6639), .B(n10237), .S(n6600), .Z(n5525) );
  NAND2_X1 U7152 ( .A1(n5525), .A2(n10228), .ZN(n5533) );
  INV_X1 U7153 ( .A(n5525), .ZN(n5526) );
  NAND2_X1 U7154 ( .A1(n5526), .A2(SI_9_), .ZN(n5527) );
  NAND2_X1 U7155 ( .A1(n6638), .A2(n5535), .ZN(n5530) );
  AOI22_X1 U7156 ( .A1(n5685), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5684), .B2(
        n5528), .ZN(n5529) );
  NAND2_X1 U7157 ( .A1(n5530), .A2(n5529), .ZN(n10039) );
  NAND2_X1 U7158 ( .A1(n7616), .A2(n10039), .ZN(n7900) );
  INV_X1 U7159 ( .A(n7616), .ZN(n7626) );
  OR2_X1 U7160 ( .A1(n10039), .A2(n7626), .ZN(n5531) );
  MUX2_X1 U7161 ( .A(n6642), .B(n10483), .S(n6600), .Z(n5550) );
  XNOR2_X1 U7162 ( .A(n5550), .B(SI_10_), .ZN(n5549) );
  XNOR2_X1 U7163 ( .A(n5554), .B(n5549), .ZN(n6641) );
  NAND2_X1 U7164 ( .A1(n6641), .A2(n5535), .ZN(n5538) );
  INV_X1 U7165 ( .A(n7343), .ZN(n5536) );
  AOI22_X1 U7166 ( .A1(n5685), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5684), .B2(
        n5536), .ZN(n5537) );
  NAND2_X1 U7167 ( .A1(n6569), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5546) );
  INV_X1 U7168 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5539) );
  OR2_X1 U7169 ( .A1(n7811), .A2(n5539), .ZN(n5545) );
  NAND2_X1 U7170 ( .A1(n5540), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5541) );
  AND2_X1 U7171 ( .A1(n5562), .A2(n5541), .ZN(n7623) );
  OR2_X1 U7172 ( .A1(n5402), .A2(n7623), .ZN(n5544) );
  INV_X1 U7173 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5542) );
  OR2_X1 U7174 ( .A1(n6572), .A2(n5542), .ZN(n5543) );
  NAND4_X1 U7175 ( .A1(n5546), .A2(n5545), .A3(n5544), .A4(n5543), .ZN(n8287)
         );
  NAND2_X1 U7176 ( .A1(n7620), .A2(n8287), .ZN(n5548) );
  NOR2_X1 U7177 ( .A1(n7620), .A2(n8287), .ZN(n5547) );
  INV_X1 U7178 ( .A(n5549), .ZN(n5553) );
  INV_X1 U7179 ( .A(n5550), .ZN(n5551) );
  NAND2_X1 U7180 ( .A1(n5551), .A2(SI_10_), .ZN(n5552) );
  MUX2_X1 U7181 ( .A(n6658), .B(n6659), .S(n6600), .Z(n5556) );
  INV_X1 U7182 ( .A(SI_11_), .ZN(n5555) );
  NAND2_X1 U7183 ( .A1(n5556), .A2(n5555), .ZN(n5569) );
  INV_X1 U7184 ( .A(n5556), .ZN(n5557) );
  NAND2_X1 U7185 ( .A1(n5557), .A2(SI_11_), .ZN(n5558) );
  NAND2_X1 U7186 ( .A1(n5569), .A2(n5558), .ZN(n5570) );
  XNOR2_X1 U7187 ( .A(n5571), .B(n5570), .ZN(n6656) );
  NAND2_X1 U7188 ( .A1(n6656), .A2(n5535), .ZN(n5560) );
  AOI22_X1 U7189 ( .A1(n5685), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5684), .B2(
        n7446), .ZN(n5559) );
  NAND2_X1 U7190 ( .A1(n5560), .A2(n5559), .ZN(n7646) );
  NAND2_X1 U7191 ( .A1(n5401), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5567) );
  OR2_X1 U7192 ( .A1(n7811), .A2(n5561), .ZN(n5566) );
  OR2_X1 U7193 ( .A1(n7807), .A2(n7536), .ZN(n5565) );
  NAND2_X1 U7194 ( .A1(n5562), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5563) );
  AND2_X1 U7195 ( .A1(n5575), .A2(n5563), .ZN(n7529) );
  OR2_X1 U7196 ( .A1(n5402), .A2(n7529), .ZN(n5564) );
  OR2_X1 U7197 ( .A1(n7646), .A2(n7629), .ZN(n7915) );
  NAND2_X1 U7198 ( .A1(n7646), .A2(n7629), .ZN(n7913) );
  NAND2_X1 U7199 ( .A1(n7915), .A2(n7913), .ZN(n7636) );
  NAND2_X1 U7200 ( .A1(n7530), .A2(n7636), .ZN(n7532) );
  NAND2_X1 U7201 ( .A1(n7646), .A2(n8162), .ZN(n5568) );
  MUX2_X1 U7202 ( .A(n6715), .B(n10225), .S(n6605), .Z(n5584) );
  XNOR2_X1 U7203 ( .A(n5584), .B(SI_12_), .ZN(n5583) );
  XNOR2_X1 U7204 ( .A(n5586), .B(n5583), .ZN(n6714) );
  NAND2_X1 U7205 ( .A1(n6714), .A2(n5535), .ZN(n5573) );
  AOI22_X1 U7206 ( .A1(n5685), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5684), .B2(
        n7662), .ZN(n5572) );
  NAND2_X1 U7207 ( .A1(n6568), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5580) );
  OR2_X1 U7208 ( .A1(n7807), .A2(n7675), .ZN(n5579) );
  NAND2_X1 U7209 ( .A1(n5575), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5576) );
  AND2_X1 U7210 ( .A1(n5591), .A2(n5576), .ZN(n8164) );
  OR2_X1 U7211 ( .A1(n5402), .A2(n8164), .ZN(n5578) );
  INV_X1 U7212 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7672) );
  OR2_X1 U7213 ( .A1(n6572), .A2(n7672), .ZN(n5577) );
  NAND4_X1 U7214 ( .A1(n5580), .A2(n5579), .A3(n5578), .A4(n5577), .ZN(n8286)
         );
  OR2_X1 U7215 ( .A1(n8166), .A2(n8286), .ZN(n5581) );
  NAND2_X1 U7216 ( .A1(n8166), .A2(n8286), .ZN(n5582) );
  INV_X1 U7217 ( .A(n5584), .ZN(n5585) );
  MUX2_X1 U7218 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6600), .Z(n5600) );
  XNOR2_X1 U7219 ( .A(n5600), .B(SI_13_), .ZN(n5597) );
  XNOR2_X1 U7220 ( .A(n5599), .B(n5597), .ZN(n6733) );
  NAND2_X1 U7221 ( .A1(n6733), .A2(n5535), .ZN(n5588) );
  AOI22_X1 U7222 ( .A1(n5685), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5684), .B2(
        n8305), .ZN(n5587) );
  NAND2_X1 U7223 ( .A1(n5401), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5596) );
  OR2_X1 U7224 ( .A1(n7811), .A2(n8302), .ZN(n5595) );
  OR2_X1 U7225 ( .A1(n7807), .A2(n8296), .ZN(n5594) );
  NAND2_X1 U7226 ( .A1(n5591), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5592) );
  AND2_X1 U7227 ( .A1(n5606), .A2(n5592), .ZN(n8226) );
  OR2_X1 U7228 ( .A1(n5402), .A2(n8226), .ZN(n5593) );
  NAND4_X1 U7229 ( .A1(n5596), .A2(n5595), .A3(n5594), .A4(n5593), .ZN(n8285)
         );
  AND2_X1 U7230 ( .A1(n8228), .A2(n8285), .ZN(n7922) );
  OR2_X1 U7231 ( .A1(n8228), .A2(n8285), .ZN(n7713) );
  INV_X1 U7232 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7233 ( .A1(n5600), .A2(SI_13_), .ZN(n5601) );
  MUX2_X1 U7234 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6605), .Z(n5616) );
  XNOR2_X1 U7235 ( .A(n5616), .B(SI_14_), .ZN(n5613) );
  XNOR2_X1 U7236 ( .A(n5615), .B(n5613), .ZN(n6823) );
  NAND2_X1 U7237 ( .A1(n6823), .A2(n5535), .ZN(n5605) );
  AOI22_X1 U7238 ( .A1(n5685), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5684), .B2(
        n5603), .ZN(n5604) );
  NAND2_X1 U7239 ( .A1(n5401), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5611) );
  OR2_X1 U7240 ( .A1(n7811), .A2(n8628), .ZN(n5610) );
  OR2_X1 U7241 ( .A1(n7807), .A2(n8571), .ZN(n5609) );
  NAND2_X1 U7242 ( .A1(n5606), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5607) );
  AND2_X1 U7243 ( .A1(n5625), .A2(n5607), .ZN(n8570) );
  OR2_X1 U7244 ( .A1(n5402), .A2(n8570), .ZN(n5608) );
  NAND4_X1 U7245 ( .A1(n5611), .A2(n5610), .A3(n5609), .A4(n5608), .ZN(n8548)
         );
  NAND2_X1 U7246 ( .A1(n8716), .A2(n8548), .ZN(n5612) );
  INV_X1 U7247 ( .A(n5613), .ZN(n5614) );
  NAND2_X1 U7248 ( .A1(n5615), .A2(n5614), .ZN(n5618) );
  NAND2_X1 U7249 ( .A1(n5616), .A2(SI_14_), .ZN(n5617) );
  MUX2_X1 U7250 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6600), .Z(n5631) );
  XNOR2_X1 U7251 ( .A(n5631), .B(SI_15_), .ZN(n5619) );
  XNOR2_X1 U7252 ( .A(n5635), .B(n5619), .ZN(n6847) );
  NAND2_X1 U7253 ( .A1(n6847), .A2(n5535), .ZN(n5622) );
  AOI22_X1 U7254 ( .A1(n5685), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5684), .B2(
        n5620), .ZN(n5621) );
  NAND2_X1 U7255 ( .A1(n5401), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5630) );
  OR2_X1 U7256 ( .A1(n7807), .A2(n8332), .ZN(n5629) );
  OR2_X1 U7257 ( .A1(n7811), .A2(n8623), .ZN(n5628) );
  NAND2_X1 U7258 ( .A1(n5625), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5626) );
  AND2_X1 U7259 ( .A1(n5640), .A2(n5626), .ZN(n8268) );
  OR2_X1 U7260 ( .A1(n5402), .A2(n8268), .ZN(n5627) );
  NAND2_X1 U7261 ( .A1(n8709), .A2(n8564), .ZN(n7942) );
  NAND2_X1 U7262 ( .A1(n7936), .A2(n7942), .ZN(n8545) );
  NOR2_X1 U7263 ( .A1(n5632), .A2(n10429), .ZN(n5634) );
  NAND2_X1 U7264 ( .A1(n5632), .A2(n10429), .ZN(n5633) );
  MUX2_X1 U7265 ( .A(n6908), .B(n6909), .S(n6605), .Z(n5646) );
  XNOR2_X1 U7266 ( .A(n5646), .B(SI_16_), .ZN(n5636) );
  XNOR2_X1 U7267 ( .A(n5647), .B(n5636), .ZN(n6907) );
  NAND2_X1 U7268 ( .A1(n6907), .A2(n5535), .ZN(n5639) );
  AOI22_X1 U7269 ( .A1(n5685), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5684), .B2(
        n5637), .ZN(n5638) );
  NAND2_X1 U7270 ( .A1(n5401), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5645) );
  OR2_X1 U7271 ( .A1(n7807), .A2(n8539), .ZN(n5644) );
  INV_X1 U7272 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8620) );
  OR2_X1 U7273 ( .A1(n7811), .A2(n8620), .ZN(n5643) );
  NAND2_X1 U7274 ( .A1(n5640), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5641) );
  AND2_X1 U7275 ( .A1(n5657), .A2(n5641), .ZN(n8540) );
  OR2_X1 U7276 ( .A1(n5402), .A2(n8540), .ZN(n5642) );
  NAND2_X1 U7277 ( .A1(n8703), .A2(n8550), .ZN(n7939) );
  INV_X1 U7278 ( .A(n8703), .ZN(n8187) );
  NAND2_X1 U7279 ( .A1(n5648), .A2(SI_16_), .ZN(n5649) );
  MUX2_X1 U7280 ( .A(n6968), .B(n10403), .S(n6600), .Z(n5651) );
  NAND2_X1 U7281 ( .A1(n5651), .A2(n5650), .ZN(n5663) );
  INV_X1 U7282 ( .A(n5651), .ZN(n5652) );
  NAND2_X1 U7283 ( .A1(n5652), .A2(SI_17_), .ZN(n5653) );
  NAND2_X1 U7284 ( .A1(n5663), .A2(n5653), .ZN(n5664) );
  XNOR2_X1 U7285 ( .A(n5665), .B(n5664), .ZN(n6966) );
  NAND2_X1 U7286 ( .A1(n6966), .A2(n5535), .ZN(n5655) );
  AOI22_X1 U7287 ( .A1(n5685), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5684), .B2(
        n8375), .ZN(n5654) );
  NAND2_X1 U7288 ( .A1(n5401), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5662) );
  OR2_X1 U7289 ( .A1(n7811), .A2(n8617), .ZN(n5661) );
  OR2_X1 U7290 ( .A1(n7807), .A2(n8367), .ZN(n5660) );
  NAND2_X1 U7291 ( .A1(n5657), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5658) );
  AND2_X1 U7292 ( .A1(n5669), .A2(n5658), .ZN(n8194) );
  OR2_X1 U7293 ( .A1(n5402), .A2(n8194), .ZN(n5659) );
  NAND2_X1 U7294 ( .A1(n8697), .A2(n8516), .ZN(n7823) );
  NAND2_X1 U7295 ( .A1(n7822), .A2(n7823), .ZN(n8523) );
  AOI22_X2 U7296 ( .A1(n8526), .A2(n8523), .B1(n8697), .B2(n8537), .ZN(n8514)
         );
  MUX2_X1 U7297 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4506), .Z(n5677) );
  XNOR2_X1 U7298 ( .A(n5677), .B(n10254), .ZN(n5676) );
  XNOR2_X1 U7299 ( .A(n5680), .B(n5676), .ZN(n7016) );
  NAND2_X1 U7300 ( .A1(n7016), .A2(n5535), .ZN(n5668) );
  AOI22_X1 U7301 ( .A1(n5685), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5684), .B2(
        n5666), .ZN(n5667) );
  NAND2_X1 U7302 ( .A1(n5669), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5670) );
  AND2_X1 U7303 ( .A1(n5690), .A2(n5670), .ZN(n8518) );
  OR2_X1 U7304 ( .A1(n5402), .A2(n8518), .ZN(n5674) );
  OR2_X1 U7305 ( .A1(n7807), .A2(n8519), .ZN(n5673) );
  INV_X1 U7306 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8615) );
  OR2_X1 U7307 ( .A1(n7811), .A2(n8615), .ZN(n5672) );
  INV_X1 U7308 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8692) );
  OR2_X1 U7309 ( .A1(n6572), .A2(n8692), .ZN(n5671) );
  NAND4_X1 U7310 ( .A1(n5674), .A2(n5673), .A3(n5672), .A4(n5671), .ZN(n8528)
         );
  NAND2_X1 U7311 ( .A1(n8614), .A2(n8528), .ZN(n5675) );
  INV_X1 U7312 ( .A(n8614), .ZN(n8252) );
  AOI22_X2 U7313 ( .A1(n8514), .A2(n5675), .B1(n8071), .B2(n8252), .ZN(n8504)
         );
  INV_X1 U7314 ( .A(n5676), .ZN(n5679) );
  NAND2_X1 U7315 ( .A1(n5677), .A2(SI_18_), .ZN(n5678) );
  MUX2_X1 U7316 ( .A(n7146), .B(n10214), .S(n6600), .Z(n5681) );
  INV_X1 U7317 ( .A(SI_19_), .ZN(n10488) );
  NAND2_X1 U7318 ( .A1(n5681), .A2(n10488), .ZN(n5700) );
  INV_X1 U7319 ( .A(n5681), .ZN(n5682) );
  NAND2_X1 U7320 ( .A1(n5682), .A2(SI_19_), .ZN(n5683) );
  NAND2_X1 U7321 ( .A1(n5700), .A2(n5683), .ZN(n5697) );
  XNOR2_X1 U7322 ( .A(n5696), .B(n5697), .ZN(n7145) );
  NAND2_X1 U7323 ( .A1(n7145), .A2(n5535), .ZN(n5687) );
  AOI22_X1 U7324 ( .A1(n5685), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n5901), .B2(
        n5684), .ZN(n5686) );
  NAND2_X1 U7325 ( .A1(n5690), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U7326 ( .A1(n5705), .A2(n5691), .ZN(n8507) );
  NAND2_X1 U7327 ( .A1(n5832), .A2(n8507), .ZN(n5695) );
  OR2_X1 U7328 ( .A1(n7807), .A2(n5268), .ZN(n5694) );
  INV_X1 U7329 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8610) );
  OR2_X1 U7330 ( .A1(n7811), .A2(n8610), .ZN(n5693) );
  INV_X1 U7331 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8686) );
  OR2_X1 U7332 ( .A1(n6572), .A2(n8686), .ZN(n5692) );
  OR2_X1 U7333 ( .A1(n8687), .A2(n8517), .ZN(n7959) );
  NAND2_X1 U7334 ( .A1(n8687), .A2(n8517), .ZN(n7958) );
  NAND2_X1 U7335 ( .A1(n7959), .A2(n7958), .ZN(n7842) );
  INV_X1 U7336 ( .A(n8517), .ZN(n8284) );
  AOI22_X2 U7337 ( .A1(n8504), .A2(n7842), .B1(n8687), .B2(n8284), .ZN(n8490)
         );
  INV_X1 U7338 ( .A(n5697), .ZN(n5698) );
  NAND2_X1 U7339 ( .A1(n5699), .A2(n5698), .ZN(n5701) );
  MUX2_X1 U7340 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6605), .Z(n5710) );
  XNOR2_X1 U7341 ( .A(n5710), .B(n10442), .ZN(n5702) );
  XNOR2_X1 U7342 ( .A(n5712), .B(n5702), .ZN(n7294) );
  NAND2_X1 U7343 ( .A1(n7294), .A2(n5535), .ZN(n5704) );
  INV_X1 U7344 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7295) );
  OR2_X1 U7345 ( .A1(n7803), .A2(n7295), .ZN(n5703) );
  NAND2_X1 U7346 ( .A1(n5705), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U7347 ( .A1(n5718), .A2(n5706), .ZN(n8496) );
  AOI22_X1 U7348 ( .A1(n8496), .A2(n5832), .B1(n5401), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5708) );
  AOI22_X1 U7349 ( .A1(n6568), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6569), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U7350 ( .A1(n8211), .A2(n8479), .ZN(n7961) );
  NAND2_X1 U7351 ( .A1(n7953), .A2(n7961), .ZN(n8489) );
  INV_X1 U7352 ( .A(n5710), .ZN(n5711) );
  MUX2_X1 U7353 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6600), .Z(n5724) );
  INV_X1 U7354 ( .A(SI_21_), .ZN(n5713) );
  XNOR2_X1 U7355 ( .A(n5724), .B(n5713), .ZN(n5714) );
  XNOR2_X1 U7356 ( .A(n5726), .B(n5714), .ZN(n7376) );
  NAND2_X1 U7357 ( .A1(n7376), .A2(n5535), .ZN(n5716) );
  INV_X1 U7358 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7377) );
  OR2_X1 U7359 ( .A1(n7803), .A2(n7377), .ZN(n5715) );
  NAND2_X1 U7360 ( .A1(n5718), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7361 ( .A1(n5732), .A2(n5719), .ZN(n8483) );
  NAND2_X1 U7362 ( .A1(n8483), .A2(n5832), .ZN(n5722) );
  AOI22_X1 U7363 ( .A1(n6568), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n6569), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U7364 ( .A1(n5401), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7365 ( .A1(n8082), .A2(n8493), .ZN(n7962) );
  NAND2_X1 U7366 ( .A1(n7954), .A2(n7962), .ZN(n8481) );
  NOR2_X1 U7367 ( .A1(n5724), .A2(SI_21_), .ZN(n5725) );
  MUX2_X1 U7368 ( .A(n7466), .B(n10415), .S(n4506), .Z(n5727) );
  INV_X1 U7369 ( .A(SI_22_), .ZN(n10279) );
  NAND2_X1 U7370 ( .A1(n5727), .A2(n10279), .ZN(n5737) );
  INV_X1 U7371 ( .A(n5727), .ZN(n5728) );
  NAND2_X1 U7372 ( .A1(n5728), .A2(SI_22_), .ZN(n5729) );
  NAND2_X1 U7373 ( .A1(n5737), .A2(n5729), .ZN(n5738) );
  XNOR2_X1 U7374 ( .A(n5739), .B(n5738), .ZN(n7464) );
  NAND2_X1 U7375 ( .A1(n7464), .A2(n5535), .ZN(n5731) );
  OR2_X1 U7376 ( .A1(n7803), .A2(n7466), .ZN(n5730) );
  NAND2_X1 U7377 ( .A1(n5732), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7378 ( .A1(n5745), .A2(n5733), .ZN(n8471) );
  NAND2_X1 U7379 ( .A1(n8471), .A2(n5832), .ZN(n5736) );
  AOI22_X1 U7380 ( .A1(n6568), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n6569), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7381 ( .A1(n5401), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U7382 ( .A1(n8470), .A2(n8480), .ZN(n7969) );
  INV_X1 U7383 ( .A(n8480), .ZN(n8283) );
  MUX2_X1 U7384 ( .A(n7513), .B(n10489), .S(n6600), .Z(n5740) );
  NAND2_X1 U7385 ( .A1(n5740), .A2(n10251), .ZN(n5755) );
  INV_X1 U7386 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U7387 ( .A1(n5741), .A2(SI_23_), .ZN(n5742) );
  XNOR2_X1 U7388 ( .A(n5754), .B(n5753), .ZN(n7511) );
  NAND2_X1 U7389 ( .A1(n7511), .A2(n5535), .ZN(n5744) );
  OR2_X1 U7390 ( .A1(n7803), .A2(n7513), .ZN(n5743) );
  NAND2_X1 U7391 ( .A1(n5745), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U7392 ( .A1(n5762), .A2(n5746), .ZN(n8462) );
  NAND2_X1 U7393 ( .A1(n8462), .A2(n5832), .ZN(n5751) );
  INV_X1 U7394 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U7395 ( .A1(n6568), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U7396 ( .A1(n6569), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5747) );
  OAI211_X1 U7397 ( .C1(n8667), .C2(n6572), .A(n5748), .B(n5747), .ZN(n5749)
         );
  INV_X1 U7398 ( .A(n5749), .ZN(n5750) );
  NOR2_X1 U7399 ( .A1(n8668), .A2(n8282), .ZN(n5752) );
  INV_X1 U7400 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7594) );
  MUX2_X1 U7401 ( .A(n7584), .B(n7594), .S(n4506), .Z(n5757) );
  INV_X1 U7402 ( .A(SI_24_), .ZN(n10289) );
  NAND2_X1 U7403 ( .A1(n5757), .A2(n10289), .ZN(n5772) );
  INV_X1 U7404 ( .A(n5757), .ZN(n5758) );
  NAND2_X1 U7405 ( .A1(n5758), .A2(SI_24_), .ZN(n5759) );
  XNOR2_X1 U7406 ( .A(n5771), .B(n5770), .ZN(n7583) );
  NOR2_X1 U7407 ( .A1(n7803), .A2(n7584), .ZN(n5760) );
  NAND2_X1 U7408 ( .A1(n5762), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7409 ( .A1(n5781), .A2(n5763), .ZN(n8448) );
  NAND2_X1 U7410 ( .A1(n8448), .A2(n5832), .ZN(n5768) );
  INV_X1 U7411 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U7412 ( .A1(n6568), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7413 ( .A1(n6569), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5764) );
  OAI211_X1 U7414 ( .C1(n8661), .C2(n6572), .A(n5765), .B(n5764), .ZN(n5766)
         );
  INV_X1 U7415 ( .A(n5766), .ZN(n5767) );
  NOR2_X1 U7416 ( .A1(n8590), .A2(n8460), .ZN(n5769) );
  INV_X1 U7417 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7685) );
  INV_X1 U7418 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7729) );
  MUX2_X1 U7419 ( .A(n7685), .B(n7729), .S(n4506), .Z(n5774) );
  INV_X1 U7420 ( .A(SI_25_), .ZN(n10409) );
  NAND2_X1 U7421 ( .A1(n5774), .A2(n10409), .ZN(n5801) );
  INV_X1 U7422 ( .A(n5774), .ZN(n5775) );
  NAND2_X1 U7423 ( .A1(n5775), .A2(SI_25_), .ZN(n5776) );
  XNOR2_X1 U7424 ( .A(n5789), .B(n5788), .ZN(n7684) );
  NAND2_X1 U7425 ( .A1(n7684), .A2(n5535), .ZN(n5778) );
  OR2_X1 U7426 ( .A1(n7803), .A2(n7685), .ZN(n5777) );
  INV_X1 U7427 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7428 ( .A1(n5781), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5782) );
  NAND2_X1 U7429 ( .A1(n5811), .A2(n5782), .ZN(n8437) );
  NAND2_X1 U7430 ( .A1(n8437), .A2(n5832), .ZN(n5787) );
  INV_X1 U7431 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U7432 ( .A1(n6569), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7433 ( .A1(n6568), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5783) );
  OAI211_X1 U7434 ( .C1(n6572), .C2(n8654), .A(n5784), .B(n5783), .ZN(n5785)
         );
  INV_X1 U7435 ( .A(n5785), .ZN(n5786) );
  NAND2_X1 U7436 ( .A1(n8655), .A2(n8446), .ZN(n7984) );
  NAND2_X1 U7437 ( .A1(n7987), .A2(n7984), .ZN(n8439) );
  INV_X1 U7438 ( .A(n8655), .ZN(n8587) );
  NAND2_X1 U7439 ( .A1(n5803), .A2(n5801), .ZN(n5793) );
  INV_X1 U7440 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7699) );
  INV_X1 U7441 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7710) );
  MUX2_X1 U7442 ( .A(n7699), .B(n7710), .S(n6600), .Z(n5790) );
  NAND2_X1 U7443 ( .A1(n5790), .A2(n10427), .ZN(n5800) );
  INV_X1 U7444 ( .A(n5790), .ZN(n5791) );
  NAND2_X1 U7445 ( .A1(n5791), .A2(SI_26_), .ZN(n5823) );
  AND2_X1 U7446 ( .A1(n5800), .A2(n5823), .ZN(n5792) );
  NOR2_X1 U7447 ( .A1(n7803), .A2(n7699), .ZN(n5794) );
  XNOR2_X1 U7448 ( .A(n5811), .B(P2_REG3_REG_26__SCAN_IN), .ZN(n8421) );
  NAND2_X1 U7449 ( .A1(n8421), .A2(n5832), .ZN(n5799) );
  INV_X1 U7450 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U7451 ( .A1(n6568), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7452 ( .A1(n6569), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5795) );
  OAI211_X1 U7453 ( .C1(n8648), .C2(n6572), .A(n5796), .B(n5795), .ZN(n5797)
         );
  INV_X1 U7454 ( .A(n5797), .ZN(n5798) );
  INV_X1 U7455 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7749) );
  MUX2_X1 U7456 ( .A(n7732), .B(n7749), .S(n6600), .Z(n5805) );
  INV_X1 U7457 ( .A(SI_27_), .ZN(n5804) );
  NAND2_X1 U7458 ( .A1(n5805), .A2(n5804), .ZN(n5826) );
  INV_X1 U7459 ( .A(n5805), .ZN(n5806) );
  NAND2_X1 U7460 ( .A1(n5806), .A2(SI_27_), .ZN(n5807) );
  NAND2_X1 U7461 ( .A1(n7731), .A2(n5535), .ZN(n5810) );
  OR2_X1 U7462 ( .A1(n7803), .A2(n7732), .ZN(n5809) );
  INV_X1 U7463 ( .A(n5811), .ZN(n5812) );
  INV_X1 U7464 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10456) );
  INV_X1 U7465 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8099) );
  INV_X1 U7466 ( .A(n5813), .ZN(n5814) );
  NAND2_X1 U7467 ( .A1(n5814), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7468 ( .A1(n5830), .A2(n5815), .ZN(n8417) );
  NAND2_X1 U7469 ( .A1(n8417), .A2(n5832), .ZN(n5820) );
  INV_X1 U7470 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U7471 ( .A1(n6569), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7472 ( .A1(n6568), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5816) );
  OAI211_X1 U7473 ( .C1(n8641), .C2(n6572), .A(n5817), .B(n5816), .ZN(n5818)
         );
  INV_X1 U7474 ( .A(n5818), .ZN(n5819) );
  INV_X1 U7475 ( .A(n8642), .ZN(n5821) );
  AND2_X1 U7476 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  MUX2_X1 U7477 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6600), .Z(n6560) );
  XNOR2_X1 U7478 ( .A(n6560), .B(n10485), .ZN(n6558) );
  NAND2_X1 U7479 ( .A1(n7791), .A2(n5535), .ZN(n5829) );
  INV_X1 U7480 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7736) );
  OR2_X1 U7481 ( .A1(n7803), .A2(n7736), .ZN(n5828) );
  NAND2_X1 U7482 ( .A1(n5830), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U7483 ( .A1(n8033), .A2(n5831), .ZN(n8139) );
  NAND2_X1 U7484 ( .A1(n8139), .A2(n5832), .ZN(n5838) );
  INV_X1 U7485 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U7486 ( .A1(n6568), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7487 ( .A1(n6569), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5833) );
  OAI211_X1 U7488 ( .C1(n5835), .C2(n6572), .A(n5834), .B(n5833), .ZN(n5836)
         );
  INV_X1 U7489 ( .A(n5836), .ZN(n5837) );
  XNOR2_X1 U7490 ( .A(n6557), .B(n5839), .ZN(n5846) );
  NAND2_X1 U7491 ( .A1(n5840), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5841) );
  MUX2_X1 U7492 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5841), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5843) );
  INV_X1 U7493 ( .A(n7852), .ZN(n6804) );
  NAND2_X1 U7494 ( .A1(n6805), .A2(n6804), .ZN(n5845) );
  NAND2_X1 U7495 ( .A1(n5901), .A2(n8027), .ZN(n5844) );
  NAND2_X1 U7496 ( .A1(n5846), .A2(n9981), .ZN(n5856) );
  XNOR2_X1 U7497 ( .A(n5847), .B(n8025), .ZN(n5853) );
  INV_X1 U7498 ( .A(n5853), .ZN(n6816) );
  OR2_X1 U7499 ( .A1(n8033), .A2(n5402), .ZN(n7814) );
  INV_X1 U7500 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7501 ( .A1(n6569), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7502 ( .A1(n6568), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5848) );
  OAI211_X1 U7503 ( .C1(n6572), .C2(n5850), .A(n5849), .B(n5848), .ZN(n5851)
         );
  INV_X1 U7504 ( .A(n5851), .ZN(n5852) );
  XNOR2_X1 U7505 ( .A(n7585), .B(P2_B_REG_SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7506 ( .A1(n5857), .A2(n7686), .ZN(n5859) );
  NAND2_X1 U7507 ( .A1(n7700), .A2(n7585), .ZN(n6626) );
  NOR2_X1 U7508 ( .A1(n7852), .A2(n7465), .ZN(n5900) );
  NAND2_X1 U7509 ( .A1(n5900), .A2(n7850), .ZN(n5860) );
  OAI21_X1 U7510 ( .B1(n6802), .B2(n5920), .A(n5914), .ZN(n5875) );
  NAND2_X1 U7511 ( .A1(n8012), .A2(n8021), .ZN(n5861) );
  NOR2_X1 U7512 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5865) );
  NOR4_X1 U7513 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5864) );
  NOR4_X1 U7514 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5863) );
  NOR4_X1 U7515 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5862) );
  NAND4_X1 U7516 ( .A1(n5865), .A2(n5864), .A3(n5863), .A4(n5862), .ZN(n5871)
         );
  NOR4_X1 U7517 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5869) );
  NOR4_X1 U7518 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5868) );
  NOR4_X1 U7519 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5867) );
  NOR4_X1 U7520 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5866) );
  NAND4_X1 U7521 ( .A1(n5869), .A2(n5868), .A3(n5867), .A4(n5866), .ZN(n5870)
         );
  NOR2_X1 U7522 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  NAND2_X1 U7523 ( .A1(n7686), .A2(n7700), .ZN(n6629) );
  NAND2_X1 U7524 ( .A1(n5915), .A2(n5913), .ZN(n5874) );
  NAND2_X1 U7525 ( .A1(n6874), .A2(n6871), .ZN(n6870) );
  NAND2_X1 U7526 ( .A1(n6870), .A2(n7858), .ZN(n9993) );
  INV_X1 U7527 ( .A(n4612), .ZN(n9994) );
  NAND2_X1 U7528 ( .A1(n9993), .A2(n9994), .ZN(n5877) );
  NAND2_X1 U7529 ( .A1(n5877), .A2(n7863), .ZN(n9973) );
  NAND2_X1 U7530 ( .A1(n9973), .A2(n9974), .ZN(n5878) );
  OR2_X1 U7531 ( .A1(n9984), .A2(n10011), .ZN(n7870) );
  NAND2_X1 U7532 ( .A1(n5878), .A2(n7870), .ZN(n6911) );
  INV_X1 U7533 ( .A(n7824), .ZN(n7875) );
  NAND2_X1 U7534 ( .A1(n6911), .A2(n7875), .ZN(n5879) );
  NAND2_X1 U7535 ( .A1(n5879), .A2(n7890), .ZN(n6973) );
  NAND2_X1 U7536 ( .A1(n8291), .A2(n7023), .ZN(n7879) );
  AND2_X1 U7537 ( .A1(n8290), .A2(n10021), .ZN(n7881) );
  OR2_X1 U7538 ( .A1(n8290), .A2(n10021), .ZN(n7882) );
  OR2_X1 U7539 ( .A1(n8291), .A2(n7023), .ZN(n7207) );
  NAND2_X1 U7540 ( .A1(n7882), .A2(n7207), .ZN(n7889) );
  INV_X1 U7541 ( .A(n7881), .ZN(n7887) );
  NAND2_X1 U7542 ( .A1(n7889), .A2(n7887), .ZN(n5880) );
  INV_X1 U7543 ( .A(n7321), .ZN(n10026) );
  OR2_X1 U7544 ( .A1(n8289), .A2(n10026), .ZN(n7898) );
  NAND2_X1 U7545 ( .A1(n8289), .A2(n10026), .ZN(n7410) );
  NAND2_X1 U7546 ( .A1(n7898), .A2(n7410), .ZN(n7829) );
  NAND2_X1 U7547 ( .A1(n8288), .A2(n10031), .ZN(n7886) );
  AND2_X1 U7548 ( .A1(n7410), .A2(n7886), .ZN(n7904) );
  OR2_X1 U7549 ( .A1(n8288), .A2(n10031), .ZN(n7899) );
  NAND2_X1 U7550 ( .A1(n7450), .A2(n7834), .ZN(n7452) );
  NAND2_X1 U7551 ( .A1(n7452), .A2(n7903), .ZN(n7497) );
  OAI21_X1 U7552 ( .B1(n7497), .B2(n7911), .A(n7908), .ZN(n7535) );
  INV_X1 U7553 ( .A(n7636), .ZN(n7836) );
  NAND2_X1 U7554 ( .A1(n7535), .A2(n7836), .ZN(n5881) );
  NAND2_X1 U7555 ( .A1(n5881), .A2(n7913), .ZN(n7669) );
  XNOR2_X1 U7556 ( .A(n8166), .B(n8050), .ZN(n7838) );
  OR2_X1 U7557 ( .A1(n8166), .A2(n8050), .ZN(n7920) );
  INV_X1 U7558 ( .A(n8285), .ZN(n8562) );
  INV_X1 U7559 ( .A(n8228), .ZN(n7925) );
  OR2_X1 U7560 ( .A1(n8716), .A2(n8223), .ZN(n7928) );
  NAND2_X1 U7561 ( .A1(n8569), .A2(n7928), .ZN(n5882) );
  NAND2_X1 U7562 ( .A1(n8716), .A2(n8223), .ZN(n7932) );
  NAND2_X1 U7563 ( .A1(n5882), .A2(n7932), .ZN(n8544) );
  INV_X1 U7564 ( .A(n8544), .ZN(n5883) );
  NAND2_X1 U7565 ( .A1(n5884), .A2(n7939), .ZN(n8524) );
  NAND2_X1 U7566 ( .A1(n8614), .A2(n8071), .ZN(n7949) );
  INV_X1 U7567 ( .A(n7961), .ZN(n5885) );
  INV_X1 U7568 ( .A(n7954), .ZN(n7963) );
  AOI21_X1 U7569 ( .B1(n8482), .B2(n7962), .A(n7963), .ZN(n8469) );
  INV_X1 U7570 ( .A(n7969), .ZN(n5886) );
  OAI21_X1 U7571 ( .B1(n8469), .B2(n5886), .A(n7968), .ZN(n8456) );
  NOR2_X1 U7572 ( .A1(n8456), .A2(n7973), .ZN(n8450) );
  NAND2_X1 U7573 ( .A1(n8662), .A2(n8460), .ZN(n7983) );
  NAND2_X1 U7574 ( .A1(n8668), .A2(n8467), .ZN(n7821) );
  NAND2_X1 U7575 ( .A1(n7983), .A2(n7821), .ZN(n7978) );
  OAI21_X1 U7576 ( .B1(n8450), .B2(n7978), .A(n7980), .ZN(n8438) );
  INV_X1 U7577 ( .A(n7987), .ZN(n5887) );
  NOR2_X1 U7578 ( .A1(n8642), .A2(n8426), .ZN(n7996) );
  XNOR2_X1 U7579 ( .A(n6567), .B(n7820), .ZN(n5926) );
  INV_X1 U7580 ( .A(n8021), .ZN(n5888) );
  NAND2_X1 U7581 ( .A1(n8012), .A2(n5888), .ZN(n6736) );
  OAI21_X1 U7582 ( .B1(n7852), .B2(n8027), .A(n7850), .ZN(n5889) );
  INV_X1 U7583 ( .A(n5889), .ZN(n5890) );
  AND2_X1 U7584 ( .A1(n10042), .A2(n5890), .ZN(n5891) );
  OAI22_X1 U7585 ( .A1(n5926), .A2(n8626), .B1(n8007), .B2(n8609), .ZN(n5892)
         );
  INV_X1 U7586 ( .A(n5892), .ZN(n5894) );
  INV_X1 U7587 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5893) );
  INV_X1 U7588 ( .A(n5903), .ZN(n5897) );
  NOR2_X1 U7589 ( .A1(n5898), .A2(n5897), .ZN(n6744) );
  NAND2_X1 U7590 ( .A1(n6744), .A2(n6746), .ZN(n6758) );
  NAND3_X1 U7591 ( .A1(n7856), .A2(n5901), .A3(n5900), .ZN(n6739) );
  AND2_X1 U7592 ( .A1(n6736), .A2(n6739), .ZN(n5902) );
  NAND3_X1 U7593 ( .A1(n6802), .A2(n5915), .A3(n5903), .ZN(n6748) );
  INV_X1 U7594 ( .A(n6746), .ZN(n5904) );
  AND2_X1 U7595 ( .A1(n8009), .A2(n10042), .ZN(n5905) );
  NAND2_X1 U7596 ( .A1(n6739), .A2(n5905), .ZN(n6753) );
  INV_X1 U7597 ( .A(n8019), .ZN(n9992) );
  NAND2_X1 U7598 ( .A1(n10040), .A2(n9992), .ZN(n8443) );
  NAND2_X1 U7599 ( .A1(n6753), .A2(n8443), .ZN(n6738) );
  NAND2_X1 U7600 ( .A1(n6755), .A2(n6738), .ZN(n5906) );
  OAI22_X1 U7601 ( .A1(n5926), .A2(n8712), .B1(n8007), .B2(n8683), .ZN(n5908)
         );
  INV_X1 U7602 ( .A(n5908), .ZN(n5910) );
  OR2_X1 U7603 ( .A1(n10048), .A2(n5835), .ZN(n5909) );
  OR2_X1 U7604 ( .A1(n6802), .A2(n5913), .ZN(n5918) );
  OR2_X1 U7605 ( .A1(n5915), .A2(n5914), .ZN(n5917) );
  NAND2_X1 U7606 ( .A1(n6802), .A2(n5915), .ZN(n5916) );
  NAND4_X1 U7607 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(n5922)
         );
  NAND2_X1 U7608 ( .A1(n5921), .A2(n9999), .ZN(n5929) );
  NAND2_X1 U7609 ( .A1(n8019), .A2(n6805), .ZN(n6872) );
  NAND2_X1 U7610 ( .A1(n7502), .A2(n6872), .ZN(n9995) );
  INV_X1 U7611 ( .A(n5922), .ZN(n5923) );
  INV_X1 U7612 ( .A(n8443), .ZN(n8566) );
  AOI22_X1 U7613 ( .A1(n8144), .A2(n8555), .B1(n8554), .B2(n8139), .ZN(n5925)
         );
  OAI21_X1 U7614 ( .B1(n5926), .B2(n8558), .A(n5096), .ZN(n5927) );
  INV_X1 U7615 ( .A(n5927), .ZN(n5928) );
  NAND2_X1 U7616 ( .A1(n5929), .A2(n5928), .ZN(P2_U3205) );
  NOR2_X1 U7617 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5930) );
  NAND3_X1 U7618 ( .A1(n6043), .A2(n6090), .A3(n5930), .ZN(n6129) );
  INV_X1 U7619 ( .A(n6129), .ZN(n5932) );
  NAND2_X1 U7620 ( .A1(n5932), .A2(n5931), .ZN(n6155) );
  NOR2_X1 U7621 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5935) );
  NAND4_X1 U7622 ( .A1(n5935), .A2(n5934), .A3(n5933), .A4(n6211), .ZN(n5936)
         );
  NOR2_X1 U7623 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5940) );
  NOR2_X1 U7624 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5939) );
  NOR2_X1 U7625 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5938) );
  NOR2_X1 U7626 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5937) );
  NAND4_X1 U7627 ( .A1(n5940), .A2(n5939), .A3(n5938), .A4(n5937), .ZN(n5943)
         );
  NAND4_X1 U7628 ( .A1(n5941), .A2(n5958), .A3(n5967), .A4(n5974), .ZN(n5942)
         );
  NAND2_X1 U7629 ( .A1(n5945), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5944) );
  MUX2_X1 U7630 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5944), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5948) );
  NAND2_X1 U7631 ( .A1(n7464), .A2(n8841), .ZN(n5952) );
  NAND2_X1 U7632 ( .A1(n6066), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5951) );
  NAND2_X1 U7633 ( .A1(n5969), .A2(n5971), .ZN(n5973) );
  INV_X1 U7634 ( .A(n5973), .ZN(n5956) );
  NAND2_X1 U7635 ( .A1(n5956), .A2(n5955), .ZN(n5962) );
  NAND2_X1 U7636 ( .A1(n5959), .A2(n5958), .ZN(n5961) );
  OR2_X1 U7637 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  NAND2_X1 U7638 ( .A1(n5961), .A2(n5960), .ZN(n6506) );
  NAND2_X1 U7639 ( .A1(n5962), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5964) );
  NOR2_X1 U7640 ( .A1(n6506), .A2(n7596), .ZN(n5965) );
  NAND2_X2 U7641 ( .A1(n6509), .A2(n5965), .ZN(n6019) );
  NAND2_X1 U7642 ( .A1(n6342), .A2(n5967), .ZN(n5968) );
  NAND2_X1 U7643 ( .A1(n5968), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6357) );
  INV_X1 U7644 ( .A(n5969), .ZN(n5970) );
  NAND2_X1 U7645 ( .A1(n5970), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7646 ( .A1(n8919), .A2(n8914), .ZN(n5981) );
  NAND2_X1 U7647 ( .A1(n6526), .A2(n5981), .ZN(n5978) );
  NAND2_X1 U7648 ( .A1(n5975), .A2(n5974), .ZN(n5976) );
  NAND2_X1 U7649 ( .A1(n5978), .A2(n6723), .ZN(n5979) );
  INV_X1 U7650 ( .A(n5981), .ZN(n7076) );
  INV_X1 U7651 ( .A(n5986), .ZN(n5983) );
  NAND2_X1 U7652 ( .A1(n5983), .A2(n5982), .ZN(n9627) );
  XNOR2_X2 U7653 ( .A(n5985), .B(n5984), .ZN(n7790) );
  NAND2_X1 U7654 ( .A1(n5986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7655 ( .A1(n8868), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5993) );
  INV_X2 U7656 ( .A(n7790), .ZN(n5989) );
  NAND2_X1 U7657 ( .A1(n4521), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5992) );
  AND2_X4 U7658 ( .A1(n5989), .A2(n5988), .ZN(n6073) );
  NAND2_X1 U7659 ( .A1(n6117), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7660 ( .A1(n6159), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7661 ( .A1(n6319), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6334) );
  XNOR2_X1 U7662 ( .A(P1_REG3_REG_22__SCAN_IN), .B(n6411), .ZN(n9481) );
  NAND2_X1 U7663 ( .A1(n6073), .A2(n9481), .ZN(n5991) );
  NAND2_X1 U7664 ( .A1(n4517), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5990) );
  NAND4_X1 U7665 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n9462)
         );
  AOI22_X1 U7666 ( .A1(n9584), .A2(n6502), .B1(n6419), .B2(n9462), .ZN(n5994)
         );
  XNOR2_X1 U7667 ( .A(n5994), .B(n4512), .ZN(n8804) );
  INV_X1 U7668 ( .A(n8804), .ZN(n6408) );
  NAND2_X1 U7669 ( .A1(n7145), .A2(n8841), .ZN(n5997) );
  AOI22_X1 U7670 ( .A1(n9357), .A2(n6360), .B1(n6066), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n5996) );
  NOR2_X1 U7671 ( .A1(n6365), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5998) );
  OR2_X1 U7672 ( .A1(n6378), .A2(n5998), .ZN(n9523) );
  INV_X1 U7673 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9524) );
  NAND2_X1 U7674 ( .A1(n4517), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7675 ( .A1(n4520), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5999) );
  OAI211_X1 U7676 ( .C1(n6074), .C2(n9524), .A(n6000), .B(n5999), .ZN(n6001)
         );
  INV_X1 U7677 ( .A(n6001), .ZN(n6002) );
  OAI21_X1 U7678 ( .B1(n9523), .B2(n6370), .A(n6002), .ZN(n9137) );
  AND2_X1 U7679 ( .A1(n9137), .A2(n6449), .ZN(n6003) );
  AOI21_X1 U7680 ( .B1(n9603), .B2(n6419), .A(n6003), .ZN(n6375) );
  INV_X2 U7681 ( .A(n4891), .ZN(n6502) );
  NAND2_X1 U7682 ( .A1(n9603), .A2(n6502), .ZN(n6005) );
  NAND2_X1 U7683 ( .A1(n9137), .A2(n6419), .ZN(n6004) );
  NAND2_X1 U7684 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  XNOR2_X1 U7685 ( .A(n6006), .B(n4512), .ZN(n6373) );
  INV_X1 U7686 ( .A(n6373), .ZN(n6374) );
  NAND2_X1 U7687 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6007) );
  XNOR2_X1 U7688 ( .A(n6007), .B(P1_IR_REG_1__SCAN_IN), .ZN(n9158) );
  INV_X1 U7689 ( .A(n9158), .ZN(n6008) );
  NAND2_X1 U7690 ( .A1(n4523), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7691 ( .A1(n6025), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6012) );
  INV_X1 U7692 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U7693 ( .A1(n6047), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6010) );
  OR2_X1 U7694 ( .A1(n6083), .A2(n9738), .ZN(n6018) );
  AND2_X1 U7695 ( .A1(n6018), .A2(n6017), .ZN(n6039) );
  NAND2_X1 U7696 ( .A1(n6038), .A2(n6039), .ZN(n6831) );
  INV_X1 U7697 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9662) );
  OR2_X1 U7698 ( .A1(n6019), .A2(n9662), .ZN(n6031) );
  INV_X1 U7699 ( .A(SI_0_), .ZN(n6021) );
  INV_X1 U7700 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6020) );
  OAI21_X1 U7701 ( .B1(n7798), .B2(n6021), .A(n6020), .ZN(n6023) );
  AND2_X1 U7702 ( .A1(n6023), .A2(n6022), .ZN(n9636) );
  INV_X1 U7703 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7704 ( .A1(n6025), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7705 ( .A1(n6073), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7706 ( .A1(n4519), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6026) );
  AND4_X2 U7707 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .ZN(n7178)
         );
  NAND3_X1 U7708 ( .A1(n6031), .A2(n6035), .A3(n6030), .ZN(n6827) );
  INV_X1 U7709 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10239) );
  INV_X1 U7710 ( .A(n7178), .ZN(n6032) );
  NAND2_X1 U7711 ( .A1(n6449), .A2(n6032), .ZN(n6033) );
  OAI211_X1 U7712 ( .C1(n10239), .C2(n6019), .A(n6034), .B(n6033), .ZN(n6826)
         );
  NAND2_X1 U7713 ( .A1(n6827), .A2(n6826), .ZN(n6037) );
  NAND2_X1 U7714 ( .A1(n6035), .A2(n6081), .ZN(n6036) );
  NAND2_X1 U7715 ( .A1(n6037), .A2(n6036), .ZN(n6834) );
  NAND2_X1 U7716 ( .A1(n6831), .A2(n6834), .ZN(n6042) );
  INV_X1 U7717 ( .A(n6038), .ZN(n6041) );
  INV_X1 U7718 ( .A(n6039), .ZN(n6040) );
  NAND2_X1 U7719 ( .A1(n6041), .A2(n6040), .ZN(n6832) );
  NAND2_X1 U7720 ( .A1(n6042), .A2(n6832), .ZN(n6852) );
  INV_X1 U7721 ( .A(n6852), .ZN(n6060) );
  NAND2_X1 U7722 ( .A1(n6066), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7723 ( .A1(n6360), .A2(n9179), .ZN(n6044) );
  NAND2_X1 U7724 ( .A1(n6046), .A2(n9745), .ZN(n6053) );
  NAND2_X1 U7725 ( .A1(n6073), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U7726 ( .A1(n6047), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7727 ( .A1(n6025), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6050) );
  INV_X1 U7728 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6048) );
  OR2_X1 U7729 ( .A1(n6074), .A2(n6048), .ZN(n6049) );
  AND4_X2 U7730 ( .A1(n6052), .A2(n6051), .A3(n6050), .A4(n6049), .ZN(n7063)
         );
  XNOR2_X1 U7731 ( .A(n6055), .B(n6054), .ZN(n6061) );
  INV_X1 U7732 ( .A(n9745), .ZN(n7101) );
  OR2_X1 U7733 ( .A1(n6450), .A2(n7101), .ZN(n6058) );
  OR2_X1 U7734 ( .A1(n4518), .A2(n7063), .ZN(n6057) );
  NAND2_X1 U7735 ( .A1(n6058), .A2(n6057), .ZN(n6062) );
  XNOR2_X1 U7736 ( .A(n6061), .B(n6062), .ZN(n6851) );
  INV_X1 U7737 ( .A(n6851), .ZN(n6059) );
  NAND2_X1 U7738 ( .A1(n6060), .A2(n6059), .ZN(n6853) );
  INV_X1 U7739 ( .A(n6061), .ZN(n6064) );
  INV_X1 U7740 ( .A(n6062), .ZN(n6063) );
  NAND2_X1 U7741 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  NAND2_X1 U7742 ( .A1(n6853), .A2(n6065), .ZN(n6884) );
  NAND2_X1 U7743 ( .A1(n6066), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6071) );
  INV_X1 U7744 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U7745 ( .A1(n6092), .A2(n6067), .ZN(n6068) );
  NAND2_X1 U7746 ( .A1(n6068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6069) );
  XNOR2_X1 U7747 ( .A(n6069), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9193) );
  NAND2_X1 U7748 ( .A1(n6360), .A2(n9193), .ZN(n6070) );
  OAI211_X1 U7749 ( .C1(n6154), .C2(n6617), .A(n6071), .B(n6070), .ZN(n7075)
         );
  INV_X1 U7750 ( .A(n7075), .ZN(n6072) );
  INV_X1 U7751 ( .A(n6083), .ZN(n6125) );
  INV_X1 U7752 ( .A(n6125), .ZN(n6450) );
  NAND2_X1 U7753 ( .A1(n4520), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6078) );
  INV_X1 U7754 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6886) );
  NAND2_X1 U7755 ( .A1(n6073), .A2(n6886), .ZN(n6077) );
  NAND2_X1 U7756 ( .A1(n6025), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7757 ( .A1(n8845), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6075) );
  OR2_X1 U7758 ( .A1(n6450), .A2(n7085), .ZN(n6079) );
  NAND2_X1 U7759 ( .A1(n6080), .A2(n6079), .ZN(n6082) );
  OR2_X1 U7760 ( .A1(n6083), .A2(n6072), .ZN(n6085) );
  OR2_X1 U7761 ( .A1(n4518), .A2(n7085), .ZN(n6084) );
  NAND2_X1 U7762 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  XNOR2_X1 U7763 ( .A(n6088), .B(n6086), .ZN(n6885) );
  INV_X1 U7764 ( .A(n6086), .ZN(n6087) );
  NAND2_X1 U7765 ( .A1(n6088), .A2(n6087), .ZN(n6089) );
  OR2_X1 U7766 ( .A1(n6090), .A2(n9626), .ZN(n6091) );
  AND2_X1 U7767 ( .A1(n6092), .A2(n6091), .ZN(n6094) );
  INV_X1 U7768 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7769 ( .A1(n6094), .A2(n6093), .ZN(n6113) );
  INV_X1 U7770 ( .A(n6094), .ZN(n6095) );
  NAND2_X1 U7771 ( .A1(n6095), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6096) );
  AOI22_X1 U7772 ( .A1(n6066), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6360), .B2(
        n9676), .ZN(n6098) );
  OR2_X1 U7773 ( .A1(n6154), .A2(n6620), .ZN(n6097) );
  NAND2_X1 U7774 ( .A1(n6098), .A2(n6097), .ZN(n9757) );
  NAND2_X1 U7775 ( .A1(n6502), .A2(n9757), .ZN(n6105) );
  NAND2_X1 U7776 ( .A1(n4521), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7777 ( .A1(n8868), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6102) );
  NOR2_X1 U7778 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6099) );
  NOR2_X1 U7779 ( .A1(n6117), .A2(n6099), .ZN(n7091) );
  NAND2_X1 U7780 ( .A1(n6073), .A2(n7091), .ZN(n6101) );
  NAND2_X1 U7781 ( .A1(n6025), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6100) );
  OR2_X1 U7783 ( .A1(n6450), .A2(n7127), .ZN(n6104) );
  NAND2_X1 U7784 ( .A1(n6105), .A2(n6104), .ZN(n6106) );
  XNOR2_X1 U7785 ( .A(n6106), .B(n4512), .ZN(n6111) );
  INV_X1 U7786 ( .A(n9757), .ZN(n7126) );
  OR2_X1 U7787 ( .A1(n6304), .A2(n7126), .ZN(n6108) );
  OR2_X1 U7788 ( .A1(n4518), .A2(n7127), .ZN(n6107) );
  NAND2_X1 U7789 ( .A1(n6108), .A2(n6107), .ZN(n6110) );
  XNOR2_X1 U7790 ( .A(n6111), .B(n6110), .ZN(n7012) );
  INV_X1 U7791 ( .A(n7012), .ZN(n6109) );
  NAND2_X1 U7792 ( .A1(n6111), .A2(n6110), .ZN(n6112) );
  NAND2_X1 U7793 ( .A1(n7010), .A2(n6112), .ZN(n7043) );
  OR2_X1 U7794 ( .A1(n6610), .A2(n6154), .ZN(n6116) );
  NAND2_X1 U7795 ( .A1(n6113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6114) );
  XNOR2_X1 U7796 ( .A(n6114), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6779) );
  AOI22_X1 U7797 ( .A1(n6066), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6360), .B2(
        n6779), .ZN(n6115) );
  NAND2_X1 U7798 ( .A1(n6116), .A2(n6115), .ZN(n7271) );
  OR2_X1 U7799 ( .A1(n9767), .A2(n6304), .ZN(n6124) );
  NAND2_X1 U7800 ( .A1(n4521), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7801 ( .A1(n8868), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6121) );
  OAI21_X1 U7802 ( .B1(n6117), .B2(P1_REG3_REG_5__SCAN_IN), .A(n6134), .ZN(
        n6118) );
  INV_X1 U7803 ( .A(n6118), .ZN(n7272) );
  NAND2_X1 U7804 ( .A1(n6073), .A2(n7272), .ZN(n6120) );
  NAND2_X1 U7805 ( .A1(n6025), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6119) );
  AND4_X2 U7806 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n7172)
         );
  OR2_X1 U7807 ( .A1(n4518), .A2(n7172), .ZN(n6123) );
  AND2_X1 U7808 ( .A1(n6124), .A2(n6123), .ZN(n7046) );
  NAND2_X1 U7809 ( .A1(n6502), .A2(n7271), .ZN(n6127) );
  NAND2_X1 U7810 ( .A1(n6127), .A2(n6126), .ZN(n6128) );
  XNOR2_X1 U7811 ( .A(n6128), .B(n6081), .ZN(n7044) );
  OR2_X1 U7812 ( .A1(n6614), .A2(n6154), .ZN(n6132) );
  NAND2_X1 U7813 ( .A1(n6129), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6130) );
  XNOR2_X1 U7814 ( .A(n6130), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6778) );
  AOI22_X1 U7815 ( .A1(n6066), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6360), .B2(
        n6778), .ZN(n6131) );
  NAND2_X1 U7816 ( .A1(n6132), .A2(n6131), .ZN(n9772) );
  NAND2_X1 U7817 ( .A1(n6502), .A2(n9772), .ZN(n6141) );
  NAND2_X1 U7818 ( .A1(n4521), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7819 ( .A1(n8868), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6138) );
  AND2_X1 U7820 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  NOR2_X1 U7821 ( .A1(n6159), .A2(n6135), .ZN(n7169) );
  NAND2_X1 U7822 ( .A1(n6073), .A2(n7169), .ZN(n6137) );
  NAND2_X1 U7823 ( .A1(n4517), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6136) );
  OR2_X1 U7824 ( .A1(n6304), .A2(n7279), .ZN(n6140) );
  NAND2_X1 U7825 ( .A1(n6141), .A2(n6140), .ZN(n6142) );
  XNOR2_X1 U7826 ( .A(n6142), .B(n6081), .ZN(n7166) );
  NAND2_X1 U7827 ( .A1(n6419), .A2(n9772), .ZN(n6144) );
  OR2_X1 U7828 ( .A1(n4518), .A2(n7279), .ZN(n6143) );
  AND2_X1 U7829 ( .A1(n6144), .A2(n6143), .ZN(n7165) );
  AOI22_X1 U7830 ( .A1(n7046), .A2(n7044), .B1(n7166), .B2(n7165), .ZN(n6145)
         );
  NAND2_X1 U7831 ( .A1(n7043), .A2(n6145), .ZN(n6153) );
  INV_X1 U7832 ( .A(n7166), .ZN(n6151) );
  INV_X1 U7833 ( .A(n7044), .ZN(n7164) );
  INV_X1 U7834 ( .A(n7046), .ZN(n6146) );
  NAND2_X1 U7835 ( .A1(n7164), .A2(n6146), .ZN(n6147) );
  NAND2_X1 U7836 ( .A1(n6147), .A2(n7165), .ZN(n6150) );
  INV_X1 U7837 ( .A(n6147), .ZN(n6149) );
  INV_X1 U7838 ( .A(n7165), .ZN(n6148) );
  AOI22_X1 U7839 ( .A1(n6151), .A2(n6150), .B1(n6149), .B2(n6148), .ZN(n6152)
         );
  NAND2_X1 U7840 ( .A1(n6156), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6157) );
  XNOR2_X1 U7841 ( .A(n6157), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6777) );
  AOI22_X1 U7842 ( .A1(n6066), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6360), .B2(
        n6777), .ZN(n6158) );
  NAND2_X1 U7843 ( .A1(n9779), .A2(n6502), .ZN(n6166) );
  NAND2_X1 U7844 ( .A1(n4521), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7845 ( .A1(n8868), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6163) );
  OR2_X1 U7846 ( .A1(n6159), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6160) );
  AND2_X1 U7847 ( .A1(n6177), .A2(n6160), .ZN(n7289) );
  NAND2_X1 U7848 ( .A1(n6073), .A2(n7289), .ZN(n6162) );
  NAND2_X1 U7849 ( .A1(n4517), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6161) );
  OR2_X1 U7850 ( .A1(n6304), .A2(n7371), .ZN(n6165) );
  NAND2_X1 U7851 ( .A1(n6166), .A2(n6165), .ZN(n6167) );
  XNOR2_X1 U7852 ( .A(n6167), .B(n6081), .ZN(n6169) );
  AOI22_X1 U7853 ( .A1(n9779), .A2(n6419), .B1(n6449), .B2(n9710), .ZN(n6168)
         );
  NAND2_X1 U7854 ( .A1(n6169), .A2(n6168), .ZN(n6172) );
  OR2_X1 U7855 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  NAND2_X1 U7856 ( .A1(n6172), .A2(n6170), .ZN(n7109) );
  INV_X1 U7857 ( .A(n7109), .ZN(n6171) );
  NAND2_X1 U7858 ( .A1(n6633), .A2(n8841), .ZN(n6175) );
  INV_X1 U7859 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7860 ( .A1(n5039), .A2(n6173), .ZN(n6213) );
  NAND2_X1 U7861 ( .A1(n6213), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6190) );
  XNOR2_X1 U7862 ( .A(n6190), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6776) );
  AOI22_X1 U7863 ( .A1(n6066), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6360), .B2(
        n6776), .ZN(n6174) );
  NAND2_X1 U7864 ( .A1(n6175), .A2(n6174), .ZN(n9720) );
  NAND2_X1 U7865 ( .A1(n9720), .A2(n6502), .ZN(n6184) );
  NAND2_X1 U7866 ( .A1(n4521), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7867 ( .A1(n8868), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7868 ( .A1(n6177), .A2(n6176), .ZN(n6178) );
  AND2_X1 U7869 ( .A1(n6195), .A2(n6178), .ZN(n9717) );
  NAND2_X1 U7870 ( .A1(n6073), .A2(n9717), .ZN(n6180) );
  NAND2_X1 U7871 ( .A1(n4517), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6179) );
  OR2_X1 U7872 ( .A1(n6450), .A2(n7361), .ZN(n6183) );
  NAND2_X1 U7873 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  XNOR2_X1 U7874 ( .A(n6185), .B(n4512), .ZN(n6187) );
  XNOR2_X1 U7875 ( .A(n6189), .B(n6187), .ZN(n7367) );
  NOR2_X1 U7876 ( .A1(n4518), .A2(n7361), .ZN(n6186) );
  AOI21_X1 U7877 ( .B1(n9720), .B2(n6419), .A(n6186), .ZN(n7368) );
  INV_X1 U7878 ( .A(n6187), .ZN(n6188) );
  NAND2_X1 U7879 ( .A1(n6189), .A2(n6188), .ZN(n7356) );
  NAND2_X1 U7880 ( .A1(n6638), .A2(n8841), .ZN(n6194) );
  NAND2_X1 U7881 ( .A1(n6190), .A2(n6211), .ZN(n6191) );
  NAND2_X1 U7882 ( .A1(n6191), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6192) );
  XNOR2_X1 U7883 ( .A(n6192), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6896) );
  AOI22_X1 U7884 ( .A1(n6066), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6360), .B2(
        n6896), .ZN(n6193) );
  NAND2_X1 U7885 ( .A1(n6194), .A2(n6193), .ZN(n7363) );
  NAND2_X1 U7886 ( .A1(n7363), .A2(n6502), .ZN(n6202) );
  NAND2_X1 U7887 ( .A1(n8868), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7888 ( .A1(n4517), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6199) );
  AND2_X1 U7889 ( .A1(n6195), .A2(n6791), .ZN(n6196) );
  NOR2_X1 U7890 ( .A1(n6223), .A2(n6196), .ZN(n7357) );
  NAND2_X1 U7891 ( .A1(n6073), .A2(n7357), .ZN(n6198) );
  NAND2_X1 U7892 ( .A1(n4521), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6197) );
  OR2_X1 U7893 ( .A1(n6304), .A2(n7524), .ZN(n6201) );
  NAND2_X1 U7894 ( .A1(n6202), .A2(n6201), .ZN(n6203) );
  XNOR2_X1 U7895 ( .A(n6203), .B(n4512), .ZN(n6206) );
  NOR2_X1 U7896 ( .A1(n4518), .A2(n7524), .ZN(n6204) );
  AOI21_X1 U7897 ( .B1(n7363), .B2(n6419), .A(n6204), .ZN(n6207) );
  XNOR2_X1 U7898 ( .A(n6206), .B(n6207), .ZN(n7355) );
  AND2_X1 U7899 ( .A1(n7356), .A2(n7355), .ZN(n6205) );
  INV_X1 U7900 ( .A(n6206), .ZN(n6208) );
  OR2_X1 U7901 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  NAND2_X1 U7902 ( .A1(n6641), .A2(n8841), .ZN(n6222) );
  INV_X1 U7903 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7904 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  NOR2_X1 U7905 ( .A1(n6213), .A2(n6212), .ZN(n6218) );
  INV_X1 U7906 ( .A(n6218), .ZN(n6214) );
  NAND2_X1 U7907 ( .A1(n6214), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6215) );
  MUX2_X1 U7908 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6215), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n6216) );
  INV_X1 U7909 ( .A(n6216), .ZN(n6220) );
  INV_X1 U7910 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7911 ( .A1(n6218), .A2(n6217), .ZN(n6256) );
  INV_X1 U7912 ( .A(n6256), .ZN(n6219) );
  AOI22_X1 U7913 ( .A1(n6066), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6360), .B2(
        n6941), .ZN(n6221) );
  NAND2_X1 U7914 ( .A1(n6222), .A2(n6221), .ZN(n7526) );
  NAND2_X1 U7915 ( .A1(n7526), .A2(n6502), .ZN(n6230) );
  NAND2_X1 U7916 ( .A1(n4521), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7917 ( .A1(n8868), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6227) );
  NOR2_X1 U7918 ( .A1(n6223), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6224) );
  OR2_X1 U7919 ( .A1(n6237), .A2(n6224), .ZN(n7140) );
  INV_X1 U7920 ( .A(n7140), .ZN(n7520) );
  NAND2_X1 U7921 ( .A1(n6073), .A2(n7520), .ZN(n6226) );
  NAND2_X1 U7922 ( .A1(n4517), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6225) );
  OR2_X1 U7923 ( .A1(n6083), .A2(n7300), .ZN(n6229) );
  NAND2_X1 U7924 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  XNOR2_X1 U7925 ( .A(n6231), .B(n6081), .ZN(n7514) );
  NOR2_X1 U7926 ( .A1(n4518), .A2(n7300), .ZN(n6232) );
  AOI21_X1 U7927 ( .B1(n7526), .B2(n6419), .A(n6232), .ZN(n7518) );
  NAND2_X1 U7928 ( .A1(n7514), .A2(n7518), .ZN(n6233) );
  NAND2_X1 U7929 ( .A1(n6656), .A2(n8841), .ZN(n6236) );
  NAND2_X1 U7930 ( .A1(n6256), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6234) );
  XNOR2_X1 U7931 ( .A(n6234), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6987) );
  AOI22_X1 U7932 ( .A1(n6066), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6360), .B2(
        n6987), .ZN(n6235) );
  NAND2_X1 U7933 ( .A1(n7569), .A2(n6502), .ZN(n6244) );
  NAND2_X1 U7934 ( .A1(n8868), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U7935 ( .A1(n4521), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6241) );
  OR2_X1 U7936 ( .A1(n6237), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6238) );
  AND2_X1 U7937 ( .A1(n6261), .A2(n6238), .ZN(n7568) );
  NAND2_X1 U7938 ( .A1(n6073), .A2(n7568), .ZN(n6240) );
  NAND2_X1 U7939 ( .A1(n4517), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6239) );
  OR2_X1 U7940 ( .A1(n6450), .A2(n7380), .ZN(n6243) );
  NAND2_X1 U7941 ( .A1(n6244), .A2(n6243), .ZN(n6245) );
  XNOR2_X1 U7942 ( .A(n6245), .B(n4512), .ZN(n6251) );
  NAND2_X1 U7943 ( .A1(n7569), .A2(n6419), .ZN(n6247) );
  OR2_X1 U7944 ( .A1(n4518), .A2(n7380), .ZN(n6246) );
  NAND2_X1 U7945 ( .A1(n6247), .A2(n6246), .ZN(n6252) );
  NAND2_X1 U7946 ( .A1(n6251), .A2(n6252), .ZN(n7562) );
  OAI21_X1 U7947 ( .B1(n7514), .B2(n7518), .A(n7562), .ZN(n6248) );
  INV_X1 U7948 ( .A(n6248), .ZN(n6249) );
  INV_X1 U7949 ( .A(n6251), .ZN(n6254) );
  INV_X1 U7950 ( .A(n6252), .ZN(n6253) );
  NAND2_X1 U7951 ( .A1(n6714), .A2(n8841), .ZN(n6259) );
  NAND2_X1 U7952 ( .A1(n6275), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6257) );
  XNOR2_X1 U7953 ( .A(n6257), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7222) );
  AOI22_X1 U7954 ( .A1(n6066), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6360), .B2(
        n7222), .ZN(n6258) );
  NAND2_X1 U7955 ( .A1(n9031), .A2(n6502), .ZN(n6268) );
  NAND2_X1 U7956 ( .A1(n8868), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7957 ( .A1(n4521), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7958 ( .A1(n6261), .A2(n6260), .ZN(n6262) );
  AND2_X1 U7959 ( .A1(n6280), .A2(n6262), .ZN(n7493) );
  NAND2_X1 U7960 ( .A1(n6073), .A2(n7493), .ZN(n6264) );
  NAND2_X1 U7961 ( .A1(n4517), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6263) );
  OR2_X1 U7962 ( .A1(n6304), .A2(n9027), .ZN(n6267) );
  NAND2_X1 U7963 ( .A1(n6268), .A2(n6267), .ZN(n6269) );
  XNOR2_X1 U7964 ( .A(n6269), .B(n4512), .ZN(n6271) );
  NOR2_X1 U7965 ( .A1(n4518), .A2(n9027), .ZN(n6270) );
  AOI21_X1 U7966 ( .B1(n9031), .B2(n6419), .A(n6270), .ZN(n6272) );
  XNOR2_X1 U7967 ( .A(n6271), .B(n6272), .ZN(n7488) );
  INV_X1 U7968 ( .A(n6271), .ZN(n6273) );
  NAND2_X1 U7969 ( .A1(n6273), .A2(n6272), .ZN(n6274) );
  NAND2_X1 U7970 ( .A1(n6733), .A2(n8841), .ZN(n6278) );
  OAI21_X1 U7971 ( .B1(n6275), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6276) );
  XNOR2_X1 U7972 ( .A(n6276), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9260) );
  AOI22_X1 U7973 ( .A1(n6066), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6360), .B2(
        n9260), .ZN(n6277) );
  NAND2_X1 U7974 ( .A1(n6278), .A2(n6277), .ZN(n7470) );
  NAND2_X1 U7975 ( .A1(n7470), .A2(n6502), .ZN(n6287) );
  NAND2_X1 U7976 ( .A1(n4521), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7977 ( .A1(n8868), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U7978 ( .A1(n6280), .A2(n6279), .ZN(n6281) );
  AND2_X1 U7979 ( .A1(n6298), .A2(n6281), .ZN(n7580) );
  NAND2_X1 U7980 ( .A1(n6073), .A2(n7580), .ZN(n6283) );
  NAND2_X1 U7981 ( .A1(n4517), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6282) );
  OR2_X1 U7982 ( .A1(n6304), .A2(n9692), .ZN(n6286) );
  NAND2_X1 U7983 ( .A1(n6287), .A2(n6286), .ZN(n6288) );
  XNOR2_X1 U7984 ( .A(n6288), .B(n4512), .ZN(n6290) );
  NOR2_X1 U7985 ( .A1(n4518), .A2(n9692), .ZN(n6289) );
  AOI21_X1 U7986 ( .B1(n7470), .B2(n6419), .A(n6289), .ZN(n6291) );
  XNOR2_X1 U7987 ( .A(n6290), .B(n6291), .ZN(n7574) );
  INV_X1 U7988 ( .A(n6290), .ZN(n6292) );
  NAND2_X1 U7989 ( .A1(n6823), .A2(n8841), .ZN(n6296) );
  OR2_X1 U7990 ( .A1(n6293), .A2(n9626), .ZN(n6294) );
  XNOR2_X1 U7991 ( .A(n6294), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9268) );
  AOI22_X1 U7992 ( .A1(n6066), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6360), .B2(
        n9268), .ZN(n6295) );
  AND2_X1 U7993 ( .A1(n6298), .A2(n6297), .ZN(n6299) );
  NOR2_X1 U7994 ( .A1(n6319), .A2(n6299), .ZN(n9697) );
  NAND2_X1 U7995 ( .A1(n9697), .A2(n6073), .ZN(n6303) );
  NAND2_X1 U7996 ( .A1(n4521), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U7997 ( .A1(n8868), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7998 ( .A1(n4517), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6300) );
  NOR2_X1 U7999 ( .A1(n6304), .A2(n7577), .ZN(n6305) );
  AOI21_X1 U8000 ( .B1(n9699), .B2(n6502), .A(n6305), .ZN(n6306) );
  XNOR2_X1 U8001 ( .A(n6306), .B(n4512), .ZN(n6310) );
  NAND2_X1 U8002 ( .A1(n9699), .A2(n6419), .ZN(n6308) );
  OR2_X1 U8003 ( .A1(n4518), .A2(n7577), .ZN(n6307) );
  NAND2_X1 U8004 ( .A1(n6308), .A2(n6307), .ZN(n7704) );
  INV_X1 U8005 ( .A(n6310), .ZN(n6311) );
  NAND2_X1 U8006 ( .A1(n6847), .A2(n8841), .ZN(n6316) );
  NAND2_X1 U8007 ( .A1(n6313), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6314) );
  XNOR2_X1 U8008 ( .A(n6314), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9281) );
  AOI22_X1 U8009 ( .A1(n6066), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6360), .B2(
        n9281), .ZN(n6315) );
  NAND2_X1 U8010 ( .A1(n7609), .A2(n6502), .ZN(n6325) );
  NAND2_X1 U8011 ( .A1(n4520), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U8012 ( .A1(n4517), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6317) );
  AND2_X1 U8013 ( .A1(n6318), .A2(n6317), .ZN(n6323) );
  OR2_X1 U8014 ( .A1(n6319), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6320) );
  AND2_X1 U8015 ( .A1(n6320), .A2(n6334), .ZN(n7760) );
  NAND2_X1 U8016 ( .A1(n7760), .A2(n6073), .ZN(n6322) );
  NAND2_X1 U8017 ( .A1(n4521), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6321) );
  OR2_X1 U8018 ( .A1(n6304), .A2(n9694), .ZN(n6324) );
  NAND2_X1 U8019 ( .A1(n6325), .A2(n6324), .ZN(n6326) );
  XNOR2_X1 U8020 ( .A(n6326), .B(n4512), .ZN(n6328) );
  NOR2_X1 U8021 ( .A1(n4518), .A2(n9694), .ZN(n6327) );
  AOI21_X1 U8022 ( .B1(n7609), .B2(n6419), .A(n6327), .ZN(n7752) );
  NAND2_X1 U8023 ( .A1(n6329), .A2(n6328), .ZN(n7751) );
  NAND2_X2 U8024 ( .A1(n7756), .A2(n7751), .ZN(n8764) );
  NAND2_X1 U8025 ( .A1(n6907), .A2(n8841), .ZN(n6332) );
  NAND2_X1 U8026 ( .A1(n4602), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6330) );
  XNOR2_X1 U8027 ( .A(n6330), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9311) );
  AOI22_X1 U8028 ( .A1(n6066), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6360), .B2(
        n9311), .ZN(n6331) );
  NAND2_X1 U8029 ( .A1(n6334), .A2(n6333), .ZN(n6335) );
  NAND2_X1 U8030 ( .A1(n6346), .A2(n6335), .ZN(n8765) );
  AOI22_X1 U8031 ( .A1(n4521), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n4517), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U8032 ( .A1(n4520), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6337) );
  OAI211_X1 U8033 ( .C1(n8765), .C2(n6370), .A(n6338), .B(n6337), .ZN(n9140)
         );
  AOI22_X1 U8034 ( .A1(n8769), .A2(n6502), .B1(n6419), .B2(n9140), .ZN(n6339)
         );
  XNOR2_X1 U8035 ( .A(n6339), .B(n4512), .ZN(n6341) );
  AOI22_X1 U8036 ( .A1(n8769), .A2(n6419), .B1(n6449), .B2(n9140), .ZN(n6340)
         );
  XNOR2_X1 U8037 ( .A(n6341), .B(n6340), .ZN(n8763) );
  NAND2_X1 U8038 ( .A1(n6966), .A2(n8841), .ZN(n6344) );
  XNOR2_X1 U8039 ( .A(n6342), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9330) );
  AOI22_X1 U8040 ( .A1(n6066), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6360), .B2(
        n9330), .ZN(n6343) );
  NAND2_X1 U8041 ( .A1(n8778), .A2(n6502), .ZN(n6351) );
  AND2_X1 U8042 ( .A1(n6346), .A2(n6345), .ZN(n6347) );
  OR2_X1 U8043 ( .A1(n6347), .A2(n6363), .ZN(n8774) );
  AOI22_X1 U8044 ( .A1(n4521), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8868), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U8045 ( .A1(n4517), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6348) );
  OAI211_X1 U8046 ( .C1(n8774), .C2(n6370), .A(n6349), .B(n6348), .ZN(n9139)
         );
  NAND2_X1 U8047 ( .A1(n9139), .A2(n6419), .ZN(n6350) );
  NAND2_X1 U8048 ( .A1(n6351), .A2(n6350), .ZN(n6352) );
  XNOR2_X1 U8049 ( .A(n6352), .B(n4512), .ZN(n6353) );
  AOI22_X1 U8050 ( .A1(n8778), .A2(n6419), .B1(n6449), .B2(n9139), .ZN(n6354)
         );
  XNOR2_X1 U8051 ( .A(n6353), .B(n6354), .ZN(n8773) );
  INV_X1 U8052 ( .A(n6353), .ZN(n6355) );
  NAND2_X1 U8053 ( .A1(n7016), .A2(n8841), .ZN(n6362) );
  OR2_X1 U8054 ( .A1(n6357), .A2(n6356), .ZN(n6358) );
  AND2_X1 U8055 ( .A1(n6359), .A2(n6358), .ZN(n9347) );
  AOI22_X1 U8056 ( .A1(n6066), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6360), .B2(
        n9347), .ZN(n6361) );
  NOR2_X1 U8057 ( .A1(n6363), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6364) );
  OR2_X1 U8058 ( .A1(n6365), .A2(n6364), .ZN(n8816) );
  INV_X1 U8059 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9324) );
  NAND2_X1 U8060 ( .A1(n4517), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6367) );
  NAND2_X1 U8061 ( .A1(n8868), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6366) );
  OAI211_X1 U8062 ( .C1(n6074), .C2(n9324), .A(n6367), .B(n6366), .ZN(n6368)
         );
  INV_X1 U8063 ( .A(n6368), .ZN(n6369) );
  AOI22_X1 U8064 ( .A1(n9608), .A2(n6046), .B1(n6419), .B2(n9138), .ZN(n6371)
         );
  XOR2_X1 U8065 ( .A(n4512), .B(n6371), .Z(n6372) );
  AOI22_X1 U8066 ( .A1(n9608), .A2(n6419), .B1(n6449), .B2(n9138), .ZN(n8814)
         );
  XOR2_X1 U8067 ( .A(n6375), .B(n6373), .Z(n8740) );
  NAND2_X1 U8068 ( .A1(n7294), .A2(n8841), .ZN(n6377) );
  NAND2_X1 U8069 ( .A1(n6066), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6376) );
  NOR2_X1 U8070 ( .A1(n6378), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6379) );
  NOR2_X1 U8071 ( .A1(n6391), .A2(n6379), .ZN(n9512) );
  INV_X1 U8072 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6382) );
  NAND2_X1 U8073 ( .A1(n4517), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6381) );
  NAND2_X1 U8074 ( .A1(n4520), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6380) );
  OAI211_X1 U8075 ( .C1(n6074), .C2(n6382), .A(n6381), .B(n6380), .ZN(n6383)
         );
  AOI21_X1 U8076 ( .B1(n9512), .B2(n6073), .A(n6383), .ZN(n9532) );
  OAI22_X1 U8077 ( .A1(n9515), .A2(n4891), .B1(n9532), .B2(n6304), .ZN(n6384)
         );
  XNOR2_X1 U8078 ( .A(n6384), .B(n4512), .ZN(n8793) );
  OAI22_X1 U8079 ( .A1(n9515), .A2(n6083), .B1(n9532), .B2(n4518), .ZN(n6386)
         );
  NAND2_X1 U8080 ( .A1(n8795), .A2(n6385), .ZN(n6388) );
  INV_X1 U8081 ( .A(n6386), .ZN(n8792) );
  NAND2_X1 U8082 ( .A1(n8793), .A2(n6386), .ZN(n6387) );
  NAND2_X1 U8083 ( .A1(n6388), .A2(n6387), .ZN(n8746) );
  NAND2_X1 U8084 ( .A1(n7376), .A2(n8841), .ZN(n6390) );
  NAND2_X1 U8085 ( .A1(n6066), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U8086 ( .A1(n9593), .A2(n6502), .ZN(n6400) );
  OR2_X1 U8087 ( .A1(n6391), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6392) );
  AND2_X1 U8088 ( .A1(n6392), .A2(n6411), .ZN(n9497) );
  NAND2_X1 U8089 ( .A1(n9497), .A2(n6073), .ZN(n6398) );
  INV_X1 U8090 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U8091 ( .A1(n4517), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6394) );
  NAND2_X1 U8092 ( .A1(n8868), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6393) );
  OAI211_X1 U8093 ( .C1(n6074), .C2(n6395), .A(n6394), .B(n6393), .ZN(n6396)
         );
  INV_X1 U8094 ( .A(n6396), .ZN(n6397) );
  NAND2_X1 U8095 ( .A1(n6398), .A2(n6397), .ZN(n9471) );
  NAND2_X1 U8096 ( .A1(n9471), .A2(n6419), .ZN(n6399) );
  NAND2_X1 U8097 ( .A1(n6400), .A2(n6399), .ZN(n6401) );
  XNOR2_X1 U8098 ( .A(n6401), .B(n4512), .ZN(n6404) );
  AOI22_X1 U8099 ( .A1(n9593), .A2(n6419), .B1(n6449), .B2(n9471), .ZN(n6402)
         );
  XNOR2_X1 U8100 ( .A(n6404), .B(n6402), .ZN(n8747) );
  INV_X1 U8101 ( .A(n6402), .ZN(n6403) );
  AOI21_X2 U8102 ( .B1(n8746), .B2(n8747), .A(n6405), .ZN(n8806) );
  INV_X1 U8103 ( .A(n8806), .ZN(n6407) );
  AOI22_X1 U8104 ( .A1(n9584), .A2(n6419), .B1(n6449), .B2(n9462), .ZN(n8803)
         );
  AOI21_X1 U8105 ( .B1(n8806), .B2(n8804), .A(n8803), .ZN(n6406) );
  NAND2_X1 U8106 ( .A1(n7511), .A2(n8841), .ZN(n6410) );
  NAND2_X1 U8107 ( .A1(n6066), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U8108 ( .A1(n4521), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6418) );
  NAND2_X1 U8109 ( .A1(n4520), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6417) );
  NOR2_X1 U8110 ( .A1(n6413), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6414) );
  NOR2_X1 U8111 ( .A1(n6426), .A2(n6414), .ZN(n9455) );
  NAND2_X1 U8112 ( .A1(n6073), .A2(n9455), .ZN(n6416) );
  NAND2_X1 U8113 ( .A1(n4517), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6415) );
  NAND4_X1 U8114 ( .A1(n6418), .A2(n6417), .A3(n6416), .A4(n6415), .ZN(n9470)
         );
  AOI22_X1 U8115 ( .A1(n9580), .A2(n6502), .B1(n6419), .B2(n9470), .ZN(n6420)
         );
  XOR2_X1 U8116 ( .A(n4512), .B(n6420), .Z(n6422) );
  OAI22_X1 U8117 ( .A1(n9457), .A2(n6083), .B1(n8809), .B2(n4518), .ZN(n6421)
         );
  NOR2_X1 U8118 ( .A1(n6422), .A2(n6421), .ZN(n6423) );
  AOI21_X1 U8119 ( .B1(n6422), .B2(n6421), .A(n6423), .ZN(n8731) );
  INV_X1 U8120 ( .A(n6423), .ZN(n8782) );
  NAND2_X1 U8121 ( .A1(n7583), .A2(n8841), .ZN(n6425) );
  NAND2_X1 U8122 ( .A1(n6066), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U8123 ( .A1(n9575), .A2(n6502), .ZN(n6433) );
  NAND2_X1 U8124 ( .A1(n4521), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U8125 ( .A1(n4520), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6430) );
  NOR2_X1 U8126 ( .A1(n6426), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6427) );
  NOR2_X1 U8127 ( .A1(n6443), .A2(n6427), .ZN(n9443) );
  NAND2_X1 U8128 ( .A1(n6073), .A2(n9443), .ZN(n6429) );
  NAND2_X1 U8129 ( .A1(n4517), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6428) );
  OR2_X1 U8130 ( .A1(n6083), .A2(n8757), .ZN(n6432) );
  NAND2_X1 U8131 ( .A1(n6433), .A2(n6432), .ZN(n6434) );
  XNOR2_X1 U8132 ( .A(n6434), .B(n6081), .ZN(n6437) );
  NOR2_X1 U8133 ( .A1(n4518), .A2(n8757), .ZN(n6435) );
  AOI21_X1 U8134 ( .B1(n9575), .B2(n6419), .A(n6435), .ZN(n6436) );
  NAND2_X1 U8135 ( .A1(n6437), .A2(n6436), .ZN(n6439) );
  OR2_X1 U8136 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  NAND2_X1 U8137 ( .A1(n6439), .A2(n6438), .ZN(n8781) );
  INV_X1 U8138 ( .A(n6439), .ZN(n6440) );
  NAND2_X1 U8139 ( .A1(n7684), .A2(n8841), .ZN(n6442) );
  NAND2_X1 U8140 ( .A1(n6066), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U8141 ( .A1(n4521), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6448) );
  NAND2_X1 U8142 ( .A1(n8868), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8143 ( .A1(n6443), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6457) );
  OAI21_X1 U8144 ( .B1(n6443), .B2(P1_REG3_REG_25__SCAN_IN), .A(n6457), .ZN(
        n6444) );
  INV_X1 U8145 ( .A(n6444), .ZN(n9428) );
  NAND2_X1 U8146 ( .A1(n6073), .A2(n9428), .ZN(n6446) );
  NAND2_X1 U8147 ( .A1(n4517), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6445) );
  AOI22_X1 U8148 ( .A1(n9570), .A2(n6419), .B1(n6449), .B2(n9449), .ZN(n6468)
         );
  NAND2_X1 U8149 ( .A1(n9570), .A2(n6502), .ZN(n6452) );
  OR2_X1 U8150 ( .A1(n6450), .A2(n8787), .ZN(n6451) );
  NAND2_X1 U8151 ( .A1(n6452), .A2(n6451), .ZN(n6453) );
  XNOR2_X1 U8152 ( .A(n6453), .B(n4512), .ZN(n6470) );
  XOR2_X1 U8153 ( .A(n6468), .B(n6470), .Z(n8753) );
  NOR2_X2 U8154 ( .A1(n8754), .A2(n8753), .ZN(n8828) );
  NAND2_X1 U8155 ( .A1(n7698), .A2(n8841), .ZN(n6455) );
  NAND2_X1 U8156 ( .A1(n6066), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U8157 ( .A1(n4521), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U8158 ( .A1(n4520), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6462) );
  INV_X1 U8159 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U8160 ( .A1(n6456), .A2(n6457), .ZN(n6459) );
  INV_X1 U8161 ( .A(n6457), .ZN(n6458) );
  NAND2_X1 U8162 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n6458), .ZN(n6493) );
  AND2_X1 U8163 ( .A1(n6459), .A2(n6493), .ZN(n9415) );
  NAND2_X1 U8164 ( .A1(n6073), .A2(n9415), .ZN(n6461) );
  NAND2_X1 U8165 ( .A1(n4517), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6460) );
  NOR2_X1 U8166 ( .A1(n4518), .A2(n8756), .ZN(n6464) );
  AOI21_X1 U8167 ( .B1(n9565), .B2(n6419), .A(n6464), .ZN(n6472) );
  NAND2_X1 U8168 ( .A1(n9565), .A2(n6046), .ZN(n6466) );
  OR2_X1 U8169 ( .A1(n6304), .A2(n8756), .ZN(n6465) );
  NAND2_X1 U8170 ( .A1(n6466), .A2(n6465), .ZN(n6467) );
  XNOR2_X1 U8171 ( .A(n6467), .B(n4512), .ZN(n6474) );
  XOR2_X1 U8172 ( .A(n6472), .B(n6474), .Z(n8826) );
  INV_X1 U8173 ( .A(n6468), .ZN(n6469) );
  NOR2_X1 U8174 ( .A1(n6470), .A2(n6469), .ZN(n8827) );
  INV_X1 U8175 ( .A(n6472), .ZN(n6473) );
  NAND2_X1 U8176 ( .A1(n7731), .A2(n8841), .ZN(n6476) );
  NAND2_X1 U8177 ( .A1(n6066), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U8178 ( .A1(n9560), .A2(n6502), .ZN(n6482) );
  NAND2_X1 U8179 ( .A1(n4521), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U8180 ( .A1(n8868), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6479) );
  XNOR2_X1 U8181 ( .A(n6493), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9404) );
  NAND2_X1 U8182 ( .A1(n4523), .A2(n9404), .ZN(n6478) );
  NAND2_X1 U8183 ( .A1(n4517), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6477) );
  OR2_X1 U8184 ( .A1(n6083), .A2(n8835), .ZN(n6481) );
  NAND2_X1 U8185 ( .A1(n6482), .A2(n6481), .ZN(n6483) );
  XNOR2_X1 U8186 ( .A(n6483), .B(n6081), .ZN(n6486) );
  NOR2_X1 U8187 ( .A1(n4518), .A2(n8835), .ZN(n6484) );
  AOI21_X1 U8188 ( .B1(n9560), .B2(n6419), .A(n6484), .ZN(n6485) );
  NAND2_X1 U8189 ( .A1(n6486), .A2(n6485), .ZN(n6549) );
  OAI21_X1 U8190 ( .B1(n6486), .B2(n6485), .A(n6549), .ZN(n6592) );
  NAND2_X1 U8191 ( .A1(n7791), .A2(n8841), .ZN(n6488) );
  NAND2_X1 U8192 ( .A1(n6066), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U8193 ( .A1(n9554), .A2(n6419), .ZN(n6500) );
  NAND2_X1 U8194 ( .A1(n4521), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6498) );
  NAND2_X1 U8195 ( .A1(n4520), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6497) );
  INV_X1 U8196 ( .A(n6493), .ZN(n6490) );
  AND2_X1 U8197 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6489) );
  NAND2_X1 U8198 ( .A1(n6490), .A2(n6489), .ZN(n6542) );
  INV_X1 U8199 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6492) );
  INV_X1 U8200 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6491) );
  OAI21_X1 U8201 ( .B1(n6493), .B2(n6492), .A(n6491), .ZN(n6494) );
  NAND2_X1 U8202 ( .A1(n6073), .A2(n7773), .ZN(n6496) );
  NAND2_X1 U8203 ( .A1(n4517), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6495) );
  OR2_X1 U8204 ( .A1(n4518), .A2(n9379), .ZN(n6499) );
  NAND2_X1 U8205 ( .A1(n6500), .A2(n6499), .ZN(n6501) );
  XNOR2_X1 U8206 ( .A(n6501), .B(n6081), .ZN(n6505) );
  NAND2_X1 U8207 ( .A1(n9554), .A2(n6502), .ZN(n6503) );
  OAI21_X1 U8208 ( .B1(n9379), .B2(n6083), .A(n6503), .ZN(n6504) );
  XNOR2_X1 U8209 ( .A(n6505), .B(n6504), .ZN(n6528) );
  INV_X1 U8210 ( .A(n6528), .ZN(n6550) );
  NAND2_X1 U8211 ( .A1(n6506), .A2(P1_B_REG_SCAN_IN), .ZN(n6508) );
  INV_X1 U8212 ( .A(n7596), .ZN(n6507) );
  MUX2_X1 U8213 ( .A(n6508), .B(P1_B_REG_SCAN_IN), .S(n6507), .Z(n6510) );
  NAND2_X1 U8214 ( .A1(n6510), .A2(n6509), .ZN(n6644) );
  INV_X1 U8215 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10424) );
  INV_X1 U8216 ( .A(n6509), .ZN(n7712) );
  INV_X1 U8217 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10399) );
  AND2_X1 U8218 ( .A1(n6506), .A2(n7712), .ZN(n6646) );
  NOR4_X1 U8219 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6519) );
  NOR4_X1 U8220 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6518) );
  INV_X1 U8221 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10247) );
  INV_X1 U8222 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9734) );
  INV_X1 U8223 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9733) );
  INV_X1 U8224 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9732) );
  NAND4_X1 U8225 ( .A1(n10247), .A2(n9734), .A3(n9733), .A4(n9732), .ZN(n6516)
         );
  NOR4_X1 U8226 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6514) );
  NOR4_X1 U8227 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6513) );
  NOR4_X1 U8228 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6512) );
  NOR4_X1 U8229 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6511) );
  NAND4_X1 U8230 ( .A1(n6514), .A2(n6513), .A3(n6512), .A4(n6511), .ZN(n6515)
         );
  NOR4_X1 U8231 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6516), .A4(n6515), .ZN(n6517) );
  NAND3_X1 U8232 ( .A1(n6519), .A2(n6518), .A3(n6517), .ZN(n6520) );
  NAND2_X1 U8233 ( .A1(n6521), .A2(n6520), .ZN(n6720) );
  NAND3_X1 U8234 ( .A1(n9543), .A2(n7055), .A3(n6720), .ZN(n6541) );
  NAND2_X1 U8235 ( .A1(n6522), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6524) );
  OR2_X1 U8236 ( .A1(n6541), .A2(n6533), .ZN(n6530) );
  NAND2_X1 U8237 ( .A1(n6525), .A2(n8881), .ZN(n7072) );
  INV_X1 U8238 ( .A(n6526), .ZN(n8955) );
  NAND2_X1 U8239 ( .A1(n9828), .A2(n7068), .ZN(n6527) );
  NAND3_X1 U8240 ( .A1(n6550), .A2(n8830), .A3(n6549), .ZN(n6555) );
  NAND2_X1 U8241 ( .A1(n6593), .A2(n6529), .ZN(n6554) );
  INV_X1 U8242 ( .A(n6530), .ZN(n6532) );
  OR2_X1 U8243 ( .A1(n7072), .A2(n8914), .ZN(n7071) );
  INV_X1 U8244 ( .A(n7071), .ZN(n6531) );
  INV_X1 U8245 ( .A(n6541), .ZN(n6535) );
  OR2_X1 U8246 ( .A1(n7068), .A2(n6526), .ZN(n6722) );
  OR2_X1 U8247 ( .A1(n6533), .A2(n6722), .ZN(n6539) );
  NOR2_X1 U8248 ( .A1(n6539), .A2(n7793), .ZN(n6534) );
  INV_X1 U8249 ( .A(n6717), .ZN(n6536) );
  NAND2_X1 U8250 ( .A1(n6541), .A2(n6536), .ZN(n6538) );
  OR2_X1 U8251 ( .A1(n7068), .A2(n8955), .ZN(n6718) );
  AND3_X1 U8252 ( .A1(n6019), .A2(n7509), .A3(n6718), .ZN(n6537) );
  NAND2_X1 U8253 ( .A1(n6538), .A2(n6537), .ZN(n6828) );
  NAND2_X1 U8254 ( .A1(n8837), .A2(n7773), .ZN(n6548) );
  INV_X1 U8255 ( .A(n6539), .ZN(n9127) );
  NAND2_X1 U8256 ( .A1(n9127), .A2(n7793), .ZN(n6540) );
  NAND2_X1 U8257 ( .A1(n4521), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8258 ( .A1(n4520), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6545) );
  INV_X1 U8259 ( .A(n6542), .ZN(n9388) );
  NAND2_X1 U8260 ( .A1(n6073), .A2(n9388), .ZN(n6544) );
  NAND2_X1 U8261 ( .A1(n4517), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6543) );
  NAND4_X1 U8262 ( .A1(n6546), .A2(n6545), .A3(n6544), .A4(n6543), .ZN(n9135)
         );
  AOI22_X1 U8263 ( .A1(n8796), .A2(n9135), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6547) );
  OAI211_X1 U8264 ( .C1(n8835), .C2(n8798), .A(n6548), .B(n6547), .ZN(n6552)
         );
  NOR3_X1 U8265 ( .A1(n6550), .A2(n8823), .A3(n6549), .ZN(n6551) );
  AOI211_X1 U8266 ( .C1(n9554), .C2(n8821), .A(n6552), .B(n6551), .ZN(n6553)
         );
  OAI211_X1 U8267 ( .C1(n6593), .C2(n6555), .A(n6554), .B(n6553), .ZN(P1_U3220) );
  NAND2_X1 U8268 ( .A1(n8007), .A2(n8101), .ZN(n6556) );
  NAND2_X1 U8269 ( .A1(n6559), .A2(n6558), .ZN(n6563) );
  INV_X1 U8270 ( .A(n6560), .ZN(n6561) );
  NAND2_X1 U8271 ( .A1(n6561), .A2(n10485), .ZN(n6562) );
  NAND2_X1 U8272 ( .A1(n6563), .A2(n6562), .ZN(n7783) );
  INV_X1 U8273 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8040) );
  INV_X1 U8274 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10410) );
  MUX2_X1 U8275 ( .A(n8040), .B(n10410), .S(n6600), .Z(n7782) );
  XNOR2_X1 U8276 ( .A(n7785), .B(SI_29_), .ZN(n8864) );
  NAND2_X1 U8277 ( .A1(n8864), .A2(n5535), .ZN(n6565) );
  OR2_X1 U8278 ( .A1(n7803), .A2(n8040), .ZN(n6564) );
  NAND2_X1 U8279 ( .A1(n6565), .A2(n6564), .ZN(n6584) );
  NAND2_X1 U8280 ( .A1(n6584), .A2(n8142), .ZN(n7816) );
  XNOR2_X1 U8281 ( .A(n6566), .B(n8005), .ZN(n6580) );
  XNOR2_X1 U8282 ( .A(n7806), .B(n4704), .ZN(n6581) );
  INV_X1 U8283 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6573) );
  NAND2_X1 U8284 ( .A1(n6568), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U8285 ( .A1(n6569), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6570) );
  OAI211_X1 U8286 ( .C1(n6573), .C2(n6572), .A(n6571), .B(n6570), .ZN(n6574)
         );
  INV_X1 U8287 ( .A(n6574), .ZN(n6575) );
  NAND2_X1 U8288 ( .A1(n7814), .A2(n6575), .ZN(n8279) );
  NAND2_X1 U8289 ( .A1(n6576), .A2(P2_B_REG_SCAN_IN), .ZN(n6577) );
  AND2_X1 U8290 ( .A1(n9983), .A2(n6577), .ZN(n8399) );
  AOI22_X1 U8291 ( .A1(n8410), .A2(n9986), .B1(n8279), .B2(n8399), .ZN(n6578)
         );
  OAI21_X1 U8292 ( .B1(n6581), .B2(n7502), .A(n6578), .ZN(n6579) );
  INV_X1 U8293 ( .A(n6581), .ZN(n6583) );
  NAND2_X1 U8294 ( .A1(n6587), .A2(n10048), .ZN(n6586) );
  INV_X1 U8295 ( .A(n6584), .ZN(n8035) );
  NAND2_X1 U8296 ( .A1(n6586), .A2(n5093), .ZN(P2_U3456) );
  INV_X1 U8297 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6588) );
  NOR2_X1 U8298 ( .A1(n10064), .A2(n6588), .ZN(n6589) );
  AOI22_X1 U8299 ( .A1(n8832), .A2(n9434), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6594) );
  OAI21_X1 U8300 ( .B1(n9379), .B2(n8834), .A(n6594), .ZN(n6595) );
  AOI21_X1 U8301 ( .B1(n9404), .B2(n8837), .A(n6595), .ZN(n6597) );
  INV_X1 U8302 ( .A(n9560), .ZN(n9407) );
  NAND2_X1 U8303 ( .A1(n9560), .A2(n8821), .ZN(n6596) );
  INV_X1 U8304 ( .A(n6019), .ZN(n6599) );
  AND2_X1 U8305 ( .A1(n6600), .A2(P1_U3086), .ZN(n7508) );
  INV_X2 U8306 ( .A(n7508), .ZN(n9634) );
  AND2_X1 U8307 ( .A1(n7798), .A2(P1_U3086), .ZN(n9629) );
  AOI22_X1 U8308 ( .A1(n9629), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9158), .ZN(n6601) );
  OAI21_X1 U8309 ( .B1(n6606), .B2(n9634), .A(n6601), .ZN(P1_U3354) );
  INV_X1 U8310 ( .A(n9179), .ZN(n6782) );
  INV_X1 U8311 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6602) );
  INV_X2 U8312 ( .A(n9629), .ZN(n9632) );
  OAI222_X1 U8313 ( .A1(n6782), .A2(P1_U3086), .B1(n9634), .B2(n6612), .C1(
        n6602), .C2(n9632), .ZN(P1_U3353) );
  INV_X1 U8314 ( .A(n9193), .ZN(n6784) );
  OAI222_X1 U8315 ( .A1(n6784), .A2(P1_U3086), .B1(n9634), .B2(n6617), .C1(
        n6603), .C2(n9632), .ZN(P1_U3352) );
  INV_X1 U8316 ( .A(n9676), .ZN(n6785) );
  INV_X1 U8317 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6604) );
  OAI222_X1 U8318 ( .A1(n6785), .A2(P1_U3086), .B1(n9634), .B2(n6620), .C1(
        n6604), .C2(n9632), .ZN(P1_U3351) );
  NAND2_X1 U8319 ( .A1(n4506), .A2(P2_U3151), .ZN(n8039) );
  AND2_X1 U8320 ( .A1(n7798), .A2(P2_U3151), .ZN(n7733) );
  INV_X2 U8321 ( .A(n7733), .ZN(n8729) );
  OAI222_X1 U8322 ( .A1(n8039), .A2(n6607), .B1(n8729), .B2(n6606), .C1(
        P2_U3151), .C2(n6678), .ZN(P2_U3294) );
  INV_X1 U8323 ( .A(n6778), .ZN(n9211) );
  INV_X1 U8324 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6608) );
  OAI222_X1 U8325 ( .A1(n9211), .A2(P1_U3086), .B1(n9634), .B2(n6614), .C1(
        n6608), .C2(n9632), .ZN(P1_U3349) );
  INV_X1 U8326 ( .A(n6779), .ZN(n9198) );
  OAI222_X1 U8327 ( .A1(n9198), .A2(P1_U3086), .B1(n9634), .B2(n6610), .C1(
        n4638), .C2(n9632), .ZN(P1_U3350) );
  INV_X1 U8328 ( .A(n8039), .ZN(n6734) );
  INV_X1 U8329 ( .A(n6734), .ZN(n8723) );
  OAI222_X1 U8330 ( .A1(n8723), .A2(n6611), .B1(n8729), .B2(n6610), .C1(
        P2_U3151), .C2(n6609), .ZN(P2_U3290) );
  OAI222_X1 U8331 ( .A1(n8723), .A2(n6613), .B1(n8729), .B2(n6612), .C1(
        P2_U3151), .C2(n4513), .ZN(P2_U3293) );
  OAI222_X1 U8332 ( .A1(n8723), .A2(n6615), .B1(n8729), .B2(n6614), .C1(
        P2_U3151), .C2(n9912), .ZN(P2_U3289) );
  OAI222_X1 U8333 ( .A1(n8723), .A2(n6618), .B1(n8729), .B2(n6617), .C1(
        P2_U3151), .C2(n6616), .ZN(P2_U3292) );
  OAI222_X1 U8334 ( .A1(n8723), .A2(n6621), .B1(n8729), .B2(n6620), .C1(
        P2_U3151), .C2(n6619), .ZN(P2_U3291) );
  INV_X1 U8335 ( .A(n6777), .ZN(n9224) );
  INV_X1 U8336 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6622) );
  OAI222_X1 U8337 ( .A1(n9224), .A2(P1_U3086), .B1(n9634), .B2(n6623), .C1(
        n6622), .C2(n9632), .ZN(P1_U3348) );
  OAI222_X1 U8338 ( .A1(n8723), .A2(n6624), .B1(n8729), .B2(n6623), .C1(
        P2_U3151), .C2(n9930), .ZN(P2_U3288) );
  INV_X1 U8339 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6628) );
  INV_X1 U8340 ( .A(n6626), .ZN(n6627) );
  AOI22_X1 U8341 ( .A1(n6637), .A2(n6628), .B1(n6631), .B2(n6627), .ZN(
        P2_U3376) );
  INV_X1 U8342 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6632) );
  INV_X1 U8343 ( .A(n6629), .ZN(n6630) );
  AOI22_X1 U8344 ( .A1(n6637), .A2(n6632), .B1(n6631), .B2(n6630), .ZN(
        P2_U3377) );
  INV_X1 U8345 ( .A(n6776), .ZN(n9237) );
  INV_X1 U8346 ( .A(n6633), .ZN(n6635) );
  OAI222_X1 U8347 ( .A1(n9237), .A2(P1_U3086), .B1(n9634), .B2(n6635), .C1(
        n6634), .C2(n9632), .ZN(P1_U3347) );
  OAI222_X1 U8348 ( .A1(n8723), .A2(n6636), .B1(n8729), .B2(n6635), .C1(
        P2_U3151), .C2(n9956), .ZN(P2_U3287) );
  AND2_X1 U8349 ( .A1(n6637), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8350 ( .A1(n6637), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8351 ( .A1(n6637), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8352 ( .A1(n6637), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8353 ( .A1(n6637), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8354 ( .A1(n6637), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8355 ( .A1(n6637), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8356 ( .A1(n6637), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8357 ( .A1(n6637), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8358 ( .A1(n6637), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8359 ( .A1(n6637), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8360 ( .A1(n6637), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8361 ( .A1(n6637), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8362 ( .A1(n6637), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8363 ( .A1(n6637), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8364 ( .A1(n6637), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8365 ( .A1(n6637), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8366 ( .A1(n6637), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8367 ( .A1(n6637), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8368 ( .A1(n6637), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8369 ( .A1(n6637), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8370 ( .A1(n6637), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8371 ( .A1(n6637), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8372 ( .A1(n6637), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8373 ( .A1(n6637), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8374 ( .A1(n6637), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8375 ( .A1(n6637), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8376 ( .A1(n6637), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8377 ( .A1(n6637), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8378 ( .A1(n6637), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8379 ( .A(n6638), .ZN(n6640) );
  OAI222_X1 U8380 ( .A1(n8729), .A2(n6640), .B1(n7196), .B2(P2_U3151), .C1(
        n6639), .C2(n8723), .ZN(P2_U3286) );
  INV_X1 U8381 ( .A(n6896), .ZN(n6794) );
  OAI222_X1 U8382 ( .A1(P1_U3086), .A2(n6794), .B1(n9634), .B2(n6640), .C1(
        n10237), .C2(n9632), .ZN(P1_U3346) );
  INV_X1 U8383 ( .A(n6641), .ZN(n6643) );
  OAI222_X1 U8384 ( .A1(n8729), .A2(n6643), .B1(n7343), .B2(P2_U3151), .C1(
        n6642), .C2(n8723), .ZN(P2_U3285) );
  INV_X1 U8385 ( .A(n6941), .ZN(n6906) );
  OAI222_X1 U8386 ( .A1(P1_U3086), .A2(n6906), .B1(n9634), .B2(n6643), .C1(
        n10483), .C2(n9632), .ZN(P1_U3345) );
  OR2_X1 U8387 ( .A1(n9735), .A2(n10399), .ZN(n6645) );
  OAI21_X1 U8388 ( .B1(n9731), .B2(n6646), .A(n6645), .ZN(P1_U3440) );
  MUX2_X1 U8389 ( .A(n6659), .B(n7629), .S(P2_U3893), .Z(n6647) );
  INV_X1 U8390 ( .A(n6647), .ZN(P2_U3502) );
  INV_X1 U8391 ( .A(n7509), .ZN(n6648) );
  OR2_X1 U8392 ( .A1(n6019), .A2(n6648), .ZN(n6649) );
  NAND2_X1 U8393 ( .A1(n6649), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6763) );
  INV_X1 U8394 ( .A(n7068), .ZN(n8912) );
  NAND2_X1 U8395 ( .A1(n7509), .A2(n8912), .ZN(n6651) );
  NAND2_X1 U8396 ( .A1(n6651), .A2(n6650), .ZN(n6762) );
  INV_X1 U8397 ( .A(n6762), .ZN(n6652) );
  OR2_X1 U8398 ( .A1(n6763), .A2(n6652), .ZN(n9338) );
  NOR2_X1 U8399 ( .A1(n9675), .A2(P1_U3973), .ZN(P1_U3085) );
  MUX2_X1 U8400 ( .A(n10237), .B(n7616), .S(P2_U3893), .Z(n6653) );
  INV_X1 U8401 ( .A(n6653), .ZN(P2_U3500) );
  NAND2_X1 U8402 ( .A1(n9731), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6654) );
  OAI21_X1 U8403 ( .B1(n9731), .B2(n6655), .A(n6654), .ZN(P1_U3439) );
  INV_X1 U8404 ( .A(n6656), .ZN(n6660) );
  OAI222_X1 U8405 ( .A1(n8723), .A2(n6658), .B1(n8729), .B2(n6660), .C1(
        P2_U3151), .C2(n6657), .ZN(P2_U3284) );
  INV_X1 U8406 ( .A(n6987), .ZN(n6981) );
  OAI222_X1 U8407 ( .A1(n6981), .A2(P1_U3086), .B1(n9634), .B2(n6660), .C1(
        n6659), .C2(n9632), .ZN(P1_U3344) );
  INV_X1 U8408 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6676) );
  NOR2_X1 U8409 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10223), .ZN(n6933) );
  INV_X1 U8410 ( .A(n6661), .ZN(n6663) );
  INV_X1 U8411 ( .A(n6662), .ZN(n6704) );
  AOI21_X1 U8412 ( .B1(n5404), .B2(n6663), .A(n6704), .ZN(n6668) );
  INV_X1 U8413 ( .A(n6664), .ZN(n6666) );
  INV_X1 U8414 ( .A(n6665), .ZN(n6698) );
  AOI21_X1 U8415 ( .B1(n5403), .B2(n6666), .A(n6698), .ZN(n6667) );
  OAI22_X1 U8416 ( .A1(n6668), .A2(n9953), .B1(n9948), .B2(n6667), .ZN(n6669)
         );
  AOI211_X1 U8417 ( .C1(n6670), .C2(n9915), .A(n6933), .B(n6669), .ZN(n6675)
         );
  OAI21_X1 U8418 ( .B1(n6672), .B2(n6671), .A(n6691), .ZN(n6673) );
  NAND2_X1 U8419 ( .A1(n6673), .A2(n9964), .ZN(n6674) );
  OAI211_X1 U8420 ( .C1(n6676), .C2(n9969), .A(n6675), .B(n6674), .ZN(P2_U3185) );
  XNOR2_X1 U8421 ( .A(n6677), .B(n9866), .ZN(n6689) );
  OAI22_X1 U8422 ( .A1(n9957), .A2(n6678), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6879), .ZN(n6687) );
  AOI21_X1 U8423 ( .B1(n10050), .B2(n6680), .A(n6679), .ZN(n6685) );
  AOI21_X1 U8424 ( .B1(n6683), .B2(n6682), .A(n6681), .ZN(n6684) );
  OAI22_X1 U8425 ( .A1(n6685), .A2(n9953), .B1(n9948), .B2(n6684), .ZN(n6686)
         );
  AOI211_X1 U8426 ( .C1(n9933), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6687), .B(
        n6686), .ZN(n6688) );
  OAI21_X1 U8427 ( .B1(n7442), .B2(n6689), .A(n6688), .ZN(P2_U3183) );
  INV_X1 U8428 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6713) );
  AND2_X1 U8429 ( .A1(n6691), .A2(n6690), .ZN(n6694) );
  OAI211_X1 U8430 ( .C1(n6694), .C2(n6693), .A(n9964), .B(n6692), .ZN(n6712)
         );
  NOR2_X1 U8431 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10269), .ZN(n6958) );
  INV_X1 U8432 ( .A(n6695), .ZN(n6696) );
  NOR3_X1 U8433 ( .A1(n6698), .A2(n6697), .A3(n6696), .ZN(n6699) );
  NOR2_X1 U8434 ( .A1(n6700), .A2(n6699), .ZN(n6708) );
  INV_X1 U8435 ( .A(n6701), .ZN(n6702) );
  NOR3_X1 U8436 ( .A1(n6704), .A2(n6703), .A3(n6702), .ZN(n6705) );
  INV_X1 U8437 ( .A(n9953), .ZN(n7435) );
  OAI21_X1 U8438 ( .B1(n6706), .B2(n6705), .A(n7435), .ZN(n6707) );
  OAI21_X1 U8439 ( .B1(n6708), .B2(n9948), .A(n6707), .ZN(n6709) );
  AOI211_X1 U8440 ( .C1(n6710), .C2(n9915), .A(n6958), .B(n6709), .ZN(n6711)
         );
  OAI211_X1 U8441 ( .C1(n6713), .C2(n9969), .A(n6712), .B(n6711), .ZN(P2_U3186) );
  INV_X1 U8442 ( .A(n6714), .ZN(n6732) );
  OAI222_X1 U8443 ( .A1(n8729), .A2(n6732), .B1(n6716), .B2(P2_U3151), .C1(
        n6715), .C2(n8039), .ZN(P2_U3283) );
  OR2_X1 U8444 ( .A1(n7055), .A2(n6717), .ZN(n6721) );
  NAND3_X1 U8445 ( .A1(n6720), .A2(n6719), .A3(n6718), .ZN(n7054) );
  INV_X1 U8446 ( .A(n9543), .ZN(n7056) );
  INV_X1 U8447 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6731) );
  INV_X1 U8448 ( .A(n7233), .ZN(n7186) );
  NAND2_X1 U8449 ( .A1(n6722), .A2(n7072), .ZN(n7237) );
  INV_X1 U8450 ( .A(n7237), .ZN(n6725) );
  NAND2_X1 U8451 ( .A1(n6723), .A2(n6526), .ZN(n6724) );
  NAND2_X1 U8452 ( .A1(n6725), .A2(n6724), .ZN(n7311) );
  OR2_X1 U8453 ( .A1(n6726), .A2(n6525), .ZN(n6727) );
  NAND2_X1 U8454 ( .A1(n8919), .A2(n4510), .ZN(n9118) );
  NAND2_X2 U8455 ( .A1(n6727), .A2(n9118), .ZN(n9491) );
  OR2_X1 U8456 ( .A1(n7233), .A2(n7178), .ZN(n8920) );
  NAND2_X1 U8457 ( .A1(n7178), .A2(n7233), .ZN(n7060) );
  AND2_X1 U8458 ( .A1(n8920), .A2(n7060), .ZN(n8883) );
  INV_X1 U8459 ( .A(n8883), .ZN(n6728) );
  OAI21_X1 U8460 ( .B1(n9824), .B2(n9491), .A(n6728), .ZN(n6729) );
  INV_X1 U8461 ( .A(n4509), .ZN(n9152) );
  INV_X1 U8462 ( .A(n7793), .ZN(n9173) );
  NAND2_X1 U8463 ( .A1(n9152), .A2(n9708), .ZN(n7236) );
  OAI211_X1 U8464 ( .C1(n7072), .C2(n7186), .A(n6729), .B(n7236), .ZN(n9611)
         );
  NAND2_X1 U8465 ( .A1(n9836), .A2(n9611), .ZN(n6730) );
  OAI21_X1 U8466 ( .B1(n9836), .B2(n6731), .A(n6730), .ZN(P1_U3453) );
  INV_X1 U8467 ( .A(n7222), .ZN(n6982) );
  OAI222_X1 U8468 ( .A1(P1_U3086), .A2(n6982), .B1(n9634), .B2(n6732), .C1(
        n10225), .C2(n9632), .ZN(P1_U3343) );
  INV_X1 U8469 ( .A(n6733), .ZN(n6795) );
  AOI22_X1 U8470 ( .A1(n8305), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n6734), .ZN(n6735) );
  OAI21_X1 U8471 ( .B1(n6795), .B2(n8729), .A(n6735), .ZN(P2_U3282) );
  INV_X1 U8472 ( .A(n6736), .ZN(n6839) );
  AND2_X1 U8473 ( .A1(n6755), .A2(n6839), .ZN(n6817) );
  INV_X1 U8474 ( .A(n6817), .ZN(n6737) );
  INV_X1 U8475 ( .A(n6738), .ZN(n6743) );
  INV_X1 U8476 ( .A(n6739), .ZN(n6754) );
  INV_X1 U8477 ( .A(n6740), .ZN(n6741) );
  AOI21_X1 U8478 ( .B1(n6748), .B2(n6754), .A(n6741), .ZN(n6742) );
  OAI21_X1 U8479 ( .B1(n6744), .B2(n6743), .A(n6742), .ZN(n6745) );
  NAND2_X1 U8480 ( .A1(n6745), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6750) );
  NAND2_X1 U8481 ( .A1(n6839), .A2(n6746), .ZN(n8026) );
  INV_X1 U8482 ( .A(n8026), .ZN(n6747) );
  NAND2_X1 U8483 ( .A1(n6748), .A2(n6747), .ZN(n6749) );
  NAND2_X1 U8484 ( .A1(n6750), .A2(n6749), .ZN(n6932) );
  NOR2_X1 U8485 ( .A1(n6932), .A2(n6751), .ZN(n6869) );
  INV_X1 U8486 ( .A(n6869), .ZN(n6752) );
  NAND2_X1 U8487 ( .A1(n6752), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6761) );
  OR2_X1 U8488 ( .A1(n6758), .A2(n6753), .ZN(n6757) );
  NAND2_X1 U8489 ( .A1(n6755), .A2(n6754), .ZN(n6756) );
  NAND2_X1 U8490 ( .A1(n8293), .A2(n6846), .ZN(n7853) );
  NAND2_X1 U8491 ( .A1(n7857), .A2(n7853), .ZN(n7826) );
  OR2_X1 U8492 ( .A1(n6758), .A2(n10042), .ZN(n6759) );
  AOI22_X1 U8493 ( .A1(n8244), .A2(n7826), .B1(n6808), .B2(n8236), .ZN(n6760)
         );
  OAI211_X1 U8494 ( .C1(n4879), .C2(n8271), .A(n6761), .B(n6760), .ZN(P2_U3172) );
  INV_X1 U8495 ( .A(n9666), .ZN(n6774) );
  NOR2_X1 U8496 ( .A1(n7793), .A2(n4522), .ZN(n9176) );
  INV_X1 U8497 ( .A(n9672), .ZN(n9327) );
  NOR2_X1 U8498 ( .A1(n6896), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6765) );
  AOI21_X1 U8499 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6896), .A(n6765), .ZN(
        n6773) );
  INV_X1 U8500 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6767) );
  NAND2_X1 U8501 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9174) );
  NOR2_X1 U8502 ( .A1(n9154), .A2(n9174), .ZN(n9153) );
  AOI21_X1 U8503 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n9158), .A(n9153), .ZN(
        n9167) );
  MUX2_X1 U8504 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6048), .S(n9179), .Z(n6766)
         );
  INV_X1 U8505 ( .A(n6766), .ZN(n9166) );
  NOR2_X1 U8506 ( .A1(n9167), .A2(n9166), .ZN(n9165) );
  MUX2_X1 U8507 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6767), .S(n9193), .Z(n9185)
         );
  INV_X1 U8508 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6768) );
  MUX2_X1 U8509 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6768), .S(n9676), .Z(n9668)
         );
  INV_X1 U8510 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6769) );
  AOI22_X1 U8511 ( .A1(n6779), .A2(n6769), .B1(P1_REG2_REG_5__SCAN_IN), .B2(
        n9198), .ZN(n9202) );
  AOI21_X1 U8512 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6779), .A(n9201), .ZN(
        n9216) );
  INV_X1 U8513 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7157) );
  AOI22_X1 U8514 ( .A1(n6778), .A2(n7157), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n9211), .ZN(n9215) );
  NOR2_X1 U8515 ( .A1(n9216), .A2(n9215), .ZN(n9214) );
  INV_X1 U8516 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6770) );
  AOI22_X1 U8517 ( .A1(n6777), .A2(n6770), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9224), .ZN(n9228) );
  INV_X1 U8518 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6771) );
  AOI22_X1 U8519 ( .A1(n6776), .A2(n6771), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n9237), .ZN(n9241) );
  NAND2_X1 U8520 ( .A1(n6773), .A2(n6772), .ZN(n6892) );
  OAI21_X1 U8521 ( .B1(n6773), .B2(n6772), .A(n6892), .ZN(n6790) );
  NAND2_X1 U8522 ( .A1(n6774), .A2(n4522), .ZN(n9351) );
  INV_X1 U8523 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6775) );
  MUX2_X1 U8524 ( .A(n6775), .B(P1_REG1_REG_9__SCAN_IN), .S(n6896), .Z(n6787)
         );
  INV_X1 U8525 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9850) );
  MUX2_X1 U8526 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n9850), .S(n6776), .Z(n9245)
         );
  INV_X1 U8527 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9848) );
  MUX2_X1 U8528 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9848), .S(n6777), .Z(n9232)
         );
  INV_X1 U8529 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9846) );
  MUX2_X1 U8530 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n9846), .S(n6778), .Z(n9219)
         );
  INV_X1 U8531 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9844) );
  MUX2_X1 U8532 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9844), .S(n6779), .Z(n9206)
         );
  INV_X1 U8533 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9842) );
  INV_X1 U8534 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9840) );
  INV_X1 U8535 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9838) );
  MUX2_X1 U8536 ( .A(n9838), .B(P1_REG1_REG_2__SCAN_IN), .S(n9179), .Z(n9168)
         );
  INV_X1 U8537 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6780) );
  MUX2_X1 U8538 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6780), .S(n9158), .Z(n9160)
         );
  AND2_X1 U8539 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9161) );
  NAND2_X1 U8540 ( .A1(n9160), .A2(n9161), .ZN(n9159) );
  NAND2_X1 U8541 ( .A1(n9158), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6781) );
  AND2_X1 U8542 ( .A1(n9159), .A2(n6781), .ZN(n9169) );
  NOR2_X1 U8543 ( .A1(n9168), .A2(n9169), .ZN(n9191) );
  NOR2_X1 U8544 ( .A1(n6782), .A2(n9838), .ZN(n9186) );
  MUX2_X1 U8545 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9840), .S(n9193), .Z(n6783)
         );
  OAI21_X1 U8546 ( .B1(n9191), .B2(n9186), .A(n6783), .ZN(n9189) );
  OAI21_X1 U8547 ( .B1(n9840), .B2(n6784), .A(n9189), .ZN(n9681) );
  MUX2_X1 U8548 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n9842), .S(n9676), .Z(n9680)
         );
  NAND2_X1 U8549 ( .A1(n9681), .A2(n9680), .ZN(n9678) );
  OAI21_X1 U8550 ( .B1(n9842), .B2(n6785), .A(n9678), .ZN(n9207) );
  NAND2_X1 U8551 ( .A1(n9206), .A2(n9207), .ZN(n9205) );
  OAI21_X1 U8552 ( .B1(n9198), .B2(n9844), .A(n9205), .ZN(n9220) );
  NAND2_X1 U8553 ( .A1(n9219), .A2(n9220), .ZN(n9218) );
  OAI21_X1 U8554 ( .B1(n9211), .B2(n9846), .A(n9218), .ZN(n9233) );
  NAND2_X1 U8555 ( .A1(n9232), .A2(n9233), .ZN(n9231) );
  OAI21_X1 U8556 ( .B1(n9224), .B2(n9848), .A(n9231), .ZN(n9246) );
  NAND2_X1 U8557 ( .A1(n9245), .A2(n9246), .ZN(n9244) );
  OAI21_X1 U8558 ( .B1(n9237), .B2(n9850), .A(n9244), .ZN(n6786) );
  NOR2_X1 U8559 ( .A1(n6787), .A2(n6786), .ZN(n6897) );
  AOI21_X1 U8560 ( .B1(n6787), .B2(n6786), .A(n6897), .ZN(n6788) );
  NOR2_X1 U8561 ( .A1(n9351), .A2(n6788), .ZN(n6789) );
  AOI21_X1 U8562 ( .B1(n9327), .B2(n6790), .A(n6789), .ZN(n6793) );
  NOR2_X1 U8563 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6791), .ZN(n7358) );
  AOI21_X1 U8564 ( .B1(n9675), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7358), .ZN(
        n6792) );
  OAI211_X1 U8565 ( .C1(n6794), .C2(n9354), .A(n6793), .B(n6792), .ZN(P1_U3252) );
  INV_X1 U8566 ( .A(n9260), .ZN(n9255) );
  INV_X1 U8567 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10277) );
  OAI222_X1 U8568 ( .A1(n9255), .A2(P1_U3086), .B1(n9634), .B2(n6795), .C1(
        n10277), .C2(n9632), .ZN(P1_U3342) );
  NAND2_X1 U8569 ( .A1(n8292), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6796) );
  OAI21_X1 U8570 ( .B1(n8493), .B2(n8292), .A(n6796), .ZN(P2_U3512) );
  NOR2_X1 U8571 ( .A1(n4879), .A2(n8565), .ZN(n6842) );
  INV_X1 U8572 ( .A(n6842), .ZN(n6798) );
  OAI21_X1 U8573 ( .B1(n9981), .B2(n10035), .A(n7826), .ZN(n6797) );
  OAI211_X1 U8574 ( .C1(n10042), .C2(n6846), .A(n6798), .B(n6797), .ZN(n6800)
         );
  NAND2_X1 U8575 ( .A1(n6800), .A2(n10048), .ZN(n6799) );
  OAI21_X1 U8576 ( .B1(n5376), .B2(n10048), .A(n6799), .ZN(P2_U3390) );
  NAND2_X1 U8577 ( .A1(n6800), .A2(n10064), .ZN(n6801) );
  OAI21_X1 U8578 ( .B1(n10064), .B2(n9865), .A(n6801), .ZN(P2_U3459) );
  NOR2_X1 U8579 ( .A1(n6802), .A2(n6805), .ZN(n6803) );
  AND2_X1 U8580 ( .A1(n6809), .A2(n7857), .ZN(n6815) );
  NAND2_X1 U8581 ( .A1(n6811), .A2(n4879), .ZN(n6861) );
  NAND2_X1 U8582 ( .A1(n6861), .A2(n6812), .ZN(n6814) );
  INV_X1 U8583 ( .A(n6862), .ZN(n6813) );
  AOI21_X1 U8584 ( .B1(n6815), .B2(n6814), .A(n6813), .ZN(n6822) );
  INV_X1 U8585 ( .A(n8293), .ZN(n6818) );
  OAI22_X1 U8586 ( .A1(n8256), .A2(n6818), .B1(n8276), .B2(n10002), .ZN(n6820)
         );
  NOR2_X1 U8587 ( .A1(n6869), .A2(n6879), .ZN(n6819) );
  AOI211_X1 U8588 ( .C1(n8258), .C2(n5398), .A(n6820), .B(n6819), .ZN(n6821)
         );
  OAI21_X1 U8589 ( .B1(n8264), .B2(n6822), .A(n6821), .ZN(P2_U3162) );
  INV_X1 U8590 ( .A(n9268), .ZN(n9272) );
  INV_X1 U8591 ( .A(n6823), .ZN(n6824) );
  INV_X1 U8592 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10430) );
  OAI222_X1 U8593 ( .A1(n9272), .A2(P1_U3086), .B1(n9634), .B2(n6824), .C1(
        n10430), .C2(n9632), .ZN(P1_U3341) );
  INV_X1 U8594 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6825) );
  OAI222_X1 U8595 ( .A1(n8723), .A2(n6825), .B1(n8729), .B2(n6824), .C1(
        P2_U3151), .C2(n8320), .ZN(P2_U3281) );
  XNOR2_X1 U8596 ( .A(n6827), .B(n6826), .ZN(n9172) );
  NOR2_X1 U8597 ( .A1(n6828), .A2(P1_U3086), .ZN(n6856) );
  INV_X1 U8598 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7235) );
  OAI22_X1 U8599 ( .A1(n6856), .A2(n7235), .B1(n4509), .B2(n8834), .ZN(n6829)
         );
  AOI21_X1 U8600 ( .B1(n7233), .B2(n8821), .A(n6829), .ZN(n6830) );
  OAI21_X1 U8601 ( .B1(n8823), .B2(n9172), .A(n6830), .ZN(P1_U3232) );
  NAND2_X1 U8602 ( .A1(n6831), .A2(n6832), .ZN(n6833) );
  XOR2_X1 U8603 ( .A(n6834), .B(n6833), .Z(n6838) );
  INV_X1 U8604 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9156) );
  INV_X1 U8605 ( .A(n7063), .ZN(n9151) );
  AOI22_X1 U8606 ( .A1(n8832), .A2(n6032), .B1(n8796), .B2(n9151), .ZN(n6835)
         );
  OAI21_X1 U8607 ( .B1(n6856), .B2(n9156), .A(n6835), .ZN(n6836) );
  AOI21_X1 U8608 ( .B1(n6016), .B2(n8821), .A(n6836), .ZN(n6837) );
  OAI21_X1 U8609 ( .B1(n6838), .B2(n8823), .A(n6837), .ZN(P1_U3222) );
  INV_X1 U8610 ( .A(n7826), .ZN(n6840) );
  NOR3_X1 U8611 ( .A1(n6840), .A2(n6839), .A3(n10040), .ZN(n6841) );
  AOI211_X1 U8612 ( .C1(n8554), .C2(P2_REG3_REG_0__SCAN_IN), .A(n6842), .B(
        n6841), .ZN(n6843) );
  MUX2_X1 U8613 ( .A(n6844), .B(n6843), .S(n9999), .Z(n6845) );
  OAI21_X1 U8614 ( .B1(n9975), .B2(n6846), .A(n6845), .ZN(P2_U3233) );
  INV_X1 U8615 ( .A(n6847), .ZN(n6849) );
  INV_X1 U8616 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6848) );
  OAI222_X1 U8617 ( .A1(n4712), .A2(P1_U3086), .B1(n9634), .B2(n6849), .C1(
        n6848), .C2(n9632), .ZN(P1_U3340) );
  INV_X1 U8618 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6850) );
  OAI222_X1 U8619 ( .A1(n8039), .A2(n6850), .B1(n8729), .B2(n6849), .C1(
        P2_U3151), .C2(n8341), .ZN(P2_U3280) );
  INV_X1 U8620 ( .A(n6853), .ZN(n6854) );
  AOI21_X1 U8621 ( .B1(n6851), .B2(n6852), .A(n6854), .ZN(n6859) );
  INV_X1 U8622 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7100) );
  INV_X1 U8623 ( .A(n7085), .ZN(n9150) );
  AOI22_X1 U8624 ( .A1(n8832), .A2(n9152), .B1(n8796), .B2(n9150), .ZN(n6855)
         );
  OAI21_X1 U8625 ( .B1(n6856), .B2(n7100), .A(n6855), .ZN(n6857) );
  AOI21_X1 U8626 ( .B1(n9745), .B2(n8821), .A(n6857), .ZN(n6858) );
  OAI21_X1 U8627 ( .B1(n6859), .B2(n8823), .A(n6858), .ZN(P1_U3237) );
  XNOR2_X1 U8628 ( .A(n4514), .B(n6860), .ZN(n6923) );
  XNOR2_X1 U8629 ( .A(n6923), .B(n5398), .ZN(n6864) );
  NAND2_X1 U8630 ( .A1(n6862), .A2(n6861), .ZN(n6863) );
  OAI21_X1 U8631 ( .B1(n6864), .B2(n6863), .A(n6925), .ZN(n6865) );
  NAND2_X1 U8632 ( .A1(n6865), .A2(n8244), .ZN(n6868) );
  OAI22_X1 U8633 ( .A1(n8256), .A2(n4879), .B1(n8276), .B2(n9989), .ZN(n6866)
         );
  AOI21_X1 U8634 ( .B1(n8258), .B2(n9984), .A(n6866), .ZN(n6867) );
  OAI211_X1 U8635 ( .C1(n6869), .C2(n10468), .A(n6868), .B(n6867), .ZN(
        P2_U3177) );
  OAI21_X1 U8636 ( .B1(n6874), .B2(n6871), .A(n6870), .ZN(n10005) );
  INV_X1 U8637 ( .A(n10005), .ZN(n6883) );
  NOR2_X1 U8638 ( .A1(n5088), .A2(n6872), .ZN(n8037) );
  INV_X1 U8639 ( .A(n8037), .ZN(n7507) );
  XNOR2_X1 U8640 ( .A(n6873), .B(n6874), .ZN(n6878) );
  INV_X1 U8641 ( .A(n7502), .ZN(n6875) );
  NAND2_X1 U8642 ( .A1(n10005), .A2(n6875), .ZN(n6877) );
  AOI22_X1 U8643 ( .A1(n9986), .A2(n8293), .B1(n5398), .B2(n9983), .ZN(n6876)
         );
  OAI211_X1 U8644 ( .C1(n6878), .C2(n8561), .A(n6877), .B(n6876), .ZN(n10003)
         );
  NAND2_X1 U8645 ( .A1(n10003), .A2(n9999), .ZN(n6882) );
  OAI22_X1 U8646 ( .A1(n9975), .A2(n10002), .B1(n9990), .B2(n6879), .ZN(n6880)
         );
  AOI21_X1 U8647 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n5088), .A(n6880), .ZN(
        n6881) );
  OAI211_X1 U8648 ( .C1(n6883), .C2(n7507), .A(n6882), .B(n6881), .ZN(P2_U3232) );
  XOR2_X1 U8649 ( .A(n6884), .B(n6885), .Z(n6891) );
  NAND2_X1 U8650 ( .A1(n8837), .A2(n6886), .ZN(n6888) );
  INV_X1 U8651 ( .A(n7127), .ZN(n9149) );
  NOR2_X1 U8652 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6886), .ZN(n9192) );
  AOI21_X1 U8653 ( .B1(n8796), .B2(n9149), .A(n9192), .ZN(n6887) );
  OAI211_X1 U8654 ( .C1(n8798), .C2(n7063), .A(n6888), .B(n6887), .ZN(n6889)
         );
  AOI21_X1 U8655 ( .B1(n7075), .B2(n8821), .A(n6889), .ZN(n6890) );
  OAI21_X1 U8656 ( .B1(n6891), .B2(n8823), .A(n6890), .ZN(P1_U3218) );
  OAI21_X1 U8657 ( .B1(n6896), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6892), .ZN(
        n6895) );
  INV_X1 U8658 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6893) );
  MUX2_X1 U8659 ( .A(n6893), .B(P1_REG2_REG_10__SCAN_IN), .S(n6941), .Z(n6894)
         );
  NOR2_X1 U8660 ( .A1(n6894), .A2(n6895), .ZN(n6940) );
  AOI211_X1 U8661 ( .C1(n6895), .C2(n6894), .A(n6940), .B(n9672), .ZN(n6903)
         );
  OR2_X1 U8662 ( .A1(n6896), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6899) );
  INV_X1 U8663 ( .A(n6897), .ZN(n6898) );
  NAND2_X1 U8664 ( .A1(n6899), .A2(n6898), .ZN(n6901) );
  INV_X1 U8665 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9853) );
  MUX2_X1 U8666 ( .A(n9853), .B(P1_REG1_REG_10__SCAN_IN), .S(n6941), .Z(n6900)
         );
  NOR2_X1 U8667 ( .A1(n6900), .A2(n6901), .ZN(n6939) );
  AOI211_X1 U8668 ( .C1(n6901), .C2(n6900), .A(n6939), .B(n9351), .ZN(n6902)
         );
  NOR2_X1 U8669 ( .A1(n6903), .A2(n6902), .ZN(n6905) );
  AND2_X1 U8670 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7521) );
  AOI21_X1 U8671 ( .B1(n9675), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7521), .ZN(
        n6904) );
  OAI211_X1 U8672 ( .C1(n6906), .C2(n9354), .A(n6905), .B(n6904), .ZN(P1_U3253) );
  INV_X1 U8673 ( .A(n6907), .ZN(n6910) );
  OAI222_X1 U8674 ( .A1(n8729), .A2(n6910), .B1(n8354), .B2(P2_U3151), .C1(
        n6908), .C2(n8723), .ZN(P2_U3279) );
  INV_X1 U8675 ( .A(n9311), .ZN(n9303) );
  OAI222_X1 U8676 ( .A1(P1_U3086), .A2(n9303), .B1(n9634), .B2(n6910), .C1(
        n6909), .C2(n9632), .ZN(P1_U3339) );
  XNOR2_X1 U8677 ( .A(n6911), .B(n7824), .ZN(n10015) );
  INV_X1 U8678 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6917) );
  OAI21_X1 U8679 ( .B1(n6913), .B2(n7824), .A(n6912), .ZN(n6916) );
  NAND2_X1 U8680 ( .A1(n9984), .A2(n9986), .ZN(n6914) );
  OAI21_X1 U8681 ( .B1(n7039), .B2(n8565), .A(n6914), .ZN(n6915) );
  AOI21_X1 U8682 ( .B1(n6916), .B2(n9981), .A(n6915), .ZN(n10019) );
  MUX2_X1 U8683 ( .A(n6917), .B(n10019), .S(n9999), .Z(n6920) );
  INV_X1 U8684 ( .A(n6962), .ZN(n6918) );
  AOI22_X1 U8685 ( .A1(n8555), .A2(n6959), .B1(n8554), .B2(n6918), .ZN(n6919)
         );
  OAI211_X1 U8686 ( .C1(n8558), .C2(n10015), .A(n6920), .B(n6919), .ZN(
        P2_U3229) );
  NAND2_X1 U8687 ( .A1(n8292), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6921) );
  OAI21_X1 U8688 ( .B1(n8446), .B2(n8292), .A(n6921), .ZN(P2_U3516) );
  XNOR2_X1 U8689 ( .A(n4511), .B(n10011), .ZN(n6950) );
  XNOR2_X1 U8690 ( .A(n6950), .B(n9984), .ZN(n6929) );
  INV_X1 U8691 ( .A(n5398), .ZN(n6922) );
  NAND2_X1 U8692 ( .A1(n6923), .A2(n6922), .ZN(n6924) );
  INV_X1 U8693 ( .A(n6952), .ZN(n6927) );
  AOI211_X1 U8694 ( .C1(n6929), .C2(n6928), .A(n8264), .B(n6927), .ZN(n6938)
         );
  OR2_X1 U8695 ( .A1(n6930), .A2(P2_U3151), .ZN(n8030) );
  INV_X1 U8696 ( .A(n8030), .ZN(n6931) );
  AOI21_X1 U8697 ( .B1(n8236), .B2(n6934), .A(n6933), .ZN(n6936) );
  AOI22_X1 U8698 ( .A1(n8258), .A2(n9971), .B1(n8269), .B2(n5398), .ZN(n6935)
         );
  OAI211_X1 U8699 ( .C1(n8247), .C2(P2_REG3_REG_3__SCAN_IN), .A(n6936), .B(
        n6935), .ZN(n6937) );
  OR2_X1 U8700 ( .A1(n6938), .A2(n6937), .ZN(P2_U3158) );
  INV_X1 U8701 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9855) );
  MUX2_X1 U8702 ( .A(n9855), .B(P1_REG1_REG_11__SCAN_IN), .S(n6987), .Z(n6978)
         );
  AOI21_X1 U8703 ( .B1(n6941), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6939), .ZN(
        n6979) );
  XOR2_X1 U8704 ( .A(n6978), .B(n6979), .Z(n6946) );
  NAND2_X1 U8705 ( .A1(n6987), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6942) );
  OAI21_X1 U8706 ( .B1(n6987), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6942), .ZN(
        n6943) );
  NOR2_X1 U8707 ( .A1(n6944), .A2(n6943), .ZN(n6986) );
  AOI211_X1 U8708 ( .C1(n6944), .C2(n6943), .A(n6986), .B(n9672), .ZN(n6945)
         );
  AOI21_X1 U8709 ( .B1(n9679), .B2(n6946), .A(n6945), .ZN(n6949) );
  NAND2_X1 U8710 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n7565) );
  INV_X1 U8711 ( .A(n7565), .ZN(n6947) );
  AOI21_X1 U8712 ( .B1(n9675), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n6947), .ZN(
        n6948) );
  OAI211_X1 U8713 ( .C1(n6981), .C2(n9354), .A(n6949), .B(n6948), .ZN(P1_U3254) );
  NAND2_X1 U8714 ( .A1(n6950), .A2(n9984), .ZN(n6951) );
  XNOR2_X1 U8715 ( .A(n4514), .B(n6959), .ZN(n6953) );
  INV_X1 U8716 ( .A(n9971), .ZN(n6972) );
  NAND2_X1 U8717 ( .A1(n6953), .A2(n6972), .ZN(n6998) );
  INV_X1 U8718 ( .A(n6953), .ZN(n6954) );
  NAND2_X1 U8719 ( .A1(n6954), .A2(n9971), .ZN(n6955) );
  AND2_X1 U8720 ( .A1(n6998), .A2(n6955), .ZN(n6956) );
  OAI21_X1 U8721 ( .B1(n6957), .B2(n6956), .A(n6995), .ZN(n6964) );
  AOI21_X1 U8722 ( .B1(n8236), .B2(n6959), .A(n6958), .ZN(n6961) );
  AOI22_X1 U8723 ( .A1(n8258), .A2(n8291), .B1(n8269), .B2(n9984), .ZN(n6960)
         );
  OAI211_X1 U8724 ( .C1(n8247), .C2(n6962), .A(n6961), .B(n6960), .ZN(n6963)
         );
  AOI21_X1 U8725 ( .B1(n6964), .B2(n8244), .A(n6963), .ZN(n6965) );
  INV_X1 U8726 ( .A(n6965), .ZN(P2_U3170) );
  INV_X1 U8727 ( .A(n6966), .ZN(n6969) );
  OAI222_X1 U8728 ( .A1(n8039), .A2(n6968), .B1(n8729), .B2(n6969), .C1(
        P2_U3151), .C2(n6967), .ZN(P2_U3278) );
  INV_X1 U8729 ( .A(n9330), .ZN(n9309) );
  OAI222_X1 U8730 ( .A1(n9632), .A2(n10403), .B1(n9634), .B2(n6969), .C1(n9309), .C2(P1_U3086), .ZN(P1_U3338) );
  XNOR2_X1 U8731 ( .A(n7039), .B(n7023), .ZN(n7827) );
  XNOR2_X1 U8732 ( .A(n6970), .B(n7827), .ZN(n6971) );
  OAI222_X1 U8733 ( .A1(n8565), .A2(n7331), .B1(n8563), .B2(n6972), .C1(n6971), 
        .C2(n8561), .ZN(n7018) );
  INV_X1 U8734 ( .A(n7018), .ZN(n6977) );
  XNOR2_X1 U8735 ( .A(n6973), .B(n7827), .ZN(n7019) );
  NOR2_X1 U8736 ( .A1(n9975), .A2(n7023), .ZN(n6975) );
  OAI22_X1 U8737 ( .A1(n9999), .A2(n9890), .B1(n7003), .B2(n9990), .ZN(n6974)
         );
  AOI211_X1 U8738 ( .C1(n7019), .C2(n9977), .A(n6975), .B(n6974), .ZN(n6976)
         );
  OAI21_X1 U8739 ( .B1(n6977), .B2(n5088), .A(n6976), .ZN(P2_U3228) );
  OR2_X1 U8740 ( .A1(n6979), .A2(n6978), .ZN(n6980) );
  OAI21_X1 U8741 ( .B1(n9855), .B2(n6981), .A(n6980), .ZN(n6984) );
  INV_X1 U8742 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9857) );
  AOI22_X1 U8743 ( .A1(n7222), .A2(n9857), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n6982), .ZN(n6983) );
  NOR2_X1 U8744 ( .A1(n6984), .A2(n6983), .ZN(n7224) );
  AOI21_X1 U8745 ( .B1(n6984), .B2(n6983), .A(n7224), .ZN(n6994) );
  NOR2_X1 U8746 ( .A1(n7222), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6985) );
  AOI21_X1 U8747 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n7222), .A(n6985), .ZN(
        n6989) );
  AOI21_X1 U8748 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6987), .A(n6986), .ZN(
        n6988) );
  NAND2_X1 U8749 ( .A1(n6989), .A2(n6988), .ZN(n7218) );
  OAI21_X1 U8750 ( .B1(n6989), .B2(n6988), .A(n7218), .ZN(n6990) );
  NAND2_X1 U8751 ( .A1(n6990), .A2(n9327), .ZN(n6993) );
  INV_X1 U8752 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10100) );
  NAND2_X1 U8753 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n7489) );
  OAI21_X1 U8754 ( .B1(n9338), .B2(n10100), .A(n7489), .ZN(n6991) );
  AOI21_X1 U8755 ( .B1(n9677), .B2(n7222), .A(n6991), .ZN(n6992) );
  OAI211_X1 U8756 ( .C1(n6994), .C2(n9351), .A(n6993), .B(n6992), .ZN(P1_U3255) );
  NAND2_X1 U8757 ( .A1(n6995), .A2(n6998), .ZN(n6996) );
  XNOR2_X1 U8758 ( .A(n4514), .B(n7023), .ZN(n7029) );
  XNOR2_X1 U8759 ( .A(n7029), .B(n7039), .ZN(n6997) );
  INV_X1 U8760 ( .A(n6997), .ZN(n6999) );
  NAND3_X1 U8761 ( .A1(n6995), .A2(n6999), .A3(n6998), .ZN(n7000) );
  AOI21_X1 U8762 ( .B1(n7032), .B2(n7000), .A(n8264), .ZN(n7005) );
  INV_X1 U8763 ( .A(n7023), .ZN(n7020) );
  NOR2_X1 U8764 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5437), .ZN(n9895) );
  AOI21_X1 U8765 ( .B1(n8236), .B2(n7020), .A(n9895), .ZN(n7002) );
  AOI22_X1 U8766 ( .A1(n8258), .A2(n8290), .B1(n8269), .B2(n9971), .ZN(n7001)
         );
  OAI211_X1 U8767 ( .C1(n8247), .C2(n7003), .A(n7002), .B(n7001), .ZN(n7004)
         );
  OR2_X1 U8768 ( .A1(n7005), .A2(n7004), .ZN(P2_U3167) );
  NAND2_X1 U8769 ( .A1(n8837), .A2(n7091), .ZN(n7008) );
  INV_X1 U8770 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7006) );
  NOR2_X1 U8771 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7006), .ZN(n9674) );
  AOI21_X1 U8772 ( .B1(n8832), .B2(n9150), .A(n9674), .ZN(n7007) );
  OAI211_X1 U8773 ( .C1(n7172), .C2(n8834), .A(n7008), .B(n7007), .ZN(n7014)
         );
  INV_X1 U8774 ( .A(n7010), .ZN(n7011) );
  AOI211_X1 U8775 ( .C1(n7012), .C2(n7009), .A(n8823), .B(n7011), .ZN(n7013)
         );
  AOI211_X1 U8776 ( .C1(n9757), .C2(n8821), .A(n7014), .B(n7013), .ZN(n7015)
         );
  INV_X1 U8777 ( .A(n7015), .ZN(P1_U3230) );
  INV_X1 U8778 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10401) );
  INV_X1 U8779 ( .A(n7016), .ZN(n7027) );
  INV_X1 U8780 ( .A(n9347), .ZN(n7017) );
  OAI222_X1 U8781 ( .A1(n9632), .A2(n10401), .B1(n9634), .B2(n7027), .C1(
        P1_U3086), .C2(n7017), .ZN(P1_U3337) );
  AOI21_X1 U8782 ( .B1(n10035), .B2(n7019), .A(n7018), .ZN(n7026) );
  AOI22_X1 U8783 ( .A1(n8629), .A2(n7020), .B1(n10062), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7021) );
  OAI21_X1 U8784 ( .B1(n7026), .B2(n10062), .A(n7021), .ZN(P2_U3464) );
  INV_X1 U8785 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7022) );
  OAI22_X1 U8786 ( .A1(n8683), .A2(n7023), .B1(n7022), .B2(n10048), .ZN(n7024)
         );
  INV_X1 U8787 ( .A(n7024), .ZN(n7025) );
  OAI21_X1 U8788 ( .B1(n7026), .B2(n10049), .A(n7025), .ZN(P2_U3405) );
  INV_X1 U8789 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7028) );
  OAI222_X1 U8790 ( .A1(n8039), .A2(n7028), .B1(n8391), .B2(P2_U3151), .C1(
        n8729), .C2(n7027), .ZN(P2_U3277) );
  INV_X1 U8791 ( .A(n7029), .ZN(n7030) );
  NAND2_X1 U8792 ( .A1(n7030), .A2(n7039), .ZN(n7031) );
  NAND2_X1 U8793 ( .A1(n7032), .A2(n7031), .ZN(n7033) );
  XNOR2_X1 U8794 ( .A(n4514), .B(n10021), .ZN(n7318) );
  XNOR2_X1 U8795 ( .A(n7318), .B(n8290), .ZN(n7034) );
  AOI21_X1 U8796 ( .B1(n7033), .B2(n7034), .A(n8264), .ZN(n7037) );
  INV_X1 U8797 ( .A(n7033), .ZN(n7036) );
  INV_X1 U8798 ( .A(n7034), .ZN(n7035) );
  NAND2_X1 U8799 ( .A1(n7037), .A2(n7320), .ZN(n7042) );
  INV_X1 U8800 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7038) );
  NOR2_X1 U8801 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7038), .ZN(n9913) );
  OAI22_X1 U8802 ( .A1(n8256), .A2(n7039), .B1(n8276), .B2(n10021), .ZN(n7040)
         );
  AOI211_X1 U8803 ( .C1(n8258), .C2(n8289), .A(n9913), .B(n7040), .ZN(n7041)
         );
  OAI211_X1 U8804 ( .C1(n7213), .C2(n8247), .A(n7042), .B(n7041), .ZN(P2_U3179) );
  XNOR2_X1 U8805 ( .A(n7044), .B(n7043), .ZN(n7045) );
  NAND2_X1 U8806 ( .A1(n7045), .A2(n7046), .ZN(n7163) );
  OAI21_X1 U8807 ( .B1(n7046), .B2(n7045), .A(n7163), .ZN(n7052) );
  NOR2_X1 U8808 ( .A1(n8840), .A2(n9767), .ZN(n7051) );
  NAND2_X1 U8809 ( .A1(n8837), .A2(n7272), .ZN(n7049) );
  INV_X1 U8810 ( .A(n7279), .ZN(n9147) );
  INV_X1 U8811 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7047) );
  NOR2_X1 U8812 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7047), .ZN(n9200) );
  AOI21_X1 U8813 ( .B1(n8796), .B2(n9147), .A(n9200), .ZN(n7048) );
  OAI211_X1 U8814 ( .C1(n8798), .C2(n7127), .A(n7049), .B(n7048), .ZN(n7050)
         );
  AOI211_X1 U8815 ( .C1(n7052), .C2(n8830), .A(n7051), .B(n7050), .ZN(n7053)
         );
  INV_X1 U8816 ( .A(n7053), .ZN(P1_U3227) );
  INV_X1 U8817 ( .A(n7054), .ZN(n7057) );
  NAND3_X1 U8818 ( .A1(n7057), .A2(n7056), .A3(n7055), .ZN(n7058) );
  XNOR2_X2 U8819 ( .A(n7059), .B(n9738), .ZN(n8880) );
  INV_X1 U8820 ( .A(n7060), .ZN(n7177) );
  NAND2_X1 U8821 ( .A1(n8880), .A2(n7177), .ZN(n7176) );
  NAND2_X1 U8822 ( .A1(n4509), .A2(n6016), .ZN(n7061) );
  NAND2_X1 U8823 ( .A1(n7176), .A2(n7061), .ZN(n8975) );
  NAND2_X1 U8824 ( .A1(n7063), .A2(n9745), .ZN(n8976) );
  INV_X1 U8825 ( .A(n8976), .ZN(n7062) );
  OR2_X1 U8826 ( .A1(n8975), .A2(n7062), .ZN(n8973) );
  NAND2_X1 U8827 ( .A1(n8973), .A2(n8974), .ZN(n7064) );
  OR2_X1 U8828 ( .A1(n7085), .A2(n7075), .ZN(n8991) );
  NAND2_X1 U8829 ( .A1(n7085), .A2(n7075), .ZN(n8982) );
  NAND2_X1 U8830 ( .A1(n7064), .A2(n8884), .ZN(n7067) );
  INV_X1 U8831 ( .A(n8974), .ZN(n7065) );
  NOR2_X1 U8832 ( .A1(n8884), .A2(n7065), .ZN(n7066) );
  NAND2_X1 U8833 ( .A1(n8973), .A2(n7066), .ZN(n7088) );
  NAND2_X1 U8834 ( .A1(n7067), .A2(n7088), .ZN(n7070) );
  OAI22_X1 U8835 ( .A1(n7063), .A2(n9691), .B1(n7127), .B2(n9693), .ZN(n7069)
         );
  AOI21_X1 U8836 ( .B1(n7070), .B2(n9491), .A(n7069), .ZN(n9752) );
  OAI211_X1 U8837 ( .C1(n4731), .C2(n6072), .A(n9722), .B(n7090), .ZN(n9751)
         );
  NOR2_X1 U8838 ( .A1(n9484), .A2(n9751), .ZN(n7074) );
  OAI22_X1 U8839 ( .A1(n9534), .A2(n6767), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9522), .ZN(n7073) );
  AOI211_X1 U8840 ( .C1(n9719), .C2(n7075), .A(n7074), .B(n7073), .ZN(n7083)
         );
  NAND2_X1 U8841 ( .A1(n7076), .A2(n9357), .ZN(n7077) );
  OR2_X1 U8842 ( .A1(n9730), .A2(n7311), .ZN(n7078) );
  NAND2_X1 U8843 ( .A1(n7059), .A2(n9738), .ZN(n7079) );
  NAND2_X1 U8844 ( .A1(n7097), .A2(n7096), .ZN(n7081) );
  NAND2_X1 U8845 ( .A1(n7063), .A2(n7101), .ZN(n7080) );
  NAND2_X1 U8846 ( .A1(n7081), .A2(n7080), .ZN(n7084) );
  XNOR2_X1 U8847 ( .A(n7084), .B(n8884), .ZN(n9754) );
  NAND2_X1 U8848 ( .A1(n9486), .A2(n9754), .ZN(n7082) );
  OAI211_X1 U8849 ( .C1(n9730), .C2(n9752), .A(n7083), .B(n7082), .ZN(P1_U3290) );
  NAND2_X1 U8850 ( .A1(n7084), .A2(n8884), .ZN(n7087) );
  NAND2_X1 U8851 ( .A1(n7085), .A2(n6072), .ZN(n7086) );
  NAND2_X1 U8852 ( .A1(n7087), .A2(n7086), .ZN(n7125) );
  OR2_X1 U8853 ( .A1(n7127), .A2(n9757), .ZN(n8983) );
  NAND2_X1 U8854 ( .A1(n7127), .A2(n9757), .ZN(n8926) );
  NAND2_X1 U8855 ( .A1(n8983), .A2(n8926), .ZN(n8885) );
  INV_X1 U8856 ( .A(n8885), .ZN(n8980) );
  XNOR2_X1 U8857 ( .A(n7125), .B(n8980), .ZN(n9761) );
  NAND2_X1 U8858 ( .A1(n7088), .A2(n8982), .ZN(n7117) );
  XNOR2_X1 U8859 ( .A(n7117), .B(n8980), .ZN(n7089) );
  INV_X1 U8860 ( .A(n7172), .ZN(n9148) );
  AOI222_X1 U8861 ( .A1(n9491), .A2(n7089), .B1(n9148), .B2(n9708), .C1(n9150), 
        .C2(n9711), .ZN(n9760) );
  MUX2_X1 U8862 ( .A(n6768), .B(n9760), .S(n9534), .Z(n7095) );
  AOI211_X1 U8863 ( .C1(n9757), .C2(n7090), .A(n9541), .B(n7270), .ZN(n9756)
         );
  INV_X1 U8864 ( .A(n7091), .ZN(n7092) );
  OAI22_X1 U8865 ( .A1(n9521), .A2(n7126), .B1(n9522), .B2(n7092), .ZN(n7093)
         );
  AOI21_X1 U8866 ( .B1(n9726), .B2(n9756), .A(n7093), .ZN(n7094) );
  OAI211_X1 U8867 ( .C1(n9537), .C2(n9761), .A(n7095), .B(n7094), .ZN(P1_U3289) );
  INV_X1 U8868 ( .A(n7096), .ZN(n8882) );
  XNOR2_X1 U8869 ( .A(n7097), .B(n8882), .ZN(n9748) );
  OAI211_X1 U8870 ( .C1(n7184), .C2(n7101), .A(n9722), .B(n7098), .ZN(n7099)
         );
  INV_X1 U8871 ( .A(n7099), .ZN(n9744) );
  OAI22_X1 U8872 ( .A1(n9521), .A2(n7101), .B1(n7100), .B2(n9522), .ZN(n7102)
         );
  AOI21_X1 U8873 ( .B1(n9726), .B2(n9744), .A(n7102), .ZN(n7105) );
  XNOR2_X1 U8874 ( .A(n8975), .B(n8882), .ZN(n7103) );
  AOI222_X1 U8875 ( .A1(n9491), .A2(n7103), .B1(n9150), .B2(n9708), .C1(n9152), 
        .C2(n9711), .ZN(n9747) );
  MUX2_X1 U8876 ( .A(n6048), .B(n9747), .S(n9534), .Z(n7104) );
  OAI211_X1 U8877 ( .C1(n9537), .C2(n9748), .A(n7105), .B(n7104), .ZN(P1_U3291) );
  INV_X1 U8878 ( .A(n7107), .ZN(n7108) );
  AOI21_X1 U8879 ( .B1(n7109), .B2(n7106), .A(n7108), .ZN(n7115) );
  NAND2_X1 U8880 ( .A1(n8837), .A2(n7289), .ZN(n7112) );
  INV_X1 U8881 ( .A(n7361), .ZN(n9146) );
  INV_X1 U8882 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7110) );
  NOR2_X1 U8883 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7110), .ZN(n9226) );
  AOI21_X1 U8884 ( .B1(n8796), .B2(n9146), .A(n9226), .ZN(n7111) );
  OAI211_X1 U8885 ( .C1(n8798), .C2(n7279), .A(n7112), .B(n7111), .ZN(n7113)
         );
  AOI21_X1 U8886 ( .B1(n9779), .B2(n8821), .A(n7113), .ZN(n7114) );
  OAI21_X1 U8887 ( .B1(n7115), .B2(n8823), .A(n7114), .ZN(P1_U3213) );
  NAND2_X1 U8888 ( .A1(n9720), .A2(n7361), .ZN(n9008) );
  NAND2_X1 U8889 ( .A1(n9779), .A2(n7371), .ZN(n7245) );
  NAND2_X1 U8890 ( .A1(n9008), .A2(n7245), .ZN(n9001) );
  OR2_X1 U8891 ( .A1(n9720), .A2(n7361), .ZN(n8989) );
  AND2_X1 U8892 ( .A1(n9001), .A2(n8989), .ZN(n7246) );
  NAND2_X1 U8893 ( .A1(n7246), .A2(n9010), .ZN(n7116) );
  NAND2_X1 U8894 ( .A1(n7363), .A2(n7524), .ZN(n9021) );
  NAND2_X1 U8895 ( .A1(n7116), .A2(n9021), .ZN(n7120) );
  AND2_X1 U8896 ( .A1(n9772), .A2(n7279), .ZN(n8996) );
  NAND2_X1 U8897 ( .A1(n7117), .A2(n8980), .ZN(n7118) );
  NAND2_X1 U8898 ( .A1(n7118), .A2(n8926), .ZN(n7265) );
  OR2_X1 U8899 ( .A1(n7271), .A2(n7172), .ZN(n8997) );
  NAND2_X1 U8900 ( .A1(n7172), .A2(n7271), .ZN(n8984) );
  NAND2_X1 U8901 ( .A1(n7265), .A2(n8889), .ZN(n7119) );
  INV_X1 U8902 ( .A(n7120), .ZN(n7121) );
  NAND2_X1 U8903 ( .A1(n9010), .A2(n8989), .ZN(n9006) );
  NOR2_X1 U8904 ( .A1(n9772), .A2(n7279), .ZN(n7242) );
  NOR2_X1 U8905 ( .A1(n9779), .A2(n7371), .ZN(n8987) );
  OR3_X1 U8906 ( .A1(n9006), .A2(n7242), .A3(n8987), .ZN(n8879) );
  NAND2_X1 U8907 ( .A1(n7121), .A2(n8879), .ZN(n8928) );
  OR2_X1 U8908 ( .A1(n7526), .A2(n7300), .ZN(n9014) );
  NAND2_X1 U8909 ( .A1(n7526), .A2(n7300), .ZN(n9012) );
  OAI21_X1 U8910 ( .B1(n7122), .B2(n8890), .A(n7307), .ZN(n7124) );
  OAI22_X1 U8911 ( .A1(n7380), .A2(n9693), .B1(n7524), .B2(n9691), .ZN(n7123)
         );
  AOI21_X1 U8912 ( .B1(n7124), .B2(n9491), .A(n7123), .ZN(n9802) );
  NAND2_X1 U8913 ( .A1(n7125), .A2(n8885), .ZN(n7129) );
  NAND2_X1 U8914 ( .A1(n7127), .A2(n7126), .ZN(n7128) );
  NAND2_X1 U8915 ( .A1(n7129), .A2(n7128), .ZN(n7267) );
  INV_X1 U8916 ( .A(n8889), .ZN(n7268) );
  NAND2_X1 U8917 ( .A1(n7267), .A2(n7268), .ZN(n7131) );
  NAND2_X1 U8918 ( .A1(n9767), .A2(n7172), .ZN(n7130) );
  NAND2_X1 U8919 ( .A1(n7131), .A2(n7130), .ZN(n7153) );
  OR2_X1 U8920 ( .A1(n7242), .A2(n8996), .ZN(n7154) );
  NAND2_X1 U8921 ( .A1(n7153), .A2(n7154), .ZN(n7133) );
  OR2_X1 U8922 ( .A1(n9772), .A2(n9147), .ZN(n7132) );
  NAND2_X1 U8923 ( .A1(n7133), .A2(n7132), .ZN(n7282) );
  XNOR2_X1 U8924 ( .A(n9779), .B(n9710), .ZN(n9000) );
  INV_X1 U8925 ( .A(n9000), .ZN(n7283) );
  NAND2_X1 U8926 ( .A1(n7282), .A2(n7283), .ZN(n7135) );
  OR2_X1 U8927 ( .A1(n9779), .A2(n9710), .ZN(n7134) );
  NAND2_X1 U8928 ( .A1(n7135), .A2(n7134), .ZN(n9704) );
  NAND2_X1 U8929 ( .A1(n8989), .A2(n9008), .ZN(n9706) );
  NAND2_X1 U8930 ( .A1(n9704), .A2(n9706), .ZN(n7137) );
  OR2_X1 U8931 ( .A1(n9720), .A2(n9146), .ZN(n7136) );
  NAND2_X1 U8932 ( .A1(n7137), .A2(n7136), .ZN(n7249) );
  NAND2_X1 U8933 ( .A1(n9010), .A2(n9021), .ZN(n7250) );
  NAND2_X1 U8934 ( .A1(n7249), .A2(n7250), .ZN(n7139) );
  INV_X1 U8935 ( .A(n7524), .ZN(n9709) );
  OR2_X1 U8936 ( .A1(n7363), .A2(n9709), .ZN(n7138) );
  NAND2_X1 U8937 ( .A1(n7139), .A2(n7138), .ZN(n7299) );
  INV_X1 U8938 ( .A(n8890), .ZN(n7298) );
  XNOR2_X1 U8939 ( .A(n7299), .B(n7298), .ZN(n9804) );
  NAND2_X1 U8940 ( .A1(n9804), .A2(n9486), .ZN(n7144) );
  OAI22_X1 U8941 ( .A1(n9534), .A2(n6893), .B1(n7140), .B2(n9522), .ZN(n7142)
         );
  NAND2_X1 U8942 ( .A1(n7270), .A2(n9767), .ZN(n7269) );
  OR2_X1 U8943 ( .A1(n7269), .A2(n9772), .ZN(n7286) );
  INV_X1 U8944 ( .A(n9720), .ZN(n9787) );
  INV_X1 U8945 ( .A(n7363), .ZN(n9795) );
  OAI211_X1 U8946 ( .C1(n4608), .C2(n4741), .A(n9722), .B(n7312), .ZN(n9801)
         );
  NOR2_X1 U8947 ( .A1(n9801), .A2(n9484), .ZN(n7141) );
  AOI211_X1 U8948 ( .C1(n9719), .C2(n7526), .A(n7142), .B(n7141), .ZN(n7143)
         );
  OAI211_X1 U8949 ( .C1(n9730), .C2(n9802), .A(n7144), .B(n7143), .ZN(P1_U3283) );
  INV_X1 U8950 ( .A(n7145), .ZN(n7147) );
  OAI222_X1 U8951 ( .A1(n8039), .A2(n7146), .B1(n8729), .B2(n7147), .C1(n7850), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U8952 ( .A1(n6726), .A2(P1_U3086), .B1(n9634), .B2(n7147), .C1(
        n10214), .C2(n9632), .ZN(P1_U3336) );
  INV_X1 U8953 ( .A(n7154), .ZN(n7148) );
  XNOR2_X1 U8954 ( .A(n7243), .B(n7148), .ZN(n7149) );
  NAND2_X1 U8955 ( .A1(n7149), .A2(n9491), .ZN(n7152) );
  OAI22_X1 U8956 ( .A1(n7172), .A2(n9691), .B1(n7371), .B2(n9693), .ZN(n7150)
         );
  INV_X1 U8957 ( .A(n7150), .ZN(n7151) );
  NAND2_X1 U8958 ( .A1(n7152), .A2(n7151), .ZN(n9777) );
  INV_X1 U8959 ( .A(n9777), .ZN(n7162) );
  XNOR2_X1 U8960 ( .A(n7153), .B(n7154), .ZN(n9771) );
  AOI21_X1 U8961 ( .B1(n7269), .B2(n9772), .A(n9541), .ZN(n7155) );
  NAND2_X1 U8962 ( .A1(n7155), .A2(n7286), .ZN(n9773) );
  INV_X1 U8963 ( .A(n7169), .ZN(n7156) );
  OAI22_X1 U8964 ( .A1(n9534), .A2(n7157), .B1(n7156), .B2(n9522), .ZN(n7158)
         );
  AOI21_X1 U8965 ( .B1(n9719), .B2(n9772), .A(n7158), .ZN(n7159) );
  OAI21_X1 U8966 ( .B1(n9484), .B2(n9773), .A(n7159), .ZN(n7160) );
  AOI21_X1 U8967 ( .B1(n9486), .B2(n9771), .A(n7160), .ZN(n7161) );
  OAI21_X1 U8968 ( .B1(n7162), .B2(n9730), .A(n7161), .ZN(P1_U3287) );
  OAI21_X1 U8969 ( .B1(n7164), .B2(n7043), .A(n7163), .ZN(n7168) );
  XNOR2_X1 U8970 ( .A(n7166), .B(n7165), .ZN(n7167) );
  XNOR2_X1 U8971 ( .A(n7168), .B(n7167), .ZN(n7175) );
  NAND2_X1 U8972 ( .A1(n8837), .A2(n7169), .ZN(n7171) );
  AND2_X1 U8973 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9213) );
  AOI21_X1 U8974 ( .B1(n8796), .B2(n9710), .A(n9213), .ZN(n7170) );
  OAI211_X1 U8975 ( .C1(n8798), .C2(n7172), .A(n7171), .B(n7170), .ZN(n7173)
         );
  AOI21_X1 U8976 ( .B1(n9772), .B2(n8821), .A(n7173), .ZN(n7174) );
  OAI21_X1 U8977 ( .B1(n7175), .B2(n8823), .A(n7174), .ZN(P1_U3239) );
  OAI21_X1 U8978 ( .B1(n7177), .B2(n8880), .A(n7176), .ZN(n7183) );
  OAI22_X1 U8979 ( .A1(n7063), .A2(n9693), .B1(n7178), .B2(n9691), .ZN(n7182)
         );
  XNOR2_X1 U8980 ( .A(n8880), .B(n7179), .ZN(n9742) );
  INV_X1 U8981 ( .A(n9742), .ZN(n7180) );
  NOR2_X1 U8982 ( .A1(n7180), .A2(n7311), .ZN(n7181) );
  AOI211_X1 U8983 ( .C1(n9491), .C2(n7183), .A(n7182), .B(n7181), .ZN(n9739)
         );
  INV_X1 U8984 ( .A(n7317), .ZN(n9727) );
  INV_X1 U8985 ( .A(n7184), .ZN(n7185) );
  OAI211_X1 U8986 ( .C1(n9738), .C2(n7186), .A(n7185), .B(n9722), .ZN(n9737)
         );
  OAI22_X1 U8987 ( .A1(n9534), .A2(n6009), .B1(n9156), .B2(n9522), .ZN(n7187)
         );
  AOI21_X1 U8988 ( .B1(n9719), .B2(n6016), .A(n7187), .ZN(n7188) );
  OAI21_X1 U8989 ( .B1(n9484), .B2(n9737), .A(n7188), .ZN(n7189) );
  AOI21_X1 U8990 ( .B1(n9727), .B2(n9742), .A(n7189), .ZN(n7190) );
  OAI21_X1 U8991 ( .B1(n9730), .B2(n9739), .A(n7190), .ZN(P1_U3292) );
  AOI21_X1 U8992 ( .B1(n7460), .B2(n7192), .A(n4503), .ZN(n7205) );
  AOI21_X1 U8993 ( .B1(n10060), .B2(n7194), .A(n7193), .ZN(n7195) );
  NOR2_X1 U8994 ( .A1(n7195), .A2(n9953), .ZN(n7203) );
  NOR2_X1 U8995 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5514), .ZN(n7543) );
  INV_X1 U8996 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10087) );
  OAI22_X1 U8997 ( .A1(n9957), .A2(n7196), .B1(n9969), .B2(n10087), .ZN(n7202)
         );
  AOI21_X1 U8998 ( .B1(n7199), .B2(n7198), .A(n7197), .ZN(n7200) );
  NOR2_X1 U8999 ( .A1(n7200), .A2(n7442), .ZN(n7201) );
  NOR4_X1 U9000 ( .A1(n7203), .A2(n7543), .A3(n7202), .A4(n7201), .ZN(n7204)
         );
  OAI21_X1 U9001 ( .B1(n7205), .B2(n9948), .A(n7204), .ZN(P2_U3191) );
  NAND2_X1 U9002 ( .A1(n8292), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7206) );
  OAI21_X1 U9003 ( .B1(n8142), .B2(n8292), .A(n7206), .ZN(P2_U3520) );
  NAND2_X1 U9004 ( .A1(n7208), .A2(n7207), .ZN(n7209) );
  XNOR2_X1 U9005 ( .A(n7331), .B(n7215), .ZN(n7831) );
  XNOR2_X1 U9006 ( .A(n7209), .B(n7831), .ZN(n10023) );
  INV_X1 U9007 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7212) );
  XNOR2_X1 U9008 ( .A(n7210), .B(n7831), .ZN(n7211) );
  AOI222_X1 U9009 ( .A1(n9981), .A2(n7211), .B1(n8289), .B2(n9983), .C1(n8291), 
        .C2(n9986), .ZN(n10020) );
  MUX2_X1 U9010 ( .A(n7212), .B(n10020), .S(n9999), .Z(n7217) );
  INV_X1 U9011 ( .A(n7213), .ZN(n7214) );
  AOI22_X1 U9012 ( .A1(n8555), .A2(n7215), .B1(n8554), .B2(n7214), .ZN(n7216)
         );
  OAI211_X1 U9013 ( .C1(n10023), .C2(n8558), .A(n7217), .B(n7216), .ZN(
        P2_U3227) );
  OAI21_X1 U9014 ( .B1(n7222), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7218), .ZN(
        n7221) );
  NAND2_X1 U9015 ( .A1(n9260), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7219) );
  OAI21_X1 U9016 ( .B1(n9260), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7219), .ZN(
        n7220) );
  NOR2_X1 U9017 ( .A1(n7220), .A2(n7221), .ZN(n9259) );
  AOI211_X1 U9018 ( .C1(n7221), .C2(n7220), .A(n9259), .B(n9672), .ZN(n7232)
         );
  NOR2_X1 U9019 ( .A1(n7222), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7223) );
  NOR2_X1 U9020 ( .A1(n7224), .A2(n7223), .ZN(n7227) );
  INV_X1 U9021 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7225) );
  MUX2_X1 U9022 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7225), .S(n9260), .Z(n7226)
         );
  NAND2_X1 U9023 ( .A1(n7226), .A2(n7227), .ZN(n9254) );
  OAI211_X1 U9024 ( .C1(n7227), .C2(n7226), .A(n9679), .B(n9254), .ZN(n7230)
         );
  NAND2_X1 U9025 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n7575) );
  INV_X1 U9026 ( .A(n7575), .ZN(n7228) );
  AOI21_X1 U9027 ( .B1(n9675), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7228), .ZN(
        n7229) );
  OAI211_X1 U9028 ( .C1(n9354), .C2(n9255), .A(n7230), .B(n7229), .ZN(n7231)
         );
  OR2_X1 U9029 ( .A1(n7232), .A2(n7231), .ZN(P1_U3256) );
  NAND2_X1 U9030 ( .A1(n9726), .A2(n9722), .ZN(n9365) );
  INV_X1 U9031 ( .A(n9365), .ZN(n7234) );
  OAI21_X1 U9032 ( .B1(n7234), .B2(n9719), .A(n7233), .ZN(n7241) );
  NOR2_X1 U9033 ( .A1(n9522), .A2(n7235), .ZN(n7239) );
  OAI21_X1 U9034 ( .B1(n8883), .B2(n7237), .A(n7236), .ZN(n7238) );
  OAI21_X1 U9035 ( .B1(n7239), .B2(n7238), .A(n9534), .ZN(n7240) );
  OAI211_X1 U9036 ( .C1(n9534), .C2(n6024), .A(n7241), .B(n7240), .ZN(P1_U3293) );
  INV_X1 U9037 ( .A(n7242), .ZN(n8999) );
  NAND2_X1 U9038 ( .A1(n7243), .A2(n8999), .ZN(n7244) );
  INV_X1 U9039 ( .A(n8996), .ZN(n8985) );
  NAND2_X1 U9040 ( .A1(n7244), .A2(n8985), .ZN(n7278) );
  NAND2_X1 U9041 ( .A1(n7278), .A2(n9000), .ZN(n7277) );
  AND2_X1 U9042 ( .A1(n7277), .A2(n7245), .ZN(n9707) );
  NOR2_X1 U9043 ( .A1(n9707), .A2(n9706), .ZN(n9705) );
  NOR2_X1 U9044 ( .A1(n9705), .A2(n7246), .ZN(n7247) );
  XNOR2_X1 U9045 ( .A(n7247), .B(n7250), .ZN(n7248) );
  AOI22_X1 U9046 ( .A1(n7248), .A2(n9491), .B1(n9711), .B2(n9146), .ZN(n9796)
         );
  XNOR2_X1 U9047 ( .A(n7249), .B(n7250), .ZN(n9799) );
  XNOR2_X1 U9048 ( .A(n9721), .B(n9795), .ZN(n7251) );
  OAI22_X1 U9049 ( .A1(n7251), .A2(n9541), .B1(n7300), .B2(n9693), .ZN(n9793)
         );
  NAND2_X1 U9050 ( .A1(n9793), .A2(n9726), .ZN(n7253) );
  AOI22_X1 U9051 ( .A1(n9730), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7357), .B2(
        n9718), .ZN(n7252) );
  OAI211_X1 U9052 ( .C1(n9795), .C2(n9521), .A(n7253), .B(n7252), .ZN(n7254)
         );
  AOI21_X1 U9053 ( .B1(n9799), .B2(n9486), .A(n7254), .ZN(n7255) );
  OAI21_X1 U9054 ( .B1(n9796), .B2(n9730), .A(n7255), .ZN(P1_U3284) );
  NAND2_X1 U9055 ( .A1(n7256), .A2(n7829), .ZN(n7257) );
  NAND2_X1 U9056 ( .A1(n7411), .A2(n7257), .ZN(n10027) );
  INV_X1 U9057 ( .A(n7829), .ZN(n7896) );
  XNOR2_X1 U9058 ( .A(n7258), .B(n7896), .ZN(n7259) );
  NAND2_X1 U9059 ( .A1(n7259), .A2(n9981), .ZN(n7261) );
  AOI22_X1 U9060 ( .A1(n8290), .A2(n9986), .B1(n9983), .B2(n8288), .ZN(n7260)
         );
  OAI211_X1 U9061 ( .C1(n7502), .C2(n10027), .A(n7261), .B(n7260), .ZN(n10029)
         );
  NAND2_X1 U9062 ( .A1(n10029), .A2(n9999), .ZN(n7264) );
  OAI22_X1 U9063 ( .A1(n9999), .A2(n9929), .B1(n7327), .B2(n9990), .ZN(n7262)
         );
  AOI21_X1 U9064 ( .B1(n8555), .B2(n7321), .A(n7262), .ZN(n7263) );
  OAI211_X1 U9065 ( .C1(n10027), .C2(n7507), .A(n7264), .B(n7263), .ZN(
        P2_U3226) );
  XNOR2_X1 U9066 ( .A(n7265), .B(n8889), .ZN(n7266) );
  AOI222_X1 U9067 ( .A1(n9491), .A2(n7266), .B1(n9147), .B2(n9708), .C1(n9149), 
        .C2(n9711), .ZN(n9766) );
  XNOR2_X1 U9068 ( .A(n7267), .B(n7268), .ZN(n9769) );
  OAI211_X1 U9069 ( .C1(n7270), .C2(n9767), .A(n9722), .B(n7269), .ZN(n9765)
         );
  NAND2_X1 U9070 ( .A1(n9719), .A2(n7271), .ZN(n7274) );
  AOI22_X1 U9071 ( .A1(n9730), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7272), .B2(
        n9718), .ZN(n7273) );
  OAI211_X1 U9072 ( .C1(n9765), .C2(n9484), .A(n7274), .B(n7273), .ZN(n7275)
         );
  AOI21_X1 U9073 ( .B1(n9486), .B2(n9769), .A(n7275), .ZN(n7276) );
  OAI21_X1 U9074 ( .B1(n9766), .B2(n9730), .A(n7276), .ZN(P1_U3288) );
  OAI21_X1 U9075 ( .B1(n7278), .B2(n9000), .A(n7277), .ZN(n7281) );
  OAI22_X1 U9076 ( .A1(n7279), .A2(n9691), .B1(n7361), .B2(n9693), .ZN(n7280)
         );
  AOI21_X1 U9077 ( .B1(n7281), .B2(n9491), .A(n7280), .ZN(n7285) );
  XNOR2_X1 U9078 ( .A(n7282), .B(n7283), .ZN(n9782) );
  INV_X1 U9079 ( .A(n7311), .ZN(n9716) );
  NAND2_X1 U9080 ( .A1(n9782), .A2(n9716), .ZN(n7284) );
  AND2_X1 U9081 ( .A1(n7285), .A2(n7284), .ZN(n9784) );
  NAND2_X1 U9082 ( .A1(n7286), .A2(n9779), .ZN(n7287) );
  NAND2_X1 U9083 ( .A1(n7287), .A2(n9722), .ZN(n7288) );
  OR2_X1 U9084 ( .A1(n7288), .A2(n9724), .ZN(n9780) );
  NAND2_X1 U9085 ( .A1(n9719), .A2(n9779), .ZN(n7291) );
  AOI22_X1 U9086 ( .A1(n9730), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7289), .B2(
        n9718), .ZN(n7290) );
  OAI211_X1 U9087 ( .C1(n9780), .C2(n9484), .A(n7291), .B(n7290), .ZN(n7292)
         );
  AOI21_X1 U9088 ( .B1(n9782), .B2(n9727), .A(n7292), .ZN(n7293) );
  OAI21_X1 U9089 ( .B1(n9784), .B2(n9730), .A(n7293), .ZN(P1_U3286) );
  INV_X1 U9090 ( .A(n7294), .ZN(n7297) );
  OAI222_X1 U9091 ( .A1(n8729), .A2(n7297), .B1(P2_U3151), .B2(n7852), .C1(
        n7295), .C2(n8723), .ZN(P2_U3275) );
  INV_X1 U9092 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7296) );
  OAI222_X1 U9093 ( .A1(P1_U3086), .A2(n8914), .B1(n9634), .B2(n7297), .C1(
        n7296), .C2(n9632), .ZN(P1_U3335) );
  NAND2_X1 U9094 ( .A1(n7299), .A2(n7298), .ZN(n7302) );
  INV_X1 U9095 ( .A(n7300), .ZN(n9145) );
  OR2_X1 U9096 ( .A1(n7526), .A2(n9145), .ZN(n7301) );
  NAND2_X1 U9097 ( .A1(n7302), .A2(n7301), .ZN(n7379) );
  OR2_X1 U9098 ( .A1(n7569), .A2(n7380), .ZN(n9015) );
  NAND2_X1 U9099 ( .A1(n7569), .A2(n7380), .ZN(n9017) );
  XNOR2_X1 U9100 ( .A(n7303), .B(n8894), .ZN(n9806) );
  INV_X1 U9101 ( .A(n9027), .ZN(n9143) );
  AOI22_X1 U9102 ( .A1(n9708), .A2(n9143), .B1(n9145), .B2(n9711), .ZN(n7310)
         );
  INV_X1 U9103 ( .A(n7307), .ZN(n7304) );
  INV_X1 U9104 ( .A(n9012), .ZN(n7305) );
  INV_X1 U9105 ( .A(n8894), .ZN(n7378) );
  OAI21_X1 U9106 ( .B1(n7304), .B2(n7305), .A(n7378), .ZN(n7308) );
  NAND2_X1 U9107 ( .A1(n7307), .A2(n7306), .ZN(n7382) );
  NAND3_X1 U9108 ( .A1(n7308), .A2(n7382), .A3(n9491), .ZN(n7309) );
  OAI211_X1 U9109 ( .C1(n9806), .C2(n7311), .A(n7310), .B(n7309), .ZN(n9810)
         );
  NAND2_X1 U9110 ( .A1(n9810), .A2(n9534), .ZN(n7316) );
  AOI211_X1 U9111 ( .C1(n7569), .C2(n7312), .A(n9541), .B(n7397), .ZN(n9807)
         );
  INV_X1 U9112 ( .A(n7569), .ZN(n9809) );
  AOI22_X1 U9113 ( .A1(n9730), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7568), .B2(
        n9718), .ZN(n7313) );
  OAI21_X1 U9114 ( .B1(n9809), .B2(n9521), .A(n7313), .ZN(n7314) );
  AOI21_X1 U9115 ( .B1(n9807), .B2(n9726), .A(n7314), .ZN(n7315) );
  OAI211_X1 U9116 ( .C1(n9806), .C2(n7317), .A(n7316), .B(n7315), .ZN(P1_U3282) );
  NAND2_X1 U9117 ( .A1(n7318), .A2(n8290), .ZN(n7319) );
  XNOR2_X1 U9118 ( .A(n4514), .B(n7321), .ZN(n7322) );
  INV_X1 U9119 ( .A(n8289), .ZN(n7421) );
  NAND2_X1 U9120 ( .A1(n7322), .A2(n7421), .ZN(n7424) );
  INV_X1 U9121 ( .A(n7322), .ZN(n7323) );
  NAND2_X1 U9122 ( .A1(n7323), .A2(n8289), .ZN(n7324) );
  AND2_X1 U9123 ( .A1(n7424), .A2(n7324), .ZN(n7325) );
  OAI21_X1 U9124 ( .B1(n7326), .B2(n7325), .A(n7422), .ZN(n7334) );
  NOR2_X1 U9125 ( .A1(n8276), .A2(n10026), .ZN(n7333) );
  NOR2_X1 U9126 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5482), .ZN(n9934) );
  AOI21_X1 U9127 ( .B1(n8258), .B2(n8288), .A(n9934), .ZN(n7330) );
  INV_X1 U9128 ( .A(n7327), .ZN(n7328) );
  NAND2_X1 U9129 ( .A1(n8273), .A2(n7328), .ZN(n7329) );
  OAI211_X1 U9130 ( .C1(n8256), .C2(n7331), .A(n7330), .B(n7329), .ZN(n7332)
         );
  AOI211_X1 U9131 ( .C1(n7334), .C2(n8244), .A(n7333), .B(n7332), .ZN(n7335)
         );
  INV_X1 U9132 ( .A(n7335), .ZN(P2_U3153) );
  AOI21_X1 U9133 ( .B1(n7338), .B2(n7337), .A(n7336), .ZN(n7352) );
  AOI21_X1 U9134 ( .B1(n7341), .B2(n7340), .A(n7339), .ZN(n7342) );
  NOR2_X1 U9135 ( .A1(n7342), .A2(n9953), .ZN(n7350) );
  INV_X1 U9136 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10470) );
  NOR2_X1 U9137 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10470), .ZN(n7625) );
  INV_X1 U9138 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10091) );
  OAI22_X1 U9139 ( .A1(n9957), .A2(n7343), .B1(n9969), .B2(n10091), .ZN(n7349)
         );
  AOI21_X1 U9140 ( .B1(n7346), .B2(n7345), .A(n7344), .ZN(n7347) );
  NOR2_X1 U9141 ( .A1(n7347), .A2(n7442), .ZN(n7348) );
  NOR4_X1 U9142 ( .A1(n7350), .A2(n7625), .A3(n7349), .A4(n7348), .ZN(n7351)
         );
  OAI21_X1 U9143 ( .B1(n7352), .B2(n9948), .A(n7351), .ZN(P2_U3192) );
  NAND2_X1 U9144 ( .A1(n7353), .A2(n8830), .ZN(n7366) );
  AOI21_X1 U9145 ( .B1(n7354), .B2(n7356), .A(n7355), .ZN(n7365) );
  NAND2_X1 U9146 ( .A1(n8837), .A2(n7357), .ZN(n7360) );
  AOI21_X1 U9147 ( .B1(n8796), .B2(n9145), .A(n7358), .ZN(n7359) );
  OAI211_X1 U9148 ( .C1(n8798), .C2(n7361), .A(n7360), .B(n7359), .ZN(n7362)
         );
  AOI21_X1 U9149 ( .B1(n7363), .B2(n8821), .A(n7362), .ZN(n7364) );
  OAI21_X1 U9150 ( .B1(n7366), .B2(n7365), .A(n7364), .ZN(P1_U3231) );
  OAI21_X1 U9151 ( .B1(n7368), .B2(n7367), .A(n7354), .ZN(n7374) );
  NOR2_X1 U9152 ( .A1(n8840), .A2(n9787), .ZN(n7373) );
  NAND2_X1 U9153 ( .A1(n8837), .A2(n9717), .ZN(n7370) );
  AND2_X1 U9154 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9239) );
  AOI21_X1 U9155 ( .B1(n8796), .B2(n9709), .A(n9239), .ZN(n7369) );
  OAI211_X1 U9156 ( .C1(n8798), .C2(n7371), .A(n7370), .B(n7369), .ZN(n7372)
         );
  AOI211_X1 U9157 ( .C1(n7374), .C2(n8830), .A(n7373), .B(n7372), .ZN(n7375)
         );
  INV_X1 U9158 ( .A(n7375), .ZN(P1_U3221) );
  INV_X1 U9159 ( .A(n7376), .ZN(n7394) );
  OAI222_X1 U9160 ( .A1(n8729), .A2(n7394), .B1(P2_U3151), .B2(n7856), .C1(
        n7377), .C2(n8723), .ZN(P2_U3274) );
  INV_X1 U9161 ( .A(n7380), .ZN(n9144) );
  OR2_X1 U9162 ( .A1(n7569), .A2(n9144), .ZN(n7381) );
  OR2_X1 U9163 ( .A1(n9031), .A2(n9027), .ZN(n8933) );
  NAND2_X1 U9164 ( .A1(n9031), .A2(n9027), .ZN(n9018) );
  OR2_X1 U9165 ( .A1(n7470), .A2(n9692), .ZN(n9041) );
  NAND2_X1 U9166 ( .A1(n7470), .A2(n9692), .ZN(n9043) );
  XNOR2_X1 U9167 ( .A(n7469), .B(n7468), .ZN(n9825) );
  INV_X1 U9168 ( .A(n9825), .ZN(n7393) );
  AND2_X1 U9169 ( .A1(n9043), .A2(n9018), .ZN(n7383) );
  NAND2_X1 U9170 ( .A1(n7402), .A2(n9018), .ZN(n7384) );
  NAND2_X1 U9171 ( .A1(n7384), .A2(n7468), .ZN(n7385) );
  OAI211_X1 U9172 ( .C1(n7476), .C2(n4766), .A(n7385), .B(n9491), .ZN(n7388)
         );
  OAI22_X1 U9173 ( .A1(n7577), .A2(n9693), .B1(n9027), .B2(n9691), .ZN(n7386)
         );
  INV_X1 U9174 ( .A(n7386), .ZN(n7387) );
  NAND2_X1 U9175 ( .A1(n7388), .A2(n7387), .ZN(n9823) );
  INV_X1 U9176 ( .A(n7470), .ZN(n9821) );
  INV_X1 U9177 ( .A(n9031), .ZN(n9816) );
  OAI211_X1 U9178 ( .C1(n9821), .C2(n7398), .A(n9722), .B(n9698), .ZN(n9820)
         );
  AOI22_X1 U9179 ( .A1(n9730), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7580), .B2(
        n9718), .ZN(n7390) );
  NAND2_X1 U9180 ( .A1(n7470), .A2(n9719), .ZN(n7389) );
  OAI211_X1 U9181 ( .C1(n9820), .C2(n9484), .A(n7390), .B(n7389), .ZN(n7391)
         );
  AOI21_X1 U9182 ( .B1(n9823), .B2(n9534), .A(n7391), .ZN(n7392) );
  OAI21_X1 U9183 ( .B1(n7393), .B2(n9537), .A(n7392), .ZN(P1_U3280) );
  INV_X1 U9184 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10413) );
  OAI222_X1 U9185 ( .A1(P1_U3086), .A2(n8881), .B1(n9634), .B2(n7394), .C1(
        n10413), .C2(n9632), .ZN(P1_U3334) );
  XNOR2_X1 U9186 ( .A(n7395), .B(n7396), .ZN(n9818) );
  OAI21_X1 U9187 ( .B1(n7397), .B2(n9816), .A(n9722), .ZN(n7399) );
  OR2_X1 U9188 ( .A1(n7399), .A2(n7398), .ZN(n9814) );
  AOI22_X1 U9189 ( .A1(n9730), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7493), .B2(
        n9718), .ZN(n7401) );
  NAND2_X1 U9190 ( .A1(n9031), .A2(n9719), .ZN(n7400) );
  OAI211_X1 U9191 ( .C1(n9814), .C2(n9484), .A(n7401), .B(n7400), .ZN(n7406)
         );
  OAI21_X1 U9192 ( .B1(n7403), .B2(n8893), .A(n7402), .ZN(n7404) );
  INV_X1 U9193 ( .A(n9692), .ZN(n9142) );
  AOI222_X1 U9194 ( .A1(n9491), .A2(n7404), .B1(n9142), .B2(n9708), .C1(n9144), 
        .C2(n9711), .ZN(n9815) );
  NOR2_X1 U9195 ( .A1(n9815), .A2(n9730), .ZN(n7405) );
  AOI211_X1 U9196 ( .C1(n9486), .C2(n9818), .A(n7406), .B(n7405), .ZN(n7407)
         );
  INV_X1 U9197 ( .A(n7407), .ZN(P1_U3281) );
  NAND2_X1 U9198 ( .A1(n7899), .A2(n7886), .ZN(n7830) );
  XOR2_X1 U9199 ( .A(n7408), .B(n7830), .Z(n7409) );
  OAI222_X1 U9200 ( .A1(n8565), .A2(n7616), .B1(n8563), .B2(n7421), .C1(n8561), 
        .C2(n7409), .ZN(n10032) );
  INV_X1 U9201 ( .A(n10032), .ZN(n7416) );
  NAND2_X1 U9202 ( .A1(n7411), .A2(n7410), .ZN(n7412) );
  XNOR2_X1 U9203 ( .A(n7412), .B(n7830), .ZN(n10034) );
  NOR2_X1 U9204 ( .A1(n9975), .A2(n10031), .ZN(n7414) );
  OAI22_X1 U9205 ( .A1(n9999), .A2(n5282), .B1(n7417), .B2(n9990), .ZN(n7413)
         );
  AOI211_X1 U9206 ( .C1(n10034), .C2(n9977), .A(n7414), .B(n7413), .ZN(n7415)
         );
  OAI21_X1 U9207 ( .B1(n7416), .B2(n5088), .A(n7415), .ZN(P2_U3225) );
  AND2_X1 U9208 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9959) );
  AOI21_X1 U9209 ( .B1(n8258), .B2(n7626), .A(n9959), .ZN(n7420) );
  INV_X1 U9210 ( .A(n7417), .ZN(n7418) );
  NAND2_X1 U9211 ( .A1(n8273), .A2(n7418), .ZN(n7419) );
  OAI211_X1 U9212 ( .C1(n8256), .C2(n7421), .A(n7420), .B(n7419), .ZN(n7428)
         );
  XNOR2_X1 U9213 ( .A(n4511), .B(n10031), .ZN(n7546) );
  XNOR2_X1 U9214 ( .A(n7546), .B(n7547), .ZN(n7423) );
  INV_X1 U9215 ( .A(n7423), .ZN(n7425) );
  NAND3_X1 U9216 ( .A1(n7422), .A2(n7425), .A3(n7424), .ZN(n7426) );
  AOI21_X1 U9217 ( .B1(n7550), .B2(n7426), .A(n8264), .ZN(n7427) );
  AOI211_X1 U9218 ( .C1(n7429), .C2(n8236), .A(n7428), .B(n7427), .ZN(n7430)
         );
  INV_X1 U9219 ( .A(n7430), .ZN(P2_U3161) );
  AOI21_X1 U9220 ( .B1(n7432), .B2(n7536), .A(n7431), .ZN(n7449) );
  INV_X1 U9221 ( .A(n7433), .ZN(n7434) );
  NOR2_X1 U9222 ( .A1(n7434), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7437) );
  OAI21_X1 U9223 ( .B1(n7437), .B2(n7436), .A(n7435), .ZN(n7448) );
  INV_X1 U9224 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10095) );
  NOR2_X1 U9225 ( .A1(n9969), .A2(n10095), .ZN(n7445) );
  AOI21_X1 U9226 ( .B1(n7440), .B2(n7439), .A(n7438), .ZN(n7443) );
  INV_X1 U9227 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10389) );
  NOR2_X1 U9228 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10389), .ZN(n7640) );
  INV_X1 U9229 ( .A(n7640), .ZN(n7441) );
  OAI21_X1 U9230 ( .B1(n7443), .B2(n7442), .A(n7441), .ZN(n7444) );
  AOI211_X1 U9231 ( .C1(n7446), .C2(n9915), .A(n7445), .B(n7444), .ZN(n7447)
         );
  OAI211_X1 U9232 ( .C1(n7449), .C2(n9948), .A(n7448), .B(n7447), .ZN(P2_U3193) );
  OR2_X1 U9233 ( .A1(n7450), .A2(n7834), .ZN(n7451) );
  NAND2_X1 U9234 ( .A1(n7452), .A2(n7451), .ZN(n10036) );
  INV_X1 U9235 ( .A(n7453), .ZN(n7456) );
  INV_X1 U9236 ( .A(n7834), .ZN(n7455) );
  OAI21_X1 U9237 ( .B1(n7456), .B2(n7455), .A(n7454), .ZN(n7457) );
  NAND2_X1 U9238 ( .A1(n7457), .A2(n9981), .ZN(n7459) );
  AOI22_X1 U9239 ( .A1(n9986), .A2(n8288), .B1(n8287), .B2(n9983), .ZN(n7458)
         );
  OAI211_X1 U9240 ( .C1(n7502), .C2(n10036), .A(n7459), .B(n7458), .ZN(n10037)
         );
  NAND2_X1 U9241 ( .A1(n10037), .A2(n9999), .ZN(n7463) );
  OAI22_X1 U9242 ( .A1(n9999), .A2(n7460), .B1(n7541), .B2(n9990), .ZN(n7461)
         );
  AOI21_X1 U9243 ( .B1(n8555), .B2(n10039), .A(n7461), .ZN(n7462) );
  OAI211_X1 U9244 ( .C1(n10036), .C2(n7507), .A(n7463), .B(n7462), .ZN(
        P2_U3224) );
  INV_X1 U9245 ( .A(n7464), .ZN(n7467) );
  OAI222_X1 U9246 ( .A1(n8039), .A2(n7466), .B1(n8729), .B2(n7467), .C1(n7465), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U9247 ( .A1(n6525), .A2(P1_U3086), .B1(n9634), .B2(n7467), .C1(
        n10415), .C2(n9632), .ZN(P1_U3333) );
  NAND2_X1 U9248 ( .A1(n7469), .A2(n7468), .ZN(n7472) );
  OR2_X1 U9249 ( .A1(n7470), .A2(n9142), .ZN(n7471) );
  NAND2_X1 U9250 ( .A1(n7472), .A2(n7471), .ZN(n9686) );
  NOR2_X1 U9251 ( .A1(n9699), .A2(n9141), .ZN(n7473) );
  OR2_X2 U9252 ( .A1(n9686), .A2(n7473), .ZN(n7475) );
  NAND2_X1 U9253 ( .A1(n9699), .A2(n9141), .ZN(n7474) );
  OR2_X1 U9254 ( .A1(n7609), .A2(n9694), .ZN(n9046) );
  NAND2_X1 U9255 ( .A1(n7609), .A2(n9694), .ZN(n9047) );
  XNOR2_X1 U9256 ( .A(n7608), .B(n8899), .ZN(n9653) );
  INV_X1 U9257 ( .A(n9653), .ZN(n7486) );
  OR2_X1 U9258 ( .A1(n9699), .A2(n7577), .ZN(n9045) );
  NAND2_X1 U9259 ( .A1(n9699), .A2(n7577), .ZN(n9044) );
  NAND2_X1 U9260 ( .A1(n9045), .A2(n9044), .ZN(n9687) );
  OAI211_X1 U9261 ( .C1(n7477), .C2(n8899), .A(n7600), .B(n9491), .ZN(n7479)
         );
  AOI22_X1 U9262 ( .A1(n9141), .A2(n9711), .B1(n9140), .B2(n9708), .ZN(n7478)
         );
  NAND2_X1 U9263 ( .A1(n7479), .A2(n7478), .ZN(n9652) );
  OAI211_X1 U9264 ( .C1(n7480), .C2(n7481), .A(n9722), .B(n7604), .ZN(n9650)
         );
  AOI22_X1 U9265 ( .A1(n9730), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7760), .B2(
        n9718), .ZN(n7483) );
  NAND2_X1 U9266 ( .A1(n7609), .A2(n9719), .ZN(n7482) );
  OAI211_X1 U9267 ( .C1(n9650), .C2(n9484), .A(n7483), .B(n7482), .ZN(n7484)
         );
  AOI21_X1 U9268 ( .B1(n9652), .B2(n9534), .A(n7484), .ZN(n7485) );
  OAI21_X1 U9269 ( .B1(n7486), .B2(n9537), .A(n7485), .ZN(P1_U3278) );
  XOR2_X1 U9270 ( .A(n7487), .B(n7488), .Z(n7495) );
  NAND2_X1 U9271 ( .A1(n8832), .A2(n9144), .ZN(n7490) );
  OAI211_X1 U9272 ( .C1(n9692), .C2(n8834), .A(n7490), .B(n7489), .ZN(n7492)
         );
  NOR2_X1 U9273 ( .A1(n9816), .A2(n8840), .ZN(n7491) );
  AOI211_X1 U9274 ( .C1(n8837), .C2(n7493), .A(n7492), .B(n7491), .ZN(n7494)
         );
  OAI21_X1 U9275 ( .B1(n7495), .B2(n8823), .A(n7494), .ZN(P1_U3224) );
  INV_X1 U9276 ( .A(n7908), .ZN(n7496) );
  NOR2_X1 U9277 ( .A1(n7911), .A2(n7496), .ZN(n7835) );
  XNOR2_X1 U9278 ( .A(n7497), .B(n7835), .ZN(n10045) );
  XOR2_X1 U9279 ( .A(n7835), .B(n7498), .Z(n7499) );
  NAND2_X1 U9280 ( .A1(n7499), .A2(n9981), .ZN(n7501) );
  AOI22_X1 U9281 ( .A1(n9986), .A2(n7626), .B1(n8162), .B2(n9983), .ZN(n7500)
         );
  OAI211_X1 U9282 ( .C1(n10045), .C2(n7502), .A(n7501), .B(n7500), .ZN(n10047)
         );
  NAND2_X1 U9283 ( .A1(n10047), .A2(n9999), .ZN(n7506) );
  INV_X1 U9284 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7503) );
  OAI22_X1 U9285 ( .A1(n9999), .A2(n7503), .B1(n7623), .B2(n9990), .ZN(n7504)
         );
  AOI21_X1 U9286 ( .B1(n8555), .B2(n7620), .A(n7504), .ZN(n7505) );
  OAI211_X1 U9287 ( .C1(n10045), .C2(n7507), .A(n7506), .B(n7505), .ZN(
        P2_U3223) );
  NAND2_X1 U9288 ( .A1(n7511), .A2(n7508), .ZN(n7510) );
  OR2_X1 U9289 ( .A1(n7509), .A2(P1_U3086), .ZN(n9131) );
  OAI211_X1 U9290 ( .C1(n10489), .C2(n9632), .A(n7510), .B(n9131), .ZN(
        P1_U3332) );
  NAND2_X1 U9291 ( .A1(n7511), .A2(n7733), .ZN(n7512) );
  OAI211_X1 U9292 ( .C1(n7513), .C2(n8723), .A(n7512), .B(n8030), .ZN(P2_U3272) );
  INV_X1 U9293 ( .A(n7514), .ZN(n7515) );
  NOR2_X1 U9294 ( .A1(n7516), .A2(n7515), .ZN(n7559) );
  AOI21_X1 U9295 ( .B1(n7516), .B2(n7515), .A(n7559), .ZN(n7517) );
  NAND2_X1 U9296 ( .A1(n7517), .A2(n7518), .ZN(n7561) );
  OAI21_X1 U9297 ( .B1(n7518), .B2(n7517), .A(n7561), .ZN(n7519) );
  NAND2_X1 U9298 ( .A1(n7519), .A2(n8830), .ZN(n7528) );
  NAND2_X1 U9299 ( .A1(n8837), .A2(n7520), .ZN(n7523) );
  AOI21_X1 U9300 ( .B1(n8796), .B2(n9144), .A(n7521), .ZN(n7522) );
  OAI211_X1 U9301 ( .C1(n8798), .C2(n7524), .A(n7523), .B(n7522), .ZN(n7525)
         );
  AOI21_X1 U9302 ( .B1(n7526), .B2(n8821), .A(n7525), .ZN(n7527) );
  NAND2_X1 U9303 ( .A1(n7528), .A2(n7527), .ZN(P1_U3217) );
  INV_X1 U9304 ( .A(n7529), .ZN(n7641) );
  OR2_X1 U9305 ( .A1(n7530), .A2(n7636), .ZN(n7531) );
  NAND3_X1 U9306 ( .A1(n7532), .A2(n9981), .A3(n7531), .ZN(n7534) );
  AOI22_X1 U9307 ( .A1(n9986), .A2(n8287), .B1(n8286), .B2(n9983), .ZN(n7533)
         );
  NAND2_X1 U9308 ( .A1(n7534), .A2(n7533), .ZN(n7589) );
  AOI21_X1 U9309 ( .B1(n8554), .B2(n7641), .A(n7589), .ZN(n7540) );
  XNOR2_X1 U9310 ( .A(n7535), .B(n7836), .ZN(n7591) );
  INV_X1 U9311 ( .A(n7646), .ZN(n7537) );
  OAI22_X1 U9312 ( .A1(n7537), .A2(n9975), .B1(n7536), .B2(n9999), .ZN(n7538)
         );
  AOI21_X1 U9313 ( .B1(n7591), .B2(n9977), .A(n7538), .ZN(n7539) );
  OAI21_X1 U9314 ( .B1(n7540), .B2(n5088), .A(n7539), .ZN(P2_U3222) );
  INV_X1 U9315 ( .A(n7541), .ZN(n7542) );
  NAND2_X1 U9316 ( .A1(n8273), .A2(n7542), .ZN(n7545) );
  AOI21_X1 U9317 ( .B1(n8269), .B2(n8288), .A(n7543), .ZN(n7544) );
  OAI211_X1 U9318 ( .C1(n7644), .C2(n8271), .A(n7545), .B(n7544), .ZN(n7557)
         );
  XNOR2_X1 U9319 ( .A(n4514), .B(n10039), .ZN(n7617) );
  XNOR2_X1 U9320 ( .A(n7617), .B(n7616), .ZN(n7555) );
  INV_X1 U9321 ( .A(n7546), .ZN(n7548) );
  NAND2_X1 U9322 ( .A1(n7548), .A2(n7547), .ZN(n7549) );
  NAND2_X1 U9323 ( .A1(n7550), .A2(n7549), .ZN(n7554) );
  INV_X1 U9324 ( .A(n7554), .ZN(n7552) );
  INV_X1 U9325 ( .A(n7619), .ZN(n7553) );
  AOI211_X1 U9326 ( .C1(n7555), .C2(n7554), .A(n8264), .B(n7553), .ZN(n7556)
         );
  AOI211_X1 U9327 ( .C1(n10039), .C2(n8236), .A(n7557), .B(n7556), .ZN(n7558)
         );
  INV_X1 U9328 ( .A(n7558), .ZN(P2_U3171) );
  INV_X1 U9329 ( .A(n7559), .ZN(n7560) );
  NAND2_X1 U9330 ( .A1(n7561), .A2(n7560), .ZN(n7564) );
  NAND2_X1 U9331 ( .A1(n5099), .A2(n7562), .ZN(n7563) );
  XNOR2_X1 U9332 ( .A(n7564), .B(n7563), .ZN(n7572) );
  NAND2_X1 U9333 ( .A1(n8832), .A2(n9145), .ZN(n7566) );
  OAI211_X1 U9334 ( .C1(n9027), .C2(n8834), .A(n7566), .B(n7565), .ZN(n7567)
         );
  AOI21_X1 U9335 ( .B1(n7568), .B2(n8837), .A(n7567), .ZN(n7571) );
  NAND2_X1 U9336 ( .A1(n8821), .A2(n7569), .ZN(n7570) );
  OAI211_X1 U9337 ( .C1(n7572), .C2(n8823), .A(n7571), .B(n7570), .ZN(P1_U3236) );
  XOR2_X1 U9338 ( .A(n7573), .B(n7574), .Z(n7582) );
  NAND2_X1 U9339 ( .A1(n8832), .A2(n9143), .ZN(n7576) );
  OAI211_X1 U9340 ( .C1(n7577), .C2(n8834), .A(n7576), .B(n7575), .ZN(n7579)
         );
  NOR2_X1 U9341 ( .A1(n9821), .A2(n8840), .ZN(n7578) );
  AOI211_X1 U9342 ( .C1(n8837), .C2(n7580), .A(n7579), .B(n7578), .ZN(n7581)
         );
  OAI21_X1 U9343 ( .B1(n7582), .B2(n8823), .A(n7581), .ZN(P1_U3234) );
  INV_X1 U9344 ( .A(n7583), .ZN(n7595) );
  OAI222_X1 U9345 ( .A1(n8729), .A2(n7595), .B1(P2_U3151), .B2(n7585), .C1(
        n7584), .C2(n8723), .ZN(P2_U3271) );
  MUX2_X1 U9346 ( .A(n7589), .B(P2_REG0_REG_11__SCAN_IN), .S(n10049), .Z(n7586) );
  INV_X1 U9347 ( .A(n7586), .ZN(n7588) );
  INV_X1 U9348 ( .A(n8712), .ZN(n8718) );
  AOI22_X1 U9349 ( .A1(n7591), .A2(n8718), .B1(n8717), .B2(n7646), .ZN(n7587)
         );
  NAND2_X1 U9350 ( .A1(n7588), .A2(n7587), .ZN(P2_U3423) );
  MUX2_X1 U9351 ( .A(n7589), .B(P2_REG1_REG_11__SCAN_IN), .S(n10062), .Z(n7590) );
  INV_X1 U9352 ( .A(n7590), .ZN(n7593) );
  INV_X1 U9353 ( .A(n8626), .ZN(n8630) );
  AOI22_X1 U9354 ( .A1(n7591), .A2(n8630), .B1(n8629), .B2(n7646), .ZN(n7592)
         );
  NAND2_X1 U9355 ( .A1(n7593), .A2(n7592), .ZN(P2_U3470) );
  OAI222_X1 U9356 ( .A1(n7596), .A2(P1_U3086), .B1(n9634), .B2(n7595), .C1(
        n7594), .C2(n9632), .ZN(P1_U3331) );
  INV_X1 U9357 ( .A(n7600), .ZN(n7597) );
  INV_X1 U9358 ( .A(n9046), .ZN(n7598) );
  INV_X1 U9359 ( .A(n9140), .ZN(n7758) );
  OR2_X1 U9360 ( .A1(n8769), .A2(n7758), .ZN(n9050) );
  NAND2_X1 U9361 ( .A1(n8769), .A2(n7758), .ZN(n9048) );
  OAI21_X1 U9362 ( .B1(n7597), .B2(n7598), .A(n7611), .ZN(n7601) );
  NOR2_X1 U9363 ( .A1(n7611), .A2(n7598), .ZN(n7599) );
  NAND2_X1 U9364 ( .A1(n7600), .A2(n7599), .ZN(n7687) );
  NAND2_X1 U9365 ( .A1(n7601), .A2(n7687), .ZN(n7602) );
  AOI222_X1 U9366 ( .A1(n9491), .A2(n7602), .B1(n9139), .B2(n9708), .C1(n5016), 
        .C2(n9711), .ZN(n9644) );
  INV_X1 U9367 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7603) );
  OAI22_X1 U9368 ( .A1(n9534), .A2(n7603), .B1(n8765), .B2(n9522), .ZN(n7607)
         );
  INV_X1 U9369 ( .A(n8769), .ZN(n9645) );
  OAI211_X1 U9370 ( .C1(n9645), .C2(n7605), .A(n9722), .B(n7692), .ZN(n9643)
         );
  NOR2_X1 U9371 ( .A1(n9643), .A2(n9484), .ZN(n7606) );
  AOI211_X1 U9372 ( .C1(n9719), .C2(n8769), .A(n7607), .B(n7606), .ZN(n7615)
         );
  AND2_X1 U9373 ( .A1(n7610), .A2(n8898), .ZN(n9642) );
  INV_X1 U9374 ( .A(n9642), .ZN(n7613) );
  INV_X1 U9375 ( .A(n7610), .ZN(n7612) );
  NAND3_X1 U9376 ( .A1(n7613), .A2(n9647), .A3(n9486), .ZN(n7614) );
  OAI211_X1 U9377 ( .C1(n9644), .C2(n9730), .A(n7615), .B(n7614), .ZN(P1_U3277) );
  OR2_X1 U9378 ( .A1(n7617), .A2(n7616), .ZN(n7618) );
  XNOR2_X1 U9379 ( .A(n7620), .B(n4511), .ZN(n7621) );
  NAND2_X1 U9380 ( .A1(n7622), .A2(n7621), .ZN(n7638) );
  OAI21_X1 U9381 ( .B1(n7622), .B2(n7621), .A(n7638), .ZN(n7632) );
  NOR2_X1 U9382 ( .A1(n8276), .A2(n10043), .ZN(n7631) );
  INV_X1 U9383 ( .A(n7623), .ZN(n7624) );
  NAND2_X1 U9384 ( .A1(n8273), .A2(n7624), .ZN(n7628) );
  AOI21_X1 U9385 ( .B1(n8269), .B2(n7626), .A(n7625), .ZN(n7627) );
  OAI211_X1 U9386 ( .C1(n7629), .C2(n8271), .A(n7628), .B(n7627), .ZN(n7630)
         );
  AOI211_X1 U9387 ( .C1(n7632), .C2(n8244), .A(n7631), .B(n7630), .ZN(n7633)
         );
  INV_X1 U9388 ( .A(n7633), .ZN(P2_U3157) );
  INV_X1 U9389 ( .A(n7634), .ZN(n7635) );
  NAND2_X1 U9390 ( .A1(n7635), .A2(n7644), .ZN(n7639) );
  XNOR2_X1 U9391 ( .A(n7636), .B(n8136), .ZN(n8046) );
  AND2_X1 U9392 ( .A1(n7639), .A2(n8046), .ZN(n7637) );
  NAND2_X1 U9393 ( .A1(n7638), .A2(n7637), .ZN(n8049) );
  NAND2_X1 U9394 ( .A1(n8049), .A2(n8244), .ZN(n7649) );
  AOI21_X1 U9395 ( .B1(n7638), .B2(n7639), .A(n8046), .ZN(n7648) );
  AOI21_X1 U9396 ( .B1(n8258), .B2(n8286), .A(n7640), .ZN(n7643) );
  NAND2_X1 U9397 ( .A1(n8273), .A2(n7641), .ZN(n7642) );
  OAI211_X1 U9398 ( .C1(n8256), .C2(n7644), .A(n7643), .B(n7642), .ZN(n7645)
         );
  AOI21_X1 U9399 ( .B1(n7646), .B2(n8236), .A(n7645), .ZN(n7647) );
  OAI21_X1 U9400 ( .B1(n7649), .B2(n7648), .A(n7647), .ZN(P2_U3176) );
  INV_X1 U9401 ( .A(n7650), .ZN(n7652) );
  NAND2_X1 U9402 ( .A1(n7652), .A2(n7651), .ZN(n7653) );
  XNOR2_X1 U9403 ( .A(n7654), .B(n7653), .ZN(n7667) );
  AOI21_X1 U9404 ( .B1(n4605), .B2(n7656), .A(n7655), .ZN(n7657) );
  NOR2_X1 U9405 ( .A1(n7657), .A2(n9948), .ZN(n7666) );
  AOI21_X1 U9406 ( .B1(n4596), .B2(n7659), .A(n7658), .ZN(n7664) );
  NOR2_X1 U9407 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7660), .ZN(n8161) );
  INV_X1 U9408 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10099) );
  NOR2_X1 U9409 ( .A1(n9969), .A2(n10099), .ZN(n7661) );
  AOI211_X1 U9410 ( .C1(n7662), .C2(n9915), .A(n8161), .B(n7661), .ZN(n7663)
         );
  OAI21_X1 U9411 ( .B1(n7664), .B2(n9953), .A(n7663), .ZN(n7665) );
  AOI211_X1 U9412 ( .C1(n7667), .C2(n9964), .A(n7666), .B(n7665), .ZN(n7668)
         );
  INV_X1 U9413 ( .A(n7668), .ZN(P2_U3194) );
  XNOR2_X1 U9414 ( .A(n7669), .B(n7838), .ZN(n7683) );
  INV_X1 U9415 ( .A(n7838), .ZN(n7918) );
  XNOR2_X1 U9416 ( .A(n7670), .B(n7918), .ZN(n7671) );
  AOI222_X1 U9417 ( .A1(n9981), .A2(n7671), .B1(n8285), .B2(n9983), .C1(n8162), 
        .C2(n9986), .ZN(n7679) );
  MUX2_X1 U9418 ( .A(n7672), .B(n7679), .S(n10048), .Z(n7674) );
  NAND2_X1 U9419 ( .A1(n8717), .A2(n8166), .ZN(n7673) );
  OAI211_X1 U9420 ( .C1(n7683), .C2(n8712), .A(n7674), .B(n7673), .ZN(P2_U3426) );
  MUX2_X1 U9421 ( .A(n7675), .B(n7679), .S(n9999), .Z(n7678) );
  INV_X1 U9422 ( .A(n8164), .ZN(n7676) );
  AOI22_X1 U9423 ( .A1(n8166), .A2(n8555), .B1(n8554), .B2(n7676), .ZN(n7677)
         );
  OAI211_X1 U9424 ( .C1(n7683), .C2(n8558), .A(n7678), .B(n7677), .ZN(P2_U3221) );
  MUX2_X1 U9425 ( .A(n7680), .B(n7679), .S(n10064), .Z(n7682) );
  NAND2_X1 U9426 ( .A1(n8166), .A2(n8629), .ZN(n7681) );
  OAI211_X1 U9427 ( .C1(n7683), .C2(n8626), .A(n7682), .B(n7681), .ZN(P2_U3471) );
  INV_X1 U9428 ( .A(n7684), .ZN(n7730) );
  OAI222_X1 U9429 ( .A1(n8729), .A2(n7730), .B1(P2_U3151), .B2(n7686), .C1(
        n7685), .C2(n8039), .ZN(P2_U3270) );
  OR2_X1 U9430 ( .A1(n8778), .A2(n5025), .ZN(n8938) );
  NAND2_X1 U9431 ( .A1(n8778), .A2(n5025), .ZN(n8940) );
  XNOR2_X1 U9432 ( .A(n7742), .B(n8900), .ZN(n7690) );
  NAND2_X1 U9433 ( .A1(n9138), .A2(n9708), .ZN(n7688) );
  OAI21_X1 U9434 ( .B1(n7758), .B2(n9691), .A(n7688), .ZN(n7689) );
  AOI21_X1 U9435 ( .B1(n7690), .B2(n9491), .A(n7689), .ZN(n9638) );
  NAND2_X1 U9436 ( .A1(n8769), .A2(n9140), .ZN(n7691) );
  XNOR2_X1 U9437 ( .A(n7737), .B(n8900), .ZN(n9641) );
  NAND2_X1 U9438 ( .A1(n9641), .A2(n9486), .ZN(n7697) );
  INV_X1 U9439 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9321) );
  OAI22_X1 U9440 ( .A1(n9534), .A2(n9321), .B1(n8774), .B2(n9522), .ZN(n7695)
         );
  INV_X1 U9441 ( .A(n7692), .ZN(n7693) );
  INV_X1 U9442 ( .A(n8778), .ZN(n9639) );
  OAI211_X1 U9443 ( .C1(n7693), .C2(n9639), .A(n9722), .B(n4592), .ZN(n9637)
         );
  NOR2_X1 U9444 ( .A1(n9637), .A2(n9484), .ZN(n7694) );
  AOI211_X1 U9445 ( .C1(n9719), .C2(n8778), .A(n7695), .B(n7694), .ZN(n7696)
         );
  OAI211_X1 U9446 ( .C1(n9730), .C2(n9638), .A(n7697), .B(n7696), .ZN(P1_U3276) );
  INV_X1 U9447 ( .A(n7698), .ZN(n7711) );
  OAI222_X1 U9448 ( .A1(n8729), .A2(n7711), .B1(P2_U3151), .B2(n7700), .C1(
        n7699), .C2(n8039), .ZN(P2_U3269) );
  NAND2_X1 U9449 ( .A1(n7702), .A2(n7701), .ZN(n7703) );
  XOR2_X1 U9450 ( .A(n7704), .B(n7703), .Z(n7709) );
  NAND2_X1 U9451 ( .A1(n8837), .A2(n9697), .ZN(n7706) );
  AND2_X1 U9452 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9251) );
  AOI21_X1 U9453 ( .B1(n8796), .B2(n5016), .A(n9251), .ZN(n7705) );
  OAI211_X1 U9454 ( .C1(n8798), .C2(n9692), .A(n7706), .B(n7705), .ZN(n7707)
         );
  AOI21_X1 U9455 ( .B1(n9699), .B2(n8821), .A(n7707), .ZN(n7708) );
  OAI21_X1 U9456 ( .B1(n7709), .B2(n8823), .A(n7708), .ZN(P1_U3215) );
  OAI222_X1 U9457 ( .A1(n7712), .A2(P1_U3086), .B1(n9634), .B2(n7711), .C1(
        n7710), .C2(n9632), .ZN(P1_U3329) );
  INV_X1 U9458 ( .A(n7922), .ZN(n7714) );
  AND2_X1 U9459 ( .A1(n7714), .A2(n7713), .ZN(n7839) );
  XOR2_X1 U9460 ( .A(n7839), .B(n7715), .Z(n7716) );
  AOI222_X1 U9461 ( .A1(n9981), .A2(n7716), .B1(n8548), .B2(n9983), .C1(n8286), 
        .C2(n9986), .ZN(n7725) );
  INV_X1 U9462 ( .A(n7725), .ZN(n7718) );
  OAI22_X1 U9463 ( .A1(n7925), .A2(n8443), .B1(n8226), .B2(n9990), .ZN(n7717)
         );
  OAI21_X1 U9464 ( .B1(n7718), .B2(n7717), .A(n9999), .ZN(n7721) );
  XNOR2_X1 U9465 ( .A(n7719), .B(n7839), .ZN(n7726) );
  AOI22_X1 U9466 ( .A1(n7726), .A2(n9977), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n5088), .ZN(n7720) );
  NAND2_X1 U9467 ( .A1(n7721), .A2(n7720), .ZN(P2_U3220) );
  INV_X1 U9468 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7722) );
  MUX2_X1 U9469 ( .A(n7722), .B(n7725), .S(n10048), .Z(n7724) );
  AOI22_X1 U9470 ( .A1(n7726), .A2(n8718), .B1(n8717), .B2(n8228), .ZN(n7723)
         );
  NAND2_X1 U9471 ( .A1(n7724), .A2(n7723), .ZN(P2_U3429) );
  MUX2_X1 U9472 ( .A(n8302), .B(n7725), .S(n10064), .Z(n7728) );
  AOI22_X1 U9473 ( .A1(n7726), .A2(n8630), .B1(n8629), .B2(n8228), .ZN(n7727)
         );
  NAND2_X1 U9474 ( .A1(n7728), .A2(n7727), .ZN(P2_U3472) );
  OAI222_X1 U9475 ( .A1(n6506), .A2(P1_U3086), .B1(n9634), .B2(n7730), .C1(
        n7729), .C2(n9632), .ZN(P1_U3330) );
  INV_X1 U9476 ( .A(n7731), .ZN(n7750) );
  OAI222_X1 U9477 ( .A1(n8729), .A2(n7750), .B1(n5315), .B2(P2_U3151), .C1(
        n7732), .C2(n8039), .ZN(P2_U3268) );
  NAND2_X1 U9478 ( .A1(n7791), .A2(n7733), .ZN(n7735) );
  OAI211_X1 U9479 ( .C1(n7736), .C2(n8723), .A(n7735), .B(n7734), .ZN(P2_U3267) );
  INV_X1 U9480 ( .A(n9138), .ZN(n9533) );
  OR2_X1 U9481 ( .A1(n9608), .A2(n9533), .ZN(n9527) );
  NAND2_X1 U9482 ( .A1(n9608), .A2(n9533), .ZN(n9057) );
  NAND2_X1 U9483 ( .A1(n9527), .A2(n9057), .ZN(n8902) );
  XNOR2_X1 U9484 ( .A(n7764), .B(n7744), .ZN(n9610) );
  INV_X1 U9485 ( .A(n9520), .ZN(n7739) );
  AOI211_X1 U9486 ( .C1(n9608), .C2(n4592), .A(n9541), .B(n7739), .ZN(n9606)
         );
  NOR2_X1 U9487 ( .A1(n7738), .A2(n9521), .ZN(n7741) );
  OAI22_X1 U9488 ( .A1(n9534), .A2(n9324), .B1(n8816), .B2(n9522), .ZN(n7740)
         );
  AOI211_X1 U9489 ( .C1(n9606), .C2(n9726), .A(n7741), .B(n7740), .ZN(n7748)
         );
  INV_X1 U9490 ( .A(n8900), .ZN(n9054) );
  OAI211_X1 U9491 ( .C1(n7744), .C2(n7743), .A(n9528), .B(n9491), .ZN(n7746)
         );
  AOI22_X1 U9492 ( .A1(n9137), .A2(n9708), .B1(n9711), .B2(n9139), .ZN(n7745)
         );
  NAND2_X1 U9493 ( .A1(n7746), .A2(n7745), .ZN(n9607) );
  NAND2_X1 U9494 ( .A1(n9607), .A2(n9534), .ZN(n7747) );
  OAI211_X1 U9495 ( .C1(n9610), .C2(n9537), .A(n7748), .B(n7747), .ZN(P1_U3275) );
  OAI222_X1 U9496 ( .A1(P1_U3086), .A2(n4522), .B1(n9634), .B2(n7750), .C1(
        n7749), .C2(n9632), .ZN(P1_U3328) );
  INV_X1 U9497 ( .A(n7751), .ZN(n7755) );
  OAI21_X1 U9498 ( .B1(n7753), .B2(n7755), .A(n7752), .ZN(n7754) );
  OAI211_X1 U9499 ( .C1(n7756), .C2(n7755), .A(n7754), .B(n8830), .ZN(n7762)
         );
  NAND2_X1 U9500 ( .A1(n8832), .A2(n9141), .ZN(n7757) );
  NAND2_X1 U9501 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9274) );
  OAI211_X1 U9502 ( .C1(n7758), .C2(n8834), .A(n7757), .B(n9274), .ZN(n7759)
         );
  AOI21_X1 U9503 ( .B1(n7760), .B2(n8837), .A(n7759), .ZN(n7761) );
  OAI211_X1 U9504 ( .C1(n7480), .C2(n8840), .A(n7762), .B(n7761), .ZN(P1_U3241) );
  INV_X1 U9505 ( .A(n9570), .ZN(n9430) );
  INV_X1 U9506 ( .A(n8757), .ZN(n9461) );
  NOR2_X1 U9507 ( .A1(n9608), .A2(n9138), .ZN(n7763) );
  NAND2_X1 U9508 ( .A1(n9608), .A2(n9138), .ZN(n7765) );
  OR2_X1 U9509 ( .A1(n9603), .A2(n9137), .ZN(n7766) );
  AND2_X1 U9510 ( .A1(n9515), .A2(n9532), .ZN(n7767) );
  AND2_X1 U9511 ( .A1(n9593), .A2(n9471), .ZN(n7769) );
  OR2_X1 U9512 ( .A1(n9593), .A2(n9471), .ZN(n7768) );
  XNOR2_X1 U9513 ( .A(n9584), .B(n9462), .ZN(n9474) );
  NAND2_X1 U9514 ( .A1(n9565), .A2(n8756), .ZN(n9096) );
  NAND2_X1 U9515 ( .A1(n9099), .A2(n9096), .ZN(n9410) );
  NAND2_X1 U9516 ( .A1(n9560), .A2(n8835), .ZN(n8858) );
  NAND2_X1 U9517 ( .A1(n9104), .A2(n8858), .ZN(n9401) );
  NAND2_X1 U9518 ( .A1(n9402), .A2(n9401), .ZN(n9400) );
  NAND2_X1 U9519 ( .A1(n9554), .A2(n9379), .ZN(n9371) );
  NAND2_X1 U9520 ( .A1(n9103), .A2(n9371), .ZN(n8907) );
  INV_X1 U9521 ( .A(n8907), .ZN(n7779) );
  XNOR2_X1 U9522 ( .A(n9382), .B(n7779), .ZN(n9557) );
  NAND2_X1 U9523 ( .A1(n9515), .A2(n9519), .ZN(n9509) );
  INV_X1 U9524 ( .A(n9403), .ZN(n7772) );
  INV_X1 U9525 ( .A(n9385), .ZN(n7771) );
  AOI211_X1 U9526 ( .C1(n9554), .C2(n7772), .A(n9541), .B(n7771), .ZN(n9553)
         );
  AOI22_X1 U9527 ( .A1(n9730), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n7773), .B2(
        n9718), .ZN(n7774) );
  OAI21_X1 U9528 ( .B1(n9380), .B2(n9521), .A(n7774), .ZN(n7780) );
  NAND2_X1 U9529 ( .A1(n9575), .A2(n8757), .ZN(n9090) );
  NAND2_X1 U9530 ( .A1(n9091), .A2(n9090), .ZN(n9448) );
  NAND2_X1 U9531 ( .A1(n9580), .A2(n8809), .ZN(n9446) );
  INV_X1 U9532 ( .A(n9446), .ZN(n9085) );
  NOR2_X1 U9533 ( .A1(n9448), .A2(n9085), .ZN(n7777) );
  INV_X1 U9534 ( .A(n9532), .ZN(n9136) );
  NAND2_X1 U9535 ( .A1(n9515), .A2(n9136), .ZN(n8969) );
  INV_X1 U9536 ( .A(n9137), .ZN(n9507) );
  OR2_X1 U9537 ( .A1(n9603), .A2(n9507), .ZN(n9066) );
  AND2_X1 U9538 ( .A1(n9066), .A2(n9527), .ZN(n9062) );
  NAND2_X1 U9539 ( .A1(n9528), .A2(n9062), .ZN(n7775) );
  NAND2_X1 U9540 ( .A1(n9603), .A2(n9507), .ZN(n9058) );
  INV_X1 U9541 ( .A(n8967), .ZN(n9067) );
  INV_X1 U9542 ( .A(n9471), .ZN(n9508) );
  OR2_X1 U9543 ( .A1(n9593), .A2(n9508), .ZN(n9081) );
  NAND2_X1 U9544 ( .A1(n9593), .A2(n9508), .ZN(n9072) );
  NAND2_X1 U9545 ( .A1(n9081), .A2(n9072), .ZN(n9492) );
  NAND2_X1 U9546 ( .A1(n9468), .A2(n9474), .ZN(n9467) );
  INV_X1 U9547 ( .A(n9462), .ZN(n9495) );
  NAND2_X1 U9548 ( .A1(n9584), .A2(n9495), .ZN(n8851) );
  OR2_X1 U9549 ( .A1(n9580), .A2(n8809), .ZN(n9087) );
  INV_X1 U9550 ( .A(n9091), .ZN(n7776) );
  OR2_X1 U9551 ( .A1(n9570), .A2(n8787), .ZN(n9098) );
  NAND2_X1 U9552 ( .A1(n9570), .A2(n8787), .ZN(n9095) );
  NAND2_X1 U9553 ( .A1(n9098), .A2(n9095), .ZN(n9425) );
  INV_X1 U9554 ( .A(n9425), .ZN(n9433) );
  NAND2_X1 U9555 ( .A1(n9431), .A2(n9095), .ZN(n9418) );
  INV_X1 U9556 ( .A(n9410), .ZN(n9419) );
  NAND2_X1 U9557 ( .A1(n9418), .A2(n9419), .ZN(n9417) );
  NAND2_X1 U9558 ( .A1(n9417), .A2(n9096), .ZN(n9396) );
  INV_X1 U9559 ( .A(n9401), .ZN(n9397) );
  NAND2_X1 U9560 ( .A1(n9396), .A2(n9397), .ZN(n9395) );
  NAND2_X1 U9561 ( .A1(n9395), .A2(n8858), .ZN(n7778) );
  NAND2_X1 U9562 ( .A1(n7778), .A2(n7779), .ZN(n9372) );
  OAI21_X1 U9563 ( .B1(n9557), .B2(n9537), .A(n7781), .ZN(P1_U3265) );
  INV_X1 U9564 ( .A(SI_29_), .ZN(n10227) );
  INV_X1 U9565 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10253) );
  INV_X1 U9566 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8045) );
  MUX2_X1 U9567 ( .A(n10253), .B(n8045), .S(n7798), .Z(n7787) );
  INV_X1 U9568 ( .A(SI_30_), .ZN(n7786) );
  NAND2_X1 U9569 ( .A1(n7787), .A2(n7786), .ZN(n7795) );
  INV_X1 U9570 ( .A(n7787), .ZN(n7788) );
  NAND2_X1 U9571 ( .A1(n7788), .A2(SI_30_), .ZN(n7789) );
  NAND2_X1 U9572 ( .A1(n7795), .A2(n7789), .ZN(n7796) );
  INV_X1 U9573 ( .A(n8842), .ZN(n8044) );
  INV_X1 U9574 ( .A(n7791), .ZN(n7792) );
  INV_X1 U9575 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10425) );
  OAI222_X1 U9576 ( .A1(P1_U3086), .A2(n7793), .B1(n9634), .B2(n7792), .C1(
        n10425), .C2(n9632), .ZN(P1_U3327) );
  NOR2_X1 U9577 ( .A1(n7803), .A2(n8045), .ZN(n7794) );
  OAI21_X1 U9578 ( .B1(n7797), .B2(n7796), .A(n7795), .ZN(n7802) );
  MUX2_X1 U9579 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7798), .Z(n7800) );
  INV_X1 U9580 ( .A(SI_31_), .ZN(n7799) );
  XNOR2_X1 U9581 ( .A(n7800), .B(n7799), .ZN(n7801) );
  XNOR2_X1 U9582 ( .A(n7802), .B(n7801), .ZN(n8874) );
  NAND2_X1 U9583 ( .A1(n8874), .A2(n5535), .ZN(n7805) );
  INV_X1 U9584 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8724) );
  OR2_X1 U9585 ( .A1(n7803), .A2(n8724), .ZN(n7804) );
  OAI22_X1 U9586 ( .A1(n7806), .A2(n8005), .B1(n8580), .B2(n8633), .ZN(n7818)
         );
  INV_X1 U9587 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7810) );
  NAND2_X1 U9588 ( .A1(n5401), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7809) );
  INV_X1 U9589 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8403) );
  OR2_X1 U9590 ( .A1(n7807), .A2(n8403), .ZN(n7808) );
  OAI211_X1 U9591 ( .C1(n7811), .C2(n7810), .A(n7809), .B(n7808), .ZN(n7812)
         );
  INV_X1 U9592 ( .A(n7812), .ZN(n7813) );
  INV_X1 U9593 ( .A(n8580), .ZN(n8637) );
  INV_X1 U9594 ( .A(n8279), .ZN(n7815) );
  NAND2_X1 U9595 ( .A1(n8016), .A2(n8001), .ZN(n7847) );
  INV_X1 U9596 ( .A(n8633), .ZN(n8577) );
  NOR2_X1 U9597 ( .A1(n8010), .A2(n8278), .ZN(n7817) );
  OAI22_X1 U9598 ( .A1(n7818), .A2(n7847), .B1(n8577), .B2(n7817), .ZN(n7849)
         );
  AND2_X1 U9599 ( .A1(n8633), .A2(n8278), .ZN(n8013) );
  INV_X1 U9600 ( .A(n7821), .ZN(n8449) );
  NAND2_X1 U9601 ( .A1(n7980), .A2(n7983), .ZN(n8452) );
  INV_X1 U9602 ( .A(n8489), .ZN(n8494) );
  INV_X1 U9603 ( .A(n8481), .ZN(n8476) );
  NAND2_X1 U9604 ( .A1(n8501), .A2(n7822), .ZN(n7951) );
  NAND2_X1 U9605 ( .A1(n7949), .A2(n7823), .ZN(n7945) );
  INV_X1 U9606 ( .A(n8545), .ZN(n8546) );
  NAND2_X1 U9607 ( .A1(n7928), .A2(n7932), .ZN(n8567) );
  NOR4_X1 U9608 ( .A1(n7826), .A2(n4612), .A3(n7825), .A4(n7824), .ZN(n7828)
         );
  NAND3_X1 U9609 ( .A1(n7828), .A2(n7827), .A3(n9974), .ZN(n7832) );
  NOR4_X1 U9610 ( .A1(n7832), .A2(n7831), .A3(n7830), .A4(n7829), .ZN(n7833)
         );
  NAND4_X1 U9611 ( .A1(n7836), .A2(n7835), .A3(n7834), .A4(n7833), .ZN(n7837)
         );
  NOR4_X1 U9612 ( .A1(n8567), .A2(n7839), .A3(n7838), .A4(n7837), .ZN(n7840)
         );
  NAND3_X1 U9613 ( .A1(n8535), .A2(n8546), .A3(n7840), .ZN(n7841) );
  NOR4_X1 U9614 ( .A1(n7842), .A2(n7951), .A3(n7945), .A4(n7841), .ZN(n7843)
         );
  NAND4_X1 U9615 ( .A1(n8468), .A2(n8494), .A3(n8476), .A4(n7843), .ZN(n7844)
         );
  NOR4_X1 U9616 ( .A1(n8439), .A2(n8458), .A3(n8452), .A4(n7844), .ZN(n7845)
         );
  NAND4_X1 U9617 ( .A1(n5839), .A2(n7977), .A3(n7845), .A4(n8406), .ZN(n7846)
         );
  XNOR2_X1 U9618 ( .A(n7851), .B(n7850), .ZN(n8024) );
  NAND2_X1 U9619 ( .A1(n7854), .A2(n7853), .ZN(n7855) );
  NAND2_X1 U9620 ( .A1(n7855), .A2(n7858), .ZN(n7861) );
  NAND2_X1 U9621 ( .A1(n7857), .A2(n7856), .ZN(n7860) );
  INV_X1 U9622 ( .A(n7858), .ZN(n7859) );
  AOI21_X1 U9623 ( .B1(n7861), .B2(n7860), .A(n7859), .ZN(n7862) );
  MUX2_X1 U9624 ( .A(n7862), .B(n7861), .S(n8012), .Z(n7869) );
  NAND2_X1 U9625 ( .A1(n7863), .A2(n7870), .ZN(n7866) );
  NAND2_X1 U9626 ( .A1(n9984), .A2(n10011), .ZN(n7871) );
  NAND2_X1 U9627 ( .A1(n7864), .A2(n7871), .ZN(n7865) );
  MUX2_X1 U9628 ( .A(n7866), .B(n7865), .S(n8012), .Z(n7867) );
  INV_X1 U9629 ( .A(n7867), .ZN(n7868) );
  OAI21_X1 U9630 ( .B1(n7869), .B2(n4612), .A(n7868), .ZN(n7876) );
  NAND2_X1 U9631 ( .A1(n7870), .A2(n8012), .ZN(n7873) );
  NAND3_X1 U9632 ( .A1(n7879), .A2(n7871), .A3(n8009), .ZN(n7872) );
  OAI22_X1 U9633 ( .A1(n7873), .A2(n7889), .B1(n7872), .B2(n7881), .ZN(n7874)
         );
  NAND3_X1 U9634 ( .A1(n7876), .A2(n7875), .A3(n7874), .ZN(n7897) );
  AOI21_X1 U9635 ( .B1(n7879), .B2(n7877), .A(n8009), .ZN(n7878) );
  INV_X1 U9636 ( .A(n7878), .ZN(n7885) );
  NAND2_X1 U9637 ( .A1(n7881), .A2(n8012), .ZN(n7884) );
  NAND2_X1 U9638 ( .A1(n7879), .A2(n8009), .ZN(n7880) );
  OR2_X1 U9639 ( .A1(n7881), .A2(n7880), .ZN(n7883) );
  NAND4_X1 U9640 ( .A1(n7885), .A2(n7884), .A3(n7883), .A4(n7882), .ZN(n7894)
         );
  AND2_X1 U9641 ( .A1(n7903), .A2(n7886), .ZN(n7888) );
  INV_X1 U9642 ( .A(n7888), .ZN(n7901) );
  NAND4_X1 U9643 ( .A1(n7888), .A2(n8012), .A3(n7887), .A4(n7889), .ZN(n7893)
         );
  INV_X1 U9644 ( .A(n7889), .ZN(n7891) );
  NAND3_X1 U9645 ( .A1(n7891), .A2(n8009), .A3(n7890), .ZN(n7892) );
  OAI211_X1 U9646 ( .C1(n7894), .C2(n7901), .A(n7893), .B(n7892), .ZN(n7895)
         );
  NAND4_X1 U9647 ( .A1(n7897), .A2(n7902), .A3(n7896), .A4(n7895), .ZN(n7907)
         );
  NAND2_X1 U9648 ( .A1(n7907), .A2(n7906), .ZN(n7912) );
  AND2_X1 U9649 ( .A1(n7913), .A2(n7908), .ZN(n7910) );
  INV_X1 U9650 ( .A(n7915), .ZN(n7909) );
  AOI21_X1 U9651 ( .B1(n7912), .B2(n7910), .A(n7909), .ZN(n7917) );
  NAND2_X1 U9652 ( .A1(n7912), .A2(n4630), .ZN(n7914) );
  NAND2_X1 U9653 ( .A1(n7914), .A2(n7913), .ZN(n7916) );
  NAND2_X1 U9654 ( .A1(n8166), .A2(n8050), .ZN(n7919) );
  MUX2_X1 U9655 ( .A(n7920), .B(n7919), .S(n8009), .Z(n7921) );
  NAND2_X1 U9656 ( .A1(n7923), .A2(n7922), .ZN(n7931) );
  NAND2_X1 U9657 ( .A1(n7931), .A2(n8012), .ZN(n7927) );
  INV_X1 U9658 ( .A(n7923), .ZN(n7924) );
  NAND2_X1 U9659 ( .A1(n7924), .A2(n8562), .ZN(n7926) );
  MUX2_X1 U9660 ( .A(n7927), .B(n7926), .S(n7925), .Z(n7935) );
  NOR2_X1 U9661 ( .A1(n8567), .A2(n8562), .ZN(n7930) );
  NAND2_X1 U9662 ( .A1(n7936), .A2(n7928), .ZN(n7929) );
  AOI21_X1 U9663 ( .B1(n7931), .B2(n7930), .A(n7929), .ZN(n7933) );
  MUX2_X1 U9664 ( .A(n7933), .B(n7932), .S(n8012), .Z(n7934) );
  OAI21_X1 U9665 ( .B1(n7935), .B2(n8567), .A(n7934), .ZN(n7943) );
  INV_X1 U9666 ( .A(n7942), .ZN(n7937) );
  OAI211_X1 U9667 ( .C1(n7943), .C2(n7937), .A(n7940), .B(n7936), .ZN(n7938)
         );
  INV_X1 U9668 ( .A(n8523), .ZN(n8525) );
  NAND2_X1 U9669 ( .A1(n7940), .A2(n8009), .ZN(n7941) );
  AOI21_X1 U9670 ( .B1(n7943), .B2(n7942), .A(n7941), .ZN(n7944) );
  AOI21_X1 U9671 ( .B1(n7948), .B2(n8009), .A(n7944), .ZN(n7952) );
  INV_X1 U9672 ( .A(n7945), .ZN(n7947) );
  NAND2_X1 U9673 ( .A1(n7959), .A2(n8501), .ZN(n7946) );
  OAI21_X1 U9674 ( .B1(n7952), .B2(n7951), .A(n7950), .ZN(n7960) );
  NAND3_X1 U9675 ( .A1(n7960), .A2(n7958), .A3(n7961), .ZN(n7957) );
  AND2_X1 U9676 ( .A1(n7954), .A2(n7953), .ZN(n7956) );
  INV_X1 U9677 ( .A(n7962), .ZN(n7955) );
  AOI21_X1 U9678 ( .B1(n7957), .B2(n7956), .A(n7955), .ZN(n7967) );
  OAI211_X1 U9679 ( .C1(n7960), .C2(n4852), .A(n8494), .B(n7959), .ZN(n7965)
         );
  AND2_X1 U9680 ( .A1(n7962), .A2(n7961), .ZN(n7964) );
  AOI21_X1 U9681 ( .B1(n7965), .B2(n7964), .A(n7963), .ZN(n7966) );
  MUX2_X1 U9682 ( .A(n7969), .B(n7968), .S(n8012), .Z(n7970) );
  INV_X1 U9683 ( .A(n7970), .ZN(n7971) );
  NOR2_X1 U9684 ( .A1(n8458), .A2(n7971), .ZN(n7972) );
  INV_X1 U9685 ( .A(n7994), .ZN(n7976) );
  NOR2_X1 U9686 ( .A1(n7973), .A2(n8012), .ZN(n7974) );
  NAND4_X1 U9687 ( .A1(n7982), .A2(n7974), .A3(n7987), .A4(n7980), .ZN(n7975)
         );
  INV_X1 U9688 ( .A(n7984), .ZN(n7979) );
  NOR4_X1 U9689 ( .A1(n8423), .A2(n7979), .A3(n8009), .A4(n7978), .ZN(n7993)
         );
  INV_X1 U9690 ( .A(n8406), .ZN(n8408) );
  NAND2_X1 U9691 ( .A1(n7987), .A2(n7980), .ZN(n7981) );
  NAND3_X1 U9692 ( .A1(n7981), .A2(n8012), .A3(n7984), .ZN(n7991) );
  XNOR2_X1 U9693 ( .A(n7982), .B(n8009), .ZN(n7986) );
  NAND3_X1 U9694 ( .A1(n7984), .A2(n8009), .A3(n7983), .ZN(n7985) );
  OAI211_X1 U9695 ( .C1(n8012), .C2(n7987), .A(n7986), .B(n7985), .ZN(n7990)
         );
  NAND2_X1 U9696 ( .A1(n7988), .A2(n8009), .ZN(n7989) );
  OAI211_X1 U9697 ( .C1(n8423), .C2(n7991), .A(n7990), .B(n7989), .ZN(n7992)
         );
  NAND2_X1 U9698 ( .A1(n8642), .A2(n8426), .ZN(n7998) );
  INV_X1 U9699 ( .A(n7996), .ZN(n7997) );
  MUX2_X1 U9700 ( .A(n7998), .B(n7997), .S(n8009), .Z(n7999) );
  AND2_X1 U9701 ( .A1(n4704), .A2(n7999), .ZN(n8000) );
  MUX2_X1 U9702 ( .A(n8101), .B(n8007), .S(n8009), .Z(n8006) );
  MUX2_X1 U9703 ( .A(n8101), .B(n8007), .S(n8012), .Z(n8008) );
  AOI21_X1 U9704 ( .B1(n8012), .B2(n8011), .A(n8010), .ZN(n8014) );
  INV_X1 U9705 ( .A(n8016), .ZN(n8017) );
  NAND2_X1 U9706 ( .A1(n8022), .A2(n8019), .ZN(n8020) );
  OAI21_X1 U9707 ( .B1(n8022), .B2(n8021), .A(n8020), .ZN(n8023) );
  NOR3_X1 U9708 ( .A1(n8026), .A2(n8025), .A3(n5235), .ZN(n8029) );
  OAI21_X1 U9709 ( .B1(n8030), .B2(n8027), .A(P2_B_REG_SCAN_IN), .ZN(n8028) );
  OAI22_X1 U9710 ( .A1(n8031), .A2(n8030), .B1(n8029), .B2(n8028), .ZN(
        P2_U3296) );
  NOR2_X1 U9711 ( .A1(n8033), .A2(n9990), .ZN(n8401) );
  AOI21_X1 U9712 ( .B1(n5088), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8401), .ZN(
        n8034) );
  OAI21_X1 U9713 ( .B1(n8035), .B2(n9975), .A(n8034), .ZN(n8036) );
  AOI21_X1 U9714 ( .B1(n6583), .B2(n8037), .A(n8036), .ZN(n8038) );
  OAI21_X1 U9715 ( .B1(n8032), .B2(n5088), .A(n8038), .ZN(P2_U3204) );
  INV_X1 U9716 ( .A(n8864), .ZN(n9633) );
  OAI222_X1 U9717 ( .A1(n8729), .A2(n9633), .B1(n8041), .B2(P2_U3151), .C1(
        n8040), .C2(n8039), .ZN(P2_U3266) );
  OAI222_X1 U9718 ( .A1(n8723), .A2(n8045), .B1(n8729), .B2(n8044), .C1(
        P2_U3151), .C2(n8042), .ZN(P2_U3265) );
  XNOR2_X1 U9719 ( .A(n8584), .B(n4514), .ZN(n8253) );
  INV_X1 U9720 ( .A(n8046), .ZN(n8047) );
  NAND2_X1 U9721 ( .A1(n8047), .A2(n8162), .ZN(n8048) );
  XNOR2_X1 U9722 ( .A(n8166), .B(n8136), .ZN(n8051) );
  XNOR2_X1 U9723 ( .A(n8051), .B(n8050), .ZN(n8158) );
  NAND2_X1 U9724 ( .A1(n8051), .A2(n8286), .ZN(n8052) );
  XNOR2_X1 U9725 ( .A(n8228), .B(n4514), .ZN(n8054) );
  NAND2_X1 U9726 ( .A1(n8054), .A2(n8562), .ZN(n8107) );
  INV_X1 U9727 ( .A(n8054), .ZN(n8055) );
  NAND2_X1 U9728 ( .A1(n8055), .A2(n8285), .ZN(n8056) );
  NAND2_X1 U9729 ( .A1(n8107), .A2(n8056), .ZN(n8221) );
  XNOR2_X1 U9730 ( .A(n8716), .B(n8136), .ZN(n8058) );
  XNOR2_X1 U9731 ( .A(n8058), .B(n8223), .ZN(n8108) );
  INV_X1 U9732 ( .A(n8058), .ZN(n8059) );
  NAND2_X1 U9733 ( .A1(n8059), .A2(n8223), .ZN(n8060) );
  XNOR2_X1 U9734 ( .A(n8709), .B(n8136), .ZN(n8065) );
  XNOR2_X1 U9735 ( .A(n8065), .B(n8536), .ZN(n8265) );
  INV_X1 U9736 ( .A(n8265), .ZN(n8061) );
  XNOR2_X1 U9737 ( .A(n8703), .B(n4511), .ZN(n8062) );
  NAND2_X1 U9738 ( .A1(n8062), .A2(n8550), .ZN(n8188) );
  INV_X1 U9739 ( .A(n8062), .ZN(n8063) );
  INV_X1 U9740 ( .A(n8550), .ZN(n8527) );
  NAND2_X1 U9741 ( .A1(n8063), .A2(n8527), .ZN(n8064) );
  NAND2_X1 U9742 ( .A1(n8188), .A2(n8064), .ZN(n8179) );
  AND2_X1 U9743 ( .A1(n8065), .A2(n8536), .ZN(n8178) );
  NOR2_X1 U9744 ( .A1(n8179), .A2(n8178), .ZN(n8066) );
  NAND2_X1 U9745 ( .A1(n8176), .A2(n8188), .ZN(n8070) );
  XNOR2_X1 U9746 ( .A(n8697), .B(n4514), .ZN(n8067) );
  NAND2_X1 U9747 ( .A1(n8067), .A2(n8516), .ZN(n8240) );
  INV_X1 U9748 ( .A(n8067), .ZN(n8068) );
  NAND2_X1 U9749 ( .A1(n8068), .A2(n8537), .ZN(n8069) );
  AND2_X1 U9750 ( .A1(n8240), .A2(n8069), .ZN(n8189) );
  NAND2_X1 U9751 ( .A1(n8070), .A2(n8189), .ZN(n8192) );
  NAND2_X1 U9752 ( .A1(n8192), .A2(n8240), .ZN(n8075) );
  XNOR2_X1 U9753 ( .A(n8614), .B(n4511), .ZN(n8072) );
  NAND2_X1 U9754 ( .A1(n8072), .A2(n8071), .ZN(n8124) );
  INV_X1 U9755 ( .A(n8072), .ZN(n8073) );
  NAND2_X1 U9756 ( .A1(n8073), .A2(n8528), .ZN(n8074) );
  AND2_X1 U9757 ( .A1(n8124), .A2(n8074), .ZN(n8241) );
  XNOR2_X1 U9758 ( .A(n8687), .B(n4514), .ZN(n8076) );
  NAND2_X1 U9759 ( .A1(n8076), .A2(n8517), .ZN(n8212) );
  INV_X1 U9760 ( .A(n8076), .ZN(n8077) );
  NAND2_X1 U9761 ( .A1(n8077), .A2(n8284), .ZN(n8078) );
  AND2_X1 U9762 ( .A1(n8212), .A2(n8078), .ZN(n8125) );
  XNOR2_X1 U9763 ( .A(n8211), .B(n4511), .ZN(n8079) );
  NAND2_X1 U9764 ( .A1(n8079), .A2(n8479), .ZN(n8148) );
  INV_X1 U9765 ( .A(n8079), .ZN(n8080) );
  NAND2_X1 U9766 ( .A1(n8080), .A2(n8505), .ZN(n8081) );
  AND2_X1 U9767 ( .A1(n8148), .A2(n8081), .ZN(n8213) );
  NAND2_X1 U9768 ( .A1(n8147), .A2(n8148), .ZN(n8083) );
  XNOR2_X1 U9769 ( .A(n8082), .B(n8136), .ZN(n8084) );
  XNOR2_X1 U9770 ( .A(n8084), .B(n8493), .ZN(n8149) );
  INV_X1 U9771 ( .A(n8084), .ZN(n8085) );
  NAND2_X1 U9772 ( .A1(n8085), .A2(n8493), .ZN(n8086) );
  XNOR2_X1 U9773 ( .A(n8470), .B(n4514), .ZN(n8231) );
  INV_X1 U9774 ( .A(n8231), .ZN(n8088) );
  NAND2_X1 U9775 ( .A1(n8088), .A2(n8283), .ZN(n8090) );
  AND2_X1 U9776 ( .A1(n8231), .A2(n8480), .ZN(n8089) );
  XNOR2_X1 U9777 ( .A(n8590), .B(n8136), .ZN(n8203) );
  XNOR2_X1 U9778 ( .A(n8668), .B(n8136), .ZN(n8200) );
  INV_X1 U9779 ( .A(n8200), .ZN(n8091) );
  OAI22_X1 U9780 ( .A1(n8203), .A2(n8460), .B1(n8467), .B2(n8091), .ZN(n8095)
         );
  OAI21_X1 U9781 ( .B1(n8200), .B2(n8282), .A(n8281), .ZN(n8093) );
  NOR3_X1 U9782 ( .A1(n8200), .A2(n8281), .A3(n8282), .ZN(n8092) );
  AOI21_X1 U9783 ( .B1(n8203), .B2(n8093), .A(n8092), .ZN(n8094) );
  XNOR2_X1 U9784 ( .A(n8655), .B(n8136), .ZN(n8096) );
  XNOR2_X1 U9785 ( .A(n8096), .B(n8446), .ZN(n8170) );
  INV_X1 U9786 ( .A(n8096), .ZN(n8097) );
  XNOR2_X1 U9787 ( .A(n8642), .B(n8136), .ZN(n8133) );
  XNOR2_X1 U9788 ( .A(n8133), .B(n8426), .ZN(n8134) );
  XNOR2_X1 U9789 ( .A(n8135), .B(n8134), .ZN(n8105) );
  INV_X1 U9790 ( .A(n8417), .ZN(n8100) );
  OAI22_X1 U9791 ( .A1(n8100), .A2(n8247), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8099), .ZN(n8103) );
  OAI22_X1 U9792 ( .A1(n8101), .A2(n8271), .B1(n8435), .B2(n8256), .ZN(n8102)
         );
  AOI211_X1 U9793 ( .C1(n8642), .C2(n8236), .A(n8103), .B(n8102), .ZN(n8104)
         );
  OAI21_X1 U9794 ( .B1(n8105), .B2(n8264), .A(n8104), .ZN(P2_U3154) );
  INV_X1 U9795 ( .A(n8716), .ZN(n8117) );
  INV_X1 U9796 ( .A(n8106), .ZN(n8220) );
  INV_X1 U9797 ( .A(n8107), .ZN(n8109) );
  NOR3_X1 U9798 ( .A1(n8220), .A2(n8109), .A3(n8108), .ZN(n8112) );
  INV_X1 U9799 ( .A(n8110), .ZN(n8111) );
  OAI21_X1 U9800 ( .B1(n8112), .B2(n8111), .A(n8244), .ZN(n8116) );
  NAND2_X1 U9801 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8318) );
  OAI21_X1 U9802 ( .B1(n8271), .B2(n8564), .A(n8318), .ZN(n8114) );
  NOR2_X1 U9803 ( .A1(n8247), .A2(n8570), .ZN(n8113) );
  AOI211_X1 U9804 ( .C1(n8269), .C2(n8285), .A(n8114), .B(n8113), .ZN(n8115)
         );
  OAI211_X1 U9805 ( .C1(n8117), .C2(n8276), .A(n8116), .B(n8115), .ZN(P2_U3155) );
  XNOR2_X1 U9806 ( .A(n8201), .B(n8200), .ZN(n8202) );
  XNOR2_X1 U9807 ( .A(n8202), .B(n8467), .ZN(n8122) );
  AOI22_X1 U9808 ( .A1(n8283), .A2(n8269), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8119) );
  NAND2_X1 U9809 ( .A1(n8273), .A2(n8462), .ZN(n8118) );
  OAI211_X1 U9810 ( .C1(n8460), .C2(n8271), .A(n8119), .B(n8118), .ZN(n8120)
         );
  AOI21_X1 U9811 ( .B1(n8668), .B2(n8236), .A(n8120), .ZN(n8121) );
  OAI21_X1 U9812 ( .B1(n8122), .B2(n8264), .A(n8121), .ZN(P2_U3156) );
  INV_X1 U9813 ( .A(n8687), .ZN(n8132) );
  INV_X1 U9814 ( .A(n8123), .ZN(n8245) );
  NOR3_X1 U9815 ( .A1(n8245), .A2(n4952), .A3(n8125), .ZN(n8126) );
  OAI21_X1 U9816 ( .B1(n8126), .B2(n4541), .A(n8244), .ZN(n8131) );
  NAND2_X1 U9817 ( .A1(n8269), .A2(n8528), .ZN(n8128) );
  OAI211_X1 U9818 ( .C1(n8479), .C2(n8271), .A(n8128), .B(n8127), .ZN(n8129)
         );
  AOI21_X1 U9819 ( .B1(n8507), .B2(n8273), .A(n8129), .ZN(n8130) );
  OAI211_X1 U9820 ( .C1(n8132), .C2(n8276), .A(n8131), .B(n8130), .ZN(P2_U3159) );
  AOI22_X1 U9821 ( .A1(n8135), .A2(n8134), .B1(n8133), .B2(n8280), .ZN(n8138)
         );
  XNOR2_X1 U9822 ( .A(n5839), .B(n8136), .ZN(n8137) );
  XNOR2_X1 U9823 ( .A(n8138), .B(n8137), .ZN(n8146) );
  AOI22_X1 U9824 ( .A1(n8280), .A2(n8269), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8141) );
  NAND2_X1 U9825 ( .A1(n8139), .A2(n8273), .ZN(n8140) );
  OAI211_X1 U9826 ( .C1(n8142), .C2(n8271), .A(n8141), .B(n8140), .ZN(n8143)
         );
  AOI21_X1 U9827 ( .B1(n8144), .B2(n8236), .A(n8143), .ZN(n8145) );
  OAI21_X1 U9828 ( .B1(n8146), .B2(n8264), .A(n8145), .ZN(P2_U3160) );
  INV_X1 U9829 ( .A(n8147), .ZN(n8214) );
  INV_X1 U9830 ( .A(n8148), .ZN(n8150) );
  NOR3_X1 U9831 ( .A1(n8214), .A2(n8150), .A3(n8149), .ZN(n8153) );
  INV_X1 U9832 ( .A(n8151), .ZN(n8152) );
  OAI21_X1 U9833 ( .B1(n8153), .B2(n8152), .A(n8244), .ZN(n8157) );
  OAI22_X1 U9834 ( .A1(n8480), .A2(n8271), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10467), .ZN(n8155) );
  NOR2_X1 U9835 ( .A1(n8256), .A2(n8479), .ZN(n8154) );
  AOI211_X1 U9836 ( .C1(n8483), .C2(n8273), .A(n8155), .B(n8154), .ZN(n8156)
         );
  OAI211_X1 U9837 ( .C1(n8679), .C2(n8276), .A(n8157), .B(n8156), .ZN(P2_U3163) );
  XNOR2_X1 U9838 ( .A(n8159), .B(n8158), .ZN(n8168) );
  NOR2_X1 U9839 ( .A1(n8271), .A2(n8562), .ZN(n8160) );
  AOI211_X1 U9840 ( .C1(n8269), .C2(n8162), .A(n8161), .B(n8160), .ZN(n8163)
         );
  OAI21_X1 U9841 ( .B1(n8164), .B2(n8247), .A(n8163), .ZN(n8165) );
  AOI21_X1 U9842 ( .B1(n8166), .B2(n8236), .A(n8165), .ZN(n8167) );
  OAI21_X1 U9843 ( .B1(n8168), .B2(n8264), .A(n8167), .ZN(P2_U3164) );
  XOR2_X1 U9844 ( .A(n8170), .B(n8169), .Z(n8175) );
  AOI22_X1 U9845 ( .A1(n8281), .A2(n8269), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8172) );
  NAND2_X1 U9846 ( .A1(n8437), .A2(n8273), .ZN(n8171) );
  OAI211_X1 U9847 ( .C1(n8435), .C2(n8271), .A(n8172), .B(n8171), .ZN(n8173)
         );
  AOI21_X1 U9848 ( .B1(n8655), .B2(n8236), .A(n8173), .ZN(n8174) );
  OAI21_X1 U9849 ( .B1(n8175), .B2(n8264), .A(n8174), .ZN(P2_U3165) );
  INV_X1 U9850 ( .A(n8176), .ZN(n8191) );
  INV_X1 U9851 ( .A(n8178), .ZN(n8181) );
  INV_X1 U9852 ( .A(n8179), .ZN(n8180) );
  AOI21_X1 U9853 ( .B1(n8177), .B2(n8181), .A(n8180), .ZN(n8182) );
  OAI21_X1 U9854 ( .B1(n8191), .B2(n8182), .A(n8244), .ZN(n8186) );
  NAND2_X1 U9855 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8353) );
  OAI21_X1 U9856 ( .B1(n8271), .B2(n8516), .A(n8353), .ZN(n8184) );
  NOR2_X1 U9857 ( .A1(n8247), .A2(n8540), .ZN(n8183) );
  AOI211_X1 U9858 ( .C1(n8269), .C2(n8536), .A(n8184), .B(n8183), .ZN(n8185)
         );
  OAI211_X1 U9859 ( .C1(n8187), .C2(n8276), .A(n8186), .B(n8185), .ZN(P2_U3166) );
  INV_X1 U9860 ( .A(n8697), .ZN(n8199) );
  INV_X1 U9861 ( .A(n8188), .ZN(n8190) );
  NOR3_X1 U9862 ( .A1(n8191), .A2(n8190), .A3(n8189), .ZN(n8193) );
  INV_X1 U9863 ( .A(n8192), .ZN(n8243) );
  OAI21_X1 U9864 ( .B1(n8193), .B2(n8243), .A(n8244), .ZN(n8198) );
  INV_X1 U9865 ( .A(n8194), .ZN(n8530) );
  AND2_X1 U9866 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8374) );
  AOI21_X1 U9867 ( .B1(n8258), .B2(n8528), .A(n8374), .ZN(n8195) );
  OAI21_X1 U9868 ( .B1(n8256), .B2(n8550), .A(n8195), .ZN(n8196) );
  AOI21_X1 U9869 ( .B1(n8530), .B2(n8273), .A(n8196), .ZN(n8197) );
  OAI211_X1 U9870 ( .C1(n8199), .C2(n8276), .A(n8198), .B(n8197), .ZN(P2_U3168) );
  OAI22_X1 U9871 ( .A1(n8202), .A2(n8282), .B1(n8201), .B2(n8200), .ZN(n8205)
         );
  XNOR2_X1 U9872 ( .A(n8203), .B(n8460), .ZN(n8204) );
  XNOR2_X1 U9873 ( .A(n8205), .B(n8204), .ZN(n8210) );
  NOR2_X1 U9874 ( .A1(n8467), .A2(n8256), .ZN(n8207) );
  OAI22_X1 U9875 ( .A1(n8446), .A2(n8271), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10473), .ZN(n8206) );
  AOI211_X1 U9876 ( .C1(n8448), .C2(n8273), .A(n8207), .B(n8206), .ZN(n8209)
         );
  NAND2_X1 U9877 ( .A1(n8662), .A2(n8236), .ZN(n8208) );
  NOR3_X1 U9878 ( .A1(n4541), .A2(n4951), .A3(n8213), .ZN(n8215) );
  OAI21_X1 U9879 ( .B1(n8215), .B2(n8214), .A(n8244), .ZN(n8219) );
  INV_X1 U9880 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10454) );
  OAI22_X1 U9881 ( .A1(n8493), .A2(n8271), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10454), .ZN(n8217) );
  NOR2_X1 U9882 ( .A1(n8256), .A2(n8517), .ZN(n8216) );
  AOI211_X1 U9883 ( .C1(n8496), .C2(n8273), .A(n8217), .B(n8216), .ZN(n8218)
         );
  OAI211_X1 U9884 ( .C1(n8684), .C2(n8276), .A(n8219), .B(n8218), .ZN(P2_U3173) );
  AOI21_X1 U9885 ( .B1(n8222), .B2(n8221), .A(n8220), .ZN(n8230) );
  AND2_X1 U9886 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8304) );
  NOR2_X1 U9887 ( .A1(n8271), .A2(n8223), .ZN(n8224) );
  AOI211_X1 U9888 ( .C1(n8269), .C2(n8286), .A(n8304), .B(n8224), .ZN(n8225)
         );
  OAI21_X1 U9889 ( .B1(n8226), .B2(n8247), .A(n8225), .ZN(n8227) );
  AOI21_X1 U9890 ( .B1(n8228), .B2(n8236), .A(n8227), .ZN(n8229) );
  OAI21_X1 U9891 ( .B1(n8230), .B2(n8264), .A(n8229), .ZN(P2_U3174) );
  XNOR2_X1 U9892 ( .A(n8231), .B(n8480), .ZN(n8232) );
  XNOR2_X1 U9893 ( .A(n8233), .B(n8232), .ZN(n8239) );
  INV_X1 U9894 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10268) );
  OAI22_X1 U9895 ( .A1(n8256), .A2(n8493), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10268), .ZN(n8235) );
  NOR2_X1 U9896 ( .A1(n8467), .A2(n8271), .ZN(n8234) );
  AOI211_X1 U9897 ( .C1(n8471), .C2(n8273), .A(n8235), .B(n8234), .ZN(n8238)
         );
  NAND2_X1 U9898 ( .A1(n8470), .A2(n8236), .ZN(n8237) );
  OAI211_X1 U9899 ( .C1(n8239), .C2(n8264), .A(n8238), .B(n8237), .ZN(P2_U3175) );
  INV_X1 U9900 ( .A(n8240), .ZN(n8242) );
  NOR3_X1 U9901 ( .A1(n8243), .A2(n8242), .A3(n8241), .ZN(n8246) );
  OAI21_X1 U9902 ( .B1(n8246), .B2(n8245), .A(n8244), .ZN(n8251) );
  NAND2_X1 U9903 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8390) );
  OAI21_X1 U9904 ( .B1(n8271), .B2(n8517), .A(n8390), .ZN(n8249) );
  NOR2_X1 U9905 ( .A1(n8247), .A2(n8518), .ZN(n8248) );
  AOI211_X1 U9906 ( .C1(n8269), .C2(n8537), .A(n8249), .B(n8248), .ZN(n8250)
         );
  OAI211_X1 U9907 ( .C1(n8252), .C2(n8276), .A(n8251), .B(n8250), .ZN(P2_U3178) );
  XNOR2_X1 U9908 ( .A(n8253), .B(n8435), .ZN(n8254) );
  XNOR2_X1 U9909 ( .A(n8255), .B(n8254), .ZN(n8263) );
  OAI22_X1 U9910 ( .A1(n8446), .A2(n8256), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10456), .ZN(n8257) );
  AOI21_X1 U9911 ( .B1(n8280), .B2(n8258), .A(n8257), .ZN(n8260) );
  NAND2_X1 U9912 ( .A1(n8421), .A2(n8273), .ZN(n8259) );
  OAI211_X1 U9913 ( .C1(n8584), .C2(n8276), .A(n8260), .B(n8259), .ZN(n8261)
         );
  INV_X1 U9914 ( .A(n8261), .ZN(n8262) );
  OAI21_X1 U9915 ( .B1(n8263), .B2(n8264), .A(n8262), .ZN(P2_U3180) );
  INV_X1 U9916 ( .A(n8709), .ZN(n8277) );
  AOI21_X1 U9917 ( .B1(n8266), .B2(n8265), .A(n8264), .ZN(n8267) );
  NAND2_X1 U9918 ( .A1(n8267), .A2(n8177), .ZN(n8275) );
  INV_X1 U9919 ( .A(n8268), .ZN(n8553) );
  NAND2_X1 U9920 ( .A1(n8269), .A2(n8548), .ZN(n8270) );
  NAND2_X1 U9921 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8339) );
  OAI211_X1 U9922 ( .C1(n8550), .C2(n8271), .A(n8270), .B(n8339), .ZN(n8272)
         );
  AOI21_X1 U9923 ( .B1(n8553), .B2(n8273), .A(n8272), .ZN(n8274) );
  OAI211_X1 U9924 ( .C1(n8277), .C2(n8276), .A(n8275), .B(n8274), .ZN(P2_U3181) );
  MUX2_X1 U9925 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8400), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9926 ( .A(n8279), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8292), .Z(
        P2_U3521) );
  MUX2_X1 U9927 ( .A(n8410), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8292), .Z(
        P2_U3519) );
  MUX2_X1 U9928 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8280), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9929 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8411), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9930 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8281), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9931 ( .A(n8282), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8292), .Z(
        P2_U3514) );
  MUX2_X1 U9932 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8283), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9933 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8505), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9934 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8284), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9935 ( .A(n8528), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8292), .Z(
        P2_U3509) );
  MUX2_X1 U9936 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8537), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9937 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8527), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9938 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8536), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9939 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8548), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9940 ( .A(n8285), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8292), .Z(
        P2_U3504) );
  MUX2_X1 U9941 ( .A(n8286), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8292), .Z(
        P2_U3503) );
  MUX2_X1 U9942 ( .A(n8287), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8292), .Z(
        P2_U3501) );
  MUX2_X1 U9943 ( .A(n8288), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8292), .Z(
        P2_U3499) );
  MUX2_X1 U9944 ( .A(n8289), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8292), .Z(
        P2_U3498) );
  MUX2_X1 U9945 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8290), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8291), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U9947 ( .A(n9971), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8292), .Z(
        P2_U3495) );
  MUX2_X1 U9948 ( .A(n9984), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8292), .Z(
        P2_U3494) );
  MUX2_X1 U9949 ( .A(n5398), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8292), .Z(
        P2_U3493) );
  MUX2_X1 U9950 ( .A(n9985), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8292), .Z(
        P2_U3492) );
  MUX2_X1 U9951 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n8293), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI21_X1 U9952 ( .B1(n8296), .B2(n8295), .A(n8294), .ZN(n8311) );
  OAI21_X1 U9953 ( .B1(n8299), .B2(n8298), .A(n8297), .ZN(n8300) );
  NAND2_X1 U9954 ( .A1(n8300), .A2(n9964), .ZN(n8310) );
  AOI21_X1 U9955 ( .B1(n8303), .B2(n8302), .A(n8301), .ZN(n8307) );
  AOI21_X1 U9956 ( .B1(n9915), .B2(n8305), .A(n8304), .ZN(n8306) );
  OAI21_X1 U9957 ( .B1(n9953), .B2(n8307), .A(n8306), .ZN(n8308) );
  AOI21_X1 U9958 ( .B1(n9933), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n8308), .ZN(
        n8309) );
  OAI211_X1 U9959 ( .C1(n8311), .C2(n9948), .A(n8310), .B(n8309), .ZN(P2_U3195) );
  AOI21_X1 U9960 ( .B1(n8314), .B2(n8313), .A(n8312), .ZN(n8329) );
  OAI21_X1 U9961 ( .B1(n8317), .B2(n8316), .A(n8315), .ZN(n8327) );
  NAND2_X1 U9962 ( .A1(n9933), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8319) );
  OAI211_X1 U9963 ( .C1(n9957), .C2(n8320), .A(n8319), .B(n8318), .ZN(n8326)
         );
  AOI21_X1 U9964 ( .B1(n8323), .B2(n8322), .A(n8321), .ZN(n8324) );
  NOR2_X1 U9965 ( .A1(n8324), .A2(n9948), .ZN(n8325) );
  AOI211_X1 U9966 ( .C1(n9964), .C2(n8327), .A(n8326), .B(n8325), .ZN(n8328)
         );
  OAI21_X1 U9967 ( .B1(n8329), .B2(n9953), .A(n8328), .ZN(P2_U3196) );
  AOI21_X1 U9968 ( .B1(n8332), .B2(n8331), .A(n8330), .ZN(n8346) );
  OAI21_X1 U9969 ( .B1(n8335), .B2(n8334), .A(n8333), .ZN(n8344) );
  AOI21_X1 U9970 ( .B1(n8337), .B2(n8623), .A(n8336), .ZN(n8338) );
  NOR2_X1 U9971 ( .A1(n8338), .A2(n9953), .ZN(n8343) );
  NAND2_X1 U9972 ( .A1(n9933), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8340) );
  OAI211_X1 U9973 ( .C1(n9957), .C2(n8341), .A(n8340), .B(n8339), .ZN(n8342)
         );
  AOI211_X1 U9974 ( .C1(n9964), .C2(n8344), .A(n8343), .B(n8342), .ZN(n8345)
         );
  OAI21_X1 U9975 ( .B1(n8346), .B2(n9948), .A(n8345), .ZN(P2_U3197) );
  AOI21_X1 U9976 ( .B1(n8349), .B2(n8348), .A(n8347), .ZN(n8364) );
  OAI21_X1 U9977 ( .B1(n8352), .B2(n8351), .A(n8350), .ZN(n8357) );
  OAI21_X1 U9978 ( .B1(n9957), .B2(n8354), .A(n8353), .ZN(n8356) );
  INV_X1 U9979 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10115) );
  NOR2_X1 U9980 ( .A1(n9969), .A2(n10115), .ZN(n8355) );
  AOI211_X1 U9981 ( .C1(n9964), .C2(n8357), .A(n8356), .B(n8355), .ZN(n8363)
         );
  AOI21_X1 U9982 ( .B1(n8360), .B2(n8359), .A(n8358), .ZN(n8361) );
  OR2_X1 U9983 ( .A1(n8361), .A2(n9948), .ZN(n8362) );
  OAI211_X1 U9984 ( .C1(n8364), .C2(n9953), .A(n8363), .B(n8362), .ZN(P2_U3198) );
  AOI21_X1 U9985 ( .B1(n8367), .B2(n8366), .A(n8365), .ZN(n8381) );
  OAI21_X1 U9986 ( .B1(n8370), .B2(n8369), .A(n8368), .ZN(n8380) );
  AOI21_X1 U9987 ( .B1(n9915), .B2(n8375), .A(n8374), .ZN(n8376) );
  OAI21_X1 U9988 ( .B1(n9953), .B2(n8377), .A(n8376), .ZN(n8379) );
  INV_X1 U9989 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10120) );
  NOR2_X1 U9990 ( .A1(n9969), .A2(n10120), .ZN(n8378) );
  AOI21_X1 U9991 ( .B1(n8384), .B2(n8383), .A(n8382), .ZN(n8398) );
  AND2_X1 U9992 ( .A1(n8386), .A2(n8385), .ZN(n8387) );
  AOI21_X1 U9993 ( .B1(n8387), .B2(P2_U3893), .A(n9915), .ZN(n8392) );
  INV_X1 U9994 ( .A(n8387), .ZN(n8388) );
  NAND3_X1 U9995 ( .A1(n8388), .A2(n9964), .A3(n8391), .ZN(n8389) );
  OAI211_X1 U9996 ( .C1(n8392), .C2(n8391), .A(n8390), .B(n8389), .ZN(n8396)
         );
  OAI21_X1 U9997 ( .B1(n8398), .B2(n9953), .A(n8397), .ZN(P2_U3200) );
  NAND2_X1 U9998 ( .A1(n8633), .A2(n8555), .ZN(n8402) );
  NAND2_X1 U9999 ( .A1(n8400), .A2(n8399), .ZN(n8575) );
  INV_X1 U10000 ( .A(n8575), .ZN(n8634) );
  AOI21_X1 U10001 ( .B1(n8634), .B2(n9999), .A(n8401), .ZN(n8405) );
  OAI211_X1 U10002 ( .C1(n9999), .C2(n8403), .A(n8402), .B(n8405), .ZN(
        P2_U3202) );
  NAND2_X1 U10003 ( .A1(n5088), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8404) );
  OAI211_X1 U10004 ( .C1(n8580), .C2(n9975), .A(n8405), .B(n8404), .ZN(
        P2_U3203) );
  XNOR2_X1 U10005 ( .A(n8407), .B(n8406), .ZN(n8645) );
  INV_X1 U10006 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8416) );
  XNOR2_X1 U10007 ( .A(n8409), .B(n8408), .ZN(n8415) );
  MUX2_X1 U10008 ( .A(n8416), .B(n8640), .S(n9999), .Z(n8419) );
  AOI22_X1 U10009 ( .A1(n8642), .A2(n8555), .B1(n8554), .B2(n8417), .ZN(n8418)
         );
  OAI211_X1 U10010 ( .C1(n8645), .C2(n8558), .A(n8419), .B(n8418), .ZN(
        P2_U3206) );
  XNOR2_X1 U10011 ( .A(n8420), .B(n8423), .ZN(n8652) );
  INV_X1 U10012 ( .A(n8652), .ZN(n8432) );
  INV_X1 U10013 ( .A(n8421), .ZN(n8422) );
  OAI22_X1 U10014 ( .A1(n8584), .A2(n9975), .B1(n9990), .B2(n8422), .ZN(n8431)
         );
  NOR2_X1 U10015 ( .A1(n8587), .A2(n8443), .ZN(n8436) );
  XOR2_X1 U10016 ( .A(n8439), .B(n8433), .Z(n8434) );
  OAI222_X1 U10017 ( .A1(n8565), .A2(n8435), .B1(n8563), .B2(n8460), .C1(n8561), .C2(n8434), .ZN(n8653) );
  AOI211_X1 U10018 ( .C1(n8554), .C2(n8437), .A(n8436), .B(n8653), .ZN(n8442)
         );
  XOR2_X1 U10019 ( .A(n8439), .B(n8438), .Z(n8658) );
  INV_X1 U10020 ( .A(n8658), .ZN(n8440) );
  AOI22_X1 U10021 ( .A1(n8440), .A2(n9977), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n5088), .ZN(n8441) );
  OAI21_X1 U10022 ( .B1(n8442), .B2(n5088), .A(n8441), .ZN(P2_U3208) );
  NOR2_X1 U10023 ( .A1(n8590), .A2(n8443), .ZN(n8447) );
  XNOR2_X1 U10024 ( .A(n8444), .B(n8452), .ZN(n8445) );
  OAI222_X1 U10025 ( .A1(n8563), .A2(n8467), .B1(n8565), .B2(n8446), .C1(n8445), .C2(n8561), .ZN(n8659) );
  AOI211_X1 U10026 ( .C1(n8554), .C2(n8448), .A(n8447), .B(n8659), .ZN(n8455)
         );
  NOR2_X1 U10027 ( .A1(n8450), .A2(n8449), .ZN(n8451) );
  XOR2_X1 U10028 ( .A(n8452), .B(n8451), .Z(n8665) );
  INV_X1 U10029 ( .A(n8665), .ZN(n8453) );
  AOI22_X1 U10030 ( .A1(n8453), .A2(n9977), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n5088), .ZN(n8454) );
  OAI21_X1 U10031 ( .B1(n8455), .B2(n5088), .A(n8454), .ZN(P2_U3209) );
  XOR2_X1 U10032 ( .A(n8456), .B(n8458), .Z(n8671) );
  INV_X1 U10033 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8461) );
  XOR2_X1 U10034 ( .A(n8458), .B(n8457), .Z(n8459) );
  OAI222_X1 U10035 ( .A1(n8563), .A2(n8480), .B1(n8565), .B2(n8460), .C1(n8561), .C2(n8459), .ZN(n8593) );
  INV_X1 U10036 ( .A(n8593), .ZN(n8666) );
  MUX2_X1 U10037 ( .A(n8461), .B(n8666), .S(n9999), .Z(n8464) );
  AOI22_X1 U10038 ( .A1(n8668), .A2(n8555), .B1(n8554), .B2(n8462), .ZN(n8463)
         );
  OAI211_X1 U10039 ( .C1(n8671), .C2(n8558), .A(n8464), .B(n8463), .ZN(
        P2_U3210) );
  XOR2_X1 U10040 ( .A(n8468), .B(n8465), .Z(n8466) );
  OAI222_X1 U10041 ( .A1(n8563), .A2(n8493), .B1(n8565), .B2(n8467), .C1(n8561), .C2(n8466), .ZN(n8597) );
  INV_X1 U10042 ( .A(n8597), .ZN(n8475) );
  XNOR2_X1 U10043 ( .A(n8469), .B(n8468), .ZN(n8598) );
  INV_X1 U10044 ( .A(n8470), .ZN(n8675) );
  AOI22_X1 U10045 ( .A1(n5088), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8471), .B2(
        n8554), .ZN(n8472) );
  OAI21_X1 U10046 ( .B1(n8675), .B2(n9975), .A(n8472), .ZN(n8473) );
  AOI21_X1 U10047 ( .B1(n8598), .B2(n9977), .A(n8473), .ZN(n8474) );
  OAI21_X1 U10048 ( .B1(n8475), .B2(n5088), .A(n8474), .ZN(P2_U3211) );
  XNOR2_X1 U10049 ( .A(n8477), .B(n8476), .ZN(n8478) );
  OAI222_X1 U10050 ( .A1(n8565), .A2(n8480), .B1(n8563), .B2(n8479), .C1(n8561), .C2(n8478), .ZN(n8601) );
  INV_X1 U10051 ( .A(n8601), .ZN(n8487) );
  XNOR2_X1 U10052 ( .A(n8482), .B(n8481), .ZN(n8602) );
  AOI22_X1 U10053 ( .A1(n5088), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8554), .B2(
        n8483), .ZN(n8484) );
  OAI21_X1 U10054 ( .B1(n8679), .B2(n9975), .A(n8484), .ZN(n8485) );
  AOI21_X1 U10055 ( .B1(n8602), .B2(n9977), .A(n8485), .ZN(n8486) );
  OAI21_X1 U10056 ( .B1(n8487), .B2(n5088), .A(n8486), .ZN(P2_U3212) );
  OAI21_X1 U10057 ( .B1(n8490), .B2(n8489), .A(n8488), .ZN(n8491) );
  INV_X1 U10058 ( .A(n8491), .ZN(n8492) );
  OAI222_X1 U10059 ( .A1(n8565), .A2(n8493), .B1(n8563), .B2(n8517), .C1(n8561), .C2(n8492), .ZN(n8605) );
  INV_X1 U10060 ( .A(n8605), .ZN(n8500) );
  XNOR2_X1 U10061 ( .A(n8495), .B(n8494), .ZN(n8606) );
  AOI22_X1 U10062 ( .A1(n5088), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8554), .B2(
        n8496), .ZN(n8497) );
  OAI21_X1 U10063 ( .B1(n8684), .B2(n9975), .A(n8497), .ZN(n8498) );
  AOI21_X1 U10064 ( .B1(n8606), .B2(n9977), .A(n8498), .ZN(n8499) );
  OAI21_X1 U10065 ( .B1(n8500), .B2(n5088), .A(n8499), .ZN(P2_U3213) );
  AOI21_X1 U10066 ( .B1(n8512), .B2(n8501), .A(n8503), .ZN(n8502) );
  NOR2_X1 U10067 ( .A1(n4595), .A2(n8502), .ZN(n8690) );
  XNOR2_X1 U10068 ( .A(n8504), .B(n8503), .ZN(n8506) );
  AOI222_X1 U10069 ( .A1(n9981), .A2(n8506), .B1(n8528), .B2(n9986), .C1(n8505), .C2(n9983), .ZN(n8685) );
  MUX2_X1 U10070 ( .A(n5268), .B(n8685), .S(n9999), .Z(n8509) );
  AOI22_X1 U10071 ( .A1(n8687), .A2(n8555), .B1(n8554), .B2(n8507), .ZN(n8508)
         );
  OAI211_X1 U10072 ( .C1(n8690), .C2(n8558), .A(n8509), .B(n8508), .ZN(
        P2_U3214) );
  OR2_X1 U10073 ( .A1(n8510), .A2(n8513), .ZN(n8511) );
  NAND2_X1 U10074 ( .A1(n8512), .A2(n8511), .ZN(n8694) );
  XNOR2_X1 U10075 ( .A(n8514), .B(n8513), .ZN(n8515) );
  OAI222_X1 U10076 ( .A1(n8565), .A2(n8517), .B1(n8563), .B2(n8516), .C1(n8515), .C2(n8561), .ZN(n8613) );
  NAND2_X1 U10077 ( .A1(n8613), .A2(n9999), .ZN(n8522) );
  OAI22_X1 U10078 ( .A1(n9999), .A2(n8519), .B1(n8518), .B2(n9990), .ZN(n8520)
         );
  AOI21_X1 U10079 ( .B1(n8614), .B2(n8555), .A(n8520), .ZN(n8521) );
  OAI211_X1 U10080 ( .C1(n8694), .C2(n8558), .A(n8522), .B(n8521), .ZN(
        P2_U3215) );
  XNOR2_X1 U10081 ( .A(n8524), .B(n8523), .ZN(n8700) );
  XNOR2_X1 U10082 ( .A(n8526), .B(n8525), .ZN(n8529) );
  AOI222_X1 U10083 ( .A1(n9981), .A2(n8529), .B1(n8528), .B2(n9983), .C1(n8527), .C2(n9986), .ZN(n8695) );
  MUX2_X1 U10084 ( .A(n8367), .B(n8695), .S(n9999), .Z(n8532) );
  AOI22_X1 U10085 ( .A1(n8697), .A2(n8555), .B1(n8554), .B2(n8530), .ZN(n8531)
         );
  OAI211_X1 U10086 ( .C1(n8700), .C2(n8558), .A(n8532), .B(n8531), .ZN(
        P2_U3216) );
  XNOR2_X1 U10087 ( .A(n8533), .B(n8535), .ZN(n8706) );
  XOR2_X1 U10088 ( .A(n8534), .B(n8535), .Z(n8538) );
  AOI222_X1 U10089 ( .A1(n9981), .A2(n8538), .B1(n8537), .B2(n9983), .C1(n8536), .C2(n9986), .ZN(n8701) );
  MUX2_X1 U10090 ( .A(n8539), .B(n8701), .S(n9999), .Z(n8543) );
  INV_X1 U10091 ( .A(n8540), .ZN(n8541) );
  AOI22_X1 U10092 ( .A1(n8703), .A2(n8555), .B1(n8554), .B2(n8541), .ZN(n8542)
         );
  OAI211_X1 U10093 ( .C1(n8706), .C2(n8558), .A(n8543), .B(n8542), .ZN(
        P2_U3217) );
  XNOR2_X1 U10094 ( .A(n8544), .B(n8545), .ZN(n8713) );
  XNOR2_X1 U10095 ( .A(n8547), .B(n8546), .ZN(n8552) );
  NAND2_X1 U10096 ( .A1(n8548), .A2(n9986), .ZN(n8549) );
  OAI21_X1 U10097 ( .B1(n8550), .B2(n8565), .A(n8549), .ZN(n8551) );
  AOI21_X1 U10098 ( .B1(n8552), .B2(n9981), .A(n8551), .ZN(n8707) );
  MUX2_X1 U10099 ( .A(n8332), .B(n8707), .S(n9999), .Z(n8557) );
  AOI22_X1 U10100 ( .A1(n8709), .A2(n8555), .B1(n8554), .B2(n8553), .ZN(n8556)
         );
  OAI211_X1 U10101 ( .C1(n8713), .C2(n8558), .A(n8557), .B(n8556), .ZN(
        P2_U3218) );
  XOR2_X1 U10102 ( .A(n8559), .B(n8567), .Z(n8560) );
  OAI222_X1 U10103 ( .A1(n8565), .A2(n8564), .B1(n8563), .B2(n8562), .C1(n8561), .C2(n8560), .ZN(n8627) );
  AOI21_X1 U10104 ( .B1(n8566), .B2(n8716), .A(n8627), .ZN(n8574) );
  INV_X1 U10105 ( .A(n8567), .ZN(n8568) );
  XNOR2_X1 U10106 ( .A(n8569), .B(n8568), .ZN(n8719) );
  OAI22_X1 U10107 ( .A1(n9999), .A2(n8571), .B1(n8570), .B2(n9990), .ZN(n8572)
         );
  AOI21_X1 U10108 ( .B1(n8719), .B2(n9977), .A(n8572), .ZN(n8573) );
  OAI21_X1 U10109 ( .B1(n8574), .B2(n5088), .A(n8573), .ZN(P2_U3219) );
  NOR2_X1 U10110 ( .A1(n8575), .A2(n10062), .ZN(n8578) );
  AOI21_X1 U10111 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10062), .A(n8578), .ZN(
        n8576) );
  OAI21_X1 U10112 ( .B1(n8577), .B2(n8609), .A(n8576), .ZN(P2_U3490) );
  AOI21_X1 U10113 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10062), .A(n8578), .ZN(
        n8579) );
  OAI21_X1 U10114 ( .B1(n8580), .B2(n8609), .A(n8579), .ZN(P2_U3489) );
  NAND2_X1 U10115 ( .A1(n8642), .A2(n8629), .ZN(n8582) );
  OAI211_X1 U10116 ( .C1(n8645), .C2(n8626), .A(n8583), .B(n8582), .ZN(
        P2_U3486) );
  MUX2_X1 U10117 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8646), .S(n10064), .Z(
        n8586) );
  OAI22_X1 U10118 ( .A1(n8652), .A2(n8626), .B1(n8584), .B2(n8609), .ZN(n8585)
         );
  OR2_X1 U10119 ( .A1(n8586), .A2(n8585), .ZN(P2_U3485) );
  MUX2_X1 U10120 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8653), .S(n10064), .Z(
        n8589) );
  OAI22_X1 U10121 ( .A1(n8658), .A2(n8626), .B1(n8587), .B2(n8609), .ZN(n8588)
         );
  OR2_X1 U10122 ( .A1(n8589), .A2(n8588), .ZN(P2_U3484) );
  MUX2_X1 U10123 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8659), .S(n10064), .Z(
        n8592) );
  OAI22_X1 U10124 ( .A1(n8665), .A2(n8626), .B1(n8590), .B2(n8609), .ZN(n8591)
         );
  OR2_X1 U10125 ( .A1(n8592), .A2(n8591), .ZN(P2_U3483) );
  MUX2_X1 U10126 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8593), .S(n10064), .Z(
        n8596) );
  OAI22_X1 U10127 ( .A1(n8671), .A2(n8626), .B1(n8594), .B2(n8609), .ZN(n8595)
         );
  OR2_X1 U10128 ( .A1(n8596), .A2(n8595), .ZN(P2_U3482) );
  INV_X1 U10129 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8599) );
  AOI21_X1 U10130 ( .B1(n10035), .B2(n8598), .A(n8597), .ZN(n8672) );
  MUX2_X1 U10131 ( .A(n8599), .B(n8672), .S(n10064), .Z(n8600) );
  OAI21_X1 U10132 ( .B1(n8675), .B2(n8609), .A(n8600), .ZN(P2_U3481) );
  INV_X1 U10133 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8603) );
  AOI21_X1 U10134 ( .B1(n8602), .B2(n10035), .A(n8601), .ZN(n8676) );
  MUX2_X1 U10135 ( .A(n8603), .B(n8676), .S(n10064), .Z(n8604) );
  OAI21_X1 U10136 ( .B1(n8679), .B2(n8609), .A(n8604), .ZN(P2_U3480) );
  INV_X1 U10137 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8607) );
  AOI21_X1 U10138 ( .B1(n8606), .B2(n10035), .A(n8605), .ZN(n8680) );
  MUX2_X1 U10139 ( .A(n8607), .B(n8680), .S(n10064), .Z(n8608) );
  OAI21_X1 U10140 ( .B1(n8684), .B2(n8609), .A(n8608), .ZN(P2_U3479) );
  MUX2_X1 U10141 ( .A(n8610), .B(n8685), .S(n10064), .Z(n8612) );
  NAND2_X1 U10142 ( .A1(n8687), .A2(n8629), .ZN(n8611) );
  OAI211_X1 U10143 ( .C1(n8690), .C2(n8626), .A(n8612), .B(n8611), .ZN(
        P2_U3478) );
  AOI21_X1 U10144 ( .B1(n10040), .B2(n8614), .A(n8613), .ZN(n8691) );
  MUX2_X1 U10145 ( .A(n8615), .B(n8691), .S(n10064), .Z(n8616) );
  OAI21_X1 U10146 ( .B1(n8626), .B2(n8694), .A(n8616), .ZN(P2_U3477) );
  MUX2_X1 U10147 ( .A(n8617), .B(n8695), .S(n10064), .Z(n8619) );
  NAND2_X1 U10148 ( .A1(n8697), .A2(n8629), .ZN(n8618) );
  OAI211_X1 U10149 ( .C1(n8626), .C2(n8700), .A(n8619), .B(n8618), .ZN(
        P2_U3476) );
  MUX2_X1 U10150 ( .A(n8620), .B(n8701), .S(n10064), .Z(n8622) );
  NAND2_X1 U10151 ( .A1(n8703), .A2(n8629), .ZN(n8621) );
  OAI211_X1 U10152 ( .C1(n8706), .C2(n8626), .A(n8622), .B(n8621), .ZN(
        P2_U3475) );
  MUX2_X1 U10153 ( .A(n8623), .B(n8707), .S(n10064), .Z(n8625) );
  NAND2_X1 U10154 ( .A1(n8709), .A2(n8629), .ZN(n8624) );
  OAI211_X1 U10155 ( .C1(n8626), .C2(n8713), .A(n8625), .B(n8624), .ZN(
        P2_U3474) );
  INV_X1 U10156 ( .A(n8627), .ZN(n8714) );
  MUX2_X1 U10157 ( .A(n8628), .B(n8714), .S(n10064), .Z(n8632) );
  AOI22_X1 U10158 ( .A1(n8719), .A2(n8630), .B1(n8629), .B2(n8716), .ZN(n8631)
         );
  NAND2_X1 U10159 ( .A1(n8632), .A2(n8631), .ZN(P2_U3473) );
  INV_X1 U10160 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U10161 ( .A1(n8633), .A2(n8717), .ZN(n8635) );
  NAND2_X1 U10162 ( .A1(n8634), .A2(n10048), .ZN(n8638) );
  OAI211_X1 U10163 ( .C1(n8636), .C2(n10048), .A(n8635), .B(n8638), .ZN(
        P2_U3458) );
  NAND2_X1 U10164 ( .A1(n8637), .A2(n8717), .ZN(n8639) );
  OAI211_X1 U10165 ( .C1(n6573), .C2(n10048), .A(n8639), .B(n8638), .ZN(
        P2_U3457) );
  MUX2_X1 U10166 ( .A(n8641), .B(n8640), .S(n10048), .Z(n8644) );
  NAND2_X1 U10167 ( .A1(n8642), .A2(n8717), .ZN(n8643) );
  OAI211_X1 U10168 ( .C1(n8645), .C2(n8712), .A(n8644), .B(n8643), .ZN(
        P2_U3454) );
  INV_X1 U10169 ( .A(n8646), .ZN(n8647) );
  MUX2_X1 U10170 ( .A(n8648), .B(n8647), .S(n10048), .Z(n8651) );
  NAND2_X1 U10171 ( .A1(n8649), .A2(n8717), .ZN(n8650) );
  OAI211_X1 U10172 ( .C1(n8652), .C2(n8712), .A(n8651), .B(n8650), .ZN(
        P2_U3453) );
  NAND2_X1 U10173 ( .A1(n8655), .A2(n8717), .ZN(n8656) );
  OAI211_X1 U10174 ( .C1(n8658), .C2(n8712), .A(n8657), .B(n8656), .ZN(
        P2_U3452) );
  INV_X1 U10175 ( .A(n8659), .ZN(n8660) );
  MUX2_X1 U10176 ( .A(n8661), .B(n8660), .S(n10048), .Z(n8664) );
  NAND2_X1 U10177 ( .A1(n8662), .A2(n8717), .ZN(n8663) );
  OAI211_X1 U10178 ( .C1(n8665), .C2(n8712), .A(n8664), .B(n8663), .ZN(
        P2_U3451) );
  MUX2_X1 U10179 ( .A(n8667), .B(n8666), .S(n10048), .Z(n8670) );
  NAND2_X1 U10180 ( .A1(n8668), .A2(n8717), .ZN(n8669) );
  OAI211_X1 U10181 ( .C1(n8671), .C2(n8712), .A(n8670), .B(n8669), .ZN(
        P2_U3450) );
  INV_X1 U10182 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8673) );
  MUX2_X1 U10183 ( .A(n8673), .B(n8672), .S(n10048), .Z(n8674) );
  OAI21_X1 U10184 ( .B1(n8675), .B2(n8683), .A(n8674), .ZN(P2_U3449) );
  INV_X1 U10185 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8677) );
  MUX2_X1 U10186 ( .A(n8677), .B(n8676), .S(n10048), .Z(n8678) );
  OAI21_X1 U10187 ( .B1(n8679), .B2(n8683), .A(n8678), .ZN(P2_U3448) );
  INV_X1 U10188 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8681) );
  MUX2_X1 U10189 ( .A(n8681), .B(n8680), .S(n10048), .Z(n8682) );
  OAI21_X1 U10190 ( .B1(n8684), .B2(n8683), .A(n8682), .ZN(P2_U3447) );
  MUX2_X1 U10191 ( .A(n8686), .B(n8685), .S(n10048), .Z(n8689) );
  NAND2_X1 U10192 ( .A1(n8687), .A2(n8717), .ZN(n8688) );
  OAI211_X1 U10193 ( .C1(n8690), .C2(n8712), .A(n8689), .B(n8688), .ZN(
        P2_U3446) );
  MUX2_X1 U10194 ( .A(n8692), .B(n8691), .S(n10048), .Z(n8693) );
  OAI21_X1 U10195 ( .B1(n8694), .B2(n8712), .A(n8693), .ZN(P2_U3444) );
  INV_X1 U10196 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8696) );
  MUX2_X1 U10197 ( .A(n8696), .B(n8695), .S(n10048), .Z(n8699) );
  NAND2_X1 U10198 ( .A1(n8697), .A2(n8717), .ZN(n8698) );
  OAI211_X1 U10199 ( .C1(n8700), .C2(n8712), .A(n8699), .B(n8698), .ZN(
        P2_U3441) );
  INV_X1 U10200 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8702) );
  MUX2_X1 U10201 ( .A(n8702), .B(n8701), .S(n10048), .Z(n8705) );
  NAND2_X1 U10202 ( .A1(n8703), .A2(n8717), .ZN(n8704) );
  OAI211_X1 U10203 ( .C1(n8706), .C2(n8712), .A(n8705), .B(n8704), .ZN(
        P2_U3438) );
  INV_X1 U10204 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8708) );
  MUX2_X1 U10205 ( .A(n8708), .B(n8707), .S(n10048), .Z(n8711) );
  NAND2_X1 U10206 ( .A1(n8709), .A2(n8717), .ZN(n8710) );
  OAI211_X1 U10207 ( .C1(n8713), .C2(n8712), .A(n8711), .B(n8710), .ZN(
        P2_U3435) );
  INV_X1 U10208 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8715) );
  MUX2_X1 U10209 ( .A(n8715), .B(n8714), .S(n10048), .Z(n8721) );
  AOI22_X1 U10210 ( .A1(n8719), .A2(n8718), .B1(n8717), .B2(n8716), .ZN(n8720)
         );
  NAND2_X1 U10211 ( .A1(n8721), .A2(n8720), .ZN(P2_U3432) );
  INV_X1 U10212 ( .A(n8874), .ZN(n9631) );
  NAND3_X1 U10213 ( .A1(n8722), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8725) );
  OAI22_X1 U10214 ( .A1(n8726), .A2(n8725), .B1(n8724), .B2(n8723), .ZN(n8727)
         );
  INV_X1 U10215 ( .A(n8727), .ZN(n8728) );
  OAI21_X1 U10216 ( .B1(n9631), .B2(n8729), .A(n8728), .ZN(P2_U3264) );
  MUX2_X1 U10217 ( .A(n8730), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10218 ( .B1(n8731), .B2(n4583), .A(n8783), .ZN(n8732) );
  NAND2_X1 U10219 ( .A1(n8732), .A2(n8830), .ZN(n8737) );
  INV_X1 U10220 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8733) );
  OAI22_X1 U10221 ( .A1(n8834), .A2(n8757), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8733), .ZN(n8735) );
  NOR2_X1 U10222 ( .A1(n8798), .A2(n9495), .ZN(n8734) );
  AOI211_X1 U10223 ( .C1(n8837), .C2(n9455), .A(n8735), .B(n8734), .ZN(n8736)
         );
  OAI211_X1 U10224 ( .C1(n9457), .C2(n8840), .A(n8737), .B(n8736), .ZN(
        P1_U3216) );
  AOI21_X1 U10225 ( .B1(n8740), .B2(n8739), .A(n8738), .ZN(n8745) );
  INV_X1 U10226 ( .A(n8837), .ZN(n8817) );
  NAND2_X1 U10227 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9343) );
  OAI21_X1 U10228 ( .B1(n9532), .B2(n8834), .A(n9343), .ZN(n8741) );
  AOI21_X1 U10229 ( .B1(n8832), .B2(n9138), .A(n8741), .ZN(n8742) );
  OAI21_X1 U10230 ( .B1(n9523), .B2(n8817), .A(n8742), .ZN(n8743) );
  AOI21_X1 U10231 ( .B1(n9603), .B2(n8821), .A(n8743), .ZN(n8744) );
  OAI21_X1 U10232 ( .B1(n8745), .B2(n8823), .A(n8744), .ZN(P1_U3219) );
  XNOR2_X1 U10233 ( .A(n8746), .B(n8747), .ZN(n8752) );
  AOI22_X1 U10234 ( .A1(n9136), .A2(n8832), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8749) );
  NAND2_X1 U10235 ( .A1(n8837), .A2(n9497), .ZN(n8748) );
  OAI211_X1 U10236 ( .C1(n9495), .C2(n8834), .A(n8749), .B(n8748), .ZN(n8750)
         );
  AOI21_X1 U10237 ( .B1(n9593), .B2(n8821), .A(n8750), .ZN(n8751) );
  OAI21_X1 U10238 ( .B1(n8752), .B2(n8823), .A(n8751), .ZN(P1_U3223) );
  AOI21_X1 U10239 ( .B1(n8754), .B2(n8753), .A(n8828), .ZN(n8762) );
  INV_X1 U10240 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8755) );
  OAI22_X1 U10241 ( .A1(n8834), .A2(n8756), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8755), .ZN(n8759) );
  NOR2_X1 U10242 ( .A1(n8798), .A2(n8757), .ZN(n8758) );
  AOI211_X1 U10243 ( .C1(n8837), .C2(n9428), .A(n8759), .B(n8758), .ZN(n8761)
         );
  NAND2_X1 U10244 ( .A1(n9570), .A2(n8821), .ZN(n8760) );
  OAI211_X1 U10245 ( .C1(n8762), .C2(n8823), .A(n8761), .B(n8760), .ZN(
        P1_U3225) );
  XOR2_X1 U10246 ( .A(n8764), .B(n8763), .Z(n8771) );
  NOR2_X1 U10247 ( .A1(n8817), .A2(n8765), .ZN(n8768) );
  NAND2_X1 U10248 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U10249 ( .A1(n8796), .A2(n9139), .ZN(n8766) );
  OAI211_X1 U10250 ( .C1(n8798), .C2(n9694), .A(n9293), .B(n8766), .ZN(n8767)
         );
  AOI211_X1 U10251 ( .C1(n8769), .C2(n8821), .A(n8768), .B(n8767), .ZN(n8770)
         );
  OAI21_X1 U10252 ( .B1(n8771), .B2(n8823), .A(n8770), .ZN(P1_U3226) );
  XOR2_X1 U10253 ( .A(n8772), .B(n8773), .Z(n8780) );
  NOR2_X1 U10254 ( .A1(n8817), .A2(n8774), .ZN(n8777) );
  NAND2_X1 U10255 ( .A1(n8832), .A2(n9140), .ZN(n8775) );
  NAND2_X1 U10256 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9314) );
  OAI211_X1 U10257 ( .C1(n9533), .C2(n8834), .A(n8775), .B(n9314), .ZN(n8776)
         );
  AOI211_X1 U10258 ( .C1(n8778), .C2(n8821), .A(n8777), .B(n8776), .ZN(n8779)
         );
  OAI21_X1 U10259 ( .B1(n8780), .B2(n8823), .A(n8779), .ZN(P1_U3228) );
  AND3_X1 U10260 ( .A1(n8783), .A2(n8782), .A3(n8781), .ZN(n8784) );
  OAI21_X1 U10261 ( .B1(n8785), .B2(n8784), .A(n8830), .ZN(n8791) );
  INV_X1 U10262 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8786) );
  OAI22_X1 U10263 ( .A1(n8834), .A2(n8787), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8786), .ZN(n8789) );
  NOR2_X1 U10264 ( .A1(n8798), .A2(n8809), .ZN(n8788) );
  AOI211_X1 U10265 ( .C1(n8837), .C2(n9443), .A(n8789), .B(n8788), .ZN(n8790)
         );
  OAI211_X1 U10266 ( .C1(n9445), .C2(n8840), .A(n8791), .B(n8790), .ZN(
        P1_U3229) );
  XNOR2_X1 U10267 ( .A(n8793), .B(n8792), .ZN(n8794) );
  XNOR2_X1 U10268 ( .A(n8795), .B(n8794), .ZN(n8802) );
  AOI22_X1 U10269 ( .A1(n9471), .A2(n8796), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n8797) );
  OAI21_X1 U10270 ( .B1(n9507), .B2(n8798), .A(n8797), .ZN(n8800) );
  NOR2_X1 U10271 ( .A1(n9515), .A2(n8840), .ZN(n8799) );
  AOI211_X1 U10272 ( .C1(n8837), .C2(n9512), .A(n8800), .B(n8799), .ZN(n8801)
         );
  OAI21_X1 U10273 ( .B1(n8802), .B2(n8823), .A(n8801), .ZN(P1_U3233) );
  XNOR2_X1 U10274 ( .A(n8804), .B(n8803), .ZN(n8805) );
  XNOR2_X1 U10275 ( .A(n8806), .B(n8805), .ZN(n8812) );
  AOI22_X1 U10276 ( .A1(n9471), .A2(n8832), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8808) );
  NAND2_X1 U10277 ( .A1(n8837), .A2(n9481), .ZN(n8807) );
  OAI211_X1 U10278 ( .C1(n8809), .C2(n8834), .A(n8808), .B(n8807), .ZN(n8810)
         );
  AOI21_X1 U10279 ( .B1(n9584), .B2(n8821), .A(n8810), .ZN(n8811) );
  OAI21_X1 U10280 ( .B1(n8812), .B2(n8823), .A(n8811), .ZN(P1_U3235) );
  NAND2_X1 U10281 ( .A1(n4929), .A2(n8813), .ZN(n8815) );
  XNOR2_X1 U10282 ( .A(n8815), .B(n8814), .ZN(n8824) );
  NOR2_X1 U10283 ( .A1(n8817), .A2(n8816), .ZN(n8820) );
  NAND2_X1 U10284 ( .A1(n8832), .A2(n9139), .ZN(n8818) );
  NAND2_X1 U10285 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9336) );
  OAI211_X1 U10286 ( .C1(n9507), .C2(n8834), .A(n8818), .B(n9336), .ZN(n8819)
         );
  AOI211_X1 U10287 ( .C1(n9608), .C2(n8821), .A(n8820), .B(n8819), .ZN(n8822)
         );
  OAI21_X1 U10288 ( .B1(n8824), .B2(n8823), .A(n8822), .ZN(P1_U3238) );
  OAI21_X1 U10289 ( .B1(n8828), .B2(n8827), .A(n8826), .ZN(n8829) );
  NAND3_X1 U10290 ( .A1(n8831), .A2(n8830), .A3(n8829), .ZN(n8839) );
  AOI22_X1 U10291 ( .A1(n8832), .A2(n9449), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8833) );
  OAI21_X1 U10292 ( .B1(n8835), .B2(n8834), .A(n8833), .ZN(n8836) );
  AOI21_X1 U10293 ( .B1(n9415), .B2(n8837), .A(n8836), .ZN(n8838) );
  OAI211_X1 U10294 ( .C1(n7770), .C2(n8840), .A(n8839), .B(n8838), .ZN(
        P1_U3240) );
  NAND2_X1 U10295 ( .A1(n8842), .A2(n8841), .ZN(n8844) );
  NAND2_X1 U10296 ( .A1(n6066), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U10297 ( .A1(n4520), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n8848) );
  NAND2_X1 U10298 ( .A1(n4521), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n8847) );
  NAND2_X1 U10299 ( .A1(n4517), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8846) );
  NAND3_X1 U10300 ( .A1(n8848), .A2(n8847), .A3(n8846), .ZN(n9133) );
  INV_X1 U10301 ( .A(n9104), .ZN(n8850) );
  INV_X1 U10302 ( .A(n9099), .ZN(n8849) );
  NOR2_X1 U10303 ( .A1(n8850), .A2(n8849), .ZN(n8862) );
  NAND2_X1 U10304 ( .A1(n9072), .A2(n8967), .ZN(n9078) );
  NAND2_X1 U10305 ( .A1(n9446), .A2(n8851), .ZN(n9074) );
  INV_X1 U10306 ( .A(n9090), .ZN(n8852) );
  AOI211_X1 U10307 ( .C1(n9081), .C2(n9078), .A(n9074), .B(n8852), .ZN(n8857)
         );
  OR2_X1 U10308 ( .A1(n9584), .A2(n9495), .ZN(n8853) );
  NAND2_X1 U10309 ( .A1(n9087), .A2(n8853), .ZN(n9084) );
  NAND2_X1 U10310 ( .A1(n9084), .A2(n9446), .ZN(n8854) );
  NAND2_X1 U10311 ( .A1(n9091), .A2(n8854), .ZN(n8855) );
  NAND2_X1 U10312 ( .A1(n8855), .A2(n9090), .ZN(n8856) );
  NAND2_X1 U10313 ( .A1(n9098), .A2(n8856), .ZN(n8860) );
  OAI21_X1 U10314 ( .B1(n8857), .B2(n8860), .A(n9095), .ZN(n8859) );
  NAND2_X1 U10315 ( .A1(n9371), .A2(n8858), .ZN(n9105) );
  AOI21_X1 U10316 ( .B1(n8862), .B2(n8859), .A(n9105), .ZN(n8944) );
  INV_X1 U10317 ( .A(n9096), .ZN(n8863) );
  NAND2_X1 U10318 ( .A1(n9081), .A2(n8969), .ZN(n9071) );
  OAI21_X1 U10319 ( .B1(n8860), .B2(n9071), .A(n9096), .ZN(n8861) );
  AND2_X1 U10320 ( .A1(n8862), .A2(n8861), .ZN(n8943) );
  OAI21_X1 U10321 ( .B1(n8863), .B2(n9505), .A(n8943), .ZN(n8867) );
  NAND2_X1 U10322 ( .A1(n8864), .A2(n8841), .ZN(n8866) );
  NAND2_X1 U10323 ( .A1(n6066), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8865) );
  INV_X1 U10324 ( .A(n9135), .ZN(n8872) );
  NAND2_X1 U10325 ( .A1(n9109), .A2(n9103), .ZN(n8917) );
  AOI21_X1 U10326 ( .B1(n8944), .B2(n8867), .A(n8917), .ZN(n8873) );
  NAND2_X1 U10327 ( .A1(n8868), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U10328 ( .A1(n4521), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U10329 ( .A1(n4517), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8869) );
  AND3_X1 U10330 ( .A1(n8871), .A2(n8870), .A3(n8869), .ZN(n9375) );
  NAND2_X1 U10331 ( .A1(n9359), .A2(n9375), .ZN(n8878) );
  NAND2_X1 U10332 ( .A1(n9549), .A2(n8872), .ZN(n9110) );
  NAND2_X1 U10333 ( .A1(n8878), .A2(n9110), .ZN(n8947) );
  INV_X1 U10334 ( .A(n9375), .ZN(n9134) );
  NAND2_X1 U10335 ( .A1(n9133), .A2(n9134), .ZN(n9113) );
  OAI22_X1 U10336 ( .A1(n8873), .A2(n8947), .B1(n9359), .B2(n9113), .ZN(n8877)
         );
  NAND2_X1 U10337 ( .A1(n8874), .A2(n8841), .ZN(n8876) );
  NAND2_X1 U10338 ( .A1(n6066), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8875) );
  AND2_X1 U10339 ( .A1(n9362), .A2(n9133), .ZN(n9119) );
  INV_X1 U10340 ( .A(n9119), .ZN(n9114) );
  OAI211_X1 U10341 ( .C1(n9547), .C2(n9133), .A(n8877), .B(n9114), .ZN(n8911)
         );
  NAND2_X1 U10342 ( .A1(n6726), .A2(n4510), .ZN(n8957) );
  OR2_X1 U10343 ( .A1(n9359), .A2(n9375), .ZN(n8950) );
  NAND2_X1 U10344 ( .A1(n8950), .A2(n8878), .ZN(n8910) );
  NAND2_X1 U10345 ( .A1(n9109), .A2(n9110), .ZN(n9383) );
  INV_X1 U10346 ( .A(n8879), .ZN(n8888) );
  NAND4_X1 U10347 ( .A1(n8883), .A2(n8882), .A3(n8881), .A4(n8880), .ZN(n8886)
         );
  NOR3_X1 U10348 ( .A1(n8886), .A2(n8885), .A3(n8884), .ZN(n8887) );
  NAND4_X1 U10349 ( .A1(n8890), .A2(n8889), .A3(n8888), .A4(n8887), .ZN(n8891)
         );
  NOR2_X1 U10350 ( .A1(n8891), .A2(n8918), .ZN(n8892) );
  NAND4_X1 U10351 ( .A1(n8895), .A2(n8894), .A3(n8893), .A4(n8892), .ZN(n8896)
         );
  NOR2_X1 U10352 ( .A1(n8896), .A2(n9687), .ZN(n8897) );
  NAND4_X1 U10353 ( .A1(n8900), .A2(n8899), .A3(n8898), .A4(n8897), .ZN(n8901)
         );
  NOR2_X1 U10354 ( .A1(n8902), .A2(n8901), .ZN(n8903) );
  NAND3_X1 U10355 ( .A1(n9504), .A2(n9529), .A3(n8903), .ZN(n8904) );
  NOR2_X1 U10356 ( .A1(n9492), .A2(n8904), .ZN(n8905) );
  NAND3_X1 U10357 ( .A1(n9460), .A2(n8905), .A3(n9474), .ZN(n8906) );
  OR3_X1 U10358 ( .A1(n9425), .A2(n8906), .A3(n9448), .ZN(n8908) );
  NOR4_X1 U10359 ( .A1(n9119), .A2(n8910), .A3(n9383), .A4(n8909), .ZN(n8913)
         );
  AOI211_X1 U10360 ( .C1(n8912), .C2(n8911), .A(n8957), .B(n8913), .ZN(n8961)
         );
  INV_X1 U10361 ( .A(n9133), .ZN(n9361) );
  NAND2_X1 U10362 ( .A1(n9539), .A2(n9361), .ZN(n9122) );
  NOR2_X1 U10363 ( .A1(n6726), .A2(n4510), .ZN(n8956) );
  INV_X1 U10364 ( .A(n8917), .ZN(n8949) );
  NAND2_X1 U10365 ( .A1(n9047), .A2(n9044), .ZN(n9035) );
  INV_X1 U10366 ( .A(n8918), .ZN(n8931) );
  INV_X1 U10367 ( .A(n8973), .ZN(n8922) );
  OAI211_X1 U10368 ( .C1(n4509), .C2(n6016), .A(n8920), .B(n8919), .ZN(n8921)
         );
  NAND2_X1 U10369 ( .A1(n8974), .A2(n8991), .ZN(n8971) );
  AOI21_X1 U10370 ( .B1(n8922), .B2(n8921), .A(n8971), .ZN(n8923) );
  INV_X1 U10371 ( .A(n8923), .ZN(n8925) );
  INV_X1 U10372 ( .A(n8983), .ZN(n8924) );
  AOI21_X1 U10373 ( .B1(n8925), .B2(n8982), .A(n8924), .ZN(n8927) );
  NAND2_X1 U10374 ( .A1(n8984), .A2(n8926), .ZN(n8992) );
  OAI21_X1 U10375 ( .B1(n8927), .B2(n8992), .A(n8997), .ZN(n8930) );
  INV_X1 U10376 ( .A(n9014), .ZN(n9020) );
  INV_X1 U10377 ( .A(n8928), .ZN(n8929) );
  AOI211_X1 U10378 ( .C1(n8931), .C2(n8930), .A(n9020), .B(n8929), .ZN(n8932)
         );
  NAND2_X1 U10379 ( .A1(n9017), .A2(n9012), .ZN(n9025) );
  NOR2_X1 U10380 ( .A1(n8932), .A2(n9025), .ZN(n8934) );
  NAND2_X1 U10381 ( .A1(n8933), .A2(n9015), .ZN(n9023) );
  OAI211_X1 U10382 ( .C1(n8934), .C2(n9023), .A(n9018), .B(n9043), .ZN(n8937)
         );
  AND2_X1 U10383 ( .A1(n9045), .A2(n9041), .ZN(n8935) );
  OR2_X1 U10384 ( .A1(n9035), .A2(n8935), .ZN(n8936) );
  AND2_X1 U10385 ( .A1(n8936), .A2(n9046), .ZN(n9037) );
  OAI21_X1 U10386 ( .B1(n9035), .B2(n8937), .A(n9037), .ZN(n8939) );
  INV_X1 U10387 ( .A(n9050), .ZN(n9039) );
  NAND2_X1 U10388 ( .A1(n9527), .A2(n8938), .ZN(n9056) );
  AOI211_X1 U10389 ( .C1(n9048), .C2(n8939), .A(n9039), .B(n9056), .ZN(n8941)
         );
  NAND2_X1 U10390 ( .A1(n9057), .A2(n8940), .ZN(n9061) );
  OAI21_X1 U10391 ( .B1(n8941), .B2(n9061), .A(n9062), .ZN(n8942) );
  AND3_X1 U10392 ( .A1(n9096), .A2(n9058), .A3(n8942), .ZN(n8946) );
  INV_X1 U10393 ( .A(n8943), .ZN(n8945) );
  OAI21_X1 U10394 ( .B1(n8946), .B2(n8945), .A(n8944), .ZN(n8948) );
  AOI21_X1 U10395 ( .B1(n8949), .B2(n8948), .A(n8947), .ZN(n8952) );
  INV_X1 U10396 ( .A(n8950), .ZN(n8951) );
  OAI21_X1 U10397 ( .B1(n8952), .B2(n8951), .A(n9114), .ZN(n8953) );
  NAND2_X1 U10398 ( .A1(n8953), .A2(n9122), .ZN(n8954) );
  MUX2_X1 U10399 ( .A(n8956), .B(n8955), .S(n8954), .Z(n8959) );
  OAI22_X1 U10400 ( .A1(n9122), .A2(n8957), .B1(n9116), .B2(n9118), .ZN(n8958)
         );
  NOR4_X1 U10401 ( .A1(n8961), .A2(n8960), .A3(n8959), .A4(n8958), .ZN(n9126)
         );
  INV_X1 U10402 ( .A(n9383), .ZN(n9374) );
  INV_X1 U10403 ( .A(n9095), .ZN(n8962) );
  NAND2_X1 U10404 ( .A1(n9099), .A2(n8962), .ZN(n8963) );
  NAND3_X1 U10405 ( .A1(n8963), .A2(n9116), .A3(n9096), .ZN(n8966) );
  NAND2_X1 U10406 ( .A1(n9105), .A2(n4644), .ZN(n8965) );
  NAND3_X1 U10407 ( .A1(n9104), .A2(n4644), .A3(n9099), .ZN(n8964) );
  OAI211_X1 U10408 ( .C1(n9105), .C2(n8966), .A(n8965), .B(n8964), .ZN(n9102)
         );
  NAND2_X1 U10409 ( .A1(n8967), .A2(n4742), .ZN(n8968) );
  NAND2_X1 U10410 ( .A1(n8968), .A2(n9116), .ZN(n8970) );
  NAND2_X1 U10411 ( .A1(n8970), .A2(n8969), .ZN(n9069) );
  INV_X1 U10412 ( .A(n8971), .ZN(n8972) );
  NAND2_X1 U10413 ( .A1(n8973), .A2(n8972), .ZN(n8979) );
  NAND2_X1 U10414 ( .A1(n8975), .A2(n8974), .ZN(n8977) );
  NAND3_X1 U10415 ( .A1(n8977), .A2(n8982), .A3(n8976), .ZN(n8978) );
  MUX2_X1 U10416 ( .A(n8979), .B(n8978), .S(n9116), .Z(n8981) );
  NAND2_X1 U10417 ( .A1(n8986), .A2(n9000), .ZN(n8990) );
  INV_X1 U10418 ( .A(n8987), .ZN(n8988) );
  INV_X1 U10419 ( .A(n8991), .ZN(n8994) );
  INV_X1 U10420 ( .A(n8992), .ZN(n8993) );
  OAI21_X1 U10421 ( .B1(n8995), .B2(n8994), .A(n8993), .ZN(n8998) );
  AOI21_X1 U10422 ( .B1(n8998), .B2(n8997), .A(n8996), .ZN(n9004) );
  NAND2_X1 U10423 ( .A1(n9000), .A2(n8999), .ZN(n9003) );
  INV_X1 U10424 ( .A(n9001), .ZN(n9002) );
  OAI21_X1 U10425 ( .B1(n9004), .B2(n9003), .A(n9002), .ZN(n9005) );
  INV_X1 U10426 ( .A(n9006), .ZN(n9007) );
  MUX2_X1 U10427 ( .A(n9008), .B(n9007), .S(n9116), .Z(n9009) );
  INV_X1 U10428 ( .A(n9021), .ZN(n9011) );
  NAND2_X1 U10429 ( .A1(n9013), .A2(n9012), .ZN(n9016) );
  NAND3_X1 U10430 ( .A1(n9016), .A2(n9015), .A3(n9014), .ZN(n9019) );
  NAND4_X1 U10431 ( .A1(n9019), .A2(n4644), .A3(n9018), .A4(n9017), .ZN(n9034)
         );
  AOI21_X1 U10432 ( .B1(n9022), .B2(n9021), .A(n9020), .ZN(n9026) );
  INV_X1 U10433 ( .A(n9023), .ZN(n9024) );
  OAI211_X1 U10434 ( .C1(n9026), .C2(n9025), .A(n9024), .B(n9116), .ZN(n9033)
         );
  NOR2_X1 U10435 ( .A1(n9027), .A2(n9116), .ZN(n9030) );
  NAND2_X1 U10436 ( .A1(n9027), .A2(n9116), .ZN(n9028) );
  NAND2_X1 U10437 ( .A1(n9031), .A2(n9028), .ZN(n9029) );
  OAI21_X1 U10438 ( .B1(n9031), .B2(n9030), .A(n9029), .ZN(n9032) );
  NAND3_X1 U10439 ( .A1(n9034), .A2(n9033), .A3(n9032), .ZN(n9042) );
  INV_X1 U10440 ( .A(n9035), .ZN(n9036) );
  NAND3_X1 U10441 ( .A1(n9042), .A2(n9036), .A3(n9043), .ZN(n9038) );
  NAND2_X1 U10442 ( .A1(n9038), .A2(n9037), .ZN(n9040) );
  AOI21_X1 U10443 ( .B1(n9040), .B2(n9048), .A(n9039), .ZN(n9053) );
  INV_X1 U10444 ( .A(n9048), .ZN(n9049) );
  AOI21_X1 U10445 ( .B1(n9051), .B2(n9050), .A(n9049), .ZN(n9052) );
  MUX2_X1 U10446 ( .A(n9053), .B(n9052), .S(n9116), .Z(n9055) );
  OR2_X1 U10447 ( .A1(n9055), .A2(n9054), .ZN(n9065) );
  INV_X1 U10448 ( .A(n9056), .ZN(n9060) );
  NAND2_X1 U10449 ( .A1(n9058), .A2(n9057), .ZN(n9059) );
  INV_X1 U10450 ( .A(n9061), .ZN(n9064) );
  INV_X1 U10451 ( .A(n9062), .ZN(n9063) );
  INV_X1 U10452 ( .A(n9066), .ZN(n9068) );
  OAI22_X1 U10453 ( .A1(n9069), .A2(n9068), .B1(n4644), .B2(n9067), .ZN(n9070)
         );
  INV_X1 U10454 ( .A(n9071), .ZN(n9073) );
  AOI21_X1 U10455 ( .B1(n9080), .B2(n9073), .A(n4752), .ZN(n9077) );
  INV_X1 U10456 ( .A(n9474), .ZN(n9076) );
  INV_X1 U10457 ( .A(n9074), .ZN(n9075) );
  OAI21_X1 U10458 ( .B1(n9077), .B2(n9076), .A(n9075), .ZN(n9086) );
  INV_X1 U10459 ( .A(n9078), .ZN(n9079) );
  NAND2_X1 U10460 ( .A1(n9080), .A2(n9079), .ZN(n9082) );
  NAND2_X1 U10461 ( .A1(n9082), .A2(n9081), .ZN(n9083) );
  NOR2_X1 U10462 ( .A1(n9087), .A2(n4644), .ZN(n9088) );
  NOR2_X1 U10463 ( .A1(n9448), .A2(n9088), .ZN(n9089) );
  MUX2_X1 U10464 ( .A(n9091), .B(n9090), .S(n9116), .Z(n9092) );
  NAND2_X1 U10465 ( .A1(n9093), .A2(n9092), .ZN(n9100) );
  INV_X1 U10466 ( .A(n9098), .ZN(n9094) );
  NAND3_X1 U10467 ( .A1(n9096), .A2(n4644), .A3(n9095), .ZN(n9097) );
  NAND4_X1 U10468 ( .A1(n9100), .A2(n9116), .A3(n9099), .A4(n9098), .ZN(n9101)
         );
  OAI21_X1 U10469 ( .B1(n9105), .B2(n9104), .A(n9103), .ZN(n9106) );
  NAND2_X1 U10470 ( .A1(n9106), .A2(n9116), .ZN(n9107) );
  NAND2_X1 U10471 ( .A1(n9374), .A2(n9108), .ZN(n9112) );
  MUX2_X1 U10472 ( .A(n9110), .B(n9109), .S(n9116), .Z(n9111) );
  NAND2_X1 U10473 ( .A1(n9112), .A2(n9111), .ZN(n9115) );
  INV_X1 U10474 ( .A(n9118), .ZN(n9117) );
  NAND3_X1 U10475 ( .A1(n9120), .A2(n9357), .A3(n9117), .ZN(n9125) );
  INV_X1 U10476 ( .A(n6525), .ZN(n9129) );
  AOI211_X1 U10477 ( .C1(n9119), .C2(n9357), .A(n9129), .B(n9118), .ZN(n9124)
         );
  OAI21_X1 U10478 ( .B1(n9122), .B2(n6726), .A(n9121), .ZN(n9123) );
  NAND2_X1 U10479 ( .A1(n9127), .A2(n9176), .ZN(n9128) );
  OAI211_X1 U10480 ( .C1(n9129), .C2(n9131), .A(n9128), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9130) );
  OAI21_X1 U10481 ( .B1(n9132), .B2(n9131), .A(n9130), .ZN(P1_U3242) );
  MUX2_X1 U10482 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9133), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10483 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9134), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10484 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9135), .S(P1_U3973), .Z(
        P1_U3583) );
  INV_X1 U10485 ( .A(n9379), .ZN(n9398) );
  MUX2_X1 U10486 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9398), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10487 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9420), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10488 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9434), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10489 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9449), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10490 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9461), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10491 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9470), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10492 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9462), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10493 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9471), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10494 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9136), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10495 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9137), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10496 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9138), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10497 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9139), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10498 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9140), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10499 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n5016), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10500 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9141), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10501 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9142), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10502 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9143), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10503 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9144), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10504 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9145), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10505 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9709), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10506 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9146), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10507 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9710), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10508 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9147), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10509 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9148), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10510 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9149), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10511 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9150), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10512 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9151), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10513 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9152), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10514 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6032), .S(P1_U3973), .Z(
        P1_U3554) );
  AOI211_X1 U10515 ( .C1(n9174), .C2(n9154), .A(n9153), .B(n9672), .ZN(n9155)
         );
  INV_X1 U10516 ( .A(n9155), .ZN(n9164) );
  INV_X1 U10517 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10066) );
  OAI22_X1 U10518 ( .A1(n9338), .A2(n10066), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9156), .ZN(n9157) );
  AOI21_X1 U10519 ( .B1(n9677), .B2(n9158), .A(n9157), .ZN(n9163) );
  OAI211_X1 U10520 ( .C1(n9161), .C2(n9160), .A(n9679), .B(n9159), .ZN(n9162)
         );
  NAND3_X1 U10521 ( .A1(n9164), .A2(n9163), .A3(n9162), .ZN(P1_U3244) );
  AOI211_X1 U10522 ( .C1(n9167), .C2(n9166), .A(n9165), .B(n9672), .ZN(n9171)
         );
  AOI211_X1 U10523 ( .C1(n9169), .C2(n9168), .A(n9191), .B(n9351), .ZN(n9170)
         );
  NOR2_X1 U10524 ( .A1(n9171), .A2(n9170), .ZN(n9182) );
  AOI22_X1 U10525 ( .A1(n9675), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9181) );
  NAND3_X1 U10526 ( .A1(n9172), .A2(n9173), .A3(n4522), .ZN(n9178) );
  OAI21_X1 U10527 ( .B1(n4522), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9173), .ZN(
        n9661) );
  INV_X1 U10528 ( .A(n9174), .ZN(n9175) );
  AOI22_X1 U10529 ( .A1(n10239), .A2(n9661), .B1(n9176), .B2(n9175), .ZN(n9177) );
  NAND3_X1 U10530 ( .A1(n9178), .A2(P1_U3973), .A3(n9177), .ZN(n9684) );
  NAND2_X1 U10531 ( .A1(n9677), .A2(n9179), .ZN(n9180) );
  NAND4_X1 U10532 ( .A1(n9182), .A2(n9181), .A3(n9684), .A4(n9180), .ZN(
        P1_U3245) );
  OAI211_X1 U10533 ( .C1(n9185), .C2(n9184), .A(n9327), .B(n9183), .ZN(n9197)
         );
  MUX2_X1 U10534 ( .A(n9840), .B(P1_REG1_REG_3__SCAN_IN), .S(n9193), .Z(n9188)
         );
  INV_X1 U10535 ( .A(n9186), .ZN(n9187) );
  NAND2_X1 U10536 ( .A1(n9188), .A2(n9187), .ZN(n9190) );
  OAI211_X1 U10537 ( .C1(n9191), .C2(n9190), .A(n9679), .B(n9189), .ZN(n9196)
         );
  AOI21_X1 U10538 ( .B1(n9675), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n9192), .ZN(
        n9195) );
  NAND2_X1 U10539 ( .A1(n9677), .A2(n9193), .ZN(n9194) );
  NAND4_X1 U10540 ( .A1(n9197), .A2(n9196), .A3(n9195), .A4(n9194), .ZN(
        P1_U3246) );
  NOR2_X1 U10541 ( .A1(n9354), .A2(n9198), .ZN(n9199) );
  AOI211_X1 U10542 ( .C1(n9675), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9200), .B(
        n9199), .ZN(n9210) );
  AOI211_X1 U10543 ( .C1(n9203), .C2(n9202), .A(n9201), .B(n9672), .ZN(n9204)
         );
  INV_X1 U10544 ( .A(n9204), .ZN(n9209) );
  OAI211_X1 U10545 ( .C1(n9207), .C2(n9206), .A(n9679), .B(n9205), .ZN(n9208)
         );
  NAND3_X1 U10546 ( .A1(n9210), .A2(n9209), .A3(n9208), .ZN(P1_U3248) );
  NOR2_X1 U10547 ( .A1(n9354), .A2(n9211), .ZN(n9212) );
  AOI211_X1 U10548 ( .C1(n9675), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9213), .B(
        n9212), .ZN(n9223) );
  AOI211_X1 U10549 ( .C1(n9216), .C2(n9215), .A(n9214), .B(n9672), .ZN(n9217)
         );
  INV_X1 U10550 ( .A(n9217), .ZN(n9222) );
  OAI211_X1 U10551 ( .C1(n9220), .C2(n9219), .A(n9679), .B(n9218), .ZN(n9221)
         );
  NAND3_X1 U10552 ( .A1(n9223), .A2(n9222), .A3(n9221), .ZN(P1_U3249) );
  NOR2_X1 U10553 ( .A1(n9354), .A2(n9224), .ZN(n9225) );
  AOI211_X1 U10554 ( .C1(n9675), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n9226), .B(
        n9225), .ZN(n9236) );
  AOI211_X1 U10555 ( .C1(n9229), .C2(n9228), .A(n9227), .B(n9672), .ZN(n9230)
         );
  INV_X1 U10556 ( .A(n9230), .ZN(n9235) );
  OAI211_X1 U10557 ( .C1(n9233), .C2(n9232), .A(n9679), .B(n9231), .ZN(n9234)
         );
  NAND3_X1 U10558 ( .A1(n9236), .A2(n9235), .A3(n9234), .ZN(P1_U3250) );
  NOR2_X1 U10559 ( .A1(n9354), .A2(n9237), .ZN(n9238) );
  AOI211_X1 U10560 ( .C1(n9675), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9239), .B(
        n9238), .ZN(n9249) );
  AOI211_X1 U10561 ( .C1(n9242), .C2(n9241), .A(n9240), .B(n9672), .ZN(n9243)
         );
  INV_X1 U10562 ( .A(n9243), .ZN(n9248) );
  OAI211_X1 U10563 ( .C1(n9246), .C2(n9245), .A(n9679), .B(n9244), .ZN(n9247)
         );
  NAND3_X1 U10564 ( .A1(n9249), .A2(n9248), .A3(n9247), .ZN(P1_U3251) );
  NOR2_X1 U10565 ( .A1(n9354), .A2(n9272), .ZN(n9250) );
  AOI211_X1 U10566 ( .C1(n9675), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n9251), .B(
        n9250), .ZN(n9266) );
  OR2_X1 U10567 ( .A1(n9268), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9253) );
  NAND2_X1 U10568 ( .A1(n9268), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9252) );
  AND2_X1 U10569 ( .A1(n9253), .A2(n9252), .ZN(n9257) );
  OAI21_X1 U10570 ( .B1(n9255), .B2(n7225), .A(n9254), .ZN(n9256) );
  NAND2_X1 U10571 ( .A1(n9257), .A2(n9256), .ZN(n9271) );
  OAI211_X1 U10572 ( .C1(n9257), .C2(n9256), .A(n9679), .B(n9271), .ZN(n9265)
         );
  NAND2_X1 U10573 ( .A1(n9268), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9258) );
  OAI21_X1 U10574 ( .B1(n9268), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9258), .ZN(
        n9262) );
  AOI211_X1 U10575 ( .C1(n9262), .C2(n9261), .A(n9267), .B(n9672), .ZN(n9263)
         );
  INV_X1 U10576 ( .A(n9263), .ZN(n9264) );
  NAND3_X1 U10577 ( .A1(n9266), .A2(n9265), .A3(n9264), .ZN(P1_U3257) );
  INV_X1 U10578 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9269) );
  NOR2_X1 U10579 ( .A1(n9269), .A2(n9270), .ZN(n9288) );
  AOI211_X1 U10580 ( .C1(n9270), .C2(n9269), .A(n9288), .B(n9672), .ZN(n9279)
         );
  INV_X1 U10581 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9861) );
  OAI21_X1 U10582 ( .B1(n9861), .B2(n9272), .A(n9271), .ZN(n9280) );
  XNOR2_X1 U10583 ( .A(n4712), .B(n9280), .ZN(n9273) );
  NAND2_X1 U10584 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9273), .ZN(n9282) );
  OAI211_X1 U10585 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9273), .A(n9679), .B(
        n9282), .ZN(n9277) );
  INV_X1 U10586 ( .A(n9274), .ZN(n9275) );
  AOI21_X1 U10587 ( .B1(n9675), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9275), .ZN(
        n9276) );
  OAI211_X1 U10588 ( .C1(n9354), .C2(n4712), .A(n9277), .B(n9276), .ZN(n9278)
         );
  OR2_X1 U10589 ( .A1(n9279), .A2(n9278), .ZN(P1_U3258) );
  NAND2_X1 U10590 ( .A1(n9281), .A2(n9280), .ZN(n9283) );
  NAND2_X1 U10591 ( .A1(n9283), .A2(n9282), .ZN(n9286) );
  INV_X1 U10592 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9649) );
  NOR2_X1 U10593 ( .A1(n9311), .A2(n9649), .ZN(n9284) );
  AOI21_X1 U10594 ( .B1(n9311), .B2(n9649), .A(n9284), .ZN(n9285) );
  NOR2_X1 U10595 ( .A1(n9285), .A2(n9286), .ZN(n9302) );
  AOI21_X1 U10596 ( .B1(n9286), .B2(n9285), .A(n9302), .ZN(n9298) );
  NOR2_X1 U10597 ( .A1(n9287), .A2(n4712), .ZN(n9289) );
  AOI22_X1 U10598 ( .A1(n9311), .A2(n7603), .B1(P1_REG2_REG_16__SCAN_IN), .B2(
        n9303), .ZN(n9290) );
  AOI211_X1 U10599 ( .C1(n9291), .C2(n9290), .A(n9310), .B(n9672), .ZN(n9292)
         );
  INV_X1 U10600 ( .A(n9292), .ZN(n9297) );
  INV_X1 U10601 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9294) );
  OAI21_X1 U10602 ( .B1(n9338), .B2(n9294), .A(n9293), .ZN(n9295) );
  AOI21_X1 U10603 ( .B1(n9677), .B2(n9311), .A(n9295), .ZN(n9296) );
  OAI211_X1 U10604 ( .C1(n9298), .C2(n9351), .A(n9297), .B(n9296), .ZN(
        P1_U3259) );
  INV_X1 U10605 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9299) );
  OR2_X1 U10606 ( .A1(n9330), .A2(n9299), .ZN(n9301) );
  NAND2_X1 U10607 ( .A1(n9330), .A2(n9299), .ZN(n9300) );
  NAND2_X1 U10608 ( .A1(n9301), .A2(n9300), .ZN(n9306) );
  AOI21_X1 U10609 ( .B1(n9303), .B2(n9649), .A(n9302), .ZN(n9304) );
  INV_X1 U10610 ( .A(n9304), .ZN(n9305) );
  NAND2_X1 U10611 ( .A1(n9306), .A2(n9305), .ZN(n9332) );
  OAI21_X1 U10612 ( .B1(n9306), .B2(n9305), .A(n9332), .ZN(n9307) );
  AOI22_X1 U10613 ( .A1(n9679), .A2(n9307), .B1(n9677), .B2(n9330), .ZN(n9318)
         );
  NOR2_X1 U10614 ( .A1(n9309), .A2(n9321), .ZN(n9308) );
  AOI21_X1 U10615 ( .B1(n9321), .B2(n9309), .A(n9308), .ZN(n9313) );
  NAND2_X1 U10616 ( .A1(n9320), .A2(n9313), .ZN(n9312) );
  OAI21_X1 U10617 ( .B1(n9313), .B2(n9320), .A(n9312), .ZN(n9316) );
  INV_X1 U10618 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10119) );
  OAI21_X1 U10619 ( .B1(n9338), .B2(n10119), .A(n9314), .ZN(n9315) );
  AOI21_X1 U10620 ( .B1(n9327), .B2(n9316), .A(n9315), .ZN(n9317) );
  NAND2_X1 U10621 ( .A1(n9318), .A2(n9317), .ZN(P1_U3260) );
  OR2_X1 U10622 ( .A1(n9330), .A2(n9319), .ZN(n9323) );
  NAND2_X1 U10623 ( .A1(n9321), .A2(n9320), .ZN(n9322) );
  OR2_X1 U10624 ( .A1(n9347), .A2(n9324), .ZN(n9326) );
  NAND2_X1 U10625 ( .A1(n9347), .A2(n9324), .ZN(n9325) );
  NAND2_X1 U10626 ( .A1(n9326), .A2(n9325), .ZN(n9328) );
  NAND2_X1 U10627 ( .A1(n9328), .A2(n9329), .ZN(n9345) );
  OAI211_X1 U10628 ( .C1(n9329), .C2(n9328), .A(n9327), .B(n9345), .ZN(n9342)
         );
  XNOR2_X1 U10629 ( .A(n9347), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9334) );
  OR2_X1 U10630 ( .A1(n9330), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9331) );
  NAND2_X1 U10631 ( .A1(n9332), .A2(n9331), .ZN(n9333) );
  OR2_X1 U10632 ( .A1(n9334), .A2(n9333), .ZN(n9349) );
  NAND2_X1 U10633 ( .A1(n9334), .A2(n9333), .ZN(n9335) );
  NAND3_X1 U10634 ( .A1(n9679), .A2(n9349), .A3(n9335), .ZN(n9341) );
  INV_X1 U10635 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9337) );
  OAI21_X1 U10636 ( .B1(n9338), .B2(n9337), .A(n9336), .ZN(n9339) );
  AOI21_X1 U10637 ( .B1(n9677), .B2(n9347), .A(n9339), .ZN(n9340) );
  NAND3_X1 U10638 ( .A1(n9342), .A2(n9341), .A3(n9340), .ZN(P1_U3261) );
  INV_X1 U10639 ( .A(n9343), .ZN(n9358) );
  NAND2_X1 U10640 ( .A1(n9347), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9344) );
  NAND2_X1 U10641 ( .A1(n9345), .A2(n9344), .ZN(n9346) );
  XNOR2_X1 U10642 ( .A(n9346), .B(n9524), .ZN(n9356) );
  INV_X1 U10643 ( .A(n9356), .ZN(n9352) );
  NAND2_X1 U10644 ( .A1(n9347), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9348) );
  NAND2_X1 U10645 ( .A1(n9349), .A2(n9348), .ZN(n9350) );
  XNOR2_X1 U10646 ( .A(n9350), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9353) );
  NAND2_X1 U10647 ( .A1(n9679), .A2(n9353), .ZN(n9355) );
  XNOR2_X1 U10648 ( .A(n9362), .B(n9366), .ZN(n9542) );
  INV_X1 U10649 ( .A(P1_B_REG_SCAN_IN), .ZN(n9360) );
  OAI21_X1 U10650 ( .B1(n4522), .B2(n9360), .A(n9708), .ZN(n9376) );
  NOR2_X1 U10651 ( .A1(n9376), .A2(n9361), .ZN(n9538) );
  INV_X1 U10652 ( .A(n9538), .ZN(n9545) );
  NOR2_X1 U10653 ( .A1(n9730), .A2(n9545), .ZN(n9369) );
  NOR2_X1 U10654 ( .A1(n9362), .A2(n9521), .ZN(n9363) );
  AOI211_X1 U10655 ( .C1(n9730), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9369), .B(
        n9363), .ZN(n9364) );
  OAI21_X1 U10656 ( .B1(n9542), .B2(n9365), .A(n9364), .ZN(P1_U3263) );
  OAI211_X1 U10657 ( .C1(n9547), .C2(n4734), .A(n9367), .B(n9722), .ZN(n9546)
         );
  NOR2_X1 U10658 ( .A1(n9547), .A2(n9521), .ZN(n9368) );
  AOI211_X1 U10659 ( .C1(n9730), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9369), .B(
        n9368), .ZN(n9370) );
  OAI21_X1 U10660 ( .B1(n9484), .B2(n9546), .A(n9370), .ZN(P1_U3264) );
  NAND2_X1 U10661 ( .A1(n9372), .A2(n9371), .ZN(n9373) );
  XNOR2_X1 U10662 ( .A(n9374), .B(n9373), .ZN(n9378) );
  OAI22_X1 U10663 ( .A1(n9376), .A2(n9375), .B1(n9379), .B2(n9691), .ZN(n9377)
         );
  AOI21_X1 U10664 ( .B1(n9378), .B2(n9491), .A(n9377), .ZN(n9551) );
  NAND2_X1 U10665 ( .A1(n9554), .A2(n9398), .ZN(n9381) );
  INV_X1 U10666 ( .A(n9552), .ZN(n9393) );
  INV_X1 U10667 ( .A(n9549), .ZN(n9391) );
  AOI21_X1 U10668 ( .B1(n9549), .B2(n9385), .A(n9541), .ZN(n9387) );
  NAND2_X1 U10669 ( .A1(n9548), .A2(n9726), .ZN(n9390) );
  AOI22_X1 U10670 ( .A1(n9730), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9388), .B2(
        n9718), .ZN(n9389) );
  OAI211_X1 U10671 ( .C1(n9391), .C2(n9521), .A(n9390), .B(n9389), .ZN(n9392)
         );
  AOI21_X1 U10672 ( .B1(n9393), .B2(n9486), .A(n9392), .ZN(n9394) );
  OAI21_X1 U10673 ( .B1(n9551), .B2(n9730), .A(n9394), .ZN(P1_U3356) );
  OAI21_X1 U10674 ( .B1(n9397), .B2(n9396), .A(n9395), .ZN(n9399) );
  AOI222_X1 U10675 ( .A1(n9491), .A2(n9399), .B1(n9398), .B2(n9708), .C1(n9434), .C2(n9711), .ZN(n9562) );
  OAI21_X1 U10676 ( .B1(n9402), .B2(n9401), .A(n9400), .ZN(n9558) );
  AOI211_X1 U10677 ( .C1(n9560), .C2(n9413), .A(n9541), .B(n9403), .ZN(n9559)
         );
  NAND2_X1 U10678 ( .A1(n9559), .A2(n9726), .ZN(n9406) );
  AOI22_X1 U10679 ( .A1(n9730), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9404), .B2(
        n9718), .ZN(n9405) );
  OAI211_X1 U10680 ( .C1(n9407), .C2(n9521), .A(n9406), .B(n9405), .ZN(n9408)
         );
  AOI21_X1 U10681 ( .B1(n9558), .B2(n9486), .A(n9408), .ZN(n9409) );
  OAI21_X1 U10682 ( .B1(n9730), .B2(n9562), .A(n9409), .ZN(P1_U3266) );
  XNOR2_X1 U10683 ( .A(n9411), .B(n9410), .ZN(n9568) );
  INV_X1 U10684 ( .A(n9413), .ZN(n9414) );
  AOI211_X1 U10685 ( .C1(n9565), .C2(n9427), .A(n9541), .B(n9414), .ZN(n9564)
         );
  AOI22_X1 U10686 ( .A1(n9730), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9415), .B2(
        n9718), .ZN(n9416) );
  OAI21_X1 U10687 ( .B1(n7770), .B2(n9521), .A(n9416), .ZN(n9423) );
  OAI21_X1 U10688 ( .B1(n9419), .B2(n9418), .A(n9417), .ZN(n9421) );
  AOI222_X1 U10689 ( .A1(n9491), .A2(n9421), .B1(n9420), .B2(n9708), .C1(n9449), .C2(n9711), .ZN(n9567) );
  NOR2_X1 U10690 ( .A1(n9567), .A2(n9730), .ZN(n9422) );
  AOI211_X1 U10691 ( .C1(n9564), .C2(n9726), .A(n9423), .B(n9422), .ZN(n9424)
         );
  OAI21_X1 U10692 ( .B1(n9568), .B2(n9537), .A(n9424), .ZN(P1_U3267) );
  XNOR2_X1 U10693 ( .A(n9426), .B(n9425), .ZN(n9573) );
  AOI211_X1 U10694 ( .C1(n9570), .C2(n9440), .A(n9541), .B(n9412), .ZN(n9569)
         );
  AOI22_X1 U10695 ( .A1(n9730), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9428), .B2(
        n9718), .ZN(n9429) );
  OAI21_X1 U10696 ( .B1(n9430), .B2(n9521), .A(n9429), .ZN(n9437) );
  OAI21_X1 U10697 ( .B1(n9433), .B2(n9432), .A(n9431), .ZN(n9435) );
  AOI222_X1 U10698 ( .A1(n9491), .A2(n9435), .B1(n9434), .B2(n9708), .C1(n9461), .C2(n9711), .ZN(n9572) );
  NOR2_X1 U10699 ( .A1(n9572), .A2(n9730), .ZN(n9436) );
  AOI211_X1 U10700 ( .C1(n9569), .C2(n9726), .A(n9437), .B(n9436), .ZN(n9438)
         );
  OAI21_X1 U10701 ( .B1(n9573), .B2(n9537), .A(n9438), .ZN(P1_U3268) );
  XNOR2_X1 U10702 ( .A(n9439), .B(n9448), .ZN(n9578) );
  INV_X1 U10703 ( .A(n9454), .ZN(n9442) );
  INV_X1 U10704 ( .A(n9440), .ZN(n9441) );
  AOI211_X1 U10705 ( .C1(n9575), .C2(n9442), .A(n9541), .B(n9441), .ZN(n9574)
         );
  AOI22_X1 U10706 ( .A1(n9730), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9443), .B2(
        n9718), .ZN(n9444) );
  OAI21_X1 U10707 ( .B1(n9445), .B2(n9521), .A(n9444), .ZN(n9452) );
  NAND2_X1 U10708 ( .A1(n9458), .A2(n9446), .ZN(n9447) );
  XOR2_X1 U10709 ( .A(n9448), .B(n9447), .Z(n9450) );
  AOI222_X1 U10710 ( .A1(n9491), .A2(n9450), .B1(n9449), .B2(n9708), .C1(n9470), .C2(n9711), .ZN(n9577) );
  NOR2_X1 U10711 ( .A1(n9577), .A2(n9730), .ZN(n9451) );
  AOI211_X1 U10712 ( .C1(n9574), .C2(n9726), .A(n9452), .B(n9451), .ZN(n9453)
         );
  OAI21_X1 U10713 ( .B1(n9537), .B2(n9578), .A(n9453), .ZN(P1_U3269) );
  XNOR2_X1 U10714 ( .A(n4549), .B(n9460), .ZN(n9583) );
  AOI211_X1 U10715 ( .C1(n9580), .C2(n9479), .A(n9541), .B(n9454), .ZN(n9579)
         );
  AOI22_X1 U10716 ( .A1(n9730), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9455), .B2(
        n9718), .ZN(n9456) );
  OAI21_X1 U10717 ( .B1(n9457), .B2(n9521), .A(n9456), .ZN(n9465) );
  OAI21_X1 U10718 ( .B1(n9460), .B2(n9459), .A(n9458), .ZN(n9463) );
  AOI222_X1 U10719 ( .A1(n9491), .A2(n9463), .B1(n9462), .B2(n9711), .C1(n9461), .C2(n9708), .ZN(n9582) );
  NOR2_X1 U10720 ( .A1(n9582), .A2(n9730), .ZN(n9464) );
  AOI211_X1 U10721 ( .C1(n9579), .C2(n9726), .A(n9465), .B(n9464), .ZN(n9466)
         );
  OAI21_X1 U10722 ( .B1(n9537), .B2(n9583), .A(n9466), .ZN(P1_U3270) );
  OAI21_X1 U10723 ( .B1(n9468), .B2(n9474), .A(n9467), .ZN(n9469) );
  NAND2_X1 U10724 ( .A1(n9469), .A2(n9491), .ZN(n9473) );
  AOI22_X1 U10725 ( .A1(n9471), .A2(n9711), .B1(n9708), .B2(n9470), .ZN(n9472)
         );
  NAND2_X1 U10726 ( .A1(n9473), .A2(n9472), .ZN(n9588) );
  INV_X1 U10727 ( .A(n9588), .ZN(n9489) );
  AND2_X1 U10728 ( .A1(n9475), .A2(n9474), .ZN(n9477) );
  OR2_X1 U10729 ( .A1(n9477), .A2(n9476), .ZN(n9590) );
  INV_X1 U10730 ( .A(n9590), .ZN(n9487) );
  AOI21_X1 U10731 ( .B1(n9584), .B2(n9496), .A(n9541), .ZN(n9480) );
  NAND2_X1 U10732 ( .A1(n9480), .A2(n9479), .ZN(n9585) );
  AOI22_X1 U10733 ( .A1(n9730), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9718), .B2(
        n9481), .ZN(n9483) );
  NAND2_X1 U10734 ( .A1(n9584), .A2(n9719), .ZN(n9482) );
  OAI211_X1 U10735 ( .C1(n9585), .C2(n9484), .A(n9483), .B(n9482), .ZN(n9485)
         );
  AOI21_X1 U10736 ( .B1(n9487), .B2(n9486), .A(n9485), .ZN(n9488) );
  OAI21_X1 U10737 ( .B1(n9730), .B2(n9489), .A(n9488), .ZN(P1_U3271) );
  XNOR2_X1 U10738 ( .A(n9490), .B(n9492), .ZN(n9595) );
  INV_X1 U10739 ( .A(n9491), .ZN(n9713) );
  AOI21_X1 U10740 ( .B1(n9493), .B2(n9492), .A(n4560), .ZN(n9494) );
  OAI222_X1 U10741 ( .A1(n9693), .A2(n9495), .B1(n9691), .B2(n9532), .C1(n9713), .C2(n9494), .ZN(n9591) );
  INV_X1 U10742 ( .A(n9593), .ZN(n9500) );
  AOI211_X1 U10743 ( .C1(n9593), .C2(n9509), .A(n9541), .B(n9478), .ZN(n9592)
         );
  NAND2_X1 U10744 ( .A1(n9592), .A2(n9726), .ZN(n9499) );
  AOI22_X1 U10745 ( .A1(n9730), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9497), .B2(
        n9718), .ZN(n9498) );
  OAI211_X1 U10746 ( .C1(n9500), .C2(n9521), .A(n9499), .B(n9498), .ZN(n9501)
         );
  AOI21_X1 U10747 ( .B1(n9591), .B2(n9534), .A(n9501), .ZN(n9502) );
  OAI21_X1 U10748 ( .B1(n9537), .B2(n9595), .A(n9502), .ZN(P1_U3272) );
  XNOR2_X1 U10749 ( .A(n9503), .B(n9504), .ZN(n9600) );
  XOR2_X1 U10750 ( .A(n9505), .B(n9504), .Z(n9506) );
  OAI222_X1 U10751 ( .A1(n9693), .A2(n9508), .B1(n9691), .B2(n9507), .C1(n9506), .C2(n9713), .ZN(n9596) );
  INV_X1 U10752 ( .A(n9515), .ZN(n9598) );
  INV_X1 U10753 ( .A(n9519), .ZN(n9511) );
  INV_X1 U10754 ( .A(n9509), .ZN(n9510) );
  AOI211_X1 U10755 ( .C1(n9598), .C2(n9511), .A(n9541), .B(n9510), .ZN(n9597)
         );
  NAND2_X1 U10756 ( .A1(n9597), .A2(n9726), .ZN(n9514) );
  AOI22_X1 U10757 ( .A1(n9730), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9512), .B2(
        n9718), .ZN(n9513) );
  OAI211_X1 U10758 ( .C1(n9515), .C2(n9521), .A(n9514), .B(n9513), .ZN(n9516)
         );
  AOI21_X1 U10759 ( .B1(n9596), .B2(n9534), .A(n9516), .ZN(n9517) );
  OAI21_X1 U10760 ( .B1(n9600), .B2(n9537), .A(n9517), .ZN(P1_U3273) );
  XOR2_X1 U10761 ( .A(n9518), .B(n9529), .Z(n9605) );
  AOI211_X1 U10762 ( .C1(n9603), .C2(n9520), .A(n9541), .B(n9519), .ZN(n9602)
         );
  NOR2_X1 U10763 ( .A1(n4742), .A2(n9521), .ZN(n9526) );
  OAI22_X1 U10764 ( .A1(n9534), .A2(n9524), .B1(n9523), .B2(n9522), .ZN(n9525)
         );
  AOI211_X1 U10765 ( .C1(n9602), .C2(n9726), .A(n9526), .B(n9525), .ZN(n9536)
         );
  NAND2_X1 U10766 ( .A1(n9528), .A2(n9527), .ZN(n9530) );
  XNOR2_X1 U10767 ( .A(n9530), .B(n9529), .ZN(n9531) );
  OAI222_X1 U10768 ( .A1(n9691), .A2(n9533), .B1(n9693), .B2(n9532), .C1(n9713), .C2(n9531), .ZN(n9601) );
  NAND2_X1 U10769 ( .A1(n9601), .A2(n9534), .ZN(n9535) );
  OAI211_X1 U10770 ( .C1(n9605), .C2(n9537), .A(n9536), .B(n9535), .ZN(
        P1_U3274) );
  AOI21_X1 U10771 ( .B1(n9539), .B2(n9758), .A(n9538), .ZN(n9540) );
  OAI21_X1 U10772 ( .B1(n9542), .B2(n9541), .A(n9540), .ZN(n9612) );
  MUX2_X1 U10773 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9612), .S(n9863), .Z(
        P1_U3553) );
  OAI211_X1 U10774 ( .C1(n9547), .C2(n9828), .A(n9546), .B(n9545), .ZN(n9613)
         );
  MUX2_X1 U10775 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9613), .S(n9863), .Z(
        P1_U3552) );
  AOI21_X1 U10776 ( .B1(n9758), .B2(n9549), .A(n9548), .ZN(n9550) );
  OAI211_X1 U10777 ( .C1(n9552), .C2(n9762), .A(n9551), .B(n9550), .ZN(n9614)
         );
  MUX2_X1 U10778 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9614), .S(n9863), .Z(
        P1_U3551) );
  AOI21_X1 U10779 ( .B1(n9758), .B2(n9554), .A(n9553), .ZN(n9555) );
  OAI211_X1 U10780 ( .C1(n9557), .C2(n9762), .A(n9556), .B(n9555), .ZN(n9615)
         );
  MUX2_X1 U10781 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9615), .S(n9863), .Z(
        P1_U3550) );
  INV_X1 U10782 ( .A(n9558), .ZN(n9563) );
  AOI21_X1 U10783 ( .B1(n9758), .B2(n9560), .A(n9559), .ZN(n9561) );
  OAI211_X1 U10784 ( .C1(n9563), .C2(n9762), .A(n9562), .B(n9561), .ZN(n9616)
         );
  MUX2_X1 U10785 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9616), .S(n9863), .Z(
        P1_U3549) );
  AOI21_X1 U10786 ( .B1(n9758), .B2(n9565), .A(n9564), .ZN(n9566) );
  OAI211_X1 U10787 ( .C1(n9568), .C2(n9762), .A(n9567), .B(n9566), .ZN(n9617)
         );
  MUX2_X1 U10788 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9617), .S(n9863), .Z(
        P1_U3548) );
  AOI21_X1 U10789 ( .B1(n9758), .B2(n9570), .A(n9569), .ZN(n9571) );
  OAI211_X1 U10790 ( .C1(n9573), .C2(n9762), .A(n9572), .B(n9571), .ZN(n9618)
         );
  MUX2_X1 U10791 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9618), .S(n9863), .Z(
        P1_U3547) );
  AOI21_X1 U10792 ( .B1(n9758), .B2(n9575), .A(n9574), .ZN(n9576) );
  OAI211_X1 U10793 ( .C1(n9578), .C2(n9762), .A(n9577), .B(n9576), .ZN(n9619)
         );
  MUX2_X1 U10794 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9619), .S(n9863), .Z(
        P1_U3546) );
  AOI21_X1 U10795 ( .B1(n9758), .B2(n9580), .A(n9579), .ZN(n9581) );
  OAI211_X1 U10796 ( .C1(n9583), .C2(n9762), .A(n9582), .B(n9581), .ZN(n9620)
         );
  MUX2_X1 U10797 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9620), .S(n9863), .Z(
        P1_U3545) );
  INV_X1 U10798 ( .A(n9584), .ZN(n9586) );
  OAI21_X1 U10799 ( .B1(n9586), .B2(n9828), .A(n9585), .ZN(n9587) );
  NOR2_X1 U10800 ( .A1(n9588), .A2(n9587), .ZN(n9589) );
  OAI21_X1 U10801 ( .B1(n9590), .B2(n9762), .A(n9589), .ZN(n9621) );
  MUX2_X1 U10802 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9621), .S(n9863), .Z(
        P1_U3544) );
  AOI211_X1 U10803 ( .C1(n9758), .C2(n9593), .A(n9592), .B(n9591), .ZN(n9594)
         );
  OAI21_X1 U10804 ( .B1(n9762), .B2(n9595), .A(n9594), .ZN(n9622) );
  MUX2_X1 U10805 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9622), .S(n9863), .Z(
        P1_U3543) );
  AOI211_X1 U10806 ( .C1(n9758), .C2(n9598), .A(n9597), .B(n9596), .ZN(n9599)
         );
  OAI21_X1 U10807 ( .B1(n9762), .B2(n9600), .A(n9599), .ZN(n9623) );
  MUX2_X1 U10808 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9623), .S(n9863), .Z(
        P1_U3542) );
  AOI211_X1 U10809 ( .C1(n9758), .C2(n9603), .A(n9602), .B(n9601), .ZN(n9604)
         );
  OAI21_X1 U10810 ( .B1(n9605), .B2(n9762), .A(n9604), .ZN(n9624) );
  MUX2_X1 U10811 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9624), .S(n9863), .Z(
        P1_U3541) );
  AOI211_X1 U10812 ( .C1(n9758), .C2(n9608), .A(n9607), .B(n9606), .ZN(n9609)
         );
  OAI21_X1 U10813 ( .B1(n9610), .B2(n9762), .A(n9609), .ZN(n9625) );
  MUX2_X1 U10814 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9625), .S(n9863), .Z(
        P1_U3540) );
  MUX2_X1 U10815 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9611), .S(n9863), .Z(
        P1_U3522) );
  MUX2_X1 U10816 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9612), .S(n9836), .Z(
        P1_U3521) );
  MUX2_X1 U10817 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9613), .S(n9836), .Z(
        P1_U3520) );
  MUX2_X1 U10818 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9614), .S(n9836), .Z(
        P1_U3519) );
  MUX2_X1 U10819 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9615), .S(n9836), .Z(
        P1_U3518) );
  MUX2_X1 U10820 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9616), .S(n9836), .Z(
        P1_U3517) );
  MUX2_X1 U10821 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9617), .S(n9836), .Z(
        P1_U3516) );
  MUX2_X1 U10822 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9618), .S(n9836), .Z(
        P1_U3515) );
  MUX2_X1 U10823 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9619), .S(n9836), .Z(
        P1_U3514) );
  MUX2_X1 U10824 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9620), .S(n9836), .Z(
        P1_U3513) );
  MUX2_X1 U10825 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9621), .S(n9836), .Z(
        P1_U3512) );
  MUX2_X1 U10826 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9622), .S(n9836), .Z(
        P1_U3511) );
  MUX2_X1 U10827 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9623), .S(n9836), .Z(
        P1_U3510) );
  MUX2_X1 U10828 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9624), .S(n9836), .Z(
        P1_U3509) );
  MUX2_X1 U10829 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9625), .S(n9836), .Z(
        P1_U3507) );
  NOR4_X1 U10830 ( .A1(n9627), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9626), .ZN(n9628) );
  AOI21_X1 U10831 ( .B1(n9629), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9628), .ZN(
        n9630) );
  OAI21_X1 U10832 ( .B1(n9631), .B2(n9634), .A(n9630), .ZN(P1_U3324) );
  OAI222_X1 U10833 ( .A1(P1_U3086), .A2(n9635), .B1(n9634), .B2(n9633), .C1(
        n10410), .C2(n9632), .ZN(P1_U3326) );
  MUX2_X1 U10834 ( .A(n9636), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  OAI211_X1 U10835 ( .C1(n9639), .C2(n9828), .A(n9638), .B(n9637), .ZN(n9640)
         );
  AOI21_X1 U10836 ( .B1(n9641), .B2(n9824), .A(n9640), .ZN(n9656) );
  AOI22_X1 U10837 ( .A1(n9863), .A2(n9656), .B1(n9299), .B2(n9860), .ZN(
        P1_U3539) );
  NOR2_X1 U10838 ( .A1(n9642), .A2(n9762), .ZN(n9648) );
  OAI211_X1 U10839 ( .C1(n9645), .C2(n9828), .A(n9644), .B(n9643), .ZN(n9646)
         );
  AOI21_X1 U10840 ( .B1(n9648), .B2(n9647), .A(n9646), .ZN(n9658) );
  AOI22_X1 U10841 ( .A1(n9863), .A2(n9658), .B1(n9649), .B2(n9860), .ZN(
        P1_U3538) );
  OAI21_X1 U10842 ( .B1(n7480), .B2(n9828), .A(n9650), .ZN(n9651) );
  AOI211_X1 U10843 ( .C1(n9653), .C2(n9824), .A(n9652), .B(n9651), .ZN(n9660)
         );
  INV_X1 U10844 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9654) );
  AOI22_X1 U10845 ( .A1(n9863), .A2(n9660), .B1(n9654), .B2(n9860), .ZN(
        P1_U3537) );
  INV_X1 U10846 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9655) );
  AOI22_X1 U10847 ( .A1(n9836), .A2(n9656), .B1(n9655), .B2(n9834), .ZN(
        P1_U3504) );
  INV_X1 U10848 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9657) );
  AOI22_X1 U10849 ( .A1(n9836), .A2(n9658), .B1(n9657), .B2(n9834), .ZN(
        P1_U3501) );
  INV_X1 U10850 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9659) );
  AOI22_X1 U10851 ( .A1(n9836), .A2(n9660), .B1(n9659), .B2(n9834), .ZN(
        P1_U3498) );
  XNOR2_X1 U10852 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10853 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U10854 ( .B1(n4522), .B2(n9662), .A(n9661), .ZN(n9663) );
  XNOR2_X1 U10855 ( .A(n9663), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9667) );
  AOI22_X1 U10856 ( .A1(n9675), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9665) );
  OAI21_X1 U10857 ( .B1(n9667), .B2(n9666), .A(n9665), .ZN(P1_U3243) );
  NOR2_X1 U10858 ( .A1(n9669), .A2(n9668), .ZN(n9670) );
  NOR3_X1 U10859 ( .A1(n9672), .A2(n9671), .A3(n9670), .ZN(n9673) );
  AOI211_X1 U10860 ( .C1(n9675), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9674), .B(
        n9673), .ZN(n9685) );
  NAND2_X1 U10861 ( .A1(n9677), .A2(n9676), .ZN(n9683) );
  OAI211_X1 U10862 ( .C1(n9681), .C2(n9680), .A(n9679), .B(n9678), .ZN(n9682)
         );
  NAND4_X1 U10863 ( .A1(n9685), .A2(n9684), .A3(n9683), .A4(n9682), .ZN(
        P1_U3247) );
  XNOR2_X1 U10864 ( .A(n9686), .B(n9687), .ZN(n9832) );
  NAND2_X1 U10865 ( .A1(n9688), .A2(n9687), .ZN(n9689) );
  AOI21_X1 U10866 ( .B1(n9690), .B2(n9689), .A(n9713), .ZN(n9696) );
  OAI22_X1 U10867 ( .A1(n9694), .A2(n9693), .B1(n9692), .B2(n9691), .ZN(n9695)
         );
  AOI211_X1 U10868 ( .C1(n9832), .C2(n9716), .A(n9696), .B(n9695), .ZN(n9829)
         );
  AOI222_X1 U10869 ( .A1(n9699), .A2(n9719), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n9730), .C1(n9718), .C2(n9697), .ZN(n9703) );
  INV_X1 U10870 ( .A(n9698), .ZN(n9700) );
  OAI211_X1 U10871 ( .C1(n9700), .C2(n4728), .A(n9722), .B(n4730), .ZN(n9827)
         );
  INV_X1 U10872 ( .A(n9827), .ZN(n9701) );
  AOI22_X1 U10873 ( .A1(n9832), .A2(n9727), .B1(n9726), .B2(n9701), .ZN(n9702)
         );
  OAI211_X1 U10874 ( .C1(n9730), .C2(n9829), .A(n9703), .B(n9702), .ZN(
        P1_U3279) );
  XNOR2_X1 U10875 ( .A(n9704), .B(n9706), .ZN(n9791) );
  AOI21_X1 U10876 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9714) );
  AOI22_X1 U10877 ( .A1(n9711), .A2(n9710), .B1(n9709), .B2(n9708), .ZN(n9712)
         );
  OAI21_X1 U10878 ( .B1(n9714), .B2(n9713), .A(n9712), .ZN(n9715) );
  AOI21_X1 U10879 ( .B1(n9716), .B2(n9791), .A(n9715), .ZN(n9788) );
  AOI222_X1 U10880 ( .A1(n9720), .A2(n9719), .B1(P1_REG2_REG_8__SCAN_IN), .B2(
        n9730), .C1(n9718), .C2(n9717), .ZN(n9729) );
  INV_X1 U10881 ( .A(n9721), .ZN(n9723) );
  OAI211_X1 U10882 ( .C1(n9787), .C2(n9724), .A(n9723), .B(n9722), .ZN(n9786)
         );
  INV_X1 U10883 ( .A(n9786), .ZN(n9725) );
  AOI22_X1 U10884 ( .A1(n9791), .A2(n9727), .B1(n9726), .B2(n9725), .ZN(n9728)
         );
  OAI211_X1 U10885 ( .C1(n9730), .C2(n9788), .A(n9729), .B(n9728), .ZN(
        P1_U3285) );
  AND2_X1 U10886 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9731), .ZN(P1_U3294) );
  AND2_X1 U10887 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9731), .ZN(P1_U3295) );
  AND2_X1 U10888 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9731), .ZN(P1_U3296) );
  AND2_X1 U10889 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9731), .ZN(P1_U3297) );
  AND2_X1 U10890 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9731), .ZN(P1_U3298) );
  AND2_X1 U10891 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9731), .ZN(P1_U3299) );
  AND2_X1 U10892 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9731), .ZN(P1_U3300) );
  AND2_X1 U10893 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9731), .ZN(P1_U3301) );
  AND2_X1 U10894 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9731), .ZN(P1_U3302) );
  AND2_X1 U10895 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9731), .ZN(P1_U3303) );
  AND2_X1 U10896 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9731), .ZN(P1_U3304) );
  AND2_X1 U10897 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9731), .ZN(P1_U3305) );
  AND2_X1 U10898 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9731), .ZN(P1_U3306) );
  AND2_X1 U10899 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9731), .ZN(P1_U3307) );
  AND2_X1 U10900 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9731), .ZN(P1_U3308) );
  AND2_X1 U10901 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9731), .ZN(P1_U3309) );
  AND2_X1 U10902 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9731), .ZN(P1_U3310) );
  AND2_X1 U10903 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9731), .ZN(P1_U3311) );
  AND2_X1 U10904 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9731), .ZN(P1_U3312) );
  AND2_X1 U10905 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9731), .ZN(P1_U3313) );
  AND2_X1 U10906 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9731), .ZN(P1_U3314) );
  AND2_X1 U10907 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9731), .ZN(P1_U3315) );
  AND2_X1 U10908 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9731), .ZN(P1_U3316) );
  AND2_X1 U10909 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9731), .ZN(P1_U3317) );
  AND2_X1 U10910 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9731), .ZN(P1_U3318) );
  AND2_X1 U10911 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9731), .ZN(P1_U3319) );
  NOR2_X1 U10912 ( .A1(n9735), .A2(n9732), .ZN(P1_U3320) );
  NOR2_X1 U10913 ( .A1(n9735), .A2(n10247), .ZN(P1_U3321) );
  NOR2_X1 U10914 ( .A1(n9735), .A2(n9733), .ZN(P1_U3322) );
  NOR2_X1 U10915 ( .A1(n9735), .A2(n9734), .ZN(P1_U3323) );
  INV_X1 U10916 ( .A(n9736), .ZN(n9833) );
  OAI21_X1 U10917 ( .B1(n9738), .B2(n9828), .A(n9737), .ZN(n9741) );
  INV_X1 U10918 ( .A(n9739), .ZN(n9740) );
  AOI211_X1 U10919 ( .C1(n9833), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9837)
         );
  INV_X1 U10920 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9743) );
  AOI22_X1 U10921 ( .A1(n9836), .A2(n9837), .B1(n9743), .B2(n9834), .ZN(
        P1_U3456) );
  AOI21_X1 U10922 ( .B1(n9758), .B2(n9745), .A(n9744), .ZN(n9746) );
  OAI211_X1 U10923 ( .C1(n9762), .C2(n9748), .A(n9747), .B(n9746), .ZN(n9749)
         );
  INV_X1 U10924 ( .A(n9749), .ZN(n9839) );
  INV_X1 U10925 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9750) );
  AOI22_X1 U10926 ( .A1(n9836), .A2(n9839), .B1(n9750), .B2(n9834), .ZN(
        P1_U3459) );
  OAI211_X1 U10927 ( .C1(n6072), .C2(n9828), .A(n9752), .B(n9751), .ZN(n9753)
         );
  AOI21_X1 U10928 ( .B1(n9824), .B2(n9754), .A(n9753), .ZN(n9841) );
  INV_X1 U10929 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9755) );
  AOI22_X1 U10930 ( .A1(n9836), .A2(n9841), .B1(n9755), .B2(n9834), .ZN(
        P1_U3462) );
  AOI21_X1 U10931 ( .B1(n9758), .B2(n9757), .A(n9756), .ZN(n9759) );
  OAI211_X1 U10932 ( .C1(n9762), .C2(n9761), .A(n9760), .B(n9759), .ZN(n9763)
         );
  INV_X1 U10933 ( .A(n9763), .ZN(n9843) );
  INV_X1 U10934 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9764) );
  AOI22_X1 U10935 ( .A1(n9836), .A2(n9843), .B1(n9764), .B2(n9834), .ZN(
        P1_U3465) );
  OAI211_X1 U10936 ( .C1(n9767), .C2(n9828), .A(n9766), .B(n9765), .ZN(n9768)
         );
  AOI21_X1 U10937 ( .B1(n9824), .B2(n9769), .A(n9768), .ZN(n9845) );
  INV_X1 U10938 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9770) );
  AOI22_X1 U10939 ( .A1(n9836), .A2(n9845), .B1(n9770), .B2(n9834), .ZN(
        P1_U3468) );
  AND2_X1 U10940 ( .A1(n9771), .A2(n9824), .ZN(n9776) );
  INV_X1 U10941 ( .A(n9772), .ZN(n9774) );
  OAI21_X1 U10942 ( .B1(n9774), .B2(n9828), .A(n9773), .ZN(n9775) );
  NOR3_X1 U10943 ( .A1(n9777), .A2(n9776), .A3(n9775), .ZN(n9847) );
  INV_X1 U10944 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U10945 ( .A1(n9836), .A2(n9847), .B1(n9778), .B2(n9834), .ZN(
        P1_U3471) );
  OAI21_X1 U10946 ( .B1(n4740), .B2(n9828), .A(n9780), .ZN(n9781) );
  AOI21_X1 U10947 ( .B1(n9782), .B2(n9833), .A(n9781), .ZN(n9783) );
  AND2_X1 U10948 ( .A1(n9784), .A2(n9783), .ZN(n9849) );
  INV_X1 U10949 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9785) );
  AOI22_X1 U10950 ( .A1(n9836), .A2(n9849), .B1(n9785), .B2(n9834), .ZN(
        P1_U3474) );
  OAI21_X1 U10951 ( .B1(n9787), .B2(n9828), .A(n9786), .ZN(n9790) );
  INV_X1 U10952 ( .A(n9788), .ZN(n9789) );
  AOI211_X1 U10953 ( .C1(n9833), .C2(n9791), .A(n9790), .B(n9789), .ZN(n9851)
         );
  INV_X1 U10954 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9792) );
  AOI22_X1 U10955 ( .A1(n9836), .A2(n9851), .B1(n9792), .B2(n9834), .ZN(
        P1_U3477) );
  INV_X1 U10956 ( .A(n9793), .ZN(n9794) );
  OAI21_X1 U10957 ( .B1(n9795), .B2(n9828), .A(n9794), .ZN(n9798) );
  INV_X1 U10958 ( .A(n9796), .ZN(n9797) );
  AOI211_X1 U10959 ( .C1(n9824), .C2(n9799), .A(n9798), .B(n9797), .ZN(n9852)
         );
  INV_X1 U10960 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9800) );
  AOI22_X1 U10961 ( .A1(n9836), .A2(n9852), .B1(n9800), .B2(n9834), .ZN(
        P1_U3480) );
  OAI211_X1 U10962 ( .C1(n4741), .C2(n9828), .A(n9802), .B(n9801), .ZN(n9803)
         );
  AOI21_X1 U10963 ( .B1(n9804), .B2(n9824), .A(n9803), .ZN(n9854) );
  INV_X1 U10964 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9805) );
  AOI22_X1 U10965 ( .A1(n9836), .A2(n9854), .B1(n9805), .B2(n9834), .ZN(
        P1_U3483) );
  INV_X1 U10966 ( .A(n9806), .ZN(n9812) );
  INV_X1 U10967 ( .A(n9807), .ZN(n9808) );
  OAI21_X1 U10968 ( .B1(n9809), .B2(n9828), .A(n9808), .ZN(n9811) );
  AOI211_X1 U10969 ( .C1(n9833), .C2(n9812), .A(n9811), .B(n9810), .ZN(n9856)
         );
  INV_X1 U10970 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9813) );
  AOI22_X1 U10971 ( .A1(n9836), .A2(n9856), .B1(n9813), .B2(n9834), .ZN(
        P1_U3486) );
  OAI211_X1 U10972 ( .C1(n9816), .C2(n9828), .A(n9815), .B(n9814), .ZN(n9817)
         );
  AOI21_X1 U10973 ( .B1(n9824), .B2(n9818), .A(n9817), .ZN(n9858) );
  INV_X1 U10974 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9819) );
  AOI22_X1 U10975 ( .A1(n9836), .A2(n9858), .B1(n9819), .B2(n9834), .ZN(
        P1_U3489) );
  OAI21_X1 U10976 ( .B1(n9821), .B2(n9828), .A(n9820), .ZN(n9822) );
  AOI211_X1 U10977 ( .C1(n9825), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9859)
         );
  INV_X1 U10978 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9826) );
  AOI22_X1 U10979 ( .A1(n9836), .A2(n9859), .B1(n9826), .B2(n9834), .ZN(
        P1_U3492) );
  OAI21_X1 U10980 ( .B1(n4728), .B2(n9828), .A(n9827), .ZN(n9831) );
  INV_X1 U10981 ( .A(n9829), .ZN(n9830) );
  AOI211_X1 U10982 ( .C1(n9833), .C2(n9832), .A(n9831), .B(n9830), .ZN(n9862)
         );
  INV_X1 U10983 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9835) );
  AOI22_X1 U10984 ( .A1(n9836), .A2(n9862), .B1(n9835), .B2(n9834), .ZN(
        P1_U3495) );
  AOI22_X1 U10985 ( .A1(n9863), .A2(n9837), .B1(n6780), .B2(n9860), .ZN(
        P1_U3523) );
  AOI22_X1 U10986 ( .A1(n9863), .A2(n9839), .B1(n9838), .B2(n9860), .ZN(
        P1_U3524) );
  AOI22_X1 U10987 ( .A1(n9863), .A2(n9841), .B1(n9840), .B2(n9860), .ZN(
        P1_U3525) );
  AOI22_X1 U10988 ( .A1(n9863), .A2(n9843), .B1(n9842), .B2(n9860), .ZN(
        P1_U3526) );
  AOI22_X1 U10989 ( .A1(n9863), .A2(n9845), .B1(n9844), .B2(n9860), .ZN(
        P1_U3527) );
  AOI22_X1 U10990 ( .A1(n9863), .A2(n9847), .B1(n9846), .B2(n9860), .ZN(
        P1_U3528) );
  AOI22_X1 U10991 ( .A1(n9863), .A2(n9849), .B1(n9848), .B2(n9860), .ZN(
        P1_U3529) );
  AOI22_X1 U10992 ( .A1(n9863), .A2(n9851), .B1(n9850), .B2(n9860), .ZN(
        P1_U3530) );
  AOI22_X1 U10993 ( .A1(n9863), .A2(n9852), .B1(n6775), .B2(n9860), .ZN(
        P1_U3531) );
  AOI22_X1 U10994 ( .A1(n9863), .A2(n9854), .B1(n9853), .B2(n9860), .ZN(
        P1_U3532) );
  AOI22_X1 U10995 ( .A1(n9863), .A2(n9856), .B1(n9855), .B2(n9860), .ZN(
        P1_U3533) );
  AOI22_X1 U10996 ( .A1(n9863), .A2(n9858), .B1(n9857), .B2(n9860), .ZN(
        P1_U3534) );
  AOI22_X1 U10997 ( .A1(n9863), .A2(n9859), .B1(n7225), .B2(n9860), .ZN(
        P1_U3535) );
  AOI22_X1 U10998 ( .A1(n9863), .A2(n9862), .B1(n9861), .B2(n9860), .ZN(
        P1_U3536) );
  INV_X1 U10999 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U11000 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(n9915), .B1(n9933), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n9870) );
  NOR2_X1 U11001 ( .A1(n5324), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9864) );
  AOI211_X1 U11002 ( .C1(n5315), .C2(n9865), .A(P2_IR_REG_0__SCAN_IN), .B(
        n9864), .ZN(n9867) );
  OAI22_X1 U11003 ( .A1(n9868), .A2(n9964), .B1(n9867), .B2(n9866), .ZN(n9869)
         );
  OAI211_X1 U11004 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10457), .A(n9870), .B(
        n9869), .ZN(P2_U3182) );
  OAI22_X1 U11005 ( .A1(n9957), .A2(n4513), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10468), .ZN(n9881) );
  AOI21_X1 U11006 ( .B1(n9874), .B2(n9873), .A(n9872), .ZN(n9879) );
  AOI21_X1 U11007 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9878) );
  OAI22_X1 U11008 ( .A1(n9879), .A2(n9953), .B1(n9948), .B2(n9878), .ZN(n9880)
         );
  AOI211_X1 U11009 ( .C1(n9933), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n9881), .B(
        n9880), .ZN(n9886) );
  XOR2_X1 U11010 ( .A(n9883), .B(n9882), .Z(n9884) );
  NAND2_X1 U11011 ( .A1(n9884), .A2(n9964), .ZN(n9885) );
  NAND2_X1 U11012 ( .A1(n9886), .A2(n9885), .ZN(P2_U3184) );
  INV_X1 U11013 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9902) );
  AOI21_X1 U11014 ( .B1(n9889), .B2(n9888), .A(n9887), .ZN(n9893) );
  AOI21_X1 U11015 ( .B1(n9891), .B2(n9890), .A(n4609), .ZN(n9892) );
  OAI22_X1 U11016 ( .A1(n9893), .A2(n9953), .B1(n9892), .B2(n9948), .ZN(n9894)
         );
  AOI211_X1 U11017 ( .C1(n9896), .C2(n9915), .A(n9895), .B(n9894), .ZN(n9901)
         );
  XOR2_X1 U11018 ( .A(n9898), .B(n9897), .Z(n9899) );
  NAND2_X1 U11019 ( .A1(n9899), .A2(n9964), .ZN(n9900) );
  OAI211_X1 U11020 ( .C1(n9902), .C2(n9969), .A(n9901), .B(n9900), .ZN(
        P2_U3187) );
  INV_X1 U11021 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U11022 ( .A1(n9904), .A2(n9903), .ZN(n9905) );
  AND2_X1 U11023 ( .A1(n9906), .A2(n9905), .ZN(n9918) );
  NAND2_X1 U11024 ( .A1(n9908), .A2(n9907), .ZN(n9909) );
  AND2_X1 U11025 ( .A1(n9910), .A2(n9909), .ZN(n9911) );
  OR2_X1 U11026 ( .A1(n9948), .A2(n9911), .ZN(n9917) );
  INV_X1 U11027 ( .A(n9912), .ZN(n9914) );
  AOI21_X1 U11028 ( .B1(n9915), .B2(n9914), .A(n9913), .ZN(n9916) );
  OAI211_X1 U11029 ( .C1(n9953), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9919)
         );
  INV_X1 U11030 ( .A(n9919), .ZN(n9925) );
  OAI21_X1 U11031 ( .B1(n9922), .B2(n9921), .A(n9920), .ZN(n9923) );
  NAND2_X1 U11032 ( .A1(n9923), .A2(n9964), .ZN(n9924) );
  OAI211_X1 U11033 ( .C1(n9926), .C2(n9969), .A(n9925), .B(n9924), .ZN(
        P2_U3188) );
  AOI21_X1 U11034 ( .B1(n9929), .B2(n9928), .A(n9927), .ZN(n9931) );
  OAI22_X1 U11035 ( .A1(n9931), .A2(n9948), .B1(n9957), .B2(n9930), .ZN(n9932)
         );
  AOI21_X1 U11036 ( .B1(n9933), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n9932), .ZN(
        n9945) );
  INV_X1 U11037 ( .A(n9934), .ZN(n9944) );
  OAI21_X1 U11038 ( .B1(n9937), .B2(n9936), .A(n9935), .ZN(n9938) );
  NAND2_X1 U11039 ( .A1(n9938), .A2(n9964), .ZN(n9943) );
  AOI21_X1 U11040 ( .B1(n9940), .B2(n10057), .A(n9939), .ZN(n9941) );
  OR2_X1 U11041 ( .A1(n9953), .A2(n9941), .ZN(n9942) );
  NAND4_X1 U11042 ( .A1(n9945), .A2(n9944), .A3(n9943), .A4(n9942), .ZN(
        P2_U3189) );
  INV_X1 U11043 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10083) );
  NAND2_X1 U11044 ( .A1(n9947), .A2(n9946), .ZN(n9949) );
  AOI21_X1 U11045 ( .B1(n9950), .B2(n9949), .A(n9948), .ZN(n9961) );
  NAND2_X1 U11046 ( .A1(n9952), .A2(n9951), .ZN(n9954) );
  AOI21_X1 U11047 ( .B1(n9955), .B2(n9954), .A(n9953), .ZN(n9960) );
  NOR2_X1 U11048 ( .A1(n9957), .A2(n9956), .ZN(n9958) );
  NOR4_X1 U11049 ( .A1(n9961), .A2(n9960), .A3(n9959), .A4(n9958), .ZN(n9968)
         );
  NOR2_X1 U11050 ( .A1(n9963), .A2(n9962), .ZN(n9965) );
  OAI21_X1 U11051 ( .B1(n9966), .B2(n9965), .A(n9964), .ZN(n9967) );
  OAI211_X1 U11052 ( .C1(n10083), .C2(n9969), .A(n9968), .B(n9967), .ZN(
        P2_U3190) );
  XOR2_X1 U11053 ( .A(n9970), .B(n9974), .Z(n9972) );
  AOI222_X1 U11054 ( .A1(n9981), .A2(n9972), .B1(n9971), .B2(n9983), .C1(n5398), .C2(n9986), .ZN(n10010) );
  XNOR2_X1 U11055 ( .A(n9973), .B(n9974), .ZN(n10013) );
  OAI22_X1 U11056 ( .A1(n9975), .A2(n10011), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9990), .ZN(n9976) );
  AOI21_X1 U11057 ( .B1(n10013), .B2(n9977), .A(n9976), .ZN(n9978) );
  OAI221_X1 U11058 ( .B1(n5088), .B2(n10010), .C1(n9999), .C2(n5403), .A(n9978), .ZN(P2_U3230) );
  XNOR2_X1 U11059 ( .A(n4612), .B(n9979), .ZN(n9982) );
  NAND2_X1 U11060 ( .A1(n9982), .A2(n9981), .ZN(n9988) );
  AOI22_X1 U11061 ( .A1(n9986), .A2(n9985), .B1(n9984), .B2(n9983), .ZN(n9987)
         );
  NAND2_X1 U11062 ( .A1(n9988), .A2(n9987), .ZN(n10007) );
  INV_X1 U11063 ( .A(n10007), .ZN(n9998) );
  NOR2_X1 U11064 ( .A1(n9989), .A2(n10042), .ZN(n10008) );
  NOR2_X1 U11065 ( .A1(n9990), .A2(n10468), .ZN(n9991) );
  AOI21_X1 U11066 ( .B1(n10008), .B2(n9992), .A(n9991), .ZN(n9997) );
  XNOR2_X1 U11067 ( .A(n9993), .B(n9994), .ZN(n10009) );
  NAND2_X1 U11068 ( .A1(n10009), .A2(n9995), .ZN(n9996) );
  AND3_X1 U11069 ( .A1(n9998), .A2(n9997), .A3(n9996), .ZN(n10000) );
  AOI22_X1 U11070 ( .A1(n5088), .A2(n10001), .B1(n10000), .B2(n9999), .ZN(
        P2_U3231) );
  INV_X1 U11071 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10006) );
  NOR2_X1 U11072 ( .A1(n10002), .A2(n10042), .ZN(n10004) );
  AOI211_X1 U11073 ( .C1(n6582), .C2(n10005), .A(n10004), .B(n10003), .ZN(
        n10051) );
  AOI22_X1 U11074 ( .A1(n10049), .A2(n10006), .B1(n10051), .B2(n10048), .ZN(
        P2_U3393) );
  AOI211_X1 U11075 ( .C1(n10009), .C2(n10035), .A(n10008), .B(n10007), .ZN(
        n10053) );
  AOI22_X1 U11076 ( .A1(n10049), .A2(n5385), .B1(n10053), .B2(n10048), .ZN(
        P2_U3396) );
  INV_X1 U11077 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10014) );
  OAI21_X1 U11078 ( .B1(n10011), .B2(n10042), .A(n10010), .ZN(n10012) );
  AOI21_X1 U11079 ( .B1(n10035), .B2(n10013), .A(n10012), .ZN(n10054) );
  AOI22_X1 U11080 ( .A1(n10049), .A2(n10014), .B1(n10054), .B2(n10048), .ZN(
        P2_U3399) );
  INV_X1 U11081 ( .A(n10035), .ZN(n10022) );
  OR2_X1 U11082 ( .A1(n10015), .A2(n10022), .ZN(n10018) );
  OR2_X1 U11083 ( .A1(n10016), .A2(n10042), .ZN(n10017) );
  AOI22_X1 U11084 ( .A1(n10049), .A2(n5421), .B1(n10055), .B2(n10048), .ZN(
        P2_U3402) );
  INV_X1 U11085 ( .A(n10020), .ZN(n10025) );
  OAI22_X1 U11086 ( .A1(n10023), .A2(n10022), .B1(n10021), .B2(n10042), .ZN(
        n10024) );
  NOR2_X1 U11087 ( .A1(n10025), .A2(n10024), .ZN(n10056) );
  AOI22_X1 U11088 ( .A1(n10049), .A2(n5453), .B1(n10056), .B2(n10048), .ZN(
        P2_U3408) );
  INV_X1 U11089 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10030) );
  OAI22_X1 U11090 ( .A1(n10027), .A2(n10044), .B1(n10026), .B2(n10042), .ZN(
        n10028) );
  NOR2_X1 U11091 ( .A1(n10029), .A2(n10028), .ZN(n10058) );
  AOI22_X1 U11092 ( .A1(n10049), .A2(n10030), .B1(n10058), .B2(n10048), .ZN(
        P2_U3411) );
  NOR2_X1 U11093 ( .A1(n10031), .A2(n10042), .ZN(n10033) );
  AOI211_X1 U11094 ( .C1(n10035), .C2(n10034), .A(n10033), .B(n10032), .ZN(
        n10059) );
  AOI22_X1 U11095 ( .A1(n10049), .A2(n5500), .B1(n10059), .B2(n10048), .ZN(
        P2_U3414) );
  INV_X1 U11096 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10041) );
  NOR2_X1 U11097 ( .A1(n10036), .A2(n10044), .ZN(n10038) );
  AOI211_X1 U11098 ( .C1(n10040), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10061) );
  AOI22_X1 U11099 ( .A1(n10049), .A2(n10041), .B1(n10061), .B2(n10048), .ZN(
        P2_U3417) );
  OAI22_X1 U11100 ( .A1(n10045), .A2(n10044), .B1(n10043), .B2(n10042), .ZN(
        n10046) );
  NOR2_X1 U11101 ( .A1(n10047), .A2(n10046), .ZN(n10063) );
  AOI22_X1 U11102 ( .A1(n10049), .A2(n5542), .B1(n10063), .B2(n10048), .ZN(
        P2_U3420) );
  AOI22_X1 U11103 ( .A1(n10064), .A2(n10051), .B1(n10050), .B2(n10062), .ZN(
        P2_U3460) );
  AOI22_X1 U11104 ( .A1(n10064), .A2(n10053), .B1(n10052), .B2(n10062), .ZN(
        P2_U3461) );
  AOI22_X1 U11105 ( .A1(n10064), .A2(n10054), .B1(n5404), .B2(n10062), .ZN(
        P2_U3462) );
  AOI22_X1 U11106 ( .A1(n10064), .A2(n10055), .B1(n5424), .B2(n10062), .ZN(
        P2_U3463) );
  AOI22_X1 U11107 ( .A1(n10064), .A2(n10056), .B1(n5456), .B2(n10062), .ZN(
        P2_U3465) );
  AOI22_X1 U11108 ( .A1(n10064), .A2(n10058), .B1(n10057), .B2(n10062), .ZN(
        P2_U3466) );
  AOI22_X1 U11109 ( .A1(n10064), .A2(n10059), .B1(n5497), .B2(n10062), .ZN(
        P2_U3467) );
  AOI22_X1 U11110 ( .A1(n10064), .A2(n10061), .B1(n10060), .B2(n10062), .ZN(
        P2_U3468) );
  AOI22_X1 U11111 ( .A1(n10064), .A2(n10063), .B1(n5539), .B2(n10062), .ZN(
        P2_U3469) );
  AOI21_X1 U11112 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10070) );
  NAND2_X1 U11113 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10065) );
  NOR2_X1 U11114 ( .A1(n10066), .A2(n10065), .ZN(n10068) );
  NOR2_X1 U11115 ( .A1(n10070), .A2(n10068), .ZN(n10067) );
  XOR2_X1 U11116 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10067), .Z(ADD_1068_U5) );
  XOR2_X1 U11117 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11118 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10117) );
  NOR2_X1 U11119 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10114) );
  NOR2_X1 U11120 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10110) );
  NOR2_X1 U11121 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10106) );
  NOR2_X1 U11122 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10102) );
  NOR2_X1 U11123 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10098) );
  NOR2_X1 U11124 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10094) );
  NOR2_X1 U11125 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10090) );
  NOR2_X1 U11126 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10086) );
  NOR2_X1 U11127 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10082) );
  NOR2_X1 U11128 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10080) );
  NOR2_X1 U11129 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10078) );
  NOR2_X1 U11130 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10076) );
  NAND2_X1 U11131 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10074) );
  XOR2_X1 U11132 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10528) );
  NAND2_X1 U11133 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10072) );
  NOR2_X1 U11134 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10068), .ZN(n10069) );
  NOR2_X1 U11135 ( .A1(n10070), .A2(n10069), .ZN(n10518) );
  XOR2_X1 U11136 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10517) );
  NAND2_X1 U11137 ( .A1(n10518), .A2(n10517), .ZN(n10071) );
  NAND2_X1 U11138 ( .A1(n10072), .A2(n10071), .ZN(n10527) );
  NAND2_X1 U11139 ( .A1(n10528), .A2(n10527), .ZN(n10073) );
  NAND2_X1 U11140 ( .A1(n10074), .A2(n10073), .ZN(n10530) );
  XNOR2_X1 U11141 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10529) );
  NOR2_X1 U11142 ( .A1(n10530), .A2(n10529), .ZN(n10075) );
  NOR2_X1 U11143 ( .A1(n10076), .A2(n10075), .ZN(n10520) );
  XNOR2_X1 U11144 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10519) );
  NOR2_X1 U11145 ( .A1(n10520), .A2(n10519), .ZN(n10077) );
  NOR2_X1 U11146 ( .A1(n10078), .A2(n10077), .ZN(n10526) );
  XNOR2_X1 U11147 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P2_ADDR_REG_6__SCAN_IN), 
        .ZN(n10525) );
  NOR2_X1 U11148 ( .A1(n10526), .A2(n10525), .ZN(n10079) );
  NOR2_X1 U11149 ( .A1(n10080), .A2(n10079), .ZN(n10522) );
  XNOR2_X1 U11150 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10521) );
  NOR2_X1 U11151 ( .A1(n10522), .A2(n10521), .ZN(n10081) );
  NOR2_X1 U11152 ( .A1(n10082), .A2(n10081), .ZN(n10524) );
  INV_X1 U11153 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U11154 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10084), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n10083), .ZN(n10523) );
  NOR2_X1 U11155 ( .A1(n10524), .A2(n10523), .ZN(n10085) );
  NOR2_X1 U11156 ( .A1(n10086), .A2(n10085), .ZN(n10516) );
  INV_X1 U11157 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10088) );
  AOI22_X1 U11158 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10088), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n10087), .ZN(n10515) );
  NOR2_X1 U11159 ( .A1(n10516), .A2(n10515), .ZN(n10089) );
  NOR2_X1 U11160 ( .A1(n10090), .A2(n10089), .ZN(n10137) );
  INV_X1 U11161 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10092) );
  AOI22_X1 U11162 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n10092), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n10091), .ZN(n10136) );
  NOR2_X1 U11163 ( .A1(n10137), .A2(n10136), .ZN(n10093) );
  NOR2_X1 U11164 ( .A1(n10094), .A2(n10093), .ZN(n10135) );
  INV_X1 U11165 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10096) );
  AOI22_X1 U11166 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10096), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n10095), .ZN(n10134) );
  NOR2_X1 U11167 ( .A1(n10135), .A2(n10134), .ZN(n10097) );
  NOR2_X1 U11168 ( .A1(n10098), .A2(n10097), .ZN(n10133) );
  AOI22_X1 U11169 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n10100), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n10099), .ZN(n10132) );
  NOR2_X1 U11170 ( .A1(n10133), .A2(n10132), .ZN(n10101) );
  NOR2_X1 U11171 ( .A1(n10102), .A2(n10101), .ZN(n10131) );
  INV_X1 U11172 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10104) );
  INV_X1 U11173 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U11174 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n10104), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n10103), .ZN(n10130) );
  NOR2_X1 U11175 ( .A1(n10131), .A2(n10130), .ZN(n10105) );
  NOR2_X1 U11176 ( .A1(n10106), .A2(n10105), .ZN(n10129) );
  INV_X1 U11177 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10108) );
  INV_X1 U11178 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U11179 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n10108), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n10107), .ZN(n10128) );
  NOR2_X1 U11180 ( .A1(n10129), .A2(n10128), .ZN(n10109) );
  NOR2_X1 U11181 ( .A1(n10110), .A2(n10109), .ZN(n10127) );
  INV_X1 U11182 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10112) );
  INV_X1 U11183 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U11184 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n10112), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n10111), .ZN(n10126) );
  NOR2_X1 U11185 ( .A1(n10127), .A2(n10126), .ZN(n10113) );
  NOR2_X1 U11186 ( .A1(n10114), .A2(n10113), .ZN(n10125) );
  AOI22_X1 U11187 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9294), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n10115), .ZN(n10124) );
  NOR2_X1 U11188 ( .A1(n10125), .A2(n10124), .ZN(n10116) );
  NOR2_X1 U11189 ( .A1(n10117), .A2(n10116), .ZN(n10123) );
  AOI22_X1 U11190 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n10119), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n10120), .ZN(n10122) );
  NOR2_X1 U11191 ( .A1(n10123), .A2(n10122), .ZN(n10118) );
  AOI21_X1 U11192 ( .B1(n10120), .B2(n10119), .A(n10118), .ZN(n10138) );
  NAND2_X1 U11193 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10138), .ZN(n10139) );
  OAI21_X1 U11194 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10138), .A(n10139), 
        .ZN(n10121) );
  XNOR2_X1 U11195 ( .A(n10121), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  XNOR2_X1 U11196 ( .A(n10123), .B(n10122), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11197 ( .A(n10125), .B(n10124), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11198 ( .A(n10127), .B(n10126), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11199 ( .A(n10129), .B(n10128), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11200 ( .A(n10131), .B(n10130), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11201 ( .A(n10133), .B(n10132), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11202 ( .A(n10135), .B(n10134), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11203 ( .A(n10137), .B(n10136), .ZN(ADD_1068_U63) );
  XOR2_X1 U11204 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n10514) );
  INV_X1 U11205 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10141) );
  NOR2_X1 U11206 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10138), .ZN(n10140) );
  OAI21_X1 U11207 ( .B1(n10141), .B2(n10140), .A(n10139), .ZN(n10512) );
  OAI22_X1 U11208 ( .A1(P2_RD_REG_SCAN_IN), .A2(keyinput_g33), .B1(
        keyinput_g100), .B2(P1_IR_REG_10__SCAN_IN), .ZN(n10142) );
  AOI221_X1 U11209 ( .B1(P2_RD_REG_SCAN_IN), .B2(keyinput_g33), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_g100), .A(n10142), .ZN(n10149) );
  OAI22_X1 U11210 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(keyinput_g79), .B1(
        keyinput_g86), .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n10143) );
  AOI221_X1 U11211 ( .B1(P2_DATAO_REG_17__SCAN_IN), .B2(keyinput_g79), .C1(
        P2_DATAO_REG_10__SCAN_IN), .C2(keyinput_g86), .A(n10143), .ZN(n10148)
         );
  OAI22_X1 U11212 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(keyinput_g70), .B1(
        keyinput_g12), .B2(SI_20_), .ZN(n10144) );
  AOI221_X1 U11213 ( .B1(P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_g70), .C1(
        SI_20_), .C2(keyinput_g12), .A(n10144), .ZN(n10147) );
  OAI22_X1 U11214 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_g38), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .ZN(n10145) );
  AOI221_X1 U11215 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .C1(
        keyinput_g88), .C2(P2_DATAO_REG_8__SCAN_IN), .A(n10145), .ZN(n10146)
         );
  NAND4_X1 U11216 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10177) );
  OAI22_X1 U11217 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(keyinput_g78), .B1(
        keyinput_g54), .B2(P2_REG3_REG_0__SCAN_IN), .ZN(n10150) );
  AOI221_X1 U11218 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(keyinput_g78), .C1(
        P2_REG3_REG_0__SCAN_IN), .C2(keyinput_g54), .A(n10150), .ZN(n10157) );
  OAI22_X1 U11219 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        keyinput_g124), .B2(P1_D_REG_2__SCAN_IN), .ZN(n10151) );
  AOI221_X1 U11220 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        P1_D_REG_2__SCAN_IN), .C2(keyinput_g124), .A(n10151), .ZN(n10156) );
  OAI22_X1 U11221 ( .A1(SI_25_), .A2(keyinput_g7), .B1(P1_IR_REG_18__SCAN_IN), 
        .B2(keyinput_g108), .ZN(n10152) );
  AOI221_X1 U11222 ( .B1(SI_25_), .B2(keyinput_g7), .C1(keyinput_g108), .C2(
        P1_IR_REG_18__SCAN_IN), .A(n10152), .ZN(n10155) );
  OAI22_X1 U11223 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(keyinput_g43), .B1(
        keyinput_g21), .B2(SI_11_), .ZN(n10153) );
  AOI221_X1 U11224 ( .B1(P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .C1(
        SI_11_), .C2(keyinput_g21), .A(n10153), .ZN(n10154) );
  NAND4_X1 U11225 ( .A1(n10157), .A2(n10156), .A3(n10155), .A4(n10154), .ZN(
        n10176) );
  OAI22_X1 U11226 ( .A1(SI_21_), .A2(keyinput_g11), .B1(keyinput_g18), .B2(
        SI_14_), .ZN(n10158) );
  AOI221_X1 U11227 ( .B1(SI_21_), .B2(keyinput_g11), .C1(SI_14_), .C2(
        keyinput_g18), .A(n10158), .ZN(n10165) );
  OAI22_X1 U11228 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(keyinput_g41), .B1(
        keyinput_g46), .B2(P2_REG3_REG_12__SCAN_IN), .ZN(n10159) );
  AOI221_X1 U11229 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_g46), .A(n10159), .ZN(n10164)
         );
  OAI22_X1 U11230 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_g51), .B1(
        P1_IR_REG_12__SCAN_IN), .B2(keyinput_g102), .ZN(n10160) );
  AOI221_X1 U11231 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_g51), .C1(
        keyinput_g102), .C2(P1_IR_REG_12__SCAN_IN), .A(n10160), .ZN(n10163) );
  OAI22_X1 U11232 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        P1_D_REG_3__SCAN_IN), .B2(keyinput_g125), .ZN(n10161) );
  AOI221_X1 U11233 ( .B1(P2_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        keyinput_g125), .C2(P1_D_REG_3__SCAN_IN), .A(n10161), .ZN(n10162) );
  NAND4_X1 U11234 ( .A1(n10165), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        n10175) );
  OAI22_X1 U11235 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_g103), .B1(
        keyinput_g127), .B2(P1_D_REG_5__SCAN_IN), .ZN(n10166) );
  AOI221_X1 U11236 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_g103), .C1(
        P1_D_REG_5__SCAN_IN), .C2(keyinput_g127), .A(n10166), .ZN(n10173) );
  OAI22_X1 U11237 ( .A1(P2_B_REG_SCAN_IN), .A2(keyinput_g64), .B1(keyinput_g94), .B2(P1_IR_REG_4__SCAN_IN), .ZN(n10167) );
  AOI221_X1 U11238 ( .B1(P2_B_REG_SCAN_IN), .B2(keyinput_g64), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_g94), .A(n10167), .ZN(n10172) );
  OAI22_X1 U11239 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(
        keyinput_g74), .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n10168) );
  AOI221_X1 U11240 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        P2_DATAO_REG_22__SCAN_IN), .C2(keyinput_g74), .A(n10168), .ZN(n10171)
         );
  OAI22_X1 U11241 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(
        keyinput_g0), .B2(P2_WR_REG_SCAN_IN), .ZN(n10169) );
  AOI221_X1 U11242 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        P2_WR_REG_SCAN_IN), .C2(keyinput_g0), .A(n10169), .ZN(n10170) );
  NAND4_X1 U11243 ( .A1(n10173), .A2(n10172), .A3(n10171), .A4(n10170), .ZN(
        n10174) );
  NOR4_X1 U11244 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n10510) );
  OAI22_X1 U11245 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_g45), .B1(SI_8_), .B2(keyinput_g24), .ZN(n10178) );
  AOI221_X1 U11246 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .C1(
        keyinput_g24), .C2(SI_8_), .A(n10178), .ZN(n10185) );
  OAI22_X1 U11247 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        keyinput_g109), .B2(P1_IR_REG_19__SCAN_IN), .ZN(n10179) );
  AOI221_X1 U11248 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput_g109), .A(n10179), .ZN(n10184) );
  OAI22_X1 U11249 ( .A1(SI_28_), .A2(keyinput_g4), .B1(SI_27_), .B2(
        keyinput_g5), .ZN(n10180) );
  AOI221_X1 U11250 ( .B1(SI_28_), .B2(keyinput_g4), .C1(keyinput_g5), .C2(
        SI_27_), .A(n10180), .ZN(n10183) );
  OAI22_X1 U11251 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_g34), .B1(
        keyinput_g91), .B2(P1_IR_REG_1__SCAN_IN), .ZN(n10181) );
  AOI221_X1 U11252 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .C1(
        P1_IR_REG_1__SCAN_IN), .C2(keyinput_g91), .A(n10181), .ZN(n10182) );
  NAND4_X1 U11253 ( .A1(n10185), .A2(n10184), .A3(n10183), .A4(n10182), .ZN(
        n10313) );
  AOI22_X1 U11254 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_g65), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n10186) );
  OAI221_X1 U11255 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_g65), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n10186), .ZN(n10193)
         );
  AOI22_X1 U11256 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput_g99), .B1(SI_5_), 
        .B2(keyinput_g27), .ZN(n10187) );
  OAI221_X1 U11257 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput_g99), .C1(SI_5_), 
        .C2(keyinput_g27), .A(n10187), .ZN(n10192) );
  AOI22_X1 U11258 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput_g115), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_g80), .ZN(n10188) );
  OAI221_X1 U11259 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput_g115), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_g80), .A(n10188), .ZN(n10191)
         );
  AOI22_X1 U11260 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(keyinput_g56), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n10189) );
  OAI221_X1 U11261 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n10189), .ZN(n10190)
         );
  NOR4_X1 U11262 ( .A1(n10193), .A2(n10192), .A3(n10191), .A4(n10190), .ZN(
        n10211) );
  AOI22_X1 U11263 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(keyinput_g112), .B1(SI_2_), 
        .B2(keyinput_g30), .ZN(n10194) );
  OAI221_X1 U11264 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(keyinput_g112), .C1(SI_2_), .C2(keyinput_g30), .A(n10194), .ZN(n10201) );
  AOI22_X1 U11265 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_g104), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_g85), .ZN(n10195) );
  OAI221_X1 U11266 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_g104), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_g85), .A(n10195), .ZN(n10200)
         );
  AOI22_X1 U11267 ( .A1(P1_D_REG_1__SCAN_IN), .A2(keyinput_g123), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .ZN(n10196) );
  OAI221_X1 U11268 ( .B1(P1_D_REG_1__SCAN_IN), .B2(keyinput_g123), .C1(
        P2_REG3_REG_2__SCAN_IN), .C2(keyinput_g59), .A(n10196), .ZN(n10199) );
  AOI22_X1 U11269 ( .A1(SI_6_), .A2(keyinput_g26), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(keyinput_g68), .ZN(n10197) );
  OAI221_X1 U11270 ( .B1(SI_6_), .B2(keyinput_g26), .C1(
        P2_DATAO_REG_28__SCAN_IN), .C2(keyinput_g68), .A(n10197), .ZN(n10198)
         );
  NOR4_X1 U11271 ( .A1(n10201), .A2(n10200), .A3(n10199), .A4(n10198), .ZN(
        n10210) );
  OAI22_X1 U11272 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_g72), .B1(
        SI_7_), .B2(keyinput_g25), .ZN(n10202) );
  AOI221_X1 U11273 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_g72), .C1(
        keyinput_g25), .C2(SI_7_), .A(n10202), .ZN(n10208) );
  OAI22_X1 U11274 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(keyinput_g69), .B1(
        P1_IR_REG_30__SCAN_IN), .B2(keyinput_g120), .ZN(n10203) );
  AOI221_X1 U11275 ( .B1(P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_g69), .C1(
        keyinput_g120), .C2(P1_IR_REG_30__SCAN_IN), .A(n10203), .ZN(n10207) );
  OAI22_X1 U11276 ( .A1(SI_15_), .A2(keyinput_g17), .B1(P1_IR_REG_27__SCAN_IN), 
        .B2(keyinput_g117), .ZN(n10204) );
  AOI221_X1 U11277 ( .B1(SI_15_), .B2(keyinput_g17), .C1(keyinput_g117), .C2(
        P1_IR_REG_27__SCAN_IN), .A(n10204), .ZN(n10206) );
  XNOR2_X1 U11278 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput_g119), .ZN(n10205)
         );
  AND4_X1 U11279 ( .A1(n10208), .A2(n10207), .A3(n10206), .A4(n10205), .ZN(
        n10209) );
  NAND3_X1 U11280 ( .A1(n10211), .A2(n10210), .A3(n10209), .ZN(n10312) );
  AOI22_X1 U11281 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput_g110), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .ZN(n10212) );
  OAI221_X1 U11282 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput_g110), .C1(
        P2_DATAO_REG_14__SCAN_IN), .C2(keyinput_g82), .A(n10212), .ZN(n10221)
         );
  AOI22_X1 U11283 ( .A1(n5482), .A2(keyinput_g35), .B1(keyinput_g77), .B2(
        n10214), .ZN(n10213) );
  OAI221_X1 U11284 ( .B1(n5482), .B2(keyinput_g35), .C1(n10214), .C2(
        keyinput_g77), .A(n10213), .ZN(n10220) );
  AOI22_X1 U11285 ( .A1(SI_30_), .A2(keyinput_g2), .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .ZN(n10215) );
  OAI221_X1 U11286 ( .B1(SI_30_), .B2(keyinput_g2), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_g48), .A(n10215), .ZN(n10219)
         );
  XNOR2_X1 U11287 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_g114), .ZN(n10217)
         );
  XNOR2_X1 U11288 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_g71), .ZN(n10216) );
  NAND2_X1 U11289 ( .A1(n10217), .A2(n10216), .ZN(n10218) );
  NOR4_X1 U11290 ( .A1(n10221), .A2(n10220), .A3(n10219), .A4(n10218), .ZN(
        n10262) );
  AOI22_X1 U11291 ( .A1(n10223), .A2(keyinput_g40), .B1(keyinput_g116), .B2(
        n5941), .ZN(n10222) );
  OAI221_X1 U11292 ( .B1(n10223), .B2(keyinput_g40), .C1(n5941), .C2(
        keyinput_g116), .A(n10222), .ZN(n10234) );
  AOI22_X1 U11293 ( .A1(n5514), .A2(keyinput_g53), .B1(keyinput_g84), .B2(
        n10225), .ZN(n10224) );
  OAI221_X1 U11294 ( .B1(n5514), .B2(keyinput_g53), .C1(n10225), .C2(
        keyinput_g84), .A(n10224), .ZN(n10233) );
  AOI22_X1 U11295 ( .A1(n10228), .A2(keyinput_g23), .B1(n10227), .B2(
        keyinput_g3), .ZN(n10226) );
  OAI221_X1 U11296 ( .B1(n10228), .B2(keyinput_g23), .C1(n10227), .C2(
        keyinput_g3), .A(n10226), .ZN(n10232) );
  XOR2_X1 U11297 ( .A(n5946), .B(keyinput_g118), .Z(n10230) );
  XNOR2_X1 U11298 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10229) );
  NAND2_X1 U11299 ( .A1(n10230), .A2(n10229), .ZN(n10231) );
  NOR4_X1 U11300 ( .A1(n10234), .A2(n10233), .A3(n10232), .A4(n10231), .ZN(
        n10261) );
  AOI22_X1 U11301 ( .A1(n10456), .A2(keyinput_g62), .B1(keyinput_g113), .B2(
        n6523), .ZN(n10235) );
  OAI221_X1 U11302 ( .B1(n10456), .B2(keyinput_g62), .C1(n6523), .C2(
        keyinput_g113), .A(n10235), .ZN(n10245) );
  INV_X1 U11303 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U11304 ( .A1(n10471), .A2(keyinput_g93), .B1(n10237), .B2(
        keyinput_g87), .ZN(n10236) );
  OAI221_X1 U11305 ( .B1(n10471), .B2(keyinput_g93), .C1(n10237), .C2(
        keyinput_g87), .A(n10236), .ZN(n10244) );
  INV_X1 U11306 ( .A(SI_12_), .ZN(n10443) );
  AOI22_X1 U11307 ( .A1(n10443), .A2(keyinput_g20), .B1(keyinput_g90), .B2(
        n10239), .ZN(n10238) );
  OAI221_X1 U11308 ( .B1(n10443), .B2(keyinput_g20), .C1(n10239), .C2(
        keyinput_g90), .A(n10238), .ZN(n10243) );
  XOR2_X1 U11309 ( .A(n5967), .B(keyinput_g107), .Z(n10241) );
  XNOR2_X1 U11310 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g96), .ZN(n10240) );
  NAND2_X1 U11311 ( .A1(n10241), .A2(n10240), .ZN(n10242) );
  NOR4_X1 U11312 ( .A1(n10245), .A2(n10244), .A3(n10243), .A4(n10242), .ZN(
        n10260) );
  AOI22_X1 U11313 ( .A1(n10248), .A2(keyinput_g50), .B1(keyinput_g126), .B2(
        n10247), .ZN(n10246) );
  OAI221_X1 U11314 ( .B1(n10248), .B2(keyinput_g50), .C1(n10247), .C2(
        keyinput_g126), .A(n10246), .ZN(n10258) );
  AOI22_X1 U11315 ( .A1(n10489), .A2(keyinput_g73), .B1(keyinput_g122), .B2(
        n10424), .ZN(n10249) );
  OAI221_X1 U11316 ( .B1(n10489), .B2(keyinput_g73), .C1(n10424), .C2(
        keyinput_g122), .A(n10249), .ZN(n10257) );
  AOI22_X1 U11317 ( .A1(n10454), .A2(keyinput_g55), .B1(keyinput_g9), .B2(
        n10251), .ZN(n10250) );
  OAI221_X1 U11318 ( .B1(n10454), .B2(keyinput_g55), .C1(n10251), .C2(
        keyinput_g9), .A(n10250), .ZN(n10256) );
  AOI22_X1 U11319 ( .A1(n10254), .A2(keyinput_g14), .B1(keyinput_g66), .B2(
        n10253), .ZN(n10252) );
  OAI221_X1 U11320 ( .B1(n10254), .B2(keyinput_g14), .C1(n10253), .C2(
        keyinput_g66), .A(n10252), .ZN(n10255) );
  NOR4_X1 U11321 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10259) );
  NAND4_X1 U11322 ( .A1(n10262), .A2(n10261), .A3(n10260), .A4(n10259), .ZN(
        n10311) );
  INV_X1 U11323 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n10486) );
  AOI22_X1 U11324 ( .A1(n10470), .A2(keyinput_g39), .B1(keyinput_g95), .B2(
        n10486), .ZN(n10263) );
  OAI221_X1 U11325 ( .B1(n10470), .B2(keyinput_g39), .C1(n10486), .C2(
        keyinput_g95), .A(n10263), .ZN(n10275) );
  INV_X1 U11326 ( .A(SI_13_), .ZN(n10265) );
  AOI22_X1 U11327 ( .A1(n10266), .A2(keyinput_g28), .B1(n10265), .B2(
        keyinput_g19), .ZN(n10264) );
  OAI221_X1 U11328 ( .B1(n10266), .B2(keyinput_g28), .C1(n10265), .C2(
        keyinput_g19), .A(n10264), .ZN(n10274) );
  AOI22_X1 U11329 ( .A1(n10269), .A2(keyinput_g52), .B1(n10268), .B2(
        keyinput_g57), .ZN(n10267) );
  OAI221_X1 U11330 ( .B1(n10269), .B2(keyinput_g52), .C1(n10268), .C2(
        keyinput_g57), .A(n10267), .ZN(n10273) );
  XNOR2_X1 U11331 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_g105), .ZN(n10271)
         );
  XNOR2_X1 U11332 ( .A(SI_19_), .B(keyinput_g13), .ZN(n10270) );
  NAND2_X1 U11333 ( .A1(n10271), .A2(n10270), .ZN(n10272) );
  NOR4_X1 U11334 ( .A1(n10275), .A2(n10274), .A3(n10273), .A4(n10272), .ZN(
        n10309) );
  AOI22_X1 U11335 ( .A1(n7799), .A2(keyinput_g1), .B1(n10277), .B2(
        keyinput_g83), .ZN(n10276) );
  OAI221_X1 U11336 ( .B1(n7799), .B2(keyinput_g1), .C1(n10277), .C2(
        keyinput_g83), .A(n10276), .ZN(n10286) );
  INV_X1 U11337 ( .A(SI_3_), .ZN(n10390) );
  AOI22_X1 U11338 ( .A1(n10279), .A2(keyinput_g10), .B1(keyinput_g29), .B2(
        n10390), .ZN(n10278) );
  OAI221_X1 U11339 ( .B1(n10279), .B2(keyinput_g10), .C1(n10390), .C2(
        keyinput_g29), .A(n10278), .ZN(n10285) );
  XNOR2_X1 U11340 ( .A(SI_0_), .B(keyinput_g32), .ZN(n10283) );
  XNOR2_X1 U11341 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_g37), .ZN(n10282)
         );
  XNOR2_X1 U11342 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_g121), .ZN(n10281)
         );
  XNOR2_X1 U11343 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_g36), .ZN(n10280)
         );
  NAND4_X1 U11344 ( .A1(n10283), .A2(n10282), .A3(n10281), .A4(n10280), .ZN(
        n10284) );
  NOR3_X1 U11345 ( .A1(n10286), .A2(n10285), .A3(n10284), .ZN(n10308) );
  INV_X1 U11346 ( .A(SI_16_), .ZN(n10397) );
  AOI22_X1 U11347 ( .A1(n10397), .A2(keyinput_g16), .B1(n5779), .B2(
        keyinput_g47), .ZN(n10287) );
  OAI221_X1 U11348 ( .B1(n10397), .B2(keyinput_g16), .C1(n5779), .C2(
        keyinput_g47), .A(n10287), .ZN(n10296) );
  AOI22_X1 U11349 ( .A1(n10427), .A2(keyinput_g6), .B1(keyinput_g8), .B2(
        n10289), .ZN(n10288) );
  OAI221_X1 U11350 ( .B1(n10427), .B2(keyinput_g6), .C1(n10289), .C2(
        keyinput_g8), .A(n10288), .ZN(n10295) );
  XNOR2_X1 U11351 ( .A(SI_17_), .B(keyinput_g15), .ZN(n10293) );
  XNOR2_X1 U11352 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_g111), .ZN(n10292)
         );
  XNOR2_X1 U11353 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g97), .ZN(n10291) );
  XNOR2_X1 U11354 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_g89), .ZN(n10290)
         );
  NAND4_X1 U11355 ( .A1(n10293), .A2(n10292), .A3(n10291), .A4(n10290), .ZN(
        n10294) );
  NOR3_X1 U11356 ( .A1(n10296), .A2(n10295), .A3(n10294), .ZN(n10307) );
  INV_X1 U11357 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U11358 ( .A1(n10458), .A2(keyinput_g98), .B1(n10410), .B2(
        keyinput_g67), .ZN(n10297) );
  OAI221_X1 U11359 ( .B1(n10458), .B2(keyinput_g98), .C1(n10410), .C2(
        keyinput_g67), .A(n10297), .ZN(n10305) );
  XOR2_X1 U11360 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_g44), .Z(n10304) );
  XNOR2_X1 U11361 ( .A(keyinput_g92), .B(n6067), .ZN(n10303) );
  XNOR2_X1 U11362 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_g101), .ZN(n10301)
         );
  XNOR2_X1 U11363 ( .A(SI_10_), .B(keyinput_g22), .ZN(n10300) );
  XNOR2_X1 U11364 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_g106), .ZN(n10299)
         );
  XNOR2_X1 U11365 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_g76), .ZN(n10298) );
  NAND4_X1 U11366 ( .A1(n10301), .A2(n10300), .A3(n10299), .A4(n10298), .ZN(
        n10302) );
  NOR4_X1 U11367 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n10306) );
  NAND4_X1 U11368 ( .A1(n10309), .A2(n10308), .A3(n10307), .A4(n10306), .ZN(
        n10310) );
  NOR4_X1 U11369 ( .A1(n10313), .A2(n10312), .A3(n10311), .A4(n10310), .ZN(
        n10509) );
  XOR2_X1 U11370 ( .A(SI_6_), .B(keyinput_f26), .Z(n10320) );
  AOI22_X1 U11371 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(keyinput_f117), .B1(
        P1_IR_REG_4__SCAN_IN), .B2(keyinput_f94), .ZN(n10314) );
  OAI221_X1 U11372 ( .B1(P1_IR_REG_27__SCAN_IN), .B2(keyinput_f117), .C1(
        P1_IR_REG_4__SCAN_IN), .C2(keyinput_f94), .A(n10314), .ZN(n10319) );
  AOI22_X1 U11373 ( .A1(keyinput_f0), .A2(P2_WR_REG_SCAN_IN), .B1(SI_31_), 
        .B2(keyinput_f1), .ZN(n10315) );
  OAI221_X1 U11374 ( .B1(keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .C1(SI_31_), 
        .C2(keyinput_f1), .A(n10315), .ZN(n10318) );
  AOI22_X1 U11375 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_f108), .B1(SI_13_), .B2(keyinput_f19), .ZN(n10316) );
  OAI221_X1 U11376 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_f108), .C1(
        SI_13_), .C2(keyinput_f19), .A(n10316), .ZN(n10317) );
  NOR4_X1 U11377 ( .A1(n10320), .A2(n10319), .A3(n10318), .A4(n10317), .ZN(
        n10348) );
  AOI22_X1 U11378 ( .A1(P1_D_REG_4__SCAN_IN), .A2(keyinput_f126), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput_f110), .ZN(n10321) );
  OAI221_X1 U11379 ( .B1(P1_D_REG_4__SCAN_IN), .B2(keyinput_f126), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput_f110), .A(n10321), .ZN(n10328) );
  AOI22_X1 U11380 ( .A1(SI_22_), .A2(keyinput_f10), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n10322) );
  OAI221_X1 U11381 ( .B1(SI_22_), .B2(keyinput_f10), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n10322), .ZN(n10327)
         );
  AOI22_X1 U11382 ( .A1(P1_D_REG_2__SCAN_IN), .A2(keyinput_f124), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(keyinput_f70), .ZN(n10323) );
  OAI221_X1 U11383 ( .B1(P1_D_REG_2__SCAN_IN), .B2(keyinput_f124), .C1(
        P2_DATAO_REG_26__SCAN_IN), .C2(keyinput_f70), .A(n10323), .ZN(n10326)
         );
  AOI22_X1 U11384 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(keyinput_f89), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .ZN(n10324) );
  OAI221_X1 U11385 ( .B1(P2_DATAO_REG_7__SCAN_IN), .B2(keyinput_f89), .C1(
        P2_REG3_REG_7__SCAN_IN), .C2(keyinput_f35), .A(n10324), .ZN(n10325) );
  NOR4_X1 U11386 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10347) );
  AOI22_X1 U11387 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_f113), .B1(
        P2_REG3_REG_4__SCAN_IN), .B2(keyinput_f52), .ZN(n10329) );
  OAI221_X1 U11388 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput_f113), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n10329), .ZN(n10336) );
  AOI22_X1 U11389 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n10330) );
  OAI221_X1 U11390 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n10330), .ZN(n10335)
         );
  AOI22_X1 U11391 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(keyinput_f48), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .ZN(n10331) );
  OAI221_X1 U11392 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_f36), .A(n10331), .ZN(n10334)
         );
  AOI22_X1 U11393 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(keyinput_f90), .B1(SI_29_), 
        .B2(keyinput_f3), .ZN(n10332) );
  OAI221_X1 U11394 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(keyinput_f90), .C1(SI_29_), 
        .C2(keyinput_f3), .A(n10332), .ZN(n10333) );
  NOR4_X1 U11395 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n10346) );
  AOI22_X1 U11396 ( .A1(SI_30_), .A2(keyinput_f2), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput_f80), .ZN(n10337) );
  OAI221_X1 U11397 ( .B1(SI_30_), .B2(keyinput_f2), .C1(
        P2_DATAO_REG_16__SCAN_IN), .C2(keyinput_f80), .A(n10337), .ZN(n10344)
         );
  AOI22_X1 U11398 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput_f116), .B1(SI_21_), .B2(keyinput_f11), .ZN(n10338) );
  OAI221_X1 U11399 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput_f116), .C1(
        SI_21_), .C2(keyinput_f11), .A(n10338), .ZN(n10343) );
  AOI22_X1 U11400 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput_f118), .B1(SI_23_), .B2(keyinput_f9), .ZN(n10339) );
  OAI221_X1 U11401 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput_f118), .C1(
        SI_23_), .C2(keyinput_f9), .A(n10339), .ZN(n10342) );
  AOI22_X1 U11402 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(keyinput_f100), .B1(SI_24_), .B2(keyinput_f8), .ZN(n10340) );
  OAI221_X1 U11403 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(keyinput_f100), .C1(
        SI_24_), .C2(keyinput_f8), .A(n10340), .ZN(n10341) );
  NOR4_X1 U11404 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10345) );
  NAND4_X1 U11405 ( .A1(n10348), .A2(n10347), .A3(n10346), .A4(n10345), .ZN(
        n10503) );
  AOI22_X1 U11406 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput_f125), .B1(
        P2_REG3_REG_8__SCAN_IN), .B2(keyinput_f43), .ZN(n10349) );
  OAI221_X1 U11407 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput_f125), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_f43), .A(n10349), .ZN(n10356) );
  AOI22_X1 U11408 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(keyinput_f88), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(keyinput_f85), .ZN(n10350) );
  OAI221_X1 U11409 ( .B1(P2_DATAO_REG_8__SCAN_IN), .B2(keyinput_f88), .C1(
        P2_DATAO_REG_11__SCAN_IN), .C2(keyinput_f85), .A(n10350), .ZN(n10355)
         );
  AOI22_X1 U11410 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_f107), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n10351) );
  OAI221_X1 U11411 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_f107), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n10351), .ZN(n10354)
         );
  AOI22_X1 U11412 ( .A1(P1_D_REG_5__SCAN_IN), .A2(keyinput_f127), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .ZN(n10352) );
  OAI221_X1 U11413 ( .B1(P1_D_REG_5__SCAN_IN), .B2(keyinput_f127), .C1(
        P2_REG3_REG_1__SCAN_IN), .C2(keyinput_f44), .A(n10352), .ZN(n10353) );
  NOR4_X1 U11414 ( .A1(n10356), .A2(n10355), .A3(n10354), .A4(n10353), .ZN(
        n10384) );
  AOI22_X1 U11415 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n10357) );
  OAI221_X1 U11416 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n10357), .ZN(n10364)
         );
  AOI22_X1 U11417 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(keyinput_f66), .B1(
        P1_IR_REG_22__SCAN_IN), .B2(keyinput_f112), .ZN(n10358) );
  OAI221_X1 U11418 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .C1(
        P1_IR_REG_22__SCAN_IN), .C2(keyinput_f112), .A(n10358), .ZN(n10363) );
  AOI22_X1 U11419 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_f103), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(keyinput_f84), .ZN(n10359) );
  OAI221_X1 U11420 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_f103), .C1(
        P2_DATAO_REG_12__SCAN_IN), .C2(keyinput_f84), .A(n10359), .ZN(n10362)
         );
  AOI22_X1 U11421 ( .A1(SI_4_), .A2(keyinput_f28), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(keyinput_f83), .ZN(n10360) );
  OAI221_X1 U11422 ( .B1(SI_4_), .B2(keyinput_f28), .C1(
        P2_DATAO_REG_13__SCAN_IN), .C2(keyinput_f83), .A(n10360), .ZN(n10361)
         );
  NOR4_X1 U11423 ( .A1(n10364), .A2(n10363), .A3(n10362), .A4(n10361), .ZN(
        n10383) );
  AOI22_X1 U11424 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput_f119), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .ZN(n10365) );
  OAI221_X1 U11425 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput_f119), .C1(
        P2_REG3_REG_17__SCAN_IN), .C2(keyinput_f50), .A(n10365), .ZN(n10372)
         );
  AOI22_X1 U11426 ( .A1(SI_18_), .A2(keyinput_f14), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n10366) );
  OAI221_X1 U11427 ( .B1(SI_18_), .B2(keyinput_f14), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n10366), .ZN(n10371)
         );
  AOI22_X1 U11428 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(keyinput_f120), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(keyinput_f77), .ZN(n10367) );
  OAI221_X1 U11429 ( .B1(P1_IR_REG_30__SCAN_IN), .B2(keyinput_f120), .C1(
        P2_DATAO_REG_19__SCAN_IN), .C2(keyinput_f77), .A(n10367), .ZN(n10370)
         );
  AOI22_X1 U11430 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(keyinput_f102), .B1(SI_27_), .B2(keyinput_f5), .ZN(n10368) );
  OAI221_X1 U11431 ( .B1(P1_IR_REG_12__SCAN_IN), .B2(keyinput_f102), .C1(
        SI_27_), .C2(keyinput_f5), .A(n10368), .ZN(n10369) );
  NOR4_X1 U11432 ( .A1(n10372), .A2(n10371), .A3(n10370), .A4(n10369), .ZN(
        n10382) );
  AOI22_X1 U11433 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(keyinput_f72), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(keyinput_f69), .ZN(n10373) );
  OAI221_X1 U11434 ( .B1(P2_DATAO_REG_24__SCAN_IN), .B2(keyinput_f72), .C1(
        P2_DATAO_REG_27__SCAN_IN), .C2(keyinput_f69), .A(n10373), .ZN(n10380)
         );
  AOI22_X1 U11435 ( .A1(SI_1_), .A2(keyinput_f31), .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .ZN(n10374) );
  OAI221_X1 U11436 ( .B1(SI_1_), .B2(keyinput_f31), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_f56), .A(n10374), .ZN(n10379)
         );
  AOI22_X1 U11437 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(keyinput_f114), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(keyinput_f71), .ZN(n10375) );
  OAI221_X1 U11438 ( .B1(P1_IR_REG_24__SCAN_IN), .B2(keyinput_f114), .C1(
        P2_DATAO_REG_25__SCAN_IN), .C2(keyinput_f71), .A(n10375), .ZN(n10378)
         );
  AOI22_X1 U11439 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(keyinput_f115), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .ZN(n10376) );
  OAI221_X1 U11440 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(keyinput_f115), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n10376), .ZN(n10377) );
  NOR4_X1 U11441 ( .A1(n10380), .A2(n10379), .A3(n10378), .A4(n10377), .ZN(
        n10381) );
  NAND4_X1 U11442 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10502) );
  AOI22_X1 U11443 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput_f91), .B1(SI_7_), 
        .B2(keyinput_f25), .ZN(n10385) );
  OAI221_X1 U11444 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput_f91), .C1(SI_7_), 
        .C2(keyinput_f25), .A(n10385), .ZN(n10394) );
  AOI22_X1 U11445 ( .A1(SI_11_), .A2(keyinput_f21), .B1(SI_17_), .B2(
        keyinput_f15), .ZN(n10386) );
  OAI221_X1 U11446 ( .B1(SI_11_), .B2(keyinput_f21), .C1(SI_17_), .C2(
        keyinput_f15), .A(n10386), .ZN(n10393) );
  AOI22_X1 U11447 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_f65), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n10387) );
  OAI221_X1 U11448 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_f65), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n10387), .ZN(n10392)
         );
  AOI22_X1 U11449 ( .A1(n10390), .A2(keyinput_f29), .B1(n10389), .B2(
        keyinput_f58), .ZN(n10388) );
  OAI221_X1 U11450 ( .B1(n10390), .B2(keyinput_f29), .C1(n10389), .C2(
        keyinput_f58), .A(n10388), .ZN(n10391) );
  NOR4_X1 U11451 ( .A1(n10394), .A2(n10393), .A3(n10392), .A4(n10391), .ZN(
        n10440) );
  INV_X1 U11452 ( .A(SI_14_), .ZN(n10396) );
  AOI22_X1 U11453 ( .A1(n10397), .A2(keyinput_f16), .B1(keyinput_f18), .B2(
        n10396), .ZN(n10395) );
  OAI221_X1 U11454 ( .B1(n10397), .B2(keyinput_f16), .C1(n10396), .C2(
        keyinput_f18), .A(n10395), .ZN(n10407) );
  AOI22_X1 U11455 ( .A1(n6210), .A2(keyinput_f99), .B1(keyinput_f123), .B2(
        n10399), .ZN(n10398) );
  OAI221_X1 U11456 ( .B1(n6210), .B2(keyinput_f99), .C1(n10399), .C2(
        keyinput_f123), .A(n10398), .ZN(n10406) );
  AOI22_X1 U11457 ( .A1(n10401), .A2(keyinput_f78), .B1(keyinput_f109), .B2(
        n5953), .ZN(n10400) );
  OAI221_X1 U11458 ( .B1(n10401), .B2(keyinput_f78), .C1(n5953), .C2(
        keyinput_f109), .A(n10400), .ZN(n10405) );
  AOI22_X1 U11459 ( .A1(n5367), .A2(keyinput_f33), .B1(keyinput_f79), .B2(
        n10403), .ZN(n10402) );
  OAI221_X1 U11460 ( .B1(n5367), .B2(keyinput_f33), .C1(n10403), .C2(
        keyinput_f79), .A(n10402), .ZN(n10404) );
  NOR4_X1 U11461 ( .A1(n10407), .A2(n10406), .A3(n10405), .A4(n10404), .ZN(
        n10439) );
  AOI22_X1 U11462 ( .A1(n10410), .A2(keyinput_f67), .B1(keyinput_f7), .B2(
        n10409), .ZN(n10408) );
  OAI221_X1 U11463 ( .B1(n10410), .B2(keyinput_f67), .C1(n10409), .C2(
        keyinput_f7), .A(n10408), .ZN(n10422) );
  INV_X1 U11464 ( .A(SI_10_), .ZN(n10412) );
  AOI22_X1 U11465 ( .A1(n10413), .A2(keyinput_f75), .B1(keyinput_f22), .B2(
        n10412), .ZN(n10411) );
  OAI221_X1 U11466 ( .B1(n10413), .B2(keyinput_f75), .C1(n10412), .C2(
        keyinput_f22), .A(n10411), .ZN(n10421) );
  AOI22_X1 U11467 ( .A1(n10416), .A2(keyinput_f24), .B1(n10415), .B2(
        keyinput_f74), .ZN(n10414) );
  OAI221_X1 U11468 ( .B1(n10416), .B2(keyinput_f24), .C1(n10415), .C2(
        keyinput_f74), .A(n10414), .ZN(n10420) );
  XNOR2_X1 U11469 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput_f111), .ZN(n10418)
         );
  XNOR2_X1 U11470 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_f97), .ZN(n10417) );
  NAND2_X1 U11471 ( .A1(n10418), .A2(n10417), .ZN(n10419) );
  NOR4_X1 U11472 ( .A1(n10422), .A2(n10421), .A3(n10420), .A4(n10419), .ZN(
        n10438) );
  AOI22_X1 U11473 ( .A1(n10425), .A2(keyinput_f68), .B1(keyinput_f122), .B2(
        n10424), .ZN(n10423) );
  OAI221_X1 U11474 ( .B1(n10425), .B2(keyinput_f68), .C1(n10424), .C2(
        keyinput_f122), .A(n10423), .ZN(n10436) );
  AOI22_X1 U11475 ( .A1(n5437), .A2(keyinput_f49), .B1(keyinput_f6), .B2(
        n10427), .ZN(n10426) );
  OAI221_X1 U11476 ( .B1(n5437), .B2(keyinput_f49), .C1(n10427), .C2(
        keyinput_f6), .A(n10426), .ZN(n10435) );
  AOI22_X1 U11477 ( .A1(n10430), .A2(keyinput_f82), .B1(n10429), .B2(
        keyinput_f17), .ZN(n10428) );
  OAI221_X1 U11478 ( .B1(n10430), .B2(keyinput_f82), .C1(n10429), .C2(
        keyinput_f17), .A(n10428), .ZN(n10434) );
  XNOR2_X1 U11479 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_f105), .ZN(n10432)
         );
  XNOR2_X1 U11480 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_f87), .ZN(n10431)
         );
  NAND2_X1 U11481 ( .A1(n10432), .A2(n10431), .ZN(n10433) );
  NOR4_X1 U11482 ( .A1(n10436), .A2(n10435), .A3(n10434), .A4(n10433), .ZN(
        n10437) );
  NAND4_X1 U11483 ( .A1(n10440), .A2(n10439), .A3(n10438), .A4(n10437), .ZN(
        n10501) );
  AOI22_X1 U11484 ( .A1(n10443), .A2(keyinput_f20), .B1(n10442), .B2(
        keyinput_f12), .ZN(n10441) );
  OAI221_X1 U11485 ( .B1(n10443), .B2(keyinput_f20), .C1(n10442), .C2(
        keyinput_f12), .A(n10441), .ZN(n10452) );
  XOR2_X1 U11486 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput_f101), .Z(n10451) );
  INV_X1 U11487 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10444) );
  XNOR2_X1 U11488 ( .A(keyinput_f38), .B(n10444), .ZN(n10450) );
  XNOR2_X1 U11489 ( .A(SI_9_), .B(keyinput_f23), .ZN(n10448) );
  XNOR2_X1 U11490 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_f106), .ZN(n10447)
         );
  XNOR2_X1 U11491 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(keyinput_f76), .ZN(n10446) );
  XNOR2_X1 U11492 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_f104), .ZN(n10445)
         );
  NAND4_X1 U11493 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        n10449) );
  NOR4_X1 U11494 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10499) );
  AOI22_X1 U11495 ( .A1(n10454), .A2(keyinput_f55), .B1(keyinput_f53), .B2(
        n5514), .ZN(n10453) );
  OAI221_X1 U11496 ( .B1(n10454), .B2(keyinput_f55), .C1(n5514), .C2(
        keyinput_f53), .A(n10453), .ZN(n10465) );
  AOI22_X1 U11497 ( .A1(n10457), .A2(keyinput_f54), .B1(n10456), .B2(
        keyinput_f62), .ZN(n10455) );
  OAI221_X1 U11498 ( .B1(n10457), .B2(keyinput_f54), .C1(n10456), .C2(
        keyinput_f62), .A(n10455), .ZN(n10464) );
  XOR2_X1 U11499 ( .A(n10458), .B(keyinput_f98), .Z(n10462) );
  XOR2_X1 U11500 ( .A(n5779), .B(keyinput_f47), .Z(n10461) );
  XNOR2_X1 U11501 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_f121), .ZN(n10460)
         );
  XNOR2_X1 U11502 ( .A(SI_2_), .B(keyinput_f30), .ZN(n10459) );
  NAND4_X1 U11503 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n10463) );
  NOR3_X1 U11504 ( .A1(n10465), .A2(n10464), .A3(n10463), .ZN(n10498) );
  AOI22_X1 U11505 ( .A1(n10468), .A2(keyinput_f59), .B1(n10467), .B2(
        keyinput_f45), .ZN(n10466) );
  OAI221_X1 U11506 ( .B1(n10468), .B2(keyinput_f59), .C1(n10467), .C2(
        keyinput_f45), .A(n10466), .ZN(n10481) );
  AOI22_X1 U11507 ( .A1(n10471), .A2(keyinput_f93), .B1(n10470), .B2(
        keyinput_f39), .ZN(n10469) );
  OAI221_X1 U11508 ( .B1(n10471), .B2(keyinput_f93), .C1(n10470), .C2(
        keyinput_f39), .A(n10469), .ZN(n10480) );
  AOI22_X1 U11509 ( .A1(n10474), .A2(keyinput_f27), .B1(n10473), .B2(
        keyinput_f51), .ZN(n10472) );
  OAI221_X1 U11510 ( .B1(n10474), .B2(keyinput_f27), .C1(n10473), .C2(
        keyinput_f51), .A(n10472), .ZN(n10479) );
  INV_X1 U11511 ( .A(P2_B_REG_SCAN_IN), .ZN(n10475) );
  XOR2_X1 U11512 ( .A(n10475), .B(keyinput_f64), .Z(n10477) );
  XNOR2_X1 U11513 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_f96), .ZN(n10476) );
  NAND2_X1 U11514 ( .A1(n10477), .A2(n10476), .ZN(n10478) );
  NOR4_X1 U11515 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10497) );
  AOI22_X1 U11516 ( .A1(n6067), .A2(keyinput_f92), .B1(n10483), .B2(
        keyinput_f86), .ZN(n10482) );
  OAI221_X1 U11517 ( .B1(n6067), .B2(keyinput_f92), .C1(n10483), .C2(
        keyinput_f86), .A(n10482), .ZN(n10495) );
  AOI22_X1 U11518 ( .A1(n10486), .A2(keyinput_f95), .B1(n10485), .B2(
        keyinput_f4), .ZN(n10484) );
  OAI221_X1 U11519 ( .B1(n10486), .B2(keyinput_f95), .C1(n10485), .C2(
        keyinput_f4), .A(n10484), .ZN(n10494) );
  AOI22_X1 U11520 ( .A1(n10489), .A2(keyinput_f73), .B1(keyinput_f13), .B2(
        n10488), .ZN(n10487) );
  OAI221_X1 U11521 ( .B1(n10489), .B2(keyinput_f73), .C1(n10488), .C2(
        keyinput_f13), .A(n10487), .ZN(n10493) );
  XNOR2_X1 U11522 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput_f34), .ZN(n10491) );
  XNOR2_X1 U11523 ( .A(SI_0_), .B(keyinput_f32), .ZN(n10490) );
  NAND2_X1 U11524 ( .A1(n10491), .A2(n10490), .ZN(n10492) );
  NOR4_X1 U11525 ( .A1(n10495), .A2(n10494), .A3(n10493), .A4(n10492), .ZN(
        n10496) );
  NAND4_X1 U11526 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(
        n10500) );
  OR4_X1 U11527 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10505) );
  AOI21_X1 U11528 ( .B1(keyinput_f81), .B2(n10505), .A(keyinput_g81), .ZN(
        n10507) );
  INV_X1 U11529 ( .A(keyinput_f81), .ZN(n10504) );
  AOI21_X1 U11530 ( .B1(n10505), .B2(n10504), .A(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n10506) );
  AOI22_X1 U11531 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n10507), .B1(
        keyinput_g81), .B2(n10506), .ZN(n10508) );
  AOI21_X1 U11532 ( .B1(n10510), .B2(n10509), .A(n10508), .ZN(n10511) );
  XNOR2_X1 U11533 ( .A(n10512), .B(n10511), .ZN(n10513) );
  XNOR2_X1 U11534 ( .A(n10514), .B(n10513), .ZN(ADD_1068_U4) );
  XNOR2_X1 U11535 ( .A(n10516), .B(n10515), .ZN(ADD_1068_U47) );
  XOR2_X1 U11536 ( .A(n10518), .B(n10517), .Z(ADD_1068_U54) );
  XNOR2_X1 U11537 ( .A(n10520), .B(n10519), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11538 ( .A(n10522), .B(n10521), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11539 ( .A(n10524), .B(n10523), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11540 ( .A(n10526), .B(n10525), .ZN(ADD_1068_U50) );
  XOR2_X1 U11541 ( .A(n10528), .B(n10527), .Z(ADD_1068_U53) );
  XNOR2_X1 U11542 ( .A(n10530), .B(n10529), .ZN(ADD_1068_U52) );
  AND4_X1 U7782 ( .A1(n6103), .A2(n6102), .A3(n6101), .A4(n6100), .ZN(n7127)
         );
  NAND2_X1 U5182 ( .A1(n6805), .A2(n8027), .ZN(n8009) );
  AND2_X1 U6458 ( .A1(n6952), .A2(n6951), .ZN(n6957) );
  CLKBUF_X2 U5009 ( .A(n6056), .Z(n4518) );
  NAND2_X2 U5044 ( .A1(n5989), .A2(n9635), .ZN(n6074) );
  XNOR2_X1 U5127 ( .A(n5356), .B(n5355), .ZN(n8041) );
  CLKBUF_X1 U5234 ( .A(n9871), .Z(n4513) );
  AND2_X1 U5236 ( .A1(n5347), .A2(n5346), .ZN(n10533) );
endmodule

