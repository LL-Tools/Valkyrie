

module b20_C_gen_AntiSAT_k_128_2 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4352, n4353, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10232;

  MUX2_X1 U4857 ( .A(n8414), .B(n8413), .S(n8545), .Z(n8417) );
  INV_X1 U4858 ( .A(n5450), .ZN(n8329) );
  AOI21_X1 U4859 ( .B1(n8394), .B2(n8545), .A(n4497), .ZN(n4496) );
  BUF_X1 U4860 ( .A(n9638), .Z(n4352) );
  XNOR2_X1 U4861 ( .A(n5107), .B(n5105), .ZN(n5596) );
  OAI21_X1 U4862 ( .B1(n5616), .B2(n4414), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5135) );
  CLKBUF_X1 U4863 ( .A(n10232), .Z(P2_U3893) );
  NOR2_X1 U4864 ( .A1(n6382), .A2(n6380), .ZN(n10232) );
  INV_X1 U4866 ( .A(n9120), .ZN(n9429) );
  INV_X1 U4867 ( .A(n8331), .ZN(n5423) );
  INV_X1 U4869 ( .A(n7923), .ZN(n6081) );
  INV_X1 U4870 ( .A(n9238), .ZN(n9438) );
  INV_X1 U4871 ( .A(n8070), .ZN(n7926) );
  NAND2_X1 U4872 ( .A1(n8958), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U4873 ( .A1(n6514), .A2(n7912), .ZN(n5889) );
  NAND2_X2 U4874 ( .A1(n6269), .A2(n8095), .ZN(n7923) );
  NAND2_X1 U4875 ( .A1(n6789), .A2(n5793), .ZN(n6956) );
  OAI211_X1 U4876 ( .C1(n7923), .C2(n9151), .A(n5767), .B(n5766), .ZN(n9083)
         );
  OAI21_X1 U4877 ( .B1(n4906), .B2(n4554), .A(n4552), .ZN(n9269) );
  OAI21_X1 U4878 ( .B1(n5709), .B2(n4382), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5710) );
  NAND2_X1 U4880 ( .A1(n5695), .A2(n5694), .ZN(n8063) );
  BUF_X2 U4881 ( .A(n5758), .Z(n6072) );
  OAI21_X2 U4882 ( .B1(n8817), .B2(n8867), .A(n8799), .ZN(n5436) );
  AOI21_X1 U4883 ( .B1(n4976), .B2(n6938), .A(n4415), .ZN(n7183) );
  INV_X4 U4884 ( .A(n8336), .ZN(n5193) );
  OAI211_X2 U4885 ( .C1(n9079), .C2(n4569), .A(n4567), .B(n6791), .ZN(n6789)
         );
  NOR2_X2 U4886 ( .A1(n4388), .A2(n4582), .ZN(n4581) );
  OAI222_X1 U4887 ( .A1(n7225), .A2(P2_U3151), .B1(n8205), .B2(n6420), .C1(
        n6419), .C2(n8968), .ZN(P2_U3288) );
  OAI222_X1 U4888 ( .A1(n9536), .A2(n6418), .B1(n7754), .B2(n6420), .C1(
        P1_U3086), .C2(n6486), .ZN(P1_U3348) );
  NAND2_X4 U4889 ( .A1(n5889), .A2(n5888), .ZN(n9660) );
  OAI21_X2 U4890 ( .B1(n5684), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6044) );
  BUF_X4 U4891 ( .A(n6072), .Z(n6435) );
  OAI21_X1 U4892 ( .B1(n6420), .B2(n5765), .A(n5856), .ZN(n9638) );
  NOR2_X2 U4893 ( .A1(n7684), .A2(n7685), .ZN(n7691) );
  AOI21_X2 U4894 ( .B1(n8788), .B2(n4729), .A(n4725), .ZN(n4724) );
  OAI21_X2 U4895 ( .B1(n8287), .B2(n8808), .A(n5436), .ZN(n8788) );
  NAND2_X2 U4896 ( .A1(n5030), .A2(n5029), .ZN(n5310) );
  CLKBUF_X3 U4897 ( .A(n6770), .Z(n4353) );
  OAI211_X1 U4898 ( .C1(n5207), .C2(n4384), .A(n5219), .B(n4360), .ZN(n6770)
         );
  NAND2_X1 U4901 ( .A1(n9065), .A2(n9064), .ZN(n9063) );
  NOR2_X1 U4902 ( .A1(n9003), .A2(n9005), .ZN(n9004) );
  NAND2_X1 U4903 ( .A1(n8405), .A2(n8400), .ZN(n8356) );
  INV_X2 U4904 ( .A(n4473), .ZN(n8170) );
  NAND2_X1 U4905 ( .A1(n4521), .A2(n5027), .ZN(n5285) );
  INV_X1 U4906 ( .A(n9639), .ZN(n6896) );
  NAND2_X2 U4907 ( .A1(n8384), .A2(n8387), .ZN(n6878) );
  NAND4_X1 U4908 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n9598)
         );
  INV_X4 U4909 ( .A(n5214), .ZN(n5601) );
  INV_X2 U4910 ( .A(n5784), .ZN(n6082) );
  NAND2_X1 U4911 ( .A1(n8063), .A2(n8072), .ZN(n6340) );
  XNOR2_X1 U4912 ( .A(n5135), .B(n5134), .ZN(n8206) );
  AOI21_X1 U4913 ( .B1(n9063), .B2(n9067), .A(n8975), .ZN(n9033) );
  NOR2_X1 U4914 ( .A1(n4390), .A2(n4530), .ZN(n4529) );
  OAI21_X1 U4915 ( .B1(n9343), .B2(n9335), .A(n7863), .ZN(n9321) );
  AOI21_X1 U4916 ( .B1(n7983), .B2(n6355), .A(n6354), .ZN(n9343) );
  OAI21_X1 U4917 ( .B1(n9823), .B2(n4947), .A(n4946), .ZN(n8676) );
  NAND2_X1 U4918 ( .A1(n8649), .A2(n4948), .ZN(n4946) );
  NAND2_X1 U4919 ( .A1(n8764), .A2(n5471), .ZN(n8756) );
  NAND2_X1 U4920 ( .A1(n7777), .A2(n6002), .ZN(n4593) );
  NAND2_X1 U4921 ( .A1(n7600), .A2(n7599), .ZN(n7598) );
  NAND2_X1 U4922 ( .A1(n5405), .A2(n5404), .ZN(n7734) );
  AND2_X1 U4923 ( .A1(n7430), .A2(n7836), .ZN(n7600) );
  NAND2_X1 U4924 ( .A1(n4742), .A2(n4741), .ZN(n7704) );
  NAND2_X1 U4925 ( .A1(n7294), .A2(n7293), .ZN(n7296) );
  AOI21_X1 U4926 ( .B1(n4548), .B2(n4549), .A(n4413), .ZN(n4547) );
  OR2_X1 U4927 ( .A1(n5317), .A2(n7154), .ZN(n7265) );
  NAND2_X1 U4928 ( .A1(n5675), .A2(n5674), .ZN(n7292) );
  AND2_X1 U4929 ( .A1(n5314), .A2(n5313), .ZN(n9909) );
  NAND2_X2 U4930 ( .A1(n5871), .A2(n5870), .ZN(n6310) );
  NAND2_X1 U4931 ( .A1(n7819), .A2(n7804), .ZN(n7817) );
  AND3_X1 U4932 ( .A1(n5290), .A2(n5289), .A3(n5288), .ZN(n9903) );
  XNOR2_X1 U4933 ( .A(n5285), .B(n5284), .ZN(n6420) );
  CLKBUF_X1 U4934 ( .A(n4473), .Z(n4456) );
  NAND2_X2 U4935 ( .A1(n4998), .A2(n6674), .ZN(n4473) );
  INV_X2 U4936 ( .A(n9393), .ZN(n9571) );
  AND2_X1 U4937 ( .A1(n6700), .A2(n6703), .ZN(n6727) );
  NAND2_X1 U4938 ( .A1(n6878), .A2(n6881), .ZN(n9848) );
  NAND4_X1 U4939 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(n9639)
         );
  NAND2_X1 U4940 ( .A1(n8663), .A2(n8375), .ZN(n4998) );
  NAND4_X1 U4941 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n9127)
         );
  NAND4_X2 U4942 ( .A1(n4810), .A2(n4809), .A3(n4808), .A4(n4807), .ZN(n9599)
         );
  NAND4_X1 U4943 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n8585)
         );
  OAI211_X1 U4944 ( .C1(n7923), .C2(n9159), .A(n5785), .B(n4898), .ZN(n9609)
         );
  INV_X2 U4945 ( .A(n6220), .ZN(n6433) );
  AND3_X1 U4946 ( .A1(n5210), .A2(n5209), .A3(n5208), .ZN(n9861) );
  AND2_X2 U4947 ( .A1(n8126), .A2(n8206), .ZN(n5214) );
  NAND2_X1 U4948 ( .A1(n7923), .A2(n7922), .ZN(n5765) );
  NAND2_X1 U4949 ( .A1(n6763), .A2(n6607), .ZN(n6608) );
  AND2_X1 U4950 ( .A1(n8006), .A2(n8064), .ZN(n5722) );
  AND2_X1 U4951 ( .A1(n6263), .A2(n5683), .ZN(n8072) );
  OR2_X2 U4952 ( .A1(n5708), .A2(n7720), .ZN(n6273) );
  NAND2_X1 U4953 ( .A1(n5700), .A2(n5699), .ZN(n8064) );
  NAND2_X1 U4954 ( .A1(n5707), .A2(n4374), .ZN(n7720) );
  XNOR2_X1 U4955 ( .A(n5696), .B(P1_IR_REG_21__SCAN_IN), .ZN(n8006) );
  AND2_X1 U4956 ( .A1(n5691), .A2(n5690), .ZN(n5695) );
  NOR2_X1 U4957 ( .A1(n5616), .A2(n4488), .ZN(n4487) );
  OAI21_X1 U4958 ( .B1(n5706), .B2(n4416), .A(n4370), .ZN(n5707) );
  NAND2_X1 U4959 ( .A1(n5699), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5696) );
  OR2_X1 U4960 ( .A1(n5697), .A2(n9527), .ZN(n5698) );
  NAND2_X1 U4961 ( .A1(n5697), .A2(n5679), .ZN(n5699) );
  NAND2_X2 U4962 ( .A1(n7917), .A2(P1_U3086), .ZN(n9536) );
  INV_X1 U4963 ( .A(n5011), .ZN(n5004) );
  NAND2_X1 U4964 ( .A1(n4371), .A2(n4753), .ZN(n4488) );
  BUF_X1 U4965 ( .A(n5671), .Z(n5854) );
  AND2_X2 U4966 ( .A1(n4533), .A2(n4532), .ZN(n5011) );
  NOR2_X1 U4967 ( .A1(n5221), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n4952) );
  AND4_X1 U4968 ( .A1(n5663), .A2(n5662), .A3(n5680), .A4(n5676), .ZN(n4365)
         );
  CLKBUF_X2 U4969 ( .A(n5184), .Z(n5207) );
  INV_X1 U4970 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4654) );
  INV_X2 U4971 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4563) );
  NOR2_X1 U4972 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5093) );
  NOR2_X1 U4973 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5095) );
  INV_X1 U4974 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6062) );
  INV_X1 U4975 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5680) );
  INV_X4 U4976 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U4977 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5663) );
  OR2_X1 U4978 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  NAND4_X2 U4979 ( .A1(n4862), .A2(n4861), .A3(n4860), .A4(n4859), .ZN(n5661)
         );
  OAI21_X1 U4980 ( .B1(n9033), .B2(n4485), .A(n4465), .ZN(n4464) );
  BUF_X4 U4981 ( .A(n6172), .Z(n4356) );
  INV_X1 U4982 ( .A(n8182), .ZN(n6172) );
  AOI21_X2 U4983 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n9817), .A(n9808), .ZN(
        n8647) );
  NAND2_X1 U4984 ( .A1(n7848), .A2(n8070), .ZN(n4818) );
  INV_X1 U4985 ( .A(n9409), .ZN(n4820) );
  NAND2_X1 U4986 ( .A1(n9328), .A2(n9304), .ZN(n4561) );
  XNOR2_X1 U4987 ( .A(n7904), .B(n7902), .ZN(n7901) );
  NAND2_X1 U4988 ( .A1(n4781), .A2(n4790), .ZN(n4780) );
  AND2_X1 U4989 ( .A1(n7854), .A2(n8035), .ZN(n4817) );
  INV_X1 U4990 ( .A(n8520), .ZN(n4492) );
  INV_X1 U4991 ( .A(n8736), .ZN(n5591) );
  NAND2_X1 U4992 ( .A1(n4688), .A2(n4687), .ZN(n7904) );
  AOI21_X1 U4993 ( .B1(n4690), .B2(n4692), .A(n4448), .ZN(n4687) );
  NOR2_X1 U4994 ( .A1(n5419), .A2(n4683), .ZN(n4682) );
  INV_X1 U4995 ( .A(n5059), .ZN(n4683) );
  INV_X1 U4996 ( .A(n5406), .ZN(n5058) );
  NOR2_X1 U4997 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4862) );
  AOI21_X1 U4998 ( .B1(n4666), .B2(n5048), .A(n5363), .ZN(n4665) );
  NOR2_X1 U4999 ( .A1(n5001), .A2(n4738), .ZN(n4737) );
  INV_X1 U5000 ( .A(n5483), .ZN(n4738) );
  INV_X1 U5001 ( .A(n8778), .ZN(n4733) );
  NAND2_X1 U5002 ( .A1(n4750), .A2(n5104), .ZN(n4754) );
  NOR3_X1 U5003 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n5104) );
  OAI21_X1 U5004 ( .B1(n5616), .B2(P2_IR_REG_26__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5107) );
  OR2_X1 U5005 ( .A1(n9433), .A2(n9442), .ZN(n4610) );
  NOR2_X1 U5006 ( .A1(n9312), .A2(n4398), .ZN(n4883) );
  OR2_X1 U5007 ( .A1(n9464), .A2(n9325), .ZN(n7871) );
  NAND2_X1 U5008 ( .A1(n4408), .A2(n4561), .ZN(n4558) );
  NAND2_X1 U5009 ( .A1(n9096), .A2(n9498), .ZN(n4910) );
  AND2_X1 U5010 ( .A1(n4542), .A2(n4362), .ZN(n4540) );
  NAND2_X1 U5011 ( .A1(n4422), .A2(n4362), .ZN(n4539) );
  NAND2_X1 U5012 ( .A1(n7437), .A2(n7408), .ZN(n4920) );
  NAND2_X1 U5013 ( .A1(n7946), .A2(n7833), .ZN(n4888) );
  AND2_X1 U5014 ( .A1(n7815), .A2(n8013), .ZN(n7939) );
  NAND2_X1 U5015 ( .A1(n4669), .A2(n4667), .ZN(n7916) );
  AND2_X1 U5016 ( .A1(n7905), .A2(n4668), .ZN(n4667) );
  INV_X1 U5017 ( .A(n7909), .ZN(n4668) );
  NAND2_X1 U5018 ( .A1(n4653), .A2(n5087), .ZN(n5485) );
  NAND2_X1 U5019 ( .A1(n5706), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5682) );
  INV_X1 U5020 ( .A(n4706), .ZN(n4705) );
  AOI21_X1 U5021 ( .B1(n4706), .B2(n4704), .A(n4703), .ZN(n4702) );
  INV_X1 U5022 ( .A(n5078), .ZN(n4703) );
  NAND2_X1 U5023 ( .A1(n4659), .A2(n4655), .ZN(n5390) );
  INV_X1 U5024 ( .A(n4656), .ZN(n4655) );
  OAI21_X1 U5025 ( .B1(n4661), .B2(n4657), .A(n5053), .ZN(n4656) );
  OAI21_X1 U5026 ( .B1(n5336), .B2(n5335), .A(n5045), .ZN(n5349) );
  NAND2_X1 U5027 ( .A1(n8162), .A2(n8242), .ZN(n8244) );
  NOR2_X1 U5028 ( .A1(n6941), .A2(n4977), .ZN(n4976) );
  XNOR2_X1 U5029 ( .A(n6886), .B(n4473), .ZN(n6798) );
  XNOR2_X1 U5030 ( .A(n8647), .B(n8648), .ZN(n9823) );
  AOI21_X1 U5031 ( .B1(n4377), .B2(n4758), .A(n4757), .ZN(n4756) );
  NAND2_X1 U5032 ( .A1(n8733), .A2(n4400), .ZN(n4755) );
  OR2_X1 U5033 ( .A1(n5442), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5453) );
  NAND2_X1 U5034 ( .A1(n5187), .A2(n7917), .ZN(n5450) );
  CLKBUF_X2 U5035 ( .A(n5226), .Z(n8331) );
  AOI21_X1 U5036 ( .B1(n4743), .B2(n4749), .A(n4407), .ZN(n4741) );
  NOR2_X1 U5037 ( .A1(n6583), .A2(n6842), .ZN(n6572) );
  XNOR2_X1 U5038 ( .A(n5561), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8381) );
  NAND2_X1 U5039 ( .A1(n5169), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U5040 ( .A1(n9569), .A2(n6174), .ZN(n5866) );
  NAND2_X1 U5041 ( .A1(n5929), .A2(n5930), .ZN(n5933) );
  NOR2_X1 U5042 ( .A1(n4431), .A2(n4591), .ZN(n4590) );
  INV_X1 U5043 ( .A(n6126), .ZN(n4591) );
  NAND2_X1 U5044 ( .A1(n4421), .A2(n6198), .ZN(n4864) );
  OR2_X1 U5045 ( .A1(n6272), .A2(n6406), .ZN(n6278) );
  NAND2_X1 U5046 ( .A1(n6330), .A2(n6329), .ZN(n8114) );
  OR2_X1 U5047 ( .A1(n9322), .A2(n9464), .ZN(n9302) );
  NAND2_X1 U5048 ( .A1(n9336), .A2(n4907), .ZN(n4906) );
  NAND2_X1 U5049 ( .A1(n9337), .A2(n9071), .ZN(n4907) );
  NOR2_X1 U5050 ( .A1(n9501), .A2(n9381), .ZN(n4913) );
  OR2_X1 U5051 ( .A1(n9617), .A2(n9626), .ZN(n7815) );
  NAND2_X1 U5052 ( .A1(n6379), .A2(n6273), .ZN(n6406) );
  AND2_X1 U5053 ( .A1(n8063), .A2(n8064), .ZN(n8079) );
  INV_X1 U5054 ( .A(n8120), .ZN(n4531) );
  NAND2_X1 U5055 ( .A1(n6026), .A2(n6025), .ZN(n9507) );
  NAND2_X1 U5056 ( .A1(n6361), .A2(n6360), .ZN(n9666) );
  NAND2_X1 U5057 ( .A1(n7309), .A2(n7308), .ZN(n7370) );
  NAND2_X1 U5058 ( .A1(n7306), .A2(n7307), .ZN(n7308) );
  INV_X1 U5059 ( .A(n8585), .ZN(n7307) );
  NOR2_X1 U5060 ( .A1(n9828), .A2(n8829), .ZN(n9827) );
  AOI21_X1 U5061 ( .B1(n9100), .B2(n4436), .A(n4853), .ZN(n4570) );
  AND2_X1 U5062 ( .A1(n9100), .A2(n4372), .ZN(n8197) );
  INV_X1 U5063 ( .A(n9119), .ZN(n9084) );
  AND2_X1 U5064 ( .A1(n8393), .A2(n8554), .ZN(n4497) );
  MUX2_X1 U5065 ( .A(n8386), .B(n8385), .S(n8554), .Z(n8396) );
  NAND2_X1 U5066 ( .A1(n7797), .A2(n7926), .ZN(n4815) );
  NOR2_X1 U5067 ( .A1(n4800), .A2(n4799), .ZN(n4798) );
  INV_X1 U5068 ( .A(n7815), .ZN(n4800) );
  INV_X1 U5069 ( .A(n7818), .ZN(n4797) );
  NAND2_X1 U5070 ( .A1(n7822), .A2(n8070), .ZN(n4801) );
  AOI21_X1 U5071 ( .B1(n4790), .B2(n4789), .A(n7926), .ZN(n4788) );
  INV_X1 U5072 ( .A(n8023), .ZN(n4789) );
  NAND2_X1 U5073 ( .A1(n4418), .A2(n7834), .ZN(n4792) );
  NAND2_X1 U5074 ( .A1(n4780), .A2(n4788), .ZN(n4787) );
  NAND2_X1 U5075 ( .A1(n4782), .A2(n4381), .ZN(n4785) );
  NAND2_X1 U5076 ( .A1(n4784), .A2(n4783), .ZN(n7842) );
  INV_X1 U5077 ( .A(n7796), .ZN(n4816) );
  NAND2_X1 U5078 ( .A1(n7850), .A2(n4481), .ZN(n4779) );
  INV_X1 U5079 ( .A(n7861), .ZN(n4777) );
  NOR2_X1 U5080 ( .A1(n4806), .A2(n4805), .ZN(n4804) );
  NAND2_X1 U5081 ( .A1(n7986), .A2(n8070), .ZN(n4805) );
  INV_X1 U5082 ( .A(n8606), .ZN(n4516) );
  OR2_X1 U5083 ( .A1(n8585), .A2(n9903), .ZN(n8424) );
  INV_X1 U5084 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5155) );
  INV_X1 U5085 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5376) );
  INV_X1 U5086 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5676) );
  AND2_X1 U5087 ( .A1(n4678), .A2(n5164), .ZN(n4676) );
  INV_X1 U5088 ( .A(SI_17_), .ZN(n5062) );
  INV_X1 U5089 ( .A(n4662), .ZN(n4661) );
  AND2_X1 U5090 ( .A1(n4701), .A2(n4997), .ZN(n4700) );
  NAND2_X1 U5091 ( .A1(n5309), .A2(n5036), .ZN(n4701) );
  INV_X1 U5092 ( .A(n8144), .ZN(n4967) );
  NAND2_X1 U5093 ( .A1(n8294), .A2(n8150), .ZN(n8152) );
  NOR2_X1 U5094 ( .A1(n8142), .A2(n4973), .ZN(n4972) );
  INV_X1 U5095 ( .A(n8139), .ZN(n4973) );
  NAND2_X1 U5096 ( .A1(n8558), .A2(n8543), .ZN(n4670) );
  NOR2_X1 U5097 ( .A1(n8552), .A2(n4673), .ZN(n4672) );
  NAND2_X1 U5098 ( .A1(n4387), .A2(n8375), .ZN(n4673) );
  INV_X1 U5099 ( .A(n4670), .ZN(n8347) );
  OR2_X1 U5100 ( .A1(n8542), .A2(n8541), .ZN(n8553) );
  NAND2_X1 U5101 ( .A1(n4510), .A2(n4509), .ZN(n7465) );
  NAND2_X1 U5102 ( .A1(n7320), .A2(n7464), .ZN(n4509) );
  NAND2_X1 U5103 ( .A1(n4513), .A2(n4394), .ZN(n4510) );
  OAI21_X1 U5104 ( .B1(n7505), .B2(n4519), .A(n4517), .ZN(n8603) );
  OR2_X1 U5105 ( .A1(n4834), .A2(n4518), .ZN(n4517) );
  NAND2_X1 U5106 ( .A1(n4376), .A2(n7581), .ZN(n4519) );
  INV_X1 U5107 ( .A(n7581), .ZN(n4518) );
  OR2_X1 U5108 ( .A1(n5413), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U5109 ( .A1(n5119), .A2(n10158), .ZN(n5413) );
  INV_X1 U5110 ( .A(n5397), .ZN(n5119) );
  OR2_X1 U5111 ( .A1(n7191), .A2(n5315), .ZN(n7266) );
  AND2_X1 U5112 ( .A1(n4635), .A2(n8415), .ZN(n4634) );
  NAND2_X1 U5113 ( .A1(n7250), .A2(n4636), .ZN(n4635) );
  AND2_X1 U5114 ( .A1(n5316), .A2(n7150), .ZN(n7154) );
  NAND2_X1 U5115 ( .A1(n8424), .A2(n7160), .ZN(n8416) );
  INV_X1 U5116 ( .A(n8405), .ZN(n4617) );
  NOR2_X1 U5117 ( .A1(n4617), .A2(n8401), .ZN(n4616) );
  OR2_X1 U5118 ( .A1(n9837), .A2(n9861), .ZN(n8390) );
  OR2_X1 U5119 ( .A1(n6675), .A2(n9872), .ZN(n8384) );
  NOR2_X1 U5120 ( .A1(n4385), .A2(n4767), .ZN(n4766) );
  NAND2_X1 U5121 ( .A1(n8327), .A2(n5591), .ZN(n4770) );
  INV_X1 U5122 ( .A(n4648), .ZN(n4646) );
  NAND2_X1 U5123 ( .A1(n4737), .A2(n4735), .ZN(n4734) );
  INV_X1 U5124 ( .A(n5000), .ZN(n4735) );
  OR2_X1 U5125 ( .A1(n8907), .A2(n8158), .ZN(n8523) );
  INV_X1 U5126 ( .A(n4640), .ZN(n4639) );
  OR2_X1 U5127 ( .A1(n8260), .A2(n8269), .ZN(n8471) );
  NOR2_X1 U5128 ( .A1(n5581), .A2(n4627), .ZN(n4626) );
  INV_X1 U5129 ( .A(n8465), .ZN(n4627) );
  NOR2_X1 U5130 ( .A1(n5387), .A2(n4744), .ZN(n4743) );
  INV_X1 U5131 ( .A(n4746), .ZN(n4744) );
  NAND2_X1 U5132 ( .A1(n7266), .A2(n5318), .ZN(n5333) );
  AND2_X1 U5133 ( .A1(n7267), .A2(n7265), .ZN(n5318) );
  NOR2_X1 U5134 ( .A1(n4723), .A2(n4719), .ZN(n4718) );
  INV_X1 U5135 ( .A(n5346), .ZN(n4723) );
  NAND2_X1 U5136 ( .A1(n5346), .A2(n4722), .ZN(n4721) );
  INV_X1 U5137 ( .A(n5334), .ZN(n4722) );
  NAND2_X1 U5138 ( .A1(n8572), .A2(n8381), .ZN(n8545) );
  INV_X1 U5139 ( .A(n8566), .ZN(n6673) );
  OR2_X1 U5140 ( .A1(n6901), .A2(n6902), .ZN(n4585) );
  NAND2_X1 U5141 ( .A1(n6901), .A2(n6902), .ZN(n4584) );
  NAND2_X1 U5142 ( .A1(n8079), .A2(n7593), .ZN(n4586) );
  INV_X1 U5143 ( .A(n5722), .ZN(n5701) );
  INV_X1 U5144 ( .A(n4584), .ZN(n4583) );
  INV_X1 U5145 ( .A(n9271), .ZN(n4885) );
  AOI21_X1 U5146 ( .B1(n4903), .B2(n4901), .A(n4417), .ZN(n4900) );
  INV_X1 U5147 ( .A(n6322), .ZN(n4901) );
  NOR2_X1 U5148 ( .A1(n4902), .A2(n4556), .ZN(n4555) );
  INV_X1 U5149 ( .A(n4558), .ZN(n4556) );
  INV_X1 U5150 ( .A(n4903), .ZN(n4902) );
  INV_X1 U5151 ( .A(n9289), .ZN(n4880) );
  NOR2_X1 U5152 ( .A1(n9479), .A2(n4601), .ZN(n4600) );
  INV_X1 U5153 ( .A(n4602), .ZN(n4601) );
  OR2_X1 U5154 ( .A1(n9494), .A2(n9498), .ZN(n7854) );
  NAND2_X1 U5155 ( .A1(n7821), .A2(n7804), .ZN(n6350) );
  AND2_X1 U5156 ( .A1(n7055), .A2(n6304), .ZN(n6306) );
  AND2_X1 U5157 ( .A1(n7937), .A2(n7815), .ZN(n4896) );
  OR2_X1 U5158 ( .A1(n6896), .A2(n9577), .ZN(n7818) );
  NAND2_X1 U5159 ( .A1(n4899), .A2(n9609), .ZN(n7809) );
  INV_X1 U5160 ( .A(n9598), .ZN(n4899) );
  NAND2_X1 U5161 ( .A1(n8008), .A2(n6344), .ZN(n7021) );
  AOI21_X1 U5162 ( .B1(n6405), .B2(n6252), .A(n6411), .ZN(n6741) );
  INV_X1 U5163 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U5164 ( .A1(n5682), .A2(n5681), .ZN(n6263) );
  OR2_X1 U5165 ( .A1(n5076), .A2(n10148), .ZN(n4709) );
  NOR2_X1 U5166 ( .A1(n5060), .A2(n4686), .ZN(n4685) );
  INV_X1 U5167 ( .A(n5056), .ZN(n4686) );
  AOI21_X1 U5168 ( .B1(n4700), .B2(n4698), .A(n4697), .ZN(n4696) );
  INV_X1 U5169 ( .A(n5040), .ZN(n4697) );
  INV_X1 U5170 ( .A(n5036), .ZN(n4698) );
  INV_X1 U5171 ( .A(n4700), .ZN(n4699) );
  NAND2_X1 U5172 ( .A1(n5285), .A2(n5284), .ZN(n5030) );
  OAI21_X1 U5173 ( .B1(n5004), .B2(n5003), .A(n5002), .ZN(n5008) );
  INV_X1 U5174 ( .A(SI_10_), .ZN(n10038) );
  NAND2_X1 U5175 ( .A1(n8153), .A2(n8508), .ZN(n4987) );
  NAND2_X1 U5176 ( .A1(n8314), .A2(n4964), .ZN(n4963) );
  INV_X1 U5177 ( .A(n8163), .ZN(n4964) );
  INV_X1 U5178 ( .A(n8314), .ZN(n4965) );
  AND2_X1 U5179 ( .A1(n8163), .A2(n8161), .ZN(n8242) );
  NAND2_X1 U5180 ( .A1(n8252), .A2(n8133), .ZN(n8265) );
  NAND2_X1 U5181 ( .A1(n8132), .A2(n8269), .ZN(n8133) );
  OR2_X1 U5182 ( .A1(n8152), .A2(n8151), .ZN(n8274) );
  NAND2_X1 U5183 ( .A1(n8140), .A2(n4972), .ZN(n4971) );
  OR2_X1 U5184 ( .A1(n7615), .A2(n7614), .ZN(n7616) );
  NAND2_X1 U5185 ( .A1(n8265), .A2(n8264), .ZN(n8263) );
  AND2_X1 U5186 ( .A1(n5102), .A2(n4983), .ZN(n4982) );
  INV_X1 U5187 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5102) );
  INV_X1 U5188 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4983) );
  OR2_X1 U5189 ( .A1(n5429), .A2(n5178), .ZN(n5180) );
  AND2_X1 U5190 ( .A1(n6833), .A2(n4934), .ZN(n4933) );
  XNOR2_X1 U5191 ( .A(n7465), .B(n7466), .ZN(n7506) );
  NOR2_X1 U5192 ( .A1(n7506), .A2(n7451), .ZN(n7505) );
  AND2_X1 U5193 ( .A1(n4928), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4925) );
  INV_X1 U5194 ( .A(n9784), .ZN(n4832) );
  OAI21_X1 U5195 ( .B1(n8591), .B2(n4941), .A(n4940), .ZN(n9808) );
  NAND2_X1 U5196 ( .A1(n4944), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4941) );
  INV_X1 U5197 ( .A(n9809), .ZN(n4944) );
  OR2_X1 U5198 ( .A1(n8591), .A2(n8590), .ZN(n4943) );
  NAND2_X1 U5199 ( .A1(n4948), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4947) );
  INV_X1 U5200 ( .A(n8651), .ZN(n4948) );
  AND2_X1 U5201 ( .A1(n8483), .A2(n8484), .ZN(n8803) );
  INV_X1 U5202 ( .A(n8578), .ZN(n7756) );
  NAND2_X1 U5203 ( .A1(n7284), .A2(n8430), .ZN(n4630) );
  NAND2_X1 U5204 ( .A1(n5333), .A2(n7274), .ZN(n7269) );
  NAND2_X1 U5205 ( .A1(n7014), .A2(n8356), .ZN(n4716) );
  NOR2_X1 U5206 ( .A1(n6403), .A2(n4713), .ZN(n4712) );
  NAND2_X1 U5207 ( .A1(n8663), .A2(n8566), .ZN(n8562) );
  NAND2_X1 U5208 ( .A1(n6382), .A2(n6587), .ZN(n6842) );
  OR2_X1 U5209 ( .A1(n8528), .A2(n4396), .ZN(n8725) );
  AOI21_X1 U5210 ( .B1(n8492), .B2(n8524), .A(n4649), .ZN(n4648) );
  INV_X1 U5211 ( .A(n8523), .ZN(n4649) );
  NOR2_X1 U5212 ( .A1(n4651), .A2(n5590), .ZN(n4650) );
  INV_X1 U5213 ( .A(n4652), .ZN(n4651) );
  INV_X1 U5214 ( .A(n8725), .ZN(n8723) );
  AND2_X1 U5215 ( .A1(n8505), .A2(n8506), .ZN(n4652) );
  OR2_X1 U5216 ( .A1(n8754), .A2(n8491), .ZN(n5589) );
  AND2_X1 U5217 ( .A1(n5475), .A2(n5474), .ZN(n8512) );
  INV_X1 U5218 ( .A(n4730), .ZN(n4729) );
  OAI21_X1 U5219 ( .B1(n4731), .B2(n4733), .A(n5460), .ZN(n4730) );
  INV_X1 U5220 ( .A(n4724), .ZN(n8764) );
  INV_X1 U5221 ( .A(n4726), .ZN(n4725) );
  AOI21_X1 U5222 ( .B1(n4729), .B2(n4731), .A(n4727), .ZN(n4726) );
  NAND2_X1 U5223 ( .A1(n8777), .A2(n4732), .ZN(n4731) );
  NAND2_X1 U5224 ( .A1(n8352), .A2(n4733), .ZN(n4732) );
  AOI21_X1 U5225 ( .B1(n8788), .B2(n4733), .A(n4731), .ZN(n4728) );
  NOR2_X1 U5226 ( .A1(n8485), .A2(n4641), .ZN(n4640) );
  NOR2_X1 U5227 ( .A1(n8788), .A2(n8352), .ZN(n8789) );
  NAND2_X1 U5228 ( .A1(n8804), .A2(n8803), .ZN(n8802) );
  NAND2_X1 U5229 ( .A1(n5163), .A2(n5162), .ZN(n8867) );
  AOI22_X1 U5230 ( .A1(n7734), .A2(n8368), .B1(n8826), .B2(n8260), .ZN(n8825)
         );
  AND2_X1 U5231 ( .A1(n8811), .A2(n8475), .ZN(n8824) );
  AOI21_X1 U5232 ( .B1(n4626), .B2(n4624), .A(n4623), .ZN(n4622) );
  INV_X1 U5233 ( .A(n8466), .ZN(n4624) );
  INV_X1 U5234 ( .A(n8471), .ZN(n4623) );
  INV_X1 U5235 ( .A(n8454), .ZN(n4749) );
  AOI21_X1 U5236 ( .B1(n8454), .B2(n4748), .A(n4747), .ZN(n4746) );
  INV_X1 U5237 ( .A(n5362), .ZN(n4748) );
  INV_X1 U5238 ( .A(n8457), .ZN(n4747) );
  INV_X1 U5239 ( .A(n8703), .ZN(n9853) );
  AND2_X1 U5240 ( .A1(n8454), .A2(n8457), .ZN(n8367) );
  NAND2_X1 U5241 ( .A1(n6676), .A2(n8554), .ZN(n8703) );
  NAND2_X1 U5242 ( .A1(n5361), .A2(n5360), .ZN(n7548) );
  AND3_X1 U5243 ( .A1(n5244), .A2(n5243), .A3(n5242), .ZN(n9889) );
  OR2_X1 U5244 ( .A1(n6845), .A2(n6842), .ZN(n6677) );
  XNOR2_X1 U5245 ( .A(n5106), .B(n5130), .ZN(n5595) );
  OR2_X1 U5246 ( .A1(n5131), .A2(n5133), .ZN(n5106) );
  AND3_X1 U5247 ( .A1(n5153), .A2(n4752), .A3(n4751), .ZN(n5131) );
  INV_X1 U5248 ( .A(n5596), .ZN(n8664) );
  NAND2_X1 U5249 ( .A1(n5609), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5611) );
  INV_X1 U5250 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5610) );
  INV_X1 U5251 ( .A(n7779), .ZN(n6001) );
  NOR2_X1 U5252 ( .A1(n6403), .A2(n7917), .ZN(n4595) );
  OR2_X1 U5253 ( .A1(n7923), .A2(n6459), .ZN(n4596) );
  OR2_X1 U5254 ( .A1(n5873), .A2(n5872), .ZN(n5891) );
  NOR2_X1 U5255 ( .A1(n7238), .A2(n5937), .ZN(n4993) );
  INV_X1 U5256 ( .A(n8079), .ZN(n6341) );
  NAND2_X1 U5257 ( .A1(n4434), .A2(n9108), .ZN(n9107) );
  NAND2_X1 U5258 ( .A1(n6072), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U5259 ( .A1(n4890), .A2(n4891), .ZN(n5684) );
  AOI21_X1 U5260 ( .B1(n4874), .B2(n6357), .A(n4873), .ZN(n4872) );
  INV_X1 U5261 ( .A(n7986), .ZN(n4873) );
  OR2_X1 U5262 ( .A1(n9243), .A2(n4877), .ZN(n4923) );
  NAND2_X1 U5263 ( .A1(n6237), .A2(n6236), .ZN(n9433) );
  OAI21_X1 U5264 ( .B1(n6324), .B2(n6323), .A(n4991), .ZN(n9256) );
  NOR2_X1 U5265 ( .A1(n9281), .A2(n9262), .ZN(n6323) );
  INV_X1 U5266 ( .A(n9269), .ZN(n6324) );
  INV_X1 U5267 ( .A(n9447), .ZN(n9430) );
  AND2_X1 U5268 ( .A1(n9289), .A2(n4391), .ZN(n4903) );
  NAND2_X1 U5269 ( .A1(n9321), .A2(n4883), .ZN(n4881) );
  AOI21_X1 U5270 ( .B1(n4883), .B2(n6356), .A(n7873), .ZN(n4882) );
  NAND2_X1 U5271 ( .A1(n4557), .A2(n4558), .ZN(n9301) );
  NAND2_X1 U5272 ( .A1(n4906), .A2(n4559), .ZN(n4557) );
  INV_X1 U5273 ( .A(n9469), .ZN(n9325) );
  NAND2_X1 U5274 ( .A1(n9479), .A2(n9468), .ZN(n4905) );
  AOI21_X1 U5275 ( .B1(n4909), .B2(n4435), .A(n4908), .ZN(n9336) );
  NOR2_X1 U5276 ( .A1(n9483), .A2(n9362), .ZN(n4908) );
  INV_X1 U5277 ( .A(n9355), .ZN(n4909) );
  NAND2_X1 U5278 ( .A1(n4423), .A2(n4910), .ZN(n4548) );
  NAND2_X1 U5279 ( .A1(n4910), .A2(n4550), .ZN(n4549) );
  INV_X1 U5280 ( .A(n4913), .ZN(n4550) );
  AND2_X1 U5281 ( .A1(n7982), .A2(n8039), .ZN(n9372) );
  INV_X1 U5282 ( .A(n9395), .ZN(n4914) );
  AOI21_X1 U5283 ( .B1(n6318), .B2(n7609), .A(n4919), .ZN(n7657) );
  AOI21_X1 U5284 ( .B1(n4543), .B2(n4393), .A(n4538), .ZN(n4919) );
  OAI21_X1 U5285 ( .B1(n4539), .B2(n7609), .A(n9121), .ZN(n4538) );
  NAND2_X1 U5286 ( .A1(n4886), .A2(n4887), .ZN(n7432) );
  AOI21_X1 U5287 ( .B1(n4364), .B2(n4888), .A(n7840), .ZN(n4887) );
  OR2_X1 U5288 ( .A1(n9696), .A2(n9686), .ZN(n4544) );
  INV_X1 U5289 ( .A(n7947), .ZN(n4542) );
  OR2_X1 U5290 ( .A1(n6352), .A2(n4888), .ZN(n7425) );
  NAND2_X1 U5291 ( .A1(n7112), .A2(n6314), .ZN(n4534) );
  NAND2_X1 U5292 ( .A1(n6346), .A2(n7939), .ZN(n6965) );
  OAI21_X1 U5293 ( .B1(n6923), .B2(n6924), .A(n6298), .ZN(n7023) );
  NAND2_X1 U5294 ( .A1(n6929), .A2(n6343), .ZN(n7022) );
  NAND2_X1 U5295 ( .A1(n6923), .A2(n6930), .ZN(n6929) );
  NOR2_X1 U5296 ( .A1(n9127), .A2(n6925), .ZN(n6930) );
  NAND2_X1 U5297 ( .A1(n5722), .A2(n8108), .ZN(n6971) );
  NAND2_X1 U5298 ( .A1(n8114), .A2(n9708), .ZN(n4597) );
  INV_X1 U5299 ( .A(n9262), .ZN(n9439) );
  NAND2_X1 U5300 ( .A1(n6186), .A2(n6185), .ZN(n9456) );
  NAND2_X1 U5301 ( .A1(n6046), .A2(n6045), .ZN(n9501) );
  NAND2_X1 U5302 ( .A1(n7995), .A2(n6452), .ZN(n9705) );
  INV_X1 U5303 ( .A(n9705), .ZN(n9659) );
  INV_X1 U5304 ( .A(n9703), .ZN(n9695) );
  INV_X1 U5305 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5664) );
  INV_X1 U5306 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5665) );
  XNOR2_X1 U5307 ( .A(n7921), .B(n7920), .ZN(n8957) );
  NAND2_X1 U5308 ( .A1(n4669), .A2(n7905), .ZN(n7910) );
  AND2_X1 U5309 ( .A1(n5679), .A2(n5680), .ZN(n4869) );
  AND2_X1 U5310 ( .A1(n4710), .A2(n4708), .ZN(n4706) );
  INV_X1 U5311 ( .A(n5446), .ZN(n4710) );
  NAND2_X1 U5312 ( .A1(n5439), .A2(n4709), .ZN(n4707) );
  NAND2_X1 U5313 ( .A1(n5076), .A2(n10148), .ZN(n4708) );
  OAI21_X1 U5314 ( .B1(n5057), .B2(n4681), .A(n4678), .ZN(n5165) );
  NAND2_X1 U5315 ( .A1(n5057), .A2(n5056), .ZN(n5408) );
  OAI21_X1 U5316 ( .B1(n5349), .B2(n4664), .A(n4662), .ZN(n5375) );
  AOI21_X1 U5317 ( .B1(n4917), .B2(n5255), .A(n4410), .ZN(n4916) );
  OR3_X1 U5318 ( .A1(n5625), .A2(n7772), .A3(n5619), .ZN(n6382) );
  INV_X1 U5319 ( .A(n5187), .ZN(n6384) );
  AOI21_X1 U5320 ( .B1(n6852), .B2(n6851), .A(n6850), .ZN(n6854) );
  AND2_X1 U5321 ( .A1(n6849), .A2(n6848), .ZN(n6850) );
  XNOR2_X1 U5322 ( .A(n6798), .B(n6675), .ZN(n6800) );
  INV_X1 U5323 ( .A(n6886), .ZN(n9872) );
  AND2_X1 U5324 ( .A1(n5445), .A2(n5444), .ZN(n8236) );
  AND2_X1 U5325 ( .A1(n5495), .A2(n5494), .ZN(n8514) );
  NAND2_X1 U5326 ( .A1(n6854), .A2(n6853), .ZN(n6938) );
  NAND2_X1 U5327 ( .A1(n9854), .A2(n4979), .ZN(n4978) );
  AND4_X1 U5328 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n7674)
         );
  AOI21_X1 U5329 ( .B1(n7370), .B2(n7369), .A(n4992), .ZN(n7372) );
  INV_X1 U5330 ( .A(n8817), .ZN(n8287) );
  NAND2_X1 U5331 ( .A1(n6575), .A2(n9862), .ZN(n8309) );
  INV_X1 U5332 ( .A(n4479), .ZN(n4478) );
  OAI21_X1 U5333 ( .B1(n8567), .B2(n8566), .A(n4480), .ZN(n4479) );
  AOI21_X1 U5334 ( .B1(n8563), .B2(n8561), .A(n8571), .ZN(n4480) );
  INV_X1 U5335 ( .A(n8490), .ZN(n8781) );
  INV_X1 U5336 ( .A(n8236), .ZN(n8800) );
  INV_X1 U5337 ( .A(n7674), .ZN(n8582) );
  NAND4_X1 U5338 ( .A1(n5266), .A2(n5265), .A3(n5264), .A4(n5263), .ZN(n8586)
         );
  NAND4_X2 U5339 ( .A1(n5237), .A2(n5236), .A3(n5235), .A4(n5234), .ZN(n9838)
         );
  NAND2_X1 U5340 ( .A1(n4513), .A2(n4357), .ZN(n4512) );
  XNOR2_X1 U5341 ( .A(n8641), .B(n8642), .ZN(n8591) );
  INV_X1 U5342 ( .A(n4507), .ZN(n8619) );
  NOR2_X1 U5343 ( .A1(n4711), .A2(n4389), .ZN(n4612) );
  AOI21_X1 U5344 ( .B1(n8198), .B2(n8329), .A(n5558), .ZN(n8697) );
  NAND2_X1 U5345 ( .A1(n5537), .A2(n5536), .ZN(n8709) );
  INV_X1 U5346 ( .A(n9862), .ZN(n9843) );
  NAND2_X1 U5347 ( .A1(n4612), .A2(n4995), .ZN(n5655) );
  OR2_X1 U5348 ( .A1(n8692), .A2(n9873), .ZN(n4995) );
  NAND2_X1 U5349 ( .A1(n5465), .A2(n5464), .ZN(n8925) );
  NAND2_X1 U5350 ( .A1(n5452), .A2(n5451), .ZN(n8931) );
  NAND2_X1 U5351 ( .A1(n6145), .A2(n6144), .ZN(n9464) );
  NAND2_X1 U5352 ( .A1(n6654), .A2(n7912), .ZN(n5940) );
  NAND2_X1 U5353 ( .A1(n4463), .A2(n5810), .ZN(n6976) );
  OR2_X1 U5354 ( .A1(n6393), .A2(n5765), .ZN(n4463) );
  NAND2_X1 U5355 ( .A1(n9031), .A2(n4486), .ZN(n4485) );
  INV_X1 U5356 ( .A(n9034), .ZN(n4465) );
  INV_X1 U5357 ( .A(n9032), .ZN(n4486) );
  INV_X1 U5358 ( .A(n9039), .ZN(n4471) );
  NAND2_X1 U5359 ( .A1(n4571), .A2(n4397), .ZN(n9100) );
  AND2_X1 U5360 ( .A1(n6268), .A2(n9402), .ZN(n9119) );
  NOR2_X2 U5361 ( .A1(n6278), .A2(n6266), .ZN(n9109) );
  OR2_X1 U5362 ( .A1(n8000), .A2(n8108), .ZN(n4826) );
  INV_X1 U5363 ( .A(n4823), .ZN(n4822) );
  OAI21_X1 U5364 ( .B1(n8065), .B2(n6359), .A(n8067), .ZN(n4823) );
  NOR2_X1 U5365 ( .A1(n4392), .A2(n4454), .ZN(n4453) );
  NAND2_X1 U5366 ( .A1(n4922), .A2(n4921), .ZN(n6339) );
  AOI21_X1 U5367 ( .B1(n4359), .B2(n4877), .A(n4395), .ZN(n4921) );
  AND2_X1 U5368 ( .A1(n8086), .A2(n6371), .ZN(n8120) );
  AOI21_X1 U5369 ( .B1(n6368), .B2(n9666), .A(n6367), .ZN(n8123) );
  NAND2_X1 U5370 ( .A1(n4989), .A2(n4450), .ZN(n6367) );
  AOI21_X1 U5371 ( .B1(n4813), .B2(n7809), .A(n7926), .ZN(n4812) );
  INV_X1 U5372 ( .A(n8008), .ZN(n4813) );
  INV_X1 U5373 ( .A(n7809), .ZN(n4814) );
  OAI21_X1 U5374 ( .B1(n8396), .B2(n8395), .A(n4496), .ZN(n8398) );
  AOI21_X1 U5375 ( .B1(n7816), .B2(n4798), .A(n4797), .ZN(n4796) );
  NAND2_X1 U5376 ( .A1(n4782), .A2(n4402), .ZN(n4783) );
  NAND2_X1 U5377 ( .A1(n4787), .A2(n4785), .ZN(n7835) );
  OR2_X1 U5378 ( .A1(n8458), .A2(n8457), .ZN(n4494) );
  NOR2_X1 U5379 ( .A1(n4483), .A2(n4482), .ZN(n4481) );
  NAND2_X1 U5380 ( .A1(n7852), .A2(n7926), .ZN(n4482) );
  INV_X1 U5381 ( .A(n8039), .ZN(n4483) );
  NAND2_X1 U5382 ( .A1(n4816), .A2(n7809), .ZN(n8011) );
  INV_X1 U5383 ( .A(n7866), .ZN(n4775) );
  NAND2_X1 U5384 ( .A1(n8519), .A2(n4490), .ZN(n4489) );
  AND2_X1 U5385 ( .A1(n8518), .A2(n4491), .ZN(n4490) );
  NAND2_X1 U5386 ( .A1(n4492), .A2(n8743), .ZN(n4491) );
  INV_X1 U5387 ( .A(n7987), .ZN(n4806) );
  INV_X1 U5388 ( .A(n6350), .ZN(n7942) );
  INV_X1 U5389 ( .A(n4691), .ZN(n4690) );
  OAI21_X1 U5390 ( .B1(n5531), .B2(n4692), .A(n5552), .ZN(n4691) );
  INV_X1 U5391 ( .A(n5535), .ZN(n4692) );
  INV_X1 U5392 ( .A(n8700), .ZN(n4759) );
  OR2_X1 U5393 ( .A1(n8357), .A2(n7250), .ZN(n7149) );
  NAND2_X1 U5394 ( .A1(n4982), .A2(n5103), .ZN(n4981) );
  INV_X1 U5395 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5157) );
  AND2_X1 U5396 ( .A1(n4356), .A2(n5768), .ZN(n4572) );
  NAND2_X1 U5397 ( .A1(n6161), .A2(n9083), .ZN(n4575) );
  INV_X1 U5398 ( .A(n4709), .ZN(n4704) );
  NAND2_X1 U5399 ( .A1(n4664), .A2(n4658), .ZN(n4657) );
  INV_X1 U5400 ( .A(n5374), .ZN(n4658) );
  NOR2_X1 U5401 ( .A1(n4661), .A2(n5374), .ZN(n4660) );
  INV_X1 U5402 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4562) );
  INV_X1 U5403 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4564) );
  INV_X1 U5404 ( .A(SI_18_), .ZN(n10162) );
  INV_X1 U5405 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10158) );
  INV_X1 U5406 ( .A(SI_9_), .ZN(n10188) );
  NAND2_X1 U5407 ( .A1(n7693), .A2(n4960), .ZN(n4958) );
  NAND2_X1 U5408 ( .A1(n6760), .A2(n6618), .ZN(n4501) );
  NAND2_X1 U5409 ( .A1(n4501), .A2(n9745), .ZN(n6621) );
  NAND2_X1 U5410 ( .A1(n4937), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4936) );
  OAI21_X1 U5411 ( .B1(n6725), .B2(n4504), .A(n4502), .ZN(n6821) );
  AOI21_X1 U5412 ( .B1(n6711), .B2(n6690), .A(n4503), .ZN(n4502) );
  INV_X1 U5413 ( .A(n6712), .ZN(n4503) );
  AND2_X1 U5414 ( .A1(n9765), .A2(n4836), .ZN(n7318) );
  NAND2_X1 U5415 ( .A1(n9772), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n4836) );
  INV_X1 U5416 ( .A(n4831), .ZN(n4514) );
  NAND2_X1 U5417 ( .A1(n4516), .A2(n4831), .ZN(n4515) );
  NAND2_X1 U5418 ( .A1(n9800), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4831) );
  INV_X1 U5419 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5158) );
  AND2_X1 U5420 ( .A1(n4762), .A2(n4759), .ZN(n4758) );
  NOR2_X1 U5421 ( .A1(n8892), .A2(n8539), .ZN(n4757) );
  INV_X1 U5422 ( .A(n5245), .ZN(n4715) );
  OR2_X1 U5423 ( .A1(n8895), .A2(n8702), .ZN(n8530) );
  INV_X1 U5424 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5629) );
  NOR2_X1 U5425 ( .A1(n5365), .A2(n5156), .ZN(n5409) );
  INV_X1 U5426 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5391) );
  NAND2_X1 U5427 ( .A1(n4475), .A2(n4474), .ZN(n5365) );
  INV_X1 U5428 ( .A(n5350), .ZN(n4475) );
  INV_X1 U5429 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5154) );
  OR2_X1 U5430 ( .A1(n5296), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5311) );
  NOR2_X1 U5431 ( .A1(n8996), .A2(n4866), .ZN(n4865) );
  OAI211_X1 U5432 ( .C1(n4356), .C2(n4575), .A(n4466), .B(n4573), .ZN(n5773)
         );
  NAND2_X1 U5433 ( .A1(n8182), .A2(n4574), .ZN(n4573) );
  NAND2_X1 U5434 ( .A1(n4572), .A2(n4575), .ZN(n4466) );
  INV_X1 U5435 ( .A(n5768), .ZN(n4574) );
  AND2_X1 U5436 ( .A1(n6068), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6085) );
  NOR2_X1 U5437 ( .A1(n6048), .A2(n6047), .ZN(n6068) );
  AND2_X1 U5438 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n6280), .ZN(n6281) );
  OR2_X1 U5439 ( .A1(n6164), .A2(n8977), .ZN(n6187) );
  NOR2_X1 U5440 ( .A1(n9483), .A2(n9488), .ZN(n4602) );
  NOR2_X1 U5441 ( .A1(n5987), .A2(n5986), .ZN(n6009) );
  OR2_X1 U5442 ( .A1(n9507), .A2(n9497), .ZN(n7846) );
  INV_X1 U5443 ( .A(n7845), .ZN(n8032) );
  OR2_X1 U5444 ( .A1(n7609), .A2(n9704), .ZN(n7841) );
  INV_X1 U5445 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5964) );
  OR2_X1 U5446 ( .A1(n5965), .A2(n5964), .ZN(n5987) );
  INV_X1 U5447 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5941) );
  OR2_X1 U5448 ( .A1(n5942), .A2(n5941), .ZN(n5965) );
  AND2_X1 U5449 ( .A1(n5890), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5714) );
  NOR2_X1 U5450 ( .A1(n9670), .A2(n7292), .ZN(n4605) );
  NAND2_X1 U5451 ( .A1(n7833), .A2(n7831), .ZN(n7944) );
  AND2_X1 U5452 ( .A1(n6347), .A2(n6350), .ZN(n8019) );
  OR2_X1 U5453 ( .A1(n9660), .A2(n7241), .ZN(n7823) );
  INV_X1 U5454 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5872) );
  OR2_X1 U5455 ( .A1(n4352), .A2(n6919), .ZN(n7819) );
  AND2_X1 U5456 ( .A1(n7810), .A2(n7813), .ZN(n7938) );
  NOR2_X1 U5457 ( .A1(n7027), .A2(n9083), .ZN(n6989) );
  INV_X1 U5458 ( .A(n7022), .ZN(n4462) );
  AND2_X1 U5459 ( .A1(n9561), .A2(n6369), .ZN(n7101) );
  NAND2_X1 U5460 ( .A1(n7901), .A2(SI_29_), .ZN(n4669) );
  NAND2_X1 U5461 ( .A1(n4404), .A2(n4365), .ZN(n4996) );
  INV_X1 U5462 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5662) );
  INV_X1 U5463 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5679) );
  INV_X1 U5464 ( .A(SI_23_), .ZN(n5085) );
  AND4_X1 U5465 ( .A1(n5692), .A2(n5685), .A3(n5677), .A4(n5676), .ZN(n5678)
         );
  INV_X1 U5466 ( .A(SI_20_), .ZN(n10148) );
  AOI21_X1 U5467 ( .B1(n4678), .B2(n4366), .A(n4409), .ZN(n4677) );
  INV_X1 U5468 ( .A(n4682), .ZN(n4681) );
  AOI21_X1 U5469 ( .B1(n4680), .B2(n4682), .A(n4679), .ZN(n4678) );
  INV_X1 U5470 ( .A(n5066), .ZN(n4679) );
  INV_X1 U5471 ( .A(n4685), .ZN(n4680) );
  INV_X1 U5472 ( .A(n4665), .ZN(n4664) );
  AOI21_X1 U5473 ( .B1(n4665), .B2(n4663), .A(n4411), .ZN(n4662) );
  INV_X1 U5474 ( .A(n5048), .ZN(n4663) );
  INV_X1 U5475 ( .A(n5348), .ZN(n4666) );
  OR2_X1 U5476 ( .A1(n5909), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U5477 ( .A1(n4694), .A2(n4693), .ZN(n5336) );
  AOI21_X1 U5478 ( .B1(n4363), .B2(n4699), .A(n4412), .ZN(n4693) );
  AND2_X1 U5479 ( .A1(n5255), .A2(n5239), .ZN(n4915) );
  INV_X1 U5480 ( .A(n5022), .ZN(n4917) );
  INV_X1 U5481 ( .A(SI_26_), .ZN(n10149) );
  AOI21_X1 U5482 ( .B1(n4970), .B2(n4968), .A(n4967), .ZN(n4966) );
  INV_X1 U5483 ( .A(n4970), .ZN(n4969) );
  INV_X1 U5484 ( .A(n4972), .ZN(n4968) );
  AND2_X1 U5485 ( .A1(n8241), .A2(n8156), .ZN(n8275) );
  NOR2_X1 U5486 ( .A1(n8284), .A2(n4975), .ZN(n4970) );
  OR2_X1 U5487 ( .A1(n7691), .A2(n4958), .ZN(n7724) );
  XNOR2_X1 U5488 ( .A(n4473), .B(n9861), .ZN(n6848) );
  INV_X1 U5489 ( .A(n4958), .ZN(n4957) );
  INV_X1 U5490 ( .A(n7723), .ZN(n4955) );
  AND2_X1 U5491 ( .A1(n7757), .A2(n7756), .ZN(n7758) );
  NOR2_X1 U5492 ( .A1(n4671), .A2(n4670), .ZN(n8376) );
  NAND2_X1 U5493 ( .A1(n4674), .A2(n4672), .ZN(n4671) );
  AND2_X1 U5494 ( .A1(n8555), .A2(n8554), .ZN(n4495) );
  INV_X1 U5495 ( .A(n5200), .ZN(n5545) );
  INV_X1 U5496 ( .A(n5429), .ZN(n5598) );
  OR2_X1 U5497 ( .A1(n5601), .A2(n5233), .ZN(n5234) );
  OAI21_X1 U5498 ( .B1(n6641), .B2(n6616), .A(n6617), .ZN(n6647) );
  NAND2_X1 U5499 ( .A1(n4830), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6645) );
  INV_X1 U5500 ( .A(n6647), .ZN(n4830) );
  OR2_X1 U5501 ( .A1(n6644), .A2(n5178), .ZN(n6642) );
  XNOR2_X1 U5502 ( .A(n4353), .B(n9870), .ZN(n6762) );
  NAND2_X1 U5503 ( .A1(n6645), .A2(n6617), .ZN(n6761) );
  NAND2_X1 U5504 ( .A1(n4499), .A2(n6621), .ZN(n9741) );
  NAND2_X1 U5505 ( .A1(n4500), .A2(n4938), .ZN(n4499) );
  INV_X1 U5506 ( .A(n4501), .ZN(n4500) );
  NAND2_X1 U5507 ( .A1(n4498), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9743) );
  INV_X1 U5508 ( .A(n9741), .ZN(n4498) );
  NAND2_X1 U5509 ( .A1(n4935), .A2(n6612), .ZN(n9753) );
  INV_X1 U5510 ( .A(n4936), .ZN(n4935) );
  AND2_X1 U5511 ( .A1(n4827), .A2(n6711), .ZN(n6725) );
  NAND2_X1 U5512 ( .A1(n4829), .A2(n4828), .ZN(n4827) );
  INV_X1 U5513 ( .A(n6710), .ZN(n4829) );
  NAND2_X1 U5514 ( .A1(n6725), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U5515 ( .A1(n4506), .A2(n4934), .ZN(n4505) );
  INV_X1 U5516 ( .A(n6822), .ZN(n4506) );
  OAI21_X1 U5517 ( .B1(n7211), .B2(n7210), .A(n9766), .ZN(n9771) );
  NAND2_X1 U5518 ( .A1(n9768), .A2(n4931), .ZN(n9769) );
  AND2_X1 U5519 ( .A1(n4932), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4931) );
  AND2_X1 U5520 ( .A1(n9771), .A2(n4949), .ZN(n7322) );
  NAND2_X1 U5521 ( .A1(n9772), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4949) );
  XNOR2_X1 U5522 ( .A(n7318), .B(n7323), .ZN(n7216) );
  AND2_X1 U5523 ( .A1(n7444), .A2(n7443), .ZN(n7445) );
  NAND2_X1 U5524 ( .A1(n4927), .A2(n4457), .ZN(n4926) );
  NAND2_X1 U5525 ( .A1(n7575), .A2(n4443), .ZN(n4924) );
  AND2_X1 U5526 ( .A1(n4930), .A2(n4929), .ZN(n9792) );
  NAND2_X1 U5527 ( .A1(n4458), .A2(n4457), .ZN(n4929) );
  NAND2_X1 U5528 ( .A1(n7575), .A2(n7574), .ZN(n4458) );
  XNOR2_X1 U5529 ( .A(n8616), .B(n8642), .ZN(n8609) );
  NOR2_X1 U5530 ( .A1(n9803), .A2(n9802), .ZN(n9801) );
  INV_X1 U5531 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5166) );
  OR2_X1 U5532 ( .A1(n9801), .A2(n4508), .ZN(n4507) );
  NOR2_X1 U5533 ( .A1(n8646), .A2(n7738), .ZN(n4508) );
  NOR2_X1 U5534 ( .A1(n9823), .A2(n9824), .ZN(n9822) );
  NAND2_X1 U5535 ( .A1(n5128), .A2(n5127), .ZN(n5505) );
  NAND2_X1 U5536 ( .A1(n5126), .A2(n10060), .ZN(n5490) );
  INV_X1 U5537 ( .A(n5488), .ZN(n5126) );
  OR2_X1 U5538 ( .A1(n5476), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U5539 ( .A1(n5125), .A2(n5124), .ZN(n5466) );
  INV_X1 U5540 ( .A(n5453), .ZN(n5125) );
  INV_X1 U5541 ( .A(n5173), .ZN(n5123) );
  INV_X1 U5542 ( .A(n5426), .ZN(n5121) );
  OR2_X1 U5543 ( .A1(n5381), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5397) );
  OR2_X1 U5544 ( .A1(n5326), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U5545 ( .A1(n4633), .A2(n4631), .ZN(n7286) );
  AOI21_X1 U5546 ( .B1(n4634), .B2(n8416), .A(n4632), .ZN(n4631) );
  INV_X1 U5547 ( .A(n8425), .ZN(n4632) );
  NAND2_X1 U5548 ( .A1(n8419), .A2(n8426), .ZN(n8361) );
  OR2_X1 U5549 ( .A1(n5260), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U5550 ( .A1(n5573), .A2(n8410), .ZN(n7248) );
  NAND2_X1 U5551 ( .A1(n7248), .A2(n7250), .ZN(n7247) );
  NAND2_X1 U5552 ( .A1(n5571), .A2(n4616), .ZN(n4615) );
  NAND2_X1 U5553 ( .A1(n5571), .A2(n8399), .ZN(n7010) );
  NAND2_X1 U5554 ( .A1(n5570), .A2(n8390), .ZN(n9841) );
  NAND2_X1 U5555 ( .A1(n5569), .A2(n4951), .ZN(n6879) );
  INV_X1 U5556 ( .A(n6571), .ZN(n4951) );
  NAND2_X1 U5557 ( .A1(n5626), .A2(n6412), .ZN(n6868) );
  AND2_X1 U5558 ( .A1(n8684), .A2(n8683), .ZN(n8880) );
  NAND2_X1 U5559 ( .A1(n4766), .A2(n4761), .ZN(n4760) );
  OR2_X1 U5560 ( .A1(n4385), .A2(n4769), .ZN(n4765) );
  AND2_X1 U5561 ( .A1(n5530), .A2(n4770), .ZN(n4769) );
  INV_X1 U5562 ( .A(n4766), .ZN(n4762) );
  XNOR2_X1 U5563 ( .A(n8709), .B(n8717), .ZN(n8700) );
  AND2_X1 U5564 ( .A1(n4764), .A2(n4770), .ZN(n4763) );
  NAND2_X1 U5565 ( .A1(n4761), .A2(n5512), .ZN(n4764) );
  OAI21_X1 U5566 ( .B1(n5589), .B2(n4645), .A(n4642), .ZN(n8714) );
  AOI21_X1 U5567 ( .B1(n4644), .B2(n4643), .A(n4396), .ZN(n4642) );
  INV_X1 U5568 ( .A(n4650), .ZN(n4643) );
  INV_X1 U5569 ( .A(n4737), .ZN(n4736) );
  NAND2_X1 U5570 ( .A1(n4638), .A2(n8501), .ZN(n4637) );
  NAND2_X1 U5571 ( .A1(n4639), .A2(n8499), .ZN(n4638) );
  NAND2_X1 U5572 ( .A1(n4621), .A2(n4619), .ZN(n8812) );
  AOI21_X1 U5573 ( .B1(n4622), .B2(n4625), .A(n4620), .ZN(n4619) );
  INV_X1 U5574 ( .A(n8475), .ZN(n4620) );
  NOR2_X1 U5575 ( .A1(n8435), .A2(n8440), .ZN(n4629) );
  AND2_X1 U5576 ( .A1(n8447), .A2(n8448), .ZN(n8445) );
  NAND2_X1 U5577 ( .A1(n4717), .A2(n4720), .ZN(n7545) );
  AND2_X1 U5578 ( .A1(n4721), .A2(n5347), .ZN(n4720) );
  NAND2_X1 U5579 ( .A1(n7596), .A2(n8375), .ZN(n9913) );
  INV_X1 U5580 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4985) );
  INV_X1 U5581 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5134) );
  XNOR2_X1 U5582 ( .A(n5617), .B(P2_IR_REG_26__SCAN_IN), .ZN(n5620) );
  XNOR2_X1 U5583 ( .A(n5628), .B(n5629), .ZN(n6843) );
  INV_X1 U5584 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5092) );
  INV_X1 U5585 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5272) );
  CLKBUF_X1 U5586 ( .A(n5221), .Z(n5222) );
  INV_X1 U5587 ( .A(n6912), .ZN(n4858) );
  NAND2_X1 U5588 ( .A1(n5770), .A2(n5771), .ZN(n5775) );
  INV_X1 U5589 ( .A(n5773), .ZN(n5770) );
  NAND2_X1 U5590 ( .A1(n6904), .A2(n4585), .ZN(n4580) );
  NAND2_X1 U5591 ( .A1(n6519), .A2(n6520), .ZN(n4844) );
  NAND2_X1 U5592 ( .A1(n9057), .A2(n6126), .ZN(n8995) );
  NAND2_X1 U5593 ( .A1(n8995), .A2(n8996), .ZN(n8994) );
  INV_X1 U5594 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6047) );
  NOR2_X1 U5595 ( .A1(n4849), .A2(n4848), .ZN(n4847) );
  INV_X1 U5596 ( .A(n9108), .ZN(n4848) );
  AND2_X1 U5597 ( .A1(n6183), .A2(n6182), .ZN(n9032) );
  AOI21_X1 U5598 ( .B1(n9057), .B2(n4590), .A(n4361), .ZN(n9034) );
  AND2_X1 U5599 ( .A1(n5904), .A2(n4579), .ZN(n4578) );
  NAND2_X1 U5600 ( .A1(n6085), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U5601 ( .A1(n8994), .A2(n6143), .ZN(n8970) );
  AND2_X1 U5602 ( .A1(n6176), .A2(n6175), .ZN(n9064) );
  NAND2_X1 U5603 ( .A1(n9078), .A2(n9079), .ZN(n9077) );
  INV_X1 U5604 ( .A(n5848), .ZN(n4856) );
  OR2_X1 U5605 ( .A1(n7593), .A2(n7932), .ZN(n6274) );
  NAND2_X1 U5606 ( .A1(n5861), .A2(n5863), .ZN(n4454) );
  NAND2_X1 U5607 ( .A1(n7914), .A2(n7913), .ZN(n8087) );
  NOR2_X1 U5608 ( .A1(n8087), .A2(n8086), .ZN(n9222) );
  NOR2_X1 U5609 ( .A1(n9424), .A2(n4607), .ZN(n4606) );
  OR2_X1 U5610 ( .A1(n4610), .A2(n9281), .ZN(n4607) );
  OR2_X1 U5611 ( .A1(n8114), .A2(n9233), .ZN(n8086) );
  NAND2_X1 U5612 ( .A1(n8044), .A2(n9255), .ZN(n4876) );
  OAI21_X1 U5613 ( .B1(n4524), .B2(n4523), .A(n4871), .ZN(n9230) );
  AOI21_X1 U5614 ( .B1(n4872), .B2(n4875), .A(n9229), .ZN(n4871) );
  INV_X1 U5615 ( .A(n4872), .ZN(n4523) );
  NOR2_X1 U5616 ( .A1(n9456), .A2(n9302), .ZN(n9293) );
  OR2_X1 U5617 ( .A1(n4884), .A2(n4369), .ZN(n4525) );
  AOI21_X1 U5618 ( .B1(n4555), .B2(n4560), .A(n4553), .ZN(n4552) );
  INV_X1 U5619 ( .A(n4555), .ZN(n4554) );
  INV_X1 U5620 ( .A(n4900), .ZN(n4553) );
  NOR2_X1 U5621 ( .A1(n9328), .A2(n4599), .ZN(n4598) );
  INV_X1 U5622 ( .A(n4600), .ZN(n4599) );
  INV_X1 U5623 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8998) );
  NAND2_X1 U5624 ( .A1(n9364), .A2(n4602), .ZN(n9350) );
  NAND2_X1 U5625 ( .A1(n9364), .A2(n9370), .ZN(n9365) );
  NOR2_X1 U5626 ( .A1(n7662), .A2(n9507), .ZN(n9396) );
  AND2_X1 U5627 ( .A1(n8035), .A2(n7851), .ZN(n9409) );
  INV_X1 U5628 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6027) );
  OR2_X1 U5629 ( .A1(n6028), .A2(n6027), .ZN(n6048) );
  NAND2_X1 U5630 ( .A1(n7598), .A2(n7841), .ZN(n7659) );
  AND2_X1 U5631 ( .A1(n7846), .A2(n8032), .ZN(n7952) );
  OR2_X1 U5632 ( .A1(n7602), .A2(n7609), .ZN(n7662) );
  INV_X1 U5633 ( .A(n4540), .ZN(n4537) );
  NAND2_X1 U5634 ( .A1(n4467), .A2(n7948), .ZN(n7430) );
  AND2_X1 U5635 ( .A1(n7101), .A2(n4603), .ZN(n7438) );
  AND2_X1 U5636 ( .A1(n7413), .A2(n4368), .ZN(n4603) );
  AND2_X1 U5637 ( .A1(n7834), .A2(n4375), .ZN(n7946) );
  INV_X1 U5638 ( .A(n7946), .ZN(n7417) );
  NAND2_X1 U5639 ( .A1(n7101), .A2(n4605), .ZN(n7419) );
  NAND2_X1 U5640 ( .A1(n7101), .A2(n7100), .ZN(n7171) );
  NAND2_X1 U5641 ( .A1(n6965), .A2(n4894), .ZN(n4893) );
  NOR2_X1 U5642 ( .A1(n6350), .A2(n4895), .ZN(n4894) );
  INV_X1 U5643 ( .A(n4896), .ZN(n4895) );
  OR2_X1 U5644 ( .A1(n8019), .A2(n8017), .ZN(n4892) );
  NAND2_X1 U5645 ( .A1(n7823), .A2(n7828), .ZN(n7121) );
  NOR2_X1 U5646 ( .A1(n9563), .A2(n6310), .ZN(n9561) );
  AND2_X1 U5647 ( .A1(n6307), .A2(n6308), .ZN(n4535) );
  NAND2_X1 U5648 ( .A1(n6970), .A2(n6309), .ZN(n4536) );
  NAND2_X1 U5649 ( .A1(n6306), .A2(n7939), .ZN(n6307) );
  NAND2_X1 U5650 ( .A1(n6965), .A2(n4896), .ZN(n7060) );
  NOR2_X1 U5651 ( .A1(n7043), .A2(n6976), .ZN(n9583) );
  INV_X1 U5652 ( .A(n7939), .ZN(n7053) );
  INV_X1 U5653 ( .A(n7938), .ZN(n7040) );
  INV_X1 U5654 ( .A(n9581), .ZN(n9562) );
  NAND2_X1 U5655 ( .A1(n6300), .A2(n6299), .ZN(n6986) );
  AND2_X1 U5656 ( .A1(n7808), .A2(n8008), .ZN(n7796) );
  NAND2_X1 U5657 ( .A1(n7796), .A2(n6987), .ZN(n7035) );
  OR2_X1 U5658 ( .A1(n6220), .A2(n5776), .ZN(n5779) );
  INV_X1 U5659 ( .A(n7021), .ZN(n7934) );
  OR2_X1 U5660 ( .A1(n6743), .A2(n6742), .ZN(n6748) );
  INV_X1 U5661 ( .A(n6274), .ZN(n7995) );
  NAND2_X1 U5662 ( .A1(n5860), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4809) );
  NAND2_X1 U5663 ( .A1(n7924), .A2(n7923), .ZN(n9416) );
  NAND2_X1 U5664 ( .A1(n6215), .A2(n6214), .ZN(n9442) );
  INV_X1 U5665 ( .A(n9678), .ZN(n9708) );
  OR2_X1 U5666 ( .A1(n5784), .A2(n6385), .ZN(n4898) );
  NAND2_X1 U5667 ( .A1(n6744), .A2(n6341), .ZN(n9678) );
  AND2_X1 U5668 ( .A1(n7593), .A2(n7932), .ZN(n6744) );
  AND2_X1 U5669 ( .A1(n6249), .A2(n6250), .ZN(n6405) );
  INV_X1 U5670 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9525) );
  XNOR2_X1 U5671 ( .A(n7901), .B(n5557), .ZN(n8198) );
  INV_X1 U5672 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9526) );
  XNOR2_X1 U5673 ( .A(n5702), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6250) );
  XNOR2_X1 U5674 ( .A(n5703), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U5675 ( .A1(n4374), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U5676 ( .A1(n9527), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4867) );
  NAND2_X1 U5677 ( .A1(n4868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4870) );
  NAND2_X1 U5678 ( .A1(n5083), .A2(n5082), .ZN(n5473) );
  OR2_X1 U5679 ( .A1(n5462), .A2(n5461), .ZN(n5083) );
  XNOR2_X1 U5680 ( .A(n6265), .B(n6264), .ZN(n6398) );
  INV_X1 U5681 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6264) );
  OR2_X1 U5682 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  NOR2_X1 U5683 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5692) );
  AND2_X1 U5684 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5686) );
  AND2_X1 U5685 ( .A1(n9527), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U5686 ( .A1(n4684), .A2(n5059), .ZN(n5420) );
  NAND2_X1 U5687 ( .A1(n5057), .A2(n4685), .ZN(n4684) );
  AND2_X1 U5688 ( .A1(n6006), .A2(n5684), .ZN(n7382) );
  XNOR2_X1 U5689 ( .A(n5349), .B(n5348), .ZN(n6654) );
  NAND2_X1 U5690 ( .A1(n4695), .A2(n4696), .ZN(n5320) );
  OR2_X1 U5691 ( .A1(n5310), .A2(n4699), .ZN(n4695) );
  OAI21_X1 U5692 ( .B1(n5310), .B2(n5309), .A(n5036), .ZN(n4528) );
  XNOR2_X1 U5693 ( .A(n5008), .B(n5005), .ZN(n5189) );
  INV_X1 U5694 ( .A(SI_11_), .ZN(n10206) );
  AND2_X1 U5695 ( .A1(n5520), .A2(n5519), .ZN(n8216) );
  OAI21_X1 U5696 ( .B1(n8209), .B2(n8208), .A(n8207), .ZN(n8211) );
  NAND2_X1 U5697 ( .A1(n7724), .A2(n7723), .ZN(n7760) );
  INV_X1 U5698 ( .A(n4987), .ZN(n4986) );
  NAND2_X1 U5699 ( .A1(n8274), .A2(n8153), .ZN(n8217) );
  NAND2_X1 U5700 ( .A1(n8140), .A2(n8139), .ZN(n8225) );
  NAND2_X1 U5701 ( .A1(n4962), .A2(n4961), .ZN(n8172) );
  AOI21_X1 U5702 ( .B1(n4358), .B2(n4965), .A(n4438), .ZN(n4961) );
  AND4_X1 U5703 ( .A1(n5295), .A2(n5294), .A3(n5293), .A4(n5292), .ZN(n7614)
         );
  NAND2_X1 U5704 ( .A1(n4971), .A2(n4974), .ZN(n8283) );
  AND4_X1 U5705 ( .A1(n5433), .A2(n5432), .A3(n5431), .A4(n5430), .ZN(n8307)
         );
  AND3_X1 U5706 ( .A1(n5277), .A2(n5276), .A3(n5275), .ZN(n9900) );
  INV_X1 U5707 ( .A(n4455), .ZN(n7763) );
  OAI21_X1 U5708 ( .B1(n7691), .B2(n4956), .A(n4954), .ZN(n4455) );
  AOI21_X1 U5709 ( .B1(n7759), .B2(n4955), .A(n7758), .ZN(n4954) );
  NAND2_X1 U5710 ( .A1(n7759), .A2(n4957), .ZN(n4956) );
  INV_X1 U5711 ( .A(n8311), .ZN(n8316) );
  XNOR2_X1 U5712 ( .A(n5560), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8572) );
  NAND2_X1 U5713 ( .A1(n4383), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5560) );
  INV_X1 U5714 ( .A(n4982), .ZN(n4980) );
  INV_X1 U5715 ( .A(n8514), .ZN(n8757) );
  INV_X1 U5716 ( .A(n7614), .ZN(n8583) );
  OR2_X1 U5717 ( .A1(n5429), .A2(n5300), .ZN(n5308) );
  NAND2_X1 U5718 ( .A1(n5214), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5203) );
  OR2_X1 U5719 ( .A1(n8336), .A2(n6889), .ZN(n5181) );
  NAND2_X1 U5720 ( .A1(n4937), .A2(n6612), .ZN(n9755) );
  NAND2_X1 U5721 ( .A1(n6701), .A2(n6702), .ZN(n6834) );
  AND3_X1 U5722 ( .A1(n7213), .A2(n4505), .A3(P2_REG2_REG_7__SCAN_IN), .ZN(
        n9763) );
  NAND2_X1 U5723 ( .A1(n7213), .A2(n4505), .ZN(n6823) );
  OAI21_X1 U5724 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9765) );
  XNOR2_X1 U5725 ( .A(n7322), .B(n7323), .ZN(n7212) );
  NOR2_X1 U5726 ( .A1(n7212), .A2(n7219), .ZN(n7324) );
  NOR2_X1 U5727 ( .A1(n7450), .A2(n7504), .ZN(n7503) );
  NAND2_X1 U5728 ( .A1(n4835), .A2(n4834), .ZN(n7582) );
  INV_X1 U5729 ( .A(n7505), .ZN(n4520) );
  INV_X1 U5730 ( .A(n4833), .ZN(n9785) );
  OR2_X1 U5731 ( .A1(n8605), .A2(n8606), .ZN(n4833) );
  INV_X1 U5732 ( .A(n4943), .ZN(n8643) );
  INV_X1 U5733 ( .A(n8644), .ZN(n4942) );
  XNOR2_X1 U5734 ( .A(n4507), .B(n9834), .ZN(n9828) );
  NAND2_X1 U5735 ( .A1(n4841), .A2(n4839), .ZN(n4838) );
  AND2_X1 U5736 ( .A1(n9833), .A2(n4840), .ZN(n4839) );
  NAND2_X1 U5737 ( .A1(n9831), .A2(n9832), .ZN(n4841) );
  OR2_X1 U5738 ( .A1(n9835), .A2(n9834), .ZN(n4840) );
  AOI21_X1 U5739 ( .B1(n8681), .B2(n9832), .A(n8680), .ZN(n4476) );
  OR2_X1 U5740 ( .A1(n8679), .A2(n9825), .ZN(n4477) );
  NOR2_X1 U5741 ( .A1(n8676), .A2(n8675), .ZN(n8678) );
  AOI21_X1 U5742 ( .B1(n8957), .B2(n8329), .A(n8328), .ZN(n8687) );
  OR2_X1 U5743 ( .A1(n8692), .A2(n8691), .ZN(n4994) );
  NAND2_X1 U5744 ( .A1(n8562), .A2(n9930), .ZN(n8742) );
  NAND2_X1 U5745 ( .A1(n7548), .A2(n5362), .ZN(n7537) );
  NAND2_X1 U5746 ( .A1(n4630), .A2(n8434), .ZN(n7361) );
  NAND2_X1 U5747 ( .A1(n7269), .A2(n5334), .ZN(n7362) );
  INV_X1 U5748 ( .A(n9909), .ZN(n7315) );
  NAND2_X1 U5749 ( .A1(n4716), .A2(n5245), .ZN(n7083) );
  NAND3_X1 U5750 ( .A1(n5192), .A2(n5191), .A3(n5190), .ZN(n6886) );
  NAND2_X1 U5751 ( .A1(n5187), .A2(n4712), .ZN(n5190) );
  OR2_X1 U5752 ( .A1(n5226), .A2(n5003), .ZN(n5192) );
  INV_X1 U5753 ( .A(n8807), .ZN(n9842) );
  NAND2_X1 U5754 ( .A1(n6574), .A2(n6573), .ZN(n9862) );
  OR2_X1 U5755 ( .A1(n6874), .A2(n8742), .ZN(n8807) );
  INV_X1 U5756 ( .A(n9868), .ZN(n9871) );
  NAND2_X1 U5757 ( .A1(n8333), .A2(n8332), .ZN(n8883) );
  INV_X1 U5758 ( .A(n8709), .ZN(n8892) );
  INV_X1 U5759 ( .A(n8216), .ZN(n8895) );
  NAND2_X1 U5760 ( .A1(n5504), .A2(n5503), .ZN(n8901) );
  NAND2_X1 U5761 ( .A1(n4647), .A2(n4648), .ZN(n8724) );
  NAND2_X1 U5762 ( .A1(n5589), .A2(n4650), .ZN(n4647) );
  AOI21_X1 U5763 ( .B1(n5589), .B2(n4652), .A(n8492), .ZN(n8732) );
  NAND2_X1 U5764 ( .A1(n4739), .A2(n5483), .ZN(n8744) );
  NAND2_X1 U5765 ( .A1(n8756), .A2(n5000), .ZN(n4739) );
  AND2_X1 U5766 ( .A1(n5589), .A2(n8506), .ZN(n8751) );
  INV_X1 U5767 ( .A(n8512), .ZN(n8919) );
  OAI21_X1 U5768 ( .B1(n8788), .B2(n4731), .A(n4729), .ZN(n8765) );
  INV_X1 U5769 ( .A(n4728), .ZN(n8780) );
  NAND2_X1 U5770 ( .A1(n8802), .A2(n4640), .ZN(n8774) );
  NAND2_X1 U5771 ( .A1(n5441), .A2(n5440), .ZN(n8937) );
  NAND2_X1 U5772 ( .A1(n8802), .A2(n8484), .ZN(n8787) );
  NAND2_X1 U5773 ( .A1(n5171), .A2(n5170), .ZN(n8944) );
  NAND2_X1 U5774 ( .A1(n4618), .A2(n4622), .ZN(n8823) );
  OR2_X1 U5775 ( .A1(n7703), .A2(n4625), .ZN(n4618) );
  NAND2_X1 U5776 ( .A1(n5412), .A2(n5411), .ZN(n8260) );
  NAND2_X1 U5777 ( .A1(n4628), .A2(n8465), .ZN(n7733) );
  NAND2_X1 U5778 ( .A1(n5396), .A2(n5395), .ZN(n7761) );
  NAND2_X1 U5779 ( .A1(n5380), .A2(n5379), .ZN(n7730) );
  NAND2_X1 U5780 ( .A1(n4745), .A2(n4746), .ZN(n7632) );
  OR2_X1 U5781 ( .A1(n7548), .A2(n4749), .ZN(n4745) );
  NAND2_X1 U5782 ( .A1(n5367), .A2(n5366), .ZN(n8451) );
  INV_X1 U5783 ( .A(n8891), .ZN(n8952) );
  INV_X1 U5784 ( .A(n8947), .ZN(n8953) );
  AND2_X1 U5785 ( .A1(n5654), .A2(n5653), .ZN(n9933) );
  INV_X2 U5786 ( .A(n9933), .ZN(n9931) );
  NAND2_X1 U5787 ( .A1(n5624), .A2(n6587), .ZN(n6421) );
  INV_X1 U5788 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U5789 ( .A1(n5612), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5614) );
  INV_X1 U5790 ( .A(n8381), .ZN(n8375) );
  NAND2_X1 U5791 ( .A1(n5564), .A2(n4386), .ZN(n8566) );
  INV_X1 U5792 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7263) );
  INV_X1 U5793 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7095) );
  INV_X1 U5794 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6983) );
  INV_X1 U5795 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6861) );
  INV_X1 U5796 ( .A(n8608), .ZN(n9800) );
  INV_X1 U5797 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6565) );
  AND2_X1 U5798 ( .A1(n6398), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6379) );
  INV_X1 U5799 ( .A(n9686), .ZN(n9706) );
  NAND2_X1 U5800 ( .A1(n5934), .A2(n5933), .ZN(n7237) );
  INV_X1 U5801 ( .A(n9100), .ZN(n6246) );
  NAND2_X1 U5802 ( .A1(n4372), .A2(n4852), .ZN(n4851) );
  AND2_X1 U5803 ( .A1(n8187), .A2(n9109), .ZN(n4852) );
  NAND2_X1 U5804 ( .A1(n7923), .A2(n4595), .ZN(n4594) );
  NAND2_X1 U5805 ( .A1(n5757), .A2(n4845), .ZN(n7788) );
  NAND2_X1 U5806 ( .A1(n4844), .A2(n5756), .ZN(n7791) );
  NAND2_X1 U5807 ( .A1(n5957), .A2(n7480), .ZN(n7485) );
  NAND2_X1 U5808 ( .A1(n4588), .A2(n4587), .ZN(n9003) );
  NAND2_X1 U5809 ( .A1(n4361), .A2(n6199), .ZN(n4587) );
  AND2_X1 U5810 ( .A1(n4590), .A2(n6199), .ZN(n4589) );
  NAND2_X1 U5811 ( .A1(n9012), .A2(n9013), .ZN(n9011) );
  NAND2_X1 U5812 ( .A1(n9107), .A2(n6023), .ZN(n9012) );
  NOR2_X1 U5813 ( .A1(n6278), .A2(n6270), .ZN(n9081) );
  NAND4_X1 U5814 ( .A1(n5878), .A2(n5877), .A3(n5876), .A4(n5875), .ZN(n9658)
         );
  NAND2_X1 U5815 ( .A1(n5741), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U5816 ( .A1(n5684), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6024) );
  INV_X1 U5817 ( .A(n9416), .ZN(n9225) );
  INV_X1 U5818 ( .A(n8087), .ZN(n9419) );
  NAND2_X1 U5819 ( .A1(n9228), .A2(n4565), .ZN(n9428) );
  NAND2_X1 U5820 ( .A1(n4566), .A2(n9231), .ZN(n4565) );
  NAND2_X1 U5821 ( .A1(n4923), .A2(n4373), .ZN(n4566) );
  NAND2_X1 U5822 ( .A1(n6223), .A2(n6222), .ZN(n9447) );
  XNOR2_X1 U5823 ( .A(n4468), .B(n4877), .ZN(n9434) );
  OR2_X1 U5824 ( .A1(n9253), .A2(n6357), .ZN(n4468) );
  AND2_X1 U5825 ( .A1(n4904), .A2(n4391), .ZN(n9290) );
  NAND2_X1 U5826 ( .A1(n4904), .A2(n4903), .ZN(n9288) );
  NAND2_X1 U5827 ( .A1(n9301), .A2(n6322), .ZN(n4904) );
  NAND2_X1 U5828 ( .A1(n4881), .A2(n4882), .ZN(n9285) );
  AOI21_X1 U5829 ( .B1(n9321), .B2(n9320), .A(n6356), .ZN(n9313) );
  NAND2_X1 U5830 ( .A1(n4906), .A2(n4905), .ZN(n9319) );
  NAND2_X1 U5831 ( .A1(n4546), .A2(n4548), .ZN(n9371) );
  OR2_X1 U5832 ( .A1(n4914), .A2(n4549), .ZN(n4546) );
  NAND2_X1 U5833 ( .A1(n6067), .A2(n6066), .ZN(n9494) );
  NAND2_X1 U5834 ( .A1(n4551), .A2(n4911), .ZN(n9377) );
  OR2_X1 U5835 ( .A1(n4914), .A2(n4913), .ZN(n4551) );
  NAND2_X1 U5836 ( .A1(n5985), .A2(n5984), .ZN(n9709) );
  NAND2_X1 U5837 ( .A1(n4541), .A2(n4544), .ZN(n7434) );
  NAND2_X1 U5838 ( .A1(n4543), .A2(n4542), .ZN(n4541) );
  NAND2_X1 U5839 ( .A1(n7425), .A2(n4375), .ZN(n7350) );
  NAND2_X1 U5840 ( .A1(n6965), .A2(n7815), .ZN(n9568) );
  NOR2_X1 U5841 ( .A1(n9571), .A2(n6972), .ZN(n9586) );
  INV_X1 U5842 ( .A(n9609), .ZN(n6991) );
  NOR2_X1 U5843 ( .A1(n9571), .A2(n9712), .ZN(n9333) );
  INV_X1 U5844 ( .A(n9585), .ZN(n9331) );
  OR2_X1 U5845 ( .A1(n9571), .A2(n9703), .ZN(n9407) );
  INV_X1 U5846 ( .A(n9740), .ZN(n9737) );
  NAND2_X1 U5847 ( .A1(n8123), .A2(n4529), .ZN(n9420) );
  NAND2_X1 U5848 ( .A1(n4531), .A2(n4597), .ZN(n4530) );
  NAND2_X1 U5849 ( .A1(n4461), .A2(n4459), .ZN(n9513) );
  INV_X1 U5850 ( .A(n4460), .ZN(n4459) );
  NAND2_X1 U5851 ( .A1(n9434), .A2(n9666), .ZN(n4461) );
  OAI21_X1 U5852 ( .B1(n9436), .B2(n9663), .A(n9435), .ZN(n4460) );
  AND2_X1 U5853 ( .A1(n7720), .A2(n7775), .ZN(n6409) );
  INV_X1 U5854 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5666) );
  XNOR2_X1 U5855 ( .A(n5553), .B(n5552), .ZN(n8964) );
  NAND2_X1 U5856 ( .A1(n4689), .A2(n5535), .ZN(n5553) );
  INV_X1 U5857 ( .A(n6250), .ZN(n7775) );
  INV_X1 U5858 ( .A(n6247), .ZN(n7755) );
  NAND2_X1 U5859 ( .A1(n4707), .A2(n4706), .ZN(n5449) );
  NAND2_X1 U5860 ( .A1(n4707), .A2(n4708), .ZN(n5447) );
  INV_X1 U5861 ( .A(n8006), .ZN(n7932) );
  INV_X1 U5862 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6984) );
  INV_X1 U5863 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U5864 ( .A1(n4918), .A2(n5022), .ZN(n5254) );
  NAND2_X1 U5865 ( .A1(n4978), .A2(n6938), .ZN(n6940) );
  INV_X1 U5866 ( .A(n4512), .ZN(n7321) );
  NAND2_X1 U5867 ( .A1(n4842), .A2(n4837), .ZN(P2_U3199) );
  OAI21_X1 U5868 ( .B1(n9827), .B2(n4843), .A(n7470), .ZN(n4842) );
  NOR2_X1 U5869 ( .A1(n9830), .A2(n4838), .ZN(n4837) );
  AND2_X1 U5870 ( .A1(n9828), .A2(n8829), .ZN(n4843) );
  AOI211_X1 U5871 ( .C1(n8668), .C2(n8656), .A(n8655), .B(n8654), .ZN(n8657)
         );
  NAND2_X1 U5872 ( .A1(n5655), .A2(n9947), .ZN(n5646) );
  NOR2_X1 U5873 ( .A1(n6295), .A2(n6294), .ZN(n6296) );
  OAI21_X1 U5874 ( .B1(n8197), .B2(n4570), .A(n9109), .ZN(n6297) );
  NOR2_X1 U5875 ( .A1(n9250), .A2(n9119), .ZN(n6295) );
  AOI211_X1 U5876 ( .C1(n9464), .C2(n9084), .A(n8979), .B(n8978), .ZN(n8980)
         );
  NOR2_X1 U5877 ( .A1(n4471), .A2(n4470), .ZN(n4469) );
  NOR2_X1 U5878 ( .A1(n9297), .A2(n9119), .ZN(n4470) );
  NAND2_X1 U5879 ( .A1(n4824), .A2(n4822), .ZN(n4821) );
  OR2_X1 U5880 ( .A1(n7323), .A2(n7318), .ZN(n4357) );
  AND2_X1 U5881 ( .A1(n8166), .A2(n4963), .ZN(n4358) );
  AND2_X1 U5882 ( .A1(n9229), .A2(n4373), .ZN(n4359) );
  NAND2_X1 U5883 ( .A1(n5133), .A2(n4945), .ZN(n4360) );
  NAND2_X1 U5884 ( .A1(n4864), .A2(n4863), .ZN(n4361) );
  INV_X1 U5885 ( .A(n8158), .ZN(n8745) );
  AND2_X1 U5886 ( .A1(n5142), .A2(n5141), .ZN(n8158) );
  NAND2_X1 U5887 ( .A1(n9709), .A2(n9694), .ZN(n4362) );
  AND2_X1 U5888 ( .A1(n4696), .A2(n5319), .ZN(n4363) );
  NOR2_X1 U5889 ( .A1(n6353), .A2(n4791), .ZN(n4364) );
  INV_X1 U5890 ( .A(n6245), .ZN(n4853) );
  OR2_X1 U5891 ( .A1(n9687), .A2(n6317), .ZN(n7834) );
  INV_X1 U5892 ( .A(n9244), .ZN(n4877) );
  AND2_X1 U5893 ( .A1(n4681), .A2(n5164), .ZN(n4366) );
  AND2_X1 U5894 ( .A1(n4788), .A2(n7838), .ZN(n4367) );
  NAND2_X1 U5895 ( .A1(n6106), .A2(n6105), .ZN(n9483) );
  NAND2_X1 U5896 ( .A1(n6008), .A2(n6007), .ZN(n7609) );
  NOR2_X1 U5897 ( .A1(n9275), .A2(n4610), .ZN(n4609) );
  AND2_X1 U5898 ( .A1(n4605), .A2(n4604), .ZN(n4368) );
  AND2_X1 U5899 ( .A1(n4882), .A2(n4880), .ZN(n4369) );
  NAND2_X1 U5900 ( .A1(n4772), .A2(n8158), .ZN(n4771) );
  INV_X1 U5901 ( .A(n4771), .ZN(n4761) );
  AND2_X1 U5902 ( .A1(n4870), .A2(n4867), .ZN(n4370) );
  AND2_X1 U5903 ( .A1(n5130), .A2(n5134), .ZN(n4371) );
  AND2_X1 U5904 ( .A1(n4853), .A2(n4436), .ZN(n4372) );
  NAND2_X1 U5905 ( .A1(n7826), .A2(n7830), .ZN(n7104) );
  INV_X1 U5906 ( .A(n7104), .ZN(n4897) );
  INV_X1 U5907 ( .A(n7937), .ZN(n4799) );
  AND2_X2 U5908 ( .A1(n5717), .A2(n9534), .ZN(n5741) );
  CLKBUF_X3 U5909 ( .A(n5741), .Z(n6434) );
  NAND2_X1 U5910 ( .A1(n9250), .A2(n9438), .ZN(n4373) );
  OR2_X1 U5911 ( .A1(n5684), .A2(n4996), .ZN(n4374) );
  NAND2_X1 U5912 ( .A1(n9687), .A2(n6317), .ZN(n4375) );
  NAND4_X2 U5913 ( .A1(n5218), .A2(n5217), .A3(n5216), .A4(n5215), .ZN(n9854)
         );
  AND2_X1 U5914 ( .A1(n6273), .A2(n5722), .ZN(n5726) );
  NAND2_X1 U5915 ( .A1(n5153), .A2(n5101), .ZN(n5562) );
  INV_X1 U5916 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5133) );
  XNOR2_X1 U5917 ( .A(n9599), .B(n7792), .ZN(n6923) );
  OR2_X1 U5918 ( .A1(n7466), .A2(n7465), .ZN(n4376) );
  AND2_X1 U5919 ( .A1(n4760), .A2(n4765), .ZN(n4377) );
  INV_X1 U5920 ( .A(n8766), .ZN(n4727) );
  AND2_X1 U5921 ( .A1(n4986), .A2(n8274), .ZN(n4378) );
  AND2_X1 U5922 ( .A1(n4369), .A2(n4881), .ZN(n4379) );
  NOR2_X1 U5923 ( .A1(n8587), .A2(n7078), .ZN(n4380) );
  AND2_X1 U5924 ( .A1(n4792), .A2(n7926), .ZN(n4381) );
  OR2_X1 U5925 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4382) );
  OR2_X1 U5926 ( .A1(n5562), .A2(n4980), .ZN(n4383) );
  OR2_X1 U5927 ( .A1(n5133), .A2(n4945), .ZN(n4384) );
  NOR2_X1 U5928 ( .A1(n8216), .A2(n8702), .ZN(n4385) );
  INV_X1 U5929 ( .A(n4875), .ZN(n4874) );
  NAND2_X1 U5930 ( .A1(n4877), .A2(n4876), .ZN(n4875) );
  OR2_X1 U5931 ( .A1(n5562), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n4386) );
  INV_X1 U5932 ( .A(n8410), .ZN(n4636) );
  INV_X1 U5933 ( .A(n7274), .ZN(n4719) );
  AND3_X1 U5934 ( .A1(n8700), .A2(n8374), .A3(n8715), .ZN(n4387) );
  AND2_X1 U5935 ( .A1(n7129), .A2(n5901), .ZN(n4388) );
  INV_X1 U5936 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8959) );
  INV_X1 U5937 ( .A(n8484), .ZN(n4641) );
  AND2_X1 U5938 ( .A1(n5566), .A2(n9851), .ZN(n4389) );
  NAND2_X1 U5939 ( .A1(n5940), .A2(n5939), .ZN(n9687) );
  INV_X1 U5940 ( .A(n9687), .ZN(n4604) );
  AND2_X1 U5941 ( .A1(n8113), .A2(n9716), .ZN(n4390) );
  NAND2_X1 U5942 ( .A1(n6321), .A2(n9325), .ZN(n4391) );
  NAND2_X1 U5943 ( .A1(n5912), .A2(n5911), .ZN(n9670) );
  AND2_X1 U5944 ( .A1(n6334), .A2(n7064), .ZN(n4392) );
  INV_X1 U5945 ( .A(n9013), .ZN(n4849) );
  NAND2_X1 U5946 ( .A1(n6328), .A2(n6327), .ZN(n9424) );
  NAND2_X1 U5947 ( .A1(n6084), .A2(n6083), .ZN(n9488) );
  INV_X1 U5948 ( .A(n9328), .ZN(n9472) );
  NAND2_X1 U5949 ( .A1(n6160), .A2(n6159), .ZN(n9328) );
  AND2_X1 U5950 ( .A1(n4540), .A2(n9542), .ZN(n4393) );
  AOI21_X1 U5951 ( .B1(n8023), .B2(n8024), .A(n4791), .ZN(n4790) );
  INV_X1 U5952 ( .A(n8743), .ZN(n8913) );
  AND2_X1 U5953 ( .A1(n5487), .A2(n5486), .ZN(n8743) );
  AND2_X1 U5954 ( .A1(n4357), .A2(n7464), .ZN(n4394) );
  AND2_X1 U5955 ( .A1(n9424), .A2(n9120), .ZN(n4395) );
  INV_X1 U5956 ( .A(n4609), .ZN(n4611) );
  AND2_X1 U5957 ( .A1(n8901), .A2(n5591), .ZN(n4396) );
  INV_X1 U5958 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4945) );
  AND2_X1 U5959 ( .A1(n6232), .A2(n6231), .ZN(n4397) );
  INV_X1 U5960 ( .A(n4608), .ZN(n9257) );
  NOR2_X1 U5961 ( .A1(n9275), .A2(n9442), .ZN(n4608) );
  INV_X1 U5962 ( .A(n4560), .ZN(n4559) );
  NAND2_X1 U5963 ( .A1(n4905), .A2(n4561), .ZN(n4560) );
  NOR2_X1 U5964 ( .A1(n9320), .A2(n6356), .ZN(n4398) );
  INV_X1 U5965 ( .A(n7948), .ZN(n7433) );
  AND2_X1 U5966 ( .A1(n8028), .A2(n7836), .ZN(n7948) );
  OR2_X1 U5967 ( .A1(n6178), .A2(n6177), .ZN(n4399) );
  AND2_X1 U5968 ( .A1(n4377), .A2(n4759), .ZN(n4400) );
  AND2_X1 U5969 ( .A1(n4943), .A2(n4942), .ZN(n4401) );
  OR2_X1 U5970 ( .A1(n7292), .A2(n7478), .ZN(n7833) );
  INV_X1 U5971 ( .A(n4912), .ZN(n4911) );
  NOR2_X1 U5972 ( .A1(n9397), .A2(n9017), .ZN(n4912) );
  AND2_X1 U5973 ( .A1(n4381), .A2(n7838), .ZN(n4402) );
  OR2_X1 U5974 ( .A1(n9456), .A2(n9461), .ZN(n7969) );
  AND2_X1 U5975 ( .A1(n4596), .A2(n4594), .ZN(n4403) );
  AND3_X1 U5976 ( .A1(n5704), .A2(n5685), .A3(n6062), .ZN(n4404) );
  INV_X1 U5977 ( .A(n4960), .ZN(n4959) );
  AND2_X1 U5978 ( .A1(n6002), .A2(n6021), .ZN(n4405) );
  INV_X1 U5979 ( .A(n4975), .ZN(n4974) );
  NOR2_X1 U5980 ( .A1(n8141), .A2(n8287), .ZN(n4975) );
  INV_X2 U5981 ( .A(n5011), .ZN(n7922) );
  INV_X1 U5982 ( .A(n5512), .ZN(n4767) );
  NAND2_X1 U5983 ( .A1(n5847), .A2(n6890), .ZN(n4406) );
  NOR2_X1 U5984 ( .A1(n7730), .A2(n8578), .ZN(n4407) );
  AND2_X1 U5985 ( .A1(n9472), .A2(n9460), .ZN(n4408) );
  AND2_X1 U5986 ( .A1(n5067), .A2(SI_18_), .ZN(n4409) );
  INV_X1 U5987 ( .A(n8563), .ZN(n4674) );
  AND2_X1 U5988 ( .A1(n5024), .A2(SI_5_), .ZN(n4410) );
  AND2_X1 U5989 ( .A1(n5049), .A2(SI_13_), .ZN(n4411) );
  AND2_X1 U5990 ( .A1(n5041), .A2(SI_10_), .ZN(n4412) );
  NOR2_X1 U5991 ( .A1(n9488), .A2(n9382), .ZN(n4413) );
  INV_X1 U5992 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5677) );
  OR2_X1 U5993 ( .A1(n4984), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4414) );
  AND2_X1 U5994 ( .A1(n7073), .A2(n7085), .ZN(n4415) );
  OR2_X1 U5995 ( .A1(n5705), .A2(n4868), .ZN(n4416) );
  INV_X1 U5996 ( .A(n4645), .ZN(n4644) );
  OR2_X1 U5997 ( .A1(n4646), .A2(n8528), .ZN(n4645) );
  NOR2_X1 U5998 ( .A1(n9297), .A2(n9461), .ZN(n4417) );
  NAND2_X1 U5999 ( .A1(n4375), .A2(n7831), .ZN(n4418) );
  NAND2_X1 U6000 ( .A1(n8913), .A2(n8757), .ZN(n4419) );
  NAND2_X1 U6001 ( .A1(n7948), .A2(n8026), .ZN(n4420) );
  OR2_X1 U6002 ( .A1(n4399), .A2(n4865), .ZN(n4421) );
  NAND2_X1 U6003 ( .A1(n4920), .A2(n4544), .ZN(n4422) );
  INV_X1 U6004 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5130) );
  INV_X1 U6005 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4868) );
  OR2_X1 U6006 ( .A1(n4912), .A2(n6319), .ZN(n4423) );
  OR2_X1 U6007 ( .A1(n9602), .A2(n9125), .ZN(n6344) );
  OR2_X1 U6008 ( .A1(n8564), .A2(n8560), .ZN(n4424) );
  AND2_X1 U6009 ( .A1(n8499), .A2(n8803), .ZN(n4425) );
  INV_X1 U6010 ( .A(n9281), .ZN(n9450) );
  NAND2_X1 U6011 ( .A1(n6201), .A2(n6200), .ZN(n9281) );
  AND2_X1 U6012 ( .A1(n7820), .A2(n7819), .ZN(n4426) );
  INV_X1 U6013 ( .A(n4375), .ZN(n4791) );
  INV_X1 U6014 ( .A(n6577), .ZN(n6875) );
  INV_X1 U6015 ( .A(n6143), .ZN(n4866) );
  NAND2_X1 U6016 ( .A1(n5105), .A2(n4985), .ZN(n4984) );
  INV_X1 U6017 ( .A(n4984), .ZN(n4753) );
  AND2_X1 U6018 ( .A1(n4477), .A2(n4476), .ZN(n4427) );
  AND2_X1 U6019 ( .A1(n8131), .A2(n8129), .ZN(n4428) );
  NAND2_X1 U6020 ( .A1(n5963), .A2(n5962), .ZN(n9696) );
  AND2_X1 U6021 ( .A1(n7834), .A2(n4786), .ZN(n4429) );
  INV_X1 U6022 ( .A(n4884), .ZN(n4879) );
  NAND2_X1 U6023 ( .A1(n4885), .A2(n7969), .ZN(n4884) );
  AND2_X1 U6024 ( .A1(n4419), .A2(n4734), .ZN(n4430) );
  NAND2_X1 U6025 ( .A1(n6198), .A2(n6143), .ZN(n4431) );
  OR2_X1 U6026 ( .A1(n6313), .A2(n7114), .ZN(n4432) );
  INV_X1 U6027 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4474) );
  INV_X1 U6028 ( .A(n6334), .ZN(n6209) );
  INV_X1 U6029 ( .A(n9745), .ZN(n4938) );
  NAND2_X1 U6030 ( .A1(n5109), .A2(n5108), .ZN(n8907) );
  INV_X1 U6031 ( .A(n8907), .ZN(n4772) );
  AND2_X1 U6032 ( .A1(n9364), .A2(n4600), .ZN(n4433) );
  INV_X1 U6033 ( .A(n8508), .ZN(n8767) );
  AND2_X1 U6034 ( .A1(n5482), .A2(n5481), .ZN(n8508) );
  AND2_X1 U6035 ( .A1(n6023), .A2(n4592), .ZN(n4434) );
  NAND2_X1 U6036 ( .A1(n6128), .A2(n6127), .ZN(n9479) );
  NAND2_X1 U6037 ( .A1(n8130), .A2(n8129), .ZN(n8251) );
  NAND2_X1 U6038 ( .A1(n6135), .A2(n6134), .ZN(n9468) );
  OR2_X1 U6039 ( .A1(n7449), .A2(n7448), .ZN(n7575) );
  INV_X1 U6040 ( .A(n7575), .ZN(n4927) );
  NAND2_X1 U6041 ( .A1(n9483), .A2(n9362), .ZN(n4435) );
  NAND2_X1 U6042 ( .A1(n6235), .A2(n6234), .ZN(n4436) );
  AND2_X1 U6043 ( .A1(n4971), .A2(n4970), .ZN(n4437) );
  INV_X1 U6044 ( .A(n9362), .ZN(n9345) );
  NAND2_X1 U6045 ( .A1(n6115), .A2(n6114), .ZN(n9362) );
  INV_X1 U6046 ( .A(n9031), .ZN(n4863) );
  AND2_X1 U6047 ( .A1(n8169), .A2(n8168), .ZN(n4438) );
  INV_X1 U6048 ( .A(n7320), .ZN(n4511) );
  OR2_X1 U6049 ( .A1(n8697), .A2(n8842), .ZN(n4439) );
  NOR2_X1 U6050 ( .A1(n7691), .A2(n4959), .ZN(n4440) );
  NOR2_X1 U6051 ( .A1(n6352), .A2(n6351), .ZN(n4441) );
  AND2_X1 U6052 ( .A1(n4833), .A2(n4832), .ZN(n4442) );
  NAND2_X2 U6053 ( .A1(n6874), .A2(n9862), .ZN(n9868) );
  OR2_X1 U6054 ( .A1(n7216), .A2(n7220), .ZN(n4513) );
  OR2_X1 U6055 ( .A1(n8072), .A2(n8063), .ZN(n8070) );
  AND2_X1 U6056 ( .A1(n4536), .A2(n4535), .ZN(n7112) );
  AND2_X1 U6057 ( .A1(n7574), .A2(n8604), .ZN(n4443) );
  AND2_X1 U6058 ( .A1(n7101), .A2(n4368), .ZN(n4444) );
  AND2_X1 U6059 ( .A1(n4584), .A2(n4580), .ZN(n4445) );
  AND2_X1 U6060 ( .A1(n4893), .A2(n4892), .ZN(n4446) );
  NAND2_X1 U6061 ( .A1(n4520), .A2(n4376), .ZN(n4835) );
  AND2_X1 U6062 ( .A1(n4512), .A2(n4511), .ZN(n4447) );
  AND2_X1 U6063 ( .A1(n5556), .A2(n5555), .ZN(n4448) );
  OR2_X1 U6064 ( .A1(n5562), .A2(n4981), .ZN(n4449) );
  INV_X1 U6065 ( .A(n9855), .ZN(n8701) );
  AND2_X1 U6066 ( .A1(n6576), .A2(n8554), .ZN(n9855) );
  AND4_X2 U6067 ( .A1(n5643), .A2(n5648), .A3(n6872), .A4(n5642), .ZN(n9947)
         );
  INV_X1 U6068 ( .A(n6711), .ZN(n4504) );
  NAND2_X1 U6069 ( .A1(n6665), .A2(n8664), .ZN(n9829) );
  NAND2_X1 U6070 ( .A1(n7931), .A2(n8090), .ZN(n4450) );
  INV_X1 U6071 ( .A(n8646), .ZN(n9817) );
  AND2_X1 U6072 ( .A1(n9768), .A2(n4932), .ZN(n4451) );
  AND2_X1 U6073 ( .A1(n4976), .A2(n6938), .ZN(n4452) );
  INV_X1 U6074 ( .A(n6730), .ZN(n4828) );
  XNOR2_X1 U6075 ( .A(n5287), .B(n5286), .ZN(n7225) );
  INV_X1 U6076 ( .A(n7467), .ZN(n4834) );
  INV_X1 U6077 ( .A(n7225), .ZN(n4934) );
  NAND2_X1 U6078 ( .A1(n6835), .A2(n7225), .ZN(n9768) );
  NAND2_X1 U6079 ( .A1(n6822), .A2(n7225), .ZN(n7213) );
  INV_X1 U6080 ( .A(n8604), .ZN(n4457) );
  OR2_X1 U6081 ( .A1(n7574), .A2(n8604), .ZN(n4928) );
  NAND3_X1 U6082 ( .A1(n6023), .A2(n4592), .A3(n4847), .ZN(n4846) );
  NAND2_X2 U6083 ( .A1(n4593), .A2(n6020), .ZN(n6023) );
  NAND2_X2 U6084 ( .A1(n5862), .A2(n4453), .ZN(n9569) );
  NAND2_X1 U6085 ( .A1(n4581), .A2(n4583), .ZN(n4579) );
  NOR2_X1 U6086 ( .A1(n4585), .A2(n4583), .ZN(n4582) );
  OAI21_X1 U6087 ( .B1(n8140), .B2(n4969), .A(n4966), .ZN(n8233) );
  AOI21_X1 U6088 ( .B1(n7683), .B2(n7682), .A(n7681), .ZN(n7684) );
  AOI21_X1 U6089 ( .B1(n7201), .B2(n8586), .A(n7200), .ZN(n7203) );
  NAND2_X1 U6090 ( .A1(n6875), .A2(n4473), .ZN(n4950) );
  NAND2_X1 U6091 ( .A1(n4522), .A2(n4916), .ZN(n5267) );
  NAND2_X1 U6092 ( .A1(n8644), .A2(n4944), .ZN(n4940) );
  AOI21_X1 U6093 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n9800), .A(n9790), .ZN(
        n8641) );
  NOR2_X1 U6094 ( .A1(n9822), .A2(n8649), .ZN(n8652) );
  NAND2_X2 U6095 ( .A1(n6103), .A2(n8987), .ZN(n8985) );
  NAND2_X1 U6096 ( .A1(n6344), .A2(n4462), .ZN(n7808) );
  INV_X1 U6097 ( .A(n4855), .ZN(n4854) );
  INV_X1 U6098 ( .A(n7432), .ZN(n4467) );
  NAND2_X1 U6099 ( .A1(n7097), .A2(n7830), .ZN(n7166) );
  NAND2_X1 U6100 ( .A1(n4406), .A2(n4856), .ZN(n6913) );
  NOR2_X1 U6101 ( .A1(n9254), .A2(n9255), .ZN(n9253) );
  NOR2_X1 U6102 ( .A1(n4527), .A2(n7104), .ZN(n4526) );
  AND2_X2 U6103 ( .A1(n6003), .A2(n5678), .ZN(n5697) );
  NAND2_X1 U6104 ( .A1(n4858), .A2(n6910), .ZN(n4857) );
  NAND2_X1 U6105 ( .A1(n4464), .A2(n9109), .ZN(n4472) );
  OR2_X2 U6106 ( .A1(n6957), .A2(n5848), .ZN(n6912) );
  NAND2_X2 U6107 ( .A1(n5997), .A2(n5996), .ZN(n6002) );
  NAND2_X1 U6108 ( .A1(n9044), .A2(n5908), .ZN(n5929) );
  OAI21_X2 U6109 ( .B1(n6956), .B2(n4857), .A(n4854), .ZN(n6904) );
  INV_X1 U6110 ( .A(n4524), .ZN(n9254) );
  NOR2_X1 U6111 ( .A1(n7166), .A2(n7944), .ZN(n6352) );
  INV_X1 U6112 ( .A(n4893), .ZN(n4527) );
  NAND2_X1 U6113 ( .A1(n4878), .A2(n4525), .ZN(n9270) );
  NAND2_X1 U6114 ( .A1(n4892), .A2(n4526), .ZN(n7097) );
  INV_X1 U6115 ( .A(n4768), .ZN(n8716) );
  AOI222_X2 U6116 ( .A1(n9851), .A2(n8718), .B1(n8736), .B2(n9855), .C1(n8717), 
        .C2(n9853), .ZN(n8893) );
  NAND2_X1 U6117 ( .A1(n4472), .A2(n4469), .ZN(P1_U3229) );
  OAI21_X1 U6118 ( .B1(n6913), .B2(n5849), .A(n6911), .ZN(n4855) );
  OAI22_X1 U6119 ( .A1(n7183), .A2(n7182), .B1(n7181), .B2(n8587), .ZN(n7184)
         );
  OR2_X2 U6120 ( .A1(n7327), .A2(n7326), .ZN(n7444) );
  NOR2_X1 U6121 ( .A1(n7324), .A2(n7325), .ZN(n7327) );
  INV_X1 U6122 ( .A(n6608), .ZN(n4939) );
  NAND2_X1 U6123 ( .A1(n6834), .A2(n6833), .ZN(n6835) );
  MUX2_X1 U6124 ( .A(n8444), .B(n8443), .S(n8554), .Z(n8446) );
  INV_X1 U6125 ( .A(n4487), .ZN(n8958) );
  OAI21_X1 U6126 ( .B1(n4489), .B2(n8522), .A(n8521), .ZN(n8526) );
  OAI22_X1 U6127 ( .A1(n8417), .A2(n8416), .B1(n8554), .B2(n8415), .ZN(n8423)
         );
  NAND3_X1 U6128 ( .A1(n4424), .A2(n8565), .A3(n4478), .ZN(n8574) );
  INV_X1 U6129 ( .A(n4978), .ZN(n4977) );
  NAND2_X1 U6130 ( .A1(n8315), .A2(n8314), .ZN(n8313) );
  INV_X1 U6131 ( .A(n6939), .ZN(n4979) );
  NAND2_X1 U6132 ( .A1(n8068), .A2(n8072), .ZN(n7961) );
  NAND3_X1 U6133 ( .A1(n7930), .A2(n7929), .A3(n8069), .ZN(n8068) );
  NAND2_X1 U6134 ( .A1(n4801), .A2(n4793), .ZN(n7829) );
  NAND2_X1 U6135 ( .A1(n4819), .A2(n4818), .ZN(n7853) );
  INV_X1 U6136 ( .A(n7832), .ZN(n4781) );
  NAND2_X1 U6137 ( .A1(n4825), .A2(n6359), .ZN(n4824) );
  NAND2_X1 U6138 ( .A1(n4795), .A2(n7821), .ZN(n4794) );
  OAI211_X1 U6139 ( .C1(n7896), .C2(n7897), .A(n7895), .B(n4803), .ZN(n4802)
         );
  NAND2_X1 U6140 ( .A1(n4484), .A2(n7875), .ZN(n7877) );
  NAND2_X1 U6141 ( .A1(n4773), .A2(n7870), .ZN(n4484) );
  NAND2_X1 U6142 ( .A1(n4794), .A2(n7926), .ZN(n4793) );
  NAND2_X1 U6143 ( .A1(n5668), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5702) );
  INV_X1 U6144 ( .A(n4802), .ZN(n7898) );
  NAND2_X1 U6145 ( .A1(n7853), .A2(n4817), .ZN(n7850) );
  NAND2_X1 U6146 ( .A1(n4821), .A2(n8085), .ZN(P1_U3242) );
  OAI21_X1 U6147 ( .B1(n4796), .B2(n7817), .A(n4426), .ZN(n4795) );
  NAND2_X1 U6148 ( .A1(n7827), .A2(n4429), .ZN(n4782) );
  NAND2_X1 U6149 ( .A1(n4811), .A2(n4815), .ZN(n7812) );
  OAI21_X1 U6150 ( .B1(n7894), .B2(n7893), .A(n4804), .ZN(n4803) );
  OAI21_X1 U6151 ( .B1(n8001), .B2(n8063), .A(n4826), .ZN(n4825) );
  AOI21_X1 U6152 ( .B1(n7849), .B2(n7926), .A(n4820), .ZN(n4819) );
  OAI211_X1 U6153 ( .C1(n6023), .C2(n4849), .A(n4846), .B(n6043), .ZN(n9024)
         );
  NAND3_X4 U6154 ( .A1(n5701), .A2(n6340), .A3(n6273), .ZN(n8182) );
  MUX2_X1 U6155 ( .A(n8482), .B(n8481), .S(n8545), .Z(n8498) );
  NAND2_X1 U6156 ( .A1(n4493), .A2(n8459), .ZN(n8464) );
  NAND2_X1 U6157 ( .A1(n8456), .A2(n4494), .ZN(n4493) );
  NAND3_X1 U6158 ( .A1(n8556), .A2(n8553), .A3(n4495), .ZN(n8557) );
  INV_X1 U6159 ( .A(n4513), .ZN(n7319) );
  OAI22_X1 U6160 ( .A1(n8605), .A2(n4515), .B1(n4832), .B2(n4514), .ZN(n8616)
         );
  NAND2_X1 U6161 ( .A1(n5267), .A2(n5268), .ZN(n4521) );
  NAND2_X1 U6162 ( .A1(n4915), .A2(n5238), .ZN(n4522) );
  OR2_X2 U6163 ( .A1(n9270), .A2(n7979), .ZN(n4524) );
  XNOR2_X2 U6164 ( .A(n4528), .B(n4997), .ZN(n6514) );
  MUX2_X1 U6165 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7917), .Z(n5024) );
  NAND3_X1 U6166 ( .A1(n4654), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4532) );
  NAND3_X1 U6167 ( .A1(n4564), .A2(n4563), .A3(n4562), .ZN(n4533) );
  NAND3_X1 U6168 ( .A1(n4534), .A2(n4432), .A3(n6315), .ZN(n7105) );
  OAI21_X1 U6169 ( .B1(n7352), .B2(n4537), .A(n4539), .ZN(n7597) );
  INV_X1 U6170 ( .A(n7352), .ZN(n4543) );
  NAND2_X1 U6171 ( .A1(n4545), .A2(n4547), .ZN(n6320) );
  NAND2_X1 U6172 ( .A1(n4914), .A2(n4548), .ZN(n4545) );
  XNOR2_X1 U6173 ( .A(n5254), .B(n5255), .ZN(n6393) );
  INV_X1 U6174 ( .A(n5775), .ZN(n4569) );
  NAND2_X1 U6175 ( .A1(n4568), .A2(n5775), .ZN(n4567) );
  INV_X1 U6176 ( .A(n9078), .ZN(n4568) );
  NAND2_X1 U6177 ( .A1(n9077), .A2(n5775), .ZN(n6790) );
  AND2_X1 U6178 ( .A1(n5774), .A2(n5775), .ZN(n9079) );
  INV_X1 U6179 ( .A(n9004), .ZN(n4571) );
  NAND2_X1 U6180 ( .A1(n8986), .A2(n8989), .ZN(n6103) );
  NAND2_X2 U6181 ( .A1(n9088), .A2(n9089), .ZN(n8986) );
  AND2_X2 U6182 ( .A1(n4576), .A2(n8989), .ZN(n9088) );
  NAND2_X1 U6183 ( .A1(n6079), .A2(n6078), .ZN(n8989) );
  OR2_X2 U6184 ( .A1(n6079), .A2(n6078), .ZN(n4576) );
  NAND2_X1 U6185 ( .A1(n4577), .A2(n4578), .ZN(n9044) );
  NAND2_X1 U6186 ( .A1(n6904), .A2(n4581), .ZN(n4577) );
  NAND2_X2 U6187 ( .A1(n6213), .A2(n8182), .ZN(n6161) );
  NAND3_X1 U6188 ( .A1(n4586), .A2(n6273), .A3(n6971), .ZN(n6213) );
  NAND2_X1 U6189 ( .A1(n9057), .A2(n4589), .ZN(n4588) );
  NAND4_X1 U6190 ( .A1(n5659), .A2(n5763), .A3(n5799), .A4(n5660), .ZN(n5671)
         );
  INV_X1 U6191 ( .A(n5671), .ZN(n4891) );
  NAND3_X1 U6192 ( .A1(n5659), .A2(n5763), .A3(n5799), .ZN(n5823) );
  NAND2_X1 U6193 ( .A1(n4405), .A2(n7777), .ZN(n4592) );
  XNOR2_X2 U6194 ( .A(n5670), .B(P1_IR_REG_27__SCAN_IN), .ZN(n8095) );
  XNOR2_X2 U6195 ( .A(n5712), .B(n9526), .ZN(n6269) );
  NAND2_X1 U6196 ( .A1(n9364), .A2(n4598), .ZN(n9322) );
  NAND2_X1 U6197 ( .A1(n9293), .A2(n4606), .ZN(n9233) );
  NAND2_X1 U6198 ( .A1(n9293), .A2(n9450), .ZN(n9275) );
  NAND2_X1 U6199 ( .A1(n4612), .A2(n4994), .ZN(n8693) );
  OAI21_X1 U6200 ( .B1(n8397), .B2(n4617), .A(n8358), .ZN(n4613) );
  INV_X1 U6201 ( .A(n4613), .ZN(n4614) );
  NAND2_X1 U6202 ( .A1(n4615), .A2(n4614), .ZN(n7086) );
  NAND2_X1 U6203 ( .A1(n7010), .A2(n8397), .ZN(n7088) );
  NAND2_X1 U6204 ( .A1(n7703), .A2(n4622), .ZN(n4621) );
  NAND2_X1 U6205 ( .A1(n7703), .A2(n8466), .ZN(n4628) );
  INV_X1 U6206 ( .A(n4626), .ZN(n4625) );
  NAND2_X1 U6207 ( .A1(n4630), .A2(n4629), .ZN(n5576) );
  NAND2_X1 U6208 ( .A1(n5573), .A2(n4634), .ZN(n4633) );
  OR2_X2 U6209 ( .A1(n5562), .A2(n4754), .ZN(n5616) );
  AOI21_X1 U6210 ( .B1(n8804), .B2(n4425), .A(n4637), .ZN(n8763) );
  NAND2_X1 U6211 ( .A1(n5485), .A2(n5484), .ZN(n5091) );
  NAND2_X1 U6212 ( .A1(n5473), .A2(n5472), .ZN(n4653) );
  NAND2_X1 U6213 ( .A1(n5349), .A2(n4660), .ZN(n4659) );
  OAI21_X1 U6214 ( .B1(n5349), .B2(n4666), .A(n5048), .ZN(n5364) );
  NAND2_X1 U6215 ( .A1(n7916), .A2(n7915), .ZN(n7921) );
  NAND2_X1 U6216 ( .A1(n5057), .A2(n4676), .ZN(n4675) );
  NAND2_X1 U6217 ( .A1(n4675), .A2(n4677), .ZN(n5152) );
  NAND2_X1 U6218 ( .A1(n5532), .A2(n4690), .ZN(n4688) );
  NAND2_X1 U6219 ( .A1(n5532), .A2(n5531), .ZN(n4689) );
  NAND2_X1 U6220 ( .A1(n5310), .A2(n4363), .ZN(n4694) );
  OAI21_X1 U6221 ( .B1(n5439), .B2(n4705), .A(n4702), .ZN(n5462) );
  NAND2_X1 U6222 ( .A1(n5607), .A2(n5606), .ZN(n4711) );
  INV_X2 U6223 ( .A(n7917), .ZN(n4713) );
  NAND2_X2 U6224 ( .A1(n5596), .A2(n5595), .ZN(n5187) );
  NAND2_X1 U6225 ( .A1(n4716), .A2(n4714), .ZN(n5259) );
  NOR2_X1 U6226 ( .A1(n4380), .A2(n4715), .ZN(n4714) );
  NAND2_X1 U6227 ( .A1(n5333), .A2(n4718), .ZN(n4717) );
  OAI21_X1 U6228 ( .B1(n8756), .B2(n4736), .A(n4430), .ZN(n4740) );
  INV_X1 U6229 ( .A(n4740), .ZN(n8735) );
  NAND2_X1 U6230 ( .A1(n7548), .A2(n4743), .ZN(n4742) );
  INV_X1 U6231 ( .A(n4981), .ZN(n4750) );
  AND2_X1 U6232 ( .A1(n5101), .A2(n4753), .ZN(n4752) );
  INV_X1 U6233 ( .A(n4754), .ZN(n4751) );
  OAI21_X1 U6234 ( .B1(n8733), .B2(n4762), .A(n4377), .ZN(n8699) );
  NAND2_X1 U6235 ( .A1(n4755), .A2(n4756), .ZN(n5559) );
  NAND2_X1 U6236 ( .A1(n8733), .A2(n4771), .ZN(n8726) );
  OAI21_X1 U6237 ( .B1(n8733), .B2(n4767), .A(n4763), .ZN(n4768) );
  NAND2_X1 U6238 ( .A1(n5259), .A2(n5258), .ZN(n7191) );
  NAND2_X1 U6239 ( .A1(n4774), .A2(n9320), .ZN(n4773) );
  NAND2_X1 U6240 ( .A1(n4776), .A2(n4775), .ZN(n4774) );
  NAND2_X1 U6241 ( .A1(n4778), .A2(n4777), .ZN(n4776) );
  OAI211_X1 U6242 ( .C1(n7857), .C2(n7926), .A(n4779), .B(n7862), .ZN(n4778)
         );
  AOI21_X1 U6243 ( .B1(n4780), .B2(n4367), .A(n4420), .ZN(n4784) );
  AND2_X1 U6244 ( .A1(n7833), .A2(n7826), .ZN(n4786) );
  NAND2_X1 U6245 ( .A1(n5758), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n4807) );
  AND2_X1 U6246 ( .A1(n8199), .A2(n9534), .ZN(n5758) );
  NAND2_X1 U6247 ( .A1(n5741), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4808) );
  NOR2_X2 U6248 ( .A1(n5717), .A2(n9534), .ZN(n5860) );
  NAND2_X1 U6249 ( .A1(n5740), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4810) );
  NOR2_X2 U6250 ( .A1(n8199), .A2(n9534), .ZN(n5740) );
  NAND2_X2 U6251 ( .A1(n5730), .A2(n4403), .ZN(n7792) );
  OAI21_X1 U6252 ( .B1(n7808), .B2(n4814), .A(n4812), .ZN(n4811) );
  NAND2_X1 U6253 ( .A1(n5667), .A2(n4990), .ZN(n5709) );
  INV_X1 U6254 ( .A(n5709), .ZN(n9531) );
  NAND2_X1 U6255 ( .A1(n6821), .A2(n6820), .ZN(n6822) );
  NAND2_X2 U6256 ( .A1(n5185), .A2(n5186), .ZN(n6641) );
  NAND4_X1 U6257 ( .A1(n4845), .A2(n4844), .A3(n5756), .A4(n5757), .ZN(n7789)
         );
  NAND2_X1 U6258 ( .A1(n5739), .A2(n5738), .ZN(n5757) );
  NAND2_X1 U6259 ( .A1(n5737), .A2(n5736), .ZN(n4845) );
  NAND2_X1 U6260 ( .A1(n5998), .A2(n6002), .ZN(n7776) );
  NAND2_X2 U6261 ( .A1(n4850), .A2(n5998), .ZN(n7777) );
  AND2_X2 U6262 ( .A1(n6002), .A2(n6001), .ZN(n4850) );
  OR2_X1 U6263 ( .A1(n6246), .A2(n4851), .ZN(n8195) );
  NAND3_X1 U6264 ( .A1(n7296), .A2(n7297), .A3(n7482), .ZN(n5957) );
  INV_X1 U6265 ( .A(n5933), .ZN(n7294) );
  NAND3_X1 U6266 ( .A1(n5934), .A2(n5933), .A3(n4993), .ZN(n7297) );
  NOR2_X2 U6267 ( .A1(n5854), .A2(n5661), .ZN(n6003) );
  NOR2_X2 U6268 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4859) );
  NOR2_X2 U6269 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4860) );
  NOR2_X2 U6270 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4861) );
  NAND2_X1 U6271 ( .A1(n5697), .A2(n4869), .ZN(n5706) );
  OAI21_X1 U6272 ( .B1(n9254), .B2(n4875), .A(n4872), .ZN(n9232) );
  NAND3_X1 U6273 ( .A1(n9321), .A2(n4883), .A3(n4879), .ZN(n4878) );
  NAND2_X1 U6274 ( .A1(n6352), .A2(n4364), .ZN(n4886) );
  NOR2_X2 U6275 ( .A1(n5661), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n4890) );
  INV_X1 U6276 ( .A(n4996), .ZN(n4889) );
  NAND4_X1 U6277 ( .A1(n4890), .A2(n5664), .A3(n4889), .A4(n4891), .ZN(n5668)
         );
  NAND2_X1 U6278 ( .A1(n5238), .A2(n5239), .ZN(n4918) );
  NAND2_X1 U6279 ( .A1(n9243), .A2(n4359), .ZN(n4922) );
  NAND2_X1 U6280 ( .A1(n4923), .A2(n4359), .ZN(n9228) );
  NAND3_X1 U6281 ( .A1(n4926), .A2(n4928), .A3(n4924), .ZN(n7577) );
  NAND3_X1 U6282 ( .A1(n4926), .A2(n4925), .A3(n4924), .ZN(n4930) );
  INV_X1 U6283 ( .A(n4930), .ZN(n8588) );
  NAND2_X1 U6284 ( .A1(n6834), .A2(n4933), .ZN(n4932) );
  NAND2_X1 U6285 ( .A1(n4936), .A2(n6612), .ZN(n6610) );
  NAND2_X1 U6286 ( .A1(n4939), .A2(n4938), .ZN(n4937) );
  NAND2_X1 U6287 ( .A1(n6608), .A2(n9745), .ZN(n6612) );
  AND2_X1 U6288 ( .A1(n6571), .A2(n4950), .ZN(n6799) );
  NOR2_X1 U6289 ( .A1(n5096), .A2(n5222), .ZN(n5321) );
  AND2_X2 U6290 ( .A1(n4953), .A2(n4952), .ZN(n5153) );
  INV_X1 U6291 ( .A(n5096), .ZN(n4953) );
  NAND2_X1 U6292 ( .A1(n8130), .A2(n4428), .ZN(n8252) );
  NAND2_X1 U6293 ( .A1(n7692), .A2(n8580), .ZN(n4960) );
  NAND2_X1 U6294 ( .A1(n8244), .A2(n8163), .ZN(n8315) );
  OAI21_X1 U6295 ( .B1(n8244), .B2(n4965), .A(n4358), .ZN(n8210) );
  NAND2_X1 U6296 ( .A1(n8244), .A2(n4358), .ZN(n4962) );
  NAND2_X1 U6297 ( .A1(n8274), .A2(n4987), .ZN(n8157) );
  NAND2_X1 U6298 ( .A1(n5693), .A2(n5692), .ZN(n5694) );
  OAI21_X1 U6299 ( .B1(n5199), .B2(n5007), .A(n5748), .ZN(n5188) );
  OAI21_X1 U6300 ( .B1(n9277), .B2(n6209), .A(n6208), .ZN(n9262) );
  OR2_X1 U6301 ( .A1(n9324), .A2(n6209), .ZN(n6169) );
  OR2_X1 U6302 ( .A1(n9339), .A2(n6209), .ZN(n6135) );
  INV_X1 U6303 ( .A(n5716), .ZN(n5717) );
  AND2_X1 U6304 ( .A1(n4713), .A2(P2_U3151), .ZN(n6683) );
  OR2_X1 U6305 ( .A1(n6312), .A2(n7817), .ZN(n9550) );
  NAND4_X2 U6306 ( .A1(n5182), .A2(n5181), .A3(n5180), .A4(n5179), .ZN(n6675)
         );
  OR2_X1 U6307 ( .A1(n5200), .A2(n6667), .ZN(n5195) );
  NAND2_X1 U6308 ( .A1(n9378), .A2(n7854), .ZN(n9360) );
  NAND2_X1 U6309 ( .A1(n9872), .A2(n6675), .ZN(n8387) );
  NAND2_X2 U6310 ( .A1(n6727), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6726) );
  INV_X2 U6311 ( .A(n5765), .ZN(n7912) );
  NAND4_X2 U6312 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n9125)
         );
  NAND4_X4 U6313 ( .A1(n5798), .A2(n5797), .A3(n5796), .A4(n5795), .ZN(n9124)
         );
  OR2_X2 U6314 ( .A1(n6209), .A2(n6958), .ZN(n5798) );
  OAI21_X1 U6315 ( .B1(n8714), .B2(n8713), .A(n8530), .ZN(n8698) );
  OR2_X1 U6316 ( .A1(n7761), .A2(n8577), .ZN(n4988) );
  XNOR2_X1 U6317 ( .A(n5614), .B(n5613), .ZN(n5625) );
  XNOR2_X1 U6318 ( .A(n5611), .B(n5610), .ZN(n5619) );
  OAI22_X1 U6319 ( .A1(n6800), .A2(n6799), .B1(n6798), .B2(n6675), .ZN(n6852)
         );
  NAND2_X1 U6320 ( .A1(n9120), .A2(n9659), .ZN(n4989) );
  AND2_X1 U6321 ( .A1(n5666), .A2(n5665), .ZN(n4990) );
  OR2_X1 U6322 ( .A1(n9450), .A2(n9439), .ZN(n4991) );
  AND2_X1 U6323 ( .A1(n7368), .A2(n7367), .ZN(n4992) );
  INV_X1 U6324 ( .A(n5458), .ZN(n8793) );
  AND3_X1 U6325 ( .A1(n5457), .A2(n5456), .A3(n5455), .ZN(n5458) );
  INV_X1 U6326 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5124) );
  INV_X1 U6327 ( .A(n8702), .ZN(n8168) );
  AND2_X1 U6328 ( .A1(n5040), .A2(n5039), .ZN(n4997) );
  INV_X1 U6329 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5120) );
  INV_X1 U6330 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5114) );
  INV_X1 U6331 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9527) );
  AND2_X1 U6332 ( .A1(n4713), .A2(P1_U3086), .ZN(n7628) );
  INV_X1 U6333 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5117) );
  INV_X1 U6334 ( .A(n8269), .ZN(n8826) );
  AND4_X1 U6335 ( .A1(n5418), .A2(n5417), .A3(n5416), .A4(n5415), .ZN(n8269)
         );
  INV_X1 U6336 ( .A(n8931), .ZN(n5459) );
  INV_X1 U6337 ( .A(n5726), .ZN(n5734) );
  NAND2_X1 U6338 ( .A1(n6748), .A2(n9402), .ZN(n9393) );
  AND2_X2 U6339 ( .A1(n6561), .A2(n6375), .ZN(n9719) );
  OR2_X1 U6340 ( .A1(n8697), .A2(n8891), .ZN(n4999) );
  INV_X1 U6341 ( .A(n8974), .ZN(n6178) );
  OR2_X1 U6342 ( .A1(n8512), .A2(n8508), .ZN(n5000) );
  AND2_X1 U6343 ( .A1(n8743), .A2(n8514), .ZN(n5001) );
  INV_X1 U6344 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5098) );
  INV_X1 U6345 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5103) );
  OR2_X1 U6346 ( .A1(n5624), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5621) );
  NAND2_X1 U6347 ( .A1(n8512), .A2(n8508), .ZN(n5483) );
  INV_X1 U6348 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5061) );
  AND2_X1 U6349 ( .A1(n8944), .A2(n8827), .ZN(n5434) );
  INV_X1 U6350 ( .A(n5354), .ZN(n5116) );
  OR2_X1 U6351 ( .A1(n8925), .A2(n8781), .ZN(n5471) );
  INV_X1 U6352 ( .A(n8361), .ZN(n5574) );
  NAND2_X1 U6353 ( .A1(n4449), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5628) );
  NOR2_X1 U6354 ( .A1(n8973), .A2(n9064), .ZN(n6177) );
  INV_X1 U6355 ( .A(n5734), .ZN(n6174) );
  AOI21_X1 U6356 ( .B1(n9599), .B2(n8179), .A(n5735), .ZN(n5738) );
  AND3_X1 U6357 ( .A1(n8069), .A2(n7960), .A3(n8071), .ZN(n7997) );
  INV_X1 U6358 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5986) );
  INV_X1 U6359 ( .A(n9424), .ZN(n6370) );
  NOR2_X1 U6360 ( .A1(n6129), .A2(n8998), .ZN(n6146) );
  INV_X1 U6361 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5685) );
  INV_X1 U6362 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5660) );
  INV_X1 U6363 ( .A(SI_30_), .ZN(n10146) );
  INV_X1 U6364 ( .A(SI_14_), .ZN(n10050) );
  INV_X1 U6365 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10040) );
  INV_X1 U6366 ( .A(n8579), .ZN(n7722) );
  INV_X1 U6367 ( .A(n8167), .ZN(n8169) );
  OR2_X1 U6368 ( .A1(n8128), .A2(n8258), .ZN(n8129) );
  INV_X1 U6369 ( .A(n8306), .ZN(n8319) );
  INV_X1 U6370 ( .A(n8206), .ZN(n5136) );
  INV_X1 U6371 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U6372 ( .A1(n5121), .A2(n5120), .ZN(n5428) );
  OR2_X1 U6373 ( .A1(n5340), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5354) );
  OR2_X1 U6374 ( .A1(n5301), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6375 ( .A1(n5187), .A2(n4713), .ZN(n5226) );
  AND2_X1 U6376 ( .A1(n8937), .A2(n8236), .ZN(n8485) );
  INV_X1 U6377 ( .A(n8445), .ZN(n5360) );
  AND2_X1 U6378 ( .A1(n7189), .A2(n8408), .ZN(n8358) );
  AND2_X1 U6379 ( .A1(n5594), .A2(n6863), .ZN(n6656) );
  NAND2_X2 U6380 ( .A1(n7923), .A2(n7917), .ZN(n5784) );
  OR2_X1 U6381 ( .A1(n6187), .A2(n9037), .ZN(n6203) );
  OR2_X1 U6382 ( .A1(n6108), .A2(n6107), .ZN(n6129) );
  NAND2_X1 U6383 ( .A1(n6896), .A2(n9577), .ZN(n7937) );
  INV_X1 U6384 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6252) );
  INV_X1 U6385 ( .A(SI_27_), .ZN(n10166) );
  INV_X1 U6386 ( .A(SI_24_), .ZN(n10058) );
  AND2_X1 U6387 ( .A1(n5687), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5688) );
  INV_X1 U6388 ( .A(SI_15_), .ZN(n10118) );
  INV_X1 U6389 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6390 ( .A1(n7721), .A2(n7722), .ZN(n7723) );
  NAND2_X1 U6391 ( .A1(n5123), .A2(n5122), .ZN(n5442) );
  INV_X1 U6392 ( .A(n8581), .ZN(n7675) );
  OR3_X1 U6393 ( .A1(n5649), .A2(n8381), .A3(n8566), .ZN(n6578) );
  OR3_X1 U6394 ( .A1(n6677), .A2(n6576), .A3(n6863), .ZN(n8321) );
  OR2_X1 U6395 ( .A1(n5538), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8685) );
  OR2_X1 U6396 ( .A1(n5466), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5476) );
  OR2_X1 U6397 ( .A1(n5428), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5173) );
  OR2_X1 U6398 ( .A1(n9838), .A2(n9889), .ZN(n8405) );
  INV_X1 U6399 ( .A(n6867), .ZN(n6866) );
  INV_X1 U6400 ( .A(n8368), .ZN(n8468) );
  INV_X1 U6401 ( .A(n8366), .ZN(n8459) );
  XNOR2_X1 U6402 ( .A(n5820), .B(n4356), .ZN(n6892) );
  INV_X1 U6403 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9037) );
  INV_X1 U6404 ( .A(n9694), .ZN(n7408) );
  INV_X1 U6405 ( .A(n9102), .ZN(n9113) );
  AND2_X1 U6406 ( .A1(n8115), .A2(n6284), .ZN(n9235) );
  NOR2_X1 U6407 ( .A1(n6203), .A2(n6202), .ZN(n6216) );
  INV_X1 U6408 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6509) );
  INV_X1 U6409 ( .A(n9446), .ZN(n9461) );
  INV_X1 U6410 ( .A(n9304), .ZN(n9460) );
  INV_X1 U6411 ( .A(n9364), .ZN(n9385) );
  INV_X1 U6412 ( .A(n9539), .ZN(n9497) );
  INV_X1 U6413 ( .A(n9121), .ZN(n9704) );
  INV_X1 U6414 ( .A(n9578), .ZN(n9369) );
  AND2_X1 U6415 ( .A1(n7838), .A2(n8026), .ZN(n7947) );
  INV_X1 U6416 ( .A(n8074), .ZN(n6360) );
  OR2_X1 U6417 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  INV_X1 U6418 ( .A(n8321), .ZN(n8303) );
  NAND2_X1 U6419 ( .A1(n8231), .A2(n8147), .ZN(n8294) );
  NAND2_X1 U6420 ( .A1(n6847), .A2(n6846), .ZN(n8323) );
  AND2_X1 U6421 ( .A1(n5529), .A2(n5528), .ZN(n8702) );
  AND3_X1 U6422 ( .A1(n5470), .A2(n5469), .A3(n5468), .ZN(n8490) );
  AND4_X1 U6423 ( .A1(n5359), .A2(n5358), .A3(n5357), .A4(n5356), .ZN(n7673)
         );
  INV_X1 U6424 ( .A(n9783), .ZN(n9818) );
  AND2_X1 U6425 ( .A1(P2_U3893), .A2(n5595), .ZN(n9832) );
  INV_X1 U6426 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7579) );
  AND2_X1 U6427 ( .A1(n5572), .A2(n8410), .ZN(n8357) );
  INV_X1 U6428 ( .A(n8833), .ZN(n9845) );
  INV_X1 U6429 ( .A(n8842), .ZN(n8875) );
  AND2_X1 U6430 ( .A1(n9947), .A2(n9919), .ZN(n8876) );
  OR2_X1 U6431 ( .A1(n5622), .A2(n6868), .ZN(n5648) );
  OR2_X1 U6432 ( .A1(n8476), .A2(n8353), .ZN(n8814) );
  INV_X1 U6433 ( .A(n9913), .ZN(n9930) );
  NAND2_X1 U6434 ( .A1(n7013), .A2(n9873), .ZN(n9919) );
  OR2_X1 U6435 ( .A1(n6677), .A2(n6581), .ZN(n5653) );
  INV_X1 U6436 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5240) );
  INV_X1 U6437 ( .A(n9112), .ZN(n9058) );
  OR2_X1 U6438 ( .A1(n6406), .A2(n6373), .ZN(n9402) );
  OR2_X1 U6439 ( .A1(n6204), .A2(n6216), .ZN(n9277) );
  NAND2_X1 U6440 ( .A1(n6169), .A2(n6168), .ZN(n9304) );
  INV_X1 U6441 ( .A(n7530), .ZN(n9204) );
  OR2_X1 U6442 ( .A1(n6476), .A2(n6475), .ZN(n7530) );
  INV_X1 U6443 ( .A(n9165), .ZN(n9211) );
  AND2_X1 U6444 ( .A1(n6744), .A2(n8064), .ZN(n9581) );
  OAI22_X1 U6445 ( .A1(n7657), .A2(n7952), .B1(n9022), .B2(n9497), .ZN(n9395)
         );
  AOI21_X1 U6446 ( .B1(n6405), .B2(n6251), .A(n6409), .ZN(n6742) );
  INV_X1 U6447 ( .A(n9666), .ZN(n9712) );
  INV_X1 U6448 ( .A(n9716), .ZN(n9663) );
  NAND2_X1 U6449 ( .A1(n9647), .A2(n9654), .ZN(n9716) );
  NOR2_X1 U6450 ( .A1(n6741), .A2(n6374), .ZN(n6561) );
  NAND2_X1 U6451 ( .A1(n6843), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6380) );
  AND2_X1 U6452 ( .A1(n6570), .A2(n6569), .ZN(n8311) );
  NAND2_X1 U6453 ( .A1(n5544), .A2(n5543), .ZN(n8717) );
  OR2_X1 U6454 ( .A1(P2_U3150), .A2(n6631), .ZN(n9783) );
  NAND2_X1 U6455 ( .A1(n6665), .A2(n8631), .ZN(n9825) );
  AND2_X1 U6456 ( .A1(n6633), .A2(n6632), .ZN(n9835) );
  AND2_X1 U6457 ( .A1(n7158), .A2(n7157), .ZN(n9912) );
  NAND2_X1 U6458 ( .A1(n9868), .A2(n9860), .ZN(n8833) );
  AND2_X1 U6459 ( .A1(n4439), .A2(n5644), .ZN(n5645) );
  INV_X1 U6460 ( .A(n8876), .ZN(n8874) );
  INV_X1 U6461 ( .A(n9947), .ZN(n9945) );
  AND2_X1 U6462 ( .A1(n4999), .A2(n5656), .ZN(n5657) );
  OR2_X1 U6463 ( .A1(n9933), .A2(n9925), .ZN(n8947) );
  AND3_X1 U6464 ( .A1(n9924), .A2(n9923), .A3(n9922), .ZN(n9944) );
  AND3_X1 U6465 ( .A1(n9881), .A2(n9880), .A3(n9879), .ZN(n9935) );
  INV_X1 U6466 ( .A(n6380), .ZN(n6587) );
  INV_X1 U6467 ( .A(n5620), .ZN(n7772) );
  INV_X1 U6468 ( .A(n8668), .ZN(n8650) );
  INV_X1 U6469 ( .A(n7214), .ZN(n9772) );
  AND2_X1 U6470 ( .A1(n6425), .A2(n6400), .ZN(n9215) );
  INV_X1 U6471 ( .A(n9501), .ZN(n9397) );
  INV_X1 U6472 ( .A(n9109), .ZN(n9075) );
  AND3_X1 U6473 ( .A1(n6337), .A2(n6336), .A3(n6335), .ZN(n9421) );
  NAND2_X1 U6474 ( .A1(n6194), .A2(n6193), .ZN(n9446) );
  INV_X1 U6475 ( .A(P1_U3973), .ZN(n9126) );
  OR2_X1 U6476 ( .A1(n6476), .A2(n9138), .ZN(n9165) );
  OR2_X1 U6477 ( .A1(n6476), .A2(n6452), .ZN(n9189) );
  INV_X1 U6478 ( .A(n9586), .ZN(n9414) );
  AND2_X2 U6479 ( .A1(n6561), .A2(n6742), .ZN(n9740) );
  NAND2_X1 U6480 ( .A1(n9717), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6376) );
  INV_X1 U6481 ( .A(n9719), .ZN(n9717) );
  AND2_X1 U6482 ( .A1(n7775), .A2(n7755), .ZN(n6411) );
  INV_X1 U6483 ( .A(n8072), .ZN(n7593) );
  INV_X1 U6484 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7262) );
  INV_X1 U6485 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6860) );
  AND2_X2 U6486 ( .A1(n6379), .A2(n6378), .ZN(P1_U3973) );
  NAND2_X1 U6487 ( .A1(n5004), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5002) );
  INV_X1 U6488 ( .A(SI_1_), .ZN(n5005) );
  NAND2_X1 U6489 ( .A1(n5011), .A2(SI_0_), .ZN(n5199) );
  INV_X1 U6490 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5007) );
  AND2_X1 U6491 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U6492 ( .A1(n7922), .A2(n5006), .ZN(n5748) );
  NAND2_X1 U6493 ( .A1(n5189), .A2(n5188), .ZN(n5010) );
  NAND2_X1 U6494 ( .A1(n5008), .A2(SI_1_), .ZN(n5009) );
  NAND2_X1 U6495 ( .A1(n5010), .A2(n5009), .ZN(n5205) );
  MUX2_X1 U6496 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n5004), .Z(n5013) );
  INV_X1 U6497 ( .A(SI_2_), .ZN(n5012) );
  XNOR2_X1 U6498 ( .A(n5013), .B(n5012), .ZN(n5206) );
  NAND2_X1 U6499 ( .A1(n5205), .A2(n5206), .ZN(n5015) );
  NAND2_X1 U6500 ( .A1(n5013), .A2(SI_2_), .ZN(n5014) );
  NAND2_X1 U6501 ( .A1(n5015), .A2(n5014), .ZN(n5224) );
  MUX2_X1 U6502 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7922), .Z(n5017) );
  INV_X1 U6503 ( .A(SI_3_), .ZN(n5016) );
  XNOR2_X1 U6504 ( .A(n5017), .B(n5016), .ZN(n5225) );
  NAND2_X1 U6505 ( .A1(n5224), .A2(n5225), .ZN(n5019) );
  NAND2_X1 U6506 ( .A1(n5017), .A2(SI_3_), .ZN(n5018) );
  NAND2_X1 U6507 ( .A1(n5019), .A2(n5018), .ZN(n5238) );
  MUX2_X1 U6508 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7922), .Z(n5021) );
  INV_X1 U6509 ( .A(SI_4_), .ZN(n5020) );
  XNOR2_X1 U6510 ( .A(n5021), .B(n5020), .ZN(n5239) );
  NAND2_X1 U6511 ( .A1(n5021), .A2(SI_4_), .ZN(n5022) );
  INV_X1 U6512 ( .A(SI_5_), .ZN(n5023) );
  XNOR2_X1 U6513 ( .A(n5024), .B(n5023), .ZN(n5255) );
  MUX2_X1 U6514 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7922), .Z(n5026) );
  INV_X1 U6515 ( .A(SI_6_), .ZN(n5025) );
  XNOR2_X1 U6516 ( .A(n5026), .B(n5025), .ZN(n5268) );
  NAND2_X1 U6517 ( .A1(n5026), .A2(SI_6_), .ZN(n5027) );
  MUX2_X1 U6518 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7922), .Z(n5028) );
  INV_X1 U6519 ( .A(SI_7_), .ZN(n10184) );
  XNOR2_X1 U6520 ( .A(n5028), .B(n10184), .ZN(n5284) );
  NAND2_X1 U6521 ( .A1(n5028), .A2(SI_7_), .ZN(n5029) );
  INV_X1 U6522 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6441) );
  INV_X1 U6523 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5031) );
  MUX2_X1 U6524 ( .A(n6441), .B(n5031), .S(n7922), .Z(n5033) );
  INV_X1 U6525 ( .A(SI_8_), .ZN(n5032) );
  NAND2_X1 U6526 ( .A1(n5033), .A2(n5032), .ZN(n5036) );
  INV_X1 U6527 ( .A(n5033), .ZN(n5034) );
  NAND2_X1 U6528 ( .A1(n5034), .A2(SI_8_), .ZN(n5035) );
  NAND2_X1 U6529 ( .A1(n5036), .A2(n5035), .ZN(n5309) );
  INV_X1 U6530 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6517) );
  INV_X1 U6531 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6516) );
  MUX2_X1 U6532 ( .A(n6517), .B(n6516), .S(n7922), .Z(n5037) );
  NAND2_X1 U6533 ( .A1(n5037), .A2(n10188), .ZN(n5040) );
  INV_X1 U6534 ( .A(n5037), .ZN(n5038) );
  NAND2_X1 U6535 ( .A1(n5038), .A2(SI_9_), .ZN(n5039) );
  MUX2_X1 U6536 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n7922), .Z(n5041) );
  XNOR2_X1 U6537 ( .A(n5041), .B(n10038), .ZN(n5319) );
  MUX2_X1 U6538 ( .A(n6565), .B(n6564), .S(n4713), .Z(n5042) );
  NAND2_X1 U6539 ( .A1(n5042), .A2(n10206), .ZN(n5045) );
  INV_X1 U6540 ( .A(n5042), .ZN(n5043) );
  NAND2_X1 U6541 ( .A1(n5043), .A2(SI_11_), .ZN(n5044) );
  NAND2_X1 U6542 ( .A1(n5045), .A2(n5044), .ZN(n5335) );
  MUX2_X1 U6543 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7922), .Z(n5047) );
  INV_X1 U6544 ( .A(SI_12_), .ZN(n5046) );
  XNOR2_X1 U6545 ( .A(n5047), .B(n5046), .ZN(n5348) );
  NAND2_X1 U6546 ( .A1(n5047), .A2(SI_12_), .ZN(n5048) );
  MUX2_X1 U6547 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7922), .Z(n5049) );
  XNOR2_X1 U6548 ( .A(n5049), .B(SI_13_), .ZN(n5363) );
  MUX2_X1 U6549 ( .A(n6861), .B(n6860), .S(n4713), .Z(n5050) );
  NAND2_X1 U6550 ( .A1(n5050), .A2(n10050), .ZN(n5053) );
  INV_X1 U6551 ( .A(n5050), .ZN(n5051) );
  NAND2_X1 U6552 ( .A1(n5051), .A2(SI_14_), .ZN(n5052) );
  NAND2_X1 U6553 ( .A1(n5053), .A2(n5052), .ZN(n5374) );
  MUX2_X1 U6554 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4713), .Z(n5388) );
  NAND2_X1 U6555 ( .A1(n5388), .A2(SI_15_), .ZN(n5054) );
  NAND2_X1 U6556 ( .A1(n5390), .A2(n5054), .ZN(n5057) );
  INV_X1 U6557 ( .A(n5388), .ZN(n5055) );
  NAND2_X1 U6558 ( .A1(n5055), .A2(n10118), .ZN(n5056) );
  MUX2_X1 U6559 ( .A(n6983), .B(n6984), .S(n4713), .Z(n5406) );
  NOR2_X1 U6560 ( .A1(n5058), .A2(SI_16_), .ZN(n5060) );
  NAND2_X1 U6561 ( .A1(n5058), .A2(SI_16_), .ZN(n5059) );
  MUX2_X1 U6562 ( .A(n7095), .B(n5061), .S(n4713), .Z(n5063) );
  NAND2_X1 U6563 ( .A1(n5063), .A2(n5062), .ZN(n5066) );
  INV_X1 U6564 ( .A(n5063), .ZN(n5064) );
  NAND2_X1 U6565 ( .A1(n5064), .A2(SI_17_), .ZN(n5065) );
  NAND2_X1 U6566 ( .A1(n5066), .A2(n5065), .ZN(n5419) );
  MUX2_X1 U6567 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4713), .Z(n5067) );
  XNOR2_X1 U6568 ( .A(n5067), .B(n10162), .ZN(n5164) );
  INV_X1 U6569 ( .A(n5152), .ZN(n5073) );
  MUX2_X1 U6570 ( .A(n7263), .B(n7262), .S(n4713), .Z(n5069) );
  INV_X1 U6571 ( .A(SI_19_), .ZN(n5068) );
  NAND2_X1 U6572 ( .A1(n5069), .A2(n5068), .ZN(n5074) );
  INV_X1 U6573 ( .A(n5069), .ZN(n5070) );
  NAND2_X1 U6574 ( .A1(n5070), .A2(SI_19_), .ZN(n5071) );
  NAND2_X1 U6575 ( .A1(n5074), .A2(n5071), .ZN(n5151) );
  INV_X1 U6576 ( .A(n5151), .ZN(n5072) );
  NAND2_X1 U6577 ( .A1(n5073), .A2(n5072), .ZN(n5075) );
  NAND2_X1 U6578 ( .A1(n5075), .A2(n5074), .ZN(n5439) );
  MUX2_X1 U6579 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n4713), .Z(n5437) );
  INV_X1 U6580 ( .A(n5437), .ZN(n5076) );
  MUX2_X1 U6581 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n4713), .Z(n5077) );
  NAND2_X1 U6582 ( .A1(n5077), .A2(SI_21_), .ZN(n5078) );
  OAI21_X1 U6583 ( .B1(n5077), .B2(SI_21_), .A(n5078), .ZN(n5446) );
  MUX2_X1 U6584 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n4713), .Z(n5079) );
  XNOR2_X1 U6585 ( .A(n5079), .B(SI_22_), .ZN(n5461) );
  INV_X1 U6586 ( .A(n5079), .ZN(n5081) );
  INV_X1 U6587 ( .A(SI_22_), .ZN(n5080) );
  NAND2_X1 U6588 ( .A1(n5081), .A2(n5080), .ZN(n5082) );
  MUX2_X1 U6589 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n4713), .Z(n5084) );
  XNOR2_X1 U6590 ( .A(n5084), .B(n5085), .ZN(n5472) );
  INV_X1 U6591 ( .A(n5084), .ZN(n5086) );
  NAND2_X1 U6592 ( .A1(n5086), .A2(n5085), .ZN(n5087) );
  MUX2_X1 U6593 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4713), .Z(n5088) );
  XNOR2_X1 U6594 ( .A(n5088), .B(n10058), .ZN(n5484) );
  INV_X1 U6595 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6596 ( .A1(n5089), .A2(n10058), .ZN(n5090) );
  NAND2_X1 U6597 ( .A1(n5091), .A2(n5090), .ZN(n5497) );
  MUX2_X1 U6598 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n4713), .Z(n5498) );
  INV_X1 U6599 ( .A(SI_25_), .ZN(n5499) );
  XNOR2_X1 U6600 ( .A(n5498), .B(n5499), .ZN(n5496) );
  XNOR2_X1 U6601 ( .A(n5497), .B(n5496), .ZN(n7750) );
  NOR2_X1 U6602 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5094) );
  NAND4_X1 U6603 ( .A1(n5094), .A2(n5093), .A3(n5092), .A4(n5240), .ZN(n5096)
         );
  NOR2_X2 U6604 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5184) );
  NAND2_X1 U6605 ( .A1(n5184), .A2(n5095), .ZN(n5221) );
  NOR2_X1 U6606 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5097) );
  NAND4_X1 U6607 ( .A1(n5097), .A2(n5376), .A3(n5158), .A4(n4474), .ZN(n5100)
         );
  NAND4_X1 U6608 ( .A1(n5155), .A2(n5154), .A3(n5157), .A4(n5098), .ZN(n5099)
         );
  NOR2_X1 U6609 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  INV_X1 U6610 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U6611 ( .A1(n7750), .A2(n8329), .ZN(n5109) );
  INV_X1 U6612 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7751) );
  OR2_X1 U6613 ( .A1(n8331), .A2(n7751), .ZN(n5108) );
  INV_X1 U6614 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9844) );
  INV_X1 U6615 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6616 ( .A1(n9844), .A2(n5110), .ZN(n5246) );
  INV_X1 U6617 ( .A(n5246), .ZN(n5112) );
  INV_X1 U6618 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6619 ( .A1(n5112), .A2(n5111), .ZN(n5260) );
  INV_X1 U6620 ( .A(n5278), .ZN(n5113) );
  NAND2_X1 U6621 ( .A1(n5113), .A2(n10163), .ZN(n5301) );
  INV_X1 U6622 ( .A(n5303), .ZN(n5115) );
  NAND2_X1 U6623 ( .A1(n5115), .A2(n5114), .ZN(n5326) );
  NAND2_X1 U6624 ( .A1(n5116), .A2(n10040), .ZN(n5368) );
  INV_X1 U6625 ( .A(n5368), .ZN(n5118) );
  NAND2_X1 U6626 ( .A1(n5118), .A2(n5117), .ZN(n5381) );
  INV_X1 U6627 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5122) );
  INV_X1 U6628 ( .A(n5490), .ZN(n5128) );
  INV_X1 U6629 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6630 ( .A1(n5490), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6631 ( .A1(n5505), .A2(n5129), .ZN(n8739) );
  XNOR2_X2 U6632 ( .A(n5132), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5137) );
  NAND2_X2 U6633 ( .A1(n5137), .A2(n5136), .ZN(n5200) );
  NAND2_X1 U6634 ( .A1(n8739), .A2(n5545), .ZN(n5142) );
  INV_X1 U6635 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8906) );
  INV_X1 U6636 ( .A(n5137), .ZN(n8126) );
  OR2_X2 U6637 ( .A1(n5137), .A2(n8206), .ZN(n5429) );
  NAND2_X1 U6638 ( .A1(n5598), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5139) );
  NAND2_X2 U6639 ( .A1(n5137), .A2(n8206), .ZN(n8336) );
  NAND2_X1 U6640 ( .A1(n5193), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5138) );
  OAI211_X1 U6641 ( .C1(n8906), .C2(n5601), .A(n5139), .B(n5138), .ZN(n5140)
         );
  INV_X1 U6642 ( .A(n5140), .ZN(n5141) );
  NAND2_X1 U6643 ( .A1(n5173), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6644 ( .A1(n5442), .A2(n5143), .ZN(n8805) );
  NAND2_X1 U6645 ( .A1(n5545), .A2(n8805), .ZN(n5150) );
  INV_X1 U6646 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n5144) );
  OR2_X1 U6647 ( .A1(n5429), .A2(n5144), .ZN(n5149) );
  INV_X1 U6648 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5145) );
  OR2_X1 U6649 ( .A1(n8336), .A2(n5145), .ZN(n5148) );
  INV_X1 U6650 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n5146) );
  OR2_X1 U6651 ( .A1(n5601), .A2(n5146), .ZN(n5147) );
  NAND4_X1 U6652 ( .A1(n5150), .A2(n5149), .A3(n5148), .A4(n5147), .ZN(n8817)
         );
  XNOR2_X1 U6653 ( .A(n5152), .B(n5151), .ZN(n7261) );
  NAND2_X1 U6654 ( .A1(n7261), .A2(n8329), .ZN(n5163) );
  NAND2_X1 U6655 ( .A1(n5153), .A2(n5154), .ZN(n5350) );
  NAND3_X1 U6656 ( .A1(n5376), .A2(n5391), .A3(n5155), .ZN(n5156) );
  NAND2_X1 U6657 ( .A1(n5409), .A2(n5157), .ZN(n5421) );
  INV_X1 U6658 ( .A(n5421), .ZN(n5159) );
  NAND2_X1 U6659 ( .A1(n5159), .A2(n5158), .ZN(n5160) );
  NAND2_X1 U6660 ( .A1(n5160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5167) );
  NAND2_X1 U6661 ( .A1(n5167), .A2(n5166), .ZN(n5169) );
  XNOR2_X2 U6662 ( .A(n5161), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8663) );
  AOI22_X1 U6663 ( .A1(n5423), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8663), .B2(
        n6384), .ZN(n5162) );
  INV_X1 U6664 ( .A(n8867), .ZN(n8808) );
  XNOR2_X1 U6665 ( .A(n5165), .B(n5164), .ZN(n7108) );
  NAND2_X1 U6666 ( .A1(n7108), .A2(n8329), .ZN(n5171) );
  OR2_X1 U6667 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  AND2_X1 U6668 ( .A1(n5169), .A2(n5168), .ZN(n8668) );
  AOI22_X1 U6669 ( .A1(n5423), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6384), .B2(
        n8668), .ZN(n5170) );
  INV_X1 U6670 ( .A(n8944), .ZN(n5582) );
  NAND2_X1 U6671 ( .A1(n5428), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5172) );
  NAND2_X1 U6672 ( .A1(n5173), .A2(n5172), .ZN(n8820) );
  NAND2_X1 U6673 ( .A1(n5545), .A2(n8820), .ZN(n5177) );
  INV_X1 U6674 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8819) );
  OR2_X1 U6675 ( .A1(n8336), .A2(n8819), .ZN(n5176) );
  INV_X1 U6676 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8943) );
  OR2_X1 U6677 ( .A1(n5601), .A2(n8943), .ZN(n5175) );
  INV_X1 U6678 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8871) );
  OR2_X1 U6679 ( .A1(n5429), .A2(n8871), .ZN(n5174) );
  NAND4_X1 U6680 ( .A1(n5177), .A2(n5176), .A3(n5175), .A4(n5174), .ZN(n8827)
         );
  INV_X1 U6681 ( .A(n8827), .ZN(n8137) );
  NAND2_X1 U6682 ( .A1(n5214), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5182) );
  INV_X1 U6683 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6889) );
  INV_X1 U6684 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5178) );
  INV_X1 U6685 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6640) );
  OR2_X1 U6686 ( .A1(n5200), .A2(n6640), .ZN(n5179) );
  NAND2_X1 U6687 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5183) );
  MUX2_X1 U6688 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5183), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5186) );
  INV_X1 U6689 ( .A(n5207), .ZN(n5185) );
  OR2_X1 U6690 ( .A1(n5187), .A2(n6641), .ZN(n5191) );
  XNOR2_X1 U6691 ( .A(n5189), .B(n5188), .ZN(n6403) );
  NAND2_X1 U6692 ( .A1(n5214), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U6693 ( .A1(n5193), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5196) );
  INV_X1 U6694 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6667) );
  INV_X1 U6695 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6604) );
  OR2_X1 U6696 ( .A1(n5429), .A2(n6604), .ZN(n5194) );
  NAND4_X1 U6697 ( .A1(n5197), .A2(n5196), .A3(n5195), .A4(n5194), .ZN(n5567)
         );
  CLKBUF_X1 U6698 ( .A(n5567), .Z(n5198) );
  XNOR2_X1 U6699 ( .A(n5199), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8969) );
  MUX2_X1 U6700 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8969), .S(n5187), .Z(n6577) );
  NAND2_X1 U6701 ( .A1(n5198), .A2(n6577), .ZN(n6881) );
  OR2_X1 U6702 ( .A1(n6675), .A2(n6886), .ZN(n9847) );
  NAND2_X1 U6703 ( .A1(n9848), .A2(n9847), .ZN(n5211) );
  NAND2_X1 U6704 ( .A1(n5193), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5204) );
  INV_X1 U6705 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6603) );
  OR2_X1 U6706 ( .A1(n5429), .A2(n6603), .ZN(n5202) );
  INV_X1 U6707 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9863) );
  OR2_X1 U6708 ( .A1(n5200), .A2(n9863), .ZN(n5201) );
  NAND4_X2 U6709 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n9837)
         );
  XNOR2_X1 U6710 ( .A(n5205), .B(n5206), .ZN(n6401) );
  OR2_X1 U6711 ( .A1(n5450), .A2(n6401), .ZN(n5210) );
  INV_X1 U6712 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6388) );
  OR2_X1 U6713 ( .A1(n5226), .A2(n6388), .ZN(n5209) );
  NAND2_X1 U6714 ( .A1(n5207), .A2(n4945), .ZN(n5219) );
  OR2_X1 U6715 ( .A1(n5187), .A2(n4353), .ZN(n5208) );
  NAND2_X1 U6716 ( .A1(n9837), .A2(n9861), .ZN(n8392) );
  NAND2_X1 U6717 ( .A1(n8390), .A2(n8392), .ZN(n8354) );
  NAND2_X1 U6718 ( .A1(n5211), .A2(n8354), .ZN(n9850) );
  INV_X1 U6719 ( .A(n9861), .ZN(n5212) );
  OR2_X1 U6720 ( .A1(n9837), .A2(n5212), .ZN(n5213) );
  NAND2_X1 U6721 ( .A1(n9850), .A2(n5213), .ZN(n9836) );
  NAND2_X1 U6722 ( .A1(n5214), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5218) );
  OR2_X1 U6723 ( .A1(n5200), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5217) );
  INV_X1 U6724 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6598) );
  OR2_X1 U6725 ( .A1(n8336), .A2(n6598), .ZN(n5216) );
  INV_X1 U6726 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6597) );
  OR2_X1 U6727 ( .A1(n5429), .A2(n6597), .ZN(n5215) );
  NAND2_X1 U6728 ( .A1(n5219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5220) );
  MUX2_X1 U6729 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5220), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5223) );
  NAND2_X1 U6730 ( .A1(n5223), .A2(n5222), .ZN(n9745) );
  XNOR2_X1 U6731 ( .A(n5224), .B(n5225), .ZN(n6387) );
  OR2_X1 U6732 ( .A1(n5450), .A2(n6387), .ZN(n5228) );
  INV_X1 U6733 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6386) );
  OR2_X1 U6734 ( .A1(n5226), .A2(n6386), .ZN(n5227) );
  OAI211_X1 U6735 ( .C1(n5187), .C2(n9745), .A(n5228), .B(n5227), .ZN(n9883)
         );
  NAND2_X1 U6736 ( .A1(n9854), .A2(n9883), .ZN(n5229) );
  NAND2_X1 U6737 ( .A1(n9836), .A2(n5229), .ZN(n5231) );
  OR2_X1 U6738 ( .A1(n9854), .A2(n9883), .ZN(n5230) );
  NAND2_X1 U6739 ( .A1(n5231), .A2(n5230), .ZN(n7014) );
  NAND2_X1 U6740 ( .A1(n5193), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5237) );
  INV_X1 U6741 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6609) );
  OR2_X1 U6742 ( .A1(n5429), .A2(n6609), .ZN(n5236) );
  NAND2_X1 U6743 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5232) );
  AND2_X1 U6744 ( .A1(n5246), .A2(n5232), .ZN(n6942) );
  OR2_X1 U6745 ( .A1(n5200), .A2(n6942), .ZN(n5235) );
  INV_X1 U6746 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5233) );
  XNOR2_X1 U6747 ( .A(n5238), .B(n5239), .ZN(n6390) );
  OR2_X1 U6748 ( .A1(n5450), .A2(n6390), .ZN(n5244) );
  INV_X1 U6749 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6389) );
  OR2_X1 U6750 ( .A1(n5226), .A2(n6389), .ZN(n5243) );
  NAND2_X1 U6751 ( .A1(n5222), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5241) );
  XNOR2_X1 U6752 ( .A(n5241), .B(n5240), .ZN(n6707) );
  OR2_X1 U6753 ( .A1(n5187), .A2(n6707), .ZN(n5242) );
  NAND2_X1 U6754 ( .A1(n9838), .A2(n9889), .ZN(n8400) );
  INV_X1 U6755 ( .A(n9889), .ZN(n7018) );
  OR2_X1 U6756 ( .A1(n9838), .A2(n7018), .ZN(n5245) );
  NAND2_X1 U6757 ( .A1(n5214), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5251) );
  INV_X1 U6758 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6689) );
  OR2_X1 U6759 ( .A1(n5429), .A2(n6689), .ZN(n5250) );
  INV_X1 U6760 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6690) );
  OR2_X1 U6761 ( .A1(n8336), .A2(n6690), .ZN(n5249) );
  NAND2_X1 U6762 ( .A1(n5246), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5247) );
  AND2_X1 U6763 ( .A1(n5260), .A2(n5247), .ZN(n7090) );
  OR2_X1 U6764 ( .A1(n5200), .A2(n7090), .ZN(n5248) );
  NAND4_X1 U6765 ( .A1(n5251), .A2(n5250), .A3(n5249), .A4(n5248), .ZN(n8587)
         );
  OR2_X1 U6766 ( .A1(n5222), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5269) );
  NAND2_X1 U6767 ( .A1(n5269), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5253) );
  INV_X1 U6768 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5252) );
  XNOR2_X1 U6769 ( .A(n5253), .B(n5252), .ZN(n6730) );
  OR2_X1 U6770 ( .A1(n5450), .A2(n6393), .ZN(n5257) );
  INV_X1 U6771 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6392) );
  OR2_X1 U6772 ( .A1(n8331), .A2(n6392), .ZN(n5256) );
  OAI211_X1 U6773 ( .C1(n5187), .C2(n6730), .A(n5257), .B(n5256), .ZN(n7078)
         );
  NAND2_X1 U6774 ( .A1(n8587), .A2(n7078), .ZN(n5258) );
  NAND2_X1 U6775 ( .A1(n5598), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5266) );
  INV_X1 U6776 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7195) );
  OR2_X1 U6777 ( .A1(n8336), .A2(n7195), .ZN(n5265) );
  NAND2_X1 U6778 ( .A1(n5260), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5261) );
  AND2_X1 U6779 ( .A1(n5278), .A2(n5261), .ZN(n7177) );
  OR2_X1 U6780 ( .A1(n5200), .A2(n7177), .ZN(n5264) );
  INV_X1 U6781 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5262) );
  OR2_X1 U6782 ( .A1(n5601), .A2(n5262), .ZN(n5263) );
  XNOR2_X1 U6783 ( .A(n5267), .B(n5268), .ZN(n6396) );
  OR2_X1 U6784 ( .A1(n5450), .A2(n6396), .ZN(n5277) );
  INV_X1 U6785 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6397) );
  OR2_X1 U6786 ( .A1(n8331), .A2(n6397), .ZN(n5276) );
  NOR2_X1 U6787 ( .A1(n5269), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5273) );
  NOR2_X1 U6788 ( .A1(n5273), .A2(n5133), .ZN(n5270) );
  MUX2_X1 U6789 ( .A(n5270), .B(n5133), .S(n5272), .Z(n5271) );
  INV_X1 U6790 ( .A(n5271), .ZN(n5274) );
  NAND2_X1 U6791 ( .A1(n5273), .A2(n5272), .ZN(n5296) );
  NAND2_X1 U6792 ( .A1(n5274), .A2(n5296), .ZN(n6832) );
  OR2_X1 U6793 ( .A1(n5187), .A2(n6832), .ZN(n5275) );
  OR2_X1 U6794 ( .A1(n8586), .A2(n9900), .ZN(n5572) );
  NAND2_X1 U6795 ( .A1(n8586), .A2(n9900), .ZN(n8410) );
  NAND2_X1 U6796 ( .A1(n5214), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5283) );
  INV_X1 U6797 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6827) );
  OR2_X1 U6798 ( .A1(n5429), .A2(n6827), .ZN(n5282) );
  INV_X1 U6799 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6828) );
  OR2_X1 U6800 ( .A1(n8336), .A2(n6828), .ZN(n5281) );
  NAND2_X1 U6801 ( .A1(n5278), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5279) );
  AND2_X1 U6802 ( .A1(n5301), .A2(n5279), .ZN(n7256) );
  OR2_X1 U6803 ( .A1(n5200), .A2(n7256), .ZN(n5280) );
  OR2_X1 U6804 ( .A1(n6420), .A2(n5450), .ZN(n5290) );
  INV_X1 U6805 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6419) );
  OR2_X1 U6806 ( .A1(n8331), .A2(n6419), .ZN(n5289) );
  NAND2_X1 U6807 ( .A1(n5296), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5287) );
  INV_X1 U6808 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5286) );
  OR2_X1 U6809 ( .A1(n5187), .A2(n7225), .ZN(n5288) );
  NAND2_X1 U6810 ( .A1(n8585), .A2(n9903), .ZN(n7160) );
  INV_X1 U6811 ( .A(n8416), .ZN(n7250) );
  NAND2_X1 U6812 ( .A1(n5214), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5295) );
  INV_X1 U6813 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7219) );
  OR2_X1 U6814 ( .A1(n5429), .A2(n7219), .ZN(n5294) );
  INV_X1 U6815 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7220) );
  OR2_X1 U6816 ( .A1(n8336), .A2(n7220), .ZN(n5293) );
  NAND2_X1 U6817 ( .A1(n5303), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5291) );
  AND2_X1 U6818 ( .A1(n5326), .A2(n5291), .ZN(n7287) );
  OR2_X1 U6819 ( .A1(n5200), .A2(n7287), .ZN(n5292) );
  NAND2_X1 U6820 ( .A1(n6514), .A2(n8329), .ZN(n5299) );
  OAI21_X1 U6821 ( .B1(n5311), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5297) );
  XNOR2_X1 U6822 ( .A(n5297), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7323) );
  AOI22_X1 U6823 ( .A1(n5423), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6384), .B2(
        n7323), .ZN(n5298) );
  NAND2_X1 U6824 ( .A1(n5299), .A2(n5298), .ZN(n7378) );
  OR2_X1 U6825 ( .A1(n7614), .A2(n7378), .ZN(n8419) );
  NAND2_X1 U6826 ( .A1(n7614), .A2(n7378), .ZN(n8426) );
  INV_X1 U6827 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5300) );
  OR2_X1 U6828 ( .A1(n8336), .A2(n7215), .ZN(n5307) );
  NAND2_X1 U6829 ( .A1(n5301), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5302) );
  AND2_X1 U6830 ( .A1(n5303), .A2(n5302), .ZN(n7310) );
  OR2_X1 U6831 ( .A1(n5200), .A2(n7310), .ZN(n5306) );
  INV_X1 U6832 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5304) );
  OR2_X1 U6833 ( .A1(n5601), .A2(n5304), .ZN(n5305) );
  NAND4_X1 U6834 ( .A1(n5308), .A2(n5307), .A3(n5306), .A4(n5305), .ZN(n8584)
         );
  XNOR2_X1 U6835 ( .A(n5310), .B(n5309), .ZN(n6430) );
  NAND2_X1 U6836 ( .A1(n6430), .A2(n8329), .ZN(n5314) );
  NAND2_X1 U6837 ( .A1(n5311), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5312) );
  XNOR2_X1 U6838 ( .A(n5312), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7214) );
  AOI22_X1 U6839 ( .A1(n5423), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6384), .B2(
        n7214), .ZN(n5313) );
  NAND2_X1 U6840 ( .A1(n8584), .A2(n7315), .ZN(n7279) );
  NAND2_X1 U6841 ( .A1(n8361), .A2(n7279), .ZN(n5317) );
  OR2_X1 U6842 ( .A1(n7149), .A2(n5317), .ZN(n5315) );
  OR2_X1 U6843 ( .A1(n7378), .A2(n8583), .ZN(n7267) );
  OR2_X1 U6844 ( .A1(n8584), .A2(n9909), .ZN(n8425) );
  NAND2_X1 U6845 ( .A1(n8584), .A2(n9909), .ZN(n8418) );
  NAND2_X1 U6846 ( .A1(n8425), .A2(n8418), .ZN(n8360) );
  INV_X1 U6847 ( .A(n9903), .ZN(n7258) );
  OR2_X1 U6848 ( .A1(n8585), .A2(n7258), .ZN(n7151) );
  AND2_X1 U6849 ( .A1(n8360), .A2(n7151), .ZN(n5316) );
  INV_X1 U6850 ( .A(n9900), .ZN(n7197) );
  OR2_X1 U6851 ( .A1(n8586), .A2(n7197), .ZN(n7249) );
  OR2_X1 U6852 ( .A1(n7250), .A2(n7249), .ZN(n7150) );
  XNOR2_X1 U6853 ( .A(n5320), .B(n5319), .ZN(n6524) );
  NAND2_X1 U6854 ( .A1(n6524), .A2(n8329), .ZN(n5325) );
  NOR2_X1 U6855 ( .A1(n5321), .A2(n5133), .ZN(n5322) );
  MUX2_X1 U6856 ( .A(n5133), .B(n5322), .S(P2_IR_REG_10__SCAN_IN), .Z(n5323)
         );
  OR2_X1 U6857 ( .A1(n5323), .A2(n5153), .ZN(n7463) );
  INV_X1 U6858 ( .A(n7463), .ZN(n7338) );
  AOI22_X1 U6859 ( .A1(n5423), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6384), .B2(
        n7338), .ZN(n5324) );
  NAND2_X1 U6860 ( .A1(n5325), .A2(n5324), .ZN(n9921) );
  NAND2_X1 U6861 ( .A1(n5598), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5332) );
  INV_X1 U6862 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7331) );
  OR2_X1 U6863 ( .A1(n8336), .A2(n7331), .ZN(n5331) );
  NAND2_X1 U6864 ( .A1(n5326), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5327) );
  AND2_X1 U6865 ( .A1(n5340), .A2(n5327), .ZN(n7619) );
  OR2_X1 U6866 ( .A1(n5200), .A2(n7619), .ZN(n5330) );
  INV_X1 U6867 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5328) );
  OR2_X1 U6868 ( .A1(n5601), .A2(n5328), .ZN(n5329) );
  OR2_X1 U6869 ( .A1(n9921), .A2(n7674), .ZN(n8438) );
  NAND2_X1 U6870 ( .A1(n9921), .A2(n7674), .ZN(n8434) );
  NAND2_X1 U6871 ( .A1(n8438), .A2(n8434), .ZN(n7274) );
  OR2_X1 U6872 ( .A1(n9921), .A2(n8582), .ZN(n5334) );
  XNOR2_X1 U6873 ( .A(n5336), .B(n5335), .ZN(n6563) );
  NAND2_X1 U6874 ( .A1(n6563), .A2(n8329), .ZN(n5339) );
  OR2_X1 U6875 ( .A1(n5153), .A2(n5133), .ZN(n5337) );
  XNOR2_X1 U6876 ( .A(n5337), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7466) );
  AOI22_X1 U6877 ( .A1(n5423), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6384), .B2(
        n7466), .ZN(n5338) );
  NAND2_X1 U6878 ( .A1(n5339), .A2(n5338), .ZN(n9929) );
  NAND2_X1 U6879 ( .A1(n5214), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5345) );
  INV_X1 U6880 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7450) );
  OR2_X1 U6881 ( .A1(n5429), .A2(n7450), .ZN(n5344) );
  INV_X1 U6882 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7451) );
  OR2_X1 U6883 ( .A1(n8336), .A2(n7451), .ZN(n5343) );
  NAND2_X1 U6884 ( .A1(n5340), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5341) );
  AND2_X1 U6885 ( .A1(n5354), .A2(n5341), .ZN(n7653) );
  OR2_X1 U6886 ( .A1(n5200), .A2(n7653), .ZN(n5342) );
  NAND4_X1 U6887 ( .A1(n5345), .A2(n5344), .A3(n5343), .A4(n5342), .ZN(n8581)
         );
  NAND2_X1 U6888 ( .A1(n9929), .A2(n8581), .ZN(n5346) );
  OR2_X1 U6889 ( .A1(n9929), .A2(n8581), .ZN(n5347) );
  INV_X1 U6890 ( .A(n7545), .ZN(n5361) );
  NAND2_X1 U6891 ( .A1(n6654), .A2(n8329), .ZN(n5353) );
  NAND2_X1 U6892 ( .A1(n5350), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5351) );
  XNOR2_X1 U6893 ( .A(n5351), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7580) );
  AOI22_X1 U6894 ( .A1(n5423), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6384), .B2(
        n7580), .ZN(n5352) );
  NAND2_X1 U6895 ( .A1(n5353), .A2(n5352), .ZN(n7688) );
  NAND2_X1 U6896 ( .A1(n5214), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5359) );
  INV_X1 U6897 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7566) );
  OR2_X1 U6898 ( .A1(n5429), .A2(n7566), .ZN(n5358) );
  OR2_X1 U6899 ( .A1(n8336), .A2(n7579), .ZN(n5357) );
  NAND2_X1 U6900 ( .A1(n5354), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5355) );
  AND2_X1 U6901 ( .A1(n5368), .A2(n5355), .ZN(n7672) );
  OR2_X1 U6902 ( .A1(n5200), .A2(n7672), .ZN(n5356) );
  OR2_X1 U6903 ( .A1(n7688), .A2(n7673), .ZN(n8447) );
  NAND2_X1 U6904 ( .A1(n7688), .A2(n7673), .ZN(n8448) );
  INV_X1 U6905 ( .A(n7673), .ZN(n8580) );
  NAND2_X1 U6906 ( .A1(n7688), .A2(n8580), .ZN(n5362) );
  XNOR2_X1 U6907 ( .A(n5364), .B(n5363), .ZN(n6682) );
  NAND2_X1 U6908 ( .A1(n6682), .A2(n8329), .ZN(n5367) );
  NAND2_X1 U6909 ( .A1(n5365), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5377) );
  XNOR2_X1 U6910 ( .A(n5377), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8604) );
  AOI22_X1 U6911 ( .A1(n5423), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6384), .B2(
        n8604), .ZN(n5366) );
  NAND2_X1 U6912 ( .A1(n5214), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5373) );
  INV_X1 U6913 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7576) );
  OR2_X1 U6914 ( .A1(n5429), .A2(n7576), .ZN(n5372) );
  INV_X1 U6915 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7584) );
  OR2_X1 U6916 ( .A1(n8336), .A2(n7584), .ZN(n5371) );
  NAND2_X1 U6917 ( .A1(n5368), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5369) );
  AND2_X1 U6918 ( .A1(n5381), .A2(n5369), .ZN(n7695) );
  OR2_X1 U6919 ( .A1(n5200), .A2(n7695), .ZN(n5370) );
  NAND4_X1 U6920 ( .A1(n5373), .A2(n5372), .A3(n5371), .A4(n5370), .ZN(n8579)
         );
  OR2_X1 U6921 ( .A1(n8451), .A2(n8579), .ZN(n8454) );
  NAND2_X1 U6922 ( .A1(n8451), .A2(n8579), .ZN(n8457) );
  XNOR2_X1 U6923 ( .A(n5375), .B(n5374), .ZN(n6859) );
  NAND2_X1 U6924 ( .A1(n6859), .A2(n8329), .ZN(n5380) );
  NAND2_X1 U6925 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  NAND2_X1 U6926 ( .A1(n5378), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5392) );
  XNOR2_X1 U6927 ( .A(n5392), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8608) );
  AOI22_X1 U6928 ( .A1(n5423), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6384), .B2(
        n8608), .ZN(n5379) );
  NAND2_X1 U6929 ( .A1(n5214), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5386) );
  INV_X1 U6930 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8589) );
  OR2_X1 U6931 ( .A1(n5429), .A2(n8589), .ZN(n5385) );
  INV_X1 U6932 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8607) );
  OR2_X1 U6933 ( .A1(n8336), .A2(n8607), .ZN(n5384) );
  NAND2_X1 U6934 ( .A1(n5381), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5382) );
  AND2_X1 U6935 ( .A1(n5397), .A2(n5382), .ZN(n7728) );
  OR2_X1 U6936 ( .A1(n5200), .A2(n7728), .ZN(n5383) );
  NAND4_X1 U6937 ( .A1(n5386), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(n8578)
         );
  AND2_X1 U6938 ( .A1(n7730), .A2(n8578), .ZN(n5387) );
  INV_X1 U6939 ( .A(n7704), .ZN(n5403) );
  XNOR2_X1 U6940 ( .A(n5388), .B(n10118), .ZN(n5389) );
  XNOR2_X1 U6941 ( .A(n5390), .B(n5389), .ZN(n6950) );
  NAND2_X1 U6942 ( .A1(n6950), .A2(n8329), .ZN(n5396) );
  NAND2_X1 U6943 ( .A1(n5392), .A2(n5391), .ZN(n5393) );
  NAND2_X1 U6944 ( .A1(n5393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U6945 ( .A(n5394), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8642) );
  AOI22_X1 U6946 ( .A1(n5423), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6384), .B2(
        n8642), .ZN(n5395) );
  NAND2_X1 U6947 ( .A1(n5214), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5402) );
  INV_X1 U6948 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7706) );
  OR2_X1 U6949 ( .A1(n8336), .A2(n7706), .ZN(n5401) );
  INV_X1 U6950 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8590) );
  OR2_X1 U6951 ( .A1(n5429), .A2(n8590), .ZN(n5400) );
  NAND2_X1 U6952 ( .A1(n5397), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5398) );
  AND2_X1 U6953 ( .A1(n5413), .A2(n5398), .ZN(n7707) );
  OR2_X1 U6954 ( .A1(n5200), .A2(n7707), .ZN(n5399) );
  NAND4_X1 U6955 ( .A1(n5402), .A2(n5401), .A3(n5400), .A4(n5399), .ZN(n8577)
         );
  NAND2_X1 U6956 ( .A1(n5403), .A2(n4988), .ZN(n5405) );
  NAND2_X1 U6957 ( .A1(n7761), .A2(n8577), .ZN(n5404) );
  XNOR2_X1 U6958 ( .A(n5406), .B(SI_16_), .ZN(n5407) );
  XNOR2_X1 U6959 ( .A(n5408), .B(n5407), .ZN(n6982) );
  NAND2_X1 U6960 ( .A1(n6982), .A2(n8329), .ZN(n5412) );
  OR2_X1 U6961 ( .A1(n5409), .A2(n5133), .ZN(n5410) );
  XNOR2_X1 U6962 ( .A(n5410), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8646) );
  AOI22_X1 U6963 ( .A1(n5423), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6384), .B2(
        n8646), .ZN(n5411) );
  NAND2_X1 U6964 ( .A1(n5214), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5418) );
  INV_X1 U6965 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8645) );
  OR2_X1 U6966 ( .A1(n5429), .A2(n8645), .ZN(n5417) );
  INV_X1 U6967 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7738) );
  OR2_X1 U6968 ( .A1(n8336), .A2(n7738), .ZN(n5416) );
  NAND2_X1 U6969 ( .A1(n5413), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5414) );
  AND2_X1 U6970 ( .A1(n5426), .A2(n5414), .ZN(n7739) );
  OR2_X1 U6971 ( .A1(n5200), .A2(n7739), .ZN(n5415) );
  NAND2_X1 U6972 ( .A1(n8260), .A2(n8269), .ZN(n8470) );
  NAND2_X1 U6973 ( .A1(n8471), .A2(n8470), .ZN(n8368) );
  XNOR2_X1 U6974 ( .A(n5420), .B(n5419), .ZN(n7081) );
  NAND2_X1 U6975 ( .A1(n7081), .A2(n8329), .ZN(n5425) );
  NAND2_X1 U6976 ( .A1(n5421), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5422) );
  XNOR2_X1 U6977 ( .A(n5422), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8648) );
  AOI22_X1 U6978 ( .A1(n5423), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6384), .B2(
        n8648), .ZN(n5424) );
  NAND2_X1 U6979 ( .A1(n5425), .A2(n5424), .ZN(n8951) );
  NAND2_X1 U6980 ( .A1(n5214), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5433) );
  INV_X1 U6981 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8829) );
  OR2_X1 U6982 ( .A1(n8336), .A2(n8829), .ZN(n5432) );
  NAND2_X1 U6983 ( .A1(n5426), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5427) );
  AND2_X1 U6984 ( .A1(n5428), .A2(n5427), .ZN(n8267) );
  OR2_X1 U6985 ( .A1(n5200), .A2(n8267), .ZN(n5431) );
  INV_X1 U6986 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9824) );
  OR2_X1 U6987 ( .A1(n5429), .A2(n9824), .ZN(n5430) );
  OR2_X1 U6988 ( .A1(n8951), .A2(n8307), .ZN(n8811) );
  NAND2_X1 U6989 ( .A1(n8951), .A2(n8307), .ZN(n8475) );
  INV_X1 U6990 ( .A(n8951), .ZN(n8273) );
  OAI22_X1 U6991 ( .A1(n8825), .A2(n8824), .B1(n8307), .B2(n8273), .ZN(n8815)
         );
  NOR2_X1 U6992 ( .A1(n8815), .A2(n5434), .ZN(n5435) );
  AOI21_X1 U6993 ( .B1(n5582), .B2(n8137), .A(n5435), .ZN(n8799) );
  XNOR2_X1 U6994 ( .A(n5437), .B(n10148), .ZN(n5438) );
  XNOR2_X1 U6995 ( .A(n5439), .B(n5438), .ZN(n7347) );
  NAND2_X1 U6996 ( .A1(n7347), .A2(n8329), .ZN(n5441) );
  INV_X1 U6997 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7359) );
  OR2_X1 U6998 ( .A1(n8331), .A2(n7359), .ZN(n5440) );
  NAND2_X1 U6999 ( .A1(n5442), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U7000 ( .A1(n5453), .A2(n5443), .ZN(n8796) );
  AOI22_X1 U7001 ( .A1(n8796), .A2(n5545), .B1(n5214), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5445) );
  AOI22_X1 U7002 ( .A1(n5598), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5193), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n5444) );
  NOR2_X1 U7003 ( .A1(n8937), .A2(n8236), .ZN(n5586) );
  NOR2_X1 U7004 ( .A1(n5586), .A2(n8485), .ZN(n8352) );
  NOR2_X1 U7005 ( .A1(n8937), .A2(n8800), .ZN(n8778) );
  NAND2_X1 U7006 ( .A1(n5447), .A2(n5446), .ZN(n5448) );
  NAND2_X1 U7007 ( .A1(n5449), .A2(n5448), .ZN(n7416) );
  OR2_X1 U7008 ( .A1(n7416), .A2(n5450), .ZN(n5452) );
  INV_X1 U7009 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7414) );
  OR2_X1 U7010 ( .A1(n8331), .A2(n7414), .ZN(n5451) );
  NAND2_X1 U7011 ( .A1(n5453), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U7012 ( .A1(n5466), .A2(n5454), .ZN(n8784) );
  NAND2_X1 U7013 ( .A1(n8784), .A2(n5545), .ZN(n5457) );
  AOI22_X1 U7014 ( .A1(n5598), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5193), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U7015 ( .A1(n5214), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5455) );
  OR2_X1 U7016 ( .A1(n8931), .A2(n5458), .ZN(n5587) );
  NAND2_X1 U7017 ( .A1(n8931), .A2(n5458), .ZN(n8501) );
  NAND2_X1 U7018 ( .A1(n5587), .A2(n8501), .ZN(n8777) );
  NAND2_X1 U7019 ( .A1(n5459), .A2(n5458), .ZN(n5460) );
  XNOR2_X1 U7020 ( .A(n5462), .B(n5461), .ZN(n7592) );
  NAND2_X1 U7021 ( .A1(n7592), .A2(n8329), .ZN(n5465) );
  INV_X1 U7022 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n5463) );
  OR2_X1 U7023 ( .A1(n8331), .A2(n5463), .ZN(n5464) );
  NAND2_X1 U7024 ( .A1(n5466), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U7025 ( .A1(n5476), .A2(n5467), .ZN(n8770) );
  NAND2_X1 U7026 ( .A1(n8770), .A2(n5545), .ZN(n5470) );
  AOI22_X1 U7027 ( .A1(n5598), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n5193), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7028 ( .A1(n5214), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5468) );
  XNOR2_X1 U7029 ( .A(n8925), .B(n8490), .ZN(n8766) );
  XNOR2_X1 U7030 ( .A(n5473), .B(n5472), .ZN(n7629) );
  NAND2_X1 U7031 ( .A1(n7629), .A2(n8329), .ZN(n5475) );
  INV_X1 U7032 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7627) );
  OR2_X1 U7033 ( .A1(n8331), .A2(n7627), .ZN(n5474) );
  NAND2_X1 U7034 ( .A1(n5476), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U7035 ( .A1(n5488), .A2(n5477), .ZN(n8760) );
  NAND2_X1 U7036 ( .A1(n8760), .A2(n5545), .ZN(n5482) );
  INV_X1 U7037 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8918) );
  NAND2_X1 U7038 ( .A1(n5598), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U7039 ( .A1(n5193), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5478) );
  OAI211_X1 U7040 ( .C1(n8918), .C2(n5601), .A(n5479), .B(n5478), .ZN(n5480)
         );
  INV_X1 U7041 ( .A(n5480), .ZN(n5481) );
  XNOR2_X1 U7042 ( .A(n5485), .B(n5484), .ZN(n7718) );
  NAND2_X1 U7043 ( .A1(n7718), .A2(n8329), .ZN(n5487) );
  INV_X1 U7044 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8124) );
  OR2_X1 U7045 ( .A1(n8331), .A2(n8124), .ZN(n5486) );
  NAND2_X1 U7046 ( .A1(n5488), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U7047 ( .A1(n5490), .A2(n5489), .ZN(n8749) );
  NAND2_X1 U7048 ( .A1(n8749), .A2(n5545), .ZN(n5495) );
  INV_X1 U7049 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U7050 ( .A1(n5193), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7051 ( .A1(n5598), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5491) );
  OAI211_X1 U7052 ( .C1(n5601), .C2(n8912), .A(n5492), .B(n5491), .ZN(n5493)
         );
  INV_X1 U7053 ( .A(n5493), .ZN(n5494) );
  NAND2_X1 U7054 ( .A1(n8907), .A2(n8158), .ZN(n8524) );
  NAND2_X1 U7055 ( .A1(n8523), .A2(n8524), .ZN(n8734) );
  NAND2_X1 U7056 ( .A1(n8735), .A2(n8734), .ZN(n8733) );
  NAND2_X1 U7057 ( .A1(n5497), .A2(n5496), .ZN(n5502) );
  INV_X1 U7058 ( .A(n5498), .ZN(n5500) );
  NAND2_X1 U7059 ( .A1(n5500), .A2(n5499), .ZN(n5501) );
  NAND2_X1 U7060 ( .A1(n5502), .A2(n5501), .ZN(n5514) );
  MUX2_X1 U7061 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n4713), .Z(n5515) );
  XNOR2_X1 U7062 ( .A(n5515), .B(n10149), .ZN(n5513) );
  XNOR2_X1 U7063 ( .A(n5514), .B(n5513), .ZN(n7770) );
  NAND2_X1 U7064 ( .A1(n7770), .A2(n8329), .ZN(n5504) );
  INV_X1 U7065 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7771) );
  OR2_X1 U7066 ( .A1(n8331), .A2(n7771), .ZN(n5503) );
  OR2_X2 U7067 ( .A1(n5505), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7068 ( .A1(n5505), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5506) );
  NAND2_X1 U7069 ( .A1(n5523), .A2(n5506), .ZN(n8729) );
  NAND2_X1 U7070 ( .A1(n8729), .A2(n5545), .ZN(n5511) );
  INV_X1 U7071 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U7072 ( .A1(n5598), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U7073 ( .A1(n5193), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5507) );
  OAI211_X1 U7074 ( .C1(n8900), .C2(n5601), .A(n5508), .B(n5507), .ZN(n5509)
         );
  INV_X1 U7075 ( .A(n5509), .ZN(n5510) );
  NAND2_X2 U7076 ( .A1(n5511), .A2(n5510), .ZN(n8736) );
  NAND2_X1 U7077 ( .A1(n8901), .A2(n8736), .ZN(n5512) );
  INV_X1 U7078 ( .A(n8901), .ZN(n8327) );
  NAND2_X1 U7079 ( .A1(n5514), .A2(n5513), .ZN(n5518) );
  INV_X1 U7080 ( .A(n5515), .ZN(n5516) );
  NAND2_X1 U7081 ( .A1(n5516), .A2(n10149), .ZN(n5517) );
  NAND2_X1 U7082 ( .A1(n5518), .A2(n5517), .ZN(n5532) );
  MUX2_X1 U7083 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n4713), .Z(n5533) );
  XNOR2_X1 U7084 ( .A(n5533), .B(n10166), .ZN(n5531) );
  XNOR2_X1 U7085 ( .A(n5532), .B(n5531), .ZN(n8094) );
  NAND2_X1 U7086 ( .A1(n8094), .A2(n8329), .ZN(n5520) );
  INV_X1 U7087 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8201) );
  OR2_X1 U7088 ( .A1(n8331), .A2(n8201), .ZN(n5519) );
  INV_X1 U7089 ( .A(n5523), .ZN(n5522) );
  INV_X1 U7090 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7091 ( .A1(n5522), .A2(n5521), .ZN(n5538) );
  NAND2_X1 U7092 ( .A1(n5523), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7093 ( .A1(n5538), .A2(n5524), .ZN(n8720) );
  NAND2_X1 U7094 ( .A1(n8720), .A2(n5545), .ZN(n5529) );
  INV_X1 U7095 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8894) );
  NAND2_X1 U7096 ( .A1(n5598), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7097 ( .A1(n5193), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5525) );
  OAI211_X1 U7098 ( .C1(n8894), .C2(n5601), .A(n5526), .B(n5525), .ZN(n5527)
         );
  INV_X1 U7099 ( .A(n5527), .ZN(n5528) );
  NAND2_X1 U7100 ( .A1(n8216), .A2(n8702), .ZN(n5530) );
  INV_X1 U7101 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U7102 ( .A1(n5534), .A2(n10166), .ZN(n5535) );
  MUX2_X1 U7103 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n4713), .Z(n5554) );
  INV_X1 U7104 ( .A(SI_28_), .ZN(n5555) );
  XNOR2_X1 U7105 ( .A(n5554), .B(n5555), .ZN(n5552) );
  NAND2_X1 U7106 ( .A1(n8964), .A2(n8329), .ZN(n5537) );
  INV_X1 U7107 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8967) );
  OR2_X1 U7108 ( .A1(n8331), .A2(n8967), .ZN(n5536) );
  NAND2_X1 U7109 ( .A1(n5538), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U7110 ( .A1(n8685), .A2(n5539), .ZN(n8708) );
  NAND2_X1 U7111 ( .A1(n8708), .A2(n5545), .ZN(n5544) );
  INV_X1 U7112 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U7113 ( .A1(n5598), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7114 ( .A1(n5193), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5540) );
  OAI211_X1 U7115 ( .C1(n8887), .C2(n5601), .A(n5541), .B(n5540), .ZN(n5542)
         );
  INV_X1 U7116 ( .A(n5542), .ZN(n5543) );
  INV_X1 U7117 ( .A(n8717), .ZN(n8539) );
  INV_X1 U7118 ( .A(n8685), .ZN(n5546) );
  NAND2_X1 U7119 ( .A1(n5546), .A2(n5545), .ZN(n8342) );
  INV_X1 U7120 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7121 ( .A1(n5193), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7122 ( .A1(n5598), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5547) );
  OAI211_X1 U7123 ( .C1(n5601), .C2(n5549), .A(n5548), .B(n5547), .ZN(n5550)
         );
  INV_X1 U7124 ( .A(n5550), .ZN(n5551) );
  NAND2_X1 U7125 ( .A1(n8342), .A2(n5551), .ZN(n8576) );
  INV_X1 U7126 ( .A(n5554), .ZN(n5556) );
  MUX2_X1 U7127 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4713), .Z(n7902) );
  INV_X1 U7128 ( .A(SI_29_), .ZN(n5557) );
  INV_X1 U7129 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8203) );
  NOR2_X1 U7130 ( .A1(n8331), .A2(n8203), .ZN(n5558) );
  XOR2_X1 U7131 ( .A(n8576), .B(n8697), .Z(n5592) );
  XNOR2_X1 U7132 ( .A(n5559), .B(n5592), .ZN(n5566) );
  NAND2_X1 U7133 ( .A1(n8663), .A2(n8572), .ZN(n5649) );
  NAND2_X1 U7134 ( .A1(n4386), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7135 ( .A1(n5562), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5563) );
  MUX2_X1 U7136 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5563), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5564) );
  NAND2_X1 U7137 ( .A1(n8381), .A2(n6673), .ZN(n5565) );
  NAND2_X2 U7138 ( .A1(n5649), .A2(n5565), .ZN(n9851) );
  INV_X1 U7139 ( .A(n6878), .ZN(n5569) );
  INV_X1 U7140 ( .A(n5567), .ZN(n5568) );
  NAND2_X1 U7141 ( .A1(n5568), .A2(n6577), .ZN(n6571) );
  NAND2_X1 U7142 ( .A1(n6879), .A2(n8384), .ZN(n9858) );
  INV_X1 U7143 ( .A(n8354), .ZN(n9859) );
  NAND2_X1 U7144 ( .A1(n9858), .A2(n9859), .ZN(n5570) );
  XNOR2_X1 U7145 ( .A(n9854), .B(n9883), .ZN(n9840) );
  NAND2_X1 U7146 ( .A1(n9841), .A2(n9840), .ZN(n5571) );
  INV_X1 U7147 ( .A(n9883), .ZN(n8391) );
  OR2_X1 U7148 ( .A1(n9854), .A2(n8391), .ZN(n8399) );
  INV_X1 U7149 ( .A(n8356), .ZN(n8397) );
  INV_X1 U7150 ( .A(n7078), .ZN(n9893) );
  OR2_X1 U7151 ( .A1(n8587), .A2(n9893), .ZN(n7189) );
  NAND2_X1 U7152 ( .A1(n8587), .A2(n9893), .ZN(n8408) );
  AND2_X1 U7153 ( .A1(n7189), .A2(n5572), .ZN(n8411) );
  NAND2_X1 U7154 ( .A1(n7086), .A2(n8411), .ZN(n5573) );
  AND2_X1 U7155 ( .A1(n8418), .A2(n7160), .ZN(n8415) );
  INV_X1 U7156 ( .A(n7286), .ZN(n5575) );
  NAND2_X1 U7157 ( .A1(n5575), .A2(n5574), .ZN(n7284) );
  AND2_X1 U7158 ( .A1(n8438), .A2(n8419), .ZN(n8430) );
  AND2_X1 U7159 ( .A1(n9929), .A2(n7675), .ZN(n8440) );
  OR2_X1 U7160 ( .A1(n9929), .A2(n7675), .ZN(n8439) );
  NAND2_X1 U7161 ( .A1(n5576), .A2(n8439), .ZN(n7543) );
  NAND2_X1 U7162 ( .A1(n7543), .A2(n8445), .ZN(n5577) );
  NAND2_X1 U7163 ( .A1(n5577), .A2(n8447), .ZN(n7540) );
  NOR2_X1 U7164 ( .A1(n8451), .A2(n7722), .ZN(n5579) );
  NAND2_X1 U7165 ( .A1(n8451), .A2(n7722), .ZN(n5578) );
  OAI21_X1 U7166 ( .B1(n7540), .B2(n5579), .A(n5578), .ZN(n7635) );
  OR2_X1 U7167 ( .A1(n7730), .A2(n7756), .ZN(n8460) );
  NAND2_X1 U7168 ( .A1(n7635), .A2(n8460), .ZN(n5580) );
  NAND2_X1 U7169 ( .A1(n7730), .A2(n7756), .ZN(n8461) );
  NAND2_X1 U7170 ( .A1(n5580), .A2(n8461), .ZN(n7703) );
  INV_X1 U7171 ( .A(n8577), .ZN(n8258) );
  OR2_X1 U7172 ( .A1(n7761), .A2(n8258), .ZN(n8466) );
  NAND2_X1 U7173 ( .A1(n7761), .A2(n8258), .ZN(n8465) );
  INV_X1 U7174 ( .A(n8470), .ZN(n5581) );
  AND2_X1 U7175 ( .A1(n5582), .A2(n8827), .ZN(n8476) );
  INV_X1 U7176 ( .A(n8476), .ZN(n5583) );
  AND2_X1 U7177 ( .A1(n5583), .A2(n8811), .ZN(n5584) );
  NAND2_X1 U7178 ( .A1(n8812), .A2(n5584), .ZN(n5585) );
  NAND2_X1 U7179 ( .A1(n8944), .A2(n8137), .ZN(n8479) );
  NAND2_X1 U7180 ( .A1(n5585), .A2(n8479), .ZN(n8804) );
  OR2_X1 U7181 ( .A1(n8867), .A2(n8287), .ZN(n8483) );
  NAND2_X1 U7182 ( .A1(n8867), .A2(n8287), .ZN(n8484) );
  INV_X1 U7183 ( .A(n5586), .ZN(n8773) );
  AND2_X1 U7184 ( .A1(n5587), .A2(n8773), .ZN(n8499) );
  INV_X1 U7185 ( .A(n8501), .ZN(n8488) );
  NAND2_X1 U7186 ( .A1(n8763), .A2(n4727), .ZN(n5588) );
  OR2_X1 U7187 ( .A1(n8925), .A2(n8490), .ZN(n8503) );
  NAND2_X1 U7188 ( .A1(n5588), .A2(n8503), .ZN(n8754) );
  NOR2_X1 U7189 ( .A1(n8919), .A2(n8508), .ZN(n8491) );
  NAND2_X1 U7190 ( .A1(n8919), .A2(n8508), .ZN(n8506) );
  NAND2_X1 U7191 ( .A1(n8913), .A2(n8514), .ZN(n8505) );
  NOR2_X1 U7192 ( .A1(n8913), .A2(n8514), .ZN(n8492) );
  INV_X1 U7193 ( .A(n8524), .ZN(n5590) );
  NOR2_X1 U7194 ( .A1(n8901), .A2(n5591), .ZN(n8528) );
  NAND2_X1 U7195 ( .A1(n8895), .A2(n8702), .ZN(n8531) );
  NAND2_X1 U7196 ( .A1(n8530), .A2(n8531), .ZN(n8713) );
  AOI22_X1 U7197 ( .A1(n8698), .A2(n8700), .B1(n8892), .B2(n8717), .ZN(n8334)
         );
  XNOR2_X1 U7198 ( .A(n8334), .B(n5592), .ZN(n5608) );
  INV_X1 U7199 ( .A(n8572), .ZN(n7596) );
  OAI21_X1 U7200 ( .B1(n8572), .B2(n8566), .A(n9913), .ZN(n5593) );
  NOR2_X1 U7201 ( .A1(n8663), .A2(n5593), .ZN(n5594) );
  OR3_X1 U7202 ( .A1(n8663), .A2(n6673), .A3(n8545), .ZN(n6863) );
  NAND2_X1 U7203 ( .A1(n5608), .A2(n6656), .ZN(n5607) );
  INV_X1 U7204 ( .A(n5595), .ZN(n8568) );
  NAND2_X1 U7205 ( .A1(n8568), .A2(n8664), .ZN(n5597) );
  NAND2_X1 U7206 ( .A1(n5187), .A2(n5597), .ZN(n6676) );
  INV_X1 U7207 ( .A(n6676), .ZN(n6576) );
  INV_X1 U7208 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7209 ( .A1(n5598), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7210 ( .A1(n5193), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5599) );
  OAI211_X1 U7211 ( .C1(n5602), .C2(n5601), .A(n5600), .B(n5599), .ZN(n5603)
         );
  INV_X1 U7212 ( .A(n5603), .ZN(n5604) );
  NAND2_X1 U7213 ( .A1(n8342), .A2(n5604), .ZN(n8575) );
  AND2_X1 U7214 ( .A1(n5187), .A2(P2_B_REG_SCAN_IN), .ZN(n5605) );
  NOR2_X1 U7215 ( .A1(n8703), .A2(n5605), .ZN(n8683) );
  AOI22_X1 U7216 ( .A1(n9855), .A2(n8717), .B1(n8575), .B2(n8683), .ZN(n5606)
         );
  INV_X1 U7217 ( .A(n5608), .ZN(n8692) );
  OR2_X1 U7218 ( .A1(n8562), .A2(n8572), .ZN(n9873) );
  NAND2_X1 U7219 ( .A1(n5628), .A2(n5629), .ZN(n5609) );
  XNOR2_X1 U7220 ( .A(n5619), .B(P2_B_REG_SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7221 ( .A1(n5611), .A2(n5610), .ZN(n5612) );
  NAND2_X1 U7222 ( .A1(n5615), .A2(n5625), .ZN(n5618) );
  NAND2_X1 U7223 ( .A1(n5616), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7224 ( .A1(n5618), .A2(n5620), .ZN(n5624) );
  NAND2_X1 U7225 ( .A1(n5619), .A2(n7772), .ZN(n6415) );
  NAND2_X1 U7226 ( .A1(n5621), .A2(n6415), .ZN(n5622) );
  NOR2_X1 U7227 ( .A1(n9873), .A2(n8381), .ZN(n6574) );
  INV_X1 U7228 ( .A(n8663), .ZN(n8673) );
  NAND3_X1 U7229 ( .A1(n8673), .A2(n8572), .A3(n6673), .ZN(n5623) );
  AND2_X1 U7230 ( .A1(n5623), .A2(n8545), .ZN(n6867) );
  OAI21_X1 U7231 ( .B1(n5622), .B2(n6574), .A(n6867), .ZN(n5643) );
  OR2_X1 U7232 ( .A1(n5624), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U7233 ( .A1(n5625), .A2(n7772), .ZN(n6412) );
  NAND2_X1 U7234 ( .A1(n8673), .A2(n8566), .ZN(n8560) );
  NAND2_X1 U7235 ( .A1(n8560), .A2(n8554), .ZN(n5627) );
  NAND2_X1 U7236 ( .A1(n5627), .A2(n6382), .ZN(n6579) );
  NOR2_X1 U7237 ( .A1(n6579), .A2(n6380), .ZN(n5641) );
  NOR2_X1 U7238 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n5633) );
  NOR4_X1 U7239 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5632) );
  NOR4_X1 U7240 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5631) );
  NOR4_X1 U7241 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n5630) );
  NAND4_X1 U7242 ( .A1(n5633), .A2(n5632), .A3(n5631), .A4(n5630), .ZN(n5639)
         );
  NOR4_X1 U7243 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5637) );
  NOR4_X1 U7244 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n5636) );
  NOR4_X1 U7245 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5635) );
  NOR4_X1 U7246 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5634) );
  NAND4_X1 U7247 ( .A1(n5637), .A2(n5636), .A3(n5635), .A4(n5634), .ZN(n5638)
         );
  NOR2_X1 U7248 ( .A1(n5639), .A2(n5638), .ZN(n5640) );
  OR2_X1 U7249 ( .A1(n5624), .A2(n5640), .ZN(n5651) );
  AND2_X1 U7250 ( .A1(n5641), .A2(n5651), .ZN(n6872) );
  NAND2_X1 U7251 ( .A1(n6868), .A2(n6866), .ZN(n5642) );
  NAND2_X1 U7252 ( .A1(n9947), .A2(n9930), .ZN(n8842) );
  NAND2_X1 U7253 ( .A1(n9945), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7254 ( .A1(n5646), .A2(n5645), .ZN(P2_U3488) );
  INV_X1 U7255 ( .A(n5651), .ZN(n5647) );
  OR2_X1 U7256 ( .A1(n5648), .A2(n5647), .ZN(n6583) );
  NAND2_X1 U7257 ( .A1(n6578), .A2(n6863), .ZN(n5650) );
  NAND2_X1 U7258 ( .A1(n6572), .A2(n5650), .ZN(n5654) );
  NAND3_X1 U7259 ( .A1(n5622), .A2(n6868), .A3(n5651), .ZN(n6845) );
  AND2_X1 U7260 ( .A1(n8545), .A2(n9913), .ZN(n5652) );
  NAND2_X1 U7261 ( .A1(n6578), .A2(n5652), .ZN(n6567) );
  AND2_X1 U7262 ( .A1(n6567), .A2(n8742), .ZN(n6581) );
  NAND2_X1 U7263 ( .A1(n5655), .A2(n9931), .ZN(n5658) );
  OR2_X1 U7264 ( .A1(n9933), .A2(n9913), .ZN(n8891) );
  OR2_X1 U7265 ( .A1(n9931), .A2(n5549), .ZN(n5656) );
  NAND2_X1 U7266 ( .A1(n5658), .A2(n5657), .ZN(P2_U3456) );
  INV_X4 U7267 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U7268 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5763) );
  NOR2_X2 U7269 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5799) );
  NOR2_X1 U7270 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5659) );
  NOR2_X2 U7271 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5704) );
  INV_X1 U7272 ( .A(n5668), .ZN(n5667) );
  NAND2_X2 U7273 ( .A1(n5709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U7274 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n5669) );
  NAND2_X1 U7275 ( .A1(n5702), .A2(n5669), .ZN(n5670) );
  NAND2_X1 U7276 ( .A1(n6563), .A2(n7912), .ZN(n5675) );
  NOR2_X1 U7277 ( .A1(n5854), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5869) );
  NOR2_X1 U7278 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5672) );
  NAND2_X1 U7279 ( .A1(n5869), .A2(n5672), .ZN(n5909) );
  NAND2_X1 U7280 ( .A1(n5938), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5673) );
  XNOR2_X1 U7281 ( .A(n5673), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6782) );
  AOI22_X1 U7282 ( .A1(n6082), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6081), .B2(
        n6782), .ZN(n5674) );
  NAND2_X1 U7283 ( .A1(n6044), .A2(n5685), .ZN(n6061) );
  NAND2_X1 U7284 ( .A1(n6061), .A2(n5686), .ZN(n5691) );
  NAND2_X1 U7285 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n5687) );
  INV_X1 U7286 ( .A(n6061), .ZN(n5693) );
  MUX2_X1 U7287 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5698), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5700) );
  NAND2_X1 U7288 ( .A1(n6250), .A2(n6247), .ZN(n5708) );
  INV_X1 U7289 ( .A(n5704), .ZN(n5705) );
  INV_X2 U7290 ( .A(n8063), .ZN(n8108) );
  NAND2_X1 U7291 ( .A1(n7292), .A2(n8184), .ZN(n5724) );
  XNOR2_X2 U7292 ( .A(n5710), .B(n9525), .ZN(n9534) );
  NAND2_X1 U7293 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5711) );
  NAND2_X1 U7294 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  XNOR2_X2 U7295 ( .A(n5713), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5716) );
  BUF_X2 U7296 ( .A(n5716), .Z(n8199) );
  BUF_X4 U7297 ( .A(n5740), .Z(n6334) );
  AND2_X1 U7298 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5794) );
  NAND2_X1 U7299 ( .A1(n5794), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5830) );
  INV_X1 U7300 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5829) );
  NOR2_X1 U7301 ( .A1(n5830), .A2(n5829), .ZN(n5828) );
  NAND2_X1 U7302 ( .A1(n5828), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5873) );
  NOR2_X1 U7303 ( .A1(n5891), .A2(n6509), .ZN(n5890) );
  NAND2_X1 U7304 ( .A1(n5714), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5942) );
  INV_X1 U7305 ( .A(n5714), .ZN(n5916) );
  INV_X1 U7306 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6553) );
  NAND2_X1 U7307 ( .A1(n5916), .A2(n6553), .ZN(n5715) );
  AND2_X1 U7308 ( .A1(n5942), .A2(n5715), .ZN(n7299) );
  NAND2_X1 U7309 ( .A1(n6334), .A2(n7299), .ZN(n5721) );
  INV_X2 U7310 ( .A(n5860), .ZN(n6220) );
  NAND2_X1 U7311 ( .A1(n6433), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5720) );
  NAND2_X1 U7312 ( .A1(n6435), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5719) );
  NAND2_X1 U7313 ( .A1(n6434), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5718) );
  NAND4_X1 U7314 ( .A1(n5721), .A2(n5720), .A3(n5719), .A4(n5718), .ZN(n9669)
         );
  NAND2_X1 U7315 ( .A1(n9669), .A2(n6174), .ZN(n5723) );
  NAND2_X1 U7316 ( .A1(n5724), .A2(n5723), .ZN(n5725) );
  XNOR2_X1 U7317 ( .A(n5725), .B(n4356), .ZN(n5924) );
  INV_X2 U7318 ( .A(n6213), .ZN(n8179) );
  AND2_X1 U7319 ( .A1(n9669), .A2(n8179), .ZN(n5727) );
  AOI21_X1 U7320 ( .B1(n7292), .B2(n4355), .A(n5727), .ZN(n5925) );
  NAND2_X1 U7321 ( .A1(n5924), .A2(n5925), .ZN(n7482) );
  INV_X2 U7322 ( .A(n5734), .ZN(n8178) );
  NAND2_X1 U7323 ( .A1(n9599), .A2(n8178), .ZN(n5732) );
  INV_X1 U7324 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U7325 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5728) );
  XNOR2_X1 U7326 ( .A(n5729), .B(n5728), .ZN(n6459) );
  INV_X1 U7327 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6404) );
  OR2_X1 U7328 ( .A1(n5784), .A2(n6404), .ZN(n5730) );
  NAND2_X1 U7329 ( .A1(n7792), .A2(n6161), .ZN(n5731) );
  NAND2_X1 U7330 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  XNOR2_X1 U7331 ( .A(n5733), .B(n4356), .ZN(n5739) );
  INV_X1 U7332 ( .A(n5739), .ZN(n5737) );
  AND2_X1 U7333 ( .A1(n7792), .A2(n5726), .ZN(n5735) );
  INV_X1 U7334 ( .A(n5738), .ZN(n5736) );
  BUF_X1 U7335 ( .A(n5740), .Z(n6285) );
  NAND2_X1 U7336 ( .A1(n6285), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U7337 ( .A1(n5860), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7338 ( .A1(n5758), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5742) );
  NAND2_X1 U7339 ( .A1(n9127), .A2(n8178), .ZN(n5751) );
  INV_X1 U7340 ( .A(SI_0_), .ZN(n5747) );
  INV_X1 U7341 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5746) );
  OAI21_X1 U7342 ( .B1(n7917), .B2(n5747), .A(n5746), .ZN(n5749) );
  AND2_X1 U7343 ( .A1(n5749), .A2(n5748), .ZN(n9538) );
  MUX2_X1 U7344 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9538), .S(n7923), .Z(n6745) );
  NAND2_X1 U7345 ( .A1(n6745), .A2(n6161), .ZN(n5750) );
  NAND2_X1 U7346 ( .A1(n5751), .A2(n5750), .ZN(n5755) );
  INV_X1 U7347 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6426) );
  NOR2_X1 U7348 ( .A1(n6273), .A2(n6426), .ZN(n5752) );
  OR2_X1 U7349 ( .A1(n5755), .A2(n5752), .ZN(n6519) );
  NAND2_X1 U7350 ( .A1(n9127), .A2(n8179), .ZN(n5754) );
  INV_X1 U7351 ( .A(n6273), .ZN(n6378) );
  AOI22_X1 U7352 ( .A1(n6745), .A2(n8178), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6378), .ZN(n5753) );
  NAND2_X1 U7353 ( .A1(n5754), .A2(n5753), .ZN(n6520) );
  OR2_X1 U7354 ( .A1(n5755), .A2(n8182), .ZN(n5756) );
  NAND2_X1 U7355 ( .A1(n7789), .A2(n5757), .ZN(n9078) );
  NAND2_X1 U7356 ( .A1(n6285), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5762) );
  NAND2_X1 U7357 ( .A1(n5860), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U7358 ( .A1(n5741), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U7359 ( .A1(n9125), .A2(n8178), .ZN(n5768) );
  OR2_X1 U7360 ( .A1(n5763), .A2(n9527), .ZN(n5801) );
  INV_X1 U7361 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U7362 ( .A1(n5801), .A2(n5764), .ZN(n5781) );
  OAI21_X1 U7363 ( .B1(n5801), .B2(n5764), .A(n5781), .ZN(n9151) );
  OR2_X1 U7364 ( .A1(n5765), .A2(n6401), .ZN(n5767) );
  INV_X1 U7365 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6402) );
  OR2_X1 U7366 ( .A1(n5784), .A2(n6402), .ZN(n5766) );
  BUF_X4 U7367 ( .A(n6161), .Z(n8184) );
  AND2_X1 U7368 ( .A1(n9083), .A2(n6174), .ZN(n5769) );
  AOI21_X1 U7369 ( .B1(n9125), .B2(n8179), .A(n5769), .ZN(n5771) );
  INV_X1 U7370 ( .A(n5771), .ZN(n5772) );
  NAND2_X1 U7371 ( .A1(n5773), .A2(n5772), .ZN(n5774) );
  INV_X1 U7372 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6792) );
  NAND2_X1 U7373 ( .A1(n6334), .A2(n6792), .ZN(n5780) );
  INV_X1 U7374 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U7375 ( .A1(n5741), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5778) );
  NAND2_X1 U7376 ( .A1(n6072), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7377 ( .A1(n9598), .A2(n8178), .ZN(n5787) );
  NAND2_X1 U7378 ( .A1(n5781), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5783) );
  INV_X1 U7379 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5782) );
  XNOR2_X1 U7380 ( .A(n5783), .B(n5782), .ZN(n9159) );
  OR2_X1 U7381 ( .A1(n5765), .A2(n6387), .ZN(n5785) );
  INV_X1 U7382 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U7383 ( .A1(n9609), .A2(n8184), .ZN(n5786) );
  NAND2_X1 U7384 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  XNOR2_X1 U7385 ( .A(n5788), .B(n8182), .ZN(n5790) );
  AND2_X1 U7386 ( .A1(n9609), .A2(n4355), .ZN(n5789) );
  AOI21_X1 U7387 ( .B1(n9598), .B2(n8179), .A(n5789), .ZN(n5791) );
  XNOR2_X1 U7388 ( .A(n5790), .B(n5791), .ZN(n6791) );
  INV_X1 U7389 ( .A(n5790), .ZN(n5792) );
  NAND2_X1 U7390 ( .A1(n5792), .A2(n5791), .ZN(n5793) );
  INV_X1 U7391 ( .A(n5794), .ZN(n5812) );
  OAI21_X1 U7392 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5812), .ZN(n6958) );
  NAND2_X1 U7393 ( .A1(n5860), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5797) );
  NAND2_X1 U7394 ( .A1(n6072), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7395 ( .A1(n5741), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7396 ( .A1(n9124), .A2(n8178), .ZN(n5805) );
  OR2_X1 U7397 ( .A1(n5799), .A2(n9527), .ZN(n5800) );
  NAND2_X1 U7398 ( .A1(n5801), .A2(n5800), .ZN(n5808) );
  XNOR2_X1 U7399 ( .A(n5808), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9178) );
  OR2_X1 U7400 ( .A1(n6390), .A2(n5765), .ZN(n5803) );
  INV_X1 U7401 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6391) );
  OR2_X1 U7402 ( .A1(n5784), .A2(n6391), .ZN(n5802) );
  OAI211_X1 U7403 ( .C1(n9178), .C2(n7923), .A(n5803), .B(n5802), .ZN(n9616)
         );
  NAND2_X1 U7404 ( .A1(n9616), .A2(n6161), .ZN(n5804) );
  NAND2_X1 U7405 ( .A1(n5805), .A2(n5804), .ZN(n5806) );
  XNOR2_X1 U7406 ( .A(n5806), .B(n4356), .ZN(n5841) );
  AND2_X1 U7407 ( .A1(n9616), .A2(n4355), .ZN(n5807) );
  AOI21_X1 U7408 ( .B1(n9124), .B2(n8179), .A(n5807), .ZN(n5842) );
  XNOR2_X1 U7409 ( .A(n5841), .B(n5842), .ZN(n6957) );
  OAI21_X1 U7410 ( .B1(n5808), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5809) );
  XNOR2_X1 U7411 ( .A(n5809), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6468) );
  AOI22_X1 U7412 ( .A1(n6082), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6081), .B2(
        n6468), .ZN(n5810) );
  NAND2_X1 U7413 ( .A1(n6976), .A2(n8184), .ZN(n5819) );
  INV_X1 U7414 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7415 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  AND2_X1 U7416 ( .A1(n5830), .A2(n5813), .ZN(n6975) );
  NAND2_X1 U7417 ( .A1(n6334), .A2(n6975), .ZN(n5817) );
  NAND2_X1 U7418 ( .A1(n5860), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U7419 ( .A1(n5741), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7420 ( .A1(n6072), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5814) );
  NAND4_X1 U7421 ( .A1(n5817), .A2(n5816), .A3(n5815), .A4(n5814), .ZN(n9617)
         );
  NAND2_X1 U7422 ( .A1(n9617), .A2(n6174), .ZN(n5818) );
  NAND2_X1 U7423 ( .A1(n5819), .A2(n5818), .ZN(n5820) );
  NAND2_X1 U7424 ( .A1(n9617), .A2(n8179), .ZN(n5822) );
  NAND2_X1 U7425 ( .A1(n6976), .A2(n6174), .ZN(n5821) );
  AND2_X1 U7426 ( .A1(n5822), .A2(n5821), .ZN(n5845) );
  AND2_X1 U7427 ( .A1(n6892), .A2(n5845), .ZN(n5848) );
  OR2_X1 U7428 ( .A1(n6396), .A2(n5765), .ZN(n5827) );
  NAND2_X1 U7429 ( .A1(n5823), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5824) );
  MUX2_X1 U7430 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5824), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5825) );
  AND2_X1 U7431 ( .A1(n5825), .A2(n5854), .ZN(n9216) );
  AOI22_X1 U7432 ( .A1(n6082), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6081), .B2(
        n9216), .ZN(n5826) );
  NAND2_X1 U7433 ( .A1(n5827), .A2(n5826), .ZN(n9577) );
  NAND2_X1 U7434 ( .A1(n9577), .A2(n8184), .ZN(n5837) );
  INV_X1 U7435 ( .A(n5828), .ZN(n5858) );
  NAND2_X1 U7436 ( .A1(n5830), .A2(n5829), .ZN(n5831) );
  AND2_X1 U7437 ( .A1(n5858), .A2(n5831), .ZN(n9572) );
  NAND2_X1 U7438 ( .A1(n6334), .A2(n9572), .ZN(n5835) );
  NAND2_X1 U7439 ( .A1(n6433), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7440 ( .A1(n6435), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7441 ( .A1(n5741), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7442 ( .A1(n9639), .A2(n6174), .ZN(n5836) );
  NAND2_X1 U7443 ( .A1(n5837), .A2(n5836), .ZN(n5838) );
  XNOR2_X1 U7444 ( .A(n5838), .B(n4356), .ZN(n5850) );
  NAND2_X1 U7445 ( .A1(n9577), .A2(n6174), .ZN(n5840) );
  NAND2_X1 U7446 ( .A1(n9639), .A2(n8179), .ZN(n5839) );
  AND2_X1 U7447 ( .A1(n5840), .A2(n5839), .ZN(n5851) );
  NAND2_X1 U7448 ( .A1(n5850), .A2(n5851), .ZN(n6910) );
  INV_X1 U7449 ( .A(n6910), .ZN(n5849) );
  INV_X1 U7450 ( .A(n5841), .ZN(n5844) );
  INV_X1 U7451 ( .A(n5842), .ZN(n5843) );
  NAND2_X1 U7452 ( .A1(n5844), .A2(n5843), .ZN(n6890) );
  INV_X1 U7453 ( .A(n6892), .ZN(n5846) );
  INV_X1 U7454 ( .A(n5845), .ZN(n6891) );
  NAND2_X1 U7455 ( .A1(n5846), .A2(n6891), .ZN(n5847) );
  INV_X1 U7456 ( .A(n5850), .ZN(n5853) );
  INV_X1 U7457 ( .A(n5851), .ZN(n5852) );
  NAND2_X1 U7458 ( .A1(n5853), .A2(n5852), .ZN(n6911) );
  NAND2_X1 U7459 ( .A1(n5854), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5855) );
  XNOR2_X1 U7460 ( .A(n5855), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6473) );
  AOI22_X1 U7461 ( .A1(n6082), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6081), .B2(
        n6473), .ZN(n5856) );
  NAND2_X1 U7462 ( .A1(n4352), .A2(n6174), .ZN(n5865) );
  INV_X1 U7463 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5857) );
  NAND2_X1 U7464 ( .A1(n5858), .A2(n5857), .ZN(n5859) );
  AND2_X1 U7465 ( .A1(n5873), .A2(n5859), .ZN(n7064) );
  NAND2_X1 U7466 ( .A1(n5860), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7467 ( .A1(n6435), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7468 ( .A1(n6434), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7469 ( .A1(n9569), .A2(n8179), .ZN(n5864) );
  NAND2_X1 U7470 ( .A1(n5865), .A2(n5864), .ZN(n6902) );
  NAND2_X1 U7471 ( .A1(n9638), .A2(n6161), .ZN(n5867) );
  NAND2_X1 U7472 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  XNOR2_X1 U7473 ( .A(n5868), .B(n8182), .ZN(n6901) );
  NAND2_X1 U7474 ( .A1(n6430), .A2(n7912), .ZN(n5871) );
  OR2_X1 U7475 ( .A1(n5869), .A2(n9527), .ZN(n5885) );
  XNOR2_X1 U7476 ( .A(n5885), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6504) );
  AOI22_X1 U7477 ( .A1(n6082), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6081), .B2(
        n6504), .ZN(n5870) );
  NAND2_X1 U7478 ( .A1(n6310), .A2(n8184), .ZN(n5880) );
  NAND2_X1 U7479 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  AND2_X1 U7480 ( .A1(n5891), .A2(n5874), .ZN(n9557) );
  NAND2_X1 U7481 ( .A1(n6334), .A2(n9557), .ZN(n5878) );
  NAND2_X1 U7482 ( .A1(n6433), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7483 ( .A1(n6434), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5876) );
  NAND2_X1 U7484 ( .A1(n6435), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U7485 ( .A1(n9658), .A2(n4355), .ZN(n5879) );
  NAND2_X1 U7486 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  XNOR2_X1 U7487 ( .A(n5881), .B(n4356), .ZN(n7129) );
  NAND2_X1 U7488 ( .A1(n6310), .A2(n6174), .ZN(n5883) );
  NAND2_X1 U7489 ( .A1(n9658), .A2(n8179), .ZN(n5882) );
  AND2_X1 U7490 ( .A1(n5883), .A2(n5882), .ZN(n5901) );
  INV_X1 U7491 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5884) );
  NAND2_X1 U7492 ( .A1(n5885), .A2(n5884), .ZN(n5886) );
  NAND2_X1 U7493 ( .A1(n5886), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5887) );
  XNOR2_X1 U7494 ( .A(n5887), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6532) );
  AOI22_X1 U7495 ( .A1(n6082), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6081), .B2(
        n6532), .ZN(n5888) );
  NAND2_X1 U7496 ( .A1(n9660), .A2(n8184), .ZN(n5898) );
  INV_X1 U7497 ( .A(n5890), .ZN(n5914) );
  NAND2_X1 U7498 ( .A1(n5891), .A2(n6509), .ZN(n5892) );
  AND2_X1 U7499 ( .A1(n5914), .A2(n5892), .ZN(n9048) );
  NAND2_X1 U7500 ( .A1(n6334), .A2(n9048), .ZN(n5896) );
  NAND2_X1 U7501 ( .A1(n6433), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U7502 ( .A1(n6435), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7503 ( .A1(n6434), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5893) );
  NAND4_X1 U7504 ( .A1(n5896), .A2(n5895), .A3(n5894), .A4(n5893), .ZN(n9553)
         );
  NAND2_X1 U7505 ( .A1(n9553), .A2(n4355), .ZN(n5897) );
  NAND2_X1 U7506 ( .A1(n5898), .A2(n5897), .ZN(n5899) );
  XNOR2_X1 U7507 ( .A(n5899), .B(n8182), .ZN(n5905) );
  AND2_X1 U7508 ( .A1(n9553), .A2(n8179), .ZN(n5900) );
  AOI21_X1 U7509 ( .B1(n9660), .B2(n4355), .A(n5900), .ZN(n5906) );
  XNOR2_X1 U7510 ( .A(n5905), .B(n5906), .ZN(n9042) );
  INV_X1 U7511 ( .A(n7129), .ZN(n5902) );
  INV_X1 U7512 ( .A(n5901), .ZN(n7131) );
  NAND2_X1 U7513 ( .A1(n5902), .A2(n7131), .ZN(n5903) );
  AND2_X1 U7514 ( .A1(n9042), .A2(n5903), .ZN(n5904) );
  INV_X1 U7515 ( .A(n5905), .ZN(n5907) );
  NAND2_X1 U7516 ( .A1(n5907), .A2(n5906), .ZN(n5908) );
  NAND2_X1 U7517 ( .A1(n6524), .A2(n7912), .ZN(n5912) );
  NAND2_X1 U7518 ( .A1(n5909), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5910) );
  XNOR2_X1 U7519 ( .A(n5910), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6547) );
  AOI22_X1 U7520 ( .A1(n6082), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6081), .B2(
        n6547), .ZN(n5911) );
  NAND2_X1 U7521 ( .A1(n9670), .A2(n8184), .ZN(n5922) );
  INV_X1 U7522 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7523 ( .A1(n5914), .A2(n5913), .ZN(n5915) );
  AND2_X1 U7524 ( .A1(n5916), .A2(n5915), .ZN(n7239) );
  NAND2_X1 U7525 ( .A1(n6334), .A2(n7239), .ZN(n5920) );
  NAND2_X1 U7526 ( .A1(n6433), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7527 ( .A1(n6434), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7528 ( .A1(n6435), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5917) );
  NAND4_X1 U7529 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(n9123)
         );
  NAND2_X1 U7530 ( .A1(n9123), .A2(n4355), .ZN(n5921) );
  NAND2_X1 U7531 ( .A1(n5922), .A2(n5921), .ZN(n5923) );
  XNOR2_X1 U7532 ( .A(n5923), .B(n4356), .ZN(n5930) );
  INV_X1 U7533 ( .A(n5924), .ZN(n5927) );
  INV_X1 U7534 ( .A(n5925), .ZN(n5926) );
  NAND2_X1 U7535 ( .A1(n5927), .A2(n5926), .ZN(n5928) );
  AND2_X1 U7536 ( .A1(n7482), .A2(n5928), .ZN(n7293) );
  INV_X1 U7537 ( .A(n5929), .ZN(n5932) );
  INV_X1 U7538 ( .A(n5930), .ZN(n5931) );
  NAND2_X1 U7539 ( .A1(n5932), .A2(n5931), .ZN(n5934) );
  NAND2_X1 U7540 ( .A1(n9670), .A2(n6174), .ZN(n5936) );
  NAND2_X1 U7541 ( .A1(n9123), .A2(n8179), .ZN(n5935) );
  NAND2_X1 U7542 ( .A1(n5936), .A2(n5935), .ZN(n7238) );
  INV_X1 U7543 ( .A(n7293), .ZN(n5937) );
  NOR2_X1 U7544 ( .A1(n5938), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5981) );
  OR2_X1 U7545 ( .A1(n5981), .A2(n9527), .ZN(n5959) );
  XNOR2_X1 U7546 ( .A(n5959), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6808) );
  AOI22_X1 U7547 ( .A1(n6082), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6081), .B2(
        n6808), .ZN(n5939) );
  NAND2_X1 U7548 ( .A1(n9687), .A2(n8184), .ZN(n5949) );
  NAND2_X1 U7549 ( .A1(n5942), .A2(n5941), .ZN(n5943) );
  AND2_X1 U7550 ( .A1(n5965), .A2(n5943), .ZN(n7475) );
  NAND2_X1 U7551 ( .A1(n6334), .A2(n7475), .ZN(n5947) );
  NAND2_X1 U7552 ( .A1(n6433), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5946) );
  NAND2_X1 U7553 ( .A1(n6434), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7554 ( .A1(n6435), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5944) );
  NAND4_X1 U7555 ( .A1(n5947), .A2(n5946), .A3(n5945), .A4(n5944), .ZN(n9122)
         );
  NAND2_X1 U7556 ( .A1(n9122), .A2(n4355), .ZN(n5948) );
  NAND2_X1 U7557 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  XNOR2_X1 U7558 ( .A(n5950), .B(n4356), .ZN(n5952) );
  AND2_X1 U7559 ( .A1(n9122), .A2(n8179), .ZN(n5951) );
  AOI21_X1 U7560 ( .B1(n9687), .B2(n4355), .A(n5951), .ZN(n5953) );
  NAND2_X1 U7561 ( .A1(n5952), .A2(n5953), .ZN(n5958) );
  INV_X1 U7562 ( .A(n5952), .ZN(n5955) );
  INV_X1 U7563 ( .A(n5953), .ZN(n5954) );
  NAND2_X1 U7564 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  AND2_X1 U7565 ( .A1(n5958), .A2(n5956), .ZN(n7480) );
  NAND2_X1 U7566 ( .A1(n7485), .A2(n5958), .ZN(n7402) );
  NAND2_X1 U7567 ( .A1(n6682), .A2(n7912), .ZN(n5963) );
  INV_X1 U7568 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U7569 ( .A1(n5959), .A2(n5979), .ZN(n5960) );
  NAND2_X1 U7570 ( .A1(n5960), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5961) );
  XNOR2_X1 U7571 ( .A(n5961), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7003) );
  AOI22_X1 U7572 ( .A1(n6082), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6081), .B2(
        n7003), .ZN(n5962) );
  NAND2_X1 U7573 ( .A1(n9696), .A2(n8184), .ZN(n5972) );
  NAND2_X1 U7574 ( .A1(n5965), .A2(n5964), .ZN(n5966) );
  AND2_X1 U7575 ( .A1(n5987), .A2(n5966), .ZN(n7406) );
  NAND2_X1 U7576 ( .A1(n6334), .A2(n7406), .ZN(n5970) );
  NAND2_X1 U7577 ( .A1(n6433), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7578 ( .A1(n6435), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7579 ( .A1(n6434), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5967) );
  NAND4_X1 U7580 ( .A1(n5970), .A2(n5969), .A3(n5968), .A4(n5967), .ZN(n9686)
         );
  NAND2_X1 U7581 ( .A1(n9686), .A2(n4355), .ZN(n5971) );
  NAND2_X1 U7582 ( .A1(n5972), .A2(n5971), .ZN(n5973) );
  XNOR2_X1 U7583 ( .A(n5973), .B(n8182), .ZN(n5975) );
  AND2_X1 U7584 ( .A1(n9686), .A2(n8179), .ZN(n5974) );
  AOI21_X1 U7585 ( .B1(n9696), .B2(n4355), .A(n5974), .ZN(n5976) );
  XNOR2_X1 U7586 ( .A(n5975), .B(n5976), .ZN(n7404) );
  NAND2_X1 U7587 ( .A1(n7402), .A2(n7404), .ZN(n7403) );
  INV_X1 U7588 ( .A(n5975), .ZN(n5977) );
  NAND2_X1 U7589 ( .A1(n5977), .A2(n5976), .ZN(n5978) );
  NAND2_X1 U7590 ( .A1(n7403), .A2(n5978), .ZN(n5997) );
  NAND2_X1 U7591 ( .A1(n6859), .A2(n7912), .ZN(n5985) );
  INV_X1 U7592 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5980) );
  NAND3_X1 U7593 ( .A1(n5981), .A2(n5980), .A3(n5979), .ZN(n5982) );
  NAND2_X1 U7594 ( .A1(n5982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7595 ( .A(n5983), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7139) );
  AOI22_X1 U7596 ( .A1(n6082), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6081), .B2(
        n7139), .ZN(n5984) );
  NAND2_X1 U7597 ( .A1(n9709), .A2(n8184), .ZN(n5994) );
  INV_X1 U7598 ( .A(n6009), .ZN(n6011) );
  NAND2_X1 U7599 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  AND2_X1 U7600 ( .A1(n6011), .A2(n5988), .ZN(n7780) );
  NAND2_X1 U7601 ( .A1(n6334), .A2(n7780), .ZN(n5992) );
  NAND2_X1 U7602 ( .A1(n6433), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5991) );
  NAND2_X1 U7603 ( .A1(n6434), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7604 ( .A1(n6435), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5989) );
  NAND4_X1 U7605 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n9694)
         );
  NAND2_X1 U7606 ( .A1(n9694), .A2(n4355), .ZN(n5993) );
  NAND2_X1 U7607 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  XNOR2_X1 U7608 ( .A(n5995), .B(n4356), .ZN(n5996) );
  NAND2_X1 U7609 ( .A1(n9709), .A2(n4355), .ZN(n6000) );
  NAND2_X1 U7610 ( .A1(n9694), .A2(n8179), .ZN(n5999) );
  NAND2_X1 U7611 ( .A1(n6000), .A2(n5999), .ZN(n7779) );
  NAND2_X1 U7612 ( .A1(n6950), .A2(n7912), .ZN(n6008) );
  INV_X1 U7613 ( .A(n6003), .ZN(n6004) );
  NAND2_X1 U7614 ( .A1(n6004), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6005) );
  MUX2_X1 U7615 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6005), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n6006) );
  AOI22_X1 U7616 ( .A1(n6082), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6081), .B2(
        n7382), .ZN(n6007) );
  NAND2_X1 U7617 ( .A1(n7609), .A2(n8184), .ZN(n6018) );
  NAND2_X1 U7618 ( .A1(n6009), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6028) );
  INV_X1 U7619 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7620 ( .A1(n6011), .A2(n6010), .ZN(n6012) );
  AND2_X1 U7621 ( .A1(n6028), .A2(n6012), .ZN(n7604) );
  NAND2_X1 U7622 ( .A1(n6334), .A2(n7604), .ZN(n6016) );
  NAND2_X1 U7623 ( .A1(n6433), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7624 ( .A1(n6435), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7625 ( .A1(n6434), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6013) );
  NAND4_X1 U7626 ( .A1(n6016), .A2(n6015), .A3(n6014), .A4(n6013), .ZN(n9121)
         );
  NAND2_X1 U7627 ( .A1(n9121), .A2(n6174), .ZN(n6017) );
  NAND2_X1 U7628 ( .A1(n6018), .A2(n6017), .ZN(n6019) );
  XNOR2_X1 U7629 ( .A(n6019), .B(n4356), .ZN(n6020) );
  INV_X1 U7630 ( .A(n6020), .ZN(n6021) );
  AND2_X1 U7631 ( .A1(n9121), .A2(n8179), .ZN(n6022) );
  AOI21_X1 U7632 ( .B1(n7609), .B2(n4355), .A(n6022), .ZN(n9108) );
  NAND2_X1 U7633 ( .A1(n6982), .A2(n7912), .ZN(n6026) );
  XNOR2_X1 U7634 ( .A(n6024), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7398) );
  AOI22_X1 U7635 ( .A1(n6082), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6081), .B2(
        n7398), .ZN(n6025) );
  NAND2_X1 U7636 ( .A1(n9507), .A2(n8184), .ZN(n6035) );
  NAND2_X1 U7637 ( .A1(n6028), .A2(n6027), .ZN(n6029) );
  AND2_X1 U7638 ( .A1(n6048), .A2(n6029), .ZN(n9015) );
  NAND2_X1 U7639 ( .A1(n6285), .A2(n9015), .ZN(n6033) );
  NAND2_X1 U7640 ( .A1(n6433), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6032) );
  NAND2_X1 U7641 ( .A1(n6434), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7642 ( .A1(n6435), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6030) );
  NAND4_X1 U7643 ( .A1(n6033), .A2(n6032), .A3(n6031), .A4(n6030), .ZN(n9539)
         );
  NAND2_X1 U7644 ( .A1(n9539), .A2(n6174), .ZN(n6034) );
  NAND2_X1 U7645 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  XNOR2_X1 U7646 ( .A(n6036), .B(n4356), .ZN(n6038) );
  AND2_X1 U7647 ( .A1(n9539), .A2(n8179), .ZN(n6037) );
  AOI21_X1 U7648 ( .B1(n9507), .B2(n4355), .A(n6037), .ZN(n6039) );
  NAND2_X1 U7649 ( .A1(n6038), .A2(n6039), .ZN(n6043) );
  INV_X1 U7650 ( .A(n6038), .ZN(n6041) );
  INV_X1 U7651 ( .A(n6039), .ZN(n6040) );
  NAND2_X1 U7652 ( .A1(n6041), .A2(n6040), .ZN(n6042) );
  AND2_X1 U7653 ( .A1(n6043), .A2(n6042), .ZN(n9013) );
  NAND2_X1 U7654 ( .A1(n7081), .A2(n7912), .ZN(n6046) );
  XNOR2_X1 U7655 ( .A(n6044), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7519) );
  AOI22_X1 U7656 ( .A1(n6082), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6081), .B2(
        n7519), .ZN(n6045) );
  NAND2_X1 U7657 ( .A1(n9501), .A2(n8184), .ZN(n6054) );
  INV_X1 U7658 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n6052) );
  INV_X1 U7659 ( .A(n6068), .ZN(n6070) );
  NAND2_X1 U7660 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  NAND2_X1 U7661 ( .A1(n6070), .A2(n6049), .ZN(n9401) );
  OR2_X1 U7662 ( .A1(n9401), .A2(n6209), .ZN(n6051) );
  AOI22_X1 U7663 ( .A1(n6434), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n6435), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n6050) );
  OAI211_X1 U7664 ( .C1(n6220), .C2(n6052), .A(n6051), .B(n6050), .ZN(n9381)
         );
  NAND2_X1 U7665 ( .A1(n9381), .A2(n4355), .ZN(n6053) );
  NAND2_X1 U7666 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  XNOR2_X1 U7667 ( .A(n6055), .B(n8182), .ZN(n6057) );
  AND2_X1 U7668 ( .A1(n9381), .A2(n8179), .ZN(n6056) );
  AOI21_X1 U7669 ( .B1(n9501), .B2(n4355), .A(n6056), .ZN(n6058) );
  XNOR2_X1 U7670 ( .A(n6057), .B(n6058), .ZN(n9025) );
  NAND2_X1 U7671 ( .A1(n9024), .A2(n9025), .ZN(n9023) );
  INV_X1 U7672 ( .A(n6057), .ZN(n6059) );
  NAND2_X1 U7673 ( .A1(n6059), .A2(n6058), .ZN(n6060) );
  NAND2_X1 U7674 ( .A1(n9023), .A2(n6060), .ZN(n6079) );
  NAND2_X1 U7675 ( .A1(n7108), .A2(n7912), .ZN(n6067) );
  NAND2_X1 U7676 ( .A1(n6061), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6063) );
  OR2_X1 U7677 ( .A1(n6063), .A2(n6062), .ZN(n6065) );
  NAND2_X1 U7678 ( .A1(n6063), .A2(n6062), .ZN(n6064) );
  AND2_X1 U7679 ( .A1(n6065), .A2(n6064), .ZN(n8102) );
  AOI22_X1 U7680 ( .A1(n6082), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6081), .B2(
        n8102), .ZN(n6066) );
  NAND2_X1 U7681 ( .A1(n9494), .A2(n8184), .ZN(n6076) );
  INV_X1 U7682 ( .A(n6085), .ZN(n6087) );
  INV_X1 U7683 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7684 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  NAND2_X1 U7685 ( .A1(n6087), .A2(n6071), .ZN(n9388) );
  AOI22_X1 U7686 ( .A1(n6434), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6072), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U7687 ( .A1(n6433), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6073) );
  OAI211_X1 U7688 ( .C1(n9388), .C2(n6209), .A(n6074), .B(n6073), .ZN(n9361)
         );
  NAND2_X1 U7689 ( .A1(n9361), .A2(n6174), .ZN(n6075) );
  NAND2_X1 U7690 ( .A1(n6076), .A2(n6075), .ZN(n6077) );
  XNOR2_X1 U7691 ( .A(n6077), .B(n4356), .ZN(n6078) );
  AND2_X1 U7692 ( .A1(n9361), .A2(n8179), .ZN(n6080) );
  AOI21_X1 U7693 ( .B1(n9494), .B2(n4355), .A(n6080), .ZN(n9089) );
  NAND2_X1 U7694 ( .A1(n7261), .A2(n7912), .ZN(n6084) );
  AOI22_X1 U7695 ( .A1(n6082), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8108), .B2(
        n6081), .ZN(n6083) );
  NAND2_X1 U7696 ( .A1(n9488), .A2(n8184), .ZN(n6095) );
  INV_X1 U7697 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7698 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  NAND2_X1 U7699 ( .A1(n6108), .A2(n6088), .ZN(n8982) );
  OR2_X1 U7700 ( .A1(n8982), .A2(n6209), .ZN(n6093) );
  INV_X1 U7701 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8099) );
  NAND2_X1 U7702 ( .A1(n6434), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7703 ( .A1(n6435), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6089) );
  OAI211_X1 U7704 ( .C1(n6220), .C2(n8099), .A(n6090), .B(n6089), .ZN(n6091)
         );
  INV_X1 U7705 ( .A(n6091), .ZN(n6092) );
  NAND2_X1 U7706 ( .A1(n6093), .A2(n6092), .ZN(n9382) );
  NAND2_X1 U7707 ( .A1(n9382), .A2(n4355), .ZN(n6094) );
  NAND2_X1 U7708 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  XNOR2_X1 U7709 ( .A(n6096), .B(n4356), .ZN(n6098) );
  AND2_X1 U7710 ( .A1(n9382), .A2(n8179), .ZN(n6097) );
  AOI21_X1 U7711 ( .B1(n9488), .B2(n4355), .A(n6097), .ZN(n6099) );
  NAND2_X1 U7712 ( .A1(n6098), .A2(n6099), .ZN(n9055) );
  INV_X1 U7713 ( .A(n6098), .ZN(n6101) );
  INV_X1 U7714 ( .A(n6099), .ZN(n6100) );
  NAND2_X1 U7715 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  AND2_X1 U7716 ( .A1(n9055), .A2(n6102), .ZN(n8987) );
  NAND2_X1 U7717 ( .A1(n8985), .A2(n9055), .ZN(n6125) );
  NAND2_X1 U7718 ( .A1(n7347), .A2(n7912), .ZN(n6106) );
  INV_X1 U7719 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6104) );
  OR2_X1 U7720 ( .A1(n5784), .A2(n6104), .ZN(n6105) );
  NAND2_X1 U7721 ( .A1(n9483), .A2(n8184), .ZN(n6117) );
  INV_X1 U7722 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6107) );
  NAND2_X1 U7723 ( .A1(n6108), .A2(n6107), .ZN(n6109) );
  AND2_X1 U7724 ( .A1(n6129), .A2(n6109), .ZN(n9352) );
  NAND2_X1 U7725 ( .A1(n9352), .A2(n6334), .ZN(n6115) );
  INV_X1 U7726 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7727 ( .A1(n6435), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U7728 ( .A1(n6434), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6110) );
  OAI211_X1 U7729 ( .C1(n6220), .C2(n6112), .A(n6111), .B(n6110), .ZN(n6113)
         );
  INV_X1 U7730 ( .A(n6113), .ZN(n6114) );
  NAND2_X1 U7731 ( .A1(n9362), .A2(n4355), .ZN(n6116) );
  NAND2_X1 U7732 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  XNOR2_X1 U7733 ( .A(n6118), .B(n4356), .ZN(n6120) );
  AND2_X1 U7734 ( .A1(n9362), .A2(n8179), .ZN(n6119) );
  AOI21_X1 U7735 ( .B1(n9483), .B2(n4355), .A(n6119), .ZN(n6121) );
  NAND2_X1 U7736 ( .A1(n6120), .A2(n6121), .ZN(n6126) );
  INV_X1 U7737 ( .A(n6120), .ZN(n6123) );
  INV_X1 U7738 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7739 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  AND2_X1 U7740 ( .A1(n6126), .A2(n6124), .ZN(n9053) );
  NAND2_X2 U7741 ( .A1(n6125), .A2(n9053), .ZN(n9057) );
  OR2_X1 U7742 ( .A1(n7416), .A2(n5765), .ZN(n6128) );
  INV_X1 U7743 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7415) );
  OR2_X1 U7744 ( .A1(n5784), .A2(n7415), .ZN(n6127) );
  NAND2_X1 U7745 ( .A1(n9479), .A2(n8184), .ZN(n6137) );
  INV_X1 U7746 ( .A(n6146), .ZN(n6162) );
  NAND2_X1 U7747 ( .A1(n6129), .A2(n8998), .ZN(n6130) );
  NAND2_X1 U7748 ( .A1(n6162), .A2(n6130), .ZN(n9339) );
  INV_X1 U7749 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9338) );
  NAND2_X1 U7750 ( .A1(n6435), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7751 ( .A1(n6434), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6131) );
  OAI211_X1 U7752 ( .C1(n6220), .C2(n9338), .A(n6132), .B(n6131), .ZN(n6133)
         );
  INV_X1 U7753 ( .A(n6133), .ZN(n6134) );
  NAND2_X1 U7754 ( .A1(n9468), .A2(n4355), .ZN(n6136) );
  NAND2_X1 U7755 ( .A1(n6137), .A2(n6136), .ZN(n6138) );
  XNOR2_X1 U7756 ( .A(n6138), .B(n8182), .ZN(n6140) );
  AND2_X1 U7757 ( .A1(n9468), .A2(n8179), .ZN(n6139) );
  AOI21_X1 U7758 ( .B1(n9479), .B2(n4355), .A(n6139), .ZN(n6141) );
  XNOR2_X1 U7759 ( .A(n6140), .B(n6141), .ZN(n8996) );
  INV_X1 U7760 ( .A(n6140), .ZN(n6142) );
  NAND2_X1 U7761 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  NAND2_X1 U7762 ( .A1(n7629), .A2(n7912), .ZN(n6145) );
  INV_X1 U7763 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7631) );
  OR2_X1 U7764 ( .A1(n5784), .A2(n7631), .ZN(n6144) );
  NAND2_X1 U7765 ( .A1(n9464), .A2(n8184), .ZN(n6155) );
  NAND2_X1 U7766 ( .A1(n6146), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6164) );
  INV_X1 U7767 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8977) );
  NAND2_X1 U7768 ( .A1(n6164), .A2(n8977), .ZN(n6147) );
  NAND2_X1 U7769 ( .A1(n6187), .A2(n6147), .ZN(n9307) );
  OR2_X1 U7770 ( .A1(n9307), .A2(n6209), .ZN(n6153) );
  INV_X1 U7771 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U7772 ( .A1(n6435), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7773 ( .A1(n6434), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6148) );
  OAI211_X1 U7774 ( .C1(n6220), .C2(n6150), .A(n6149), .B(n6148), .ZN(n6151)
         );
  INV_X1 U7775 ( .A(n6151), .ZN(n6152) );
  NAND2_X1 U7776 ( .A1(n6153), .A2(n6152), .ZN(n9469) );
  NAND2_X1 U7777 ( .A1(n9469), .A2(n4355), .ZN(n6154) );
  NAND2_X1 U7778 ( .A1(n6155), .A2(n6154), .ZN(n6156) );
  XNOR2_X1 U7779 ( .A(n6156), .B(n8182), .ZN(n6180) );
  NAND2_X1 U7780 ( .A1(n9464), .A2(n8178), .ZN(n6158) );
  NAND2_X1 U7781 ( .A1(n9469), .A2(n8179), .ZN(n6157) );
  NAND2_X1 U7782 ( .A1(n6158), .A2(n6157), .ZN(n6181) );
  NAND2_X1 U7783 ( .A1(n6180), .A2(n6181), .ZN(n8974) );
  NAND2_X1 U7784 ( .A1(n7592), .A2(n7912), .ZN(n6160) );
  INV_X1 U7785 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7594) );
  OR2_X1 U7786 ( .A1(n5784), .A2(n7594), .ZN(n6159) );
  NAND2_X1 U7787 ( .A1(n9328), .A2(n8184), .ZN(n6171) );
  INV_X1 U7788 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9069) );
  NAND2_X1 U7789 ( .A1(n6162), .A2(n9069), .ZN(n6163) );
  NAND2_X1 U7790 ( .A1(n6164), .A2(n6163), .ZN(n9324) );
  INV_X1 U7791 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U7792 ( .A1(n6435), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7793 ( .A1(n6434), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6165) );
  OAI211_X1 U7794 ( .C1(n6220), .C2(n9323), .A(n6166), .B(n6165), .ZN(n6167)
         );
  INV_X1 U7795 ( .A(n6167), .ZN(n6168) );
  NAND2_X1 U7796 ( .A1(n9304), .A2(n6174), .ZN(n6170) );
  NAND2_X1 U7797 ( .A1(n6171), .A2(n6170), .ZN(n6173) );
  XNOR2_X1 U7798 ( .A(n6173), .B(n4356), .ZN(n8973) );
  NAND2_X1 U7799 ( .A1(n9328), .A2(n6174), .ZN(n6176) );
  NAND2_X1 U7800 ( .A1(n9304), .A2(n8179), .ZN(n6175) );
  INV_X1 U7801 ( .A(n8973), .ZN(n8971) );
  INV_X1 U7802 ( .A(n9064), .ZN(n6179) );
  NOR2_X1 U7803 ( .A1(n8971), .A2(n6179), .ZN(n6184) );
  INV_X1 U7804 ( .A(n6180), .ZN(n6183) );
  INV_X1 U7805 ( .A(n6181), .ZN(n6182) );
  AOI21_X1 U7806 ( .B1(n6184), .B2(n8974), .A(n9032), .ZN(n6198) );
  NAND2_X1 U7807 ( .A1(n7718), .A2(n7912), .ZN(n6186) );
  INV_X1 U7808 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7719) );
  OR2_X1 U7809 ( .A1(n5784), .A2(n7719), .ZN(n6185) );
  NAND2_X1 U7810 ( .A1(n6187), .A2(n9037), .ZN(n6188) );
  AND2_X1 U7811 ( .A1(n6203), .A2(n6188), .ZN(n9294) );
  NAND2_X1 U7812 ( .A1(n9294), .A2(n6334), .ZN(n6194) );
  INV_X1 U7813 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7814 ( .A1(n6435), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7815 ( .A1(n6434), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6189) );
  OAI211_X1 U7816 ( .C1(n6220), .C2(n6191), .A(n6190), .B(n6189), .ZN(n6192)
         );
  INV_X1 U7817 ( .A(n6192), .ZN(n6193) );
  AOI22_X1 U7818 ( .A1(n9456), .A2(n8184), .B1(n6174), .B2(n9446), .ZN(n6195)
         );
  XNOR2_X1 U7819 ( .A(n6195), .B(n8182), .ZN(n6197) );
  AOI22_X1 U7820 ( .A1(n9456), .A2(n4355), .B1(n8179), .B2(n9446), .ZN(n6196)
         );
  NAND2_X1 U7821 ( .A1(n6197), .A2(n6196), .ZN(n6199) );
  OAI21_X1 U7822 ( .B1(n6197), .B2(n6196), .A(n6199), .ZN(n9031) );
  NAND2_X1 U7823 ( .A1(n7750), .A2(n7912), .ZN(n6201) );
  INV_X1 U7824 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7752) );
  OR2_X1 U7825 ( .A1(n5784), .A2(n7752), .ZN(n6200) );
  NAND2_X1 U7826 ( .A1(n9281), .A2(n8184), .ZN(n6211) );
  INV_X1 U7827 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6202) );
  AND2_X1 U7828 ( .A1(n6203), .A2(n6202), .ZN(n6204) );
  INV_X1 U7829 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9276) );
  NAND2_X1 U7830 ( .A1(n6435), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7831 ( .A1(n6434), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6205) );
  OAI211_X1 U7832 ( .C1(n6220), .C2(n9276), .A(n6206), .B(n6205), .ZN(n6207)
         );
  INV_X1 U7833 ( .A(n6207), .ZN(n6208) );
  NAND2_X1 U7834 ( .A1(n9262), .A2(n8178), .ZN(n6210) );
  NAND2_X1 U7835 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  XNOR2_X1 U7836 ( .A(n6212), .B(n8182), .ZN(n6230) );
  OAI22_X1 U7837 ( .A1(n9450), .A2(n5734), .B1(n9439), .B2(n6213), .ZN(n6229)
         );
  XNOR2_X1 U7838 ( .A(n6230), .B(n6229), .ZN(n9005) );
  NAND2_X1 U7839 ( .A1(n7770), .A2(n7912), .ZN(n6215) );
  INV_X1 U7840 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7773) );
  OR2_X1 U7841 ( .A1(n5784), .A2(n7773), .ZN(n6214) );
  OR2_X1 U7842 ( .A1(n6216), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7843 ( .A1(n6216), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6279) );
  AND2_X1 U7844 ( .A1(n6217), .A2(n6279), .ZN(n9101) );
  NAND2_X1 U7845 ( .A1(n9101), .A2(n6334), .ZN(n6223) );
  INV_X1 U7846 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9258) );
  NAND2_X1 U7847 ( .A1(n6435), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7848 ( .A1(n6434), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6218) );
  OAI211_X1 U7849 ( .C1(n6220), .C2(n9258), .A(n6219), .B(n6218), .ZN(n6221)
         );
  INV_X1 U7850 ( .A(n6221), .ZN(n6222) );
  AND2_X1 U7851 ( .A1(n9447), .A2(n8179), .ZN(n6224) );
  AOI21_X1 U7852 ( .B1(n9442), .B2(n4355), .A(n6224), .ZN(n6233) );
  NAND2_X1 U7853 ( .A1(n9442), .A2(n8184), .ZN(n6227) );
  NAND2_X1 U7854 ( .A1(n9447), .A2(n8178), .ZN(n6226) );
  NAND2_X1 U7855 ( .A1(n6227), .A2(n6226), .ZN(n6228) );
  XNOR2_X1 U7856 ( .A(n6228), .B(n8182), .ZN(n6235) );
  XOR2_X1 U7857 ( .A(n6233), .B(n6235), .Z(n9097) );
  INV_X1 U7858 ( .A(n9097), .ZN(n6232) );
  NOR2_X1 U7859 ( .A1(n6230), .A2(n6229), .ZN(n9098) );
  INV_X1 U7860 ( .A(n9098), .ZN(n6231) );
  INV_X1 U7861 ( .A(n6233), .ZN(n6234) );
  NAND2_X1 U7862 ( .A1(n8094), .A2(n7912), .ZN(n6237) );
  INV_X1 U7863 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8096) );
  OR2_X1 U7864 ( .A1(n5784), .A2(n8096), .ZN(n6236) );
  XNOR2_X1 U7865 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n6279), .ZN(n9245) );
  NAND2_X1 U7866 ( .A1(n6334), .A2(n9245), .ZN(n6241) );
  NAND2_X1 U7867 ( .A1(n6433), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7868 ( .A1(n6434), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7869 ( .A1(n6435), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6238) );
  NAND4_X1 U7870 ( .A1(n6241), .A2(n6240), .A3(n6239), .A4(n6238), .ZN(n9238)
         );
  AOI22_X1 U7871 ( .A1(n9433), .A2(n8184), .B1(n4355), .B2(n9238), .ZN(n6242)
         );
  XNOR2_X1 U7872 ( .A(n6242), .B(n8182), .ZN(n6244) );
  AOI22_X1 U7873 ( .A1(n9433), .A2(n6174), .B1(n8179), .B2(n9238), .ZN(n6243)
         );
  NAND2_X1 U7874 ( .A1(n6244), .A2(n6243), .ZN(n8190) );
  OAI21_X1 U7875 ( .B1(n6244), .B2(n6243), .A(n8190), .ZN(n6245) );
  NAND2_X1 U7876 ( .A1(n7755), .A2(P1_B_REG_SCAN_IN), .ZN(n6248) );
  MUX2_X1 U7877 ( .A(P1_B_REG_SCAN_IN), .B(n6248), .S(n7720), .Z(n6249) );
  INV_X1 U7878 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6251) );
  NOR4_X1 U7879 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6261) );
  NOR4_X1 U7880 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6260) );
  OR4_X1 U7881 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6258) );
  NOR4_X1 U7882 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6256) );
  NOR4_X1 U7883 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6255) );
  NOR4_X1 U7884 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6254) );
  NOR4_X1 U7885 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6253) );
  NAND4_X1 U7886 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n6257)
         );
  NOR4_X1 U7887 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6258), .A4(n6257), .ZN(n6259) );
  NAND3_X1 U7888 ( .A1(n6261), .A2(n6260), .A3(n6259), .ZN(n6262) );
  NAND2_X1 U7889 ( .A1(n6405), .A2(n6262), .ZN(n6739) );
  NAND3_X1 U7890 ( .A1(n6742), .A2(n6741), .A3(n6739), .ZN(n6272) );
  NAND2_X1 U7891 ( .A1(n6263), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7892 ( .A1(n9678), .A2(n6274), .ZN(n6266) );
  INV_X1 U7893 ( .A(n9433), .ZN(n9250) );
  INV_X1 U7894 ( .A(n6278), .ZN(n6267) );
  INV_X1 U7895 ( .A(n6744), .ZN(n6753) );
  NOR2_X1 U7896 ( .A1(n6753), .A2(n8064), .ZN(n6926) );
  NAND2_X1 U7897 ( .A1(n6267), .A2(n6926), .ZN(n6268) );
  NAND2_X1 U7898 ( .A1(n9581), .A2(n8108), .ZN(n6373) );
  INV_X1 U7899 ( .A(n6269), .ZN(n6452) );
  OR2_X1 U7900 ( .A1(n9705), .A2(n6341), .ZN(n6270) );
  CLKBUF_X1 U7901 ( .A(n9081), .Z(n9116) );
  INV_X1 U7902 ( .A(n9245), .ZN(n6291) );
  NOR2_X1 U7903 ( .A1(n8064), .A2(P1_U3086), .ZN(n7348) );
  OR2_X1 U7904 ( .A1(n9678), .A2(n7348), .ZN(n6271) );
  NAND2_X1 U7905 ( .A1(n6272), .A2(n6271), .ZN(n6276) );
  OAI211_X1 U7906 ( .C1(n6274), .C2(n8079), .A(n6273), .B(n6398), .ZN(n6372)
         );
  INV_X1 U7907 ( .A(n6372), .ZN(n6275) );
  NAND2_X1 U7908 ( .A1(n6276), .A2(n6275), .ZN(n6521) );
  NAND2_X1 U7909 ( .A1(n6521), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9112) );
  NAND2_X1 U7910 ( .A1(n7995), .A2(n6269), .ZN(n9703) );
  OR2_X1 U7911 ( .A1(n9703), .A2(n6341), .ZN(n6277) );
  NOR2_X2 U7912 ( .A1(n6278), .A2(n6277), .ZN(n9102) );
  INV_X1 U7913 ( .A(n6279), .ZN(n6280) );
  NAND2_X1 U7914 ( .A1(n6281), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8115) );
  INV_X1 U7915 ( .A(n6281), .ZN(n6283) );
  INV_X1 U7916 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U7917 ( .A1(n6283), .A2(n6282), .ZN(n6284) );
  NAND2_X1 U7918 ( .A1(n6285), .A2(n9235), .ZN(n6289) );
  NAND2_X1 U7919 ( .A1(n6433), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7920 ( .A1(n6434), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7921 ( .A1(n6435), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6286) );
  NAND4_X1 U7922 ( .A1(n6289), .A2(n6288), .A3(n6287), .A4(n6286), .ZN(n9120)
         );
  AOI22_X1 U7923 ( .A1(n9102), .A2(n9120), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6290) );
  OAI21_X1 U7924 ( .B1(n6291), .B2(n9112), .A(n6290), .ZN(n6292) );
  AOI21_X1 U7925 ( .B1(n9447), .B2(n9116), .A(n6292), .ZN(n6293) );
  INV_X1 U7926 ( .A(n6293), .ZN(n6294) );
  NAND2_X1 U7927 ( .A1(n6297), .A2(n6296), .ZN(P1_U3214) );
  INV_X1 U7928 ( .A(n9456), .ZN(n9297) );
  INV_X1 U7929 ( .A(n9479), .ZN(n9337) );
  INV_X1 U7930 ( .A(n9468), .ZN(n9071) );
  INV_X1 U7931 ( .A(n9483), .ZN(n9354) );
  INV_X1 U7932 ( .A(n9382), .ZN(n9091) );
  INV_X1 U7933 ( .A(n9488), .ZN(n9370) );
  INV_X1 U7934 ( .A(n9361), .ZN(n9498) );
  INV_X1 U7935 ( .A(n9494), .ZN(n9096) );
  AND2_X1 U7936 ( .A1(n9494), .A2(n9361), .ZN(n6319) );
  INV_X1 U7937 ( .A(n9381), .ZN(n9017) );
  INV_X1 U7938 ( .A(n9709), .ZN(n7437) );
  AND2_X1 U7939 ( .A1(n9127), .A2(n6745), .ZN(n6924) );
  OR2_X1 U7940 ( .A1(n9599), .A2(n7792), .ZN(n6298) );
  INV_X1 U7941 ( .A(n9083), .ZN(n9602) );
  NAND2_X1 U7942 ( .A1(n9125), .A2(n9602), .ZN(n8008) );
  NAND2_X1 U7943 ( .A1(n7023), .A2(n7021), .ZN(n6300) );
  OR2_X1 U7944 ( .A1(n9125), .A2(n9083), .ZN(n6299) );
  NAND2_X1 U7945 ( .A1(n9598), .A2(n6991), .ZN(n7798) );
  NAND2_X1 U7946 ( .A1(n7809), .A2(n7798), .ZN(n7935) );
  NAND2_X1 U7947 ( .A1(n6986), .A2(n7935), .ZN(n6302) );
  OR2_X1 U7948 ( .A1(n9598), .A2(n9609), .ZN(n6301) );
  NAND2_X1 U7949 ( .A1(n6302), .A2(n6301), .ZN(n7041) );
  INV_X1 U7950 ( .A(n9124), .ZN(n6303) );
  NAND2_X1 U7951 ( .A1(n6303), .A2(n9616), .ZN(n7810) );
  INV_X1 U7952 ( .A(n9616), .ZN(n7047) );
  NAND2_X1 U7953 ( .A1(n9124), .A2(n7047), .ZN(n7813) );
  NAND2_X1 U7954 ( .A1(n7041), .A2(n7040), .ZN(n6970) );
  NAND2_X1 U7955 ( .A1(n6303), .A2(n7047), .ZN(n6969) );
  OR2_X1 U7956 ( .A1(n9617), .A2(n6976), .ZN(n7055) );
  OR2_X1 U7957 ( .A1(n9577), .A2(n9639), .ZN(n7057) );
  OR2_X1 U7958 ( .A1(n4352), .A2(n9569), .ZN(n6311) );
  AND2_X1 U7959 ( .A1(n7057), .A2(n6311), .ZN(n6304) );
  AND2_X1 U7960 ( .A1(n6969), .A2(n6306), .ZN(n6309) );
  INV_X1 U7961 ( .A(n6304), .ZN(n6305) );
  NAND2_X1 U7962 ( .A1(n7818), .A2(n7937), .ZN(n9579) );
  OR2_X1 U7963 ( .A1(n6305), .A2(n9579), .ZN(n6308) );
  INV_X1 U7964 ( .A(n6976), .ZN(n9626) );
  NAND2_X1 U7965 ( .A1(n9617), .A2(n9626), .ZN(n8013) );
  INV_X1 U7966 ( .A(n9658), .ZN(n7067) );
  OR2_X1 U7967 ( .A1(n6310), .A2(n7067), .ZN(n7820) );
  NAND2_X1 U7968 ( .A1(n6310), .A2(n7067), .ZN(n7803) );
  NAND2_X1 U7969 ( .A1(n7820), .A2(n7803), .ZN(n9552) );
  INV_X1 U7970 ( .A(n6311), .ZN(n6312) );
  INV_X1 U7971 ( .A(n9569), .ZN(n6919) );
  NAND2_X1 U7972 ( .A1(n4352), .A2(n6919), .ZN(n7804) );
  AND2_X1 U7973 ( .A1(n9552), .A2(n9550), .ZN(n7113) );
  INV_X1 U7974 ( .A(n9553), .ZN(n7241) );
  NAND2_X1 U7975 ( .A1(n9660), .A2(n7241), .ZN(n7828) );
  AND2_X1 U7976 ( .A1(n7113), .A2(n7121), .ZN(n6314) );
  INV_X1 U7977 ( .A(n7121), .ZN(n6313) );
  OR2_X1 U7978 ( .A1(n6310), .A2(n9658), .ZN(n7114) );
  OR2_X1 U7979 ( .A1(n9660), .A2(n9553), .ZN(n6315) );
  INV_X1 U7980 ( .A(n9123), .ZN(n7301) );
  NOR2_X1 U7981 ( .A1(n9670), .A2(n7301), .ZN(n8020) );
  INV_X1 U7982 ( .A(n8020), .ZN(n7826) );
  NAND2_X1 U7983 ( .A1(n9670), .A2(n7301), .ZN(n7830) );
  NOR2_X1 U7984 ( .A1(n9670), .A2(n9123), .ZN(n6316) );
  AOI21_X2 U7985 ( .B1(n7105), .B2(n7104), .A(n6316), .ZN(n7165) );
  INV_X1 U7986 ( .A(n9669), .ZN(n7478) );
  NAND2_X1 U7987 ( .A1(n7292), .A2(n7478), .ZN(n7831) );
  INV_X1 U7988 ( .A(n7944), .ZN(n7164) );
  OAI22_X1 U7989 ( .A1(n7165), .A2(n7164), .B1(n7292), .B2(n9669), .ZN(n7418)
         );
  INV_X1 U7990 ( .A(n9122), .ZN(n6317) );
  AOI22_X1 U7991 ( .A1(n7418), .A2(n7417), .B1(n4604), .B2(n6317), .ZN(n7352)
         );
  NOR2_X1 U7992 ( .A1(n9696), .A2(n9706), .ZN(n7840) );
  INV_X1 U7993 ( .A(n7840), .ZN(n7838) );
  NAND2_X1 U7994 ( .A1(n9696), .A2(n9706), .ZN(n8026) );
  INV_X1 U7995 ( .A(n7597), .ZN(n6318) );
  INV_X1 U7996 ( .A(n7609), .ZN(n9542) );
  AND2_X1 U7997 ( .A1(n9507), .A2(n9497), .ZN(n7845) );
  INV_X1 U7998 ( .A(n9507), .ZN(n9022) );
  OAI21_X1 U7999 ( .B1(n9091), .B2(n9370), .A(n6320), .ZN(n9355) );
  NAND2_X1 U8000 ( .A1(n9464), .A2(n9469), .ZN(n6322) );
  INV_X1 U8001 ( .A(n9464), .ZN(n6321) );
  NAND2_X1 U8002 ( .A1(n9456), .A2(n9461), .ZN(n7976) );
  NAND2_X1 U8003 ( .A1(n7969), .A2(n7976), .ZN(n9289) );
  NOR2_X1 U8004 ( .A1(n9442), .A2(n9430), .ZN(n7893) );
  INV_X1 U8005 ( .A(n7893), .ZN(n7964) );
  NAND2_X1 U8006 ( .A1(n9442), .A2(n9430), .ZN(n8044) );
  NAND2_X1 U8007 ( .A1(n7964), .A2(n8044), .ZN(n9255) );
  NAND2_X1 U8008 ( .A1(n9256), .A2(n9255), .ZN(n6326) );
  NAND2_X1 U8009 ( .A1(n9442), .A2(n9447), .ZN(n6325) );
  NAND2_X1 U8010 ( .A1(n6326), .A2(n6325), .ZN(n9243) );
  OR2_X1 U8011 ( .A1(n9433), .A2(n9438), .ZN(n7965) );
  NAND2_X1 U8012 ( .A1(n9433), .A2(n9438), .ZN(n7986) );
  NAND2_X1 U8013 ( .A1(n7965), .A2(n7986), .ZN(n9244) );
  NAND2_X1 U8014 ( .A1(n8964), .A2(n7912), .ZN(n6328) );
  INV_X1 U8015 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7787) );
  OR2_X1 U8016 ( .A1(n5784), .A2(n7787), .ZN(n6327) );
  OR2_X1 U8017 ( .A1(n9424), .A2(n9429), .ZN(n7962) );
  NAND2_X1 U8018 ( .A1(n9424), .A2(n9429), .ZN(n7987) );
  NAND2_X1 U8019 ( .A1(n7962), .A2(n7987), .ZN(n9229) );
  NAND2_X1 U8020 ( .A1(n8198), .A2(n7912), .ZN(n6330) );
  INV_X1 U8021 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8200) );
  OR2_X1 U8022 ( .A1(n5784), .A2(n8200), .ZN(n6329) );
  NAND2_X1 U8023 ( .A1(n6434), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U8024 ( .A1(n6435), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6331) );
  AND2_X1 U8025 ( .A1(n6332), .A2(n6331), .ZN(n6337) );
  INV_X1 U8026 ( .A(n8115), .ZN(n6333) );
  NAND2_X1 U8027 ( .A1(n6334), .A2(n6333), .ZN(n6336) );
  NAND2_X1 U8028 ( .A1(n6433), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6335) );
  OR2_X1 U8029 ( .A1(n8114), .A2(n9421), .ZN(n7963) );
  NAND2_X1 U8030 ( .A1(n8114), .A2(n9421), .ZN(n7990) );
  NAND2_X1 U8031 ( .A1(n7963), .A2(n7990), .ZN(n7957) );
  INV_X1 U8032 ( .A(n7957), .ZN(n6338) );
  XNOR2_X1 U8033 ( .A(n6339), .B(n6338), .ZN(n8113) );
  NAND2_X1 U8034 ( .A1(n7995), .A2(n8079), .ZN(n6752) );
  NAND2_X1 U8035 ( .A1(n6341), .A2(n6340), .ZN(n6342) );
  NAND3_X1 U8036 ( .A1(n6752), .A2(n6753), .A3(n6342), .ZN(n9647) );
  NAND2_X1 U8037 ( .A1(n7926), .A2(n8064), .ZN(n9654) );
  INV_X1 U8038 ( .A(n6745), .ZN(n6925) );
  INV_X1 U8039 ( .A(n7792), .ZN(n9593) );
  OR2_X1 U8040 ( .A1(n9599), .A2(n9593), .ZN(n6343) );
  INV_X1 U8041 ( .A(n7935), .ZN(n6987) );
  NAND2_X1 U8042 ( .A1(n7035), .A2(n7809), .ZN(n6345) );
  NAND2_X1 U8043 ( .A1(n6345), .A2(n7938), .ZN(n6963) );
  NAND2_X1 U8044 ( .A1(n6963), .A2(n7810), .ZN(n6346) );
  AND2_X1 U8045 ( .A1(n7828), .A2(n7803), .ZN(n7821) );
  INV_X1 U8046 ( .A(n7804), .ZN(n7117) );
  AND2_X1 U8047 ( .A1(n7823), .A2(n7820), .ZN(n7806) );
  INV_X1 U8048 ( .A(n7806), .ZN(n6349) );
  NAND2_X1 U8049 ( .A1(n6349), .A2(n7828), .ZN(n6347) );
  NAND2_X1 U8050 ( .A1(n7819), .A2(n7818), .ZN(n6348) );
  NOR2_X1 U8051 ( .A1(n6349), .A2(n6348), .ZN(n8017) );
  INV_X1 U8052 ( .A(n7833), .ZN(n6351) );
  INV_X1 U8053 ( .A(n8026), .ZN(n6353) );
  OR2_X1 U8054 ( .A1(n9709), .A2(n7408), .ZN(n8028) );
  NAND2_X1 U8055 ( .A1(n9709), .A2(n7408), .ZN(n7836) );
  NAND2_X1 U8056 ( .A1(n7609), .A2(n9704), .ZN(n7843) );
  NAND2_X1 U8057 ( .A1(n7841), .A2(n7843), .ZN(n7950) );
  INV_X1 U8058 ( .A(n7950), .ZN(n7599) );
  NAND2_X1 U8059 ( .A1(n7659), .A2(n7952), .ZN(n7658) );
  NAND2_X1 U8060 ( .A1(n7658), .A2(n7846), .ZN(n9410) );
  OR2_X1 U8061 ( .A1(n9501), .A2(n9017), .ZN(n8035) );
  NAND2_X1 U8062 ( .A1(n9501), .A2(n9017), .ZN(n7851) );
  NAND2_X1 U8063 ( .A1(n9410), .A2(n9409), .ZN(n9408) );
  NAND2_X1 U8064 ( .A1(n9408), .A2(n8035), .ZN(n9379) );
  NAND2_X1 U8065 ( .A1(n9494), .A2(n9498), .ZN(n7852) );
  NAND2_X1 U8066 ( .A1(n7854), .A2(n7852), .ZN(n9376) );
  INV_X1 U8067 ( .A(n9376), .ZN(n9380) );
  NAND2_X1 U8068 ( .A1(n9379), .A2(n9380), .ZN(n9378) );
  NAND2_X1 U8069 ( .A1(n9488), .A2(n9091), .ZN(n8039) );
  NAND2_X1 U8070 ( .A1(n9360), .A2(n8039), .ZN(n7983) );
  OR2_X1 U8071 ( .A1(n9483), .A2(n9345), .ZN(n7860) );
  OR2_X1 U8072 ( .A1(n9488), .A2(n9091), .ZN(n7982) );
  NAND2_X1 U8073 ( .A1(n7860), .A2(n7982), .ZN(n7858) );
  INV_X1 U8074 ( .A(n7858), .ZN(n6355) );
  NAND2_X1 U8075 ( .A1(n9483), .A2(n9345), .ZN(n7859) );
  INV_X1 U8076 ( .A(n7859), .ZN(n6354) );
  XNOR2_X1 U8077 ( .A(n9479), .B(n9468), .ZN(n9342) );
  INV_X1 U8078 ( .A(n9342), .ZN(n9335) );
  NAND2_X1 U8079 ( .A1(n9479), .A2(n9071), .ZN(n7863) );
  XNOR2_X1 U8080 ( .A(n9328), .B(n9304), .ZN(n9320) );
  NAND2_X1 U8081 ( .A1(n9328), .A2(n9460), .ZN(n7868) );
  INV_X1 U8082 ( .A(n7868), .ZN(n6356) );
  NAND2_X1 U8083 ( .A1(n9464), .A2(n9325), .ZN(n7966) );
  NAND2_X1 U8084 ( .A1(n7871), .A2(n7966), .ZN(n9312) );
  INV_X1 U8085 ( .A(n7969), .ZN(n9272) );
  OR2_X1 U8086 ( .A1(n9281), .A2(n9439), .ZN(n7972) );
  NAND2_X1 U8087 ( .A1(n9281), .A2(n9439), .ZN(n7878) );
  NAND2_X1 U8088 ( .A1(n7972), .A2(n7878), .ZN(n9271) );
  INV_X1 U8089 ( .A(n7878), .ZN(n7979) );
  INV_X1 U8090 ( .A(n8044), .ZN(n6357) );
  INV_X1 U8091 ( .A(n9229), .ZN(n9231) );
  NAND2_X1 U8092 ( .A1(n9230), .A2(n7987), .ZN(n6358) );
  XNOR2_X1 U8093 ( .A(n6358), .B(n6338), .ZN(n6368) );
  NAND2_X1 U8094 ( .A1(n8072), .A2(n8108), .ZN(n6361) );
  INV_X1 U8095 ( .A(n8064), .ZN(n6359) );
  AND2_X1 U8096 ( .A1(n6359), .A2(n8006), .ZN(n8074) );
  NAND2_X1 U8097 ( .A1(n6433), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U8098 ( .A1(n6434), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8099 ( .A1(n6435), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6362) );
  NAND3_X1 U8100 ( .A1(n6364), .A2(n6363), .A3(n6362), .ZN(n7931) );
  INV_X1 U8101 ( .A(P1_B_REG_SCAN_IN), .ZN(n6365) );
  NOR2_X1 U8102 ( .A1(n8095), .A2(n6365), .ZN(n6366) );
  NOR2_X1 U8103 ( .A1(n9703), .A2(n6366), .ZN(n8090) );
  OR2_X1 U8104 ( .A1(n7792), .A2(n6745), .ZN(n7027) );
  NAND2_X1 U8105 ( .A1(n6989), .A2(n6991), .ZN(n7042) );
  OR2_X1 U8106 ( .A1(n7042), .A2(n9616), .ZN(n7043) );
  INV_X1 U8107 ( .A(n9577), .ZN(n9632) );
  NAND2_X1 U8108 ( .A1(n9583), .A2(n9632), .ZN(n9582) );
  OR2_X1 U8109 ( .A1(n9582), .A2(n4352), .ZN(n9563) );
  INV_X1 U8110 ( .A(n9660), .ZN(n6369) );
  INV_X1 U8111 ( .A(n9670), .ZN(n7100) );
  INV_X1 U8112 ( .A(n9696), .ZN(n7413) );
  NAND2_X1 U8113 ( .A1(n7438), .A2(n7437), .ZN(n7602) );
  NAND2_X1 U8114 ( .A1(n9397), .A2(n9396), .ZN(n9399) );
  NOR2_X2 U8115 ( .A1(n9399), .A2(n9494), .ZN(n9364) );
  AOI21_X1 U8116 ( .B1(n8114), .B2(n9233), .A(n9562), .ZN(n6371) );
  NOR2_X1 U8117 ( .A1(n6372), .A2(P1_U3086), .ZN(n6740) );
  NAND3_X1 U8118 ( .A1(n6739), .A2(n6740), .A3(n6373), .ZN(n6374) );
  INV_X1 U8119 ( .A(n6742), .ZN(n6375) );
  NAND2_X1 U8120 ( .A1(n9420), .A2(n9719), .ZN(n6377) );
  NAND2_X1 U8121 ( .A1(n6377), .A2(n6376), .ZN(P1_U3519) );
  INV_X1 U8122 ( .A(n6843), .ZN(n6381) );
  OR2_X1 U8123 ( .A1(n6382), .A2(n6381), .ZN(n6592) );
  NAND2_X1 U8124 ( .A1(n6843), .A2(n8554), .ZN(n6383) );
  NAND2_X1 U8125 ( .A1(n6592), .A2(n6383), .ZN(n6626) );
  OAI21_X1 U8126 ( .B1(n6626), .B2(n6384), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  OAI222_X1 U8127 ( .A1(n9536), .A2(n6385), .B1(n7754), .B2(n6387), .C1(
        P1_U3086), .C2(n9159), .ZN(P1_U3352) );
  AND2_X1 U8128 ( .A1(n7917), .A2(P2_U3151), .ZN(n8963) );
  INV_X2 U8129 ( .A(n6683), .ZN(n8968) );
  OAI222_X1 U8130 ( .A1(n9745), .A2(P2_U3151), .B1(n8205), .B2(n6387), .C1(
        n6386), .C2(n8968), .ZN(P2_U3292) );
  OAI222_X1 U8131 ( .A1(n4353), .A2(P2_U3151), .B1(n8205), .B2(n6401), .C1(
        n6388), .C2(n8968), .ZN(P2_U3293) );
  OAI222_X1 U8132 ( .A1(n6707), .A2(P2_U3151), .B1(n8205), .B2(n6390), .C1(
        n6389), .C2(n8968), .ZN(P2_U3291) );
  INV_X2 U8133 ( .A(n8963), .ZN(n8205) );
  OAI222_X1 U8134 ( .A1(n6641), .A2(P2_U3151), .B1(n8205), .B2(n6403), .C1(
        n5003), .C2(n8968), .ZN(P2_U3294) );
  INV_X2 U8135 ( .A(n7628), .ZN(n7754) );
  OAI222_X1 U8136 ( .A1(n6391), .A2(n9536), .B1(P1_U3086), .B2(n9178), .C1(
        n7754), .C2(n6390), .ZN(P1_U3351) );
  OAI222_X1 U8137 ( .A1(n6730), .A2(P2_U3151), .B1(n8205), .B2(n6393), .C1(
        n6392), .C2(n8968), .ZN(P2_U3290) );
  INV_X1 U8138 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6394) );
  INV_X1 U8139 ( .A(n6468), .ZN(n9188) );
  OAI222_X1 U8140 ( .A1(n9536), .A2(n6394), .B1(n7754), .B2(n6393), .C1(
        P1_U3086), .C2(n9188), .ZN(P1_U3350) );
  INV_X1 U8141 ( .A(n9536), .ZN(n9529) );
  AOI22_X1 U8142 ( .A1(n9216), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9529), .ZN(n6395) );
  OAI21_X1 U8143 ( .B1(n6396), .B2(n7754), .A(n6395), .ZN(P1_U3349) );
  OAI222_X1 U8144 ( .A1(n8968), .A2(n6397), .B1(n8205), .B2(n6396), .C1(n6832), 
        .C2(P2_U3151), .ZN(P2_U3289) );
  OR2_X1 U8145 ( .A1(n6398), .A2(P1_U3086), .ZN(n8073) );
  NAND2_X1 U8146 ( .A1(n6406), .A2(n8073), .ZN(n6425) );
  NAND2_X1 U8147 ( .A1(n6398), .A2(n7995), .ZN(n6399) );
  AND2_X1 U8148 ( .A1(n6399), .A2(n7923), .ZN(n6424) );
  INV_X1 U8149 ( .A(n6424), .ZN(n6400) );
  NOR2_X1 U8150 ( .A1(n9215), .A2(P1_U3973), .ZN(P1_U3085) );
  OAI222_X1 U8151 ( .A1(n9536), .A2(n6402), .B1(n7754), .B2(n6401), .C1(
        P1_U3086), .C2(n9151), .ZN(P1_U3353) );
  OAI222_X1 U8152 ( .A1(n9536), .A2(n6404), .B1(n7754), .B2(n6403), .C1(
        P1_U3086), .C2(n6459), .ZN(P1_U3354) );
  INV_X1 U8153 ( .A(n6405), .ZN(n6407) );
  INV_X1 U8154 ( .A(n6406), .ZN(n8080) );
  NAND2_X2 U8155 ( .A1(n6407), .A2(n8080), .ZN(n9589) );
  NAND2_X1 U8156 ( .A1(n9589), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6408) );
  OAI21_X1 U8157 ( .B1(n9589), .B2(n6409), .A(n6408), .ZN(P1_U3439) );
  NAND2_X1 U8158 ( .A1(n9589), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6410) );
  OAI21_X1 U8159 ( .B1(n9589), .B2(n6411), .A(n6410), .ZN(P1_U3440) );
  INV_X1 U8160 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6414) );
  INV_X1 U8161 ( .A(n6412), .ZN(n6413) );
  AOI22_X1 U8162 ( .A1(n6421), .A2(n6414), .B1(n6413), .B2(n6587), .ZN(
        P2_U3377) );
  INV_X1 U8163 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6417) );
  INV_X1 U8164 ( .A(n6415), .ZN(n6416) );
  AOI22_X1 U8165 ( .A1(n6421), .A2(n6417), .B1(n6416), .B2(n6587), .ZN(
        P2_U3376) );
  INV_X1 U8166 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6418) );
  INV_X1 U8167 ( .A(n6473), .ZN(n6486) );
  AND2_X1 U8168 ( .A1(n6421), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8169 ( .A1(n6421), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8170 ( .A1(n6421), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8171 ( .A1(n6421), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8172 ( .A1(n6421), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8173 ( .A1(n6421), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8174 ( .A1(n6421), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8175 ( .A1(n6421), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8176 ( .A1(n6421), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8177 ( .A1(n6421), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8178 ( .A1(n6421), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8179 ( .A1(n6421), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8180 ( .A1(n6421), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8181 ( .A1(n6421), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8182 ( .A1(n6421), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8183 ( .A1(n6421), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8184 ( .A1(n6421), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8185 ( .A1(n6421), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8186 ( .A1(n6421), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8187 ( .A1(n6421), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8188 ( .A1(n6421), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8189 ( .A1(n6421), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8190 ( .A1(n6421), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8191 ( .A1(n6421), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8192 ( .A1(n6421), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8193 ( .A1(n6421), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8194 ( .A1(n6421), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8195 ( .A1(n6421), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8196 ( .A1(n6421), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8197 ( .A1(n6421), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  OAI21_X1 U8198 ( .B1(n8095), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6452), .ZN(
        n9142) );
  INV_X1 U8199 ( .A(n9142), .ZN(n6423) );
  INV_X1 U8200 ( .A(n8095), .ZN(n9138) );
  OAI21_X1 U8201 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n9138), .A(n6423), .ZN(
        n6422) );
  INV_X1 U8202 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9141) );
  MUX2_X1 U8203 ( .A(n6423), .B(n6422), .S(n9141), .Z(n6429) );
  NAND2_X1 U8204 ( .A1(n6425), .A2(n6424), .ZN(n6476) );
  NAND3_X1 U8205 ( .A1(n9211), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6426), .ZN(
        n6428) );
  AOI22_X1 U8206 ( .A1(n9215), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6427) );
  OAI211_X1 U8207 ( .C1(n6429), .C2(n6476), .A(n6428), .B(n6427), .ZN(P1_U3243) );
  INV_X1 U8208 ( .A(n6430), .ZN(n6442) );
  AOI22_X1 U8209 ( .A1(n6504), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9529), .ZN(n6431) );
  OAI21_X1 U8210 ( .B1(n6442), .B2(n7754), .A(n6431), .ZN(P1_U3347) );
  INV_X1 U8211 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U8212 ( .A1(n7931), .A2(P1_U3973), .ZN(n6432) );
  OAI21_X1 U8213 ( .B1(n8127), .B2(P1_U3973), .A(n6432), .ZN(P1_U3584) );
  INV_X1 U8214 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8215 ( .A1(n6433), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U8216 ( .A1(n6434), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8217 ( .A1(n6435), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6436) );
  NAND3_X1 U8218 ( .A1(n6438), .A2(n6437), .A3(n6436), .ZN(n8091) );
  NAND2_X1 U8219 ( .A1(n8091), .A2(P1_U3973), .ZN(n6439) );
  OAI21_X1 U8220 ( .B1(P1_U3973), .B2(n6440), .A(n6439), .ZN(P1_U3585) );
  OAI222_X1 U8221 ( .A1(n9772), .A2(P2_U3151), .B1(n8205), .B2(n6442), .C1(
        n6441), .C2(n8968), .ZN(P2_U3287) );
  INV_X1 U8222 ( .A(n9151), .ZN(n6461) );
  INV_X1 U8223 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6443) );
  MUX2_X1 U8224 ( .A(n6443), .B(P1_REG1_REG_2__SCAN_IN), .S(n9151), .Z(n6446)
         );
  INV_X1 U8225 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6444) );
  MUX2_X1 U8226 ( .A(n6444), .B(P1_REG1_REG_1__SCAN_IN), .S(n6459), .Z(n9131)
         );
  AND2_X1 U8227 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9132) );
  NAND2_X1 U8228 ( .A1(n9131), .A2(n9132), .ZN(n9146) );
  OR2_X1 U8229 ( .A1(n6459), .A2(n6444), .ZN(n9145) );
  NAND2_X1 U8230 ( .A1(n9146), .A2(n9145), .ZN(n6445) );
  NAND2_X1 U8231 ( .A1(n6446), .A2(n6445), .ZN(n9149) );
  INV_X1 U8232 ( .A(n9149), .ZN(n6447) );
  AOI21_X1 U8233 ( .B1(n6461), .B2(P1_REG1_REG_2__SCAN_IN), .A(n6447), .ZN(
        n9167) );
  INV_X1 U8234 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9722) );
  MUX2_X1 U8235 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9722), .S(n9159), .Z(n9166)
         );
  NOR2_X1 U8236 ( .A1(n9167), .A2(n9166), .ZN(n9182) );
  NOR2_X1 U8237 ( .A1(n9159), .A2(n9722), .ZN(n9177) );
  INV_X1 U8238 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6448) );
  MUX2_X1 U8239 ( .A(n6448), .B(P1_REG1_REG_4__SCAN_IN), .S(n9178), .Z(n6449)
         );
  OAI21_X1 U8240 ( .B1(n9182), .B2(n9177), .A(n6449), .ZN(n9197) );
  INV_X1 U8241 ( .A(n9178), .ZN(n6465) );
  NAND2_X1 U8242 ( .A1(n6465), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9196) );
  INV_X1 U8243 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9725) );
  MUX2_X1 U8244 ( .A(n9725), .B(P1_REG1_REG_5__SCAN_IN), .S(n6468), .Z(n9195)
         );
  AOI21_X1 U8245 ( .B1(n9197), .B2(n9196), .A(n9195), .ZN(n9213) );
  NOR2_X1 U8246 ( .A1(n9188), .A2(n9725), .ZN(n9207) );
  INV_X1 U8247 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6450) );
  MUX2_X1 U8248 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6450), .S(n9216), .Z(n6451)
         );
  OAI21_X1 U8249 ( .B1(n9213), .B2(n9207), .A(n6451), .ZN(n9210) );
  NAND2_X1 U8250 ( .A1(n9216), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6484) );
  INV_X1 U8251 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9728) );
  MUX2_X1 U8252 ( .A(n9728), .B(P1_REG1_REG_7__SCAN_IN), .S(n6473), .Z(n6483)
         );
  AOI21_X1 U8253 ( .B1(n9210), .B2(n6484), .A(n6483), .ZN(n6495) );
  AOI21_X1 U8254 ( .B1(n6473), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6495), .ZN(
        n6497) );
  INV_X1 U8255 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9730) );
  MUX2_X1 U8256 ( .A(n9730), .B(P1_REG1_REG_8__SCAN_IN), .S(n6504), .Z(n6496)
         );
  XNOR2_X1 U8257 ( .A(n6497), .B(n6496), .ZN(n6482) );
  AND2_X1 U8258 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7132) );
  INV_X1 U8259 ( .A(n6504), .ZN(n6453) );
  NOR2_X1 U8260 ( .A1(n9189), .A2(n6453), .ZN(n6454) );
  AOI211_X1 U8261 ( .C1(n9215), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n7132), .B(
        n6454), .ZN(n6481) );
  OR2_X1 U8262 ( .A1(n6504), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6456) );
  NAND2_X1 U8263 ( .A1(n6504), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6455) );
  AND2_X1 U8264 ( .A1(n6456), .A2(n6455), .ZN(n6479) );
  INV_X1 U8265 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6457) );
  MUX2_X1 U8266 ( .A(n6457), .B(P1_REG2_REG_2__SCAN_IN), .S(n9151), .Z(n9155)
         );
  INV_X1 U8267 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6458) );
  MUX2_X1 U8268 ( .A(n6458), .B(P1_REG2_REG_1__SCAN_IN), .S(n6459), .Z(n9130)
         );
  NAND2_X1 U8269 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9139) );
  INV_X1 U8270 ( .A(n9139), .ZN(n9129) );
  NAND2_X1 U8271 ( .A1(n9130), .A2(n9129), .ZN(n9128) );
  INV_X1 U8272 ( .A(n6459), .ZN(n9133) );
  NAND2_X1 U8273 ( .A1(n9133), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U8274 ( .A1(n9128), .A2(n6460), .ZN(n9154) );
  NAND2_X1 U8275 ( .A1(n9155), .A2(n9154), .ZN(n9153) );
  NAND2_X1 U8276 ( .A1(n6461), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U8277 ( .A1(n9153), .A2(n6462), .ZN(n9163) );
  MUX2_X1 U8278 ( .A(n5776), .B(P1_REG2_REG_3__SCAN_IN), .S(n9159), .Z(n9164)
         );
  NAND2_X1 U8279 ( .A1(n9163), .A2(n9164), .ZN(n9162) );
  INV_X1 U8280 ( .A(n9159), .ZN(n6463) );
  NAND2_X1 U8281 ( .A1(n6463), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U8282 ( .A1(n9162), .A2(n6464), .ZN(n9176) );
  XNOR2_X1 U8283 ( .A(n9178), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9175) );
  NAND2_X1 U8284 ( .A1(n9176), .A2(n9175), .ZN(n9174) );
  NAND2_X1 U8285 ( .A1(n6465), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U8286 ( .A1(n9174), .A2(n6466), .ZN(n9193) );
  INV_X1 U8287 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6467) );
  XNOR2_X1 U8288 ( .A(n6468), .B(n6467), .ZN(n9194) );
  NAND2_X1 U8289 ( .A1(n9193), .A2(n9194), .ZN(n9192) );
  NAND2_X1 U8290 ( .A1(n6468), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6469) );
  NAND2_X1 U8291 ( .A1(n9192), .A2(n6469), .ZN(n9205) );
  INV_X1 U8292 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6470) );
  MUX2_X1 U8293 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6470), .S(n9216), .Z(n9206)
         );
  NAND2_X1 U8294 ( .A1(n9205), .A2(n9206), .ZN(n9203) );
  NAND2_X1 U8295 ( .A1(n9216), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6471) );
  NAND2_X1 U8296 ( .A1(n9203), .A2(n6471), .ZN(n6490) );
  INV_X1 U8297 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6472) );
  XNOR2_X1 U8298 ( .A(n6473), .B(n6472), .ZN(n6491) );
  NAND2_X1 U8299 ( .A1(n6490), .A2(n6491), .ZN(n6489) );
  NAND2_X1 U8300 ( .A1(n6473), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U8301 ( .A1(n6489), .A2(n6474), .ZN(n6478) );
  AND2_X1 U8302 ( .A1(n6478), .A2(n6479), .ZN(n6503) );
  INV_X1 U8303 ( .A(n6503), .ZN(n6477) );
  OR2_X1 U8304 ( .A1(n6269), .A2(n8095), .ZN(n6475) );
  OAI211_X1 U8305 ( .C1(n6479), .C2(n6478), .A(n6477), .B(n9204), .ZN(n6480)
         );
  OAI211_X1 U8306 ( .C1(n6482), .C2(n9165), .A(n6481), .B(n6480), .ZN(P1_U3251) );
  NAND3_X1 U8307 ( .A1(n9210), .A2(n6484), .A3(n6483), .ZN(n6485) );
  NAND2_X1 U8308 ( .A1(n6485), .A2(n9211), .ZN(n6494) );
  NAND2_X1 U8309 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n6905) );
  INV_X1 U8310 ( .A(n6905), .ZN(n6488) );
  NOR2_X1 U8311 ( .A1(n9189), .A2(n6486), .ZN(n6487) );
  AOI211_X1 U8312 ( .C1(n9215), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n6488), .B(
        n6487), .ZN(n6493) );
  OAI211_X1 U8313 ( .C1(n6491), .C2(n6490), .A(n9204), .B(n6489), .ZN(n6492)
         );
  OAI211_X1 U8314 ( .C1(n6495), .C2(n6494), .A(n6493), .B(n6492), .ZN(P1_U3250) );
  NAND2_X1 U8315 ( .A1(n6504), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6499) );
  OR2_X1 U8316 ( .A1(n6497), .A2(n6496), .ZN(n6498) );
  NAND2_X1 U8317 ( .A1(n6499), .A2(n6498), .ZN(n6502) );
  INV_X1 U8318 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6500) );
  MUX2_X1 U8319 ( .A(n6500), .B(P1_REG1_REG_9__SCAN_IN), .S(n6532), .Z(n6501)
         );
  NOR2_X1 U8320 ( .A1(n6501), .A2(n6502), .ZN(n6533) );
  AOI21_X1 U8321 ( .B1(n6502), .B2(n6501), .A(n6533), .ZN(n6513) );
  AOI21_X1 U8322 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6504), .A(n6503), .ZN(
        n6507) );
  NOR2_X1 U8323 ( .A1(n6532), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6505) );
  AOI21_X1 U8324 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6532), .A(n6505), .ZN(
        n6506) );
  NAND2_X1 U8325 ( .A1(n6506), .A2(n6507), .ZN(n6529) );
  AOI221_X1 U8326 ( .B1(n6507), .B2(n6529), .C1(n6506), .C2(n6529), .A(n7530), 
        .ZN(n6508) );
  INV_X1 U8327 ( .A(n6508), .ZN(n6512) );
  NOR2_X1 U8328 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6509), .ZN(n9047) );
  INV_X1 U8329 ( .A(n6532), .ZN(n6515) );
  NOR2_X1 U8330 ( .A1(n9189), .A2(n6515), .ZN(n6510) );
  AOI211_X1 U8331 ( .C1(n9215), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n9047), .B(
        n6510), .ZN(n6511) );
  OAI211_X1 U8332 ( .C1(n6513), .C2(n9165), .A(n6512), .B(n6511), .ZN(P1_U3252) );
  INV_X1 U8333 ( .A(n6514), .ZN(n6518) );
  OAI222_X1 U8334 ( .A1(n9536), .A2(n6516), .B1(n7754), .B2(n6518), .C1(n6515), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8335 ( .A(n7323), .ZN(n7218) );
  OAI222_X1 U8336 ( .A1(P2_U3151), .A2(n7218), .B1(n8205), .B2(n6518), .C1(
        n6517), .C2(n8968), .ZN(P2_U3286) );
  XOR2_X1 U8337 ( .A(n6520), .B(n6519), .Z(n9140) );
  NAND2_X1 U8338 ( .A1(n9140), .A2(n9109), .ZN(n6523) );
  OR2_X1 U8339 ( .A1(n6521), .A2(P1_U3086), .ZN(n9082) );
  AOI22_X1 U8340 ( .A1(n9102), .A2(n9599), .B1(n9082), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6522) );
  OAI211_X1 U8341 ( .C1(n9119), .C2(n6925), .A(n6523), .B(n6522), .ZN(P1_U3232) );
  INV_X1 U8342 ( .A(n6524), .ZN(n6526) );
  INV_X1 U8343 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6525) );
  OAI222_X1 U8344 ( .A1(P2_U3151), .A2(n7463), .B1(n8205), .B2(n6526), .C1(
        n6525), .C2(n8968), .ZN(P2_U3285) );
  INV_X1 U8345 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6527) );
  INV_X1 U8346 ( .A(n6547), .ZN(n6540) );
  OAI222_X1 U8347 ( .A1(n9536), .A2(n6527), .B1(n7754), .B2(n6526), .C1(n6540), 
        .C2(P1_U3086), .ZN(P1_U3345) );
  NAND2_X1 U8348 ( .A1(n6547), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6528) );
  OAI21_X1 U8349 ( .B1(n6547), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6528), .ZN(
        n6531) );
  OAI21_X1 U8350 ( .B1(n6532), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6529), .ZN(
        n6530) );
  NOR2_X1 U8351 ( .A1(n6531), .A2(n6530), .ZN(n6543) );
  AOI211_X1 U8352 ( .C1(n6531), .C2(n6530), .A(n6543), .B(n7530), .ZN(n6542)
         );
  NOR2_X1 U8353 ( .A1(n6532), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6534) );
  NOR2_X1 U8354 ( .A1(n6534), .A2(n6533), .ZN(n6537) );
  INV_X1 U8355 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6535) );
  MUX2_X1 U8356 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6535), .S(n6547), .Z(n6536)
         );
  NAND2_X1 U8357 ( .A1(n6536), .A2(n6537), .ZN(n6548) );
  OAI211_X1 U8358 ( .C1(n6537), .C2(n6536), .A(n9211), .B(n6548), .ZN(n6539)
         );
  AND2_X1 U8359 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7243) );
  AOI21_X1 U8360 ( .B1(n9215), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7243), .ZN(
        n6538) );
  OAI211_X1 U8361 ( .C1(n9189), .C2(n6540), .A(n6539), .B(n6538), .ZN(n6541)
         );
  OR2_X1 U8362 ( .A1(n6542), .A2(n6541), .ZN(P1_U3253) );
  AOI21_X1 U8363 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n6547), .A(n6543), .ZN(
        n6546) );
  NAND2_X1 U8364 ( .A1(n6782), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6544) );
  OAI21_X1 U8365 ( .B1(n6782), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6544), .ZN(
        n6545) );
  NOR2_X1 U8366 ( .A1(n6546), .A2(n6545), .ZN(n6781) );
  AOI211_X1 U8367 ( .C1(n6546), .C2(n6545), .A(n6781), .B(n7530), .ZN(n6557)
         );
  INV_X1 U8368 ( .A(n6782), .ZN(n6776) );
  NAND2_X1 U8369 ( .A1(n6547), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U8370 ( .A1(n6549), .A2(n6548), .ZN(n6552) );
  INV_X1 U8371 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6550) );
  MUX2_X1 U8372 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6550), .S(n6782), .Z(n6551)
         );
  NAND2_X1 U8373 ( .A1(n6551), .A2(n6552), .ZN(n6775) );
  OAI211_X1 U8374 ( .C1(n6552), .C2(n6551), .A(n6775), .B(n9211), .ZN(n6555)
         );
  NOR2_X1 U8375 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6553), .ZN(n7303) );
  AOI21_X1 U8376 ( .B1(n9215), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7303), .ZN(
        n6554) );
  OAI211_X1 U8377 ( .C1(n9189), .C2(n6776), .A(n6555), .B(n6554), .ZN(n6556)
         );
  OR2_X1 U8378 ( .A1(n6557), .A2(n6556), .ZN(P1_U3254) );
  NAND2_X1 U8379 ( .A1(n9304), .A2(P1_U3973), .ZN(n6558) );
  OAI21_X1 U8380 ( .B1(n5463), .B2(P1_U3973), .A(n6558), .ZN(P1_U3576) );
  NAND2_X1 U8381 ( .A1(n9663), .A2(n9712), .ZN(n6560) );
  INV_X1 U8382 ( .A(n6930), .ZN(n6559) );
  NAND2_X1 U8383 ( .A1(n9127), .A2(n6925), .ZN(n8007) );
  AND2_X1 U8384 ( .A1(n6559), .A2(n8007), .ZN(n7933) );
  INV_X1 U8385 ( .A(n7933), .ZN(n6754) );
  AOI222_X1 U8386 ( .A1(n6560), .A2(n6754), .B1(n6745), .B2(n6744), .C1(n9599), 
        .C2(n9695), .ZN(n9591) );
  NAND2_X1 U8387 ( .A1(n9737), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6562) );
  OAI21_X1 U8388 ( .B1(n9591), .B2(n9737), .A(n6562), .ZN(P1_U3522) );
  INV_X1 U8389 ( .A(n6563), .ZN(n6566) );
  OAI222_X1 U8390 ( .A1(n9536), .A2(n6564), .B1(n7754), .B2(n6566), .C1(
        P1_U3086), .C2(n6776), .ZN(P1_U3344) );
  INV_X1 U8391 ( .A(n7466), .ZN(n7508) );
  OAI222_X1 U8392 ( .A1(n7508), .A2(P2_U3151), .B1(n8205), .B2(n6566), .C1(
        n6565), .C2(n8968), .ZN(P2_U3284) );
  INV_X1 U8393 ( .A(n6567), .ZN(n6568) );
  NAND2_X1 U8394 ( .A1(n6572), .A2(n6568), .ZN(n6570) );
  OR2_X1 U8395 ( .A1(n6677), .A2(n6578), .ZN(n6569) );
  NAND2_X1 U8396 ( .A1(n5198), .A2(n6875), .ZN(n8382) );
  NAND2_X1 U8397 ( .A1(n6571), .A2(n8382), .ZN(n8355) );
  INV_X1 U8398 ( .A(n8355), .ZN(n6591) );
  NAND2_X1 U8399 ( .A1(n6572), .A2(n9930), .ZN(n6575) );
  INV_X1 U8400 ( .A(n6842), .ZN(n6573) );
  AOI22_X1 U8401 ( .A1(n8309), .A2(n6577), .B1(n8303), .B2(n6675), .ZN(n6590)
         );
  INV_X1 U8402 ( .A(n6845), .ZN(n6588) );
  INV_X1 U8403 ( .A(n6578), .ZN(n6580) );
  AOI21_X1 U8404 ( .B1(n6845), .B2(n6580), .A(n6579), .ZN(n6585) );
  INV_X1 U8405 ( .A(n6581), .ZN(n6582) );
  NAND2_X1 U8406 ( .A1(n6583), .A2(n6582), .ZN(n6584) );
  NAND2_X1 U8407 ( .A1(n6585), .A2(n6584), .ZN(n6586) );
  NAND2_X1 U8408 ( .A1(n6586), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6847) );
  OAI211_X1 U8409 ( .C1(n6588), .C2(n6863), .A(n6847), .B(n6587), .ZN(n6803)
         );
  NAND2_X1 U8410 ( .A1(n6803), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6589) );
  OAI211_X1 U8411 ( .C1(n8311), .C2(n6591), .A(n6590), .B(n6589), .ZN(P2_U3172) );
  INV_X1 U8412 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6638) );
  INV_X1 U8413 ( .A(n6592), .ZN(n6631) );
  MUX2_X1 U8414 ( .A(n6889), .B(n5178), .S(n5596), .Z(n6593) );
  XOR2_X1 U8415 ( .A(n6641), .B(n6593), .Z(n6639) );
  INV_X1 U8416 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6615) );
  MUX2_X1 U8417 ( .A(n6615), .B(n6604), .S(n8631), .Z(n6662) );
  AND2_X1 U8418 ( .A1(n6662), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6664) );
  INV_X1 U8419 ( .A(n6641), .ZN(n6594) );
  OAI22_X1 U8420 ( .A1(n6639), .A2(n6664), .B1(n6594), .B2(n6593), .ZN(n6759)
         );
  INV_X1 U8421 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9870) );
  MUX2_X1 U8422 ( .A(n9870), .B(n6603), .S(n8631), .Z(n6595) );
  XNOR2_X1 U8423 ( .A(n6595), .B(n4353), .ZN(n6758) );
  INV_X1 U8424 ( .A(n6595), .ZN(n6596) );
  AOI22_X1 U8425 ( .A1(n6759), .A2(n6758), .B1(n4353), .B2(n6596), .ZN(n9751)
         );
  INV_X4 U8426 ( .A(n8664), .ZN(n8631) );
  MUX2_X1 U8427 ( .A(n6598), .B(n6597), .S(n8631), .Z(n6599) );
  XNOR2_X1 U8428 ( .A(n6599), .B(n9745), .ZN(n9750) );
  NAND2_X1 U8429 ( .A1(n9751), .A2(n9750), .ZN(n9749) );
  NAND2_X1 U8430 ( .A1(n6599), .A2(n4938), .ZN(n6600) );
  AND2_X1 U8431 ( .A1(n9749), .A2(n6600), .ZN(n6602) );
  MUX2_X1 U8432 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8631), .Z(n6685) );
  XOR2_X1 U8433 ( .A(n6707), .B(n6685), .Z(n6601) );
  NAND3_X1 U8434 ( .A1(n9749), .A2(n6600), .A3(n6601), .ZN(n6686) );
  OAI211_X1 U8435 ( .C1(n6602), .C2(n6601), .A(n9832), .B(n6686), .ZN(n6637)
         );
  XNOR2_X1 U8436 ( .A(n4353), .B(n6603), .ZN(n6765) );
  NOR2_X1 U8437 ( .A1(n6604), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U8438 ( .A1(n5207), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6606) );
  OAI21_X1 U8439 ( .B1(n6641), .B2(n6605), .A(n6606), .ZN(n6644) );
  NAND2_X1 U8440 ( .A1(n6642), .A2(n6606), .ZN(n6764) );
  NAND2_X1 U8441 ( .A1(n6765), .A2(n6764), .ZN(n6763) );
  NAND2_X1 U8442 ( .A1(n4353), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6607) );
  XNOR2_X1 U8443 ( .A(n6707), .B(n6609), .ZN(n6611) );
  NAND2_X1 U8444 ( .A1(n6610), .A2(n6611), .ZN(n6698) );
  INV_X1 U8445 ( .A(n6611), .ZN(n6613) );
  NAND3_X1 U8446 ( .A1(n9753), .A2(n6613), .A3(n6612), .ZN(n6614) );
  AND2_X1 U8447 ( .A1(n6698), .A2(n6614), .ZN(n6625) );
  OR2_X1 U8448 ( .A1(n5595), .A2(P2_U3151), .ZN(n8965) );
  NOR2_X1 U8449 ( .A1(n6626), .A2(n8965), .ZN(n6665) );
  NOR2_X1 U8450 ( .A1(n6615), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U8451 ( .A1(n5207), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6617) );
  NAND2_X1 U8452 ( .A1(n6762), .A2(n6761), .ZN(n6760) );
  NAND2_X1 U8453 ( .A1(n4353), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6618) );
  NAND2_X1 U8454 ( .A1(n9743), .A2(n6621), .ZN(n6619) );
  INV_X1 U8455 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7016) );
  XNOR2_X1 U8456 ( .A(n6707), .B(n7016), .ZN(n6620) );
  NAND2_X1 U8457 ( .A1(n6619), .A2(n6620), .ZN(n6709) );
  INV_X1 U8458 ( .A(n6620), .ZN(n6622) );
  NAND3_X1 U8459 ( .A1(n9743), .A2(n6622), .A3(n6621), .ZN(n6623) );
  AND2_X1 U8460 ( .A1(n6709), .A2(n6623), .ZN(n6624) );
  OAI22_X1 U8461 ( .A1(n6625), .A2(n9825), .B1(n9829), .B2(n6624), .ZN(n6635)
         );
  INV_X1 U8462 ( .A(n6626), .ZN(n6629) );
  NOR2_X1 U8463 ( .A1(n8631), .A2(P2_U3151), .ZN(n6627) );
  AND2_X1 U8464 ( .A1(n5595), .A2(n6627), .ZN(n6628) );
  NAND2_X1 U8465 ( .A1(n6629), .A2(n6628), .ZN(n6633) );
  INV_X1 U8466 ( .A(n8965), .ZN(n6630) );
  NAND2_X1 U8467 ( .A1(n6631), .A2(n6630), .ZN(n6632) );
  NAND2_X1 U8468 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6943) );
  OAI21_X1 U8469 ( .B1(n9835), .B2(n6707), .A(n6943), .ZN(n6634) );
  NOR2_X1 U8470 ( .A1(n6635), .A2(n6634), .ZN(n6636) );
  OAI211_X1 U8471 ( .C1(n6638), .C2(n9783), .A(n6637), .B(n6636), .ZN(P2_U3186) );
  XNOR2_X1 U8472 ( .A(n6639), .B(n6664), .ZN(n6653) );
  INV_X1 U8473 ( .A(n9832), .ZN(n7512) );
  OAI22_X1 U8474 ( .A1(n9835), .A2(n6641), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6640), .ZN(n6651) );
  INV_X1 U8475 ( .A(n6642), .ZN(n6643) );
  AOI21_X1 U8476 ( .B1(n5178), .B2(n6644), .A(n6643), .ZN(n6649) );
  INV_X1 U8477 ( .A(n6645), .ZN(n6646) );
  AOI21_X1 U8478 ( .B1(n6889), .B2(n6647), .A(n6646), .ZN(n6648) );
  OAI22_X1 U8479 ( .A1(n6649), .A2(n9825), .B1(n9829), .B2(n6648), .ZN(n6650)
         );
  AOI211_X1 U8480 ( .C1(n9818), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6651), .B(
        n6650), .ZN(n6652) );
  OAI21_X1 U8481 ( .B1(n6653), .B2(n7512), .A(n6652), .ZN(P2_U3183) );
  INV_X1 U8482 ( .A(n6654), .ZN(n6671) );
  AOI22_X1 U8483 ( .A1(n7580), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n6683), .ZN(n6655) );
  OAI21_X1 U8484 ( .B1(n6671), .B2(n8205), .A(n6655), .ZN(P2_U3283) );
  INV_X1 U8485 ( .A(n6656), .ZN(n7013) );
  OAI21_X1 U8486 ( .B1(n9851), .B2(n9919), .A(n8355), .ZN(n6657) );
  NAND2_X1 U8487 ( .A1(n6675), .A2(n9853), .ZN(n6864) );
  OAI211_X1 U8488 ( .C1(n6875), .C2(n9913), .A(n6657), .B(n6864), .ZN(n6659)
         );
  NAND2_X1 U8489 ( .A1(n6659), .A2(n9947), .ZN(n6658) );
  OAI21_X1 U8490 ( .B1(n9947), .B2(n6604), .A(n6658), .ZN(P2_U3459) );
  INV_X1 U8491 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U8492 ( .A1(n9931), .A2(n6659), .ZN(n6660) );
  OAI21_X1 U8493 ( .B1(n9931), .B2(n6661), .A(n6660), .ZN(P2_U3390) );
  INV_X1 U8494 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6670) );
  INV_X1 U8495 ( .A(n9835), .ZN(n8600) );
  NOR2_X1 U8496 ( .A1(n6662), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6663) );
  OAI22_X1 U8497 ( .A1(n6665), .A2(n9832), .B1(n6664), .B2(n6663), .ZN(n6666)
         );
  OAI21_X1 U8498 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6667), .A(n6666), .ZN(n6668) );
  AOI21_X1 U8499 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n8600), .A(n6668), .ZN(n6669) );
  OAI21_X1 U8500 ( .B1(n9783), .B2(n6670), .A(n6669), .ZN(P2_U3182) );
  INV_X1 U8501 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6672) );
  INV_X1 U8502 ( .A(n6808), .ZN(n6812) );
  OAI222_X1 U8503 ( .A1(n9536), .A2(n6672), .B1(n7754), .B2(n6671), .C1(n6812), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  NAND2_X1 U8504 ( .A1(n6673), .A2(n8381), .ZN(n6674) );
  XOR2_X1 U8505 ( .A(n6800), .B(n6799), .Z(n6681) );
  INV_X1 U8506 ( .A(n8309), .ZN(n8326) );
  OR3_X1 U8507 ( .A1(n6677), .A2(n6863), .A3(n6676), .ZN(n8306) );
  AOI22_X1 U8508 ( .A1(n8319), .A2(n5198), .B1(n8303), .B2(n9837), .ZN(n6678)
         );
  OAI21_X1 U8509 ( .B1(n8326), .B2(n9872), .A(n6678), .ZN(n6679) );
  AOI21_X1 U8510 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6803), .A(n6679), .ZN(
        n6680) );
  OAI21_X1 U8511 ( .B1(n6681), .B2(n8311), .A(n6680), .ZN(P2_U3162) );
  INV_X1 U8512 ( .A(n6682), .ZN(n6737) );
  AOI22_X1 U8513 ( .A1(n8604), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n6683), .ZN(n6684) );
  OAI21_X1 U8514 ( .B1(n6737), .B2(n8205), .A(n6684), .ZN(P2_U3282) );
  INV_X1 U8515 ( .A(n6707), .ZN(n6688) );
  INV_X1 U8516 ( .A(n6685), .ZN(n6687) );
  OAI21_X1 U8517 ( .B1(n6688), .B2(n6687), .A(n6686), .ZN(n6722) );
  MUX2_X1 U8518 ( .A(n6690), .B(n6689), .S(n8631), .Z(n6691) );
  XNOR2_X1 U8519 ( .A(n6691), .B(n6730), .ZN(n6723) );
  INV_X1 U8520 ( .A(n6691), .ZN(n6692) );
  AOI22_X1 U8521 ( .A1(n6722), .A2(n6723), .B1(n6692), .B2(n6730), .ZN(n6695)
         );
  MUX2_X1 U8522 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8631), .Z(n6693) );
  NOR2_X1 U8523 ( .A1(n6693), .A2(n6832), .ZN(n6824) );
  AOI21_X1 U8524 ( .B1(n6693), .B2(n6832), .A(n6824), .ZN(n6694) );
  NAND2_X1 U8525 ( .A1(n6695), .A2(n6694), .ZN(n6826) );
  OAI21_X1 U8526 ( .B1(n6695), .B2(n6694), .A(n6826), .ZN(n6696) );
  NAND2_X1 U8527 ( .A1(n6696), .A2(n9832), .ZN(n6721) );
  INV_X1 U8528 ( .A(n9825), .ZN(n7343) );
  NAND2_X1 U8529 ( .A1(n6707), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8530 ( .A1(n6698), .A2(n6697), .ZN(n6699) );
  OR2_X1 U8531 ( .A1(n6699), .A2(n6730), .ZN(n6700) );
  NAND2_X1 U8532 ( .A1(n6699), .A2(n6730), .ZN(n6703) );
  NAND2_X1 U8533 ( .A1(n6726), .A2(n6703), .ZN(n6701) );
  INV_X1 U8534 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9939) );
  MUX2_X1 U8535 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9939), .S(n6832), .Z(n6702)
         );
  INV_X1 U8536 ( .A(n6702), .ZN(n6704) );
  NAND3_X1 U8537 ( .A1(n6726), .A2(n6704), .A3(n6703), .ZN(n6705) );
  NAND2_X1 U8538 ( .A1(n6834), .A2(n6705), .ZN(n6719) );
  INV_X1 U8539 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10165) );
  NOR2_X1 U8540 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10165), .ZN(n7178) );
  INV_X1 U8541 ( .A(n7178), .ZN(n6706) );
  OAI21_X1 U8542 ( .B1(n9835), .B2(n6832), .A(n6706), .ZN(n6718) );
  INV_X1 U8543 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6716) );
  NAND2_X1 U8544 ( .A1(n6707), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U8545 ( .A1(n6709), .A2(n6708), .ZN(n6710) );
  NAND2_X1 U8546 ( .A1(n6710), .A2(n6730), .ZN(n6711) );
  MUX2_X1 U8547 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7195), .S(n6832), .Z(n6712)
         );
  NOR2_X1 U8548 ( .A1(n4504), .A2(n6712), .ZN(n6714) );
  INV_X1 U8549 ( .A(n6821), .ZN(n6713) );
  AOI21_X1 U8550 ( .B1(n6714), .B2(n6724), .A(n6713), .ZN(n6715) );
  OAI22_X1 U8551 ( .A1(n9783), .A2(n6716), .B1(n9829), .B2(n6715), .ZN(n6717)
         );
  AOI211_X1 U8552 ( .C1(n7343), .C2(n6719), .A(n6718), .B(n6717), .ZN(n6720)
         );
  NAND2_X1 U8553 ( .A1(n6721), .A2(n6720), .ZN(P2_U3188) );
  XOR2_X1 U8554 ( .A(n6723), .B(n6722), .Z(n6735) );
  INV_X1 U8555 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6733) );
  INV_X1 U8556 ( .A(n9829), .ZN(n7470) );
  OAI21_X1 U8557 ( .B1(n6725), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6724), .ZN(
        n6729) );
  OAI21_X1 U8558 ( .B1(n6727), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6726), .ZN(
        n6728) );
  AOI22_X1 U8559 ( .A1(n7470), .A2(n6729), .B1(n7343), .B2(n6728), .ZN(n6732)
         );
  AND2_X1 U8560 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7074) );
  AOI21_X1 U8561 ( .B1(n8600), .B2(n4828), .A(n7074), .ZN(n6731) );
  OAI211_X1 U8562 ( .C1(n6733), .C2(n9783), .A(n6732), .B(n6731), .ZN(n6734)
         );
  AOI21_X1 U8563 ( .B1(n6735), .B2(n9832), .A(n6734), .ZN(n6736) );
  INV_X1 U8564 ( .A(n6736), .ZN(P2_U3187) );
  INV_X1 U8565 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6738) );
  INV_X1 U8566 ( .A(n7003), .ZN(n6997) );
  OAI222_X1 U8567 ( .A1(n9536), .A2(n6738), .B1(n7754), .B2(n6737), .C1(
        P1_U3086), .C2(n6997), .ZN(P1_U3342) );
  INV_X1 U8568 ( .A(n9599), .ZN(n6757) );
  NAND3_X1 U8569 ( .A1(n6741), .A2(n6740), .A3(n6739), .ZN(n6743) );
  INV_X1 U8570 ( .A(n9402), .ZN(n9573) );
  AND2_X1 U8571 ( .A1(n6744), .A2(n8063), .ZN(n6746) );
  OAI21_X1 U8572 ( .B1(n6926), .B2(n6746), .A(n6745), .ZN(n6747) );
  NOR2_X1 U8573 ( .A1(n6748), .A2(n6747), .ZN(n6751) );
  INV_X1 U8574 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6749) );
  NOR2_X1 U8575 ( .A1(n9393), .A2(n6749), .ZN(n6750) );
  AOI211_X1 U8576 ( .C1(n9573), .C2(P1_REG3_REG_0__SCAN_IN), .A(n6751), .B(
        n6750), .ZN(n6756) );
  NAND4_X1 U8577 ( .A1(n6754), .A2(n9393), .A3(n6753), .A4(n6752), .ZN(n6755)
         );
  OAI211_X1 U8578 ( .C1(n6757), .C2(n9407), .A(n6756), .B(n6755), .ZN(P1_U3293) );
  XNOR2_X1 U8579 ( .A(n6759), .B(n6758), .ZN(n6773) );
  OAI21_X1 U8580 ( .B1(n6762), .B2(n6761), .A(n6760), .ZN(n6767) );
  OAI21_X1 U8581 ( .B1(n6765), .B2(n6764), .A(n6763), .ZN(n6766) );
  AOI22_X1 U8582 ( .A1(n7470), .A2(n6767), .B1(n7343), .B2(n6766), .ZN(n6769)
         );
  NAND2_X1 U8583 ( .A1(P2_U3151), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6768) );
  OAI211_X1 U8584 ( .C1(n9835), .C2(n4353), .A(n6769), .B(n6768), .ZN(n6771)
         );
  AOI21_X1 U8585 ( .B1(n9818), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n6771), .ZN(
        n6772) );
  OAI21_X1 U8586 ( .B1(n6773), .B2(n7512), .A(n6772), .ZN(P2_U3184) );
  INV_X1 U8587 ( .A(n9189), .ZN(n9217) );
  INV_X1 U8588 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6774) );
  MUX2_X1 U8589 ( .A(n6774), .B(P1_REG1_REG_12__SCAN_IN), .S(n6808), .Z(n6778)
         );
  OAI21_X1 U8590 ( .B1(n6776), .B2(n6550), .A(n6775), .ZN(n6777) );
  NOR2_X1 U8591 ( .A1(n6777), .A2(n6778), .ZN(n6811) );
  AOI21_X1 U8592 ( .B1(n6778), .B2(n6777), .A(n6811), .ZN(n6780) );
  NAND2_X1 U8593 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7476) );
  NAND2_X1 U8594 ( .A1(n9215), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6779) );
  OAI211_X1 U8595 ( .C1(n9165), .C2(n6780), .A(n7476), .B(n6779), .ZN(n6787)
         );
  AOI21_X1 U8596 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6782), .A(n6781), .ZN(
        n6785) );
  NOR2_X1 U8597 ( .A1(n6808), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6783) );
  AOI21_X1 U8598 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n6808), .A(n6783), .ZN(
        n6784) );
  NAND2_X1 U8599 ( .A1(n6784), .A2(n6785), .ZN(n6807) );
  AOI221_X1 U8600 ( .B1(n6785), .B2(n6807), .C1(n6784), .C2(n6807), .A(n7530), 
        .ZN(n6786) );
  AOI211_X1 U8601 ( .C1(n9217), .C2(n6808), .A(n6787), .B(n6786), .ZN(n6788)
         );
  INV_X1 U8602 ( .A(n6788), .ZN(P1_U3255) );
  OAI21_X1 U8603 ( .B1(n6791), .B2(n6790), .A(n6789), .ZN(n6796) );
  AOI22_X1 U8604 ( .A1(n9058), .A2(n6792), .B1(n9116), .B2(n9125), .ZN(n6794)
         );
  AND2_X1 U8605 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9161) );
  AOI21_X1 U8606 ( .B1(n9102), .B2(n9124), .A(n9161), .ZN(n6793) );
  OAI211_X1 U8607 ( .C1(n6991), .C2(n9119), .A(n6794), .B(n6793), .ZN(n6795)
         );
  AOI21_X1 U8608 ( .B1(n6796), .B2(n9109), .A(n6795), .ZN(n6797) );
  INV_X1 U8609 ( .A(n6797), .ZN(P1_U3218) );
  XNOR2_X1 U8610 ( .A(n6848), .B(n9837), .ZN(n6851) );
  XOR2_X1 U8611 ( .A(n6852), .B(n6851), .Z(n6805) );
  AOI22_X1 U8612 ( .A1(n8319), .A2(n6675), .B1(n8303), .B2(n9854), .ZN(n6801)
         );
  OAI21_X1 U8613 ( .B1(n8326), .B2(n9861), .A(n6801), .ZN(n6802) );
  AOI21_X1 U8614 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6803), .A(n6802), .ZN(
        n6804) );
  OAI21_X1 U8615 ( .B1(n6805), .B2(n8311), .A(n6804), .ZN(P2_U3177) );
  NAND2_X1 U8616 ( .A1(n7003), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6806) );
  OAI21_X1 U8617 ( .B1(n7003), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6806), .ZN(
        n6810) );
  OAI21_X1 U8618 ( .B1(n6808), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6807), .ZN(
        n6809) );
  NOR2_X1 U8619 ( .A1(n6810), .A2(n6809), .ZN(n7002) );
  AOI211_X1 U8620 ( .C1(n6810), .C2(n6809), .A(n7002), .B(n7530), .ZN(n6819)
         );
  AOI21_X1 U8621 ( .B1(n6812), .B2(n6774), .A(n6811), .ZN(n6815) );
  INV_X1 U8622 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6813) );
  MUX2_X1 U8623 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6813), .S(n7003), .Z(n6814)
         );
  NAND2_X1 U8624 ( .A1(n6814), .A2(n6815), .ZN(n6996) );
  OAI211_X1 U8625 ( .C1(n6815), .C2(n6814), .A(n9211), .B(n6996), .ZN(n6817)
         );
  AND2_X1 U8626 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7410) );
  AOI21_X1 U8627 ( .B1(n9215), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7410), .ZN(
        n6816) );
  OAI211_X1 U8628 ( .C1(n9189), .C2(n6997), .A(n6817), .B(n6816), .ZN(n6818)
         );
  OR2_X1 U8629 ( .A1(n6819), .A2(n6818), .ZN(P1_U3256) );
  NAND2_X1 U8630 ( .A1(n6832), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6820) );
  AOI21_X1 U8631 ( .B1(n6828), .B2(n6823), .A(n9763), .ZN(n6841) );
  INV_X1 U8632 ( .A(n6824), .ZN(n6825) );
  NAND2_X1 U8633 ( .A1(n6826), .A2(n6825), .ZN(n6830) );
  MUX2_X1 U8634 ( .A(n6828), .B(n6827), .S(n8631), .Z(n7223) );
  XNOR2_X1 U8635 ( .A(n7223), .B(n7225), .ZN(n6829) );
  NAND2_X1 U8636 ( .A1(n6830), .A2(n6829), .ZN(n7224) );
  OAI21_X1 U8637 ( .B1(n6830), .B2(n6829), .A(n7224), .ZN(n6831) );
  NAND2_X1 U8638 ( .A1(n6831), .A2(n9832), .ZN(n6840) );
  NAND2_X1 U8639 ( .A1(n6832), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6833) );
  OAI21_X1 U8640 ( .B1(n4451), .B2(P2_REG1_REG_7__SCAN_IN), .A(n9769), .ZN(
        n6838) );
  INV_X1 U8641 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n9964) );
  INV_X1 U8642 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10163) );
  NOR2_X1 U8643 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10163), .ZN(n7205) );
  AOI21_X1 U8644 ( .B1(n8600), .B2(n4934), .A(n7205), .ZN(n6836) );
  OAI21_X1 U8645 ( .B1(n9964), .B2(n9783), .A(n6836), .ZN(n6837) );
  AOI21_X1 U8646 ( .B1(n7343), .B2(n6838), .A(n6837), .ZN(n6839) );
  OAI211_X1 U8647 ( .C1(n6841), .C2(n9829), .A(n6840), .B(n6839), .ZN(P2_U3189) );
  NOR2_X1 U8648 ( .A1(n6842), .A2(n6863), .ZN(n8569) );
  OR2_X1 U8649 ( .A1(n6843), .A2(P2_U3151), .ZN(n8571) );
  INV_X1 U8650 ( .A(n8571), .ZN(n6844) );
  AOI21_X1 U8651 ( .B1(n6845), .B2(n8569), .A(n6844), .ZN(n6846) );
  INV_X1 U8652 ( .A(n8323), .ZN(n7727) );
  INV_X1 U8653 ( .A(n9837), .ZN(n6849) );
  XNOR2_X1 U8654 ( .A(n8170), .B(n9883), .ZN(n6939) );
  XNOR2_X1 U8655 ( .A(n6939), .B(n9854), .ZN(n6853) );
  OAI211_X1 U8656 ( .C1(n6854), .C2(n6853), .A(n6938), .B(n8316), .ZN(n6858)
         );
  INV_X1 U8657 ( .A(n9838), .ZN(n7085) );
  NAND2_X1 U8658 ( .A1(n8319), .A2(n9837), .ZN(n6855) );
  NAND2_X1 U8659 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3151), .ZN(n9759) );
  OAI211_X1 U8660 ( .C1(n7085), .C2(n8321), .A(n6855), .B(n9759), .ZN(n6856)
         );
  AOI21_X1 U8661 ( .B1(n9883), .B2(n8309), .A(n6856), .ZN(n6857) );
  OAI211_X1 U8662 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7727), .A(n6858), .B(
        n6857), .ZN(P2_U3158) );
  INV_X1 U8663 ( .A(n6859), .ZN(n6862) );
  INV_X1 U8664 ( .A(n7139), .ZN(n7143) );
  OAI222_X1 U8665 ( .A1(n9536), .A2(n6860), .B1(n7754), .B2(n6862), .C1(
        P1_U3086), .C2(n7143), .ZN(P1_U3341) );
  OAI222_X1 U8666 ( .A1(n9800), .A2(P2_U3151), .B1(n8205), .B2(n6862), .C1(
        n6861), .C2(n8968), .ZN(P2_U3281) );
  NAND3_X1 U8667 ( .A1(n8355), .A2(n9913), .A3(n6863), .ZN(n6865) );
  NAND2_X1 U8668 ( .A1(n6865), .A2(n6864), .ZN(n6873) );
  OR2_X1 U8669 ( .A1(n5622), .A2(n6866), .ZN(n6871) );
  OR2_X1 U8670 ( .A1(n6868), .A2(n6867), .ZN(n6870) );
  NAND2_X1 U8671 ( .A1(n5622), .A2(n6868), .ZN(n6869) );
  NAND4_X1 U8672 ( .A1(n6872), .A2(n6871), .A3(n6870), .A4(n6869), .ZN(n6874)
         );
  MUX2_X1 U8673 ( .A(n6873), .B(P2_REG2_REG_0__SCAN_IN), .S(n9871), .Z(n6877)
         );
  OAI22_X1 U8674 ( .A1(n8807), .A2(n6875), .B1(n6667), .B2(n9862), .ZN(n6876)
         );
  OR2_X1 U8675 ( .A1(n6877), .A2(n6876), .ZN(P2_U3233) );
  INV_X1 U8676 ( .A(n6879), .ZN(n6880) );
  AOI21_X1 U8677 ( .B1(n6571), .B2(n6878), .A(n6880), .ZN(n9874) );
  AOI22_X1 U8678 ( .A1(n9855), .A2(n5198), .B1(n9837), .B2(n9853), .ZN(n6884)
         );
  OAI21_X1 U8679 ( .B1(n6881), .B2(n6878), .A(n9848), .ZN(n6882) );
  NAND2_X1 U8680 ( .A1(n6882), .A2(n9851), .ZN(n6883) );
  OAI211_X1 U8681 ( .C1(n9874), .C2(n7013), .A(n6884), .B(n6883), .ZN(n9876)
         );
  OR2_X1 U8682 ( .A1(n8562), .A2(n8375), .ZN(n8691) );
  NOR2_X1 U8683 ( .A1(n9874), .A2(n8691), .ZN(n6885) );
  OAI21_X1 U8684 ( .B1(n9876), .B2(n6885), .A(n9868), .ZN(n6888) );
  AOI22_X1 U8685 ( .A1(n9842), .A2(n6886), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9843), .ZN(n6887) );
  OAI211_X1 U8686 ( .C1(n9868), .C2(n6889), .A(n6888), .B(n6887), .ZN(P2_U3232) );
  OR2_X1 U8687 ( .A1(n6956), .A2(n6957), .ZN(n6954) );
  NAND2_X1 U8688 ( .A1(n6954), .A2(n6890), .ZN(n6894) );
  XNOR2_X1 U8689 ( .A(n6892), .B(n6891), .ZN(n6893) );
  XNOR2_X1 U8690 ( .A(n6894), .B(n6893), .ZN(n6899) );
  AOI22_X1 U8691 ( .A1(n9058), .A2(n6975), .B1(n9081), .B2(n9124), .ZN(n6895)
         );
  NAND2_X1 U8692 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9187) );
  OAI211_X1 U8693 ( .C1(n6896), .C2(n9113), .A(n6895), .B(n9187), .ZN(n6897)
         );
  AOI21_X1 U8694 ( .B1(n6976), .B2(n9084), .A(n6897), .ZN(n6898) );
  OAI21_X1 U8695 ( .B1(n6899), .B2(n9075), .A(n6898), .ZN(P1_U3227) );
  NAND2_X1 U8696 ( .A1(n9126), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6900) );
  OAI21_X1 U8697 ( .B1(n9421), .B2(n9126), .A(n6900), .ZN(P1_U3583) );
  XOR2_X1 U8698 ( .A(n6902), .B(n6901), .Z(n6903) );
  XNOR2_X1 U8699 ( .A(n6904), .B(n6903), .ZN(n6909) );
  AOI22_X1 U8700 ( .A1(n9058), .A2(n7064), .B1(n9116), .B2(n9639), .ZN(n6906)
         );
  OAI211_X1 U8701 ( .C1(n7067), .C2(n9113), .A(n6906), .B(n6905), .ZN(n6907)
         );
  AOI21_X1 U8702 ( .B1(n4352), .B2(n9084), .A(n6907), .ZN(n6908) );
  OAI21_X1 U8703 ( .B1(n6909), .B2(n9075), .A(n6908), .ZN(P1_U3213) );
  NAND2_X1 U8704 ( .A1(n6911), .A2(n6910), .ZN(n6916) );
  OR2_X1 U8705 ( .A1(n6956), .A2(n6912), .ZN(n6914) );
  NAND2_X1 U8706 ( .A1(n6914), .A2(n6913), .ZN(n6915) );
  XOR2_X1 U8707 ( .A(n6916), .B(n6915), .Z(n6922) );
  AOI22_X1 U8708 ( .A1(n9058), .A2(n9572), .B1(n9081), .B2(n9617), .ZN(n6918)
         );
  AND2_X1 U8709 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9214) );
  INV_X1 U8710 ( .A(n9214), .ZN(n6917) );
  OAI211_X1 U8711 ( .C1(n6919), .C2(n9113), .A(n6918), .B(n6917), .ZN(n6920)
         );
  AOI21_X1 U8712 ( .B1(n9577), .B2(n9084), .A(n6920), .ZN(n6921) );
  OAI21_X1 U8713 ( .B1(n6922), .B2(n9075), .A(n6921), .ZN(P1_U3239) );
  XOR2_X1 U8714 ( .A(n6924), .B(n6923), .Z(n6934) );
  INV_X1 U8715 ( .A(n6934), .ZN(n9596) );
  NOR2_X1 U8716 ( .A1(n9571), .A2(n6971), .ZN(n9564) );
  NOR2_X2 U8717 ( .A1(n9571), .A2(n8108), .ZN(n9585) );
  OAI211_X1 U8718 ( .C1(n9593), .C2(n6925), .A(n9581), .B(n7027), .ZN(n9592)
         );
  INV_X1 U8719 ( .A(n6926), .ZN(n6927) );
  NOR2_X2 U8720 ( .A1(n9571), .A2(n6927), .ZN(n9578) );
  AOI22_X1 U8721 ( .A1(n9578), .A2(n7792), .B1(n9573), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6928) );
  OAI21_X1 U8722 ( .B1(n9331), .B2(n9592), .A(n6928), .ZN(n6936) );
  AOI22_X1 U8723 ( .A1(n9659), .A2(n9127), .B1(n9125), .B2(n9695), .ZN(n6933)
         );
  OAI21_X1 U8724 ( .B1(n6930), .B2(n6923), .A(n6929), .ZN(n6931) );
  NAND2_X1 U8725 ( .A1(n6931), .A2(n9666), .ZN(n6932) );
  OAI211_X1 U8726 ( .C1(n6934), .C2(n9647), .A(n6933), .B(n6932), .ZN(n9594)
         );
  MUX2_X1 U8727 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9594), .S(n9393), .Z(n6935)
         );
  AOI211_X1 U8728 ( .C1(n9596), .C2(n9564), .A(n6936), .B(n6935), .ZN(n6937)
         );
  INV_X1 U8729 ( .A(n6937), .ZN(P1_U3292) );
  XNOR2_X1 U8730 ( .A(n7018), .B(n4473), .ZN(n7072) );
  XNOR2_X1 U8731 ( .A(n7072), .B(n9838), .ZN(n6941) );
  INV_X1 U8732 ( .A(n9854), .ZN(n6944) );
  AOI21_X1 U8733 ( .B1(n6941), .B2(n6940), .A(n4452), .ZN(n6949) );
  INV_X1 U8734 ( .A(n6942), .ZN(n7017) );
  OAI21_X1 U8735 ( .B1(n6944), .B2(n8306), .A(n6943), .ZN(n6945) );
  AOI21_X1 U8736 ( .B1(n8303), .B2(n8587), .A(n6945), .ZN(n6946) );
  OAI21_X1 U8737 ( .B1(n9889), .B2(n8326), .A(n6946), .ZN(n6947) );
  AOI21_X1 U8738 ( .B1(n7017), .B2(n8323), .A(n6947), .ZN(n6948) );
  OAI21_X1 U8739 ( .B1(n6949), .B2(n8311), .A(n6948), .ZN(P2_U3170) );
  INV_X1 U8740 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6951) );
  INV_X1 U8741 ( .A(n6950), .ZN(n6953) );
  INV_X1 U8742 ( .A(n7382), .ZN(n7389) );
  OAI222_X1 U8743 ( .A1(n9536), .A2(n6951), .B1(n7754), .B2(n6953), .C1(n7389), 
        .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U8744 ( .A(n8642), .ZN(n8625) );
  INV_X1 U8745 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6952) );
  OAI222_X1 U8746 ( .A1(P2_U3151), .A2(n8625), .B1(n8205), .B2(n6953), .C1(
        n6952), .C2(n8968), .ZN(P2_U3280) );
  INV_X1 U8747 ( .A(n6954), .ZN(n6955) );
  AOI211_X1 U8748 ( .C1(n6957), .C2(n6956), .A(n9075), .B(n6955), .ZN(n6962)
         );
  INV_X1 U8749 ( .A(n6958), .ZN(n7045) );
  AOI22_X1 U8750 ( .A1(n9058), .A2(n7045), .B1(n9116), .B2(n9598), .ZN(n6960)
         );
  AND2_X1 U8751 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9173) );
  AOI21_X1 U8752 ( .B1(n9102), .B2(n9617), .A(n9173), .ZN(n6959) );
  OAI211_X1 U8753 ( .C1(n7047), .C2(n9119), .A(n6960), .B(n6959), .ZN(n6961)
         );
  OR2_X1 U8754 ( .A1(n6962), .A2(n6961), .ZN(P1_U3230) );
  NAND3_X1 U8755 ( .A1(n6963), .A2(n7810), .A3(n7053), .ZN(n6964) );
  NAND2_X1 U8756 ( .A1(n6965), .A2(n6964), .ZN(n6966) );
  NAND2_X1 U8757 ( .A1(n6966), .A2(n9666), .ZN(n6968) );
  AOI22_X1 U8758 ( .A1(n9659), .A2(n9124), .B1(n9639), .B2(n9695), .ZN(n6967)
         );
  NAND2_X1 U8759 ( .A1(n6968), .A2(n6967), .ZN(n9629) );
  INV_X1 U8760 ( .A(n9629), .ZN(n6981) );
  NAND2_X1 U8761 ( .A1(n6970), .A2(n6969), .ZN(n7054) );
  XNOR2_X1 U8762 ( .A(n7054), .B(n7053), .ZN(n9624) );
  AND2_X1 U8763 ( .A1(n9647), .A2(n6971), .ZN(n6972) );
  NAND2_X1 U8764 ( .A1(n7043), .A2(n6976), .ZN(n6973) );
  NAND2_X1 U8765 ( .A1(n6973), .A2(n9581), .ZN(n6974) );
  OR2_X1 U8766 ( .A1(n6974), .A2(n9583), .ZN(n9625) );
  AOI22_X1 U8767 ( .A1(n9571), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6975), .B2(
        n9573), .ZN(n6978) );
  NAND2_X1 U8768 ( .A1(n9578), .A2(n6976), .ZN(n6977) );
  OAI211_X1 U8769 ( .C1(n9625), .C2(n9331), .A(n6978), .B(n6977), .ZN(n6979)
         );
  AOI21_X1 U8770 ( .B1(n9624), .B2(n9586), .A(n6979), .ZN(n6980) );
  OAI21_X1 U8771 ( .B1(n6981), .B2(n9571), .A(n6980), .ZN(P1_U3288) );
  INV_X1 U8772 ( .A(n6982), .ZN(n6985) );
  OAI222_X1 U8773 ( .A1(P2_U3151), .A2(n9817), .B1(n8205), .B2(n6985), .C1(
        n6983), .C2(n8968), .ZN(P2_U3279) );
  INV_X1 U8774 ( .A(n7398), .ZN(n7386) );
  OAI222_X1 U8775 ( .A1(P1_U3086), .A2(n7386), .B1(n7754), .B2(n6985), .C1(
        n6984), .C2(n9536), .ZN(P1_U3339) );
  XNOR2_X1 U8776 ( .A(n6986), .B(n6987), .ZN(n9612) );
  OAI21_X1 U8777 ( .B1(n7796), .B2(n6987), .A(n7035), .ZN(n6988) );
  AOI222_X1 U8778 ( .A1(n9666), .A2(n6988), .B1(n9124), .B2(n9695), .C1(n9125), 
        .C2(n9659), .ZN(n9611) );
  MUX2_X1 U8779 ( .A(n5776), .B(n9611), .S(n9393), .Z(n6994) );
  INV_X1 U8780 ( .A(n6989), .ZN(n7029) );
  INV_X1 U8781 ( .A(n7042), .ZN(n6990) );
  AOI211_X1 U8782 ( .C1(n9609), .C2(n7029), .A(n9562), .B(n6990), .ZN(n9608)
         );
  OAI22_X1 U8783 ( .A1(n9369), .A2(n6991), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9402), .ZN(n6992) );
  AOI21_X1 U8784 ( .B1(n9608), .B2(n9585), .A(n6992), .ZN(n6993) );
  OAI211_X1 U8785 ( .C1(n9612), .C2(n9414), .A(n6994), .B(n6993), .ZN(P1_U3290) );
  INV_X1 U8786 ( .A(n9215), .ZN(n8112) );
  INV_X1 U8787 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7001) );
  NOR2_X1 U8788 ( .A1(n7139), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6995) );
  AOI21_X1 U8789 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n7139), .A(n6995), .ZN(
        n6999) );
  OAI21_X1 U8790 ( .B1(n6997), .B2(n6813), .A(n6996), .ZN(n6998) );
  NAND2_X1 U8791 ( .A1(n6999), .A2(n6998), .ZN(n7142) );
  OAI211_X1 U8792 ( .C1(n6999), .C2(n6998), .A(n9211), .B(n7142), .ZN(n7000)
         );
  NAND2_X1 U8793 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7781) );
  OAI211_X1 U8794 ( .C1(n8112), .C2(n7001), .A(n7000), .B(n7781), .ZN(n7008)
         );
  AOI21_X1 U8795 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7003), .A(n7002), .ZN(
        n7006) );
  NAND2_X1 U8796 ( .A1(n7139), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7004) );
  OAI21_X1 U8797 ( .B1(n7139), .B2(P1_REG2_REG_14__SCAN_IN), .A(n7004), .ZN(
        n7005) );
  NOR2_X1 U8798 ( .A1(n7006), .A2(n7005), .ZN(n7138) );
  AOI211_X1 U8799 ( .C1(n7006), .C2(n7005), .A(n7138), .B(n7530), .ZN(n7007)
         );
  AOI211_X1 U8800 ( .C1(n9217), .C2(n7139), .A(n7008), .B(n7007), .ZN(n7009)
         );
  INV_X1 U8801 ( .A(n7009), .ZN(P1_U3257) );
  INV_X1 U8802 ( .A(n7010), .ZN(n7012) );
  INV_X1 U8803 ( .A(n7088), .ZN(n7011) );
  AOI21_X1 U8804 ( .B1(n7012), .B2(n8356), .A(n7011), .ZN(n9890) );
  NAND2_X1 U8805 ( .A1(n7013), .A2(n8691), .ZN(n9860) );
  XNOR2_X1 U8806 ( .A(n7014), .B(n8356), .ZN(n7015) );
  AOI222_X1 U8807 ( .A1(n9851), .A2(n7015), .B1(n8587), .B2(n9853), .C1(n9854), 
        .C2(n9855), .ZN(n9888) );
  MUX2_X1 U8808 ( .A(n7016), .B(n9888), .S(n9868), .Z(n7020) );
  AOI22_X1 U8809 ( .A1(n9842), .A2(n7018), .B1(n9843), .B2(n7017), .ZN(n7019)
         );
  OAI211_X1 U8810 ( .C1(n9890), .C2(n8833), .A(n7020), .B(n7019), .ZN(P2_U3229) );
  XNOR2_X1 U8811 ( .A(n7022), .B(n7934), .ZN(n9606) );
  XNOR2_X1 U8812 ( .A(n7023), .B(n7934), .ZN(n9603) );
  NOR2_X1 U8813 ( .A1(n9571), .A2(n9705), .ZN(n9404) );
  INV_X1 U8814 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7024) );
  OAI22_X1 U8815 ( .A1(n9393), .A2(n6457), .B1(n7024), .B2(n9402), .ZN(n7026)
         );
  NOR2_X1 U8816 ( .A1(n9369), .A2(n9602), .ZN(n7025) );
  AOI211_X1 U8817 ( .C1(n9404), .C2(n9599), .A(n7026), .B(n7025), .ZN(n7032)
         );
  AOI21_X1 U8818 ( .B1(n7027), .B2(n9083), .A(n9562), .ZN(n7028) );
  NAND2_X1 U8819 ( .A1(n7029), .A2(n7028), .ZN(n9601) );
  INV_X1 U8820 ( .A(n9601), .ZN(n7030) );
  INV_X1 U8821 ( .A(n9407), .ZN(n9309) );
  AOI22_X1 U8822 ( .A1(n7030), .A2(n9585), .B1(n9309), .B2(n9598), .ZN(n7031)
         );
  OAI211_X1 U8823 ( .C1(n9414), .C2(n9603), .A(n7032), .B(n7031), .ZN(n7033)
         );
  AOI21_X1 U8824 ( .B1(n9333), .B2(n9606), .A(n7033), .ZN(n7034) );
  INV_X1 U8825 ( .A(n7034), .ZN(P1_U3291) );
  NAND3_X1 U8826 ( .A1(n7035), .A2(n7809), .A3(n7040), .ZN(n7036) );
  NAND2_X1 U8827 ( .A1(n6963), .A2(n7036), .ZN(n7037) );
  NAND2_X1 U8828 ( .A1(n7037), .A2(n9666), .ZN(n7039) );
  NAND2_X1 U8829 ( .A1(n9598), .A2(n9659), .ZN(n7038) );
  NAND2_X1 U8830 ( .A1(n7039), .A2(n7038), .ZN(n9622) );
  INV_X1 U8831 ( .A(n9622), .ZN(n7052) );
  XNOR2_X1 U8832 ( .A(n7041), .B(n7040), .ZN(n9615) );
  AOI21_X1 U8833 ( .B1(n7042), .B2(n9616), .A(n9562), .ZN(n7044) );
  NAND2_X1 U8834 ( .A1(n7044), .A2(n7043), .ZN(n9619) );
  AOI22_X1 U8835 ( .A1(n9571), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7045), .B2(
        n9573), .ZN(n7046) );
  OAI21_X1 U8836 ( .B1(n9369), .B2(n7047), .A(n7046), .ZN(n7048) );
  AOI21_X1 U8837 ( .B1(n9309), .B2(n9617), .A(n7048), .ZN(n7049) );
  OAI21_X1 U8838 ( .B1(n9331), .B2(n9619), .A(n7049), .ZN(n7050) );
  AOI21_X1 U8839 ( .B1(n9586), .B2(n9615), .A(n7050), .ZN(n7051) );
  OAI21_X1 U8840 ( .B1(n7052), .B2(n9571), .A(n7051), .ZN(P1_U3289) );
  NAND2_X1 U8841 ( .A1(n7054), .A2(n7053), .ZN(n7056) );
  NAND2_X1 U8842 ( .A1(n7056), .A2(n7055), .ZN(n9580) );
  NAND2_X1 U8843 ( .A1(n9580), .A2(n9579), .ZN(n7058) );
  NAND2_X1 U8844 ( .A1(n7058), .A2(n7057), .ZN(n7059) );
  XNOR2_X1 U8845 ( .A(n7059), .B(n7817), .ZN(n9645) );
  INV_X1 U8846 ( .A(n9645), .ZN(n9648) );
  NAND2_X1 U8847 ( .A1(n7060), .A2(n7818), .ZN(n7061) );
  NOR2_X1 U8848 ( .A1(n7061), .A2(n7817), .ZN(n7118) );
  AOI21_X1 U8849 ( .B1(n7817), .B2(n7061), .A(n7118), .ZN(n7062) );
  NOR2_X1 U8850 ( .A1(n7062), .A2(n9712), .ZN(n9643) );
  AOI21_X1 U8851 ( .B1(n9582), .B2(n4352), .A(n9562), .ZN(n7063) );
  NAND2_X1 U8852 ( .A1(n7063), .A2(n9563), .ZN(n9641) );
  NAND2_X1 U8853 ( .A1(n9404), .A2(n9639), .ZN(n7066) );
  AOI22_X1 U8854 ( .A1(n9571), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7064), .B2(
        n9573), .ZN(n7065) );
  OAI211_X1 U8855 ( .C1(n7067), .C2(n9407), .A(n7066), .B(n7065), .ZN(n7068)
         );
  AOI21_X1 U8856 ( .B1(n9578), .B2(n4352), .A(n7068), .ZN(n7069) );
  OAI21_X1 U8857 ( .B1(n9641), .B2(n9331), .A(n7069), .ZN(n7070) );
  AOI21_X1 U8858 ( .B1(n9643), .B2(n9393), .A(n7070), .ZN(n7071) );
  OAI21_X1 U8859 ( .B1(n9648), .B2(n9414), .A(n7071), .ZN(P1_U3286) );
  XNOR2_X1 U8860 ( .A(n4456), .B(n7078), .ZN(n7181) );
  XNOR2_X1 U8861 ( .A(n7181), .B(n8587), .ZN(n7182) );
  INV_X1 U8862 ( .A(n7072), .ZN(n7073) );
  XOR2_X1 U8863 ( .A(n7183), .B(n7182), .Z(n7080) );
  INV_X1 U8864 ( .A(n8586), .ZN(n7255) );
  AOI21_X1 U8865 ( .B1(n8319), .B2(n9838), .A(n7074), .ZN(n7075) );
  OAI21_X1 U8866 ( .B1(n7255), .B2(n8321), .A(n7075), .ZN(n7077) );
  NOR2_X1 U8867 ( .A1(n7727), .A2(n7090), .ZN(n7076) );
  AOI211_X1 U8868 ( .C1(n7078), .C2(n8309), .A(n7077), .B(n7076), .ZN(n7079)
         );
  OAI21_X1 U8869 ( .B1(n7080), .B2(n8311), .A(n7079), .ZN(P2_U3167) );
  INV_X1 U8870 ( .A(n7081), .ZN(n7096) );
  AOI22_X1 U8871 ( .A1(n7519), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9529), .ZN(n7082) );
  OAI21_X1 U8872 ( .B1(n7096), .B2(n7754), .A(n7082), .ZN(P1_U3338) );
  INV_X1 U8873 ( .A(n9851), .ZN(n7546) );
  XNOR2_X1 U8874 ( .A(n7083), .B(n8358), .ZN(n7084) );
  OAI222_X1 U8875 ( .A1(n8703), .A2(n7255), .B1(n8701), .B2(n7085), .C1(n7546), 
        .C2(n7084), .ZN(n9894) );
  INV_X1 U8876 ( .A(n9894), .ZN(n7094) );
  INV_X1 U8877 ( .A(n8358), .ZN(n7087) );
  NAND3_X1 U8878 ( .A1(n7088), .A2(n7087), .A3(n8405), .ZN(n7089) );
  NAND2_X1 U8879 ( .A1(n7086), .A2(n7089), .ZN(n9896) );
  NOR2_X1 U8880 ( .A1(n9868), .A2(n6690), .ZN(n7092) );
  OAI22_X1 U8881 ( .A1(n8807), .A2(n9893), .B1(n7090), .B2(n9862), .ZN(n7091)
         );
  AOI211_X1 U8882 ( .C1(n9896), .C2(n9845), .A(n7092), .B(n7091), .ZN(n7093)
         );
  OAI21_X1 U8883 ( .B1(n7094), .B2(n9871), .A(n7093), .ZN(P2_U3228) );
  INV_X1 U8884 ( .A(n8648), .ZN(n9834) );
  OAI222_X1 U8885 ( .A1(n9834), .A2(P2_U3151), .B1(n8205), .B2(n7096), .C1(
        n7095), .C2(n8968), .ZN(P2_U3278) );
  OAI21_X1 U8886 ( .B1(n4446), .B2(n4897), .A(n7097), .ZN(n7098) );
  AOI22_X1 U8887 ( .A1(n7098), .A2(n9666), .B1(n9659), .B2(n9553), .ZN(n9673)
         );
  AOI22_X1 U8888 ( .A1(n9571), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7239), .B2(
        n9573), .ZN(n7099) );
  OAI21_X1 U8889 ( .B1(n9407), .B2(n7478), .A(n7099), .ZN(n7103) );
  OAI211_X1 U8890 ( .C1(n7101), .C2(n7100), .A(n9581), .B(n7171), .ZN(n9671)
         );
  NOR2_X1 U8891 ( .A1(n9671), .A2(n9331), .ZN(n7102) );
  AOI211_X1 U8892 ( .C1(n9578), .C2(n9670), .A(n7103), .B(n7102), .ZN(n7107)
         );
  XNOR2_X1 U8893 ( .A(n7105), .B(n7104), .ZN(n9675) );
  NAND2_X1 U8894 ( .A1(n9675), .A2(n9586), .ZN(n7106) );
  OAI211_X1 U8895 ( .C1(n9673), .C2(n9571), .A(n7107), .B(n7106), .ZN(P1_U3283) );
  INV_X1 U8896 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7109) );
  INV_X1 U8897 ( .A(n7108), .ZN(n7111) );
  OAI222_X1 U8898 ( .A1(n8968), .A2(n7109), .B1(n8205), .B2(n7111), .C1(
        P2_U3151), .C2(n8650), .ZN(P2_U3277) );
  INV_X1 U8899 ( .A(n8102), .ZN(n7536) );
  INV_X1 U8900 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7110) );
  OAI222_X1 U8901 ( .A1(P1_U3086), .A2(n7536), .B1(n7754), .B2(n7111), .C1(
        n7110), .C2(n9536), .ZN(P1_U3337) );
  NAND2_X1 U8902 ( .A1(n7112), .A2(n7113), .ZN(n7115) );
  NAND2_X1 U8903 ( .A1(n7115), .A2(n7114), .ZN(n7116) );
  XOR2_X1 U8904 ( .A(n7121), .B(n7116), .Z(n9664) );
  NOR2_X1 U8905 ( .A1(n7118), .A2(n7117), .ZN(n9549) );
  INV_X1 U8906 ( .A(n7820), .ZN(n7119) );
  OAI21_X1 U8907 ( .B1(n9549), .B2(n7119), .A(n7803), .ZN(n7120) );
  XOR2_X1 U8908 ( .A(n7121), .B(n7120), .Z(n9667) );
  NAND2_X1 U8909 ( .A1(n9667), .A2(n9333), .ZN(n7128) );
  NAND2_X1 U8910 ( .A1(n9404), .A2(n9658), .ZN(n7123) );
  AOI22_X1 U8911 ( .A1(n9571), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9048), .B2(
        n9573), .ZN(n7122) );
  NAND2_X1 U8912 ( .A1(n7123), .A2(n7122), .ZN(n7126) );
  XNOR2_X1 U8913 ( .A(n9561), .B(n9660), .ZN(n7124) );
  AOI22_X1 U8914 ( .A1(n7124), .A2(n9581), .B1(n9695), .B2(n9123), .ZN(n9662)
         );
  NOR2_X1 U8915 ( .A1(n9662), .A2(n9331), .ZN(n7125) );
  AOI211_X1 U8916 ( .C1(n9578), .C2(n9660), .A(n7126), .B(n7125), .ZN(n7127)
         );
  OAI211_X1 U8917 ( .C1(n9664), .C2(n9414), .A(n7128), .B(n7127), .ZN(P1_U3284) );
  NAND2_X1 U8918 ( .A1(n4445), .A2(n7129), .ZN(n9040) );
  OAI21_X1 U8919 ( .B1(n4445), .B2(n7129), .A(n9040), .ZN(n7130) );
  NOR2_X1 U8920 ( .A1(n7130), .A2(n7131), .ZN(n9043) );
  AOI21_X1 U8921 ( .B1(n7131), .B2(n7130), .A(n9043), .ZN(n7137) );
  AOI22_X1 U8922 ( .A1(n9058), .A2(n9557), .B1(n9116), .B2(n9569), .ZN(n7134)
         );
  INV_X1 U8923 ( .A(n7132), .ZN(n7133) );
  OAI211_X1 U8924 ( .C1(n7241), .C2(n9113), .A(n7134), .B(n7133), .ZN(n7135)
         );
  AOI21_X1 U8925 ( .B1(n6310), .B2(n9084), .A(n7135), .ZN(n7136) );
  OAI21_X1 U8926 ( .B1(n7137), .B2(n9075), .A(n7136), .ZN(P1_U3221) );
  INV_X1 U8927 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7141) );
  AOI21_X1 U8928 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7139), .A(n7138), .ZN(
        n7390) );
  XNOR2_X1 U8929 ( .A(n7390), .B(n7389), .ZN(n7140) );
  NOR2_X1 U8930 ( .A1(n7141), .A2(n7140), .ZN(n7391) );
  AOI211_X1 U8931 ( .C1(n7141), .C2(n7140), .A(n7391), .B(n7530), .ZN(n7148)
         );
  INV_X1 U8932 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9738) );
  OAI21_X1 U8933 ( .B1(n9738), .B2(n7143), .A(n7142), .ZN(n7381) );
  XNOR2_X1 U8934 ( .A(n7389), .B(n7381), .ZN(n7144) );
  NAND2_X1 U8935 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7144), .ZN(n7383) );
  OAI211_X1 U8936 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7144), .A(n9211), .B(
        n7383), .ZN(n7146) );
  AND2_X1 U8937 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9115) );
  AOI21_X1 U8938 ( .B1(n9215), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n9115), .ZN(
        n7145) );
  OAI211_X1 U8939 ( .C1(n9189), .C2(n7389), .A(n7146), .B(n7145), .ZN(n7147)
         );
  OR2_X1 U8940 ( .A1(n7148), .A2(n7147), .ZN(P1_U3258) );
  OR2_X1 U8941 ( .A1(n7191), .A2(n7149), .ZN(n7155) );
  AND2_X1 U8942 ( .A1(n7155), .A2(n7150), .ZN(n7253) );
  NAND2_X1 U8943 ( .A1(n7253), .A2(n7151), .ZN(n7153) );
  INV_X1 U8944 ( .A(n8360), .ZN(n7152) );
  NAND2_X1 U8945 ( .A1(n7153), .A2(n7152), .ZN(n7156) );
  NAND2_X1 U8946 ( .A1(n7155), .A2(n7154), .ZN(n7280) );
  NAND3_X1 U8947 ( .A1(n7156), .A2(n9851), .A3(n7280), .ZN(n7158) );
  AOI22_X1 U8948 ( .A1(n8583), .A2(n9853), .B1(n9855), .B2(n8585), .ZN(n7157)
         );
  OAI22_X1 U8949 ( .A1(n9868), .A2(n7215), .B1(n7310), .B2(n9862), .ZN(n7159)
         );
  AOI21_X1 U8950 ( .B1(n9842), .B2(n7315), .A(n7159), .ZN(n7163) );
  NAND2_X1 U8951 ( .A1(n7247), .A2(n7160), .ZN(n7161) );
  XNOR2_X1 U8952 ( .A(n7161), .B(n8360), .ZN(n9908) );
  NAND2_X1 U8953 ( .A1(n9908), .A2(n9845), .ZN(n7162) );
  OAI211_X1 U8954 ( .C1(n9912), .C2(n9871), .A(n7163), .B(n7162), .ZN(P2_U3225) );
  XNOR2_X1 U8955 ( .A(n7165), .B(n7164), .ZN(n9682) );
  INV_X1 U8956 ( .A(n9647), .ZN(n7170) );
  XNOR2_X1 U8957 ( .A(n7166), .B(n7944), .ZN(n7168) );
  AOI22_X1 U8958 ( .A1(n9659), .A2(n9123), .B1(n9122), .B2(n9695), .ZN(n7167)
         );
  OAI21_X1 U8959 ( .B1(n7168), .B2(n9712), .A(n7167), .ZN(n7169) );
  AOI21_X1 U8960 ( .B1(n9682), .B2(n7170), .A(n7169), .ZN(n9684) );
  AOI21_X1 U8961 ( .B1(n7171), .B2(n7292), .A(n9562), .ZN(n7172) );
  NAND2_X1 U8962 ( .A1(n7172), .A2(n7419), .ZN(n9677) );
  AOI22_X1 U8963 ( .A1(n9571), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7299), .B2(
        n9573), .ZN(n7174) );
  NAND2_X1 U8964 ( .A1(n7292), .A2(n9578), .ZN(n7173) );
  OAI211_X1 U8965 ( .C1(n9677), .C2(n9331), .A(n7174), .B(n7173), .ZN(n7175)
         );
  AOI21_X1 U8966 ( .B1(n9682), .B2(n9564), .A(n7175), .ZN(n7176) );
  OAI21_X1 U8967 ( .B1(n9684), .B2(n9571), .A(n7176), .ZN(P1_U3282) );
  INV_X1 U8968 ( .A(n7177), .ZN(n7196) );
  AOI21_X1 U8969 ( .B1(n8319), .B2(n8587), .A(n7178), .ZN(n7180) );
  NAND2_X1 U8970 ( .A1(n8303), .A2(n8585), .ZN(n7179) );
  OAI211_X1 U8971 ( .C1(n8326), .C2(n9900), .A(n7180), .B(n7179), .ZN(n7187)
         );
  XNOR2_X1 U8972 ( .A(n8170), .B(n9900), .ZN(n7201) );
  XNOR2_X1 U8973 ( .A(n7201), .B(n8586), .ZN(n7185) );
  NOR2_X1 U8974 ( .A1(n7184), .A2(n7185), .ZN(n7200) );
  AOI211_X1 U8975 ( .C1(n7185), .C2(n7184), .A(n8311), .B(n7200), .ZN(n7186)
         );
  AOI211_X1 U8976 ( .C1(n7196), .C2(n8323), .A(n7187), .B(n7186), .ZN(n7188)
         );
  INV_X1 U8977 ( .A(n7188), .ZN(P2_U3179) );
  NAND2_X1 U8978 ( .A1(n7086), .A2(n7189), .ZN(n7190) );
  XOR2_X1 U8979 ( .A(n8357), .B(n7190), .Z(n9898) );
  INV_X1 U8980 ( .A(n7191), .ZN(n7193) );
  INV_X1 U8981 ( .A(n8357), .ZN(n7192) );
  OR2_X1 U8982 ( .A1(n7191), .A2(n8357), .ZN(n7251) );
  OAI21_X1 U8983 ( .B1(n7193), .B2(n7192), .A(n7251), .ZN(n7194) );
  AOI222_X1 U8984 ( .A1(n9851), .A2(n7194), .B1(n8585), .B2(n9853), .C1(n8587), 
        .C2(n9855), .ZN(n9899) );
  MUX2_X1 U8985 ( .A(n7195), .B(n9899), .S(n9868), .Z(n7199) );
  AOI22_X1 U8986 ( .A1(n9842), .A2(n7197), .B1(n9843), .B2(n7196), .ZN(n7198)
         );
  OAI211_X1 U8987 ( .C1(n8833), .C2(n9898), .A(n7199), .B(n7198), .ZN(P2_U3227) );
  XNOR2_X1 U8988 ( .A(n4456), .B(n9903), .ZN(n7306) );
  XNOR2_X1 U8989 ( .A(n7306), .B(n8585), .ZN(n7202) );
  NAND2_X1 U8990 ( .A1(n7203), .A2(n7202), .ZN(n7309) );
  OAI21_X1 U8991 ( .B1(n7203), .B2(n7202), .A(n7309), .ZN(n7204) );
  NAND2_X1 U8992 ( .A1(n7204), .A2(n8316), .ZN(n7209) );
  INV_X1 U8993 ( .A(n8584), .ZN(n7368) );
  AOI21_X1 U8994 ( .B1(n8319), .B2(n8586), .A(n7205), .ZN(n7206) );
  OAI21_X1 U8995 ( .B1(n7368), .B2(n8321), .A(n7206), .ZN(n7207) );
  AOI21_X1 U8996 ( .B1(n7258), .B2(n8309), .A(n7207), .ZN(n7208) );
  OAI211_X1 U8997 ( .C1(n7256), .C2(n7727), .A(n7209), .B(n7208), .ZN(P2_U3153) );
  INV_X1 U8998 ( .A(n9769), .ZN(n7211) );
  INV_X1 U8999 ( .A(n9768), .ZN(n7210) );
  MUX2_X1 U9000 ( .A(n5300), .B(P2_REG1_REG_8__SCAN_IN), .S(n7214), .Z(n9766)
         );
  AOI21_X1 U9001 ( .B1(n7219), .B2(n7212), .A(n7324), .ZN(n7236) );
  INV_X1 U9002 ( .A(n7213), .ZN(n9762) );
  INV_X1 U9003 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7215) );
  MUX2_X1 U9004 ( .A(n7215), .B(P2_REG2_REG_8__SCAN_IN), .S(n7214), .Z(n9761)
         );
  AOI21_X1 U9005 ( .B1(n7220), .B2(n7216), .A(n7319), .ZN(n7217) );
  NOR2_X1 U9006 ( .A1(n7217), .A2(n9829), .ZN(n7234) );
  NOR2_X1 U9007 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5114), .ZN(n7374) );
  INV_X1 U9008 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9972) );
  OAI22_X1 U9009 ( .A1(n9835), .A2(n7218), .B1(n9783), .B2(n9972), .ZN(n7233)
         );
  MUX2_X1 U9010 ( .A(n7220), .B(n7219), .S(n8631), .Z(n7222) );
  AND2_X1 U9011 ( .A1(n7222), .A2(n7323), .ZN(n7335) );
  INV_X1 U9012 ( .A(n7335), .ZN(n7221) );
  OAI21_X1 U9013 ( .B1(n7323), .B2(n7222), .A(n7221), .ZN(n7230) );
  MUX2_X1 U9014 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8631), .Z(n7227) );
  NOR2_X1 U9015 ( .A1(n7227), .A2(n9772), .ZN(n7228) );
  INV_X1 U9016 ( .A(n7223), .ZN(n7226) );
  OAI21_X1 U9017 ( .B1(n7226), .B2(n7225), .A(n7224), .ZN(n9778) );
  AOI21_X1 U9018 ( .B1(n7227), .B2(n9772), .A(n7228), .ZN(n9777) );
  AND2_X1 U9019 ( .A1(n9778), .A2(n9777), .ZN(n9780) );
  NOR2_X1 U9020 ( .A1(n7228), .A2(n9780), .ZN(n7229) );
  NOR2_X1 U9021 ( .A1(n7229), .A2(n7230), .ZN(n7334) );
  AOI21_X1 U9022 ( .B1(n7230), .B2(n7229), .A(n7334), .ZN(n7231) );
  NOR2_X1 U9023 ( .A1(n7231), .A2(n7512), .ZN(n7232) );
  NOR4_X1 U9024 ( .A1(n7234), .A2(n7374), .A3(n7233), .A4(n7232), .ZN(n7235)
         );
  OAI21_X1 U9025 ( .B1(n7236), .B2(n9825), .A(n7235), .ZN(P2_U3191) );
  NOR2_X1 U9026 ( .A1(n7237), .A2(n7238), .ZN(n7295) );
  AOI21_X1 U9027 ( .B1(n7238), .B2(n7237), .A(n7295), .ZN(n7246) );
  INV_X1 U9028 ( .A(n9081), .ZN(n9070) );
  INV_X1 U9029 ( .A(n7239), .ZN(n7240) );
  OAI22_X1 U9030 ( .A1(n9070), .A2(n7241), .B1(n7240), .B2(n9112), .ZN(n7242)
         );
  AOI211_X1 U9031 ( .C1(n9102), .C2(n9669), .A(n7243), .B(n7242), .ZN(n7245)
         );
  NAND2_X1 U9032 ( .A1(n9670), .A2(n9084), .ZN(n7244) );
  OAI211_X1 U9033 ( .C1(n7246), .C2(n9075), .A(n7245), .B(n7244), .ZN(P1_U3217) );
  OAI21_X1 U9034 ( .B1(n7248), .B2(n7250), .A(n7247), .ZN(n9904) );
  NAND3_X1 U9035 ( .A1(n7251), .A2(n7250), .A3(n7249), .ZN(n7252) );
  AND2_X1 U9036 ( .A1(n7253), .A2(n7252), .ZN(n7254) );
  OAI222_X1 U9037 ( .A1(n8703), .A2(n7368), .B1(n8701), .B2(n7255), .C1(n7546), 
        .C2(n7254), .ZN(n9906) );
  NAND2_X1 U9038 ( .A1(n9906), .A2(n9868), .ZN(n7260) );
  OAI22_X1 U9039 ( .A1(n9868), .A2(n6828), .B1(n7256), .B2(n9862), .ZN(n7257)
         );
  AOI21_X1 U9040 ( .B1(n9842), .B2(n7258), .A(n7257), .ZN(n7259) );
  OAI211_X1 U9041 ( .C1(n8833), .C2(n9904), .A(n7260), .B(n7259), .ZN(P2_U3226) );
  INV_X1 U9042 ( .A(n7261), .ZN(n7264) );
  OAI222_X1 U9043 ( .A1(n9536), .A2(n7262), .B1(n7754), .B2(n7264), .C1(n8063), 
        .C2(P1_U3086), .ZN(P1_U3336) );
  OAI222_X1 U9044 ( .A1(n8673), .A2(P2_U3151), .B1(n8205), .B2(n7264), .C1(
        n7263), .C2(n8968), .ZN(P2_U3276) );
  AND2_X1 U9045 ( .A1(n7266), .A2(n7265), .ZN(n7278) );
  NAND3_X1 U9046 ( .A1(n7278), .A2(n4719), .A3(n7267), .ZN(n7268) );
  NAND2_X1 U9047 ( .A1(n7269), .A2(n7268), .ZN(n7272) );
  NAND2_X1 U9048 ( .A1(n8581), .A2(n9853), .ZN(n7270) );
  OAI21_X1 U9049 ( .B1(n7614), .B2(n8701), .A(n7270), .ZN(n7271) );
  AOI21_X1 U9050 ( .B1(n7272), .B2(n9851), .A(n7271), .ZN(n9924) );
  OAI22_X1 U9051 ( .A1(n9868), .A2(n7331), .B1(n7619), .B2(n9862), .ZN(n7273)
         );
  AOI21_X1 U9052 ( .B1(n9842), .B2(n9921), .A(n7273), .ZN(n7277) );
  NAND2_X1 U9053 ( .A1(n7284), .A2(n8419), .ZN(n7275) );
  XNOR2_X1 U9054 ( .A(n7275), .B(n7274), .ZN(n9920) );
  NAND2_X1 U9055 ( .A1(n9920), .A2(n9845), .ZN(n7276) );
  OAI211_X1 U9056 ( .C1(n9924), .C2(n9871), .A(n7277), .B(n7276), .ZN(P2_U3223) );
  INV_X1 U9057 ( .A(n7278), .ZN(n7282) );
  AOI21_X1 U9058 ( .B1(n7280), .B2(n7279), .A(n8361), .ZN(n7281) );
  NOR2_X1 U9059 ( .A1(n7282), .A2(n7281), .ZN(n7283) );
  OAI222_X1 U9060 ( .A1(n8701), .A2(n7368), .B1(n8703), .B2(n7674), .C1(n7546), 
        .C2(n7283), .ZN(n9915) );
  INV_X1 U9061 ( .A(n9915), .ZN(n7291) );
  INV_X1 U9062 ( .A(n7284), .ZN(n7285) );
  AOI21_X1 U9063 ( .B1(n8361), .B2(n7286), .A(n7285), .ZN(n9917) );
  INV_X1 U9064 ( .A(n7378), .ZN(n9914) );
  INV_X1 U9065 ( .A(n7287), .ZN(n7373) );
  AOI22_X1 U9066 ( .A1(n9871), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n9843), .B2(
        n7373), .ZN(n7288) );
  OAI21_X1 U9067 ( .B1(n9914), .B2(n8807), .A(n7288), .ZN(n7289) );
  AOI21_X1 U9068 ( .B1(n9917), .B2(n9845), .A(n7289), .ZN(n7290) );
  OAI21_X1 U9069 ( .B1(n7291), .B2(n9871), .A(n7290), .ZN(P2_U3224) );
  INV_X1 U9070 ( .A(n7292), .ZN(n9679) );
  NOR3_X1 U9071 ( .A1(n7295), .A2(n7294), .A3(n7293), .ZN(n7298) );
  NAND2_X1 U9072 ( .A1(n7297), .A2(n7296), .ZN(n7479) );
  OAI21_X1 U9073 ( .B1(n7298), .B2(n7479), .A(n9109), .ZN(n7305) );
  INV_X1 U9074 ( .A(n7299), .ZN(n7300) );
  OAI22_X1 U9075 ( .A1(n9070), .A2(n7301), .B1(n7300), .B2(n9112), .ZN(n7302)
         );
  AOI211_X1 U9076 ( .C1(n9102), .C2(n9122), .A(n7303), .B(n7302), .ZN(n7304)
         );
  OAI211_X1 U9077 ( .C1(n9679), .C2(n9119), .A(n7305), .B(n7304), .ZN(P1_U3236) );
  XNOR2_X1 U9078 ( .A(n8170), .B(n7315), .ZN(n7367) );
  XNOR2_X1 U9079 ( .A(n7367), .B(n8584), .ZN(n7369) );
  XOR2_X1 U9080 ( .A(n7370), .B(n7369), .Z(n7317) );
  INV_X1 U9081 ( .A(n7310), .ZN(n7311) );
  NAND2_X1 U9082 ( .A1(n8323), .A2(n7311), .ZN(n7313) );
  INV_X1 U9083 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U9084 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10049), .ZN(n9774) );
  AOI21_X1 U9085 ( .B1(n8319), .B2(n8585), .A(n9774), .ZN(n7312) );
  OAI211_X1 U9086 ( .C1(n7614), .C2(n8321), .A(n7313), .B(n7312), .ZN(n7314)
         );
  AOI21_X1 U9087 ( .B1(n7315), .B2(n8309), .A(n7314), .ZN(n7316) );
  OAI21_X1 U9088 ( .B1(n7317), .B2(n8311), .A(n7316), .ZN(P2_U3161) );
  MUX2_X1 U9089 ( .A(n7331), .B(P2_REG2_REG_10__SCAN_IN), .S(n7463), .Z(n7320)
         );
  AOI21_X1 U9090 ( .B1(n7321), .B2(n7320), .A(n4447), .ZN(n7346) );
  NOR2_X1 U9091 ( .A1(n7323), .A2(n7322), .ZN(n7325) );
  INV_X1 U9092 ( .A(n7327), .ZN(n7329) );
  INV_X1 U9093 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7330) );
  MUX2_X1 U9094 ( .A(n7330), .B(P2_REG1_REG_10__SCAN_IN), .S(n7463), .Z(n7326)
         );
  INV_X1 U9095 ( .A(n7326), .ZN(n7328) );
  OAI21_X1 U9096 ( .B1(n7329), .B2(n7328), .A(n7444), .ZN(n7344) );
  MUX2_X1 U9097 ( .A(n7331), .B(n7330), .S(n8631), .Z(n7333) );
  AND2_X1 U9098 ( .A1(n7333), .A2(n7338), .ZN(n7453) );
  INV_X1 U9099 ( .A(n7453), .ZN(n7332) );
  OAI21_X1 U9100 ( .B1(n7338), .B2(n7333), .A(n7332), .ZN(n7337) );
  NOR2_X1 U9101 ( .A1(n7335), .A2(n7334), .ZN(n7336) );
  NOR2_X1 U9102 ( .A1(n7336), .A2(n7337), .ZN(n7452) );
  AOI21_X1 U9103 ( .B1(n7337), .B2(n7336), .A(n7452), .ZN(n7341) );
  INV_X1 U9104 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9976) );
  OR2_X1 U9105 ( .A1(n9783), .A2(n9976), .ZN(n7340) );
  INV_X1 U9106 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U9107 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10062), .ZN(n7618) );
  AOI21_X1 U9108 ( .B1(n8600), .B2(n7338), .A(n7618), .ZN(n7339) );
  OAI211_X1 U9109 ( .C1(n7341), .C2(n7512), .A(n7340), .B(n7339), .ZN(n7342)
         );
  AOI21_X1 U9110 ( .B1(n7344), .B2(n7343), .A(n7342), .ZN(n7345) );
  OAI21_X1 U9111 ( .B1(n7346), .B2(n9829), .A(n7345), .ZN(P2_U3192) );
  INV_X1 U9112 ( .A(n7347), .ZN(n7360) );
  AOI21_X1 U9113 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(n9529), .A(n7348), .ZN(
        n7349) );
  OAI21_X1 U9114 ( .B1(n7360), .B2(n7754), .A(n7349), .ZN(P1_U3335) );
  XNOR2_X1 U9115 ( .A(n7350), .B(n7947), .ZN(n7351) );
  AOI22_X1 U9116 ( .A1(n7351), .A2(n9666), .B1(n9659), .B2(n9122), .ZN(n9699)
         );
  XNOR2_X1 U9117 ( .A(n7352), .B(n7947), .ZN(n9701) );
  INV_X1 U9118 ( .A(n7438), .ZN(n7353) );
  OAI211_X1 U9119 ( .C1(n7413), .C2(n4444), .A(n7353), .B(n9581), .ZN(n9697)
         );
  AOI22_X1 U9120 ( .A1(n9571), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7406), .B2(
        n9573), .ZN(n7354) );
  OAI21_X1 U9121 ( .B1(n9407), .B2(n7408), .A(n7354), .ZN(n7355) );
  AOI21_X1 U9122 ( .B1(n9696), .B2(n9578), .A(n7355), .ZN(n7356) );
  OAI21_X1 U9123 ( .B1(n9697), .B2(n9331), .A(n7356), .ZN(n7357) );
  AOI21_X1 U9124 ( .B1(n9701), .B2(n9586), .A(n7357), .ZN(n7358) );
  OAI21_X1 U9125 ( .B1(n9571), .B2(n9699), .A(n7358), .ZN(P1_U3280) );
  OAI222_X1 U9126 ( .A1(P2_U3151), .A2(n8566), .B1(n8205), .B2(n7360), .C1(
        n7359), .C2(n8968), .ZN(P2_U3275) );
  INV_X1 U9127 ( .A(n8439), .ZN(n8436) );
  NOR2_X1 U9128 ( .A1(n8436), .A2(n8440), .ZN(n8363) );
  XOR2_X1 U9129 ( .A(n7361), .B(n8363), .Z(n9926) );
  XNOR2_X1 U9130 ( .A(n7362), .B(n8363), .ZN(n7363) );
  OAI222_X1 U9131 ( .A1(n8703), .A2(n7673), .B1(n8701), .B2(n7674), .C1(n7546), 
        .C2(n7363), .ZN(n9927) );
  NAND2_X1 U9132 ( .A1(n9927), .A2(n9868), .ZN(n7366) );
  OAI22_X1 U9133 ( .A1(n9868), .A2(n7451), .B1(n7653), .B2(n9862), .ZN(n7364)
         );
  AOI21_X1 U9134 ( .B1(n9929), .B2(n9842), .A(n7364), .ZN(n7365) );
  OAI211_X1 U9135 ( .C1(n8833), .C2(n9926), .A(n7366), .B(n7365), .ZN(P2_U3222) );
  XNOR2_X1 U9136 ( .A(n7378), .B(n8170), .ZN(n7615) );
  XNOR2_X1 U9137 ( .A(n7615), .B(n8583), .ZN(n7371) );
  NAND2_X1 U9138 ( .A1(n7372), .A2(n7371), .ZN(n7617) );
  OAI211_X1 U9139 ( .C1(n7372), .C2(n7371), .A(n7617), .B(n8316), .ZN(n7380)
         );
  NAND2_X1 U9140 ( .A1(n8323), .A2(n7373), .ZN(n7376) );
  AOI21_X1 U9141 ( .B1(n8319), .B2(n8584), .A(n7374), .ZN(n7375) );
  OAI211_X1 U9142 ( .C1(n7674), .C2(n8321), .A(n7376), .B(n7375), .ZN(n7377)
         );
  AOI21_X1 U9143 ( .B1(n7378), .B2(n8309), .A(n7377), .ZN(n7379) );
  NAND2_X1 U9144 ( .A1(n7380), .A2(n7379), .ZN(P2_U3171) );
  NAND2_X1 U9145 ( .A1(n7382), .A2(n7381), .ZN(n7384) );
  NAND2_X1 U9146 ( .A1(n7384), .A2(n7383), .ZN(n7388) );
  INV_X1 U9147 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7385) );
  NAND2_X1 U9148 ( .A1(n7386), .A2(n7385), .ZN(n7489) );
  OAI21_X1 U9149 ( .B1(n7386), .B2(n7385), .A(n7489), .ZN(n7387) );
  NOR2_X1 U9150 ( .A1(n7388), .A2(n7387), .ZN(n7491) );
  AOI21_X1 U9151 ( .B1(n7388), .B2(n7387), .A(n7491), .ZN(n7401) );
  AND2_X1 U9152 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9019) );
  NOR2_X1 U9153 ( .A1(n7390), .A2(n7389), .ZN(n7392) );
  NOR2_X1 U9154 ( .A1(n7392), .A2(n7391), .ZN(n7396) );
  NAND2_X1 U9155 ( .A1(n7398), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7494) );
  OR2_X1 U9156 ( .A1(n7398), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7393) );
  NAND2_X1 U9157 ( .A1(n7494), .A2(n7393), .ZN(n7395) );
  OR2_X1 U9158 ( .A1(n7396), .A2(n7395), .ZN(n7495) );
  INV_X1 U9159 ( .A(n7495), .ZN(n7394) );
  AOI211_X1 U9160 ( .C1(n7396), .C2(n7395), .A(n7394), .B(n7530), .ZN(n7397)
         );
  AOI211_X1 U9161 ( .C1(n9215), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9019), .B(
        n7397), .ZN(n7400) );
  NAND2_X1 U9162 ( .A1(n9217), .A2(n7398), .ZN(n7399) );
  OAI211_X1 U9163 ( .C1(n7401), .C2(n9165), .A(n7400), .B(n7399), .ZN(P1_U3259) );
  OAI21_X1 U9164 ( .B1(n7404), .B2(n7402), .A(n7403), .ZN(n7405) );
  NAND2_X1 U9165 ( .A1(n7405), .A2(n9109), .ZN(n7412) );
  INV_X1 U9166 ( .A(n7406), .ZN(n7407) );
  OAI22_X1 U9167 ( .A1(n9113), .A2(n7408), .B1(n7407), .B2(n9112), .ZN(n7409)
         );
  AOI211_X1 U9168 ( .C1(n9116), .C2(n9122), .A(n7410), .B(n7409), .ZN(n7411)
         );
  OAI211_X1 U9169 ( .C1(n7413), .C2(n9119), .A(n7412), .B(n7411), .ZN(P1_U3234) );
  OAI222_X1 U9170 ( .A1(P2_U3151), .A2(n8375), .B1(n8205), .B2(n7416), .C1(
        n7414), .C2(n8968), .ZN(P2_U3274) );
  OAI222_X1 U9171 ( .A1(P1_U3086), .A2(n7932), .B1(n7754), .B2(n7416), .C1(
        n7415), .C2(n9536), .ZN(P1_U3334) );
  XNOR2_X1 U9172 ( .A(n7418), .B(n7417), .ZN(n9692) );
  NAND2_X1 U9173 ( .A1(n7419), .A2(n9687), .ZN(n7420) );
  NAND2_X1 U9174 ( .A1(n7420), .A2(n9581), .ZN(n7421) );
  OR2_X1 U9175 ( .A1(n4444), .A2(n7421), .ZN(n9688) );
  AOI22_X1 U9176 ( .A1(n9571), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7475), .B2(
        n9573), .ZN(n7422) );
  OAI21_X1 U9177 ( .B1(n9407), .B2(n9706), .A(n7422), .ZN(n7423) );
  AOI21_X1 U9178 ( .B1(n9687), .B2(n9578), .A(n7423), .ZN(n7424) );
  OAI21_X1 U9179 ( .B1(n9688), .B2(n9331), .A(n7424), .ZN(n7428) );
  OAI21_X1 U9180 ( .B1(n7946), .B2(n4441), .A(n7425), .ZN(n7426) );
  AOI22_X1 U9181 ( .A1(n7426), .A2(n9666), .B1(n9659), .B2(n9669), .ZN(n9690)
         );
  NOR2_X1 U9182 ( .A1(n9690), .A2(n9571), .ZN(n7427) );
  AOI211_X1 U9183 ( .C1(n9586), .C2(n9692), .A(n7428), .B(n7427), .ZN(n7429)
         );
  INV_X1 U9184 ( .A(n7429), .ZN(P1_U3281) );
  INV_X1 U9185 ( .A(n7430), .ZN(n7431) );
  AOI21_X1 U9186 ( .B1(n7433), .B2(n7432), .A(n7431), .ZN(n9713) );
  INV_X1 U9187 ( .A(n9333), .ZN(n9268) );
  XNOR2_X1 U9188 ( .A(n7434), .B(n7433), .ZN(n9715) );
  NAND2_X1 U9189 ( .A1(n9715), .A2(n9586), .ZN(n7442) );
  NAND2_X1 U9190 ( .A1(n9404), .A2(n9686), .ZN(n7436) );
  AOI22_X1 U9191 ( .A1(n9571), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7780), .B2(
        n9573), .ZN(n7435) );
  OAI211_X1 U9192 ( .C1(n9704), .C2(n9407), .A(n7436), .B(n7435), .ZN(n7440)
         );
  OAI211_X1 U9193 ( .C1(n7438), .C2(n7437), .A(n9581), .B(n7602), .ZN(n9710)
         );
  NOR2_X1 U9194 ( .A1(n9710), .A2(n9331), .ZN(n7439) );
  AOI211_X1 U9195 ( .C1(n9578), .C2(n9709), .A(n7440), .B(n7439), .ZN(n7441)
         );
  OAI211_X1 U9196 ( .C1(n9713), .C2(n9268), .A(n7442), .B(n7441), .ZN(P1_U3279) );
  NAND2_X1 U9197 ( .A1(n7463), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7443) );
  NOR2_X1 U9198 ( .A1(n7466), .A2(n7445), .ZN(n7446) );
  XNOR2_X1 U9199 ( .A(n7466), .B(n7445), .ZN(n7504) );
  NOR2_X1 U9200 ( .A1(n7446), .A2(n7503), .ZN(n7449) );
  OR2_X1 U9201 ( .A1(n7580), .A2(n7566), .ZN(n7574) );
  NAND2_X1 U9202 ( .A1(n7580), .A2(n7566), .ZN(n7447) );
  NAND2_X1 U9203 ( .A1(n7574), .A2(n7447), .ZN(n7448) );
  AOI21_X1 U9204 ( .B1(n7449), .B2(n7448), .A(n4927), .ZN(n7474) );
  MUX2_X1 U9205 ( .A(n7451), .B(n7450), .S(n8631), .Z(n7455) );
  AND2_X1 U9206 ( .A1(n7455), .A2(n7466), .ZN(n7456) );
  NOR2_X1 U9207 ( .A1(n7453), .A2(n7452), .ZN(n7510) );
  INV_X1 U9208 ( .A(n7456), .ZN(n7454) );
  OAI21_X1 U9209 ( .B1(n7466), .B2(n7455), .A(n7454), .ZN(n7511) );
  NOR2_X1 U9210 ( .A1(n7510), .A2(n7511), .ZN(n7509) );
  NOR2_X1 U9211 ( .A1(n7456), .A2(n7509), .ZN(n7571) );
  MUX2_X1 U9212 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8631), .Z(n7458) );
  INV_X1 U9213 ( .A(n7580), .ZN(n7457) );
  AND2_X1 U9214 ( .A1(n7458), .A2(n7457), .ZN(n7569) );
  INV_X1 U9215 ( .A(n7569), .ZN(n7460) );
  MUX2_X1 U9216 ( .A(n7579), .B(n7566), .S(n8631), .Z(n7459) );
  NAND2_X1 U9217 ( .A1(n7459), .A2(n7580), .ZN(n7570) );
  NAND2_X1 U9218 ( .A1(n7460), .A2(n7570), .ZN(n7461) );
  XNOR2_X1 U9219 ( .A(n7571), .B(n7461), .ZN(n7462) );
  NAND2_X1 U9220 ( .A1(n7462), .A2(n9832), .ZN(n7473) );
  NAND2_X1 U9221 ( .A1(n7463), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7464) );
  MUX2_X1 U9222 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7579), .S(n7580), .Z(n7467)
         );
  OAI21_X1 U9223 ( .B1(n4835), .B2(n4834), .A(n7582), .ZN(n7471) );
  INV_X1 U9224 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9984) );
  NOR2_X1 U9225 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10040), .ZN(n7670) );
  AOI21_X1 U9226 ( .B1(n8600), .B2(n7580), .A(n7670), .ZN(n7468) );
  OAI21_X1 U9227 ( .B1(n9984), .B2(n9783), .A(n7468), .ZN(n7469) );
  AOI21_X1 U9228 ( .B1(n7471), .B2(n7470), .A(n7469), .ZN(n7472) );
  OAI211_X1 U9229 ( .C1(n7474), .C2(n9825), .A(n7473), .B(n7472), .ZN(P2_U3194) );
  AOI22_X1 U9230 ( .A1(n9058), .A2(n7475), .B1(n9102), .B2(n9686), .ZN(n7477)
         );
  OAI211_X1 U9231 ( .C1(n7478), .C2(n9070), .A(n7477), .B(n7476), .ZN(n7487)
         );
  INV_X1 U9232 ( .A(n7479), .ZN(n7483) );
  INV_X1 U9233 ( .A(n7480), .ZN(n7481) );
  NAND3_X1 U9234 ( .A1(n7483), .A2(n7482), .A3(n7481), .ZN(n7484) );
  AOI21_X1 U9235 ( .B1(n7485), .B2(n7484), .A(n9075), .ZN(n7486) );
  AOI211_X1 U9236 ( .C1(n9687), .C2(n9084), .A(n7487), .B(n7486), .ZN(n7488)
         );
  INV_X1 U9237 ( .A(n7488), .ZN(P1_U3224) );
  INV_X1 U9238 ( .A(n7489), .ZN(n7490) );
  NOR2_X1 U9239 ( .A1(n7491), .A2(n7490), .ZN(n7493) );
  XNOR2_X1 U9240 ( .A(n7519), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7492) );
  NOR2_X1 U9241 ( .A1(n7493), .A2(n7492), .ZN(n7522) );
  AOI21_X1 U9242 ( .B1(n7493), .B2(n7492), .A(n7522), .ZN(n7502) );
  AND2_X1 U9243 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9028) );
  AND2_X1 U9244 ( .A1(n7495), .A2(n7494), .ZN(n7498) );
  OR2_X1 U9245 ( .A1(n7519), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7525) );
  NAND2_X1 U9246 ( .A1(n7519), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7496) );
  AND2_X1 U9247 ( .A1(n7525), .A2(n7496), .ZN(n7497) );
  NAND2_X1 U9248 ( .A1(n7498), .A2(n7497), .ZN(n7526) );
  AOI221_X1 U9249 ( .B1(n7498), .B2(n7526), .C1(n7497), .C2(n7526), .A(n7530), 
        .ZN(n7499) );
  AOI211_X1 U9250 ( .C1(n9215), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9028), .B(
        n7499), .ZN(n7501) );
  NAND2_X1 U9251 ( .A1(n9217), .A2(n7519), .ZN(n7500) );
  OAI211_X1 U9252 ( .C1(n7502), .C2(n9165), .A(n7501), .B(n7500), .ZN(P1_U3260) );
  AOI21_X1 U9253 ( .B1(n7450), .B2(n7504), .A(n7503), .ZN(n7518) );
  AOI21_X1 U9254 ( .B1(n7451), .B2(n7506), .A(n7505), .ZN(n7507) );
  NOR2_X1 U9255 ( .A1(n7507), .A2(n9829), .ZN(n7516) );
  INV_X1 U9256 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10157) );
  NOR2_X1 U9257 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10157), .ZN(n7651) );
  INV_X1 U9258 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9980) );
  OAI22_X1 U9259 ( .A1(n9835), .A2(n7508), .B1(n9783), .B2(n9980), .ZN(n7515)
         );
  AOI21_X1 U9260 ( .B1(n7511), .B2(n7510), .A(n7509), .ZN(n7513) );
  NOR2_X1 U9261 ( .A1(n7513), .A2(n7512), .ZN(n7514) );
  NOR4_X1 U9262 ( .A1(n7516), .A2(n7651), .A3(n7515), .A4(n7514), .ZN(n7517)
         );
  OAI21_X1 U9263 ( .B1(n7518), .B2(n9825), .A(n7517), .ZN(P2_U3193) );
  NOR2_X1 U9264 ( .A1(n7519), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n7521) );
  XNOR2_X1 U9265 ( .A(n8102), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n7520) );
  NOR3_X1 U9266 ( .A1(n7522), .A2(n7521), .A3(n7520), .ZN(n8101) );
  INV_X1 U9267 ( .A(n8101), .ZN(n7524) );
  OAI21_X1 U9268 ( .B1(n7522), .B2(n7521), .A(n7520), .ZN(n7523) );
  NAND3_X1 U9269 ( .A1(n7524), .A2(n9211), .A3(n7523), .ZN(n7535) );
  AND2_X1 U9270 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9093) );
  NAND2_X1 U9271 ( .A1(n7526), .A2(n7525), .ZN(n7532) );
  NAND2_X1 U9272 ( .A1(n7536), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7529) );
  INV_X1 U9273 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n7527) );
  NAND2_X1 U9274 ( .A1(n8102), .A2(n7527), .ZN(n7528) );
  AND2_X1 U9275 ( .A1(n7529), .A2(n7528), .ZN(n7531) );
  NOR2_X1 U9276 ( .A1(n7532), .A2(n7531), .ZN(n8098) );
  AOI211_X1 U9277 ( .C1(n7532), .C2(n7531), .A(n8098), .B(n7530), .ZN(n7533)
         );
  AOI211_X1 U9278 ( .C1(n9215), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9093), .B(
        n7533), .ZN(n7534) );
  OAI211_X1 U9279 ( .C1(n9189), .C2(n7536), .A(n7535), .B(n7534), .ZN(P1_U3261) );
  XNOR2_X1 U9280 ( .A(n7537), .B(n8367), .ZN(n7538) );
  OAI222_X1 U9281 ( .A1(n8703), .A2(n7756), .B1(n8701), .B2(n7673), .C1(n7546), 
        .C2(n7538), .ZN(n7553) );
  INV_X1 U9282 ( .A(n8451), .ZN(n7702) );
  OAI22_X1 U9283 ( .A1(n7702), .A2(n8742), .B1(n7695), .B2(n9862), .ZN(n7539)
         );
  OAI21_X1 U9284 ( .B1(n7553), .B2(n7539), .A(n9868), .ZN(n7542) );
  XNOR2_X1 U9285 ( .A(n7540), .B(n8367), .ZN(n7558) );
  AOI22_X1 U9286 ( .A1(n7558), .A2(n9845), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n9871), .ZN(n7541) );
  NAND2_X1 U9287 ( .A1(n7542), .A2(n7541), .ZN(P2_U3220) );
  XOR2_X1 U9288 ( .A(n7543), .B(n8445), .Z(n7564) );
  INV_X1 U9289 ( .A(n7564), .ZN(n7552) );
  INV_X1 U9290 ( .A(n7672), .ZN(n7544) );
  AOI22_X1 U9291 ( .A1(n7688), .A2(n9842), .B1(n9843), .B2(n7544), .ZN(n7551)
         );
  AOI21_X1 U9292 ( .B1(n7545), .B2(n8445), .A(n7546), .ZN(n7549) );
  OAI22_X1 U9293 ( .A1(n7675), .A2(n8701), .B1(n7722), .B2(n8703), .ZN(n7547)
         );
  AOI21_X1 U9294 ( .B1(n7549), .B2(n7548), .A(n7547), .ZN(n7565) );
  MUX2_X1 U9295 ( .A(n7579), .B(n7565), .S(n9868), .Z(n7550) );
  OAI211_X1 U9296 ( .C1(n7552), .C2(n8833), .A(n7551), .B(n7550), .ZN(P2_U3221) );
  INV_X1 U9297 ( .A(n7553), .ZN(n7556) );
  MUX2_X1 U9298 ( .A(n7576), .B(n7556), .S(n9947), .Z(n7555) );
  AOI22_X1 U9299 ( .A1(n7558), .A2(n8876), .B1(n8875), .B2(n8451), .ZN(n7554)
         );
  NAND2_X1 U9300 ( .A1(n7555), .A2(n7554), .ZN(P2_U3472) );
  INV_X1 U9301 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7557) );
  MUX2_X1 U9302 ( .A(n7557), .B(n7556), .S(n9931), .Z(n7560) );
  INV_X1 U9303 ( .A(n9919), .ZN(n9925) );
  AOI22_X1 U9304 ( .A1(n7558), .A2(n8953), .B1(n8952), .B2(n8451), .ZN(n7559)
         );
  NAND2_X1 U9305 ( .A1(n7560), .A2(n7559), .ZN(P2_U3429) );
  AOI22_X1 U9306 ( .A1(n7564), .A2(n8953), .B1(n8952), .B2(n7688), .ZN(n7563)
         );
  INV_X1 U9307 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7561) );
  MUX2_X1 U9308 ( .A(n7561), .B(n7565), .S(n9931), .Z(n7562) );
  NAND2_X1 U9309 ( .A1(n7563), .A2(n7562), .ZN(P2_U3426) );
  AOI22_X1 U9310 ( .A1(n7564), .A2(n8876), .B1(n8875), .B2(n7688), .ZN(n7568)
         );
  MUX2_X1 U9311 ( .A(n7566), .B(n7565), .S(n9947), .Z(n7567) );
  NAND2_X1 U9312 ( .A1(n7568), .A2(n7567), .ZN(P2_U3471) );
  AOI21_X1 U9313 ( .B1(n7571), .B2(n7570), .A(n7569), .ZN(n7573) );
  MUX2_X1 U9314 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8631), .Z(n8593) );
  XNOR2_X1 U9315 ( .A(n8593), .B(n8604), .ZN(n7572) );
  NAND2_X1 U9316 ( .A1(n7573), .A2(n7572), .ZN(n8595) );
  OAI21_X1 U9317 ( .B1(n7573), .B2(n7572), .A(n8595), .ZN(n7590) );
  AOI21_X1 U9318 ( .B1(n7577), .B2(n7576), .A(n8588), .ZN(n7578) );
  NOR2_X1 U9319 ( .A1(n7578), .A2(n9825), .ZN(n7589) );
  INV_X1 U9320 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n9988) );
  OR2_X1 U9321 ( .A1(n7580), .A2(n7579), .ZN(n7581) );
  XNOR2_X1 U9322 ( .A(n8604), .B(n8603), .ZN(n7583) );
  NOR2_X1 U9323 ( .A1(n7584), .A2(n7583), .ZN(n8605) );
  AOI21_X1 U9324 ( .B1(n7584), .B2(n7583), .A(n8605), .ZN(n7585) );
  OR2_X1 U9325 ( .A1(n7585), .A2(n9829), .ZN(n7587) );
  NOR2_X1 U9326 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5117), .ZN(n7696) );
  AOI21_X1 U9327 ( .B1(n8600), .B2(n8604), .A(n7696), .ZN(n7586) );
  OAI211_X1 U9328 ( .C1(n9988), .C2(n9783), .A(n7587), .B(n7586), .ZN(n7588)
         );
  AOI211_X1 U9329 ( .C1(n7590), .C2(n9832), .A(n7589), .B(n7588), .ZN(n7591)
         );
  INV_X1 U9330 ( .A(n7591), .ZN(P2_U3195) );
  INV_X1 U9331 ( .A(n7592), .ZN(n7595) );
  OAI222_X1 U9332 ( .A1(n9536), .A2(n7594), .B1(n7754), .B2(n7595), .C1(
        P1_U3086), .C2(n7593), .ZN(P1_U3333) );
  OAI222_X1 U9333 ( .A1(n7596), .A2(P2_U3151), .B1(n8205), .B2(n7595), .C1(
        n8968), .C2(n5463), .ZN(P2_U3273) );
  XNOR2_X1 U9334 ( .A(n7597), .B(n7950), .ZN(n9545) );
  INV_X1 U9335 ( .A(n9545), .ZN(n7613) );
  OAI211_X1 U9336 ( .C1(n7600), .C2(n7599), .A(n9666), .B(n7598), .ZN(n7601)
         );
  INV_X1 U9337 ( .A(n7601), .ZN(n9544) );
  AOI21_X1 U9338 ( .B1(n7602), .B2(n7609), .A(n9562), .ZN(n7603) );
  NAND2_X1 U9339 ( .A1(n7603), .A2(n7662), .ZN(n9541) );
  NAND2_X1 U9340 ( .A1(n9404), .A2(n9694), .ZN(n7607) );
  INV_X1 U9341 ( .A(n7604), .ZN(n9111) );
  NOR2_X1 U9342 ( .A1(n9402), .A2(n9111), .ZN(n7605) );
  AOI21_X1 U9343 ( .B1(n9571), .B2(P1_REG2_REG_15__SCAN_IN), .A(n7605), .ZN(
        n7606) );
  OAI211_X1 U9344 ( .C1(n9497), .C2(n9407), .A(n7607), .B(n7606), .ZN(n7608)
         );
  AOI21_X1 U9345 ( .B1(n7609), .B2(n9578), .A(n7608), .ZN(n7610) );
  OAI21_X1 U9346 ( .B1(n9541), .B2(n9331), .A(n7610), .ZN(n7611) );
  AOI21_X1 U9347 ( .B1(n9544), .B2(n9393), .A(n7611), .ZN(n7612) );
  OAI21_X1 U9348 ( .B1(n7613), .B2(n9414), .A(n7612), .ZN(P1_U3278) );
  NAND2_X1 U9349 ( .A1(n7617), .A2(n7616), .ZN(n7683) );
  XNOR2_X1 U9350 ( .A(n7683), .B(n8582), .ZN(n7647) );
  XNOR2_X1 U9351 ( .A(n9921), .B(n8170), .ZN(n7678) );
  XNOR2_X1 U9352 ( .A(n7647), .B(n7678), .ZN(n7625) );
  AOI21_X1 U9353 ( .B1(n8583), .B2(n8319), .A(n7618), .ZN(n7622) );
  INV_X1 U9354 ( .A(n7619), .ZN(n7620) );
  NAND2_X1 U9355 ( .A1(n8323), .A2(n7620), .ZN(n7621) );
  OAI211_X1 U9356 ( .C1(n7675), .C2(n8321), .A(n7622), .B(n7621), .ZN(n7623)
         );
  AOI21_X1 U9357 ( .B1(n9921), .B2(n8309), .A(n7623), .ZN(n7624) );
  OAI21_X1 U9358 ( .B1(n7625), .B2(n8311), .A(n7624), .ZN(P2_U3157) );
  NAND2_X1 U9359 ( .A1(n7629), .A2(n8963), .ZN(n7626) );
  OAI211_X1 U9360 ( .C1(n7627), .C2(n8968), .A(n7626), .B(n8571), .ZN(P2_U3272) );
  NAND2_X1 U9361 ( .A1(n7629), .A2(n7628), .ZN(n7630) );
  OAI211_X1 U9362 ( .C1(n7631), .C2(n9536), .A(n7630), .B(n8073), .ZN(P1_U3332) );
  INV_X1 U9363 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7634) );
  NAND2_X1 U9364 ( .A1(n8460), .A2(n8461), .ZN(n8366) );
  XNOR2_X1 U9365 ( .A(n7632), .B(n8459), .ZN(n7633) );
  AOI222_X1 U9366 ( .A1(n9851), .A2(n7633), .B1(n8577), .B2(n9853), .C1(n8579), 
        .C2(n9855), .ZN(n7640) );
  MUX2_X1 U9367 ( .A(n7634), .B(n7640), .S(n9931), .Z(n7637) );
  XNOR2_X1 U9368 ( .A(n7635), .B(n8459), .ZN(n7644) );
  AOI22_X1 U9369 ( .A1(n7644), .A2(n8953), .B1(n8952), .B2(n7730), .ZN(n7636)
         );
  NAND2_X1 U9370 ( .A1(n7637), .A2(n7636), .ZN(P2_U3432) );
  MUX2_X1 U9371 ( .A(n8589), .B(n7640), .S(n9947), .Z(n7639) );
  AOI22_X1 U9372 ( .A1(n7644), .A2(n8876), .B1(n8875), .B2(n7730), .ZN(n7638)
         );
  NAND2_X1 U9373 ( .A1(n7639), .A2(n7638), .ZN(P2_U3473) );
  INV_X1 U9374 ( .A(n7640), .ZN(n7643) );
  INV_X1 U9375 ( .A(n7730), .ZN(n7641) );
  OAI22_X1 U9376 ( .A1(n7641), .A2(n8742), .B1(n7728), .B2(n9862), .ZN(n7642)
         );
  OAI21_X1 U9377 ( .B1(n7643), .B2(n7642), .A(n9868), .ZN(n7646) );
  AOI22_X1 U9378 ( .A1(n7644), .A2(n9845), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9871), .ZN(n7645) );
  NAND2_X1 U9379 ( .A1(n7646), .A2(n7645), .ZN(P2_U3219) );
  INV_X1 U9380 ( .A(n7678), .ZN(n7676) );
  OAI22_X1 U9381 ( .A1(n7647), .A2(n7676), .B1(n7683), .B2(n8582), .ZN(n7649)
         );
  XNOR2_X1 U9382 ( .A(n9929), .B(n8170), .ZN(n7680) );
  XNOR2_X1 U9383 ( .A(n7680), .B(n7675), .ZN(n7648) );
  XNOR2_X1 U9384 ( .A(n7649), .B(n7648), .ZN(n7656) );
  NOR2_X1 U9385 ( .A1(n7674), .A2(n8306), .ZN(n7650) );
  AOI211_X1 U9386 ( .C1(n8303), .C2(n8580), .A(n7651), .B(n7650), .ZN(n7652)
         );
  OAI21_X1 U9387 ( .B1(n7653), .B2(n7727), .A(n7652), .ZN(n7654) );
  AOI21_X1 U9388 ( .B1(n9929), .B2(n8309), .A(n7654), .ZN(n7655) );
  OAI21_X1 U9389 ( .B1(n7656), .B2(n8311), .A(n7655), .ZN(P2_U3176) );
  XNOR2_X1 U9390 ( .A(n7657), .B(n7952), .ZN(n9509) );
  OAI211_X1 U9391 ( .C1(n7659), .C2(n7952), .A(n7658), .B(n9666), .ZN(n7661)
         );
  AOI22_X1 U9392 ( .A1(n9381), .A2(n9695), .B1(n9659), .B2(n9121), .ZN(n7660)
         );
  NAND2_X1 U9393 ( .A1(n7661), .A2(n7660), .ZN(n9505) );
  NAND2_X1 U9394 ( .A1(n7662), .A2(n9507), .ZN(n7663) );
  NAND2_X1 U9395 ( .A1(n7663), .A2(n9581), .ZN(n7664) );
  NOR2_X1 U9396 ( .A1(n9396), .A2(n7664), .ZN(n9506) );
  NAND2_X1 U9397 ( .A1(n9506), .A2(n9585), .ZN(n7666) );
  AOI22_X1 U9398 ( .A1(n9571), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9015), .B2(
        n9573), .ZN(n7665) );
  OAI211_X1 U9399 ( .C1(n9022), .C2(n9369), .A(n7666), .B(n7665), .ZN(n7667)
         );
  AOI21_X1 U9400 ( .B1(n9505), .B2(n9393), .A(n7667), .ZN(n7668) );
  OAI21_X1 U9401 ( .B1(n9509), .B2(n9414), .A(n7668), .ZN(P1_U3277) );
  NOR2_X1 U9402 ( .A1(n7675), .A2(n8306), .ZN(n7669) );
  AOI211_X1 U9403 ( .C1(n8303), .C2(n8579), .A(n7670), .B(n7669), .ZN(n7671)
         );
  OAI21_X1 U9404 ( .B1(n7672), .B2(n7727), .A(n7671), .ZN(n7687) );
  XNOR2_X1 U9405 ( .A(n7688), .B(n8170), .ZN(n7690) );
  XNOR2_X1 U9406 ( .A(n7690), .B(n7673), .ZN(n7685) );
  AOI22_X1 U9407 ( .A1(n7680), .A2(n7675), .B1(n7674), .B2(n7678), .ZN(n7682)
         );
  AOI21_X1 U9408 ( .B1(n7676), .B2(n8582), .A(n8581), .ZN(n7679) );
  NAND2_X1 U9409 ( .A1(n8582), .A2(n8581), .ZN(n7677) );
  OAI22_X1 U9410 ( .A1(n7680), .A2(n7679), .B1(n7678), .B2(n7677), .ZN(n7681)
         );
  AOI211_X1 U9411 ( .C1(n7685), .C2(n7684), .A(n8311), .B(n7691), .ZN(n7686)
         );
  AOI211_X1 U9412 ( .C1(n7688), .C2(n8309), .A(n7687), .B(n7686), .ZN(n7689)
         );
  INV_X1 U9413 ( .A(n7689), .ZN(P2_U3164) );
  INV_X1 U9414 ( .A(n7690), .ZN(n7692) );
  XNOR2_X1 U9415 ( .A(n8451), .B(n8170), .ZN(n7721) );
  XNOR2_X1 U9416 ( .A(n7721), .B(n8579), .ZN(n7693) );
  OAI21_X1 U9417 ( .B1(n4440), .B2(n7693), .A(n7724), .ZN(n7694) );
  NAND2_X1 U9418 ( .A1(n7694), .A2(n8316), .ZN(n7701) );
  INV_X1 U9419 ( .A(n7695), .ZN(n7699) );
  AOI21_X1 U9420 ( .B1(n8580), .B2(n8319), .A(n7696), .ZN(n7697) );
  OAI21_X1 U9421 ( .B1(n7756), .B2(n8321), .A(n7697), .ZN(n7698) );
  AOI21_X1 U9422 ( .B1(n7699), .B2(n8323), .A(n7698), .ZN(n7700) );
  OAI211_X1 U9423 ( .C1(n7702), .C2(n8326), .A(n7701), .B(n7700), .ZN(P2_U3174) );
  XNOR2_X1 U9424 ( .A(n7761), .B(n8577), .ZN(n8463) );
  XNOR2_X1 U9425 ( .A(n7703), .B(n8463), .ZN(n7715) );
  INV_X1 U9426 ( .A(n7715), .ZN(n7710) );
  XOR2_X1 U9427 ( .A(n7704), .B(n8463), .Z(n7705) );
  AOI222_X1 U9428 ( .A1(n9851), .A2(n7705), .B1(n8826), .B2(n9853), .C1(n8578), 
        .C2(n9855), .ZN(n7714) );
  MUX2_X1 U9429 ( .A(n7706), .B(n7714), .S(n9868), .Z(n7709) );
  INV_X1 U9430 ( .A(n7707), .ZN(n7766) );
  AOI22_X1 U9431 ( .A1(n7761), .A2(n9842), .B1(n9843), .B2(n7766), .ZN(n7708)
         );
  OAI211_X1 U9432 ( .C1(n7710), .C2(n8833), .A(n7709), .B(n7708), .ZN(P2_U3218) );
  INV_X1 U9433 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7711) );
  MUX2_X1 U9434 ( .A(n7711), .B(n7714), .S(n9931), .Z(n7713) );
  AOI22_X1 U9435 ( .A1(n7715), .A2(n8953), .B1(n8952), .B2(n7761), .ZN(n7712)
         );
  NAND2_X1 U9436 ( .A1(n7713), .A2(n7712), .ZN(P2_U3435) );
  MUX2_X1 U9437 ( .A(n8590), .B(n7714), .S(n9947), .Z(n7717) );
  AOI22_X1 U9438 ( .A1(n7715), .A2(n8876), .B1(n8875), .B2(n7761), .ZN(n7716)
         );
  NAND2_X1 U9439 ( .A1(n7717), .A2(n7716), .ZN(P2_U3474) );
  INV_X1 U9440 ( .A(n7718), .ZN(n8125) );
  OAI222_X1 U9441 ( .A1(n7720), .A2(P1_U3086), .B1(n7754), .B2(n8125), .C1(
        n7719), .C2(n9536), .ZN(P1_U3331) );
  XNOR2_X1 U9442 ( .A(n7730), .B(n8170), .ZN(n7757) );
  XNOR2_X1 U9443 ( .A(n7757), .B(n8578), .ZN(n7759) );
  XOR2_X1 U9444 ( .A(n7760), .B(n7759), .Z(n7732) );
  INV_X1 U9445 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10185) );
  OAI22_X1 U9446 ( .A1(n8258), .A2(n8321), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10185), .ZN(n7725) );
  AOI21_X1 U9447 ( .B1(n8319), .B2(n8579), .A(n7725), .ZN(n7726) );
  OAI21_X1 U9448 ( .B1(n7728), .B2(n7727), .A(n7726), .ZN(n7729) );
  AOI21_X1 U9449 ( .B1(n7730), .B2(n8309), .A(n7729), .ZN(n7731) );
  OAI21_X1 U9450 ( .B1(n7732), .B2(n8311), .A(n7731), .ZN(P2_U3155) );
  XNOR2_X1 U9451 ( .A(n7733), .B(n8468), .ZN(n7747) );
  INV_X1 U9452 ( .A(n7747), .ZN(n7742) );
  XNOR2_X1 U9453 ( .A(n7734), .B(n8468), .ZN(n7737) );
  NAND2_X1 U9454 ( .A1(n8577), .A2(n9855), .ZN(n7735) );
  OAI21_X1 U9455 ( .B1(n8307), .B2(n8703), .A(n7735), .ZN(n7736) );
  AOI21_X1 U9456 ( .B1(n7737), .B2(n9851), .A(n7736), .ZN(n7746) );
  MUX2_X1 U9457 ( .A(n7738), .B(n7746), .S(n9868), .Z(n7741) );
  INV_X1 U9458 ( .A(n7739), .ZN(n8255) );
  AOI22_X1 U9459 ( .A1(n8260), .A2(n9842), .B1(n9843), .B2(n8255), .ZN(n7740)
         );
  OAI211_X1 U9460 ( .C1(n7742), .C2(n8833), .A(n7741), .B(n7740), .ZN(P2_U3217) );
  INV_X1 U9461 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7743) );
  MUX2_X1 U9462 ( .A(n7743), .B(n7746), .S(n9931), .Z(n7745) );
  AOI22_X1 U9463 ( .A1(n7747), .A2(n8953), .B1(n8952), .B2(n8260), .ZN(n7744)
         );
  NAND2_X1 U9464 ( .A1(n7745), .A2(n7744), .ZN(P2_U3438) );
  MUX2_X1 U9465 ( .A(n8645), .B(n7746), .S(n9947), .Z(n7749) );
  AOI22_X1 U9466 ( .A1(n7747), .A2(n8876), .B1(n8875), .B2(n8260), .ZN(n7748)
         );
  NAND2_X1 U9467 ( .A1(n7749), .A2(n7748), .ZN(P2_U3475) );
  INV_X1 U9468 ( .A(n7750), .ZN(n7753) );
  OAI222_X1 U9469 ( .A1(n5625), .A2(P2_U3151), .B1(n8205), .B2(n7753), .C1(
        n7751), .C2(n8968), .ZN(P2_U3270) );
  OAI222_X1 U9470 ( .A1(n7755), .A2(P1_U3086), .B1(n7754), .B2(n7753), .C1(
        n7752), .C2(n9536), .ZN(P1_U3330) );
  INV_X1 U9471 ( .A(n7761), .ZN(n7769) );
  XNOR2_X1 U9472 ( .A(n7761), .B(n8170), .ZN(n8128) );
  XNOR2_X1 U9473 ( .A(n8128), .B(n8577), .ZN(n7762) );
  NAND2_X1 U9474 ( .A1(n7763), .A2(n7762), .ZN(n8130) );
  OAI211_X1 U9475 ( .C1(n7763), .C2(n7762), .A(n8130), .B(n8316), .ZN(n7768)
         );
  NAND2_X1 U9476 ( .A1(n8319), .A2(n8578), .ZN(n7764) );
  NAND2_X1 U9477 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8601) );
  OAI211_X1 U9478 ( .C1(n8269), .C2(n8321), .A(n7764), .B(n8601), .ZN(n7765)
         );
  AOI21_X1 U9479 ( .B1(n7766), .B2(n8323), .A(n7765), .ZN(n7767) );
  OAI211_X1 U9480 ( .C1(n7769), .C2(n8326), .A(n7768), .B(n7767), .ZN(P2_U3181) );
  INV_X1 U9481 ( .A(n7770), .ZN(n7774) );
  OAI222_X1 U9482 ( .A1(n7772), .A2(P2_U3151), .B1(n8205), .B2(n7774), .C1(
        n7771), .C2(n8968), .ZN(P2_U3269) );
  OAI222_X1 U9483 ( .A1(n7775), .A2(P1_U3086), .B1(n7754), .B2(n7774), .C1(
        n7773), .C2(n9536), .ZN(P1_U3329) );
  INV_X1 U9484 ( .A(n7777), .ZN(n7778) );
  AOI21_X1 U9485 ( .B1(n7779), .B2(n7776), .A(n7778), .ZN(n7785) );
  AOI22_X1 U9486 ( .A1(n9058), .A2(n7780), .B1(n9102), .B2(n9121), .ZN(n7782)
         );
  OAI211_X1 U9487 ( .C1(n9706), .C2(n9070), .A(n7782), .B(n7781), .ZN(n7783)
         );
  AOI21_X1 U9488 ( .B1(n9709), .B2(n9084), .A(n7783), .ZN(n7784) );
  OAI21_X1 U9489 ( .B1(n7785), .B2(n9075), .A(n7784), .ZN(P1_U3215) );
  INV_X1 U9490 ( .A(n8964), .ZN(n7786) );
  OAI222_X1 U9491 ( .A1(n9536), .A2(n7787), .B1(P1_U3086), .B2(n6269), .C1(
        n7754), .C2(n7786), .ZN(P1_U3327) );
  INV_X1 U9492 ( .A(n7789), .ZN(n7790) );
  AOI21_X1 U9493 ( .B1(n7791), .B2(n7788), .A(n7790), .ZN(n7795) );
  AOI22_X1 U9494 ( .A1(n9081), .A2(n9127), .B1(n9102), .B2(n9125), .ZN(n7794)
         );
  AOI22_X1 U9495 ( .A1(n9084), .A2(n7792), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9082), .ZN(n7793) );
  OAI211_X1 U9496 ( .C1(n7795), .C2(n9075), .A(n7794), .B(n7793), .ZN(P1_U3222) );
  NAND4_X1 U9497 ( .A1(n7962), .A2(n7926), .A3(n7964), .A4(n7965), .ZN(n7897)
         );
  NAND2_X1 U9498 ( .A1(n8008), .A2(n7798), .ZN(n7797) );
  AND2_X1 U9499 ( .A1(n7798), .A2(n7813), .ZN(n8009) );
  NAND2_X1 U9500 ( .A1(n7810), .A2(n7815), .ZN(n8012) );
  AOI21_X1 U9501 ( .B1(n7812), .B2(n8009), .A(n8012), .ZN(n7800) );
  NAND2_X1 U9502 ( .A1(n7818), .A2(n8013), .ZN(n7799) );
  OAI21_X1 U9503 ( .B1(n7800), .B2(n7799), .A(n7937), .ZN(n7802) );
  INV_X1 U9504 ( .A(n7817), .ZN(n7801) );
  NAND2_X1 U9505 ( .A1(n7802), .A2(n7801), .ZN(n7805) );
  NAND3_X1 U9506 ( .A1(n7805), .A2(n7804), .A3(n7803), .ZN(n7807) );
  NAND2_X1 U9507 ( .A1(n7807), .A2(n7806), .ZN(n7822) );
  INV_X1 U9508 ( .A(n7808), .ZN(n7811) );
  OAI211_X1 U9509 ( .C1(n7812), .C2(n7811), .A(n7810), .B(n7809), .ZN(n7814)
         );
  NAND3_X1 U9510 ( .A1(n7814), .A2(n8013), .A3(n7813), .ZN(n7816) );
  INV_X1 U9511 ( .A(n7829), .ZN(n7825) );
  INV_X1 U9512 ( .A(n7823), .ZN(n7824) );
  OAI21_X1 U9513 ( .B1(n7825), .B2(n7824), .A(n7830), .ZN(n7827) );
  AOI21_X1 U9514 ( .B1(n7829), .B2(n7828), .A(n8020), .ZN(n7832) );
  NAND2_X1 U9515 ( .A1(n7831), .A2(n7830), .ZN(n8024) );
  AND2_X1 U9516 ( .A1(n7834), .A2(n7833), .ZN(n8023) );
  NAND2_X1 U9517 ( .A1(n7835), .A2(n8026), .ZN(n7837) );
  NAND2_X1 U9518 ( .A1(n7843), .A2(n7836), .ZN(n8031) );
  AOI21_X1 U9519 ( .B1(n7837), .B2(n7948), .A(n8031), .ZN(n7839) );
  OAI211_X1 U9520 ( .C1(n8031), .C2(n7838), .A(n7846), .B(n7841), .ZN(n8034)
         );
  OAI21_X1 U9521 ( .B1(n7839), .B2(n8034), .A(n8032), .ZN(n7849) );
  NAND3_X1 U9522 ( .A1(n7842), .A2(n7841), .A3(n8028), .ZN(n7844) );
  NAND2_X1 U9523 ( .A1(n7844), .A2(n7843), .ZN(n7847) );
  AOI21_X1 U9524 ( .B1(n7847), .B2(n7846), .A(n7845), .ZN(n7848) );
  AND2_X1 U9525 ( .A1(n7852), .A2(n7851), .ZN(n8004) );
  NAND2_X1 U9526 ( .A1(n7853), .A2(n8004), .ZN(n7856) );
  AND2_X1 U9527 ( .A1(n7982), .A2(n7854), .ZN(n8003) );
  NAND2_X1 U9528 ( .A1(n7859), .A2(n8039), .ZN(n7855) );
  AOI21_X1 U9529 ( .B1(n7856), .B2(n8003), .A(n7855), .ZN(n7857) );
  NAND2_X1 U9530 ( .A1(n7858), .A2(n7926), .ZN(n7862) );
  NAND2_X1 U9531 ( .A1(n7863), .A2(n7859), .ZN(n7973) );
  OR2_X1 U9532 ( .A1(n9479), .A2(n9071), .ZN(n7864) );
  NAND2_X1 U9533 ( .A1(n7864), .A2(n7860), .ZN(n8002) );
  MUX2_X1 U9534 ( .A(n7973), .B(n8002), .S(n8070), .Z(n7861) );
  INV_X1 U9535 ( .A(n7863), .ZN(n7865) );
  INV_X1 U9536 ( .A(n7864), .ZN(n7978) );
  MUX2_X1 U9537 ( .A(n7865), .B(n7978), .S(n7926), .Z(n7866) );
  OR2_X1 U9538 ( .A1(n9328), .A2(n9460), .ZN(n7867) );
  NAND2_X1 U9539 ( .A1(n7871), .A2(n7867), .ZN(n7967) );
  NAND2_X1 U9540 ( .A1(n7966), .A2(n7868), .ZN(n7974) );
  MUX2_X1 U9541 ( .A(n7967), .B(n7974), .S(n8070), .Z(n7869) );
  INV_X1 U9542 ( .A(n7869), .ZN(n7870) );
  INV_X1 U9543 ( .A(n7966), .ZN(n7873) );
  INV_X1 U9544 ( .A(n7871), .ZN(n7872) );
  MUX2_X1 U9545 ( .A(n7873), .B(n7872), .S(n8070), .Z(n7874) );
  NOR2_X1 U9546 ( .A1(n9289), .A2(n7874), .ZN(n7875) );
  MUX2_X1 U9547 ( .A(n7976), .B(n7969), .S(n7926), .Z(n7876) );
  NAND2_X1 U9548 ( .A1(n7877), .A2(n7876), .ZN(n7892) );
  INV_X1 U9549 ( .A(n7892), .ZN(n7879) );
  NAND2_X1 U9550 ( .A1(n8044), .A2(n7878), .ZN(n7891) );
  AOI21_X1 U9551 ( .B1(n7879), .B2(n7972), .A(n7891), .ZN(n7896) );
  NOR2_X1 U9552 ( .A1(n9238), .A2(n8070), .ZN(n7883) );
  NOR2_X1 U9553 ( .A1(n9120), .A2(n8070), .ZN(n7880) );
  AOI21_X1 U9554 ( .B1(n9433), .B2(n7883), .A(n7880), .ZN(n7889) );
  NAND2_X1 U9555 ( .A1(n9238), .A2(n8070), .ZN(n7882) );
  OAI22_X1 U9556 ( .A1(n9433), .A2(n7882), .B1(n9429), .B2(n7926), .ZN(n7881)
         );
  NAND2_X1 U9557 ( .A1(n6370), .A2(n7881), .ZN(n7888) );
  NOR2_X1 U9558 ( .A1(n7882), .A2(n9429), .ZN(n7886) );
  NAND2_X1 U9559 ( .A1(n7883), .A2(n9429), .ZN(n7884) );
  NAND2_X1 U9560 ( .A1(n9433), .A2(n7884), .ZN(n7885) );
  OAI21_X1 U9561 ( .B1(n9433), .B2(n7886), .A(n7885), .ZN(n7887) );
  OAI211_X1 U9562 ( .C1(n6370), .C2(n7889), .A(n7888), .B(n7887), .ZN(n7890)
         );
  INV_X1 U9563 ( .A(n7890), .ZN(n7895) );
  AOI21_X1 U9564 ( .B1(n7892), .B2(n7972), .A(n7891), .ZN(n7894) );
  OR2_X1 U9565 ( .A1(n7957), .A2(n7898), .ZN(n7900) );
  MUX2_X1 U9566 ( .A(n7990), .B(n7963), .S(n8070), .Z(n7899) );
  NAND2_X1 U9567 ( .A1(n7900), .A2(n7899), .ZN(n7927) );
  INV_X1 U9568 ( .A(n7902), .ZN(n7903) );
  OR2_X1 U9569 ( .A1(n7904), .A2(n7903), .ZN(n7905) );
  INV_X1 U9570 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9537) );
  MUX2_X1 U9571 ( .A(n9537), .B(n8127), .S(n7917), .Z(n7906) );
  NAND2_X1 U9572 ( .A1(n7906), .A2(n10146), .ZN(n7915) );
  INV_X1 U9573 ( .A(n7906), .ZN(n7907) );
  NAND2_X1 U9574 ( .A1(n7907), .A2(SI_30_), .ZN(n7908) );
  NAND2_X1 U9575 ( .A1(n7915), .A2(n7908), .ZN(n7909) );
  NAND2_X1 U9576 ( .A1(n7910), .A2(n7909), .ZN(n7911) );
  NAND2_X1 U9577 ( .A1(n7916), .A2(n7911), .ZN(n8330) );
  NAND2_X1 U9578 ( .A1(n8330), .A2(n7912), .ZN(n7914) );
  OR2_X1 U9579 ( .A1(n5784), .A2(n9537), .ZN(n7913) );
  MUX2_X1 U9580 ( .A(n8070), .B(n7927), .S(n8087), .Z(n7925) );
  MUX2_X1 U9581 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7917), .Z(n7919) );
  INV_X1 U9582 ( .A(SI_31_), .ZN(n7918) );
  XNOR2_X1 U9583 ( .A(n7919), .B(n7918), .ZN(n7920) );
  MUX2_X1 U9584 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8957), .S(n4713), .Z(n7924) );
  NAND3_X1 U9585 ( .A1(n7925), .A2(n9225), .A3(n7931), .ZN(n7930) );
  MUX2_X1 U9586 ( .A(n7927), .B(n7926), .S(n8087), .Z(n7928) );
  NAND2_X1 U9587 ( .A1(n9416), .A2(n8091), .ZN(n8071) );
  NAND2_X1 U9588 ( .A1(n8091), .A2(n7931), .ZN(n7992) );
  NAND3_X1 U9589 ( .A1(n7928), .A2(n8071), .A3(n7992), .ZN(n7929) );
  OR2_X1 U9590 ( .A1(n9416), .A2(n8091), .ZN(n8069) );
  INV_X1 U9591 ( .A(n7931), .ZN(n8060) );
  XNOR2_X1 U9592 ( .A(n8087), .B(n8060), .ZN(n7959) );
  INV_X1 U9593 ( .A(n9320), .ZN(n9318) );
  NAND4_X1 U9594 ( .A1(n7934), .A2(n7933), .A3(n6923), .A4(n7932), .ZN(n7936)
         );
  NOR2_X1 U9595 ( .A1(n7936), .A2(n7935), .ZN(n7940) );
  AND4_X1 U9596 ( .A1(n7940), .A2(n7939), .A3(n7938), .A4(n7937), .ZN(n7941)
         );
  NAND4_X1 U9597 ( .A1(n4897), .A2(n7942), .A3(n8017), .A4(n7941), .ZN(n7943)
         );
  NOR2_X1 U9598 ( .A1(n7944), .A2(n7943), .ZN(n7945) );
  NAND4_X1 U9599 ( .A1(n7948), .A2(n7947), .A3(n7946), .A4(n7945), .ZN(n7949)
         );
  NOR2_X1 U9600 ( .A1(n7950), .A2(n7949), .ZN(n7951) );
  NAND3_X1 U9601 ( .A1(n9409), .A2(n7952), .A3(n7951), .ZN(n7953) );
  NOR2_X1 U9602 ( .A1(n9376), .A2(n7953), .ZN(n7954) );
  XNOR2_X1 U9603 ( .A(n9483), .B(n9362), .ZN(n9356) );
  NAND4_X1 U9604 ( .A1(n9342), .A2(n9372), .A3(n7954), .A4(n9356), .ZN(n7955)
         );
  OR4_X1 U9605 ( .A1(n9312), .A2(n9289), .A3(n9318), .A4(n7955), .ZN(n7956) );
  OR4_X1 U9606 ( .A1(n7956), .A2(n9244), .A3(n9255), .A4(n9271), .ZN(n7958) );
  NOR4_X1 U9607 ( .A1(n7959), .A2(n7958), .A3(n7957), .A4(n9229), .ZN(n7960)
         );
  AOI21_X1 U9608 ( .B1(n7961), .B2(n8006), .A(n7997), .ZN(n8001) );
  NAND2_X1 U9609 ( .A1(n7963), .A2(n7962), .ZN(n8052) );
  AND2_X1 U9610 ( .A1(n7965), .A2(n7964), .ZN(n8048) );
  NAND2_X1 U9611 ( .A1(n7967), .A2(n7966), .ZN(n7968) );
  NAND2_X1 U9612 ( .A1(n7969), .A2(n7968), .ZN(n7970) );
  NAND2_X1 U9613 ( .A1(n7970), .A2(n7976), .ZN(n7971) );
  AND2_X1 U9614 ( .A1(n7972), .A2(n7971), .ZN(n7981) );
  INV_X1 U9615 ( .A(n7973), .ZN(n7977) );
  INV_X1 U9616 ( .A(n7974), .ZN(n7975) );
  OAI211_X1 U9617 ( .C1(n7978), .C2(n7977), .A(n7976), .B(n7975), .ZN(n7980)
         );
  AOI21_X1 U9618 ( .B1(n7981), .B2(n7980), .A(n7979), .ZN(n8050) );
  INV_X1 U9619 ( .A(n7981), .ZN(n8046) );
  NAND2_X1 U9620 ( .A1(n7983), .A2(n7982), .ZN(n9348) );
  OR3_X1 U9621 ( .A1(n8046), .A2(n8002), .A3(n9348), .ZN(n7984) );
  NAND3_X1 U9622 ( .A1(n8050), .A2(n8044), .A3(n7984), .ZN(n7985) );
  AND2_X1 U9623 ( .A1(n8048), .A2(n7985), .ZN(n7988) );
  NAND2_X1 U9624 ( .A1(n7987), .A2(n7986), .ZN(n8055) );
  NOR2_X1 U9625 ( .A1(n7988), .A2(n8055), .ZN(n7989) );
  NOR2_X1 U9626 ( .A1(n8052), .A2(n7989), .ZN(n7993) );
  NAND2_X1 U9627 ( .A1(n8087), .A2(n8060), .ZN(n7991) );
  NAND2_X1 U9628 ( .A1(n7991), .A2(n7990), .ZN(n8056) );
  OAI22_X1 U9629 ( .A1(n7993), .A2(n8056), .B1(n8087), .B2(n7992), .ZN(n7994)
         );
  OAI211_X1 U9630 ( .C1(n9419), .C2(n8091), .A(n8071), .B(n7994), .ZN(n7996)
         );
  NAND3_X1 U9631 ( .A1(n7996), .A2(n7995), .A3(n8069), .ZN(n7999) );
  INV_X1 U9632 ( .A(n7997), .ZN(n7998) );
  NAND2_X1 U9633 ( .A1(n7999), .A2(n7998), .ZN(n8000) );
  INV_X1 U9634 ( .A(n8002), .ZN(n8043) );
  INV_X1 U9635 ( .A(n8003), .ZN(n8041) );
  INV_X1 U9636 ( .A(n8004), .ZN(n8038) );
  NAND2_X1 U9637 ( .A1(n9599), .A2(n9593), .ZN(n8005) );
  AND4_X1 U9638 ( .A1(n8008), .A2(n8007), .A3(n8006), .A4(n8005), .ZN(n8010)
         );
  OAI21_X1 U9639 ( .B1(n8011), .B2(n8010), .A(n8009), .ZN(n8016) );
  INV_X1 U9640 ( .A(n8012), .ZN(n8015) );
  INV_X1 U9641 ( .A(n8013), .ZN(n8014) );
  AOI21_X1 U9642 ( .B1(n8016), .B2(n8015), .A(n8014), .ZN(n8018) );
  OAI21_X1 U9643 ( .B1(n8018), .B2(n4799), .A(n8017), .ZN(n8022) );
  INV_X1 U9644 ( .A(n8019), .ZN(n8021) );
  AOI21_X1 U9645 ( .B1(n8022), .B2(n8021), .A(n8020), .ZN(n8025) );
  OAI21_X1 U9646 ( .B1(n8025), .B2(n8024), .A(n8023), .ZN(n8027) );
  NAND3_X1 U9647 ( .A1(n8027), .A2(n8026), .A3(n4375), .ZN(n8029) );
  AND2_X1 U9648 ( .A1(n8029), .A2(n8028), .ZN(n8030) );
  NOR2_X1 U9649 ( .A1(n8031), .A2(n8030), .ZN(n8033) );
  OAI21_X1 U9650 ( .B1(n8034), .B2(n8033), .A(n8032), .ZN(n8036) );
  AND2_X1 U9651 ( .A1(n8036), .A2(n8035), .ZN(n8037) );
  NOR2_X1 U9652 ( .A1(n8038), .A2(n8037), .ZN(n8040) );
  OAI21_X1 U9653 ( .B1(n8041), .B2(n8040), .A(n8039), .ZN(n8042) );
  NAND2_X1 U9654 ( .A1(n8043), .A2(n8042), .ZN(n8045) );
  OAI21_X1 U9655 ( .B1(n8046), .B2(n8045), .A(n8044), .ZN(n8047) );
  INV_X1 U9656 ( .A(n8047), .ZN(n8051) );
  INV_X1 U9657 ( .A(n8048), .ZN(n8049) );
  AOI21_X1 U9658 ( .B1(n8051), .B2(n8050), .A(n8049), .ZN(n8054) );
  INV_X1 U9659 ( .A(n8052), .ZN(n8053) );
  OAI21_X1 U9660 ( .B1(n8055), .B2(n8054), .A(n8053), .ZN(n8058) );
  INV_X1 U9661 ( .A(n8056), .ZN(n8057) );
  NAND2_X1 U9662 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  OAI21_X1 U9663 ( .B1(n8060), .B2(n8087), .A(n8059), .ZN(n8061) );
  NAND2_X1 U9664 ( .A1(n8061), .A2(n8071), .ZN(n8062) );
  NAND2_X1 U9665 ( .A1(n8062), .A2(n8069), .ZN(n8066) );
  OR2_X1 U9666 ( .A1(n8066), .A2(n8063), .ZN(n8065) );
  AOI21_X1 U9667 ( .B1(n8066), .B2(n8079), .A(n8073), .ZN(n8067) );
  OAI21_X1 U9668 ( .B1(n8070), .B2(n8069), .A(n8068), .ZN(n8084) );
  INV_X1 U9669 ( .A(n8071), .ZN(n8076) );
  NOR2_X1 U9670 ( .A1(n8073), .A2(n8072), .ZN(n8077) );
  NAND2_X1 U9671 ( .A1(n8077), .A2(n8074), .ZN(n8075) );
  AOI21_X1 U9672 ( .B1(n8076), .B2(n8108), .A(n8075), .ZN(n8083) );
  INV_X1 U9673 ( .A(n8077), .ZN(n8078) );
  AND2_X1 U9674 ( .A1(n8078), .A2(P1_B_REG_SCAN_IN), .ZN(n8082) );
  NAND4_X1 U9675 ( .A1(n8080), .A2(n8079), .A3(n9659), .A4(n9138), .ZN(n8081)
         );
  AOI22_X1 U9676 ( .A1(n8084), .A2(n8083), .B1(n8082), .B2(n8081), .ZN(n8085)
         );
  INV_X1 U9677 ( .A(n8086), .ZN(n8089) );
  INV_X1 U9678 ( .A(n9222), .ZN(n8088) );
  OAI211_X1 U9679 ( .C1(n9419), .C2(n8089), .A(n8088), .B(n9581), .ZN(n9418)
         );
  NAND2_X1 U9680 ( .A1(n8091), .A2(n8090), .ZN(n9417) );
  NOR2_X1 U9681 ( .A1(n9571), .A2(n9417), .ZN(n9224) );
  NOR2_X1 U9682 ( .A1(n9419), .A2(n9369), .ZN(n8092) );
  AOI211_X1 U9683 ( .C1(n9571), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9224), .B(
        n8092), .ZN(n8093) );
  OAI21_X1 U9684 ( .B1(n9331), .B2(n9418), .A(n8093), .ZN(P1_U3264) );
  INV_X1 U9685 ( .A(n8094), .ZN(n8202) );
  OAI222_X1 U9686 ( .A1(n9536), .A2(n8096), .B1(P1_U3086), .B2(n8095), .C1(
        n7754), .C2(n8202), .ZN(P1_U3328) );
  AND2_X1 U9687 ( .A1(n8102), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8097) );
  OR2_X1 U9688 ( .A1(n8098), .A2(n8097), .ZN(n8100) );
  XNOR2_X1 U9689 ( .A(n8100), .B(n8099), .ZN(n8104) );
  AOI21_X1 U9690 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n8102), .A(n8101), .ZN(
        n8103) );
  XNOR2_X1 U9691 ( .A(n8103), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8105) );
  AOI22_X1 U9692 ( .A1(n8104), .A2(n9204), .B1(n9211), .B2(n8105), .ZN(n8110)
         );
  INV_X1 U9693 ( .A(n8104), .ZN(n8107) );
  OAI21_X1 U9694 ( .B1(n8105), .B2(n9165), .A(n9189), .ZN(n8106) );
  AOI21_X1 U9695 ( .B1(n8107), .B2(n9204), .A(n8106), .ZN(n8109) );
  MUX2_X1 U9696 ( .A(n8110), .B(n8109), .S(n8108), .Z(n8111) );
  NAND2_X1 U9697 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8983) );
  OAI211_X1 U9698 ( .C1(n4563), .C2(n8112), .A(n8111), .B(n8983), .ZN(P1_U3262) );
  NAND2_X1 U9699 ( .A1(n8113), .A2(n9586), .ZN(n8122) );
  NAND2_X1 U9700 ( .A1(n8114), .A2(n9578), .ZN(n8118) );
  NOR2_X1 U9701 ( .A1(n9402), .A2(n8115), .ZN(n8116) );
  AOI21_X1 U9702 ( .B1(n9571), .B2(P1_REG2_REG_29__SCAN_IN), .A(n8116), .ZN(
        n8117) );
  NAND2_X1 U9703 ( .A1(n8118), .A2(n8117), .ZN(n8119) );
  AOI21_X1 U9704 ( .B1(n8120), .B2(n9585), .A(n8119), .ZN(n8121) );
  OAI211_X1 U9705 ( .C1(n8123), .C2(n9571), .A(n8122), .B(n8121), .ZN(P1_U3356) );
  OAI222_X1 U9706 ( .A1(n5619), .A2(P2_U3151), .B1(n8205), .B2(n8125), .C1(
        n8124), .C2(n8968), .ZN(P2_U3271) );
  INV_X1 U9707 ( .A(n8330), .ZN(n9535) );
  OAI222_X1 U9708 ( .A1(n8126), .A2(P2_U3151), .B1(n8205), .B2(n9535), .C1(
        n8968), .C2(n8127), .ZN(P2_U3265) );
  XNOR2_X1 U9709 ( .A(n8260), .B(n8170), .ZN(n8132) );
  XNOR2_X1 U9710 ( .A(n8132), .B(n8269), .ZN(n8254) );
  INV_X1 U9711 ( .A(n8254), .ZN(n8131) );
  XNOR2_X1 U9712 ( .A(n8273), .B(n8170), .ZN(n8134) );
  XNOR2_X1 U9713 ( .A(n8134), .B(n8307), .ZN(n8264) );
  INV_X1 U9714 ( .A(n8134), .ZN(n8135) );
  NAND2_X1 U9715 ( .A1(n8135), .A2(n8307), .ZN(n8136) );
  NAND2_X1 U9716 ( .A1(n8263), .A2(n8136), .ZN(n8302) );
  XNOR2_X1 U9717 ( .A(n8944), .B(n8170), .ZN(n8138) );
  XNOR2_X1 U9718 ( .A(n8138), .B(n8827), .ZN(n8301) );
  NAND2_X1 U9719 ( .A1(n8302), .A2(n8301), .ZN(n8140) );
  NAND2_X1 U9720 ( .A1(n8138), .A2(n8137), .ZN(n8139) );
  XNOR2_X1 U9721 ( .A(n8867), .B(n4456), .ZN(n8223) );
  NOR2_X1 U9722 ( .A1(n8223), .A2(n8817), .ZN(n8142) );
  INV_X1 U9723 ( .A(n8223), .ZN(n8141) );
  XNOR2_X1 U9724 ( .A(n8937), .B(n8170), .ZN(n8143) );
  NAND2_X1 U9725 ( .A1(n8143), .A2(n8236), .ZN(n8144) );
  OAI21_X1 U9726 ( .B1(n8143), .B2(n8236), .A(n8144), .ZN(n8284) );
  XNOR2_X1 U9727 ( .A(n8931), .B(n8170), .ZN(n8145) );
  XNOR2_X1 U9728 ( .A(n8145), .B(n8793), .ZN(n8232) );
  NAND2_X1 U9729 ( .A1(n8233), .A2(n8232), .ZN(n8231) );
  XNOR2_X1 U9730 ( .A(n8925), .B(n8170), .ZN(n8148) );
  XNOR2_X1 U9731 ( .A(n8148), .B(n8490), .ZN(n8291) );
  INV_X1 U9732 ( .A(n8145), .ZN(n8146) );
  NOR2_X1 U9733 ( .A1(n8146), .A2(n8793), .ZN(n8292) );
  NOR2_X1 U9734 ( .A1(n8291), .A2(n8292), .ZN(n8147) );
  INV_X1 U9735 ( .A(n8148), .ZN(n8149) );
  NAND2_X1 U9736 ( .A1(n8149), .A2(n8781), .ZN(n8150) );
  XNOR2_X1 U9737 ( .A(n8512), .B(n8170), .ZN(n8151) );
  NAND2_X1 U9738 ( .A1(n8152), .A2(n8151), .ZN(n8153) );
  XNOR2_X1 U9739 ( .A(n8743), .B(n4456), .ZN(n8154) );
  NAND2_X1 U9740 ( .A1(n8154), .A2(n8514), .ZN(n8241) );
  INV_X1 U9741 ( .A(n8154), .ZN(n8155) );
  NAND2_X1 U9742 ( .A1(n8155), .A2(n8757), .ZN(n8156) );
  NAND2_X1 U9743 ( .A1(n8157), .A2(n8275), .ZN(n8240) );
  NAND2_X1 U9744 ( .A1(n8240), .A2(n8241), .ZN(n8162) );
  XNOR2_X1 U9745 ( .A(n8907), .B(n8170), .ZN(n8159) );
  NAND2_X1 U9746 ( .A1(n8159), .A2(n8158), .ZN(n8163) );
  INV_X1 U9747 ( .A(n8159), .ZN(n8160) );
  NAND2_X1 U9748 ( .A1(n8160), .A2(n8745), .ZN(n8161) );
  XNOR2_X1 U9749 ( .A(n8901), .B(n8170), .ZN(n8164) );
  XNOR2_X1 U9750 ( .A(n8164), .B(n8736), .ZN(n8314) );
  XNOR2_X1 U9751 ( .A(n8216), .B(n4456), .ZN(n8167) );
  XNOR2_X1 U9752 ( .A(n8167), .B(n8702), .ZN(n8207) );
  INV_X1 U9753 ( .A(n8164), .ZN(n8165) );
  NOR2_X1 U9754 ( .A1(n8165), .A2(n8736), .ZN(n8208) );
  NOR2_X1 U9755 ( .A1(n8207), .A2(n8208), .ZN(n8166) );
  XNOR2_X1 U9756 ( .A(n8700), .B(n8170), .ZN(n8171) );
  XNOR2_X1 U9757 ( .A(n8172), .B(n8171), .ZN(n8177) );
  INV_X1 U9758 ( .A(n8576), .ZN(n8704) );
  AOI22_X1 U9759 ( .A1(n8168), .A2(n8319), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8174) );
  NAND2_X1 U9760 ( .A1(n8708), .A2(n8323), .ZN(n8173) );
  OAI211_X1 U9761 ( .C1(n8704), .C2(n8321), .A(n8174), .B(n8173), .ZN(n8175)
         );
  AOI21_X1 U9762 ( .B1(n8709), .B2(n8309), .A(n8175), .ZN(n8176) );
  OAI21_X1 U9763 ( .B1(n8177), .B2(n8311), .A(n8176), .ZN(P2_U3160) );
  NAND2_X1 U9764 ( .A1(n9424), .A2(n8178), .ZN(n8181) );
  NAND2_X1 U9765 ( .A1(n9120), .A2(n8179), .ZN(n8180) );
  NAND2_X1 U9766 ( .A1(n8181), .A2(n8180), .ZN(n8183) );
  XNOR2_X1 U9767 ( .A(n8183), .B(n8182), .ZN(n8186) );
  AOI22_X1 U9768 ( .A1(n9424), .A2(n8184), .B1(n4355), .B2(n9120), .ZN(n8185)
         );
  XNOR2_X1 U9769 ( .A(n8186), .B(n8185), .ZN(n8187) );
  INV_X1 U9770 ( .A(n8187), .ZN(n8191) );
  NAND3_X1 U9771 ( .A1(n8191), .A2(n9109), .A3(n8190), .ZN(n8196) );
  AOI22_X1 U9772 ( .A1(n9116), .A2(n9238), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8189) );
  NAND2_X1 U9773 ( .A1(n9058), .A2(n9235), .ZN(n8188) );
  OAI211_X1 U9774 ( .C1(n9113), .C2(n9421), .A(n8189), .B(n8188), .ZN(n8193)
         );
  NOR3_X1 U9775 ( .A1(n8191), .A2(n8190), .A3(n9075), .ZN(n8192) );
  AOI211_X1 U9776 ( .C1(n9424), .C2(n9084), .A(n8193), .B(n8192), .ZN(n8194)
         );
  OAI211_X1 U9777 ( .C1(n8197), .C2(n8196), .A(n8195), .B(n8194), .ZN(P1_U3220) );
  INV_X1 U9778 ( .A(n8198), .ZN(n8204) );
  OAI222_X1 U9779 ( .A1(n9536), .A2(n8200), .B1(P1_U3086), .B2(n8199), .C1(
        n7754), .C2(n8204), .ZN(P1_U3326) );
  OAI222_X1 U9780 ( .A1(P2_U3151), .A2(n8631), .B1(n8205), .B2(n8202), .C1(
        n8201), .C2(n8968), .ZN(P2_U3268) );
  OAI222_X1 U9781 ( .A1(P2_U3151), .A2(n8206), .B1(n8205), .B2(n8204), .C1(
        n8203), .C2(n8968), .ZN(P2_U3266) );
  INV_X1 U9782 ( .A(n8313), .ZN(n8209) );
  NAND3_X1 U9783 ( .A1(n8211), .A2(n8316), .A3(n8210), .ZN(n8215) );
  AOI22_X1 U9784 ( .A1(n8736), .A2(n8319), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8212) );
  OAI21_X1 U9785 ( .B1(n8539), .B2(n8321), .A(n8212), .ZN(n8213) );
  AOI21_X1 U9786 ( .B1(n8720), .B2(n8323), .A(n8213), .ZN(n8214) );
  OAI211_X1 U9787 ( .C1(n8216), .C2(n8326), .A(n8215), .B(n8214), .ZN(P2_U3154) );
  AOI21_X1 U9788 ( .B1(n8767), .B2(n8217), .A(n4378), .ZN(n8222) );
  AOI22_X1 U9789 ( .A1(n8757), .A2(n8303), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8219) );
  NAND2_X1 U9790 ( .A1(n8323), .A2(n8760), .ZN(n8218) );
  OAI211_X1 U9791 ( .C1(n8490), .C2(n8306), .A(n8219), .B(n8218), .ZN(n8220)
         );
  AOI21_X1 U9792 ( .B1(n8919), .B2(n8309), .A(n8220), .ZN(n8221) );
  OAI21_X1 U9793 ( .B1(n8222), .B2(n8311), .A(n8221), .ZN(P2_U3156) );
  XNOR2_X1 U9794 ( .A(n8223), .B(n8817), .ZN(n8224) );
  XNOR2_X1 U9795 ( .A(n8225), .B(n8224), .ZN(n8230) );
  NAND2_X1 U9796 ( .A1(n8319), .A2(n8827), .ZN(n8226) );
  NAND2_X1 U9797 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8671) );
  OAI211_X1 U9798 ( .C1(n8236), .C2(n8321), .A(n8226), .B(n8671), .ZN(n8228)
         );
  NOR2_X1 U9799 ( .A1(n8808), .A2(n8326), .ZN(n8227) );
  AOI211_X1 U9800 ( .C1(n8805), .C2(n8323), .A(n8228), .B(n8227), .ZN(n8229)
         );
  OAI21_X1 U9801 ( .B1(n8230), .B2(n8311), .A(n8229), .ZN(P2_U3159) );
  OAI21_X1 U9802 ( .B1(n8233), .B2(n8232), .A(n8231), .ZN(n8234) );
  NAND2_X1 U9803 ( .A1(n8234), .A2(n8316), .ZN(n8239) );
  AOI22_X1 U9804 ( .A1(n8781), .A2(n8303), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8235) );
  OAI21_X1 U9805 ( .B1(n8236), .B2(n8306), .A(n8235), .ZN(n8237) );
  AOI21_X1 U9806 ( .B1(n8784), .B2(n8323), .A(n8237), .ZN(n8238) );
  OAI211_X1 U9807 ( .C1(n5459), .C2(n8326), .A(n8239), .B(n8238), .ZN(P2_U3163) );
  INV_X1 U9808 ( .A(n8240), .ZN(n8277) );
  INV_X1 U9809 ( .A(n8241), .ZN(n8243) );
  NOR3_X1 U9810 ( .A1(n8277), .A2(n8243), .A3(n8242), .ZN(n8246) );
  INV_X1 U9811 ( .A(n8244), .ZN(n8245) );
  OAI21_X1 U9812 ( .B1(n8246), .B2(n8245), .A(n8316), .ZN(n8250) );
  AOI22_X1 U9813 ( .A1(n8736), .A2(n8303), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8247) );
  OAI21_X1 U9814 ( .B1(n8514), .B2(n8306), .A(n8247), .ZN(n8248) );
  AOI21_X1 U9815 ( .B1(n8739), .B2(n8323), .A(n8248), .ZN(n8249) );
  OAI211_X1 U9816 ( .C1(n4772), .C2(n8326), .A(n8250), .B(n8249), .ZN(P2_U3165) );
  INV_X1 U9817 ( .A(n8252), .ZN(n8253) );
  AOI21_X1 U9818 ( .B1(n8254), .B2(n8251), .A(n8253), .ZN(n8262) );
  INV_X1 U9819 ( .A(n8307), .ZN(n8816) );
  AOI22_X1 U9820 ( .A1(n8816), .A2(n8303), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3151), .ZN(n8257) );
  NAND2_X1 U9821 ( .A1(n8323), .A2(n8255), .ZN(n8256) );
  OAI211_X1 U9822 ( .C1(n8258), .C2(n8306), .A(n8257), .B(n8256), .ZN(n8259)
         );
  AOI21_X1 U9823 ( .B1(n8260), .B2(n8309), .A(n8259), .ZN(n8261) );
  OAI21_X1 U9824 ( .B1(n8262), .B2(n8311), .A(n8261), .ZN(P2_U3166) );
  OAI21_X1 U9825 ( .B1(n8265), .B2(n8264), .A(n8263), .ZN(n8266) );
  NAND2_X1 U9826 ( .A1(n8266), .A2(n8316), .ZN(n8272) );
  INV_X1 U9827 ( .A(n8267), .ZN(n8830) );
  AOI22_X1 U9828 ( .A1(n8303), .A2(n8827), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8268) );
  OAI21_X1 U9829 ( .B1(n8269), .B2(n8306), .A(n8268), .ZN(n8270) );
  AOI21_X1 U9830 ( .B1(n8830), .B2(n8323), .A(n8270), .ZN(n8271) );
  OAI211_X1 U9831 ( .C1(n8273), .C2(n8326), .A(n8272), .B(n8271), .ZN(P2_U3168) );
  INV_X1 U9832 ( .A(n8274), .ZN(n8276) );
  NOR3_X1 U9833 ( .A1(n4378), .A2(n8276), .A3(n8275), .ZN(n8278) );
  OAI21_X1 U9834 ( .B1(n8278), .B2(n8277), .A(n8316), .ZN(n8282) );
  AOI22_X1 U9835 ( .A1(n8745), .A2(n8303), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8279) );
  OAI21_X1 U9836 ( .B1(n8508), .B2(n8306), .A(n8279), .ZN(n8280) );
  AOI21_X1 U9837 ( .B1(n8749), .B2(n8323), .A(n8280), .ZN(n8281) );
  OAI211_X1 U9838 ( .C1(n8743), .C2(n8326), .A(n8282), .B(n8281), .ZN(P2_U3169) );
  AOI21_X1 U9839 ( .B1(n8284), .B2(n8283), .A(n4437), .ZN(n8290) );
  AOI22_X1 U9840 ( .A1(n8793), .A2(n8303), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8286) );
  NAND2_X1 U9841 ( .A1(n8323), .A2(n8796), .ZN(n8285) );
  OAI211_X1 U9842 ( .C1(n8287), .C2(n8306), .A(n8286), .B(n8285), .ZN(n8288)
         );
  AOI21_X1 U9843 ( .B1(n8937), .B2(n8309), .A(n8288), .ZN(n8289) );
  OAI21_X1 U9844 ( .B1(n8290), .B2(n8311), .A(n8289), .ZN(P2_U3173) );
  INV_X1 U9845 ( .A(n8925), .ZN(n8300) );
  INV_X1 U9846 ( .A(n8231), .ZN(n8293) );
  OAI21_X1 U9847 ( .B1(n8293), .B2(n8292), .A(n8291), .ZN(n8295) );
  NAND3_X1 U9848 ( .A1(n8295), .A2(n8316), .A3(n8294), .ZN(n8299) );
  AOI22_X1 U9849 ( .A1(n8793), .A2(n8319), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8296) );
  OAI21_X1 U9850 ( .B1(n8508), .B2(n8321), .A(n8296), .ZN(n8297) );
  AOI21_X1 U9851 ( .B1(n8770), .B2(n8323), .A(n8297), .ZN(n8298) );
  OAI211_X1 U9852 ( .C1(n8300), .C2(n8326), .A(n8299), .B(n8298), .ZN(P2_U3175) );
  XOR2_X1 U9853 ( .A(n8302), .B(n8301), .Z(n8312) );
  AOI22_X1 U9854 ( .A1(n8303), .A2(n8817), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8305) );
  NAND2_X1 U9855 ( .A1(n8323), .A2(n8820), .ZN(n8304) );
  OAI211_X1 U9856 ( .C1(n8307), .C2(n8306), .A(n8305), .B(n8304), .ZN(n8308)
         );
  AOI21_X1 U9857 ( .B1(n8944), .B2(n8309), .A(n8308), .ZN(n8310) );
  OAI21_X1 U9858 ( .B1(n8312), .B2(n8311), .A(n8310), .ZN(P2_U3178) );
  OAI21_X1 U9859 ( .B1(n8315), .B2(n8314), .A(n8313), .ZN(n8317) );
  NAND2_X1 U9860 ( .A1(n8317), .A2(n8316), .ZN(n8325) );
  AOI22_X1 U9861 ( .A1(n8745), .A2(n8319), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8320) );
  OAI21_X1 U9862 ( .B1(n8702), .B2(n8321), .A(n8320), .ZN(n8322) );
  AOI21_X1 U9863 ( .B1(n8729), .B2(n8323), .A(n8322), .ZN(n8324) );
  OAI211_X1 U9864 ( .C1(n8327), .C2(n8326), .A(n8325), .B(n8324), .ZN(P2_U3180) );
  NAND2_X1 U9865 ( .A1(n8697), .A2(n8576), .ZN(n8349) );
  NOR2_X1 U9866 ( .A1(n8331), .A2(n6440), .ZN(n8328) );
  NAND2_X1 U9867 ( .A1(n8330), .A2(n8329), .ZN(n8333) );
  OR2_X1 U9868 ( .A1(n8331), .A2(n8127), .ZN(n8332) );
  AOI22_X1 U9869 ( .A1(n8334), .A2(n8349), .B1(n8687), .B2(n8883), .ZN(n8346)
         );
  INV_X1 U9870 ( .A(n8687), .ZN(n8879) );
  INV_X1 U9871 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U9872 ( .A1(n5214), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8338) );
  INV_X1 U9873 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8335) );
  OR2_X1 U9874 ( .A1(n8336), .A2(n8335), .ZN(n8337) );
  OAI211_X1 U9875 ( .C1(n5429), .C2(n8339), .A(n8338), .B(n8337), .ZN(n8340)
         );
  INV_X1 U9876 ( .A(n8340), .ZN(n8341) );
  NAND2_X1 U9877 ( .A1(n8342), .A2(n8341), .ZN(n8684) );
  INV_X1 U9878 ( .A(n8684), .ZN(n8348) );
  OR2_X1 U9879 ( .A1(n8879), .A2(n8348), .ZN(n8558) );
  INV_X1 U9880 ( .A(n8575), .ZN(n8344) );
  NAND2_X1 U9881 ( .A1(n8883), .A2(n8344), .ZN(n8547) );
  OR2_X1 U9882 ( .A1(n8697), .A2(n8576), .ZN(n8343) );
  AND2_X1 U9883 ( .A1(n8547), .A2(n8343), .ZN(n8543) );
  OR2_X1 U9884 ( .A1(n8883), .A2(n8344), .ZN(n8546) );
  AOI21_X1 U9885 ( .B1(n8684), .B2(n8546), .A(n8687), .ZN(n8345) );
  AOI21_X1 U9886 ( .B1(n8346), .B2(n8347), .A(n8345), .ZN(n8377) );
  AND2_X1 U9887 ( .A1(n8879), .A2(n8348), .ZN(n8563) );
  NAND2_X1 U9888 ( .A1(n8546), .A2(n8349), .ZN(n8552) );
  INV_X1 U9889 ( .A(n8505), .ZN(n8350) );
  OR2_X1 U9890 ( .A1(n8492), .A2(n8350), .ZN(n8750) );
  INV_X1 U9891 ( .A(n8506), .ZN(n8351) );
  NOR2_X1 U9892 ( .A1(n8491), .A2(n8351), .ZN(n8755) );
  INV_X1 U9893 ( .A(n8777), .ZN(n8775) );
  INV_X1 U9894 ( .A(n8352), .ZN(n8791) );
  INV_X1 U9895 ( .A(n8803), .ZN(n8371) );
  INV_X1 U9896 ( .A(n8479), .ZN(n8353) );
  NOR4_X1 U9897 ( .A1(n8356), .A2(n8355), .A3(n6878), .A4(n8354), .ZN(n8359)
         );
  NAND4_X1 U9898 ( .A1(n8359), .A2(n8358), .A3(n8357), .A4(n9840), .ZN(n8362)
         );
  NOR4_X1 U9899 ( .A1(n8362), .A2(n8361), .A3(n8360), .A4(n8416), .ZN(n8364)
         );
  NAND4_X1 U9900 ( .A1(n8364), .A2(n8445), .A3(n8363), .A4(n4719), .ZN(n8365)
         );
  NOR4_X1 U9901 ( .A1(n8368), .A2(n8367), .A3(n8366), .A4(n8365), .ZN(n8369)
         );
  NAND3_X1 U9902 ( .A1(n8824), .A2(n8369), .A3(n8463), .ZN(n8370) );
  NOR4_X1 U9903 ( .A1(n8791), .A2(n8371), .A3(n8814), .A4(n8370), .ZN(n8372)
         );
  NAND4_X1 U9904 ( .A1(n8755), .A2(n8775), .A3(n8372), .A4(n4727), .ZN(n8373)
         );
  NOR4_X1 U9905 ( .A1(n8725), .A2(n8734), .A3(n8750), .A4(n8373), .ZN(n8374)
         );
  INV_X1 U9906 ( .A(n8713), .ZN(n8715) );
  AOI21_X1 U9907 ( .B1(n8377), .B2(n8381), .A(n8376), .ZN(n8378) );
  XNOR2_X1 U9908 ( .A(n8378), .B(n8663), .ZN(n8567) );
  INV_X1 U9909 ( .A(n8560), .ZN(n8561) );
  MUX2_X1 U9910 ( .A(n8704), .B(n8545), .S(n8697), .Z(n8380) );
  OR2_X1 U9911 ( .A1(n8576), .A2(n8554), .ZN(n8379) );
  NAND2_X1 U9912 ( .A1(n8380), .A2(n8379), .ZN(n8537) );
  NAND2_X1 U9913 ( .A1(n8382), .A2(n8381), .ZN(n8389) );
  NAND3_X1 U9914 ( .A1(n8389), .A2(n6571), .A3(n8384), .ZN(n8383) );
  NAND2_X1 U9915 ( .A1(n8383), .A2(n8387), .ZN(n8386) );
  INV_X1 U9916 ( .A(n8384), .ZN(n8385) );
  NAND2_X1 U9917 ( .A1(n8387), .A2(n8572), .ZN(n8388) );
  OAI21_X1 U9918 ( .B1(n8389), .B2(n8388), .A(n9859), .ZN(n8395) );
  NAND2_X1 U9919 ( .A1(n8390), .A2(n8399), .ZN(n8394) );
  NAND2_X1 U9920 ( .A1(n9854), .A2(n8391), .ZN(n8404) );
  NAND2_X1 U9921 ( .A1(n8392), .A2(n8404), .ZN(n8393) );
  NAND2_X1 U9922 ( .A1(n8398), .A2(n8397), .ZN(n8407) );
  INV_X1 U9923 ( .A(n8399), .ZN(n8401) );
  OAI211_X1 U9924 ( .C1(n8407), .C2(n8401), .A(n8408), .B(n8400), .ZN(n8402)
         );
  NAND2_X1 U9925 ( .A1(n8402), .A2(n8411), .ZN(n8403) );
  NAND2_X1 U9926 ( .A1(n8403), .A2(n8410), .ZN(n8414) );
  INV_X1 U9927 ( .A(n8404), .ZN(n8406) );
  OAI21_X1 U9928 ( .B1(n8407), .B2(n8406), .A(n8405), .ZN(n8409) );
  NAND2_X1 U9929 ( .A1(n8409), .A2(n8408), .ZN(n8412) );
  AOI21_X1 U9930 ( .B1(n8412), .B2(n8411), .A(n4636), .ZN(n8413) );
  NAND2_X1 U9931 ( .A1(n8426), .A2(n8425), .ZN(n8421) );
  NAND2_X1 U9932 ( .A1(n8419), .A2(n8418), .ZN(n8420) );
  MUX2_X1 U9933 ( .A(n8421), .B(n8420), .S(n8554), .Z(n8422) );
  INV_X1 U9934 ( .A(n8422), .ZN(n8429) );
  NAND2_X1 U9935 ( .A1(n8423), .A2(n8429), .ZN(n8433) );
  NAND2_X1 U9936 ( .A1(n8425), .A2(n8424), .ZN(n8428) );
  NAND2_X1 U9937 ( .A1(n8434), .A2(n8426), .ZN(n8427) );
  AOI21_X1 U9938 ( .B1(n8429), .B2(n8428), .A(n8427), .ZN(n8431) );
  MUX2_X1 U9939 ( .A(n8431), .B(n8430), .S(n8545), .Z(n8432) );
  NAND2_X1 U9940 ( .A1(n8433), .A2(n8432), .ZN(n8442) );
  INV_X1 U9941 ( .A(n8434), .ZN(n8435) );
  NOR2_X1 U9942 ( .A1(n8440), .A2(n8435), .ZN(n8437) );
  AOI21_X1 U9943 ( .B1(n8442), .B2(n8437), .A(n8436), .ZN(n8444) );
  AND2_X1 U9944 ( .A1(n8439), .A2(n8438), .ZN(n8441) );
  AOI21_X1 U9945 ( .B1(n8442), .B2(n8441), .A(n8440), .ZN(n8443) );
  NAND2_X1 U9946 ( .A1(n8446), .A2(n8445), .ZN(n8450) );
  MUX2_X1 U9947 ( .A(n8448), .B(n8447), .S(n8554), .Z(n8449) );
  NAND2_X1 U9948 ( .A1(n8450), .A2(n8449), .ZN(n8455) );
  INV_X1 U9949 ( .A(n8455), .ZN(n8458) );
  MUX2_X1 U9950 ( .A(n8579), .B(n8451), .S(n8554), .Z(n8452) );
  INV_X1 U9951 ( .A(n8452), .ZN(n8453) );
  OAI21_X1 U9952 ( .B1(n8455), .B2(n8454), .A(n8453), .ZN(n8456) );
  MUX2_X1 U9953 ( .A(n8461), .B(n8460), .S(n8554), .Z(n8462) );
  NAND3_X1 U9954 ( .A1(n8464), .A2(n8463), .A3(n8462), .ZN(n8469) );
  MUX2_X1 U9955 ( .A(n8466), .B(n8465), .S(n8554), .Z(n8467) );
  NAND3_X1 U9956 ( .A1(n8469), .A2(n8468), .A3(n8467), .ZN(n8474) );
  MUX2_X1 U9957 ( .A(n8471), .B(n8470), .S(n8545), .Z(n8472) );
  AND2_X1 U9958 ( .A1(n8824), .A2(n8472), .ZN(n8473) );
  NAND2_X1 U9959 ( .A1(n8474), .A2(n8473), .ZN(n8478) );
  NAND3_X1 U9960 ( .A1(n8478), .A2(n8479), .A3(n8475), .ZN(n8477) );
  NAND3_X1 U9961 ( .A1(n8477), .A2(n8483), .A3(n5583), .ZN(n8482) );
  NAND3_X1 U9962 ( .A1(n8478), .A2(n5583), .A3(n8811), .ZN(n8480) );
  NAND2_X1 U9963 ( .A1(n8480), .A2(n8479), .ZN(n8481) );
  NAND2_X1 U9964 ( .A1(n8498), .A2(n8483), .ZN(n8487) );
  NOR2_X1 U9965 ( .A1(n8485), .A2(n4641), .ZN(n8497) );
  INV_X1 U9966 ( .A(n8499), .ZN(n8486) );
  AOI21_X1 U9967 ( .B1(n8487), .B2(n8497), .A(n8486), .ZN(n8489) );
  OAI21_X1 U9968 ( .B1(n8489), .B2(n8488), .A(n4727), .ZN(n8495) );
  NAND2_X1 U9969 ( .A1(n8925), .A2(n8490), .ZN(n8494) );
  OR3_X1 U9970 ( .A1(n8492), .A2(n8554), .A3(n8491), .ZN(n8493) );
  AOI21_X1 U9971 ( .B1(n8495), .B2(n8494), .A(n8493), .ZN(n8522) );
  NAND2_X1 U9972 ( .A1(n8767), .A2(n8554), .ZN(n8513) );
  INV_X1 U9973 ( .A(n8513), .ZN(n8496) );
  AOI22_X1 U9974 ( .A1(n8512), .A2(n8496), .B1(n8554), .B2(n8757), .ZN(n8520)
         );
  NAND2_X1 U9975 ( .A1(n8498), .A2(n8497), .ZN(n8500) );
  NAND2_X1 U9976 ( .A1(n8500), .A2(n8499), .ZN(n8502) );
  NAND3_X1 U9977 ( .A1(n8502), .A2(n4727), .A3(n8501), .ZN(n8504) );
  NAND2_X1 U9978 ( .A1(n8504), .A2(n8503), .ZN(n8507) );
  NAND4_X1 U9979 ( .A1(n8507), .A2(n8554), .A3(n8506), .A4(n8505), .ZN(n8519)
         );
  NAND2_X1 U9980 ( .A1(n8508), .A2(n8545), .ZN(n8509) );
  OAI22_X1 U9981 ( .A1(n8512), .A2(n8509), .B1(n8554), .B2(n8757), .ZN(n8517)
         );
  INV_X1 U9982 ( .A(n8509), .ZN(n8510) );
  AND2_X1 U9983 ( .A1(n8514), .A2(n8510), .ZN(n8511) );
  OR2_X1 U9984 ( .A1(n8512), .A2(n8511), .ZN(n8516) );
  OAI21_X1 U9985 ( .B1(n8514), .B2(n8513), .A(n8512), .ZN(n8515) );
  AOI22_X1 U9986 ( .A1(n8913), .A2(n8517), .B1(n8516), .B2(n8515), .ZN(n8518)
         );
  INV_X1 U9987 ( .A(n8734), .ZN(n8521) );
  MUX2_X1 U9988 ( .A(n8524), .B(n8523), .S(n8554), .Z(n8525) );
  NAND2_X1 U9989 ( .A1(n8526), .A2(n8525), .ZN(n8527) );
  NAND2_X1 U9990 ( .A1(n8527), .A2(n8723), .ZN(n8535) );
  MUX2_X1 U9991 ( .A(n4396), .B(n8528), .S(n8554), .Z(n8529) );
  NOR2_X1 U9992 ( .A1(n8713), .A2(n8529), .ZN(n8534) );
  MUX2_X1 U9993 ( .A(n8531), .B(n8530), .S(n8545), .Z(n8532) );
  INV_X1 U9994 ( .A(n8532), .ZN(n8533) );
  AOI21_X1 U9995 ( .B1(n8535), .B2(n8534), .A(n8533), .ZN(n8536) );
  NAND2_X1 U9996 ( .A1(n8537), .A2(n8536), .ZN(n8542) );
  MUX2_X1 U9997 ( .A(n8717), .B(n8709), .S(n8545), .Z(n8540) );
  NAND2_X1 U9998 ( .A1(n8537), .A2(n8540), .ZN(n8538) );
  NAND2_X1 U9999 ( .A1(n8542), .A2(n8538), .ZN(n8551) );
  NAND2_X1 U10000 ( .A1(n8551), .A2(n8539), .ZN(n8544) );
  INV_X1 U10001 ( .A(n8540), .ZN(n8541) );
  NAND3_X1 U10002 ( .A1(n8544), .A2(n8543), .A3(n8553), .ZN(n8550) );
  NAND2_X1 U10003 ( .A1(n8546), .A2(n8545), .ZN(n8548) );
  NAND2_X1 U10004 ( .A1(n8548), .A2(n8547), .ZN(n8549) );
  NAND2_X1 U10005 ( .A1(n8550), .A2(n8549), .ZN(n8559) );
  NAND2_X1 U10006 ( .A1(n8551), .A2(n8892), .ZN(n8556) );
  INV_X1 U10007 ( .A(n8552), .ZN(n8555) );
  NAND3_X1 U10008 ( .A1(n8559), .A2(n8558), .A3(n8557), .ZN(n8564) );
  INV_X1 U10009 ( .A(n8562), .ZN(n9864) );
  NAND3_X1 U10010 ( .A1(n8564), .A2(n9864), .A3(n4674), .ZN(n8565) );
  NAND3_X1 U10011 ( .A1(n8569), .A2(n8568), .A3(n8631), .ZN(n8570) );
  OAI211_X1 U10012 ( .C1(n8572), .C2(n8571), .A(n8570), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8573) );
  NAND2_X1 U10013 ( .A1(n8574), .A2(n8573), .ZN(P2_U3296) );
  MUX2_X1 U10014 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8684), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10015 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8575), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10016 ( .A(P2_U3893), .ZN(n8637) );
  MUX2_X1 U10017 ( .A(n8576), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8637), .Z(
        P2_U3520) );
  MUX2_X1 U10018 ( .A(n8717), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8637), .Z(
        P2_U3519) );
  MUX2_X1 U10019 ( .A(n8168), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8637), .Z(
        P2_U3518) );
  MUX2_X1 U10020 ( .A(n8736), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8637), .Z(
        P2_U3517) );
  MUX2_X1 U10021 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8745), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10022 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8757), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10023 ( .A(n8767), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8637), .Z(
        P2_U3514) );
  MUX2_X1 U10024 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8781), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10025 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8793), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10026 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8800), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10027 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8817), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10028 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8827), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8816), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10030 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8826), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10031 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8577), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8578), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10033 ( .A(n8579), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8637), .Z(
        P2_U3504) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8580), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10035 ( .A(n8581), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8637), .Z(
        P2_U3502) );
  MUX2_X1 U10036 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8582), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8583), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10038 ( .A(n8584), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8637), .Z(
        P2_U3499) );
  MUX2_X1 U10039 ( .A(n8585), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8637), .Z(
        P2_U3498) );
  MUX2_X1 U10040 ( .A(n8586), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8637), .Z(
        P2_U3497) );
  MUX2_X1 U10041 ( .A(n8587), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8637), .Z(
        P2_U3496) );
  MUX2_X1 U10042 ( .A(n9838), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8637), .Z(
        P2_U3495) );
  MUX2_X1 U10043 ( .A(n9854), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8637), .Z(
        P2_U3494) );
  MUX2_X1 U10044 ( .A(n9837), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8637), .Z(
        P2_U3493) );
  MUX2_X1 U10045 ( .A(n6675), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8637), .Z(
        P2_U3492) );
  MUX2_X1 U10046 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n5198), .S(P2_U3893), .Z(
        P2_U3491) );
  AOI22_X1 U10047 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8608), .B1(n9800), .B2(
        n8589), .ZN(n9791) );
  NOR2_X1 U10048 ( .A1(n9792), .A2(n9791), .ZN(n9790) );
  AOI21_X1 U10049 ( .B1(n8591), .B2(n8590), .A(n8643), .ZN(n8615) );
  MUX2_X1 U10050 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8631), .Z(n8626) );
  XNOR2_X1 U10051 ( .A(n8626), .B(n8642), .ZN(n8599) );
  MUX2_X1 U10052 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8631), .Z(n8592) );
  OR2_X1 U10053 ( .A1(n8592), .A2(n9800), .ZN(n8597) );
  XNOR2_X1 U10054 ( .A(n8592), .B(n8608), .ZN(n9788) );
  INV_X1 U10055 ( .A(n8593), .ZN(n8594) );
  NAND2_X1 U10056 ( .A1(n8604), .A2(n8594), .ZN(n8596) );
  NAND2_X1 U10057 ( .A1(n8596), .A2(n8595), .ZN(n9787) );
  NAND2_X1 U10058 ( .A1(n9788), .A2(n9787), .ZN(n9786) );
  NAND2_X1 U10059 ( .A1(n8597), .A2(n9786), .ZN(n8598) );
  NAND2_X1 U10060 ( .A1(n8599), .A2(n8598), .ZN(n8627) );
  OAI21_X1 U10061 ( .B1(n8599), .B2(n8598), .A(n8627), .ZN(n8613) );
  INV_X1 U10062 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U10063 ( .A1(n8600), .A2(n8642), .ZN(n8602) );
  OAI211_X1 U10064 ( .C1(n9994), .C2(n9783), .A(n8602), .B(n8601), .ZN(n8612)
         );
  NOR2_X1 U10065 ( .A1(n8604), .A2(n8603), .ZN(n8606) );
  AOI22_X1 U10066 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8608), .B1(n9800), .B2(
        n8607), .ZN(n9784) );
  NOR2_X1 U10067 ( .A1(n7706), .A2(n8609), .ZN(n8617) );
  AOI21_X1 U10068 ( .B1(n7706), .B2(n8609), .A(n8617), .ZN(n8610) );
  NOR2_X1 U10069 ( .A1(n8610), .A2(n9829), .ZN(n8611) );
  AOI211_X1 U10070 ( .C1(n9832), .C2(n8613), .A(n8612), .B(n8611), .ZN(n8614)
         );
  OAI21_X1 U10071 ( .B1(n8615), .B2(n9825), .A(n8614), .ZN(P2_U3197) );
  NOR2_X1 U10072 ( .A1(n8642), .A2(n8616), .ZN(n8618) );
  NOR2_X1 U10073 ( .A1(n8618), .A2(n8617), .ZN(n9803) );
  AOI22_X1 U10074 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8646), .B1(n9817), .B2(
        n7738), .ZN(n9802) );
  NOR2_X1 U10075 ( .A1(n8648), .A2(n8619), .ZN(n8620) );
  NOR2_X1 U10076 ( .A1(n8620), .A2(n9827), .ZN(n8622) );
  NAND2_X1 U10077 ( .A1(n8650), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8659) );
  OAI21_X1 U10078 ( .B1(n8650), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8659), .ZN(
        n8621) );
  NOR2_X1 U10079 ( .A1(n8622), .A2(n8621), .ZN(n8661) );
  AOI21_X1 U10080 ( .B1(n8622), .B2(n8621), .A(n8661), .ZN(n8658) );
  MUX2_X1 U10081 ( .A(n8829), .B(n9824), .S(n8631), .Z(n8623) );
  NAND2_X1 U10082 ( .A1(n8623), .A2(n8648), .ZN(n8630) );
  XNOR2_X1 U10083 ( .A(n8623), .B(n9834), .ZN(n9821) );
  MUX2_X1 U10084 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8631), .Z(n8624) );
  OR2_X1 U10085 ( .A1(n8624), .A2(n9817), .ZN(n8629) );
  XNOR2_X1 U10086 ( .A(n8624), .B(n8646), .ZN(n9806) );
  OR2_X1 U10087 ( .A1(n8626), .A2(n8625), .ZN(n8628) );
  NAND2_X1 U10088 ( .A1(n8628), .A2(n8627), .ZN(n9805) );
  NAND2_X1 U10089 ( .A1(n9806), .A2(n9805), .ZN(n9804) );
  NAND2_X1 U10090 ( .A1(n8629), .A2(n9804), .ZN(n9820) );
  NAND2_X1 U10091 ( .A1(n9821), .A2(n9820), .ZN(n9819) );
  NAND2_X1 U10092 ( .A1(n8630), .A2(n9819), .ZN(n8632) );
  MUX2_X1 U10093 ( .A(n8819), .B(n8871), .S(n8631), .Z(n8633) );
  AND2_X1 U10094 ( .A1(n8632), .A2(n8633), .ZN(n8666) );
  INV_X1 U10095 ( .A(n8666), .ZN(n8636) );
  INV_X1 U10096 ( .A(n8632), .ZN(n8635) );
  INV_X1 U10097 ( .A(n8633), .ZN(n8634) );
  NAND2_X1 U10098 ( .A1(n8635), .A2(n8634), .ZN(n8667) );
  NAND2_X1 U10099 ( .A1(n8636), .A2(n8667), .ZN(n8638) );
  OAI21_X1 U10100 ( .B1(n8638), .B2(n8637), .A(n9835), .ZN(n8656) );
  INV_X1 U10101 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10021) );
  NAND3_X1 U10102 ( .A1(n8638), .A2(n9832), .A3(n8650), .ZN(n8640) );
  INV_X1 U10103 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10027) );
  OR2_X1 U10104 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10027), .ZN(n8639) );
  OAI211_X1 U10105 ( .C1(n10021), .C2(n9783), .A(n8640), .B(n8639), .ZN(n8655)
         );
  NOR2_X1 U10106 ( .A1(n8642), .A2(n8641), .ZN(n8644) );
  AOI22_X1 U10107 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8646), .B1(n9817), .B2(
        n8645), .ZN(n9809) );
  NOR2_X1 U10108 ( .A1(n8648), .A2(n8647), .ZN(n8649) );
  NAND2_X1 U10109 ( .A1(n8650), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8674) );
  OAI21_X1 U10110 ( .B1(n8650), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8674), .ZN(
        n8651) );
  AOI21_X1 U10111 ( .B1(n8652), .B2(n8651), .A(n8676), .ZN(n8653) );
  NOR2_X1 U10112 ( .A1(n8653), .A2(n9825), .ZN(n8654) );
  OAI21_X1 U10113 ( .B1(n8658), .B2(n9829), .A(n8657), .ZN(P2_U3200) );
  INV_X1 U10114 ( .A(n8659), .ZN(n8660) );
  NOR2_X1 U10115 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  MUX2_X1 U10116 ( .A(n5145), .B(P2_REG2_REG_19__SCAN_IN), .S(n8663), .Z(n8665) );
  XNOR2_X1 U10117 ( .A(n8662), .B(n8665), .ZN(n8682) );
  XNOR2_X1 U10118 ( .A(n8663), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8677) );
  MUX2_X1 U10119 ( .A(n8677), .B(n8665), .S(n8664), .Z(n8670) );
  AOI21_X1 U10120 ( .B1(n8668), .B2(n8667), .A(n8666), .ZN(n8669) );
  XOR2_X1 U10121 ( .A(n8670), .B(n8669), .Z(n8681) );
  NAND2_X1 U10122 ( .A1(n9818), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8672) );
  OAI211_X1 U10123 ( .C1(n9835), .C2(n8673), .A(n8672), .B(n8671), .ZN(n8680)
         );
  INV_X1 U10124 ( .A(n8674), .ZN(n8675) );
  XNOR2_X1 U10125 ( .A(n8678), .B(n8677), .ZN(n8679) );
  OAI21_X1 U10126 ( .B1(n9829), .B2(n8682), .A(n4427), .ZN(P2_U3201) );
  NOR2_X1 U10127 ( .A1(n8685), .A2(n9862), .ZN(n8694) );
  AOI21_X1 U10128 ( .B1(n8880), .B2(n9868), .A(n8694), .ZN(n8689) );
  NAND2_X1 U10129 ( .A1(n9871), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8686) );
  OAI211_X1 U10130 ( .C1(n8687), .C2(n8807), .A(n8689), .B(n8686), .ZN(
        P2_U3202) );
  INV_X1 U10131 ( .A(n8883), .ZN(n8690) );
  NAND2_X1 U10132 ( .A1(n9871), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8688) );
  OAI211_X1 U10133 ( .C1(n8690), .C2(n8807), .A(n8689), .B(n8688), .ZN(
        P2_U3203) );
  NAND2_X1 U10134 ( .A1(n8693), .A2(n9868), .ZN(n8696) );
  AOI21_X1 U10135 ( .B1(n9871), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8694), .ZN(
        n8695) );
  OAI211_X1 U10136 ( .C1(n8697), .C2(n8807), .A(n8696), .B(n8695), .ZN(
        P2_U3204) );
  XOR2_X1 U10137 ( .A(n8700), .B(n8698), .Z(n8888) );
  INV_X1 U10138 ( .A(n8888), .ZN(n8712) );
  INV_X1 U10139 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8707) );
  XOR2_X1 U10140 ( .A(n8700), .B(n8699), .Z(n8706) );
  OAI22_X1 U10141 ( .A1(n8704), .A2(n8703), .B1(n8702), .B2(n8701), .ZN(n8705)
         );
  AOI21_X1 U10142 ( .B1(n8706), .B2(n9851), .A(n8705), .ZN(n8886) );
  MUX2_X1 U10143 ( .A(n8707), .B(n8886), .S(n9868), .Z(n8711) );
  AOI22_X1 U10144 ( .A1(n8709), .A2(n9842), .B1(n9843), .B2(n8708), .ZN(n8710)
         );
  OAI211_X1 U10145 ( .C1(n8712), .C2(n8833), .A(n8711), .B(n8710), .ZN(
        P2_U3205) );
  XNOR2_X1 U10146 ( .A(n8714), .B(n8713), .ZN(n8898) );
  INV_X1 U10147 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8719) );
  XNOR2_X1 U10148 ( .A(n8716), .B(n8715), .ZN(n8718) );
  MUX2_X1 U10149 ( .A(n8719), .B(n8893), .S(n9868), .Z(n8722) );
  AOI22_X1 U10150 ( .A1(n8895), .A2(n9842), .B1(n9843), .B2(n8720), .ZN(n8721)
         );
  OAI211_X1 U10151 ( .C1(n8898), .C2(n8833), .A(n8722), .B(n8721), .ZN(
        P2_U3206) );
  XNOR2_X1 U10152 ( .A(n8724), .B(n8723), .ZN(n8904) );
  INV_X1 U10153 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8728) );
  XNOR2_X1 U10154 ( .A(n8726), .B(n8725), .ZN(n8727) );
  AOI222_X1 U10155 ( .A1(n9851), .A2(n8727), .B1(n8745), .B2(n9855), .C1(n8168), .C2(n9853), .ZN(n8899) );
  MUX2_X1 U10156 ( .A(n8728), .B(n8899), .S(n9868), .Z(n8731) );
  AOI22_X1 U10157 ( .A1(n8901), .A2(n9842), .B1(n9843), .B2(n8729), .ZN(n8730)
         );
  OAI211_X1 U10158 ( .C1(n8904), .C2(n8833), .A(n8731), .B(n8730), .ZN(
        P2_U3207) );
  XNOR2_X1 U10159 ( .A(n8732), .B(n8734), .ZN(n8910) );
  OAI21_X1 U10160 ( .B1(n8735), .B2(n8734), .A(n8733), .ZN(n8737) );
  AOI222_X1 U10161 ( .A1(n9851), .A2(n8737), .B1(n8736), .B2(n9853), .C1(n8757), .C2(n9855), .ZN(n8905) );
  OAI21_X1 U10162 ( .B1(n4772), .B2(n8742), .A(n8905), .ZN(n8738) );
  NAND2_X1 U10163 ( .A1(n8738), .A2(n9868), .ZN(n8741) );
  AOI22_X1 U10164 ( .A1(n8739), .A2(n9843), .B1(n9871), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8740) );
  OAI211_X1 U10165 ( .C1(n8910), .C2(n8833), .A(n8741), .B(n8740), .ZN(
        P2_U3208) );
  NOR2_X1 U10166 ( .A1(n8743), .A2(n8742), .ZN(n8748) );
  XNOR2_X1 U10167 ( .A(n8744), .B(n8750), .ZN(n8746) );
  AOI222_X1 U10168 ( .A1(n9851), .A2(n8746), .B1(n8745), .B2(n9853), .C1(n8767), .C2(n9855), .ZN(n8911) );
  INV_X1 U10169 ( .A(n8911), .ZN(n8747) );
  AOI211_X1 U10170 ( .C1(n9843), .C2(n8749), .A(n8748), .B(n8747), .ZN(n8753)
         );
  XNOR2_X1 U10171 ( .A(n8751), .B(n8750), .ZN(n8914) );
  AOI22_X1 U10172 ( .A1(n8914), .A2(n9845), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9871), .ZN(n8752) );
  OAI21_X1 U10173 ( .B1(n8753), .B2(n9871), .A(n8752), .ZN(P2_U3209) );
  XNOR2_X1 U10174 ( .A(n8754), .B(n8755), .ZN(n8922) );
  INV_X1 U10175 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8759) );
  XOR2_X1 U10176 ( .A(n8756), .B(n8755), .Z(n8758) );
  AOI222_X1 U10177 ( .A1(n9851), .A2(n8758), .B1(n8757), .B2(n9853), .C1(n8781), .C2(n9855), .ZN(n8917) );
  MUX2_X1 U10178 ( .A(n8759), .B(n8917), .S(n9868), .Z(n8762) );
  AOI22_X1 U10179 ( .A1(n8919), .A2(n9842), .B1(n9843), .B2(n8760), .ZN(n8761)
         );
  OAI211_X1 U10180 ( .C1(n8922), .C2(n8833), .A(n8762), .B(n8761), .ZN(
        P2_U3210) );
  XNOR2_X1 U10181 ( .A(n8763), .B(n4727), .ZN(n8928) );
  INV_X1 U10182 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8769) );
  OAI21_X1 U10183 ( .B1(n8766), .B2(n8765), .A(n8764), .ZN(n8768) );
  AOI222_X1 U10184 ( .A1(n9851), .A2(n8768), .B1(n8793), .B2(n9855), .C1(n8767), .C2(n9853), .ZN(n8923) );
  MUX2_X1 U10185 ( .A(n8769), .B(n8923), .S(n9868), .Z(n8772) );
  AOI22_X1 U10186 ( .A1(n8925), .A2(n9842), .B1(n9843), .B2(n8770), .ZN(n8771)
         );
  OAI211_X1 U10187 ( .C1(n8928), .C2(n8833), .A(n8772), .B(n8771), .ZN(
        P2_U3211) );
  NAND2_X1 U10188 ( .A1(n8774), .A2(n8773), .ZN(n8776) );
  XNOR2_X1 U10189 ( .A(n8776), .B(n8775), .ZN(n8934) );
  INV_X1 U10190 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8783) );
  OR3_X1 U10191 ( .A1(n8789), .A2(n8778), .A3(n8777), .ZN(n8779) );
  NAND2_X1 U10192 ( .A1(n8780), .A2(n8779), .ZN(n8782) );
  AOI222_X1 U10193 ( .A1(n9851), .A2(n8782), .B1(n8781), .B2(n9853), .C1(n8800), .C2(n9855), .ZN(n8929) );
  MUX2_X1 U10194 ( .A(n8783), .B(n8929), .S(n9868), .Z(n8786) );
  AOI22_X1 U10195 ( .A1(n8931), .A2(n9842), .B1(n9843), .B2(n8784), .ZN(n8785)
         );
  OAI211_X1 U10196 ( .C1(n8934), .C2(n8833), .A(n8786), .B(n8785), .ZN(
        P2_U3212) );
  XNOR2_X1 U10197 ( .A(n8787), .B(n8791), .ZN(n8940) );
  INV_X1 U10198 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8795) );
  INV_X1 U10199 ( .A(n8788), .ZN(n8792) );
  INV_X1 U10200 ( .A(n8789), .ZN(n8790) );
  OAI21_X1 U10201 ( .B1(n8792), .B2(n8791), .A(n8790), .ZN(n8794) );
  AOI222_X1 U10202 ( .A1(n9851), .A2(n8794), .B1(n8793), .B2(n9853), .C1(n8817), .C2(n9855), .ZN(n8935) );
  MUX2_X1 U10203 ( .A(n8795), .B(n8935), .S(n9868), .Z(n8798) );
  AOI22_X1 U10204 ( .A1(n8937), .A2(n9842), .B1(n9843), .B2(n8796), .ZN(n8797)
         );
  OAI211_X1 U10205 ( .C1(n8940), .C2(n8833), .A(n8798), .B(n8797), .ZN(
        P2_U3213) );
  XNOR2_X1 U10206 ( .A(n8799), .B(n8803), .ZN(n8801) );
  AOI222_X1 U10207 ( .A1(n9851), .A2(n8801), .B1(n8800), .B2(n9853), .C1(n8827), .C2(n9855), .ZN(n8870) );
  OAI21_X1 U10208 ( .B1(n8804), .B2(n8803), .A(n8802), .ZN(n8868) );
  AOI22_X1 U10209 ( .A1(n9871), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9843), .B2(
        n8805), .ZN(n8806) );
  OAI21_X1 U10210 ( .B1(n8808), .B2(n8807), .A(n8806), .ZN(n8809) );
  AOI21_X1 U10211 ( .B1(n8868), .B2(n9845), .A(n8809), .ZN(n8810) );
  OAI21_X1 U10212 ( .B1(n8870), .B2(n9871), .A(n8810), .ZN(P2_U3214) );
  NAND2_X1 U10213 ( .A1(n8812), .A2(n8811), .ZN(n8813) );
  XOR2_X1 U10214 ( .A(n8814), .B(n8813), .Z(n8948) );
  XOR2_X1 U10215 ( .A(n8815), .B(n8814), .Z(n8818) );
  AOI222_X1 U10216 ( .A1(n9851), .A2(n8818), .B1(n8817), .B2(n9853), .C1(n8816), .C2(n9855), .ZN(n8942) );
  MUX2_X1 U10217 ( .A(n8819), .B(n8942), .S(n9868), .Z(n8822) );
  AOI22_X1 U10218 ( .A1(n8944), .A2(n9842), .B1(n9843), .B2(n8820), .ZN(n8821)
         );
  OAI211_X1 U10219 ( .C1(n8948), .C2(n8833), .A(n8822), .B(n8821), .ZN(
        P2_U3215) );
  XOR2_X1 U10220 ( .A(n8823), .B(n8824), .Z(n8954) );
  INV_X1 U10221 ( .A(n8954), .ZN(n8834) );
  XOR2_X1 U10222 ( .A(n8825), .B(n8824), .Z(n8828) );
  AOI222_X1 U10223 ( .A1(n9851), .A2(n8828), .B1(n8827), .B2(n9853), .C1(n8826), .C2(n9855), .ZN(n8949) );
  MUX2_X1 U10224 ( .A(n8829), .B(n8949), .S(n9868), .Z(n8832) );
  AOI22_X1 U10225 ( .A1(n8951), .A2(n9842), .B1(n9843), .B2(n8830), .ZN(n8831)
         );
  OAI211_X1 U10226 ( .C1(n8834), .C2(n8833), .A(n8832), .B(n8831), .ZN(
        P2_U3216) );
  NAND2_X1 U10227 ( .A1(n8879), .A2(n8875), .ZN(n8835) );
  NAND2_X1 U10228 ( .A1(n8880), .A2(n9947), .ZN(n8836) );
  OAI211_X1 U10229 ( .C1(n9947), .C2(n8339), .A(n8835), .B(n8836), .ZN(
        P2_U3490) );
  INV_X1 U10230 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U10231 ( .A1(n8883), .A2(n8875), .ZN(n8837) );
  OAI211_X1 U10232 ( .C1(n9947), .C2(n8838), .A(n8837), .B(n8836), .ZN(
        P2_U3489) );
  INV_X1 U10233 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8839) );
  MUX2_X1 U10234 ( .A(n8839), .B(n8886), .S(n9947), .Z(n8841) );
  NAND2_X1 U10235 ( .A1(n8888), .A2(n8876), .ZN(n8840) );
  OAI211_X1 U10236 ( .C1(n8892), .C2(n8842), .A(n8841), .B(n8840), .ZN(
        P2_U3487) );
  INV_X1 U10237 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8843) );
  MUX2_X1 U10238 ( .A(n8843), .B(n8893), .S(n9947), .Z(n8845) );
  NAND2_X1 U10239 ( .A1(n8895), .A2(n8875), .ZN(n8844) );
  OAI211_X1 U10240 ( .C1(n8874), .C2(n8898), .A(n8845), .B(n8844), .ZN(
        P2_U3486) );
  INV_X1 U10241 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8846) );
  MUX2_X1 U10242 ( .A(n8846), .B(n8899), .S(n9947), .Z(n8848) );
  NAND2_X1 U10243 ( .A1(n8901), .A2(n8875), .ZN(n8847) );
  OAI211_X1 U10244 ( .C1(n8904), .C2(n8874), .A(n8848), .B(n8847), .ZN(
        P2_U3485) );
  INV_X1 U10245 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8849) );
  MUX2_X1 U10246 ( .A(n8849), .B(n8905), .S(n9947), .Z(n8851) );
  NAND2_X1 U10247 ( .A1(n8907), .A2(n8875), .ZN(n8850) );
  OAI211_X1 U10248 ( .C1(n8910), .C2(n8874), .A(n8851), .B(n8850), .ZN(
        P2_U3484) );
  INV_X1 U10249 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8852) );
  MUX2_X1 U10250 ( .A(n8852), .B(n8911), .S(n9947), .Z(n8854) );
  AOI22_X1 U10251 ( .A1(n8914), .A2(n8876), .B1(n8875), .B2(n8913), .ZN(n8853)
         );
  NAND2_X1 U10252 ( .A1(n8854), .A2(n8853), .ZN(P2_U3483) );
  INV_X1 U10253 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8855) );
  MUX2_X1 U10254 ( .A(n8855), .B(n8917), .S(n9947), .Z(n8857) );
  NAND2_X1 U10255 ( .A1(n8919), .A2(n8875), .ZN(n8856) );
  OAI211_X1 U10256 ( .C1(n8922), .C2(n8874), .A(n8857), .B(n8856), .ZN(
        P2_U3482) );
  INV_X1 U10257 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8858) );
  MUX2_X1 U10258 ( .A(n8858), .B(n8923), .S(n9947), .Z(n8860) );
  NAND2_X1 U10259 ( .A1(n8925), .A2(n8875), .ZN(n8859) );
  OAI211_X1 U10260 ( .C1(n8928), .C2(n8874), .A(n8860), .B(n8859), .ZN(
        P2_U3481) );
  INV_X1 U10261 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8861) );
  MUX2_X1 U10262 ( .A(n8861), .B(n8929), .S(n9947), .Z(n8863) );
  NAND2_X1 U10263 ( .A1(n8931), .A2(n8875), .ZN(n8862) );
  OAI211_X1 U10264 ( .C1(n8934), .C2(n8874), .A(n8863), .B(n8862), .ZN(
        P2_U3480) );
  INV_X1 U10265 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8864) );
  MUX2_X1 U10266 ( .A(n8864), .B(n8935), .S(n9947), .Z(n8866) );
  NAND2_X1 U10267 ( .A1(n8937), .A2(n8875), .ZN(n8865) );
  OAI211_X1 U10268 ( .C1(n8874), .C2(n8940), .A(n8866), .B(n8865), .ZN(
        P2_U3479) );
  AOI22_X1 U10269 ( .A1(n8868), .A2(n9919), .B1(n9930), .B2(n8867), .ZN(n8869)
         );
  NAND2_X1 U10270 ( .A1(n8870), .A2(n8869), .ZN(n8941) );
  MUX2_X1 U10271 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8941), .S(n9947), .Z(
        P2_U3478) );
  MUX2_X1 U10272 ( .A(n8871), .B(n8942), .S(n9947), .Z(n8873) );
  NAND2_X1 U10273 ( .A1(n8944), .A2(n8875), .ZN(n8872) );
  OAI211_X1 U10274 ( .C1(n8948), .C2(n8874), .A(n8873), .B(n8872), .ZN(
        P2_U3477) );
  MUX2_X1 U10275 ( .A(n9824), .B(n8949), .S(n9947), .Z(n8878) );
  AOI22_X1 U10276 ( .A1(n8954), .A2(n8876), .B1(n8875), .B2(n8951), .ZN(n8877)
         );
  NAND2_X1 U10277 ( .A1(n8878), .A2(n8877), .ZN(P2_U3476) );
  INV_X1 U10278 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8882) );
  NAND2_X1 U10279 ( .A1(n8879), .A2(n8952), .ZN(n8881) );
  NAND2_X1 U10280 ( .A1(n8880), .A2(n9931), .ZN(n8884) );
  OAI211_X1 U10281 ( .C1(n8882), .C2(n9931), .A(n8881), .B(n8884), .ZN(
        P2_U3458) );
  NAND2_X1 U10282 ( .A1(n8883), .A2(n8952), .ZN(n8885) );
  OAI211_X1 U10283 ( .C1(n5602), .C2(n9931), .A(n8885), .B(n8884), .ZN(
        P2_U3457) );
  MUX2_X1 U10284 ( .A(n8887), .B(n8886), .S(n9931), .Z(n8890) );
  NAND2_X1 U10285 ( .A1(n8888), .A2(n8953), .ZN(n8889) );
  OAI211_X1 U10286 ( .C1(n8892), .C2(n8891), .A(n8890), .B(n8889), .ZN(
        P2_U3455) );
  MUX2_X1 U10287 ( .A(n8894), .B(n8893), .S(n9931), .Z(n8897) );
  NAND2_X1 U10288 ( .A1(n8895), .A2(n8952), .ZN(n8896) );
  OAI211_X1 U10289 ( .C1(n8898), .C2(n8947), .A(n8897), .B(n8896), .ZN(
        P2_U3454) );
  MUX2_X1 U10290 ( .A(n8900), .B(n8899), .S(n9931), .Z(n8903) );
  NAND2_X1 U10291 ( .A1(n8901), .A2(n8952), .ZN(n8902) );
  OAI211_X1 U10292 ( .C1(n8904), .C2(n8947), .A(n8903), .B(n8902), .ZN(
        P2_U3453) );
  MUX2_X1 U10293 ( .A(n8906), .B(n8905), .S(n9931), .Z(n8909) );
  NAND2_X1 U10294 ( .A1(n8907), .A2(n8952), .ZN(n8908) );
  OAI211_X1 U10295 ( .C1(n8910), .C2(n8947), .A(n8909), .B(n8908), .ZN(
        P2_U3452) );
  MUX2_X1 U10296 ( .A(n8912), .B(n8911), .S(n9931), .Z(n8916) );
  AOI22_X1 U10297 ( .A1(n8914), .A2(n8953), .B1(n8952), .B2(n8913), .ZN(n8915)
         );
  NAND2_X1 U10298 ( .A1(n8916), .A2(n8915), .ZN(P2_U3451) );
  MUX2_X1 U10299 ( .A(n8918), .B(n8917), .S(n9931), .Z(n8921) );
  NAND2_X1 U10300 ( .A1(n8919), .A2(n8952), .ZN(n8920) );
  OAI211_X1 U10301 ( .C1(n8922), .C2(n8947), .A(n8921), .B(n8920), .ZN(
        P2_U3450) );
  INV_X1 U10302 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8924) );
  MUX2_X1 U10303 ( .A(n8924), .B(n8923), .S(n9931), .Z(n8927) );
  NAND2_X1 U10304 ( .A1(n8925), .A2(n8952), .ZN(n8926) );
  OAI211_X1 U10305 ( .C1(n8928), .C2(n8947), .A(n8927), .B(n8926), .ZN(
        P2_U3449) );
  INV_X1 U10306 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8930) );
  MUX2_X1 U10307 ( .A(n8930), .B(n8929), .S(n9931), .Z(n8933) );
  NAND2_X1 U10308 ( .A1(n8931), .A2(n8952), .ZN(n8932) );
  OAI211_X1 U10309 ( .C1(n8934), .C2(n8947), .A(n8933), .B(n8932), .ZN(
        P2_U3448) );
  INV_X1 U10310 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8936) );
  MUX2_X1 U10311 ( .A(n8936), .B(n8935), .S(n9931), .Z(n8939) );
  NAND2_X1 U10312 ( .A1(n8937), .A2(n8952), .ZN(n8938) );
  OAI211_X1 U10313 ( .C1(n8940), .C2(n8947), .A(n8939), .B(n8938), .ZN(
        P2_U3447) );
  MUX2_X1 U10314 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8941), .S(n9931), .Z(
        P2_U3446) );
  MUX2_X1 U10315 ( .A(n8943), .B(n8942), .S(n9931), .Z(n8946) );
  NAND2_X1 U10316 ( .A1(n8944), .A2(n8952), .ZN(n8945) );
  OAI211_X1 U10317 ( .C1(n8948), .C2(n8947), .A(n8946), .B(n8945), .ZN(
        P2_U3444) );
  INV_X1 U10318 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8950) );
  MUX2_X1 U10319 ( .A(n8950), .B(n8949), .S(n9931), .Z(n8956) );
  AOI22_X1 U10320 ( .A1(n8954), .A2(n8953), .B1(n8952), .B2(n8951), .ZN(n8955)
         );
  NAND2_X1 U10321 ( .A1(n8956), .A2(n8955), .ZN(P2_U3441) );
  INV_X1 U10322 ( .A(n8957), .ZN(n9533) );
  NAND3_X1 U10323 ( .A1(n8959), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8960) );
  OAI22_X1 U10324 ( .A1(n8958), .A2(n8960), .B1(n6440), .B2(n8968), .ZN(n8961)
         );
  INV_X1 U10325 ( .A(n8961), .ZN(n8962) );
  OAI21_X1 U10326 ( .B1(n9533), .B2(n8205), .A(n8962), .ZN(P2_U3264) );
  NAND2_X1 U10327 ( .A1(n8964), .A2(n8963), .ZN(n8966) );
  OAI211_X1 U10328 ( .C1(n8968), .C2(n8967), .A(n8966), .B(n8965), .ZN(
        P2_U3267) );
  MUX2_X1 U10329 ( .A(n8969), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10330 ( .A(n8970), .ZN(n8972) );
  NAND2_X1 U10331 ( .A1(n8972), .A2(n8971), .ZN(n9065) );
  NAND2_X1 U10332 ( .A1(n8970), .A2(n8973), .ZN(n9067) );
  OR2_X1 U10333 ( .A1(n6178), .A2(n9032), .ZN(n8975) );
  AND3_X1 U10334 ( .A1(n9063), .A2(n9067), .A3(n8975), .ZN(n8976) );
  OAI21_X1 U10335 ( .B1(n9033), .B2(n8976), .A(n9109), .ZN(n8981) );
  OAI22_X1 U10336 ( .A1(n9460), .A2(n9070), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8977), .ZN(n8979) );
  OAI22_X1 U10337 ( .A1(n9461), .A2(n9113), .B1(n9112), .B2(n9307), .ZN(n8978)
         );
  NAND2_X1 U10338 ( .A1(n8981), .A2(n8980), .ZN(P1_U3216) );
  INV_X1 U10339 ( .A(n8982), .ZN(n9367) );
  AOI22_X1 U10340 ( .A1(n9058), .A2(n9367), .B1(n9116), .B2(n9361), .ZN(n8984)
         );
  OAI211_X1 U10341 ( .C1(n9345), .C2(n9113), .A(n8984), .B(n8983), .ZN(n8992)
         );
  INV_X1 U10342 ( .A(n8987), .ZN(n8988) );
  NAND3_X1 U10343 ( .A1(n8986), .A2(n8989), .A3(n8988), .ZN(n8990) );
  AOI21_X1 U10344 ( .B1(n8985), .B2(n8990), .A(n9075), .ZN(n8991) );
  AOI211_X1 U10345 ( .C1(n9488), .C2(n9084), .A(n8992), .B(n8991), .ZN(n8993)
         );
  INV_X1 U10346 ( .A(n8993), .ZN(P1_U3219) );
  OAI21_X1 U10347 ( .B1(n8996), .B2(n8995), .A(n8994), .ZN(n8997) );
  NAND2_X1 U10348 ( .A1(n8997), .A2(n9109), .ZN(n9002) );
  NOR2_X1 U10349 ( .A1(n9339), .A2(n9112), .ZN(n9000) );
  OAI22_X1 U10350 ( .A1(n9460), .A2(n9113), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8998), .ZN(n8999) );
  AOI211_X1 U10351 ( .C1(n9081), .C2(n9362), .A(n9000), .B(n8999), .ZN(n9001)
         );
  OAI211_X1 U10352 ( .C1(n9337), .C2(n9119), .A(n9002), .B(n9001), .ZN(
        P1_U3223) );
  AOI21_X1 U10353 ( .B1(n9003), .B2(n9005), .A(n9004), .ZN(n9010) );
  NAND2_X1 U10354 ( .A1(n9447), .A2(n9102), .ZN(n9007) );
  AOI22_X1 U10355 ( .A1(n9446), .A2(n9081), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9006) );
  OAI211_X1 U10356 ( .C1(n9112), .C2(n9277), .A(n9007), .B(n9006), .ZN(n9008)
         );
  AOI21_X1 U10357 ( .B1(n9281), .B2(n9084), .A(n9008), .ZN(n9009) );
  OAI21_X1 U10358 ( .B1(n9010), .B2(n9075), .A(n9009), .ZN(P1_U3225) );
  OAI21_X1 U10359 ( .B1(n9013), .B2(n9012), .A(n9011), .ZN(n9014) );
  NAND2_X1 U10360 ( .A1(n9014), .A2(n9109), .ZN(n9021) );
  INV_X1 U10361 ( .A(n9015), .ZN(n9016) );
  OAI22_X1 U10362 ( .A1(n9113), .A2(n9017), .B1(n9112), .B2(n9016), .ZN(n9018)
         );
  AOI211_X1 U10363 ( .C1(n9081), .C2(n9121), .A(n9019), .B(n9018), .ZN(n9020)
         );
  OAI211_X1 U10364 ( .C1(n9022), .C2(n9119), .A(n9021), .B(n9020), .ZN(
        P1_U3226) );
  OAI21_X1 U10365 ( .B1(n9025), .B2(n9024), .A(n9023), .ZN(n9026) );
  NAND2_X1 U10366 ( .A1(n9026), .A2(n9109), .ZN(n9030) );
  OAI22_X1 U10367 ( .A1(n9113), .A2(n9498), .B1(n9112), .B2(n9401), .ZN(n9027)
         );
  AOI211_X1 U10368 ( .C1(n9081), .C2(n9539), .A(n9028), .B(n9027), .ZN(n9029)
         );
  OAI211_X1 U10369 ( .C1(n9397), .C2(n9119), .A(n9030), .B(n9029), .ZN(
        P1_U3228) );
  NAND2_X1 U10370 ( .A1(n9469), .A2(n9081), .ZN(n9036) );
  NAND2_X1 U10371 ( .A1(n9294), .A2(n9058), .ZN(n9035) );
  OAI211_X1 U10372 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9037), .A(n9036), .B(
        n9035), .ZN(n9038) );
  AOI21_X1 U10373 ( .B1(n9262), .B2(n9102), .A(n9038), .ZN(n9039) );
  INV_X1 U10374 ( .A(n9040), .ZN(n9041) );
  NOR3_X1 U10375 ( .A1(n9043), .A2(n9042), .A3(n9041), .ZN(n9046) );
  INV_X1 U10376 ( .A(n9044), .ZN(n9045) );
  OAI21_X1 U10377 ( .B1(n9046), .B2(n9045), .A(n9109), .ZN(n9052) );
  AOI21_X1 U10378 ( .B1(n9102), .B2(n9123), .A(n9047), .ZN(n9051) );
  AOI22_X1 U10379 ( .A1(n9058), .A2(n9048), .B1(n9081), .B2(n9658), .ZN(n9050)
         );
  NAND2_X1 U10380 ( .A1(n9084), .A2(n9660), .ZN(n9049) );
  NAND4_X1 U10381 ( .A1(n9052), .A2(n9051), .A3(n9050), .A4(n9049), .ZN(
        P1_U3231) );
  INV_X1 U10382 ( .A(n9053), .ZN(n9054) );
  NAND3_X1 U10383 ( .A1(n8985), .A2(n9055), .A3(n9054), .ZN(n9056) );
  AOI21_X1 U10384 ( .B1(n9057), .B2(n9056), .A(n9075), .ZN(n9062) );
  AOI22_X1 U10385 ( .A1(n9468), .A2(n9102), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9060) );
  AOI22_X1 U10386 ( .A1(n9058), .A2(n9352), .B1(n9116), .B2(n9382), .ZN(n9059)
         );
  OAI211_X1 U10387 ( .C1(n9354), .C2(n9119), .A(n9060), .B(n9059), .ZN(n9061)
         );
  OR2_X1 U10388 ( .A1(n9062), .A2(n9061), .ZN(P1_U3233) );
  INV_X1 U10389 ( .A(n9063), .ZN(n9068) );
  AOI21_X1 U10390 ( .B1(n9065), .B2(n9067), .A(n9064), .ZN(n9066) );
  AOI21_X1 U10391 ( .B1(n9068), .B2(n9067), .A(n9066), .ZN(n9076) );
  OAI22_X1 U10392 ( .A1(n9325), .A2(n9113), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9069), .ZN(n9073) );
  OAI22_X1 U10393 ( .A1(n9071), .A2(n9070), .B1(n9324), .B2(n9112), .ZN(n9072)
         );
  AOI211_X1 U10394 ( .C1(n9328), .C2(n9084), .A(n9073), .B(n9072), .ZN(n9074)
         );
  OAI21_X1 U10395 ( .B1(n9076), .B2(n9075), .A(n9074), .ZN(P1_U3235) );
  OAI21_X1 U10396 ( .B1(n9079), .B2(n9078), .A(n9077), .ZN(n9080) );
  NAND2_X1 U10397 ( .A1(n9080), .A2(n9109), .ZN(n9087) );
  AOI22_X1 U10398 ( .A1(n9081), .A2(n9599), .B1(n9102), .B2(n9598), .ZN(n9086)
         );
  AOI22_X1 U10399 ( .A1(n9084), .A2(n9083), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9082), .ZN(n9085) );
  NAND3_X1 U10400 ( .A1(n9087), .A2(n9086), .A3(n9085), .ZN(P1_U3237) );
  OAI21_X1 U10401 ( .B1(n9089), .B2(n9088), .A(n8986), .ZN(n9090) );
  NAND2_X1 U10402 ( .A1(n9090), .A2(n9109), .ZN(n9095) );
  OAI22_X1 U10403 ( .A1(n9113), .A2(n9091), .B1(n9112), .B2(n9388), .ZN(n9092)
         );
  AOI211_X1 U10404 ( .C1(n9116), .C2(n9381), .A(n9093), .B(n9092), .ZN(n9094)
         );
  OAI211_X1 U10405 ( .C1(n9096), .C2(n9119), .A(n9095), .B(n9094), .ZN(
        P1_U3238) );
  INV_X1 U10406 ( .A(n9442), .ZN(n9264) );
  OAI21_X1 U10407 ( .B1(n9004), .B2(n9098), .A(n9097), .ZN(n9099) );
  NAND3_X1 U10408 ( .A1(n9100), .A2(n9109), .A3(n9099), .ZN(n9106) );
  INV_X1 U10409 ( .A(n9101), .ZN(n9259) );
  AOI22_X1 U10410 ( .A1(n9102), .A2(n9238), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9103) );
  OAI21_X1 U10411 ( .B1(n9259), .B2(n9112), .A(n9103), .ZN(n9104) );
  AOI21_X1 U10412 ( .B1(n9116), .B2(n9262), .A(n9104), .ZN(n9105) );
  OAI211_X1 U10413 ( .C1(n9264), .C2(n9119), .A(n9106), .B(n9105), .ZN(
        P1_U3240) );
  OAI21_X1 U10414 ( .B1(n4434), .B2(n9108), .A(n9107), .ZN(n9110) );
  NAND2_X1 U10415 ( .A1(n9110), .A2(n9109), .ZN(n9118) );
  OAI22_X1 U10416 ( .A1(n9113), .A2(n9497), .B1(n9112), .B2(n9111), .ZN(n9114)
         );
  AOI211_X1 U10417 ( .C1(n9116), .C2(n9694), .A(n9115), .B(n9114), .ZN(n9117)
         );
  OAI211_X1 U10418 ( .C1(n9542), .C2(n9119), .A(n9118), .B(n9117), .ZN(
        P1_U3241) );
  MUX2_X1 U10419 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9120), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10420 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9238), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10421 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9447), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10422 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9262), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10423 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9446), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10424 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9469), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10425 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9468), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10426 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9362), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10427 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9382), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10428 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9361), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10429 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9381), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10430 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9539), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10431 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9121), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10432 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9694), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10433 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9686), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10434 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9122), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10435 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9669), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10436 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9123), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9553), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10438 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9658), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10439 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9569), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10440 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9639), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10441 ( .A(n9617), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9126), .Z(
        P1_U3559) );
  MUX2_X1 U10442 ( .A(n9124), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9126), .Z(
        P1_U3558) );
  MUX2_X1 U10443 ( .A(n9598), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9126), .Z(
        P1_U3557) );
  MUX2_X1 U10444 ( .A(n9125), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9126), .Z(
        P1_U3556) );
  MUX2_X1 U10445 ( .A(n9599), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9126), .Z(
        P1_U3555) );
  MUX2_X1 U10446 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9127), .S(P1_U3973), .Z(
        P1_U3554) );
  OAI211_X1 U10447 ( .C1(n9130), .C2(n9129), .A(n9204), .B(n9128), .ZN(n9137)
         );
  OAI211_X1 U10448 ( .C1(n9132), .C2(n9131), .A(n9211), .B(n9146), .ZN(n9136)
         );
  AOI22_X1 U10449 ( .A1(n9215), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9135) );
  NAND2_X1 U10450 ( .A1(n9217), .A2(n9133), .ZN(n9134) );
  NAND4_X1 U10451 ( .A1(n9137), .A2(n9136), .A3(n9135), .A4(n9134), .ZN(
        P1_U3244) );
  MUX2_X1 U10452 ( .A(n9140), .B(n9139), .S(n9138), .Z(n9144) );
  NAND2_X1 U10453 ( .A1(n9142), .A2(n9141), .ZN(n9143) );
  OAI211_X1 U10454 ( .C1(n9144), .C2(n6269), .A(P1_U3973), .B(n9143), .ZN(
        n9186) );
  AOI22_X1 U10455 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .B1(
        P1_ADDR_REG_2__SCAN_IN), .B2(n9215), .ZN(n9158) );
  MUX2_X1 U10456 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6443), .S(n9151), .Z(n9147)
         );
  NAND3_X1 U10457 ( .A1(n9147), .A2(n9146), .A3(n9145), .ZN(n9148) );
  NAND2_X1 U10458 ( .A1(n9149), .A2(n9148), .ZN(n9150) );
  OAI22_X1 U10459 ( .A1(n9151), .A2(n9189), .B1(n9165), .B2(n9150), .ZN(n9152)
         );
  INV_X1 U10460 ( .A(n9152), .ZN(n9157) );
  OAI211_X1 U10461 ( .C1(n9155), .C2(n9154), .A(n9204), .B(n9153), .ZN(n9156)
         );
  NAND4_X1 U10462 ( .A1(n9186), .A2(n9158), .A3(n9157), .A4(n9156), .ZN(
        P1_U3245) );
  NOR2_X1 U10463 ( .A1(n9189), .A2(n9159), .ZN(n9160) );
  AOI211_X1 U10464 ( .C1(n9215), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9161), .B(
        n9160), .ZN(n9171) );
  OAI211_X1 U10465 ( .C1(n9164), .C2(n9163), .A(n9204), .B(n9162), .ZN(n9170)
         );
  AOI211_X1 U10466 ( .C1(n9167), .C2(n9166), .A(n9182), .B(n9165), .ZN(n9168)
         );
  INV_X1 U10467 ( .A(n9168), .ZN(n9169) );
  NAND3_X1 U10468 ( .A1(n9171), .A2(n9170), .A3(n9169), .ZN(P1_U3246) );
  NOR2_X1 U10469 ( .A1(n9189), .A2(n9178), .ZN(n9172) );
  AOI211_X1 U10470 ( .C1(n9215), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n9173), .B(
        n9172), .ZN(n9185) );
  OAI211_X1 U10471 ( .C1(n9176), .C2(n9175), .A(n9204), .B(n9174), .ZN(n9184)
         );
  INV_X1 U10472 ( .A(n9177), .ZN(n9180) );
  MUX2_X1 U10473 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6448), .S(n9178), .Z(n9179)
         );
  NAND2_X1 U10474 ( .A1(n9180), .A2(n9179), .ZN(n9181) );
  OAI211_X1 U10475 ( .C1(n9182), .C2(n9181), .A(n9211), .B(n9197), .ZN(n9183)
         );
  NAND4_X1 U10476 ( .A1(n9186), .A2(n9185), .A3(n9184), .A4(n9183), .ZN(
        P1_U3247) );
  INV_X1 U10477 ( .A(n9187), .ZN(n9191) );
  NOR2_X1 U10478 ( .A1(n9189), .A2(n9188), .ZN(n9190) );
  AOI211_X1 U10479 ( .C1(n9215), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n9191), .B(
        n9190), .ZN(n9202) );
  OAI211_X1 U10480 ( .C1(n9194), .C2(n9193), .A(n9204), .B(n9192), .ZN(n9201)
         );
  INV_X1 U10481 ( .A(n9213), .ZN(n9199) );
  NAND3_X1 U10482 ( .A1(n9197), .A2(n9196), .A3(n9195), .ZN(n9198) );
  NAND3_X1 U10483 ( .A1(n9211), .A2(n9199), .A3(n9198), .ZN(n9200) );
  NAND3_X1 U10484 ( .A1(n9202), .A2(n9201), .A3(n9200), .ZN(P1_U3248) );
  OAI211_X1 U10485 ( .C1(n9206), .C2(n9205), .A(n9204), .B(n9203), .ZN(n9221)
         );
  INV_X1 U10486 ( .A(n9207), .ZN(n9209) );
  MUX2_X1 U10487 ( .A(n6450), .B(P1_REG1_REG_6__SCAN_IN), .S(n9216), .Z(n9208)
         );
  NAND2_X1 U10488 ( .A1(n9209), .A2(n9208), .ZN(n9212) );
  OAI211_X1 U10489 ( .C1(n9213), .C2(n9212), .A(n9211), .B(n9210), .ZN(n9220)
         );
  AOI21_X1 U10490 ( .B1(n9215), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n9214), .ZN(
        n9219) );
  NAND2_X1 U10491 ( .A1(n9217), .A2(n9216), .ZN(n9218) );
  NAND4_X1 U10492 ( .A1(n9221), .A2(n9220), .A3(n9219), .A4(n9218), .ZN(
        P1_U3249) );
  XNOR2_X1 U10493 ( .A(n9225), .B(n9222), .ZN(n9223) );
  NAND2_X1 U10494 ( .A1(n9223), .A2(n9581), .ZN(n9415) );
  AOI21_X1 U10495 ( .B1(n9571), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9224), .ZN(
        n9227) );
  NAND2_X1 U10496 ( .A1(n9225), .A2(n9578), .ZN(n9226) );
  OAI211_X1 U10497 ( .C1(n9415), .C2(n9331), .A(n9227), .B(n9226), .ZN(
        P1_U3263) );
  OAI21_X1 U10498 ( .B1(n9232), .B2(n9231), .A(n9230), .ZN(n9425) );
  INV_X1 U10499 ( .A(n9233), .ZN(n9234) );
  AOI211_X1 U10500 ( .C1(n9424), .C2(n4611), .A(n9562), .B(n9234), .ZN(n9422)
         );
  NAND2_X1 U10501 ( .A1(n9422), .A2(n9585), .ZN(n9240) );
  AOI22_X1 U10502 ( .A1(n9571), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9235), .B2(
        n9573), .ZN(n9236) );
  OAI21_X1 U10503 ( .B1(n9407), .B2(n9421), .A(n9236), .ZN(n9237) );
  AOI21_X1 U10504 ( .B1(n9404), .B2(n9238), .A(n9237), .ZN(n9239) );
  OAI211_X1 U10505 ( .C1(n6370), .C2(n9369), .A(n9240), .B(n9239), .ZN(n9241)
         );
  AOI21_X1 U10506 ( .B1(n9425), .B2(n9333), .A(n9241), .ZN(n9242) );
  OAI21_X1 U10507 ( .B1(n9428), .B2(n9414), .A(n9242), .ZN(P1_U3265) );
  XNOR2_X1 U10508 ( .A(n9243), .B(n9244), .ZN(n9436) );
  AOI211_X1 U10509 ( .C1(n9433), .C2(n9257), .A(n9562), .B(n4609), .ZN(n9431)
         );
  NAND2_X1 U10510 ( .A1(n9431), .A2(n9585), .ZN(n9249) );
  AOI22_X1 U10511 ( .A1(n9571), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9573), .B2(
        n9245), .ZN(n9246) );
  OAI21_X1 U10512 ( .B1(n9407), .B2(n9429), .A(n9246), .ZN(n9247) );
  AOI21_X1 U10513 ( .B1(n9447), .B2(n9404), .A(n9247), .ZN(n9248) );
  OAI211_X1 U10514 ( .C1(n9250), .C2(n9369), .A(n9249), .B(n9248), .ZN(n9251)
         );
  AOI21_X1 U10515 ( .B1(n9434), .B2(n9333), .A(n9251), .ZN(n9252) );
  OAI21_X1 U10516 ( .B1(n9436), .B2(n9414), .A(n9252), .ZN(P1_U3266) );
  AOI21_X1 U10517 ( .B1(n9254), .B2(n9255), .A(n9253), .ZN(n9445) );
  XOR2_X1 U10518 ( .A(n9256), .B(n9255), .Z(n9437) );
  NAND2_X1 U10519 ( .A1(n9437), .A2(n9586), .ZN(n9267) );
  AOI211_X1 U10520 ( .C1(n9442), .C2(n9275), .A(n9562), .B(n4608), .ZN(n9440)
         );
  OAI22_X1 U10521 ( .A1(n9438), .A2(n9407), .B1(n9393), .B2(n9258), .ZN(n9261)
         );
  NOR2_X1 U10522 ( .A1(n9259), .A2(n9402), .ZN(n9260) );
  AOI211_X1 U10523 ( .C1(n9404), .C2(n9262), .A(n9261), .B(n9260), .ZN(n9263)
         );
  OAI21_X1 U10524 ( .B1(n9264), .B2(n9369), .A(n9263), .ZN(n9265) );
  AOI21_X1 U10525 ( .B1(n9440), .B2(n9585), .A(n9265), .ZN(n9266) );
  OAI211_X1 U10526 ( .C1(n9445), .C2(n9268), .A(n9267), .B(n9266), .ZN(
        P1_U3267) );
  XNOR2_X1 U10527 ( .A(n9269), .B(n9271), .ZN(n9454) );
  INV_X1 U10528 ( .A(n9270), .ZN(n9274) );
  OAI21_X1 U10529 ( .B1(n4379), .B2(n9272), .A(n9271), .ZN(n9273) );
  NAND2_X1 U10530 ( .A1(n9274), .A2(n9273), .ZN(n9452) );
  OAI211_X1 U10531 ( .C1(n9450), .C2(n9293), .A(n9581), .B(n9275), .ZN(n9449)
         );
  OAI22_X1 U10532 ( .A1(n9277), .A2(n9402), .B1(n9276), .B2(n9393), .ZN(n9278)
         );
  AOI21_X1 U10533 ( .B1(n9404), .B2(n9446), .A(n9278), .ZN(n9279) );
  OAI21_X1 U10534 ( .B1(n9430), .B2(n9407), .A(n9279), .ZN(n9280) );
  AOI21_X1 U10535 ( .B1(n9281), .B2(n9578), .A(n9280), .ZN(n9282) );
  OAI21_X1 U10536 ( .B1(n9449), .B2(n9331), .A(n9282), .ZN(n9283) );
  AOI21_X1 U10537 ( .B1(n9452), .B2(n9333), .A(n9283), .ZN(n9284) );
  OAI21_X1 U10538 ( .B1(n9454), .B2(n9414), .A(n9284), .ZN(P1_U3268) );
  AOI211_X1 U10539 ( .C1(n9289), .C2(n9285), .A(n9712), .B(n4379), .ZN(n9287)
         );
  OAI22_X1 U10540 ( .A1(n9439), .A2(n9703), .B1(n9325), .B2(n9705), .ZN(n9286)
         );
  NOR2_X1 U10541 ( .A1(n9287), .A2(n9286), .ZN(n9458) );
  OAI21_X1 U10542 ( .B1(n9290), .B2(n9289), .A(n9288), .ZN(n9459) );
  INV_X1 U10543 ( .A(n9459), .ZN(n9299) );
  NAND2_X1 U10544 ( .A1(n9456), .A2(n9302), .ZN(n9291) );
  NAND2_X1 U10545 ( .A1(n9291), .A2(n9581), .ZN(n9292) );
  NOR2_X1 U10546 ( .A1(n9293), .A2(n9292), .ZN(n9455) );
  NAND2_X1 U10547 ( .A1(n9455), .A2(n9585), .ZN(n9296) );
  AOI22_X1 U10548 ( .A1(n9294), .A2(n9573), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9571), .ZN(n9295) );
  OAI211_X1 U10549 ( .C1(n9297), .C2(n9369), .A(n9296), .B(n9295), .ZN(n9298)
         );
  AOI21_X1 U10550 ( .B1(n9299), .B2(n9586), .A(n9298), .ZN(n9300) );
  OAI21_X1 U10551 ( .B1(n9571), .B2(n9458), .A(n9300), .ZN(P1_U3269) );
  XOR2_X1 U10552 ( .A(n9312), .B(n9301), .Z(n9467) );
  AOI21_X1 U10553 ( .B1(n9322), .B2(n9464), .A(n9562), .ZN(n9303) );
  AND2_X1 U10554 ( .A1(n9303), .A2(n9302), .ZN(n9462) );
  NAND2_X1 U10555 ( .A1(n9464), .A2(n9578), .ZN(n9311) );
  NAND2_X1 U10556 ( .A1(n9304), .A2(n9404), .ZN(n9306) );
  NAND2_X1 U10557 ( .A1(n9571), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9305) );
  OAI211_X1 U10558 ( .C1(n9402), .C2(n9307), .A(n9306), .B(n9305), .ZN(n9308)
         );
  AOI21_X1 U10559 ( .B1(n9446), .B2(n9309), .A(n9308), .ZN(n9310) );
  NAND2_X1 U10560 ( .A1(n9311), .A2(n9310), .ZN(n9316) );
  XNOR2_X1 U10561 ( .A(n9313), .B(n9312), .ZN(n9314) );
  NAND2_X1 U10562 ( .A1(n9314), .A2(n9666), .ZN(n9465) );
  NOR2_X1 U10563 ( .A1(n9465), .A2(n9571), .ZN(n9315) );
  AOI211_X1 U10564 ( .C1(n9462), .C2(n9585), .A(n9316), .B(n9315), .ZN(n9317)
         );
  OAI21_X1 U10565 ( .B1(n9467), .B2(n9414), .A(n9317), .ZN(P1_U3270) );
  XNOR2_X1 U10566 ( .A(n9319), .B(n9318), .ZN(n9476) );
  XNOR2_X1 U10567 ( .A(n9321), .B(n9320), .ZN(n9474) );
  OAI211_X1 U10568 ( .C1(n9472), .C2(n4433), .A(n9581), .B(n9322), .ZN(n9471)
         );
  OAI22_X1 U10569 ( .A1(n9324), .A2(n9402), .B1(n9323), .B2(n9393), .ZN(n9327)
         );
  NOR2_X1 U10570 ( .A1(n9325), .A2(n9407), .ZN(n9326) );
  AOI211_X1 U10571 ( .C1(n9404), .C2(n9468), .A(n9327), .B(n9326), .ZN(n9330)
         );
  NAND2_X1 U10572 ( .A1(n9328), .A2(n9578), .ZN(n9329) );
  OAI211_X1 U10573 ( .C1(n9471), .C2(n9331), .A(n9330), .B(n9329), .ZN(n9332)
         );
  AOI21_X1 U10574 ( .B1(n9474), .B2(n9333), .A(n9332), .ZN(n9334) );
  OAI21_X1 U10575 ( .B1(n9476), .B2(n9414), .A(n9334), .ZN(P1_U3271) );
  XNOR2_X1 U10576 ( .A(n9336), .B(n9335), .ZN(n9481) );
  AOI211_X1 U10577 ( .C1(n9479), .C2(n9350), .A(n9562), .B(n4433), .ZN(n9478)
         );
  NOR2_X1 U10578 ( .A1(n9337), .A2(n9369), .ZN(n9341) );
  OAI22_X1 U10579 ( .A1(n9339), .A2(n9402), .B1(n9393), .B2(n9338), .ZN(n9340)
         );
  AOI211_X1 U10580 ( .C1(n9478), .C2(n9585), .A(n9341), .B(n9340), .ZN(n9347)
         );
  XNOR2_X1 U10581 ( .A(n9343), .B(n9342), .ZN(n9344) );
  OAI222_X1 U10582 ( .A1(n9703), .A2(n9460), .B1(n9705), .B2(n9345), .C1(n9712), .C2(n9344), .ZN(n9477) );
  NAND2_X1 U10583 ( .A1(n9477), .A2(n9393), .ZN(n9346) );
  OAI211_X1 U10584 ( .C1(n9481), .C2(n9414), .A(n9347), .B(n9346), .ZN(
        P1_U3272) );
  XOR2_X1 U10585 ( .A(n9348), .B(n9356), .Z(n9349) );
  AOI222_X1 U10586 ( .A1(n9666), .A2(n9349), .B1(n9468), .B2(n9695), .C1(n9382), .C2(n9659), .ZN(n9485) );
  INV_X1 U10587 ( .A(n9350), .ZN(n9351) );
  AOI211_X1 U10588 ( .C1(n9483), .C2(n9365), .A(n9351), .B(n9562), .ZN(n9482)
         );
  AOI22_X1 U10589 ( .A1(n9352), .A2(n9573), .B1(n9571), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9353) );
  OAI21_X1 U10590 ( .B1(n9354), .B2(n9369), .A(n9353), .ZN(n9358) );
  XOR2_X1 U10591 ( .A(n9356), .B(n9355), .Z(n9486) );
  NOR2_X1 U10592 ( .A1(n9486), .A2(n9414), .ZN(n9357) );
  AOI211_X1 U10593 ( .C1(n9482), .C2(n9585), .A(n9358), .B(n9357), .ZN(n9359)
         );
  OAI21_X1 U10594 ( .B1(n9571), .B2(n9485), .A(n9359), .ZN(P1_U3273) );
  XOR2_X1 U10595 ( .A(n9360), .B(n9372), .Z(n9363) );
  AOI222_X1 U10596 ( .A1(n9666), .A2(n9363), .B1(n9362), .B2(n9695), .C1(n9361), .C2(n9659), .ZN(n9490) );
  INV_X1 U10597 ( .A(n9365), .ZN(n9366) );
  AOI211_X1 U10598 ( .C1(n9488), .C2(n9385), .A(n9562), .B(n9366), .ZN(n9487)
         );
  AOI22_X1 U10599 ( .A1(n9571), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9367), .B2(
        n9573), .ZN(n9368) );
  OAI21_X1 U10600 ( .B1(n9370), .B2(n9369), .A(n9368), .ZN(n9374) );
  XOR2_X1 U10601 ( .A(n9372), .B(n9371), .Z(n9491) );
  NOR2_X1 U10602 ( .A1(n9491), .A2(n9414), .ZN(n9373) );
  AOI211_X1 U10603 ( .C1(n9487), .C2(n9585), .A(n9374), .B(n9373), .ZN(n9375)
         );
  OAI21_X1 U10604 ( .B1(n9571), .B2(n9490), .A(n9375), .ZN(P1_U3274) );
  XNOR2_X1 U10605 ( .A(n9377), .B(n9376), .ZN(n9496) );
  OAI211_X1 U10606 ( .C1(n9380), .C2(n9379), .A(n9378), .B(n9666), .ZN(n9384)
         );
  AOI22_X1 U10607 ( .A1(n9382), .A2(n9695), .B1(n9659), .B2(n9381), .ZN(n9383)
         );
  NAND2_X1 U10608 ( .A1(n9384), .A2(n9383), .ZN(n9492) );
  AOI21_X1 U10609 ( .B1(n9494), .B2(n9399), .A(n9562), .ZN(n9386) );
  AND2_X1 U10610 ( .A1(n9386), .A2(n9385), .ZN(n9493) );
  NAND2_X1 U10611 ( .A1(n9493), .A2(n9585), .ZN(n9391) );
  NAND2_X1 U10612 ( .A1(n9571), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9387) );
  OAI21_X1 U10613 ( .B1(n9402), .B2(n9388), .A(n9387), .ZN(n9389) );
  AOI21_X1 U10614 ( .B1(n9494), .B2(n9578), .A(n9389), .ZN(n9390) );
  NAND2_X1 U10615 ( .A1(n9391), .A2(n9390), .ZN(n9392) );
  AOI21_X1 U10616 ( .B1(n9492), .B2(n9393), .A(n9392), .ZN(n9394) );
  OAI21_X1 U10617 ( .B1(n9496), .B2(n9414), .A(n9394), .ZN(P1_U3275) );
  XOR2_X1 U10618 ( .A(n9409), .B(n9395), .Z(n9504) );
  OR2_X1 U10619 ( .A1(n9397), .A2(n9396), .ZN(n9398) );
  AND3_X1 U10620 ( .A1(n9399), .A2(n9398), .A3(n9581), .ZN(n9499) );
  NAND2_X1 U10621 ( .A1(n9501), .A2(n9578), .ZN(n9406) );
  NAND2_X1 U10622 ( .A1(n9571), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9400) );
  OAI21_X1 U10623 ( .B1(n9402), .B2(n9401), .A(n9400), .ZN(n9403) );
  AOI21_X1 U10624 ( .B1(n9404), .B2(n9539), .A(n9403), .ZN(n9405) );
  OAI211_X1 U10625 ( .C1(n9498), .C2(n9407), .A(n9406), .B(n9405), .ZN(n9412)
         );
  OAI211_X1 U10626 ( .C1(n9410), .C2(n9409), .A(n9666), .B(n9408), .ZN(n9502)
         );
  NOR2_X1 U10627 ( .A1(n9502), .A2(n9571), .ZN(n9411) );
  AOI211_X1 U10628 ( .C1(n9499), .C2(n9585), .A(n9412), .B(n9411), .ZN(n9413)
         );
  OAI21_X1 U10629 ( .B1(n9504), .B2(n9414), .A(n9413), .ZN(P1_U3276) );
  OAI211_X1 U10630 ( .C1(n9416), .C2(n9678), .A(n9415), .B(n9417), .ZN(n9510)
         );
  MUX2_X1 U10631 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9510), .S(n9740), .Z(
        P1_U3553) );
  OAI211_X1 U10632 ( .C1(n9419), .C2(n9678), .A(n9418), .B(n9417), .ZN(n9511)
         );
  MUX2_X1 U10633 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9511), .S(n9740), .Z(
        P1_U3552) );
  MUX2_X1 U10634 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9420), .S(n9740), .Z(
        P1_U3551) );
  OAI22_X1 U10635 ( .A1(n9438), .A2(n9705), .B1(n9421), .B2(n9703), .ZN(n9423)
         );
  AOI211_X1 U10636 ( .C1(n9708), .C2(n9424), .A(n9423), .B(n9422), .ZN(n9427)
         );
  NAND2_X1 U10637 ( .A1(n9425), .A2(n9666), .ZN(n9426) );
  OAI211_X1 U10638 ( .C1(n9428), .C2(n9663), .A(n9427), .B(n9426), .ZN(n9512)
         );
  MUX2_X1 U10639 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9512), .S(n9740), .Z(
        P1_U3550) );
  OAI22_X1 U10640 ( .A1(n9430), .A2(n9705), .B1(n9429), .B2(n9703), .ZN(n9432)
         );
  AOI211_X1 U10641 ( .C1(n9708), .C2(n9433), .A(n9432), .B(n9431), .ZN(n9435)
         );
  MUX2_X1 U10642 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9513), .S(n9740), .Z(
        P1_U3549) );
  NAND2_X1 U10643 ( .A1(n9437), .A2(n9716), .ZN(n9444) );
  OAI22_X1 U10644 ( .A1(n9439), .A2(n9705), .B1(n9438), .B2(n9703), .ZN(n9441)
         );
  AOI211_X1 U10645 ( .C1(n9708), .C2(n9442), .A(n9441), .B(n9440), .ZN(n9443)
         );
  OAI211_X1 U10646 ( .C1(n9712), .C2(n9445), .A(n9444), .B(n9443), .ZN(n9514)
         );
  MUX2_X1 U10647 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9514), .S(n9740), .Z(
        P1_U3548) );
  AOI22_X1 U10648 ( .A1(n9447), .A2(n9695), .B1(n9659), .B2(n9446), .ZN(n9448)
         );
  OAI211_X1 U10649 ( .C1(n9450), .C2(n9678), .A(n9449), .B(n9448), .ZN(n9451)
         );
  AOI21_X1 U10650 ( .B1(n9452), .B2(n9666), .A(n9451), .ZN(n9453) );
  OAI21_X1 U10651 ( .B1(n9454), .B2(n9663), .A(n9453), .ZN(n9515) );
  MUX2_X1 U10652 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9515), .S(n9740), .Z(
        P1_U3547) );
  AOI21_X1 U10653 ( .B1(n9708), .B2(n9456), .A(n9455), .ZN(n9457) );
  OAI211_X1 U10654 ( .C1(n9459), .C2(n9663), .A(n9458), .B(n9457), .ZN(n9516)
         );
  MUX2_X1 U10655 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9516), .S(n9740), .Z(
        P1_U3546) );
  OAI22_X1 U10656 ( .A1(n9461), .A2(n9703), .B1(n9460), .B2(n9705), .ZN(n9463)
         );
  AOI211_X1 U10657 ( .C1(n9708), .C2(n9464), .A(n9463), .B(n9462), .ZN(n9466)
         );
  OAI211_X1 U10658 ( .C1(n9467), .C2(n9663), .A(n9466), .B(n9465), .ZN(n9517)
         );
  MUX2_X1 U10659 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9517), .S(n9740), .Z(
        P1_U3545) );
  AOI22_X1 U10660 ( .A1(n9469), .A2(n9695), .B1(n9659), .B2(n9468), .ZN(n9470)
         );
  OAI211_X1 U10661 ( .C1(n9472), .C2(n9678), .A(n9471), .B(n9470), .ZN(n9473)
         );
  AOI21_X1 U10662 ( .B1(n9474), .B2(n9666), .A(n9473), .ZN(n9475) );
  OAI21_X1 U10663 ( .B1(n9476), .B2(n9663), .A(n9475), .ZN(n9518) );
  MUX2_X1 U10664 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9518), .S(n9740), .Z(
        P1_U3544) );
  AOI211_X1 U10665 ( .C1(n9708), .C2(n9479), .A(n9478), .B(n9477), .ZN(n9480)
         );
  OAI21_X1 U10666 ( .B1(n9481), .B2(n9663), .A(n9480), .ZN(n9519) );
  MUX2_X1 U10667 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9519), .S(n9740), .Z(
        P1_U3543) );
  AOI21_X1 U10668 ( .B1(n9708), .B2(n9483), .A(n9482), .ZN(n9484) );
  OAI211_X1 U10669 ( .C1(n9486), .C2(n9663), .A(n9485), .B(n9484), .ZN(n9520)
         );
  MUX2_X1 U10670 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9520), .S(n9740), .Z(
        P1_U3542) );
  AOI21_X1 U10671 ( .B1(n9708), .B2(n9488), .A(n9487), .ZN(n9489) );
  OAI211_X1 U10672 ( .C1(n9491), .C2(n9663), .A(n9490), .B(n9489), .ZN(n9521)
         );
  MUX2_X1 U10673 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9521), .S(n9740), .Z(
        P1_U3541) );
  AOI211_X1 U10674 ( .C1(n9708), .C2(n9494), .A(n9493), .B(n9492), .ZN(n9495)
         );
  OAI21_X1 U10675 ( .B1(n9496), .B2(n9663), .A(n9495), .ZN(n9522) );
  MUX2_X1 U10676 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9522), .S(n9740), .Z(
        P1_U3540) );
  OAI22_X1 U10677 ( .A1(n9498), .A2(n9703), .B1(n9497), .B2(n9705), .ZN(n9500)
         );
  AOI211_X1 U10678 ( .C1(n9708), .C2(n9501), .A(n9500), .B(n9499), .ZN(n9503)
         );
  OAI211_X1 U10679 ( .C1(n9504), .C2(n9663), .A(n9503), .B(n9502), .ZN(n9523)
         );
  MUX2_X1 U10680 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9523), .S(n9740), .Z(
        P1_U3539) );
  AOI211_X1 U10681 ( .C1(n9708), .C2(n9507), .A(n9506), .B(n9505), .ZN(n9508)
         );
  OAI21_X1 U10682 ( .B1(n9509), .B2(n9663), .A(n9508), .ZN(n9524) );
  MUX2_X1 U10683 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9524), .S(n9740), .Z(
        P1_U3538) );
  MUX2_X1 U10684 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9510), .S(n9719), .Z(
        P1_U3521) );
  MUX2_X1 U10685 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9511), .S(n9719), .Z(
        P1_U3520) );
  MUX2_X1 U10686 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9512), .S(n9719), .Z(
        P1_U3518) );
  MUX2_X1 U10687 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9513), .S(n9719), .Z(
        P1_U3517) );
  MUX2_X1 U10688 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9514), .S(n9719), .Z(
        P1_U3516) );
  MUX2_X1 U10689 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9515), .S(n9719), .Z(
        P1_U3515) );
  MUX2_X1 U10690 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9516), .S(n9719), .Z(
        P1_U3514) );
  MUX2_X1 U10691 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9517), .S(n9719), .Z(
        P1_U3513) );
  MUX2_X1 U10692 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9518), .S(n9719), .Z(
        P1_U3512) );
  MUX2_X1 U10693 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9519), .S(n9719), .Z(
        P1_U3511) );
  MUX2_X1 U10694 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9520), .S(n9719), .Z(
        P1_U3510) );
  MUX2_X1 U10695 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9521), .S(n9719), .Z(
        P1_U3509) );
  MUX2_X1 U10696 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9522), .S(n9719), .Z(
        P1_U3507) );
  MUX2_X1 U10697 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9523), .S(n9719), .Z(
        P1_U3504) );
  MUX2_X1 U10698 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9524), .S(n9719), .Z(
        P1_U3501) );
  NAND2_X1 U10699 ( .A1(n9526), .A2(n9525), .ZN(n9528) );
  NOR4_X1 U10700 ( .A1(n9528), .A2(P1_U3086), .A3(n9527), .A4(
        P1_IR_REG_29__SCAN_IN), .ZN(n9530) );
  AOI22_X1 U10701 ( .A1(n9531), .A2(n9530), .B1(P2_DATAO_REG_31__SCAN_IN), 
        .B2(n9529), .ZN(n9532) );
  OAI21_X1 U10702 ( .B1(n9533), .B2(n7754), .A(n9532), .ZN(P1_U3324) );
  OAI222_X1 U10703 ( .A1(n9537), .A2(n9536), .B1(n7754), .B2(n9535), .C1(
        P1_U3086), .C2(n9534), .ZN(P1_U3325) );
  MUX2_X1 U10704 ( .A(n9538), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI22_X1 U10705 ( .A1(n9659), .A2(n9694), .B1(n9539), .B2(n9695), .ZN(n9540)
         );
  OAI211_X1 U10706 ( .C1(n9542), .C2(n9678), .A(n9541), .B(n9540), .ZN(n9543)
         );
  AOI211_X1 U10707 ( .C1(n9545), .C2(n9716), .A(n9544), .B(n9543), .ZN(n9548)
         );
  INV_X1 U10708 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9546) );
  AOI22_X1 U10709 ( .A1(n9740), .A2(n9548), .B1(n9546), .B2(n9737), .ZN(
        P1_U3537) );
  INV_X1 U10710 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9547) );
  AOI22_X1 U10711 ( .A1(n9719), .A2(n9548), .B1(n9547), .B2(n9717), .ZN(
        P1_U3498) );
  XNOR2_X1 U10712 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10713 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  XNOR2_X1 U10714 ( .A(n9552), .B(n9549), .ZN(n9556) );
  AND2_X1 U10715 ( .A1(n7112), .A2(n9550), .ZN(n9551) );
  XOR2_X1 U10716 ( .A(n9552), .B(n9551), .Z(n9655) );
  AOI22_X1 U10717 ( .A1(n9659), .A2(n9569), .B1(n9553), .B2(n9695), .ZN(n9554)
         );
  OAI21_X1 U10718 ( .B1(n9655), .B2(n9647), .A(n9554), .ZN(n9555) );
  AOI21_X1 U10719 ( .B1(n9556), .B2(n9666), .A(n9555), .ZN(n9653) );
  NAND2_X1 U10720 ( .A1(n9571), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9559) );
  NAND2_X1 U10721 ( .A1(n9573), .A2(n9557), .ZN(n9558) );
  NAND2_X1 U10722 ( .A1(n9559), .A2(n9558), .ZN(n9560) );
  AOI21_X1 U10723 ( .B1(n9578), .B2(n6310), .A(n9560), .ZN(n9567) );
  INV_X1 U10724 ( .A(n9655), .ZN(n9565) );
  AOI211_X1 U10725 ( .C1(n6310), .C2(n9563), .A(n9562), .B(n9561), .ZN(n9651)
         );
  AOI22_X1 U10726 ( .A1(n9565), .A2(n9564), .B1(n9585), .B2(n9651), .ZN(n9566)
         );
  OAI211_X1 U10727 ( .C1(n9571), .C2(n9653), .A(n9567), .B(n9566), .ZN(
        P1_U3285) );
  XOR2_X1 U10728 ( .A(n9579), .B(n9568), .Z(n9570) );
  AOI222_X1 U10729 ( .A1(n9666), .A2(n9570), .B1(n9569), .B2(n9695), .C1(n9617), .C2(n9659), .ZN(n9633) );
  NAND2_X1 U10730 ( .A1(n9571), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9575) );
  NAND2_X1 U10731 ( .A1(n9573), .A2(n9572), .ZN(n9574) );
  NAND2_X1 U10732 ( .A1(n9575), .A2(n9574), .ZN(n9576) );
  AOI21_X1 U10733 ( .B1(n9578), .B2(n9577), .A(n9576), .ZN(n9588) );
  XNOR2_X1 U10734 ( .A(n9580), .B(n9579), .ZN(n9636) );
  OAI211_X1 U10735 ( .C1(n9583), .C2(n9632), .A(n9582), .B(n9581), .ZN(n9631)
         );
  INV_X1 U10736 ( .A(n9631), .ZN(n9584) );
  AOI22_X1 U10737 ( .A1(n9636), .A2(n9586), .B1(n9585), .B2(n9584), .ZN(n9587)
         );
  OAI211_X1 U10738 ( .C1(n9571), .C2(n9633), .A(n9588), .B(n9587), .ZN(
        P1_U3287) );
  AND2_X1 U10739 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9589), .ZN(P1_U3294) );
  AND2_X1 U10740 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9589), .ZN(P1_U3295) );
  AND2_X1 U10741 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9589), .ZN(P1_U3296) );
  AND2_X1 U10742 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9589), .ZN(P1_U3297) );
  AND2_X1 U10743 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9589), .ZN(P1_U3298) );
  AND2_X1 U10744 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9589), .ZN(P1_U3299) );
  AND2_X1 U10745 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9589), .ZN(P1_U3300) );
  AND2_X1 U10746 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9589), .ZN(P1_U3301) );
  AND2_X1 U10747 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9589), .ZN(P1_U3302) );
  AND2_X1 U10748 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9589), .ZN(P1_U3303) );
  AND2_X1 U10749 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9589), .ZN(P1_U3304) );
  AND2_X1 U10750 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9589), .ZN(P1_U3305) );
  AND2_X1 U10751 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9589), .ZN(P1_U3306) );
  AND2_X1 U10752 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9589), .ZN(P1_U3307) );
  AND2_X1 U10753 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9589), .ZN(P1_U3308) );
  AND2_X1 U10754 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9589), .ZN(P1_U3309) );
  AND2_X1 U10755 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9589), .ZN(P1_U3310) );
  AND2_X1 U10756 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9589), .ZN(P1_U3311) );
  AND2_X1 U10757 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9589), .ZN(P1_U3312) );
  AND2_X1 U10758 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9589), .ZN(P1_U3313) );
  AND2_X1 U10759 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9589), .ZN(P1_U3314) );
  AND2_X1 U10760 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9589), .ZN(P1_U3315) );
  AND2_X1 U10761 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9589), .ZN(P1_U3316) );
  AND2_X1 U10762 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9589), .ZN(P1_U3317) );
  AND2_X1 U10763 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9589), .ZN(P1_U3318) );
  AND2_X1 U10764 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9589), .ZN(P1_U3319) );
  AND2_X1 U10765 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9589), .ZN(P1_U3320) );
  AND2_X1 U10766 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9589), .ZN(P1_U3321) );
  AND2_X1 U10767 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9589), .ZN(P1_U3322) );
  AND2_X1 U10768 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9589), .ZN(P1_U3323) );
  INV_X1 U10769 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9590) );
  AOI22_X1 U10770 ( .A1(n9719), .A2(n9591), .B1(n9590), .B2(n9717), .ZN(
        P1_U3453) );
  INV_X1 U10771 ( .A(n9654), .ZN(n9681) );
  OAI21_X1 U10772 ( .B1(n9593), .B2(n9678), .A(n9592), .ZN(n9595) );
  AOI211_X1 U10773 ( .C1(n9681), .C2(n9596), .A(n9595), .B(n9594), .ZN(n9720)
         );
  INV_X1 U10774 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9597) );
  AOI22_X1 U10775 ( .A1(n9719), .A2(n9720), .B1(n9597), .B2(n9717), .ZN(
        P1_U3456) );
  AOI22_X1 U10776 ( .A1(n9659), .A2(n9599), .B1(n9598), .B2(n9695), .ZN(n9600)
         );
  OAI211_X1 U10777 ( .C1(n9602), .C2(n9678), .A(n9601), .B(n9600), .ZN(n9605)
         );
  NOR2_X1 U10778 ( .A1(n9603), .A2(n9663), .ZN(n9604) );
  AOI211_X1 U10779 ( .C1(n9606), .C2(n9666), .A(n9605), .B(n9604), .ZN(n9721)
         );
  INV_X1 U10780 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9607) );
  AOI22_X1 U10781 ( .A1(n9719), .A2(n9721), .B1(n9607), .B2(n9717), .ZN(
        P1_U3459) );
  AOI21_X1 U10782 ( .B1(n9708), .B2(n9609), .A(n9608), .ZN(n9610) );
  OAI211_X1 U10783 ( .C1(n9663), .C2(n9612), .A(n9611), .B(n9610), .ZN(n9613)
         );
  INV_X1 U10784 ( .A(n9613), .ZN(n9723) );
  INV_X1 U10785 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9614) );
  AOI22_X1 U10786 ( .A1(n9719), .A2(n9723), .B1(n9614), .B2(n9717), .ZN(
        P1_U3462) );
  AND2_X1 U10787 ( .A1(n9615), .A2(n9716), .ZN(n9621) );
  AOI22_X1 U10788 ( .A1(n9617), .A2(n9695), .B1(n9708), .B2(n9616), .ZN(n9618)
         );
  NAND2_X1 U10789 ( .A1(n9619), .A2(n9618), .ZN(n9620) );
  NOR3_X1 U10790 ( .A1(n9622), .A2(n9621), .A3(n9620), .ZN(n9724) );
  INV_X1 U10791 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9623) );
  AOI22_X1 U10792 ( .A1(n9719), .A2(n9724), .B1(n9623), .B2(n9717), .ZN(
        P1_U3465) );
  AND2_X1 U10793 ( .A1(n9624), .A2(n9716), .ZN(n9628) );
  OAI21_X1 U10794 ( .B1(n9626), .B2(n9678), .A(n9625), .ZN(n9627) );
  NOR3_X1 U10795 ( .A1(n9629), .A2(n9628), .A3(n9627), .ZN(n9726) );
  INV_X1 U10796 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9630) );
  AOI22_X1 U10797 ( .A1(n9719), .A2(n9726), .B1(n9630), .B2(n9717), .ZN(
        P1_U3468) );
  OAI21_X1 U10798 ( .B1(n9632), .B2(n9678), .A(n9631), .ZN(n9635) );
  INV_X1 U10799 ( .A(n9633), .ZN(n9634) );
  AOI211_X1 U10800 ( .C1(n9716), .C2(n9636), .A(n9635), .B(n9634), .ZN(n9727)
         );
  INV_X1 U10801 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9637) );
  AOI22_X1 U10802 ( .A1(n9719), .A2(n9727), .B1(n9637), .B2(n9717), .ZN(
        P1_U3471) );
  INV_X1 U10803 ( .A(n4352), .ZN(n9642) );
  AOI22_X1 U10804 ( .A1(n9659), .A2(n9639), .B1(n9658), .B2(n9695), .ZN(n9640)
         );
  OAI211_X1 U10805 ( .C1(n9642), .C2(n9678), .A(n9641), .B(n9640), .ZN(n9644)
         );
  AOI211_X1 U10806 ( .C1(n9681), .C2(n9645), .A(n9644), .B(n9643), .ZN(n9646)
         );
  OAI21_X1 U10807 ( .B1(n9648), .B2(n9647), .A(n9646), .ZN(n9649) );
  INV_X1 U10808 ( .A(n9649), .ZN(n9729) );
  INV_X1 U10809 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9650) );
  AOI22_X1 U10810 ( .A1(n9719), .A2(n9729), .B1(n9650), .B2(n9717), .ZN(
        P1_U3474) );
  AOI21_X1 U10811 ( .B1(n9708), .B2(n6310), .A(n9651), .ZN(n9652) );
  OAI211_X1 U10812 ( .C1(n9655), .C2(n9654), .A(n9653), .B(n9652), .ZN(n9656)
         );
  INV_X1 U10813 ( .A(n9656), .ZN(n9731) );
  INV_X1 U10814 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9657) );
  AOI22_X1 U10815 ( .A1(n9719), .A2(n9731), .B1(n9657), .B2(n9717), .ZN(
        P1_U3477) );
  AOI22_X1 U10816 ( .A1(n9660), .A2(n9708), .B1(n9659), .B2(n9658), .ZN(n9661)
         );
  OAI211_X1 U10817 ( .C1(n9664), .C2(n9663), .A(n9662), .B(n9661), .ZN(n9665)
         );
  AOI21_X1 U10818 ( .B1(n9667), .B2(n9666), .A(n9665), .ZN(n9732) );
  INV_X1 U10819 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9668) );
  AOI22_X1 U10820 ( .A1(n9719), .A2(n9732), .B1(n9668), .B2(n9717), .ZN(
        P1_U3480) );
  AOI22_X1 U10821 ( .A1(n9670), .A2(n9708), .B1(n9695), .B2(n9669), .ZN(n9672)
         );
  NAND3_X1 U10822 ( .A1(n9673), .A2(n9672), .A3(n9671), .ZN(n9674) );
  AOI21_X1 U10823 ( .B1(n9716), .B2(n9675), .A(n9674), .ZN(n9733) );
  INV_X1 U10824 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9676) );
  AOI22_X1 U10825 ( .A1(n9719), .A2(n9733), .B1(n9676), .B2(n9717), .ZN(
        P1_U3483) );
  OAI21_X1 U10826 ( .B1(n9679), .B2(n9678), .A(n9677), .ZN(n9680) );
  AOI21_X1 U10827 ( .B1(n9682), .B2(n9681), .A(n9680), .ZN(n9683) );
  AND2_X1 U10828 ( .A1(n9684), .A2(n9683), .ZN(n9734) );
  INV_X1 U10829 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9685) );
  AOI22_X1 U10830 ( .A1(n9719), .A2(n9734), .B1(n9685), .B2(n9717), .ZN(
        P1_U3486) );
  AOI22_X1 U10831 ( .A1(n9687), .A2(n9708), .B1(n9695), .B2(n9686), .ZN(n9689)
         );
  NAND3_X1 U10832 ( .A1(n9690), .A2(n9689), .A3(n9688), .ZN(n9691) );
  AOI21_X1 U10833 ( .B1(n9716), .B2(n9692), .A(n9691), .ZN(n9735) );
  INV_X1 U10834 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9693) );
  AOI22_X1 U10835 ( .A1(n9719), .A2(n9735), .B1(n9693), .B2(n9717), .ZN(
        P1_U3489) );
  AOI22_X1 U10836 ( .A1(n9696), .A2(n9708), .B1(n9695), .B2(n9694), .ZN(n9698)
         );
  NAND3_X1 U10837 ( .A1(n9699), .A2(n9698), .A3(n9697), .ZN(n9700) );
  AOI21_X1 U10838 ( .B1(n9716), .B2(n9701), .A(n9700), .ZN(n9736) );
  INV_X1 U10839 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9702) );
  AOI22_X1 U10840 ( .A1(n9719), .A2(n9736), .B1(n9702), .B2(n9717), .ZN(
        P1_U3492) );
  OAI22_X1 U10841 ( .A1(n9706), .A2(n9705), .B1(n9704), .B2(n9703), .ZN(n9707)
         );
  AOI21_X1 U10842 ( .B1(n9709), .B2(n9708), .A(n9707), .ZN(n9711) );
  OAI211_X1 U10843 ( .C1(n9713), .C2(n9712), .A(n9711), .B(n9710), .ZN(n9714)
         );
  AOI21_X1 U10844 ( .B1(n9716), .B2(n9715), .A(n9714), .ZN(n9739) );
  INV_X1 U10845 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9718) );
  AOI22_X1 U10846 ( .A1(n9719), .A2(n9739), .B1(n9718), .B2(n9717), .ZN(
        P1_U3495) );
  AOI22_X1 U10847 ( .A1(n9740), .A2(n9720), .B1(n6444), .B2(n9737), .ZN(
        P1_U3523) );
  AOI22_X1 U10848 ( .A1(n9740), .A2(n9721), .B1(n6443), .B2(n9737), .ZN(
        P1_U3524) );
  AOI22_X1 U10849 ( .A1(n9740), .A2(n9723), .B1(n9722), .B2(n9737), .ZN(
        P1_U3525) );
  AOI22_X1 U10850 ( .A1(n9740), .A2(n9724), .B1(n6448), .B2(n9737), .ZN(
        P1_U3526) );
  AOI22_X1 U10851 ( .A1(n9740), .A2(n9726), .B1(n9725), .B2(n9737), .ZN(
        P1_U3527) );
  AOI22_X1 U10852 ( .A1(n9740), .A2(n9727), .B1(n6450), .B2(n9737), .ZN(
        P1_U3528) );
  AOI22_X1 U10853 ( .A1(n9740), .A2(n9729), .B1(n9728), .B2(n9737), .ZN(
        P1_U3529) );
  AOI22_X1 U10854 ( .A1(n9740), .A2(n9731), .B1(n9730), .B2(n9737), .ZN(
        P1_U3530) );
  AOI22_X1 U10855 ( .A1(n9740), .A2(n9732), .B1(n6500), .B2(n9737), .ZN(
        P1_U3531) );
  AOI22_X1 U10856 ( .A1(n9740), .A2(n9733), .B1(n6535), .B2(n9737), .ZN(
        P1_U3532) );
  AOI22_X1 U10857 ( .A1(n9740), .A2(n9734), .B1(n6550), .B2(n9737), .ZN(
        P1_U3533) );
  AOI22_X1 U10858 ( .A1(n9740), .A2(n9735), .B1(n6774), .B2(n9737), .ZN(
        P1_U3534) );
  AOI22_X1 U10859 ( .A1(n9740), .A2(n9736), .B1(n6813), .B2(n9737), .ZN(
        P1_U3535) );
  AOI22_X1 U10860 ( .A1(n9740), .A2(n9739), .B1(n9738), .B2(n9737), .ZN(
        P1_U3536) );
  NAND2_X1 U10861 ( .A1(n9741), .A2(n6598), .ZN(n9742) );
  AND2_X1 U10862 ( .A1(n9743), .A2(n9742), .ZN(n9744) );
  OAI22_X1 U10863 ( .A1(n9835), .A2(n9745), .B1(n9829), .B2(n9744), .ZN(n9748)
         );
  INV_X1 U10864 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9746) );
  NOR2_X1 U10865 ( .A1(n9783), .A2(n9746), .ZN(n9747) );
  NOR2_X1 U10866 ( .A1(n9748), .A2(n9747), .ZN(n9760) );
  OAI21_X1 U10867 ( .B1(n9751), .B2(n9750), .A(n9749), .ZN(n9752) );
  NAND2_X1 U10868 ( .A1(n9752), .A2(n9832), .ZN(n9758) );
  INV_X1 U10869 ( .A(n9753), .ZN(n9754) );
  AOI21_X1 U10870 ( .B1(n6597), .B2(n9755), .A(n9754), .ZN(n9756) );
  OR2_X1 U10871 ( .A1(n9825), .A2(n9756), .ZN(n9757) );
  NAND4_X1 U10872 ( .A1(n9760), .A2(n9759), .A3(n9758), .A4(n9757), .ZN(
        P2_U3185) );
  INV_X1 U10873 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n9968) );
  OR3_X1 U10874 ( .A1(n9763), .A2(n9762), .A3(n9761), .ZN(n9764) );
  AOI21_X1 U10875 ( .B1(n9765), .B2(n9764), .A(n9829), .ZN(n9776) );
  INV_X1 U10876 ( .A(n9766), .ZN(n9767) );
  NAND3_X1 U10877 ( .A1(n9769), .A2(n9768), .A3(n9767), .ZN(n9770) );
  AOI21_X1 U10878 ( .B1(n9771), .B2(n9770), .A(n9825), .ZN(n9775) );
  NOR2_X1 U10879 ( .A1(n9835), .A2(n9772), .ZN(n9773) );
  NOR4_X1 U10880 ( .A1(n9776), .A2(n9775), .A3(n9774), .A4(n9773), .ZN(n9782)
         );
  NOR2_X1 U10881 ( .A1(n9778), .A2(n9777), .ZN(n9779) );
  OAI21_X1 U10882 ( .B1(n9780), .B2(n9779), .A(n9832), .ZN(n9781) );
  OAI211_X1 U10883 ( .C1(n9968), .C2(n9783), .A(n9782), .B(n9781), .ZN(
        P2_U3190) );
  AOI22_X1 U10884 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n9818), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3151), .ZN(n9799) );
  AOI21_X1 U10885 ( .B1(n9785), .B2(n9784), .A(n4442), .ZN(n9796) );
  OAI21_X1 U10886 ( .B1(n9788), .B2(n9787), .A(n9786), .ZN(n9789) );
  NAND2_X1 U10887 ( .A1(n9789), .A2(n9832), .ZN(n9795) );
  AOI21_X1 U10888 ( .B1(n9792), .B2(n9791), .A(n9790), .ZN(n9793) );
  OR2_X1 U10889 ( .A1(n9793), .A2(n9825), .ZN(n9794) );
  OAI211_X1 U10890 ( .C1(n9796), .C2(n9829), .A(n9795), .B(n9794), .ZN(n9797)
         );
  INV_X1 U10891 ( .A(n9797), .ZN(n9798) );
  OAI211_X1 U10892 ( .C1(n9835), .C2(n9800), .A(n9799), .B(n9798), .ZN(
        P2_U3196) );
  AOI22_X1 U10893 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9818), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(P2_U3151), .ZN(n9816) );
  AOI21_X1 U10894 ( .B1(n9803), .B2(n9802), .A(n9801), .ZN(n9813) );
  OAI21_X1 U10895 ( .B1(n9806), .B2(n9805), .A(n9804), .ZN(n9807) );
  NAND2_X1 U10896 ( .A1(n9807), .A2(n9832), .ZN(n9812) );
  AOI21_X1 U10897 ( .B1(n4401), .B2(n9809), .A(n9808), .ZN(n9810) );
  OR2_X1 U10898 ( .A1(n9810), .A2(n9825), .ZN(n9811) );
  OAI211_X1 U10899 ( .C1(n9813), .C2(n9829), .A(n9812), .B(n9811), .ZN(n9814)
         );
  INV_X1 U10900 ( .A(n9814), .ZN(n9815) );
  OAI211_X1 U10901 ( .C1(n9835), .C2(n9817), .A(n9816), .B(n9815), .ZN(
        P2_U3198) );
  AOI22_X1 U10902 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9818), .B1(
        P2_REG3_REG_17__SCAN_IN), .B2(P2_U3151), .ZN(n9833) );
  OAI21_X1 U10903 ( .B1(n9821), .B2(n9820), .A(n9819), .ZN(n9831) );
  AOI21_X1 U10904 ( .B1(n9824), .B2(n9823), .A(n9822), .ZN(n9826) );
  NOR2_X1 U10905 ( .A1(n9826), .A2(n9825), .ZN(n9830) );
  XOR2_X1 U10906 ( .A(n9836), .B(n9840), .Z(n9839) );
  AOI222_X1 U10907 ( .A1(n9851), .A2(n9839), .B1(n9838), .B2(n9853), .C1(n9837), .C2(n9855), .ZN(n9886) );
  XNOR2_X1 U10908 ( .A(n9841), .B(n9840), .ZN(n9884) );
  AOI222_X1 U10909 ( .A1(n9884), .A2(n9845), .B1(n9844), .B2(n9843), .C1(n9883), .C2(n9842), .ZN(n9846) );
  OAI221_X1 U10910 ( .B1(n9871), .B2(n9886), .C1(n9868), .C2(n6598), .A(n9846), 
        .ZN(P2_U3230) );
  NAND3_X1 U10911 ( .A1(n9848), .A2(n9859), .A3(n9847), .ZN(n9849) );
  NAND2_X1 U10912 ( .A1(n9850), .A2(n9849), .ZN(n9852) );
  NAND2_X1 U10913 ( .A1(n9852), .A2(n9851), .ZN(n9857) );
  AOI22_X1 U10914 ( .A1(n9855), .A2(n6675), .B1(n9854), .B2(n9853), .ZN(n9856)
         );
  AND2_X1 U10915 ( .A1(n9857), .A2(n9856), .ZN(n9881) );
  XNOR2_X1 U10916 ( .A(n9858), .B(n9859), .ZN(n9878) );
  NAND2_X1 U10917 ( .A1(n9878), .A2(n9860), .ZN(n9867) );
  OR2_X1 U10918 ( .A1(n9861), .A2(n9913), .ZN(n9879) );
  OAI22_X1 U10919 ( .A1(n9879), .A2(n9864), .B1(n9863), .B2(n9862), .ZN(n9865)
         );
  INV_X1 U10920 ( .A(n9865), .ZN(n9866) );
  AND3_X1 U10921 ( .A1(n9881), .A2(n9867), .A3(n9866), .ZN(n9869) );
  AOI22_X1 U10922 ( .A1(n9871), .A2(n9870), .B1(n9869), .B2(n9868), .ZN(
        P2_U3231) );
  INV_X1 U10923 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9877) );
  OAI22_X1 U10924 ( .A1(n9874), .A2(n9873), .B1(n9872), .B2(n9913), .ZN(n9875)
         );
  NOR2_X1 U10925 ( .A1(n9876), .A2(n9875), .ZN(n9934) );
  AOI22_X1 U10926 ( .A1(n9933), .A2(n9877), .B1(n9934), .B2(n9931), .ZN(
        P2_U3393) );
  INV_X1 U10927 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U10928 ( .A1(n9878), .A2(n9919), .ZN(n9880) );
  AOI22_X1 U10929 ( .A1(n9933), .A2(n9882), .B1(n9935), .B2(n9931), .ZN(
        P2_U3396) );
  INV_X1 U10930 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9887) );
  AOI22_X1 U10931 ( .A1(n9884), .A2(n9919), .B1(n9930), .B2(n9883), .ZN(n9885)
         );
  AND2_X1 U10932 ( .A1(n9886), .A2(n9885), .ZN(n9936) );
  AOI22_X1 U10933 ( .A1(n9933), .A2(n9887), .B1(n9936), .B2(n9931), .ZN(
        P2_U3399) );
  INV_X1 U10934 ( .A(n9888), .ZN(n9892) );
  OAI22_X1 U10935 ( .A1(n9890), .A2(n9925), .B1(n9889), .B2(n9913), .ZN(n9891)
         );
  NOR2_X1 U10936 ( .A1(n9892), .A2(n9891), .ZN(n9937) );
  AOI22_X1 U10937 ( .A1(n9933), .A2(n5233), .B1(n9937), .B2(n9931), .ZN(
        P2_U3402) );
  INV_X1 U10938 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9897) );
  NOR2_X1 U10939 ( .A1(n9893), .A2(n9913), .ZN(n9895) );
  AOI211_X1 U10940 ( .C1(n9919), .C2(n9896), .A(n9895), .B(n9894), .ZN(n9938)
         );
  AOI22_X1 U10941 ( .A1(n9933), .A2(n9897), .B1(n9938), .B2(n9931), .ZN(
        P2_U3405) );
  INV_X1 U10942 ( .A(n9898), .ZN(n9902) );
  OAI21_X1 U10943 ( .B1(n9900), .B2(n9913), .A(n9899), .ZN(n9901) );
  AOI21_X1 U10944 ( .B1(n9902), .B2(n9919), .A(n9901), .ZN(n9940) );
  AOI22_X1 U10945 ( .A1(n9933), .A2(n5262), .B1(n9940), .B2(n9931), .ZN(
        P2_U3408) );
  INV_X1 U10946 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9907) );
  OAI22_X1 U10947 ( .A1(n9904), .A2(n9925), .B1(n9903), .B2(n9913), .ZN(n9905)
         );
  NOR2_X1 U10948 ( .A1(n9906), .A2(n9905), .ZN(n9941) );
  AOI22_X1 U10949 ( .A1(n9933), .A2(n9907), .B1(n9941), .B2(n9931), .ZN(
        P2_U3411) );
  NAND2_X1 U10950 ( .A1(n9908), .A2(n9919), .ZN(n9911) );
  OR2_X1 U10951 ( .A1(n9909), .A2(n9913), .ZN(n9910) );
  AND3_X1 U10952 ( .A1(n9912), .A2(n9911), .A3(n9910), .ZN(n9942) );
  AOI22_X1 U10953 ( .A1(n9933), .A2(n5304), .B1(n9942), .B2(n9931), .ZN(
        P2_U3414) );
  INV_X1 U10954 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9918) );
  NOR2_X1 U10955 ( .A1(n9914), .A2(n9913), .ZN(n9916) );
  AOI211_X1 U10956 ( .C1(n9917), .C2(n9919), .A(n9916), .B(n9915), .ZN(n9943)
         );
  AOI22_X1 U10957 ( .A1(n9933), .A2(n9918), .B1(n9943), .B2(n9931), .ZN(
        P2_U3417) );
  NAND2_X1 U10958 ( .A1(n9920), .A2(n9919), .ZN(n9923) );
  NAND2_X1 U10959 ( .A1(n9921), .A2(n9930), .ZN(n9922) );
  AOI22_X1 U10960 ( .A1(n9933), .A2(n5328), .B1(n9944), .B2(n9931), .ZN(
        P2_U3420) );
  INV_X1 U10961 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9932) );
  NOR2_X1 U10962 ( .A1(n9926), .A2(n9925), .ZN(n9928) );
  AOI211_X1 U10963 ( .C1(n9930), .C2(n9929), .A(n9928), .B(n9927), .ZN(n9946)
         );
  AOI22_X1 U10964 ( .A1(n9933), .A2(n9932), .B1(n9946), .B2(n9931), .ZN(
        P2_U3423) );
  AOI22_X1 U10965 ( .A1(n9947), .A2(n9934), .B1(n5178), .B2(n9945), .ZN(
        P2_U3460) );
  AOI22_X1 U10966 ( .A1(n9947), .A2(n9935), .B1(n6603), .B2(n9945), .ZN(
        P2_U3461) );
  AOI22_X1 U10967 ( .A1(n9947), .A2(n9936), .B1(n6597), .B2(n9945), .ZN(
        P2_U3462) );
  AOI22_X1 U10968 ( .A1(n9947), .A2(n9937), .B1(n6609), .B2(n9945), .ZN(
        P2_U3463) );
  AOI22_X1 U10969 ( .A1(n9947), .A2(n9938), .B1(n6689), .B2(n9945), .ZN(
        P2_U3464) );
  AOI22_X1 U10970 ( .A1(n9947), .A2(n9940), .B1(n9939), .B2(n9945), .ZN(
        P2_U3465) );
  AOI22_X1 U10971 ( .A1(n9947), .A2(n9941), .B1(n6827), .B2(n9945), .ZN(
        P2_U3466) );
  AOI22_X1 U10972 ( .A1(n9947), .A2(n9942), .B1(n5300), .B2(n9945), .ZN(
        P2_U3467) );
  AOI22_X1 U10973 ( .A1(n9947), .A2(n9943), .B1(n7219), .B2(n9945), .ZN(
        P2_U3468) );
  AOI22_X1 U10974 ( .A1(n9947), .A2(n9944), .B1(n7330), .B2(n9945), .ZN(
        P2_U3469) );
  AOI22_X1 U10975 ( .A1(n9947), .A2(n9946), .B1(n7450), .B2(n9945), .ZN(
        P2_U3470) );
  AOI21_X1 U10976 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9953) );
  INV_X1 U10977 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9949) );
  NAND2_X1 U10978 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n9948) );
  NOR2_X1 U10979 ( .A1(n9949), .A2(n9948), .ZN(n9951) );
  NOR2_X1 U10980 ( .A1(n9953), .A2(n9951), .ZN(n9950) );
  XOR2_X1 U10981 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9950), .Z(ADD_1068_U5) );
  XOR2_X1 U10982 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U10983 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10001) );
  NOR2_X1 U10984 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9999) );
  NOR2_X1 U10985 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9997) );
  NOR2_X1 U10986 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9993) );
  NOR2_X1 U10987 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9991) );
  NOR2_X1 U10988 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9987) );
  NOR2_X1 U10989 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9983) );
  NOR2_X1 U10990 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9979) );
  NOR2_X1 U10991 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9975) );
  NOR2_X1 U10992 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9971) );
  NOR2_X1 U10993 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n9967) );
  NOR2_X1 U10994 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9963) );
  NOR2_X1 U10995 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n9961) );
  NOR2_X1 U10996 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9959) );
  NAND2_X1 U10997 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9957) );
  XOR2_X1 U10998 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10228) );
  NAND2_X1 U10999 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n9955) );
  NOR2_X1 U11000 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n9951), .ZN(n9952) );
  NOR2_X1 U11001 ( .A1(n9953), .A2(n9952), .ZN(n10216) );
  XOR2_X1 U11002 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10215) );
  NAND2_X1 U11003 ( .A1(n10216), .A2(n10215), .ZN(n9954) );
  NAND2_X1 U11004 ( .A1(n9955), .A2(n9954), .ZN(n10227) );
  NAND2_X1 U11005 ( .A1(n10228), .A2(n10227), .ZN(n9956) );
  NAND2_X1 U11006 ( .A1(n9957), .A2(n9956), .ZN(n10230) );
  XNOR2_X1 U11007 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10229) );
  NOR2_X1 U11008 ( .A1(n10230), .A2(n10229), .ZN(n9958) );
  NOR2_X1 U11009 ( .A1(n9959), .A2(n9958), .ZN(n10226) );
  XNOR2_X1 U11010 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n10225) );
  NOR2_X1 U11011 ( .A1(n10226), .A2(n10225), .ZN(n9960) );
  NOR2_X1 U11012 ( .A1(n9961), .A2(n9960), .ZN(n10224) );
  XNOR2_X1 U11013 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10223) );
  NOR2_X1 U11014 ( .A1(n10224), .A2(n10223), .ZN(n9962) );
  NOR2_X1 U11015 ( .A1(n9963), .A2(n9962), .ZN(n10222) );
  INV_X1 U11016 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9965) );
  AOI22_X1 U11017 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9965), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(n9964), .ZN(n10221) );
  NOR2_X1 U11018 ( .A1(n10222), .A2(n10221), .ZN(n9966) );
  NOR2_X1 U11019 ( .A1(n9967), .A2(n9966), .ZN(n10220) );
  INV_X1 U11020 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U11021 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9969), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n9968), .ZN(n10219) );
  NOR2_X1 U11022 ( .A1(n10220), .A2(n10219), .ZN(n9970) );
  NOR2_X1 U11023 ( .A1(n9971), .A2(n9970), .ZN(n10218) );
  INV_X1 U11024 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9973) );
  AOI22_X1 U11025 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9973), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n9972), .ZN(n10217) );
  NOR2_X1 U11026 ( .A1(n10218), .A2(n10217), .ZN(n9974) );
  NOR2_X1 U11027 ( .A1(n9975), .A2(n9974), .ZN(n10018) );
  INV_X1 U11028 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9977) );
  AOI22_X1 U11029 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n9977), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n9976), .ZN(n10017) );
  NOR2_X1 U11030 ( .A1(n10018), .A2(n10017), .ZN(n9978) );
  NOR2_X1 U11031 ( .A1(n9979), .A2(n9978), .ZN(n10016) );
  INV_X1 U11032 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9981) );
  AOI22_X1 U11033 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n9981), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n9980), .ZN(n10015) );
  NOR2_X1 U11034 ( .A1(n10016), .A2(n10015), .ZN(n9982) );
  NOR2_X1 U11035 ( .A1(n9983), .A2(n9982), .ZN(n10014) );
  INV_X1 U11036 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9985) );
  AOI22_X1 U11037 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n9985), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n9984), .ZN(n10013) );
  NOR2_X1 U11038 ( .A1(n10014), .A2(n10013), .ZN(n9986) );
  NOR2_X1 U11039 ( .A1(n9987), .A2(n9986), .ZN(n10012) );
  INV_X1 U11040 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9989) );
  AOI22_X1 U11041 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n9989), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n9988), .ZN(n10011) );
  NOR2_X1 U11042 ( .A1(n10012), .A2(n10011), .ZN(n9990) );
  NOR2_X1 U11043 ( .A1(n9991), .A2(n9990), .ZN(n10010) );
  XNOR2_X1 U11044 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10009) );
  NOR2_X1 U11045 ( .A1(n10010), .A2(n10009), .ZN(n9992) );
  NOR2_X1 U11046 ( .A1(n9993), .A2(n9992), .ZN(n10008) );
  INV_X1 U11047 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9995) );
  AOI22_X1 U11048 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9995), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n9994), .ZN(n10007) );
  NOR2_X1 U11049 ( .A1(n10008), .A2(n10007), .ZN(n9996) );
  NOR2_X1 U11050 ( .A1(n9997), .A2(n9996), .ZN(n10006) );
  XNOR2_X1 U11051 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10005) );
  NOR2_X1 U11052 ( .A1(n10006), .A2(n10005), .ZN(n9998) );
  NOR2_X1 U11053 ( .A1(n9999), .A2(n9998), .ZN(n10004) );
  XNOR2_X1 U11054 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10003) );
  NOR2_X1 U11055 ( .A1(n10004), .A2(n10003), .ZN(n10000) );
  NOR2_X1 U11056 ( .A1(n10001), .A2(n10000), .ZN(n10019) );
  NOR2_X1 U11057 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10019), .ZN(n10020) );
  AOI21_X1 U11058 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10019), .A(n10020), 
        .ZN(n10002) );
  XNOR2_X1 U11059 ( .A(n10002), .B(n10021), .ZN(ADD_1068_U55) );
  XNOR2_X1 U11060 ( .A(n10004), .B(n10003), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11061 ( .A(n10006), .B(n10005), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11062 ( .A(n10008), .B(n10007), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11063 ( .A(n10010), .B(n10009), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11064 ( .A(n10012), .B(n10011), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11065 ( .A(n10014), .B(n10013), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11066 ( .A(n10016), .B(n10015), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11067 ( .A(n10018), .B(n10017), .ZN(ADD_1068_U63) );
  NAND2_X1 U11068 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10019), .ZN(n10022) );
  AOI21_X1 U11069 ( .B1(n10022), .B2(n10021), .A(n10020), .ZN(n10024) );
  XNOR2_X1 U11070 ( .A(n4563), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n10023) );
  XNOR2_X1 U11071 ( .A(n10024), .B(n10023), .ZN(n10214) );
  AOI22_X1 U11072 ( .A1(n5120), .A2(keyinput_g50), .B1(keyinput_g54), .B2(
        n6667), .ZN(n10025) );
  OAI221_X1 U11073 ( .B1(n5120), .B2(keyinput_g50), .C1(n6667), .C2(
        keyinput_g54), .A(n10025), .ZN(n10034) );
  INV_X1 U11074 ( .A(SI_13_), .ZN(n10187) );
  AOI22_X1 U11075 ( .A1(n10027), .A2(keyinput_g60), .B1(keyinput_g19), .B2(
        n10187), .ZN(n10026) );
  OAI221_X1 U11076 ( .B1(n10027), .B2(keyinput_g60), .C1(n10187), .C2(
        keyinput_g19), .A(n10026), .ZN(n10033) );
  INV_X1 U11077 ( .A(SI_16_), .ZN(n10160) );
  AOI22_X1 U11078 ( .A1(n10160), .A2(keyinput_g16), .B1(n10149), .B2(
        keyinput_g6), .ZN(n10028) );
  OAI221_X1 U11079 ( .B1(n10160), .B2(keyinput_g16), .C1(n10149), .C2(
        keyinput_g6), .A(n10028), .ZN(n10032) );
  XNOR2_X1 U11080 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10030) );
  XNOR2_X1 U11081 ( .A(SI_5_), .B(keyinput_g27), .ZN(n10029) );
  NAND2_X1 U11082 ( .A1(n10030), .A2(n10029), .ZN(n10031) );
  NOR4_X1 U11083 ( .A1(n10034), .A2(n10033), .A3(n10032), .A4(n10031), .ZN(
        n10071) );
  INV_X1 U11084 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10142) );
  AOI22_X1 U11085 ( .A1(n5117), .A2(keyinput_g56), .B1(keyinput_g33), .B2(
        n10142), .ZN(n10035) );
  OAI221_X1 U11086 ( .B1(n5117), .B2(keyinput_g56), .C1(n10142), .C2(
        keyinput_g33), .A(n10035), .ZN(n10044) );
  AOI22_X1 U11087 ( .A1(SI_17_), .A2(keyinput_g15), .B1(
        P2_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .ZN(n10036) );
  OAI221_X1 U11088 ( .B1(SI_17_), .B2(keyinput_g15), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_g48), .A(n10036), .ZN(n10043)
         );
  INV_X1 U11089 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n10172) );
  AOI22_X1 U11090 ( .A1(n10172), .A2(keyinput_g42), .B1(keyinput_g22), .B2(
        n10038), .ZN(n10037) );
  OAI221_X1 U11091 ( .B1(n10172), .B2(keyinput_g42), .C1(n10038), .C2(
        keyinput_g22), .A(n10037), .ZN(n10042) );
  AOI22_X1 U11092 ( .A1(n10040), .A2(keyinput_g46), .B1(keyinput_g35), .B2(
        n10163), .ZN(n10039) );
  OAI221_X1 U11093 ( .B1(n10040), .B2(keyinput_g46), .C1(n10163), .C2(
        keyinput_g35), .A(n10039), .ZN(n10041) );
  NOR4_X1 U11094 ( .A1(n10044), .A2(n10043), .A3(n10042), .A4(n10041), .ZN(
        n10070) );
  AOI22_X1 U11095 ( .A1(P2_U3151), .A2(keyinput_g34), .B1(keyinput_g1), .B2(
        n7918), .ZN(n10045) );
  OAI221_X1 U11096 ( .B1(P2_U3151), .B2(keyinput_g34), .C1(n7918), .C2(
        keyinput_g1), .A(n10045), .ZN(n10056) );
  INV_X1 U11097 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10175) );
  INV_X1 U11098 ( .A(SI_21_), .ZN(n10047) );
  AOI22_X1 U11099 ( .A1(n10175), .A2(keyinput_g38), .B1(keyinput_g11), .B2(
        n10047), .ZN(n10046) );
  OAI221_X1 U11100 ( .B1(n10175), .B2(keyinput_g38), .C1(n10047), .C2(
        keyinput_g11), .A(n10046), .ZN(n10055) );
  AOI22_X1 U11101 ( .A1(n10050), .A2(keyinput_g18), .B1(n10049), .B2(
        keyinput_g43), .ZN(n10048) );
  OAI221_X1 U11102 ( .B1(n10050), .B2(keyinput_g18), .C1(n10049), .C2(
        keyinput_g43), .A(n10048), .ZN(n10054) );
  XNOR2_X1 U11103 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_g44), .ZN(n10052)
         );
  XNOR2_X1 U11104 ( .A(SI_18_), .B(keyinput_g14), .ZN(n10051) );
  NAND2_X1 U11105 ( .A1(n10052), .A2(n10051), .ZN(n10053) );
  NOR4_X1 U11106 ( .A1(n10056), .A2(n10055), .A3(n10054), .A4(n10053), .ZN(
        n10069) );
  AOI22_X1 U11107 ( .A1(n5124), .A2(keyinput_g45), .B1(keyinput_g8), .B2(
        n10058), .ZN(n10057) );
  OAI221_X1 U11108 ( .B1(n5124), .B2(keyinput_g45), .C1(n10058), .C2(
        keyinput_g8), .A(n10057), .ZN(n10067) );
  AOI22_X1 U11109 ( .A1(n10060), .A2(keyinput_g51), .B1(keyinput_g37), .B2(
        n10185), .ZN(n10059) );
  OAI221_X1 U11110 ( .B1(n10060), .B2(keyinput_g51), .C1(n10185), .C2(
        keyinput_g37), .A(n10059), .ZN(n10066) );
  AOI22_X1 U11111 ( .A1(n10062), .A2(keyinput_g39), .B1(keyinput_g61), .B2(
        n10165), .ZN(n10061) );
  OAI221_X1 U11112 ( .B1(n10062), .B2(keyinput_g39), .C1(n10165), .C2(
        keyinput_g61), .A(n10061), .ZN(n10065) );
  AOI22_X1 U11113 ( .A1(n10146), .A2(keyinput_g2), .B1(n5114), .B2(
        keyinput_g53), .ZN(n10063) );
  OAI221_X1 U11114 ( .B1(n10146), .B2(keyinput_g2), .C1(n5114), .C2(
        keyinput_g53), .A(n10063), .ZN(n10064) );
  NOR4_X1 U11115 ( .A1(n10067), .A2(n10066), .A3(n10065), .A4(n10064), .ZN(
        n10068) );
  NAND4_X1 U11116 ( .A1(n10071), .A2(n10070), .A3(n10069), .A4(n10068), .ZN(
        n10212) );
  AOI22_X1 U11117 ( .A1(SI_15_), .A2(keyinput_g17), .B1(SI_23_), .B2(
        keyinput_g9), .ZN(n10072) );
  OAI221_X1 U11118 ( .B1(SI_15_), .B2(keyinput_g17), .C1(SI_23_), .C2(
        keyinput_g9), .A(n10072), .ZN(n10079) );
  AOI22_X1 U11119 ( .A1(SI_22_), .A2(keyinput_g10), .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .ZN(n10073) );
  OAI221_X1 U11120 ( .B1(SI_22_), .B2(keyinput_g10), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_g40), .A(n10073), .ZN(n10078) );
  AOI22_X1 U11121 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_12_), .B2(keyinput_g20), .ZN(n10074) );
  OAI221_X1 U11122 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        SI_12_), .C2(keyinput_g20), .A(n10074), .ZN(n10077) );
  AOI22_X1 U11123 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n10075) );
  OAI221_X1 U11124 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_g36), .A(n10075), .ZN(n10076)
         );
  NOR4_X1 U11125 ( .A1(n10079), .A2(n10078), .A3(n10077), .A4(n10076), .ZN(
        n10106) );
  XNOR2_X1 U11126 ( .A(SI_7_), .B(keyinput_g25), .ZN(n10086) );
  AOI22_X1 U11127 ( .A1(SI_6_), .A2(keyinput_g26), .B1(n5127), .B2(
        keyinput_g47), .ZN(n10080) );
  OAI221_X1 U11128 ( .B1(SI_6_), .B2(keyinput_g26), .C1(n5127), .C2(
        keyinput_g47), .A(n10080), .ZN(n10085) );
  AOI22_X1 U11129 ( .A1(SI_4_), .A2(keyinput_g28), .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n10081) );
  OAI221_X1 U11130 ( .B1(SI_4_), .B2(keyinput_g28), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n10081), .ZN(n10084)
         );
  AOI22_X1 U11131 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_g55), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n10082) );
  OAI221_X1 U11132 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n10082), .ZN(n10083)
         );
  NOR4_X1 U11133 ( .A1(n10086), .A2(n10085), .A3(n10084), .A4(n10083), .ZN(
        n10105) );
  AOI22_X1 U11134 ( .A1(SI_2_), .A2(keyinput_g30), .B1(SI_20_), .B2(
        keyinput_g12), .ZN(n10087) );
  OAI221_X1 U11135 ( .B1(SI_2_), .B2(keyinput_g30), .C1(SI_20_), .C2(
        keyinput_g12), .A(n10087), .ZN(n10094) );
  AOI22_X1 U11136 ( .A1(SI_3_), .A2(keyinput_g29), .B1(SI_25_), .B2(
        keyinput_g7), .ZN(n10088) );
  OAI221_X1 U11137 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_25_), .C2(
        keyinput_g7), .A(n10088), .ZN(n10093) );
  AOI22_X1 U11138 ( .A1(SI_27_), .A2(keyinput_g5), .B1(SI_28_), .B2(
        keyinput_g4), .ZN(n10089) );
  OAI221_X1 U11139 ( .B1(SI_27_), .B2(keyinput_g5), .C1(SI_28_), .C2(
        keyinput_g4), .A(n10089), .ZN(n10092) );
  AOI22_X1 U11140 ( .A1(SI_0_), .A2(keyinput_g32), .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n10090) );
  OAI221_X1 U11141 ( .B1(SI_0_), .B2(keyinput_g32), .C1(
        P2_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n10090), .ZN(n10091)
         );
  NOR4_X1 U11142 ( .A1(n10094), .A2(n10093), .A3(n10092), .A4(n10091), .ZN(
        n10104) );
  AOI22_X1 U11143 ( .A1(SI_9_), .A2(keyinput_g23), .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n10095) );
  OAI221_X1 U11144 ( .B1(SI_9_), .B2(keyinput_g23), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n10095), .ZN(n10102)
         );
  AOI22_X1 U11145 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_g49), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n10096) );
  OAI221_X1 U11146 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n10096), .ZN(n10101)
         );
  AOI22_X1 U11147 ( .A1(SI_8_), .A2(keyinput_g24), .B1(P2_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_g52), .ZN(n10097) );
  OAI221_X1 U11148 ( .B1(SI_8_), .B2(keyinput_g24), .C1(P2_REG3_REG_4__SCAN_IN), .C2(keyinput_g52), .A(n10097), .ZN(n10100) );
  AOI22_X1 U11149 ( .A1(SI_19_), .A2(keyinput_g13), .B1(SI_29_), .B2(
        keyinput_g3), .ZN(n10098) );
  OAI221_X1 U11150 ( .B1(SI_19_), .B2(keyinput_g13), .C1(SI_29_), .C2(
        keyinput_g3), .A(n10098), .ZN(n10099) );
  NOR4_X1 U11151 ( .A1(n10102), .A2(n10101), .A3(n10100), .A4(n10099), .ZN(
        n10103) );
  NAND4_X1 U11152 ( .A1(n10106), .A2(n10105), .A3(n10104), .A4(n10103), .ZN(
        n10211) );
  INV_X1 U11153 ( .A(keyinput_f21), .ZN(n10204) );
  OAI22_X1 U11154 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        keyinput_f52), .B2(P2_REG3_REG_4__SCAN_IN), .ZN(n10107) );
  AOI221_X1 U11155 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        P2_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n10107), .ZN(n10124) );
  OAI22_X1 U11156 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        keyinput_f20), .B2(SI_12_), .ZN(n10108) );
  AOI221_X1 U11157 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        SI_12_), .C2(keyinput_f20), .A(n10108), .ZN(n10123) );
  AOI22_X1 U11158 ( .A1(SI_24_), .A2(keyinput_f8), .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_f48), .ZN(n10109) );
  OAI221_X1 U11159 ( .B1(SI_24_), .B2(keyinput_f8), .C1(
        P2_REG3_REG_16__SCAN_IN), .C2(keyinput_f48), .A(n10109), .ZN(n10116)
         );
  AOI22_X1 U11160 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_f59), .B1(SI_23_), .B2(keyinput_f9), .ZN(n10110) );
  OAI221_X1 U11161 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_f59), .C1(
        SI_23_), .C2(keyinput_f9), .A(n10110), .ZN(n10115) );
  AOI22_X1 U11162 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput_f53), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n10111) );
  OAI221_X1 U11163 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n10111), .ZN(n10114)
         );
  AOI22_X1 U11164 ( .A1(SI_1_), .A2(keyinput_f31), .B1(SI_25_), .B2(
        keyinput_f7), .ZN(n10112) );
  OAI221_X1 U11165 ( .B1(SI_1_), .B2(keyinput_f31), .C1(SI_25_), .C2(
        keyinput_f7), .A(n10112), .ZN(n10113) );
  NOR4_X1 U11166 ( .A1(n10116), .A2(n10115), .A3(n10114), .A4(n10113), .ZN(
        n10120) );
  OAI22_X1 U11167 ( .A1(n10118), .A2(keyinput_f17), .B1(keyinput_f10), .B2(
        SI_22_), .ZN(n10117) );
  AOI221_X1 U11168 ( .B1(n10118), .B2(keyinput_f17), .C1(SI_22_), .C2(
        keyinput_f10), .A(n10117), .ZN(n10119) );
  OAI211_X1 U11169 ( .C1(P2_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(
        n10120), .B(n10119), .ZN(n10121) );
  AOI21_X1 U11170 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .A(n10121), .ZN(n10122) );
  NAND3_X1 U11171 ( .A1(n10124), .A2(n10123), .A3(n10122), .ZN(n10203) );
  OAI22_X1 U11172 ( .A1(SI_10_), .A2(keyinput_f22), .B1(SI_31_), .B2(
        keyinput_f1), .ZN(n10125) );
  AOI221_X1 U11173 ( .B1(SI_10_), .B2(keyinput_f22), .C1(keyinput_f1), .C2(
        SI_31_), .A(n10125), .ZN(n10132) );
  OAI22_X1 U11174 ( .A1(SI_29_), .A2(keyinput_f3), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(keyinput_f54), .ZN(n10126) );
  AOI221_X1 U11175 ( .B1(SI_29_), .B2(keyinput_f3), .C1(keyinput_f54), .C2(
        P2_REG3_REG_0__SCAN_IN), .A(n10126), .ZN(n10131) );
  OAI22_X1 U11176 ( .A1(SI_19_), .A2(keyinput_f13), .B1(keyinput_f15), .B2(
        SI_17_), .ZN(n10127) );
  AOI221_X1 U11177 ( .B1(SI_19_), .B2(keyinput_f13), .C1(SI_17_), .C2(
        keyinput_f15), .A(n10127), .ZN(n10130) );
  OAI22_X1 U11178 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_f50), .B1(
        keyinput_f4), .B2(SI_28_), .ZN(n10128) );
  AOI221_X1 U11179 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .C1(
        SI_28_), .C2(keyinput_f4), .A(n10128), .ZN(n10129) );
  NAND4_X1 U11180 ( .A1(n10132), .A2(n10131), .A3(n10130), .A4(n10129), .ZN(
        n10202) );
  OAI22_X1 U11181 ( .A1(SI_21_), .A2(keyinput_f11), .B1(SI_6_), .B2(
        keyinput_f26), .ZN(n10133) );
  AOI221_X1 U11182 ( .B1(SI_21_), .B2(keyinput_f11), .C1(keyinput_f26), .C2(
        SI_6_), .A(n10133), .ZN(n10140) );
  OAI22_X1 U11183 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(
        P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n10134) );
  AOI221_X1 U11184 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        keyinput_f55), .C2(P2_REG3_REG_20__SCAN_IN), .A(n10134), .ZN(n10139)
         );
  OAI22_X1 U11185 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_f49), .B1(SI_8_), 
        .B2(keyinput_f24), .ZN(n10135) );
  AOI221_X1 U11186 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .C1(
        keyinput_f24), .C2(SI_8_), .A(n10135), .ZN(n10138) );
  OAI22_X1 U11187 ( .A1(P2_STATE_REG_SCAN_IN), .A2(keyinput_f34), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n10136) );
  AOI221_X1 U11188 ( .B1(P2_STATE_REG_SCAN_IN), .B2(keyinput_f34), .C1(
        keyinput_f46), .C2(P2_REG3_REG_12__SCAN_IN), .A(n10136), .ZN(n10137)
         );
  NAND4_X1 U11189 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10201) );
  INV_X1 U11190 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10143) );
  AOI22_X1 U11191 ( .A1(n10143), .A2(keyinput_f57), .B1(keyinput_f33), .B2(
        n10142), .ZN(n10141) );
  OAI221_X1 U11192 ( .B1(n10143), .B2(keyinput_f57), .C1(n10142), .C2(
        keyinput_f33), .A(n10141), .ZN(n10155) );
  INV_X1 U11193 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10145) );
  AOI22_X1 U11194 ( .A1(n10146), .A2(keyinput_f2), .B1(keyinput_f0), .B2(
        n10145), .ZN(n10144) );
  OAI221_X1 U11195 ( .B1(n10146), .B2(keyinput_f2), .C1(n10145), .C2(
        keyinput_f0), .A(n10144), .ZN(n10154) );
  AOI22_X1 U11196 ( .A1(n10149), .A2(keyinput_f6), .B1(keyinput_f12), .B2(
        n10148), .ZN(n10147) );
  OAI221_X1 U11197 ( .B1(n10149), .B2(keyinput_f6), .C1(n10148), .C2(
        keyinput_f12), .A(n10147), .ZN(n10153) );
  XNOR2_X1 U11198 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_f43), .ZN(n10151)
         );
  XNOR2_X1 U11199 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_f40), .ZN(n10150)
         );
  NAND2_X1 U11200 ( .A1(n10151), .A2(n10150), .ZN(n10152) );
  NOR4_X1 U11201 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n10199) );
  AOI22_X1 U11202 ( .A1(n10158), .A2(keyinput_f63), .B1(keyinput_f58), .B2(
        n10157), .ZN(n10156) );
  OAI221_X1 U11203 ( .B1(n10158), .B2(keyinput_f63), .C1(n10157), .C2(
        keyinput_f58), .A(n10156), .ZN(n10170) );
  AOI22_X1 U11204 ( .A1(SI_4_), .A2(keyinput_f28), .B1(n10160), .B2(
        keyinput_f16), .ZN(n10159) );
  OAI221_X1 U11205 ( .B1(SI_4_), .B2(keyinput_f28), .C1(n10160), .C2(
        keyinput_f16), .A(n10159), .ZN(n10169) );
  AOI22_X1 U11206 ( .A1(n10163), .A2(keyinput_f35), .B1(keyinput_f14), .B2(
        n10162), .ZN(n10161) );
  OAI221_X1 U11207 ( .B1(n10163), .B2(keyinput_f35), .C1(n10162), .C2(
        keyinput_f14), .A(n10161), .ZN(n10168) );
  AOI22_X1 U11208 ( .A1(n10166), .A2(keyinput_f5), .B1(n10165), .B2(
        keyinput_f61), .ZN(n10164) );
  OAI221_X1 U11209 ( .B1(n10166), .B2(keyinput_f5), .C1(n10165), .C2(
        keyinput_f61), .A(n10164), .ZN(n10167) );
  NOR4_X1 U11210 ( .A1(n10170), .A2(n10169), .A3(n10168), .A4(n10167), .ZN(
        n10198) );
  AOI22_X1 U11211 ( .A1(n5117), .A2(keyinput_f56), .B1(n10172), .B2(
        keyinput_f42), .ZN(n10171) );
  OAI221_X1 U11212 ( .B1(n5117), .B2(keyinput_f56), .C1(n10172), .C2(
        keyinput_f42), .A(n10171), .ZN(n10182) );
  INV_X1 U11213 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U11214 ( .A1(n10174), .A2(keyinput_f62), .B1(n5521), .B2(
        keyinput_f36), .ZN(n10173) );
  OAI221_X1 U11215 ( .B1(n10174), .B2(keyinput_f62), .C1(n5521), .C2(
        keyinput_f36), .A(n10173), .ZN(n10181) );
  XOR2_X1 U11216 ( .A(n10175), .B(keyinput_f38), .Z(n10179) );
  XNOR2_X1 U11217 ( .A(SI_5_), .B(keyinput_f27), .ZN(n10178) );
  XNOR2_X1 U11218 ( .A(SI_2_), .B(keyinput_f30), .ZN(n10177) );
  XNOR2_X1 U11219 ( .A(SI_3_), .B(keyinput_f29), .ZN(n10176) );
  NAND4_X1 U11220 ( .A1(n10179), .A2(n10178), .A3(n10177), .A4(n10176), .ZN(
        n10180) );
  NOR3_X1 U11221 ( .A1(n10182), .A2(n10181), .A3(n10180), .ZN(n10197) );
  AOI22_X1 U11222 ( .A1(n10185), .A2(keyinput_f37), .B1(keyinput_f25), .B2(
        n10184), .ZN(n10183) );
  OAI221_X1 U11223 ( .B1(n10185), .B2(keyinput_f37), .C1(n10184), .C2(
        keyinput_f25), .A(n10183), .ZN(n10195) );
  AOI22_X1 U11224 ( .A1(n10188), .A2(keyinput_f23), .B1(n10187), .B2(
        keyinput_f19), .ZN(n10186) );
  OAI221_X1 U11225 ( .B1(n10188), .B2(keyinput_f23), .C1(n10187), .C2(
        keyinput_f19), .A(n10186), .ZN(n10194) );
  XNOR2_X1 U11226 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_f39), .ZN(n10192)
         );
  XNOR2_X1 U11227 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_f44), .ZN(n10191)
         );
  XNOR2_X1 U11228 ( .A(SI_0_), .B(keyinput_f32), .ZN(n10190) );
  XNOR2_X1 U11229 ( .A(SI_14_), .B(keyinput_f18), .ZN(n10189) );
  NAND4_X1 U11230 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10193) );
  NOR3_X1 U11231 ( .A1(n10195), .A2(n10194), .A3(n10193), .ZN(n10196) );
  NAND4_X1 U11232 ( .A1(n10199), .A2(n10198), .A3(n10197), .A4(n10196), .ZN(
        n10200) );
  NOR4_X1 U11233 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10207) );
  OAI211_X1 U11234 ( .C1(n10204), .C2(n10207), .A(SI_11_), .B(keyinput_g21), 
        .ZN(n10209) );
  INV_X1 U11235 ( .A(keyinput_g21), .ZN(n10205) );
  OAI211_X1 U11236 ( .C1(n10207), .C2(keyinput_f21), .A(n10206), .B(n10205), 
        .ZN(n10208) );
  NAND2_X1 U11237 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  OAI21_X1 U11238 ( .B1(n10212), .B2(n10211), .A(n10210), .ZN(n10213) );
  XOR2_X1 U11239 ( .A(n10214), .B(n10213), .Z(ADD_1068_U4) );
  XOR2_X1 U11240 ( .A(n10216), .B(n10215), .Z(ADD_1068_U54) );
  XNOR2_X1 U11241 ( .A(n10218), .B(n10217), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11242 ( .A(n10220), .B(n10219), .ZN(ADD_1068_U48) );
  XNOR2_X1 U11243 ( .A(n10222), .B(n10221), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11244 ( .A(n10224), .B(n10223), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11245 ( .A(n10226), .B(n10225), .ZN(ADD_1068_U51) );
  XOR2_X1 U11246 ( .A(n10228), .B(n10227), .Z(ADD_1068_U53) );
  XNOR2_X1 U11247 ( .A(n10230), .B(n10229), .ZN(ADD_1068_U52) );
  INV_X2 U4865 ( .A(n8545), .ZN(n8554) );
  CLKBUF_X2 U4868 ( .A(n5726), .Z(n4355) );
  CLKBUF_X1 U4879 ( .A(n5011), .Z(n7917) );
endmodule

