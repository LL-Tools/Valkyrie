

module b22_C_AntiSAT_k_128_10 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293;

  AND2_X1 U7207 ( .A1(n7135), .A2(n9223), .ZN(n6567) );
  NAND2_X1 U7208 ( .A1(n7638), .A2(n7637), .ZN(n13314) );
  NAND2_X1 U7209 ( .A1(n8178), .A2(n8177), .ZN(n13327) );
  NAND2_X1 U7210 ( .A1(n8482), .A2(n8481), .ZN(n11820) );
  CLKBUF_X2 U7211 ( .A(n10153), .Z(n13555) );
  INV_X1 U7212 ( .A(n8210), .ZN(n8201) );
  CLKBUF_X2 U7213 ( .A(n10153), .Z(n6460) );
  INV_X2 U7214 ( .A(n13625), .ZN(n13561) );
  INV_X2 U7215 ( .A(n9499), .ZN(n10389) );
  BUF_X1 U7216 ( .A(n7773), .Z(n12785) );
  CLKBUF_X2 U7217 ( .A(n9000), .Z(n9306) );
  INV_X1 U7218 ( .A(n13780), .ZN(n10164) );
  INV_X1 U7219 ( .A(n8829), .ZN(n7333) );
  AND2_X1 U7220 ( .A1(n7694), .A2(n11929), .ZN(n7773) );
  AND2_X1 U7221 ( .A1(n8251), .A2(n8255), .ZN(n8294) );
  NAND2_X2 U7222 ( .A1(n7632), .A2(n7631), .ZN(n13454) );
  NAND2_X1 U7223 ( .A1(n6823), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6687) );
  NAND2_X2 U7224 ( .A1(n10006), .A2(n10190), .ZN(n14650) );
  OR2_X1 U7225 ( .A1(n13267), .A2(n13251), .ZN(n13249) );
  OAI21_X1 U7226 ( .B1(n11391), .B2(n7143), .A(n7142), .ZN(n11704) );
  NAND2_X2 U7227 ( .A1(n11454), .A2(n10011), .ZN(n10019) );
  NAND2_X1 U7228 ( .A1(n7569), .A2(n7568), .ZN(n7570) );
  CLKBUF_X2 U7229 ( .A(n8823), .Z(n9134) );
  AND2_X1 U7230 ( .A1(n11884), .A2(n8774), .ZN(n8824) );
  AND2_X1 U7231 ( .A1(n9337), .A2(n9479), .ZN(n9745) );
  NAND2_X1 U7232 ( .A1(n7114), .A2(n7112), .ZN(n12516) );
  AND3_X1 U7233 ( .A1(n8816), .A2(n8815), .A3(n8814), .ZN(n15031) );
  NAND2_X1 U7234 ( .A1(n8721), .A2(n8720), .ZN(n8722) );
  NAND2_X1 U7235 ( .A1(n13454), .A2(n10058), .ZN(n10053) );
  CLKBUF_X2 U7236 ( .A(n7744), .Z(n8210) );
  AND2_X1 U7237 ( .A1(n10052), .A2(n10059), .ZN(n13036) );
  OR2_X1 U7238 ( .A1(n7669), .A2(n7805), .ZN(n7673) );
  NAND2_X1 U7239 ( .A1(n13708), .A2(n13709), .ZN(n13707) );
  OAI21_X1 U7240 ( .B1(n11820), .B2(n9682), .A(n9683), .ZN(n14033) );
  OAI21_X1 U7241 ( .B1(n8628), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7286) );
  OAI22_X1 U7242 ( .A1(n14177), .A2(n14178), .B1(P1_ADDR_REG_1__SCAN_IN), .B2(
        n14179), .ZN(n14237) );
  AND3_X1 U7243 ( .A1(n8869), .A2(n8868), .A3(n8867), .ZN(n14994) );
  AND2_X1 U7244 ( .A1(n7064), .A2(n7060), .ZN(n12289) );
  NAND2_X1 U7245 ( .A1(n8764), .A2(n8763), .ZN(n11963) );
  XNOR2_X1 U7246 ( .A(n9174), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11033) );
  OAI21_X1 U7247 ( .B1(P1_DATAO_REG_18__SCAN_IN), .B2(n10777), .A(n8731), .ZN(
        n9073) );
  XNOR2_X1 U7248 ( .A(n8722), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8985) );
  INV_X1 U7249 ( .A(n12886), .ZN(n13435) );
  OR2_X1 U7250 ( .A1(n14059), .A2(n14016), .ZN(n7517) );
  NAND2_X1 U7251 ( .A1(n8444), .A2(n8443), .ZN(n14414) );
  INV_X1 U7252 ( .A(n9926), .ZN(n9925) );
  NAND2_X1 U7253 ( .A1(n8773), .A2(n12644), .ZN(n11879) );
  AOI211_X1 U7254 ( .C1(n13327), .C2(n14381), .A(n12686), .B(n12685), .ZN(
        n12687) );
  CLKBUF_X3 U7255 ( .A(n10028), .Z(n14629) );
  XOR2_X1 U7256 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n14233), .Z(n15292) );
  INV_X1 U7257 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8841) );
  NOR2_X2 U7258 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6472) );
  OAI21_X2 U7259 ( .B1(n8838), .B2(n8705), .A(n8704), .ZN(n8853) );
  NOR2_X2 U7260 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), .ZN(
        n8752) );
  XNOR2_X1 U7261 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8810) );
  NAND2_X4 U7262 ( .A1(n6895), .A2(n6766), .ZN(n7522) );
  INV_X2 U7263 ( .A(n7522), .ZN(n7524) );
  XNOR2_X2 U7264 ( .A(n6635), .B(n12836), .ZN(n10765) );
  OR2_X2 U7265 ( .A1(n11807), .A2(n11806), .ZN(n6628) );
  NAND2_X2 U7266 ( .A1(n7685), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7677) );
  INV_X2 U7267 ( .A(n11983), .ZN(n13068) );
  XNOR2_X2 U7268 ( .A(n10890), .B(n10888), .ZN(n10887) );
  NAND2_X2 U7269 ( .A1(n10868), .A2(n10867), .ZN(n10890) );
  AOI211_X2 U7270 ( .C1(n13031), .C2(n13030), .A(n13029), .B(n13028), .ZN(
        n13032) );
  AOI21_X2 U7271 ( .B1(n6744), .B2(n12977), .A(n12976), .ZN(n13031) );
  INV_X2 U7272 ( .A(n11417), .ZN(n7734) );
  NOR2_X2 U7273 ( .A1(n14276), .A2(n14275), .ZN(n14479) );
  XNOR2_X1 U7275 ( .A(n7286), .B(n8239), .ZN(n14489) );
  NOR2_X2 U7276 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n7680) );
  NOR2_X4 U7277 ( .A1(n8286), .A2(n6725), .ZN(n13788) );
  OAI21_X4 U7278 ( .B1(n13743), .B2(n13744), .A(n13509), .ZN(n13662) );
  NAND2_X2 U7279 ( .A1(n7073), .A2(n8813), .ZN(n10456) );
  AOI21_X2 U7280 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n11077), .A(n14931), .ZN(
        n11226) );
  OAI21_X2 U7281 ( .B1(n14272), .B2(n14271), .A(n14468), .ZN(n14473) );
  AOI211_X1 U7282 ( .C1(n13314), .C2(n14381), .A(n8218), .B(n8217), .ZN(n8224)
         );
  NAND2_X1 U7283 ( .A1(n7195), .A2(n7192), .ZN(n14078) );
  NAND2_X1 U7284 ( .A1(n7733), .A2(n7732), .ZN(n13322) );
  NAND2_X1 U7285 ( .A1(n6465), .A2(n6462), .ZN(n10963) );
  INV_X2 U7286 ( .A(n14987), .ZN(n14969) );
  BUF_X2 U7287 ( .A(n9134), .Z(n9231) );
  CLKBUF_X3 U7288 ( .A(n8824), .Z(n8893) );
  NAND4_X1 U7289 ( .A1(n8327), .A2(n8326), .A3(n8325), .A4(n8324), .ZN(n13777)
         );
  INV_X8 U7290 ( .A(n12852), .ZN(n6461) );
  INV_X1 U7291 ( .A(n10264), .ZN(n14659) );
  AND3_X1 U7292 ( .A1(n7035), .A2(n7743), .A3(n7034), .ZN(n10355) );
  NAND2_X1 U7293 ( .A1(n7761), .A2(n6650), .ZN(n12824) );
  INV_X1 U7295 ( .A(n9499), .ZN(n6717) );
  NAND2_X1 U7296 ( .A1(n12784), .A2(n6742), .ZN(n12814) );
  CLKBUF_X2 U7297 ( .A(n7735), .Z(n6742) );
  CLKBUF_X2 U7298 ( .A(n8279), .Z(n8550) );
  NOR2_X1 U7299 ( .A1(n11033), .A2(n9230), .ZN(n15023) );
  NOR2_X4 U7300 ( .A1(n11515), .A2(n7734), .ZN(n7737) );
  AND2_X1 U7301 ( .A1(n8546), .A2(n9925), .ZN(n8290) );
  INV_X1 U7302 ( .A(n14155), .ZN(n8251) );
  CLKBUF_X2 U7303 ( .A(n8264), .Z(n14159) );
  NAND2_X1 U7304 ( .A1(n7675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7671) );
  NAND2_X1 U7305 ( .A1(n7675), .A2(n7674), .ZN(n11515) );
  NAND2_X1 U7306 ( .A1(n7673), .A2(n7672), .ZN(n7675) );
  OR2_X1 U7307 ( .A1(n7673), .A2(n7672), .ZN(n7674) );
  INV_X8 U7308 ( .A(n7522), .ZN(n9926) );
  INV_X2 U7309 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n8241) );
  OAI21_X1 U7310 ( .B1(n7266), .B2(n7184), .A(n14724), .ZN(n7183) );
  AOI211_X1 U7311 ( .C1(n14065), .C2(n14644), .A(n13909), .B(n13908), .ZN(
        n13910) );
  AND2_X1 U7312 ( .A1(n13316), .A2(n6753), .ZN(n13399) );
  OR2_X1 U7313 ( .A1(n12354), .A2(n9472), .ZN(n7135) );
  AND2_X1 U7314 ( .A1(n6755), .A2(n6754), .ZN(n13316) );
  NAND2_X1 U7315 ( .A1(n6631), .A2(n9344), .ZN(n12354) );
  NAND2_X1 U7316 ( .A1(n13100), .A2(n11900), .ZN(n11903) );
  AND2_X1 U7317 ( .A1(n13914), .A2(n6955), .ZN(n13869) );
  NOR2_X1 U7318 ( .A1(n13090), .A2(n13089), .ZN(n13300) );
  NAND2_X1 U7319 ( .A1(n12382), .A2(n9348), .ZN(n12369) );
  AOI22_X1 U7320 ( .A1(n7470), .A2(n7473), .B1(n6510), .B2(n7477), .ZN(n7469)
         );
  NAND2_X1 U7321 ( .A1(n12395), .A2(n6533), .ZN(n12382) );
  NAND2_X1 U7322 ( .A1(n13157), .A2(n11898), .ZN(n13143) );
  NOR2_X1 U7323 ( .A1(n8688), .A2(n6484), .ZN(n6829) );
  NAND2_X1 U7324 ( .A1(n9297), .A2(n9296), .ZN(n9315) );
  AOI21_X2 U7325 ( .B1(n12783), .B2(n12782), .A(n7515), .ZN(n13022) );
  AND2_X1 U7326 ( .A1(n9655), .A2(n9671), .ZN(n12783) );
  OAI22_X1 U7327 ( .A1(n9303), .A2(n9292), .B1(P2_DATAO_REG_30__SCAN_IN), .B2(
        n11928), .ZN(n6722) );
  OR2_X1 U7328 ( .A1(n12308), .A2(n12307), .ZN(n12326) );
  INV_X1 U7329 ( .A(n7158), .ZN(n6466) );
  NAND2_X1 U7330 ( .A1(n13982), .A2(n8544), .ZN(n13973) );
  NAND2_X1 U7331 ( .A1(n13222), .A2(n11893), .ZN(n13206) );
  NOR2_X1 U7332 ( .A1(n11899), .A2(n7157), .ZN(n7156) );
  NAND2_X1 U7333 ( .A1(n13211), .A2(n6531), .ZN(n13147) );
  NAND2_X1 U7334 ( .A1(n6471), .A2(n13220), .ZN(n13222) );
  AND2_X1 U7335 ( .A1(n13927), .A2(n6521), .ZN(n7192) );
  NAND2_X1 U7336 ( .A1(n8246), .A2(n8245), .ZN(n14066) );
  OR2_X1 U7337 ( .A1(n12523), .A2(n12353), .ZN(n9473) );
  AND2_X2 U7338 ( .A1(n8200), .A2(n8199), .ZN(n13402) );
  AND2_X1 U7339 ( .A1(n9223), .A2(n9222), .ZN(n12355) );
  NAND2_X1 U7340 ( .A1(n8783), .A2(n8782), .ZN(n12523) );
  NAND2_X1 U7341 ( .A1(n6632), .A2(n9070), .ZN(n12454) );
  INV_X1 U7342 ( .A(n12946), .ZN(n13408) );
  INV_X1 U7343 ( .A(n12456), .ZN(n6632) );
  NAND2_X1 U7344 ( .A1(n7109), .A2(n7108), .ZN(n12456) );
  OAI21_X1 U7345 ( .B1(n13260), .B2(n11890), .A(n11891), .ZN(n13241) );
  NAND2_X1 U7346 ( .A1(n8585), .A2(n8584), .ZN(n13915) );
  NAND2_X1 U7347 ( .A1(n7101), .A2(n6898), .ZN(n13178) );
  NAND2_X1 U7348 ( .A1(n6464), .A2(n12913), .ZN(n13260) );
  NOR2_X1 U7349 ( .A1(n8742), .A2(n7319), .ZN(n8781) );
  AND2_X1 U7350 ( .A1(n8162), .A2(n8161), .ZN(n11844) );
  NOR2_X1 U7351 ( .A1(n14285), .A2(n14284), .ZN(n14484) );
  NAND2_X1 U7352 ( .A1(n13278), .A2(n12912), .ZN(n6464) );
  AND2_X1 U7353 ( .A1(n9131), .A2(n9130), .ZN(n12602) );
  NOR2_X1 U7354 ( .A1(n7273), .A2(n6538), .ZN(n7272) );
  NAND2_X1 U7355 ( .A1(n8147), .A2(n8146), .ZN(n13182) );
  NAND2_X1 U7356 ( .A1(n11749), .A2(n8467), .ZN(n11776) );
  OAI21_X1 U7357 ( .B1(n8158), .B2(n6609), .A(n6705), .ZN(n7729) );
  AND2_X1 U7358 ( .A1(n8009), .A2(n8022), .ZN(n6929) );
  NAND2_X1 U7359 ( .A1(n11889), .A2(n11888), .ZN(n13278) );
  AOI21_X1 U7360 ( .B1(n11704), .B2(n11703), .A(n11705), .ZN(n6476) );
  OAI21_X1 U7361 ( .B1(n12516), .B2(n9206), .A(n9422), .ZN(n11807) );
  NAND2_X1 U7362 ( .A1(n8533), .A2(n8532), .ZN(n14108) );
  NAND2_X1 U7363 ( .A1(n11389), .A2(n11388), .ZN(n11391) );
  NAND2_X1 U7364 ( .A1(n14546), .A2(n14545), .ZN(n14544) );
  OR2_X1 U7365 ( .A1(n11993), .A2(n8131), .ZN(n6897) );
  NAND2_X1 U7366 ( .A1(n7016), .A2(n7015), .ZN(n14274) );
  NAND2_X1 U7367 ( .A1(n8523), .A2(n8522), .ZN(n14113) );
  NOR2_X1 U7368 ( .A1(n14391), .A2(n7393), .ZN(n7392) );
  NAND2_X1 U7369 ( .A1(n7374), .A2(n7373), .ZN(n11632) );
  AOI21_X1 U7370 ( .B1(n11570), .B2(n11569), .A(n11568), .ZN(n11653) );
  OAI22_X1 U7371 ( .A1(n9412), .A2(n9411), .B1(n10389), .B2(n9410), .ZN(n9416)
         );
  NAND2_X1 U7372 ( .A1(n6623), .A2(n8926), .ZN(n11455) );
  AND2_X1 U7373 ( .A1(n7440), .A2(n8106), .ZN(n8087) );
  AOI21_X1 U7374 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14206), .A(n14205), .ZN(
        n14221) );
  NAND2_X1 U7375 ( .A1(n6568), .A2(n7367), .ZN(n13717) );
  AND2_X1 U7376 ( .A1(n12886), .A2(n13056), .ZN(n11705) );
  AND2_X1 U7377 ( .A1(n7981), .A2(n7980), .ZN(n12892) );
  NAND2_X1 U7378 ( .A1(n10963), .A2(n10962), .ZN(n11286) );
  OAI22_X1 U7379 ( .A1(n7570), .A2(n6701), .B1(n10421), .B2(n8045), .ZN(n8069)
         );
  OAI22_X1 U7380 ( .A1(n12838), .A2(n6900), .B1(n12839), .B2(n6899), .ZN(
        n12844) );
  XNOR2_X1 U7381 ( .A(n14264), .B(n14265), .ZN(n14296) );
  NAND2_X1 U7382 ( .A1(n8025), .A2(n8026), .ZN(n7569) );
  NAND2_X1 U7383 ( .A1(n7925), .A2(n7924), .ZN(n12875) );
  NAND2_X1 U7384 ( .A1(n14262), .A2(n14263), .ZN(n14264) );
  NAND2_X1 U7385 ( .A1(n8401), .A2(n8400), .ZN(n14453) );
  NOR2_X2 U7386 ( .A1(n10939), .A2(n14705), .ZN(n11001) );
  NAND2_X1 U7387 ( .A1(n8388), .A2(n8387), .ZN(n11381) );
  NAND2_X1 U7388 ( .A1(n7908), .A2(n7907), .ZN(n14892) );
  AND2_X1 U7389 ( .A1(n9391), .A2(n9389), .ZN(n11089) );
  INV_X1 U7390 ( .A(n12998), .ZN(n6462) );
  INV_X2 U7391 ( .A(n13248), .ZN(n13298) );
  NAND2_X1 U7392 ( .A1(n13248), .A2(n10570), .ZN(n13293) );
  AND2_X2 U7393 ( .A1(n13248), .A2(n13026), .ZN(n13288) );
  AND2_X1 U7394 ( .A1(n9377), .A2(n9378), .ZN(n15004) );
  INV_X2 U7395 ( .A(n15050), .ZN(n14334) );
  OAI211_X1 U7396 ( .C1(n7839), .C2(n6704), .A(n7547), .B(n6703), .ZN(n7451)
         );
  NOR2_X1 U7397 ( .A1(n7751), .A2(n11940), .ZN(n6743) );
  NAND3_X1 U7398 ( .A1(n7051), .A2(n7052), .A3(n6486), .ZN(n10629) );
  NAND4_X1 U7399 ( .A1(n8828), .A2(n8827), .A3(n8826), .A4(n8825), .ZN(n15033)
         );
  BUF_X2 U7400 ( .A(n8893), .Z(n6463) );
  OR2_X1 U7401 ( .A1(n9309), .A2(n8832), .ZN(n8833) );
  AND3_X1 U7402 ( .A1(n8861), .A2(n8860), .A3(n8859), .ZN(n14999) );
  NAND2_X2 U7403 ( .A1(n6779), .A2(n7336), .ZN(n10315) );
  INV_X1 U7404 ( .A(n14917), .ZN(n10311) );
  NAND2_X1 U7405 ( .A1(n8824), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8805) );
  NAND2_X1 U7406 ( .A1(n7539), .A2(n7538), .ZN(n7823) );
  INV_X4 U7407 ( .A(n13231), .ZN(n13106) );
  XNOR2_X1 U7408 ( .A(n13069), .B(n12824), .ZN(n12992) );
  XNOR2_X1 U7409 ( .A(n10355), .B(n7147), .ZN(n12991) );
  INV_X2 U7410 ( .A(n12814), .ZN(n12852) );
  AND4_X1 U7411 ( .A1(n8300), .A2(n8299), .A3(n8298), .A4(n8297), .ZN(n10847)
         );
  AND2_X1 U7412 ( .A1(n7084), .A2(n6572), .ZN(n11983) );
  AND2_X1 U7413 ( .A1(n7772), .A2(n7082), .ZN(n10566) );
  AOI21_X1 U7414 ( .B1(n13823), .B2(P1_REG1_REG_4__SCAN_IN), .A(n13821), .ZN(
        n9990) );
  INV_X1 U7415 ( .A(n13067), .ZN(n6635) );
  CLKBUF_X3 U7416 ( .A(n8294), .Z(n8606) );
  NAND4_X2 U7417 ( .A1(n7750), .A2(n7749), .A3(n7747), .A4(n7748), .ZN(n13072)
         );
  MUX2_X1 U7418 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8771), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8773) );
  INV_X2 U7419 ( .A(n8546), .ZN(n9921) );
  NAND2_X1 U7420 ( .A1(n7745), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U7421 ( .A1(n8770), .A2(n8761), .ZN(n11876) );
  MUX2_X1 U7422 ( .A(n13784), .B(n14175), .S(n8546), .Z(n14628) );
  NAND2_X2 U7423 ( .A1(n8264), .A2(n14489), .ZN(n8546) );
  NAND2_X1 U7424 ( .A1(n8623), .A2(n8622), .ZN(n11454) );
  NAND2_X1 U7425 ( .A1(n8250), .A2(n6823), .ZN(n14155) );
  NAND2_X1 U7426 ( .A1(n8204), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7427 ( .A1(n8247), .A2(n8244), .ZN(n8264) );
  MUX2_X1 U7428 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8249), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8250) );
  NAND2_X1 U7429 ( .A1(n7635), .A2(n7636), .ZN(n10058) );
  XNOR2_X1 U7430 ( .A(n8510), .B(n8509), .ZN(n13858) );
  MUX2_X1 U7431 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7634), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n7635) );
  XNOR2_X1 U7432 ( .A(n6653), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7693) );
  INV_X1 U7433 ( .A(n13449), .ZN(n7694) );
  XNOR2_X1 U7434 ( .A(n6470), .B(n6469), .ZN(n13449) );
  NAND2_X1 U7435 ( .A1(n7032), .A2(n7030), .ZN(n14181) );
  AND2_X1 U7436 ( .A1(n8858), .A2(n8889), .ZN(n10724) );
  XNOR2_X1 U7437 ( .A(n7537), .B(SI_5_), .ZN(n7803) );
  AND2_X1 U7438 ( .A1(n6646), .A2(n6918), .ZN(n7669) );
  NAND2_X1 U7439 ( .A1(n6644), .A2(n6918), .ZN(n7685) );
  OR2_X1 U7440 ( .A1(n7692), .A2(n7805), .ZN(n6470) );
  XNOR2_X1 U7441 ( .A(n8794), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10416) );
  NAND2_X1 U7442 ( .A1(n8813), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8794) );
  NOR2_X1 U7443 ( .A1(n7629), .A2(n7625), .ZN(n7202) );
  NOR2_X1 U7444 ( .A1(n7784), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7786) );
  AND2_X1 U7445 ( .A1(n8267), .A2(n8227), .ZN(n8314) );
  AND4_X1 U7446 ( .A1(n6667), .A2(n8226), .A3(n8332), .A4(n8313), .ZN(n6666)
         );
  AND2_X1 U7447 ( .A1(n6998), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14231) );
  AND2_X1 U7448 ( .A1(n8818), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8809) );
  NOR2_X1 U7449 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6667) );
  INV_X1 U7450 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9057) );
  INV_X4 U7451 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X4 U7452 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7453 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6998) );
  INV_X1 U7454 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8470) );
  NOR2_X1 U7455 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6474) );
  NOR2_X1 U7456 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n6473) );
  INV_X1 U7457 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9256) );
  INV_X1 U7458 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n8811) );
  INV_X1 U7459 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n9170) );
  INV_X1 U7460 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6469) );
  NOR2_X1 U7461 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n7622) );
  INV_X1 U7462 ( .A(n10599), .ZN(n6465) );
  OAI21_X1 U7463 ( .B1(n10597), .B2(n10596), .A(n10598), .ZN(n10599) );
  NAND2_X1 U7464 ( .A1(n10581), .A2(n10580), .ZN(n10597) );
  INV_X1 U7465 ( .A(n13120), .ZN(n7155) );
  NAND3_X1 U7466 ( .A1(n7153), .A2(n7161), .A3(n6503), .ZN(n13100) );
  NAND2_X1 U7467 ( .A1(n6466), .A2(n13120), .ZN(n6503) );
  NAND2_X1 U7468 ( .A1(n13143), .A2(n6573), .ZN(n7153) );
  INV_X2 U7469 ( .A(n7147), .ZN(n13070) );
  AND4_X2 U7470 ( .A1(n7738), .A2(n6468), .A3(n7739), .A4(n6467), .ZN(n7147)
         );
  AND4_X2 U7471 ( .A1(n7201), .A2(n7202), .A3(n6647), .A4(n7204), .ZN(n7692)
         );
  AOI21_X2 U7472 ( .B1(n13206), .B2(n11895), .A(n11894), .ZN(n13200) );
  NAND2_X1 U7473 ( .A1(n13240), .A2(n13243), .ZN(n6471) );
  NAND4_X1 U7474 ( .A1(n6474), .A2(n6473), .A3(n6472), .A4(n6654), .ZN(n7938)
         );
  AOI21_X2 U7475 ( .B1(n13608), .B2(n13680), .A(n13577), .ZN(n13684) );
  OAI22_X2 U7476 ( .A1(n8961), .A2(n8719), .B1(P2_DATAO_REG_11__SCAN_IN), .B2(
        n10037), .ZN(n8970) );
  OAI22_X2 U7477 ( .A1(n14033), .A2(n8505), .B1(n14130), .B2(n13765), .ZN(
        n14020) );
  NAND2_X2 U7478 ( .A1(n8164), .A2(n8163), .ZN(n12946) );
  NOR2_X2 U7479 ( .A1(n12223), .A2(n12224), .ZN(n12246) );
  NAND2_X2 U7480 ( .A1(n10335), .A2(n12984), .ZN(n7744) );
  NAND2_X1 U7481 ( .A1(n7465), .A2(n9557), .ZN(n7464) );
  NAND2_X1 U7482 ( .A1(n7467), .A2(n7466), .ZN(n7465) );
  NOR3_X1 U7483 ( .A1(n12901), .A2(n12900), .A3(n7208), .ZN(n6914) );
  NOR2_X1 U7484 ( .A1(n12922), .A2(n12921), .ZN(n7208) );
  NAND2_X1 U7485 ( .A1(n12955), .A2(n7234), .ZN(n7233) );
  AND2_X1 U7486 ( .A1(n9313), .A2(n11958), .ZN(n9336) );
  INV_X1 U7487 ( .A(n7558), .ZN(n6890) );
  NOR2_X1 U7488 ( .A1(n9488), .A2(n9486), .ZN(n9320) );
  OR2_X1 U7489 ( .A1(n12261), .A2(n12262), .ZN(n7070) );
  OR2_X1 U7490 ( .A1(n12050), .A2(n12428), .ZN(n9355) );
  AND2_X1 U7491 ( .A1(n12780), .A2(n8192), .ZN(n7243) );
  AOI21_X1 U7492 ( .B1(n7423), .B2(n7426), .A(n6563), .ZN(n7420) );
  NAND2_X1 U7493 ( .A1(n9768), .A2(n10661), .ZN(n7336) );
  NAND2_X1 U7494 ( .A1(n7335), .A2(n7334), .ZN(n6779) );
  INV_X1 U7495 ( .A(n7901), .ZN(n8131) );
  INV_X1 U7496 ( .A(n11515), .ZN(n13029) );
  NAND2_X1 U7497 ( .A1(n10053), .A2(n9925), .ZN(n7922) );
  OR2_X1 U7498 ( .A1(n7641), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n7645) );
  INV_X1 U7499 ( .A(n13757), .ZN(n13599) );
  INV_X1 U7500 ( .A(n12837), .ZN(n6899) );
  NOR2_X1 U7501 ( .A1(n12840), .A2(n12837), .ZN(n6900) );
  AND2_X1 U7502 ( .A1(n9553), .A2(n7468), .ZN(n7467) );
  INV_X1 U7503 ( .A(n9571), .ZN(n6734) );
  OAI21_X1 U7504 ( .B1(n9591), .B2(n7494), .A(n7491), .ZN(n9593) );
  NAND2_X1 U7505 ( .A1(n7495), .A2(n9682), .ZN(n7494) );
  NOR2_X1 U7506 ( .A1(n7493), .A2(n7492), .ZN(n7491) );
  INV_X1 U7507 ( .A(n7496), .ZN(n7495) );
  NAND2_X1 U7508 ( .A1(n7229), .A2(n12929), .ZN(n7228) );
  NAND2_X1 U7509 ( .A1(n6921), .A2(n6550), .ZN(n6920) );
  INV_X1 U7510 ( .A(n7231), .ZN(n6921) );
  MUX2_X1 U7511 ( .A(n12796), .B(n12795), .S(n6461), .Z(n12806) );
  OR2_X1 U7512 ( .A1(n9504), .A2(n13858), .ZN(n7462) );
  NAND2_X1 U7513 ( .A1(n9644), .A2(n7476), .ZN(n7475) );
  INV_X1 U7514 ( .A(n6806), .ZN(n6804) );
  NOR2_X1 U7515 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7619) );
  INV_X1 U7516 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6917) );
  INV_X1 U7517 ( .A(n9647), .ZN(n7478) );
  AOI21_X1 U7518 ( .B1(n6711), .B2(n6710), .A(n6600), .ZN(n7576) );
  INV_X1 U7519 ( .A(n8068), .ZN(n6710) );
  INV_X1 U7520 ( .A(n8069), .ZN(n6711) );
  OR2_X1 U7521 ( .A1(n7576), .A2(SI_20_), .ZN(n7440) );
  INV_X1 U7522 ( .A(n6889), .ZN(n6888) );
  OAI21_X1 U7523 ( .B1(n7959), .B2(n6890), .A(n7561), .ZN(n6889) );
  INV_X1 U7524 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8412) );
  AND2_X1 U7525 ( .A1(n9320), .A2(n9314), .ZN(n6626) );
  INV_X1 U7526 ( .A(n12542), .ZN(n9819) );
  INV_X1 U7527 ( .A(n12393), .ZN(n7446) );
  OR2_X1 U7528 ( .A1(n12406), .A2(n12416), .ZN(n9353) );
  NAND2_X1 U7529 ( .A1(n12479), .A2(n9211), .ZN(n6748) );
  NAND2_X1 U7530 ( .A1(n7118), .A2(n6543), .ZN(n11197) );
  NAND2_X1 U7531 ( .A1(n7120), .A2(n7122), .ZN(n7119) );
  AOI21_X1 U7532 ( .B1(n7133), .B2(n9472), .A(n7131), .ZN(n7130) );
  INV_X1 U7533 ( .A(n9167), .ZN(n7131) );
  NAND2_X1 U7534 ( .A1(n6778), .A2(n11764), .ZN(n6777) );
  XNOR2_X1 U7535 ( .A(n11702), .B(P3_B_REG_SCAN_IN), .ZN(n6778) );
  INV_X1 U7536 ( .A(n7290), .ZN(n7288) );
  INV_X1 U7537 ( .A(n8715), .ZN(n7292) );
  NOR2_X2 U7538 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n10404) );
  XNOR2_X1 U7539 ( .A(n8210), .B(n12849), .ZN(n7833) );
  OR2_X1 U7540 ( .A1(n13314), .A2(n12957), .ZN(n11900) );
  INV_X1 U7541 ( .A(n12987), .ZN(n7159) );
  NOR2_X1 U7542 ( .A1(n11899), .A2(n7162), .ZN(n7160) );
  INV_X1 U7543 ( .A(n11559), .ZN(n7146) );
  INV_X1 U7544 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7617) );
  INV_X1 U7545 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7616) );
  INV_X1 U7546 ( .A(n7625), .ZN(n6918) );
  AND2_X1 U7547 ( .A1(n6524), .A2(n11264), .ZN(n7379) );
  XNOR2_X1 U7548 ( .A(n13866), .B(n13864), .ZN(n9709) );
  NOR2_X1 U7549 ( .A1(n9645), .A2(n6959), .ZN(n6958) );
  NOR2_X1 U7550 ( .A1(n13927), .A2(n6845), .ZN(n6844) );
  INV_X1 U7551 ( .A(n8685), .ZN(n6845) );
  INV_X1 U7552 ( .A(n6838), .ZN(n6837) );
  OAI21_X1 U7553 ( .B1(n7253), .B2(n6839), .A(n11753), .ZN(n6838) );
  INV_X1 U7554 ( .A(n9575), .ZN(n6839) );
  NAND2_X1 U7555 ( .A1(n9504), .A2(n13858), .ZN(n9505) );
  OR2_X1 U7556 ( .A1(n14414), .A2(n13495), .ZN(n9575) );
  NAND2_X1 U7557 ( .A1(n7576), .A2(SI_20_), .ZN(n8106) );
  NAND3_X1 U7558 ( .A1(n7440), .A2(n8088), .A3(n8106), .ZN(n8086) );
  INV_X1 U7559 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8507) );
  XNOR2_X1 U7560 ( .A(n7565), .B(SI_16_), .ZN(n8011) );
  NOR2_X1 U7561 ( .A1(n7918), .A2(n7429), .ZN(n7428) );
  INV_X1 U7562 ( .A(n7553), .ZN(n7429) );
  AND2_X1 U7563 ( .A1(n7510), .A2(n7549), .ZN(n7450) );
  AND2_X2 U7564 ( .A1(n8314), .A2(n6666), .ZN(n8486) );
  INV_X1 U7565 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8226) );
  XNOR2_X1 U7566 ( .A(n7534), .B(SI_4_), .ZN(n7782) );
  OAI21_X1 U7567 ( .B1(n9882), .B2(n8818), .A(n8275), .ZN(n7741) );
  NAND2_X1 U7568 ( .A1(n9775), .A2(n10786), .ZN(n7363) );
  AOI21_X1 U7569 ( .B1(n7351), .B2(n7350), .A(n6598), .ZN(n7349) );
  NAND2_X1 U7570 ( .A1(n6812), .A2(n6488), .ZN(n7347) );
  AND2_X1 U7571 ( .A1(n7359), .A2(n7363), .ZN(n7361) );
  INV_X1 U7572 ( .A(n10651), .ZN(n7359) );
  NOR2_X1 U7573 ( .A1(n9796), .A2(n6818), .ZN(n6817) );
  INV_X1 U7574 ( .A(n9791), .ZN(n6818) );
  XNOR2_X1 U7575 ( .A(n10315), .B(n15031), .ZN(n7330) );
  AND2_X1 U7576 ( .A1(n8774), .A2(n8775), .ZN(n8823) );
  NAND2_X1 U7577 ( .A1(n6986), .A2(n6985), .ZN(n11518) );
  INV_X1 U7578 ( .A(n11230), .ZN(n6985) );
  AND2_X1 U7579 ( .A1(n6863), .A2(n6864), .ZN(n11615) );
  AOI21_X1 U7580 ( .B1(n6866), .B2(n6871), .A(n11524), .ZN(n6864) );
  OR2_X1 U7581 ( .A1(n11070), .A2(n6865), .ZN(n6863) );
  INV_X1 U7582 ( .A(n6866), .ZN(n6865) );
  OR2_X1 U7583 ( .A1(n11785), .A2(n12583), .ZN(n6763) );
  NAND2_X1 U7584 ( .A1(n7050), .A2(n7049), .ZN(n7048) );
  INV_X1 U7585 ( .A(n12212), .ZN(n7049) );
  INV_X1 U7586 ( .A(n12220), .ZN(n6992) );
  NAND2_X1 U7587 ( .A1(n7070), .A2(n6620), .ZN(n7064) );
  OR2_X1 U7588 ( .A1(n12293), .A2(n12292), .ZN(n12315) );
  OR2_X1 U7589 ( .A1(n12155), .A2(n12367), .ZN(n9223) );
  NAND2_X1 U7590 ( .A1(n12369), .A2(n12368), .ZN(n6631) );
  INV_X1 U7591 ( .A(n12364), .ZN(n12389) );
  NAND2_X1 U7592 ( .A1(n12412), .A2(n9216), .ZN(n12402) );
  NAND2_X1 U7593 ( .A1(n6630), .A2(n9355), .ZN(n12405) );
  XNOR2_X1 U7594 ( .A(n12115), .B(n12441), .ZN(n12429) );
  NAND2_X1 U7595 ( .A1(n12454), .A2(n9085), .ZN(n12443) );
  AND2_X1 U7596 ( .A1(n9437), .A2(n9434), .ZN(n12485) );
  NAND2_X1 U7597 ( .A1(n6628), .A2(n9435), .ZN(n12502) );
  NOR2_X1 U7598 ( .A1(n11456), .A2(n7435), .ZN(n7434) );
  INV_X1 U7599 ( .A(n7437), .ZN(n7435) );
  AND2_X1 U7600 ( .A1(n9271), .A2(n9270), .ZN(n10283) );
  AND2_X1 U7602 ( .A1(n7329), .A2(n7328), .ZN(n9303) );
  NAND2_X1 U7603 ( .A1(n15205), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7328) );
  OR2_X1 U7604 ( .A1(n9291), .A2(n9290), .ZN(n7329) );
  NAND2_X1 U7605 ( .A1(n8733), .A2(n8732), .ZN(n9087) );
  NAND2_X1 U7606 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11086), .ZN(n8732) );
  NAND2_X1 U7607 ( .A1(n9073), .A2(n9071), .ZN(n8733) );
  XNOR2_X1 U7608 ( .A(n9075), .B(P3_IR_REG_19__SCAN_IN), .ZN(n9767) );
  OAI21_X1 U7609 ( .B1(n9074), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9075) );
  INV_X1 U7610 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8818) );
  AOI21_X1 U7611 ( .B1(n12746), .B2(n12745), .A(n8142), .ZN(n8157) );
  AND2_X1 U7612 ( .A1(n7243), .A2(n6945), .ZN(n6944) );
  NAND2_X1 U7613 ( .A1(n6947), .A2(n8190), .ZN(n6945) );
  INV_X1 U7614 ( .A(n7242), .ZN(n7239) );
  XNOR2_X1 U7615 ( .A(n13088), .B(n13091), .ZN(n13025) );
  XNOR2_X1 U7616 ( .A(n12007), .B(n14826), .ZN(n14816) );
  INV_X1 U7617 ( .A(n13402), .ZN(n13124) );
  OR2_X1 U7618 ( .A1(n13219), .A2(n11921), .ZN(n11923) );
  NOR2_X1 U7619 ( .A1(n13386), .A2(n11398), .ZN(n11564) );
  NAND2_X1 U7620 ( .A1(n6657), .A2(n13065), .ZN(n10595) );
  NAND2_X1 U7621 ( .A1(n10338), .A2(n10337), .ZN(n13198) );
  OR2_X1 U7622 ( .A1(n6742), .A2(n13026), .ZN(n10338) );
  NAND2_X1 U7623 ( .A1(n11902), .A2(n11901), .ZN(n13308) );
  NAND2_X1 U7624 ( .A1(n13030), .A2(n6742), .ZN(n14895) );
  INV_X1 U7625 ( .A(n8295), .ZN(n8305) );
  NAND2_X1 U7626 ( .A1(n7180), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n8464) );
  NOR2_X1 U7627 ( .A1(n13790), .A2(n13791), .ZN(n13789) );
  NOR2_X1 U7628 ( .A1(n13836), .A2(n14581), .ZN(n13837) );
  NOR2_X1 U7629 ( .A1(n13850), .A2(n6966), .ZN(n6967) );
  OR2_X1 U7630 ( .A1(n13837), .A2(n8501), .ZN(n6965) );
  INV_X1 U7631 ( .A(n6959), .ZN(n6957) );
  AND2_X1 U7632 ( .A1(n8687), .A2(n8604), .ZN(n13879) );
  NOR2_X1 U7633 ( .A1(n13907), .A2(n7188), .ZN(n7187) );
  INV_X1 U7634 ( .A(n7512), .ZN(n7188) );
  NOR2_X1 U7635 ( .A1(n8678), .A2(n13766), .ZN(n7280) );
  OR2_X1 U7636 ( .A1(n14439), .A2(n14386), .ZN(n9582) );
  INV_X1 U7637 ( .A(n13858), .ZN(n14023) );
  NOR2_X1 U7638 ( .A1(n14675), .A2(n13858), .ZN(n10191) );
  NAND2_X1 U7639 ( .A1(n10202), .A2(n10013), .ZN(n14717) );
  INV_X1 U7640 ( .A(n9504), .ZN(n10202) );
  NAND2_X1 U7641 ( .A1(n14268), .A2(n14796), .ZN(n7021) );
  OAI22_X1 U7642 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14208), .B1(n14221), 
        .B2(n14207), .ZN(n14219) );
  NAND2_X1 U7643 ( .A1(n7347), .A2(n7345), .ZN(n7502) );
  AND2_X1 U7644 ( .A1(n7349), .A2(n7346), .ZN(n7345) );
  INV_X1 U7645 ( .A(n12084), .ZN(n7346) );
  NOR2_X1 U7646 ( .A1(n11057), .A2(n11058), .ZN(n11227) );
  NOR2_X1 U7647 ( .A1(n11781), .A2(n11782), .ZN(n12193) );
  AND2_X1 U7648 ( .A1(n11812), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9868) );
  OR2_X1 U7649 ( .A1(n7664), .A2(n13458), .ZN(n10057) );
  INV_X1 U7650 ( .A(n7184), .ZN(n14058) );
  NOR2_X1 U7651 ( .A1(n14476), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n14275) );
  MUX2_X1 U7652 ( .A(n9517), .B(n9516), .S(n10028), .Z(n9518) );
  AND2_X1 U7653 ( .A1(n9534), .A2(n9533), .ZN(n7480) );
  INV_X1 U7654 ( .A(n9540), .ZN(n7500) );
  NAND2_X1 U7655 ( .A1(n6718), .A2(n6716), .ZN(n6715) );
  NOR2_X1 U7656 ( .A1(n9362), .A2(n6717), .ZN(n6716) );
  NAND2_X1 U7657 ( .A1(n9363), .A2(n9184), .ZN(n6718) );
  NAND2_X1 U7658 ( .A1(n12863), .A2(n7217), .ZN(n7216) );
  OR2_X1 U7659 ( .A1(n7463), .A2(n6737), .ZN(n9559) );
  INV_X1 U7660 ( .A(n9556), .ZN(n6737) );
  OAI21_X1 U7661 ( .B1(n9552), .B2(n7467), .A(n6558), .ZN(n9558) );
  INV_X1 U7662 ( .A(n9557), .ZN(n6756) );
  NAND2_X1 U7663 ( .A1(n9565), .A2(n9566), .ZN(n9564) );
  NAND2_X1 U7664 ( .A1(n12882), .A2(n7211), .ZN(n7210) );
  NAND2_X1 U7665 ( .A1(n12885), .A2(n7212), .ZN(n7211) );
  NOR2_X1 U7666 ( .A1(n7209), .A2(n7207), .ZN(n7206) );
  INV_X1 U7667 ( .A(n12921), .ZN(n7207) );
  NOR2_X1 U7668 ( .A1(n12918), .A2(n12922), .ZN(n7209) );
  NOR2_X1 U7669 ( .A1(n12919), .A2(n12920), .ZN(n7205) );
  OAI21_X1 U7670 ( .B1(n9599), .B2(n9598), .A(n6555), .ZN(n7489) );
  INV_X1 U7671 ( .A(n12955), .ZN(n7232) );
  NAND2_X1 U7672 ( .A1(n6909), .A2(n6907), .ZN(n12948) );
  AOI21_X1 U7673 ( .B1(n6911), .B2(n6910), .A(n6908), .ZN(n6907) );
  NAND2_X1 U7674 ( .A1(n6906), .A2(n6746), .ZN(n12950) );
  AND2_X1 U7675 ( .A1(n6908), .A2(n6910), .ZN(n6746) );
  AND2_X1 U7676 ( .A1(n7233), .A2(n12952), .ZN(n7231) );
  INV_X1 U7677 ( .A(n11916), .ZN(n6640) );
  INV_X1 U7678 ( .A(n7535), .ZN(n7419) );
  INV_X1 U7679 ( .A(n7343), .ZN(n7342) );
  INV_X1 U7680 ( .A(n7340), .ZN(n6801) );
  AOI21_X1 U7681 ( .B1(n7343), .B2(n7341), .A(n9812), .ZN(n7340) );
  INV_X1 U7682 ( .A(n12110), .ZN(n7341) );
  INV_X1 U7683 ( .A(n9391), .ZN(n7122) );
  NAND2_X1 U7684 ( .A1(n12970), .A2(n12971), .ZN(n6732) );
  NAND2_X1 U7685 ( .A1(n12797), .A2(n12798), .ZN(n6733) );
  NAND2_X1 U7686 ( .A1(n13013), .A2(n11916), .ZN(n7096) );
  OR2_X1 U7687 ( .A1(n11714), .A2(n6640), .ZN(n6638) );
  OR2_X1 U7688 ( .A1(n6662), .A2(n6640), .ZN(n6639) );
  AOI21_X1 U7689 ( .B1(n7478), .B2(n7472), .A(n7471), .ZN(n7470) );
  INV_X1 U7690 ( .A(n7475), .ZN(n7472) );
  INV_X1 U7691 ( .A(n9646), .ZN(n7471) );
  NOR2_X1 U7692 ( .A1(n10017), .A2(n14628), .ZN(n9513) );
  NAND2_X1 U7693 ( .A1(n11826), .A2(n14044), .ZN(n14021) );
  NOR2_X1 U7694 ( .A1(n11827), .A2(n14423), .ZN(n11826) );
  AND2_X1 U7695 ( .A1(n7584), .A2(n7583), .ZN(n7587) );
  OR2_X1 U7696 ( .A1(n7584), .A2(n7583), .ZN(n7577) );
  AND2_X1 U7697 ( .A1(n8106), .A2(n7577), .ZN(n6891) );
  AOI21_X1 U7698 ( .B1(n7427), .B2(n7425), .A(n7424), .ZN(n7423) );
  INV_X1 U7699 ( .A(n7936), .ZN(n7424) );
  INV_X1 U7700 ( .A(n7428), .ZN(n7425) );
  INV_X1 U7701 ( .A(n7427), .ZN(n7426) );
  OAI21_X1 U7702 ( .B1(n9926), .B2(n9967), .A(n6730), .ZN(n7552) );
  NAND2_X1 U7703 ( .A1(n9926), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6730) );
  NAND2_X1 U7704 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7031), .ZN(n7030) );
  NAND2_X1 U7705 ( .A1(n14237), .A2(n14236), .ZN(n7032) );
  NAND2_X1 U7706 ( .A1(n12129), .A2(n9818), .ZN(n9823) );
  NAND2_X1 U7707 ( .A1(n9779), .A2(n15005), .ZN(n6789) );
  AND2_X1 U7708 ( .A1(n11784), .A2(n11783), .ZN(n12209) );
  INV_X1 U7709 ( .A(n12275), .ZN(n6875) );
  OR2_X1 U7710 ( .A1(n11963), .A2(n9748), .ZN(n9343) );
  AND2_X1 U7711 ( .A1(n12338), .A2(n9226), .ZN(n9228) );
  OAI21_X1 U7712 ( .B1(n12485), .B2(n9430), .A(n12470), .ZN(n7111) );
  NOR2_X1 U7713 ( .A1(n8988), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9001) );
  INV_X1 U7714 ( .A(n7116), .ZN(n7115) );
  OAI21_X1 U7715 ( .B1(n8967), .B2(n7117), .A(n14339), .ZN(n7116) );
  INV_X1 U7716 ( .A(n9409), .ZN(n7117) );
  INV_X1 U7717 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11619) );
  INV_X1 U7718 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11525) );
  AND2_X1 U7719 ( .A1(n9407), .A2(n9406), .ZN(n9325) );
  AND2_X1 U7720 ( .A1(n9343), .A2(n9342), .ZN(n11952) );
  AND2_X1 U7721 ( .A1(n8758), .A2(n7458), .ZN(n7457) );
  INV_X1 U7722 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7458) );
  AND2_X1 U7723 ( .A1(n9025), .A2(n9029), .ZN(n7365) );
  INV_X1 U7724 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9029) );
  NOR2_X1 U7725 ( .A1(n6611), .A2(n7301), .ZN(n7300) );
  NAND2_X1 U7726 ( .A1(n11906), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U7727 ( .A1(n8204), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6651) );
  AND2_X1 U7728 ( .A1(n8115), .A2(n7689), .ZN(n8149) );
  NAND2_X1 U7729 ( .A1(n11713), .A2(n13015), .ZN(n6662) );
  NOR2_X1 U7730 ( .A1(n6528), .A2(n7145), .ZN(n7144) );
  NOR2_X1 U7731 ( .A1(n11392), .A2(n7146), .ZN(n7145) );
  OR2_X1 U7732 ( .A1(n7941), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n7978) );
  OR2_X1 U7733 ( .A1(n7840), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n7858) );
  INV_X1 U7734 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7613) );
  INV_X1 U7735 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6916) );
  CLKBUF_X1 U7736 ( .A(n7786), .Z(n7787) );
  INV_X1 U7737 ( .A(n13640), .ZN(n7400) );
  INV_X1 U7738 ( .A(n13673), .ZN(n7405) );
  OAI22_X1 U7739 ( .A1(n9633), .A2(n6676), .B1(n6677), .B2(n9634), .ZN(n9637)
         );
  AND2_X1 U7740 ( .A1(n9634), .A2(n6677), .ZN(n6676) );
  INV_X1 U7741 ( .A(n9632), .ZN(n6677) );
  NAND2_X1 U7742 ( .A1(n8295), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8298) );
  INV_X1 U7743 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8236) );
  NAND2_X1 U7744 ( .A1(n14555), .A2(n13835), .ZN(n13836) );
  NAND2_X1 U7745 ( .A1(n6960), .A2(n13904), .ZN(n6959) );
  AND2_X1 U7746 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n8595), .ZN(n8596) );
  NOR2_X1 U7747 ( .A1(n14021), .A2(n14027), .ZN(n6950) );
  OR2_X1 U7748 ( .A1(n14027), .A2(n13711), .ZN(n9601) );
  AND2_X1 U7749 ( .A1(n14413), .A2(n7254), .ZN(n7253) );
  NAND2_X1 U7750 ( .A1(n7256), .A2(n9694), .ZN(n7254) );
  OR2_X1 U7751 ( .A1(n10476), .A2(n10847), .ZN(n9525) );
  NAND2_X1 U7752 ( .A1(n10476), .A2(n10847), .ZN(n9524) );
  NAND2_X1 U7753 ( .A1(n9521), .A2(n9519), .ZN(n9686) );
  NAND2_X1 U7754 ( .A1(n10028), .A2(n14652), .ZN(n8654) );
  NAND2_X1 U7755 ( .A1(n10754), .A2(n10751), .ZN(n7283) );
  NAND2_X1 U7756 ( .A1(n11454), .A2(n10202), .ZN(n10201) );
  INV_X1 U7757 ( .A(n7431), .ZN(n6698) );
  AOI21_X1 U7758 ( .B1(n6697), .B2(n7431), .A(n6696), .ZN(n6695) );
  INV_X1 U7759 ( .A(n9648), .ZN(n6697) );
  INV_X1 U7760 ( .A(n9670), .ZN(n6696) );
  NAND2_X1 U7761 ( .A1(n9649), .A2(n9648), .ZN(n7433) );
  AND2_X1 U7762 ( .A1(n9651), .A2(n7432), .ZN(n7431) );
  INV_X1 U7763 ( .A(n9653), .ZN(n7432) );
  OAI22_X1 U7764 ( .A1(n7729), .A2(n7449), .B1(n7730), .B2(n11852), .ZN(n8196)
         );
  NOR2_X1 U7765 ( .A1(n7603), .A2(SI_26_), .ZN(n7449) );
  INV_X1 U7766 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U7767 ( .A1(n7578), .A2(SI_21_), .ZN(n7583) );
  NOR2_X1 U7768 ( .A1(n7572), .A2(SI_18_), .ZN(n6701) );
  INV_X1 U7769 ( .A(n6693), .ZN(n6692) );
  OAI21_X1 U7770 ( .B1(n6884), .B2(n6694), .A(n7566), .ZN(n6693) );
  XNOR2_X1 U7771 ( .A(n7567), .B(SI_17_), .ZN(n8026) );
  NOR2_X1 U7772 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n8229) );
  NOR2_X1 U7773 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8228) );
  INV_X1 U7774 ( .A(n7822), .ZN(n7540) );
  INV_X1 U7775 ( .A(n7782), .ZN(n7533) );
  OAI21_X1 U7776 ( .B1(n7524), .B2(n9942), .A(n6709), .ZN(n7527) );
  NAND2_X1 U7777 ( .A1(n7524), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6709) );
  AOI21_X1 U7778 ( .B1(n11959), .B2(n12179), .A(n11954), .ZN(n9836) );
  AOI21_X1 U7779 ( .B1(n6798), .B2(n9835), .A(n6795), .ZN(n6794) );
  NOR2_X1 U7780 ( .A1(n9836), .A2(n6796), .ZN(n6795) );
  OR2_X1 U7781 ( .A1(n12158), .A2(n9835), .ZN(n6796) );
  AOI21_X1 U7782 ( .B1(n6814), .B2(n6811), .A(n6599), .ZN(n6810) );
  INV_X1 U7783 ( .A(n6817), .ZN(n6811) );
  OR2_X1 U7784 ( .A1(n11662), .A2(n6813), .ZN(n6812) );
  INV_X1 U7785 ( .A(n6814), .ZN(n6813) );
  AND2_X1 U7786 ( .A1(n9836), .A2(n6799), .ZN(n6798) );
  OR2_X1 U7787 ( .A1(n12158), .A2(n9835), .ZN(n6799) );
  AND2_X1 U7788 ( .A1(n12052), .A2(n6499), .ZN(n7343) );
  AND2_X1 U7789 ( .A1(n9102), .A2(n12054), .ZN(n9112) );
  AND2_X1 U7790 ( .A1(n9833), .A2(n9831), .ZN(n12075) );
  INV_X1 U7791 ( .A(n9786), .ZN(n7354) );
  AOI21_X1 U7792 ( .B1(n12043), .B2(n6807), .A(n6530), .ZN(n6806) );
  INV_X1 U7793 ( .A(n6809), .ZN(n6807) );
  OR2_X1 U7794 ( .A1(n6786), .A2(n6784), .ZN(n6783) );
  INV_X1 U7795 ( .A(n6789), .ZN(n6784) );
  AND2_X1 U7796 ( .A1(n6787), .A2(n10915), .ZN(n6786) );
  NAND2_X1 U7797 ( .A1(n6788), .A2(n6790), .ZN(n6787) );
  NAND2_X1 U7798 ( .A1(n6790), .A2(n6789), .ZN(n6785) );
  NAND2_X1 U7799 ( .A1(n9799), .A2(n12025), .ZN(n7352) );
  MUX2_X1 U7800 ( .A(n9484), .B(n9483), .S(n9499), .Z(n9487) );
  NAND2_X1 U7801 ( .A1(n9320), .A2(n7323), .ZN(n7322) );
  NOR2_X1 U7802 ( .A1(n9489), .A2(n7324), .ZN(n7323) );
  NAND2_X1 U7803 ( .A1(n9485), .A2(n7325), .ZN(n7324) );
  NOR2_X1 U7804 ( .A1(n9752), .A2(n7326), .ZN(n7325) );
  NAND2_X1 U7805 ( .A1(n6625), .A2(n6546), .ZN(n9318) );
  OAI21_X1 U7806 ( .B1(n9751), .B2(n9481), .A(n6626), .ZN(n6625) );
  NAND2_X1 U7807 ( .A1(n9316), .A2(n9315), .ZN(n9317) );
  AND4_X1 U7808 ( .A1(n8900), .A2(n8899), .A3(n8898), .A4(n8897), .ZN(n11311)
         );
  OAI21_X1 U7809 ( .B1(n10456), .B2(n10396), .A(n6501), .ZN(n10446) );
  INV_X1 U7810 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n14179) );
  NAND2_X1 U7811 ( .A1(n7079), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7077) );
  NAND2_X1 U7812 ( .A1(n7080), .A2(n11059), .ZN(n7079) );
  INV_X1 U7813 ( .A(n10679), .ZN(n7080) );
  NAND2_X1 U7814 ( .A1(n6872), .A2(n6869), .ZN(n6868) );
  NAND2_X1 U7815 ( .A1(n7072), .A2(n7071), .ZN(n11531) );
  AND2_X1 U7816 ( .A1(n6868), .A2(n6604), .ZN(n6866) );
  NAND2_X1 U7817 ( .A1(n11070), .A2(n6870), .ZN(n6867) );
  NAND2_X1 U7818 ( .A1(n11616), .A2(n11617), .ZN(n11789) );
  OR2_X1 U7819 ( .A1(n11604), .A2(n11605), .ZN(n6991) );
  NAND2_X1 U7820 ( .A1(n7081), .A2(n11614), .ZN(n11784) );
  OAI211_X1 U7821 ( .C1(n12249), .C2(n6980), .A(n6978), .B(n6977), .ZN(n12283)
         );
  NAND2_X1 U7822 ( .A1(n6981), .A2(n12296), .ZN(n6980) );
  INV_X1 U7823 ( .A(n6979), .ZN(n6978) );
  NAND2_X1 U7824 ( .A1(n7070), .A2(n7069), .ZN(n12272) );
  OR2_X1 U7825 ( .A1(n9228), .A2(n9227), .ZN(n9229) );
  INV_X1 U7826 ( .A(n9223), .ZN(n7134) );
  AND2_X1 U7827 ( .A1(n8791), .A2(n8790), .ZN(n12353) );
  AOI21_X1 U7828 ( .B1(n7444), .B2(n12401), .A(n6548), .ZN(n7443) );
  AND2_X1 U7829 ( .A1(n9351), .A2(n9350), .ZN(n12393) );
  NAND2_X1 U7830 ( .A1(n7447), .A2(n9217), .ZN(n12388) );
  NAND2_X1 U7831 ( .A1(n12402), .A2(n12404), .ZN(n7447) );
  NAND2_X1 U7832 ( .A1(n7442), .A2(n7441), .ZN(n12412) );
  AND2_X1 U7833 ( .A1(n9215), .A2(n9214), .ZN(n7441) );
  AND2_X1 U7834 ( .A1(n9355), .A2(n9354), .ZN(n12417) );
  AND4_X1 U7835 ( .A1(n9069), .A2(n9068), .A3(n9067), .A4(n9066), .ZN(n12440)
         );
  INV_X1 U7836 ( .A(n6748), .ZN(n12465) );
  NAND2_X1 U7837 ( .A1(n12465), .A2(n12464), .ZN(n12463) );
  NAND2_X1 U7838 ( .A1(n12486), .A2(n12485), .ZN(n12488) );
  NAND2_X1 U7839 ( .A1(n12494), .A2(n6534), .ZN(n12479) );
  INV_X1 U7840 ( .A(n12485), .ZN(n9210) );
  AND4_X1 U7841 ( .A1(n9006), .A2(n9005), .A3(n9004), .A4(n9003), .ZN(n12514)
         );
  AND2_X1 U7842 ( .A1(n9417), .A2(n9415), .ZN(n14339) );
  NAND2_X1 U7843 ( .A1(n8968), .A2(n8967), .ZN(n11511) );
  INV_X1 U7844 ( .A(n9325), .ZN(n11410) );
  AND4_X1 U7845 ( .A1(n8946), .A2(n8945), .A3(n8944), .A4(n8943), .ZN(n12140)
         );
  NAND2_X1 U7846 ( .A1(n9199), .A2(n7438), .ZN(n7436) );
  NOR2_X1 U7847 ( .A1(n9200), .A2(n7439), .ZN(n7438) );
  INV_X1 U7848 ( .A(n9198), .ZN(n7439) );
  OR2_X1 U7849 ( .A1(n14968), .A2(n11315), .ZN(n7437) );
  INV_X1 U7850 ( .A(n15039), .ZN(n12512) );
  AND2_X1 U7851 ( .A1(n9393), .A2(n9392), .ZN(n14965) );
  OR2_X1 U7852 ( .A1(n8878), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8894) );
  NAND2_X1 U7853 ( .A1(n9859), .A2(n10389), .ZN(n15019) );
  NAND2_X1 U7854 ( .A1(n9754), .A2(n9340), .ZN(n15039) );
  AND2_X1 U7855 ( .A1(n9845), .A2(n10389), .ZN(n15035) );
  OR2_X1 U7856 ( .A1(n8839), .A2(n9914), .ZN(n8814) );
  OAI211_X1 U7857 ( .C1(n10285), .C2(n10284), .A(n10283), .B(n10282), .ZN(
        n10287) );
  NAND2_X1 U7858 ( .A1(n9158), .A2(n9157), .ZN(n12155) );
  OR2_X1 U7859 ( .A1(n9295), .A2(n11852), .ZN(n9157) );
  NAND2_X1 U7860 ( .A1(n9145), .A2(n9144), .ZN(n12072) );
  OR2_X1 U7861 ( .A1(n9295), .A2(n15233), .ZN(n9144) );
  NAND2_X1 U7862 ( .A1(n9101), .A2(n9100), .ZN(n12050) );
  OR2_X1 U7863 ( .A1(n9295), .A2(n10880), .ZN(n9100) );
  NAND2_X1 U7864 ( .A1(n9046), .A2(n9045), .ZN(n12095) );
  AND2_X1 U7865 ( .A1(n8954), .A2(n8953), .ZN(n9789) );
  OR2_X1 U7866 ( .A1(n8822), .A2(n8803), .ZN(n8806) );
  INV_X1 U7867 ( .A(n15035), .ZN(n15017) );
  NAND2_X1 U7868 ( .A1(n6777), .A2(n6525), .ZN(n9250) );
  NAND2_X1 U7869 ( .A1(n8772), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8769) );
  NAND2_X1 U7870 ( .A1(n6752), .A2(n6627), .ZN(n8759) );
  NOR2_X1 U7871 ( .A1(n6750), .A2(n8971), .ZN(n6627) );
  NAND2_X1 U7872 ( .A1(n6751), .A2(n8762), .ZN(n6750) );
  AND2_X1 U7873 ( .A1(n7318), .A2(n8743), .ZN(n9284) );
  OAI21_X1 U7874 ( .B1(n9129), .B2(n11845), .A(n6508), .ZN(n7320) );
  INV_X1 U7875 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8755) );
  INV_X1 U7876 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8754) );
  XNOR2_X1 U7877 ( .A(n8741), .B(P2_DATAO_REG_24__SCAN_IN), .ZN(n9129) );
  NOR2_X1 U7878 ( .A1(n8738), .A2(n8737), .ZN(n9117) );
  AND2_X1 U7879 ( .A1(n8736), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8737) );
  NAND2_X1 U7880 ( .A1(n7305), .A2(n6497), .ZN(n7304) );
  NOR2_X1 U7881 ( .A1(n9098), .A2(n7307), .ZN(n7306) );
  INV_X1 U7882 ( .A(n7308), .ZN(n7307) );
  NAND2_X1 U7883 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n15251), .ZN(n7308) );
  NAND2_X1 U7884 ( .A1(n9087), .A2(n9086), .ZN(n8734) );
  AND2_X1 U7885 ( .A1(n9178), .A2(n9177), .ZN(n9338) );
  AOI21_X1 U7886 ( .B1(n6601), .B2(n8730), .A(n7312), .ZN(n7311) );
  INV_X1 U7887 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9025) );
  AND2_X1 U7888 ( .A1(n6577), .A2(n8749), .ZN(n6820) );
  AND2_X1 U7889 ( .A1(n10037), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8719) );
  AOI21_X1 U7890 ( .B1(n7291), .B2(n8714), .A(n6492), .ZN(n7290) );
  INV_X1 U7891 ( .A(n8918), .ZN(n7295) );
  INV_X1 U7892 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U7893 ( .A1(n7314), .A2(n7313), .ZN(n8888) );
  AND2_X1 U7894 ( .A1(n8711), .A2(n8709), .ZN(n7313) );
  NAND2_X1 U7895 ( .A1(n8708), .A2(n8707), .ZN(n8865) );
  XNOR2_X1 U7896 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8864) );
  INV_X1 U7897 ( .A(n10404), .ZN(n8813) );
  NAND2_X1 U7898 ( .A1(n8811), .A2(n7076), .ZN(n7075) );
  INV_X1 U7899 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7076) );
  NOR2_X1 U7900 ( .A1(n10910), .A2(n7245), .ZN(n7244) );
  INV_X1 U7901 ( .A(n7821), .ZN(n7245) );
  OR2_X1 U7902 ( .A1(n8193), .A2(n8194), .ZN(n7242) );
  NAND2_X1 U7903 ( .A1(n8174), .A2(n12727), .ZN(n6948) );
  NOR2_X1 U7904 ( .A1(n8216), .A2(n12759), .ZN(n7241) );
  NOR2_X1 U7905 ( .A1(n7237), .A2(n7243), .ZN(n7236) );
  NAND2_X1 U7906 ( .A1(n8149), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8179) );
  INV_X1 U7907 ( .A(n11540), .ZN(n6937) );
  NAND2_X1 U7908 ( .A1(n6933), .A2(n6939), .ZN(n6930) );
  OR2_X1 U7909 ( .A1(n8000), .A2(n11836), .ZN(n8018) );
  AND2_X1 U7910 ( .A1(n13038), .A2(n13029), .ZN(n10052) );
  AND2_X1 U7911 ( .A1(n7699), .A2(n7698), .ZN(n12956) );
  NAND2_X1 U7912 ( .A1(n14755), .A2(n14756), .ZN(n14754) );
  NAND2_X1 U7913 ( .A1(n10090), .A2(n10091), .ZN(n10112) );
  NAND2_X1 U7914 ( .A1(n10306), .A2(n6624), .ZN(n10540) );
  NOR2_X1 U7915 ( .A1(n12005), .A2(n6617), .ZN(n12007) );
  NOR2_X1 U7916 ( .A1(n14816), .A2(n14815), .ZN(n14814) );
  OR2_X1 U7917 ( .A1(n7678), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n8028) );
  AND2_X1 U7918 ( .A1(n11900), .A2(n11885), .ZN(n13112) );
  INV_X1 U7919 ( .A(n13314), .ZN(n13111) );
  OAI21_X1 U7920 ( .B1(n7097), .B2(n6892), .A(n6559), .ZN(n13121) );
  NOR2_X1 U7921 ( .A1(n13322), .A2(n13046), .ZN(n6892) );
  OAI21_X1 U7922 ( .B1(n13151), .B2(n7099), .A(n7098), .ZN(n7097) );
  AND2_X1 U7923 ( .A1(n13327), .A2(n13047), .ZN(n7099) );
  NAND2_X1 U7924 ( .A1(n7044), .A2(n12772), .ZN(n7098) );
  NAND2_X1 U7925 ( .A1(n13327), .A2(n12772), .ZN(n7162) );
  NAND2_X1 U7926 ( .A1(n13162), .A2(n7100), .ZN(n13151) );
  NAND2_X1 U7927 ( .A1(n12946), .A2(n13048), .ZN(n7100) );
  OAI21_X1 U7928 ( .B1(n13200), .B2(n7168), .A(n7166), .ZN(n7518) );
  NAND2_X1 U7929 ( .A1(n7166), .A2(n7168), .ZN(n7165) );
  AND2_X1 U7930 ( .A1(n6643), .A2(n6642), .ZN(n13164) );
  NAND2_X1 U7931 ( .A1(n13412), .A2(n12730), .ZN(n6642) );
  NAND2_X1 U7932 ( .A1(n13178), .A2(n13179), .ZN(n6643) );
  NAND2_X1 U7933 ( .A1(n13190), .A2(n6512), .ZN(n7103) );
  NAND2_X1 U7934 ( .A1(n11923), .A2(n6506), .ZN(n7104) );
  AND2_X1 U7935 ( .A1(n11896), .A2(n11887), .ZN(n13201) );
  INV_X1 U7936 ( .A(n13016), .ZN(n13210) );
  AOI21_X1 U7937 ( .B1(n7093), .B2(n7091), .A(n7090), .ZN(n7089) );
  INV_X1 U7938 ( .A(n7093), .ZN(n7092) );
  INV_X1 U7939 ( .A(n12990), .ZN(n7090) );
  NAND2_X1 U7940 ( .A1(n7095), .A2(n13266), .ZN(n13265) );
  AND2_X1 U7941 ( .A1(n12912), .A2(n12913), .ZN(n13283) );
  NAND2_X1 U7942 ( .A1(n6662), .A2(n11714), .ZN(n11715) );
  OR2_X1 U7943 ( .A1(n11715), .A2(n13013), .ZN(n11917) );
  NAND2_X1 U7944 ( .A1(n11654), .A2(n12886), .ZN(n11710) );
  NAND2_X1 U7945 ( .A1(n6649), .A2(n11402), .ZN(n11570) );
  NAND2_X1 U7946 ( .A1(n11401), .A2(n11400), .ZN(n6649) );
  NAND2_X1 U7947 ( .A1(n11393), .A2(n11392), .ZN(n11560) );
  NAND2_X1 U7948 ( .A1(n6648), .A2(n10959), .ZN(n11036) );
  NAND2_X1 U7949 ( .A1(n11133), .A2(n11132), .ZN(n6648) );
  NAND2_X1 U7950 ( .A1(n11135), .A2(n13002), .ZN(n11134) );
  NAND2_X1 U7951 ( .A1(n10594), .A2(n10593), .ZN(n10956) );
  NAND2_X1 U7952 ( .A1(n9890), .A2(n7901), .ZN(n7250) );
  NAND2_X1 U7953 ( .A1(n10612), .A2(n12994), .ZN(n6636) );
  INV_X1 U7954 ( .A(n9943), .ZN(n6727) );
  NAND2_X1 U7955 ( .A1(n10574), .A2(n10573), .ZN(n10833) );
  NAND2_X1 U7956 ( .A1(n6723), .A2(n12800), .ZN(n13088) );
  NAND2_X1 U7957 ( .A1(n13440), .A2(n12782), .ZN(n6723) );
  NAND2_X1 U7958 ( .A1(n13314), .A2(n14891), .ZN(n6775) );
  NAND2_X1 U7959 ( .A1(n8114), .A2(n8113), .ZN(n13212) );
  OR2_X1 U7960 ( .A1(n11557), .A2(n8131), .ZN(n8114) );
  NAND2_X1 U7961 ( .A1(n7962), .A2(n7961), .ZN(n13386) );
  INV_X1 U7962 ( .A(n8131), .ZN(n12782) );
  AND2_X1 U7963 ( .A1(n10336), .A2(n14895), .ZN(n14851) );
  CLKBUF_X1 U7964 ( .A(n10335), .Z(n10336) );
  INV_X1 U7965 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7203) );
  AND2_X1 U7966 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n7628) );
  OR2_X1 U7967 ( .A1(n7665), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n7641) );
  INV_X1 U7968 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n7670) );
  INV_X1 U7969 ( .A(n7678), .ZN(n6644) );
  AND2_X1 U7970 ( .A1(n11847), .A2(n14162), .ZN(n6767) );
  AOI21_X1 U7971 ( .B1(n13597), .B2(n13595), .A(n13624), .ZN(n7387) );
  INV_X1 U7972 ( .A(n7387), .ZN(n7384) );
  NAND2_X1 U7973 ( .A1(n11262), .A2(n11261), .ZN(n7380) );
  XNOR2_X1 U7974 ( .A(n6688), .B(n13561), .ZN(n10156) );
  NAND2_X1 U7975 ( .A1(n10152), .A2(n10151), .ZN(n6688) );
  AND3_X1 U7976 ( .A1(n14159), .A2(n9993), .A3(n6459), .ZN(n6683) );
  AND2_X1 U7977 ( .A1(n13671), .A2(n7410), .ZN(n7409) );
  NAND2_X1 U7978 ( .A1(n13663), .A2(n13673), .ZN(n7410) );
  NAND2_X1 U7979 ( .A1(n7380), .A2(n7379), .ZN(n11332) );
  AND2_X1 U7980 ( .A1(n11331), .A2(n7376), .ZN(n7375) );
  NAND2_X1 U7981 ( .A1(n7379), .A2(n7377), .ZN(n7376) );
  INV_X1 U7982 ( .A(n11261), .ZN(n7377) );
  INV_X1 U7983 ( .A(n7379), .ZN(n7378) );
  NAND2_X1 U7984 ( .A1(n11637), .A2(n6540), .ZN(n11681) );
  NAND2_X1 U7985 ( .A1(n11632), .A2(n11631), .ZN(n11637) );
  NAND2_X1 U7986 ( .A1(n13717), .A2(n11015), .ZN(n13718) );
  AOI21_X1 U7987 ( .B1(n7392), .B2(n7390), .A(n7389), .ZN(n7388) );
  INV_X1 U7988 ( .A(n7392), .ZN(n7391) );
  INV_X1 U7989 ( .A(n13486), .ZN(n7390) );
  XNOR2_X1 U7990 ( .A(n7452), .B(n14023), .ZN(n9706) );
  NAND2_X1 U7991 ( .A1(n6851), .A2(n8255), .ZN(n6850) );
  AND2_X1 U7992 ( .A1(n14155), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6851) );
  AND2_X1 U7993 ( .A1(n13788), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6970) );
  OR2_X1 U7994 ( .A1(n13801), .A2(n13800), .ZN(n6969) );
  OR2_X1 U7995 ( .A1(n9997), .A2(n9996), .ZN(n6972) );
  AND2_X1 U7996 ( .A1(n11428), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6974) );
  NOR2_X1 U7997 ( .A1(n14513), .A2(n14514), .ZN(n14515) );
  AND2_X1 U7998 ( .A1(n14525), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6975) );
  XNOR2_X1 U7999 ( .A(n13839), .B(n8458), .ZN(n11866) );
  NAND2_X1 U8000 ( .A1(n11866), .A2(n14445), .ZN(n13841) );
  NAND2_X1 U8001 ( .A1(n9676), .A2(n9675), .ZN(n13866) );
  INV_X1 U8002 ( .A(n13755), .ZN(n13628) );
  INV_X1 U8003 ( .A(n13879), .ZN(n13883) );
  NAND2_X1 U8004 ( .A1(n13904), .A2(n13634), .ZN(n7189) );
  OR2_X1 U8005 ( .A1(n14070), .A2(n13599), .ZN(n7512) );
  OAI211_X1 U8006 ( .C1(n13923), .C2(n8686), .A(n6841), .B(n13907), .ZN(n13895) );
  NAND2_X1 U8007 ( .A1(n6843), .A2(n6842), .ZN(n6841) );
  NOR2_X1 U8008 ( .A1(n8686), .A2(n6847), .ZN(n6842) );
  OR2_X1 U8009 ( .A1(n13660), .A2(n8583), .ZN(n7513) );
  NAND2_X1 U8010 ( .A1(n13913), .A2(n13912), .ZN(n13911) );
  NAND2_X1 U8011 ( .A1(n14095), .A2(n7193), .ZN(n7195) );
  NOR2_X1 U8012 ( .A1(n8683), .A2(n7194), .ZN(n7193) );
  INV_X1 U8013 ( .A(n8566), .ZN(n7194) );
  NOR2_X1 U8014 ( .A1(n13942), .A2(n7268), .ZN(n7267) );
  INV_X1 U8015 ( .A(n8682), .ZN(n7268) );
  OAI21_X1 U8016 ( .B1(n13971), .B2(n13972), .A(n6827), .ZN(n13957) );
  NAND2_X1 U8017 ( .A1(n6828), .A2(n13642), .ZN(n6827) );
  OAI21_X1 U8018 ( .B1(n14001), .B2(n7271), .A(n7269), .ZN(n13971) );
  AOI21_X1 U8019 ( .B1(n7272), .B2(n7270), .A(n6544), .ZN(n7269) );
  INV_X1 U8020 ( .A(n7272), .ZN(n7271) );
  INV_X1 U8021 ( .A(n8680), .ZN(n7270) );
  NAND2_X1 U8022 ( .A1(n13999), .A2(n7198), .ZN(n13982) );
  AND2_X1 U8023 ( .A1(n7273), .A2(n8531), .ZN(n7198) );
  NAND2_X1 U8024 ( .A1(n8521), .A2(n7199), .ZN(n13999) );
  NOR2_X1 U8025 ( .A1(n13996), .A2(n7200), .ZN(n7199) );
  INV_X1 U8026 ( .A(n8520), .ZN(n7200) );
  NAND2_X1 U8027 ( .A1(n7274), .A2(n13996), .ZN(n14003) );
  INV_X1 U8028 ( .A(n14001), .ZN(n7274) );
  AND2_X1 U8029 ( .A1(n9601), .A2(n9600), .ZN(n14017) );
  NAND2_X1 U8030 ( .A1(n7280), .A2(n7278), .ZN(n7277) );
  OR2_X1 U8031 ( .A1(n14423), .A2(n7279), .ZN(n7278) );
  AOI21_X1 U8032 ( .B1(n6837), .B2(n6839), .A(n6493), .ZN(n6836) );
  OAI21_X1 U8033 ( .B1(n7255), .B2(n6839), .A(n6837), .ZN(n11752) );
  NAND2_X1 U8034 ( .A1(n14410), .A2(n6541), .ZN(n11749) );
  AND4_X1 U8035 ( .A1(n8453), .A2(n8452), .A3(n8451), .A4(n8450), .ZN(n13495)
         );
  NAND2_X1 U8036 ( .A1(n7255), .A2(n7253), .ZN(n14406) );
  NAND2_X1 U8037 ( .A1(n8438), .A2(n7196), .ZN(n14410) );
  NOR2_X1 U8038 ( .A1(n14413), .A2(n7197), .ZN(n7196) );
  INV_X1 U8039 ( .A(n8437), .ZN(n7197) );
  AND2_X1 U8040 ( .A1(n9575), .A2(n9574), .ZN(n14413) );
  NAND2_X1 U8041 ( .A1(n11213), .A2(n8673), .ZN(n11344) );
  NAND2_X1 U8042 ( .A1(n11344), .A2(n11343), .ZN(n11342) );
  AOI21_X1 U8043 ( .B1(n10996), .B2(n7173), .A(n6551), .ZN(n7171) );
  NAND2_X1 U8044 ( .A1(n10934), .A2(n7284), .ZN(n10999) );
  NOR2_X1 U8045 ( .A1(n10996), .A2(n7285), .ZN(n7284) );
  INV_X1 U8046 ( .A(n8670), .ZN(n7285) );
  NAND2_X1 U8047 ( .A1(n7283), .A2(n7281), .ZN(n10696) );
  NOR2_X1 U8048 ( .A1(n10691), .A2(n7282), .ZN(n7281) );
  INV_X1 U8049 ( .A(n8666), .ZN(n7282) );
  NAND2_X1 U8050 ( .A1(n10696), .A2(n6848), .ZN(n10934) );
  AND2_X1 U8051 ( .A1(n10932), .A2(n8668), .ZN(n6848) );
  AND2_X1 U8052 ( .A1(n9510), .A2(n8654), .ZN(n14624) );
  NAND2_X1 U8053 ( .A1(n8559), .A2(n8558), .ZN(n14093) );
  INV_X1 U8054 ( .A(n14044), .ZN(n14130) );
  MUX2_X1 U8055 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8243), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n8244) );
  AND2_X1 U8056 ( .A1(n7591), .A2(n7590), .ZN(n8129) );
  INV_X1 U8057 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U8058 ( .A1(n8622), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8620) );
  AND2_X1 U8059 ( .A1(n8086), .A2(n8091), .ZN(n11416) );
  NAND2_X1 U8060 ( .A1(n6886), .A2(n6884), .ZN(n8010) );
  INV_X1 U8061 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U8062 ( .A1(n7422), .A2(n7427), .ZN(n7937) );
  NAND2_X1 U8063 ( .A1(n7899), .A2(n7428), .ZN(n7422) );
  OR2_X1 U8064 ( .A1(n8316), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n8331) );
  INV_X1 U8065 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8313) );
  XNOR2_X1 U8066 ( .A(n7527), .B(SI_2_), .ZN(n7757) );
  INV_X1 U8067 ( .A(n7523), .ZN(n7251) );
  BUF_X1 U8068 ( .A(n8314), .Z(n6725) );
  NAND2_X1 U8069 ( .A1(n14295), .A2(n14294), .ZN(n7002) );
  NAND2_X1 U8070 ( .A1(n14301), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7026) );
  INV_X1 U8071 ( .A(n7026), .ZN(n7023) );
  OR2_X1 U8072 ( .A1(n14301), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7027) );
  NAND2_X1 U8073 ( .A1(n14474), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7015) );
  NAND2_X1 U8074 ( .A1(n7012), .A2(n7014), .ZN(n7011) );
  NAND2_X1 U8075 ( .A1(n7007), .A2(n7006), .ZN(n7005) );
  NAND2_X1 U8076 ( .A1(n14277), .A2(n6490), .ZN(n7004) );
  NAND2_X1 U8077 ( .A1(n6999), .A2(n14313), .ZN(n14318) );
  OAI21_X1 U8078 ( .B1(n14314), .B2(n14315), .A(P2_ADDR_REG_17__SCAN_IN), .ZN(
        n6999) );
  NAND2_X1 U8079 ( .A1(n11148), .A2(n11147), .ZN(n11146) );
  NAND2_X1 U8080 ( .A1(n6812), .A2(n6810), .ZN(n12024) );
  NAND2_X1 U8081 ( .A1(n7356), .A2(n7353), .ZN(n11662) );
  AND2_X1 U8082 ( .A1(n11663), .A2(n7355), .ZN(n7353) );
  NAND2_X1 U8083 ( .A1(n11310), .A2(n11309), .ZN(n11308) );
  AND3_X1 U8084 ( .A1(n9095), .A2(n9094), .A3(n9093), .ZN(n12441) );
  AND2_X1 U8085 ( .A1(n9166), .A2(n9165), .ZN(n12367) );
  OR2_X1 U8086 ( .A1(n9802), .A2(n12500), .ZN(n9803) );
  INV_X1 U8087 ( .A(n12379), .ZN(n12352) );
  INV_X1 U8088 ( .A(n7362), .ZN(n7360) );
  AND2_X1 U8089 ( .A1(n7362), .A2(n10365), .ZN(n7358) );
  NAND2_X1 U8090 ( .A1(n9090), .A2(n9089), .ZN(n12115) );
  OR2_X1 U8091 ( .A1(n9088), .A2(n10659), .ZN(n9089) );
  NAND2_X1 U8092 ( .A1(n9110), .A2(n9109), .ZN(n12406) );
  AND4_X1 U8093 ( .A1(n8959), .A2(n8958), .A3(n8957), .A4(n8956), .ZN(n14347)
         );
  AND4_X1 U8094 ( .A1(n9084), .A2(n9083), .A3(n9082), .A4(n9081), .ZN(n12427)
         );
  NAND2_X1 U8095 ( .A1(n9139), .A2(n9138), .ZN(n12364) );
  INV_X1 U8096 ( .A(n12441), .ZN(n12182) );
  INV_X1 U8097 ( .A(n12427), .ZN(n12452) );
  AOI21_X1 U8098 ( .B1(n10637), .B2(n10638), .A(n6862), .ZN(n10707) );
  AND2_X1 U8099 ( .A1(n10504), .A2(n10647), .ZN(n6862) );
  OAI22_X1 U8100 ( .A1(n10707), .A2(n10708), .B1(n10505), .B2(n10525), .ZN(
        n10621) );
  OR2_X1 U8101 ( .A1(n11227), .A2(n11228), .ZN(n6986) );
  OR2_X1 U8102 ( .A1(n12193), .A2(n12194), .ZN(n6993) );
  INV_X1 U8103 ( .A(n7050), .ZN(n12213) );
  INV_X1 U8104 ( .A(n7048), .ZN(n12234) );
  XNOR2_X1 U8105 ( .A(n12245), .B(n12260), .ZN(n12223) );
  OR2_X1 U8106 ( .A1(n12249), .A2(n12250), .ZN(n12282) );
  NAND2_X1 U8107 ( .A1(n7062), .A2(n7063), .ZN(n7061) );
  AND2_X1 U8108 ( .A1(n7068), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7063) );
  INV_X1 U8109 ( .A(n12321), .ZN(n6761) );
  NAND2_X1 U8110 ( .A1(n12315), .A2(n12314), .ZN(n6762) );
  NAND2_X1 U8111 ( .A1(n6879), .A2(n6613), .ZN(n6740) );
  NAND2_X1 U8112 ( .A1(n6880), .A2(n14922), .ZN(n6879) );
  OAI21_X1 U8113 ( .B1(n11883), .B2(n9305), .A(n9304), .ZN(n14355) );
  AND2_X1 U8114 ( .A1(n9254), .A2(n9253), .ZN(n12639) );
  NOR2_X1 U8115 ( .A1(n14374), .A2(n6771), .ZN(n7246) );
  INV_X1 U8116 ( .A(n7974), .ZN(n6771) );
  NOR2_X1 U8117 ( .A1(n12730), .A2(n13106), .ZN(n6924) );
  NAND2_X1 U8118 ( .A1(n9918), .A2(n7901), .ZN(n6928) );
  OAI21_X1 U8119 ( .B1(n13227), .B2(n8167), .A(n8100), .ZN(n12928) );
  NAND2_X1 U8120 ( .A1(n6655), .A2(n7832), .ZN(n13065) );
  AOI21_X1 U8121 ( .B1(n12785), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6656), .ZN(
        n6655) );
  NAND2_X1 U8122 ( .A1(n7831), .A2(n7830), .ZN(n6656) );
  CLKBUF_X2 U8123 ( .A(P2_U3947), .Z(n13071) );
  NAND2_X1 U8124 ( .A1(n10129), .A2(n10130), .ZN(n10210) );
  NOR2_X1 U8125 ( .A1(n11439), .A2(n11438), .ZN(n11738) );
  AND2_X1 U8126 ( .A1(n10089), .A2(n10060), .ZN(n14805) );
  NAND2_X1 U8127 ( .A1(n13307), .A2(n13288), .ZN(n6759) );
  INV_X1 U8128 ( .A(n11927), .ZN(n7106) );
  AND2_X1 U8129 ( .A1(n7710), .A2(n7709), .ZN(n13105) );
  OR2_X1 U8130 ( .A1(n13315), .A2(n13238), .ZN(n6660) );
  INV_X1 U8131 ( .A(n13118), .ZN(n6754) );
  NAND2_X1 U8132 ( .A1(n14835), .A2(n7686), .ZN(n13226) );
  OAI22_X1 U8133 ( .A1(n14828), .A2(P2_D_REG_1__SCAN_IN), .B1(n7662), .B2(
        n13461), .ZN(n14834) );
  OAI21_X1 U8134 ( .B1(n14828), .B2(P2_D_REG_0__SCAN_IN), .A(n7649), .ZN(
        n14831) );
  XNOR2_X1 U8135 ( .A(n7647), .B(n7646), .ZN(n13458) );
  INV_X1 U8136 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n7646) );
  OAI21_X1 U8137 ( .B1(n7645), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7647) );
  INV_X1 U8138 ( .A(n12979), .ZN(n13026) );
  XNOR2_X1 U8139 ( .A(n6689), .B(n13597), .ZN(n13598) );
  NAND2_X1 U8140 ( .A1(n13728), .A2(n13596), .ZN(n6689) );
  OR2_X1 U8141 ( .A1(n11557), .A2(n8312), .ZN(n8533) );
  NAND2_X1 U8142 ( .A1(n7261), .A2(n7259), .ZN(n10876) );
  NAND2_X1 U8143 ( .A1(n9674), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7261) );
  AND2_X1 U8144 ( .A1(n7262), .A2(n7260), .ZN(n7259) );
  NAND2_X1 U8145 ( .A1(n9921), .A2(n13823), .ZN(n7260) );
  NAND2_X1 U8146 ( .A1(n13617), .A2(n13542), .ZN(n13693) );
  NAND2_X1 U8147 ( .A1(n8430), .A2(n8429), .ZN(n11733) );
  INV_X1 U8148 ( .A(n13751), .ZN(n14395) );
  NAND2_X1 U8149 ( .A1(n8460), .A2(n8459), .ZN(n14439) );
  NAND2_X1 U8150 ( .A1(n7180), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U8151 ( .A1(n7180), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8564) );
  AOI22_X1 U8152 ( .A1(n7180), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n9659), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n8495) );
  NAND2_X1 U8153 ( .A1(n7180), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U8154 ( .A1(n8295), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n8284) );
  INV_X1 U8155 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7520) );
  AND2_X1 U8156 ( .A1(n6965), .A2(n6964), .ZN(n13838) );
  INV_X1 U8157 ( .A(n14576), .ZN(n14558) );
  NAND2_X1 U8158 ( .A1(n13873), .A2(n13872), .ZN(n14052) );
  AND2_X1 U8159 ( .A1(n13871), .A2(n14617), .ZN(n13872) );
  OR2_X1 U8160 ( .A1(n6477), .A2(n6956), .ZN(n13871) );
  NAND2_X1 U8161 ( .A1(n7185), .A2(n14057), .ZN(n7266) );
  OAI211_X1 U8162 ( .C1(n13877), .C2(n6834), .A(n6832), .B(n6830), .ZN(n7184)
         );
  OR2_X1 U8163 ( .A1(n9703), .A2(n14608), .ZN(n6834) );
  AND2_X1 U8164 ( .A1(n6833), .A2(n6608), .ZN(n6832) );
  NAND2_X1 U8165 ( .A1(n6686), .A2(n6549), .ZN(n6685) );
  NAND2_X1 U8166 ( .A1(n8616), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8510) );
  NAND2_X1 U8167 ( .A1(n7007), .A2(n7009), .ZN(n7013) );
  AND2_X1 U8168 ( .A1(n7008), .A2(n7013), .ZN(n14482) );
  NAND2_X1 U8169 ( .A1(n14277), .A2(n14810), .ZN(n7008) );
  INV_X1 U8170 ( .A(n14481), .ZN(n7012) );
  MUX2_X1 U8171 ( .A(n10264), .B(n13780), .S(n9541), .Z(n9520) );
  NAND2_X1 U8172 ( .A1(n6569), .A2(n6489), .ZN(n6668) );
  NAND2_X1 U8173 ( .A1(n7226), .A2(n12834), .ZN(n7225) );
  NAND2_X1 U8174 ( .A1(n6678), .A2(n7499), .ZN(n9544) );
  NAND2_X1 U8175 ( .A1(n9539), .A2(n7500), .ZN(n7499) );
  OR2_X1 U8176 ( .A1(n9359), .A2(n9230), .ZN(n9360) );
  NAND2_X1 U8177 ( .A1(n12848), .A2(n7214), .ZN(n7213) );
  NAND2_X1 U8178 ( .A1(n12851), .A2(n7215), .ZN(n7214) );
  NAND2_X1 U8179 ( .A1(n9551), .A2(n9554), .ZN(n7466) );
  NAND2_X1 U8180 ( .A1(n6715), .A2(n6714), .ZN(n9367) );
  NAND2_X1 U8181 ( .A1(n9184), .A2(n6717), .ZN(n6714) );
  NAND2_X1 U8182 ( .A1(n6903), .A2(n6902), .ZN(n12867) );
  NAND2_X1 U8183 ( .A1(n12862), .A2(n12864), .ZN(n6902) );
  AND2_X1 U8184 ( .A1(n9562), .A2(n6675), .ZN(n6674) );
  INV_X1 U8185 ( .A(n9560), .ZN(n6675) );
  NAND2_X1 U8186 ( .A1(n12874), .A2(n7222), .ZN(n7221) );
  NAND2_X1 U8187 ( .A1(n12867), .A2(n12868), .ZN(n6901) );
  AOI21_X1 U8188 ( .B1(n9572), .B2(n9573), .A(n6734), .ZN(n6769) );
  AND2_X1 U8189 ( .A1(n12891), .A2(n12907), .ZN(n12908) );
  NOR2_X1 U8190 ( .A1(n7498), .A2(n7497), .ZN(n7496) );
  INV_X1 U8191 ( .A(n9590), .ZN(n7497) );
  INV_X1 U8192 ( .A(n9589), .ZN(n7498) );
  NOR2_X1 U8193 ( .A1(n6595), .A2(n9684), .ZN(n7493) );
  INV_X1 U8194 ( .A(n9592), .ZN(n7492) );
  AOI21_X1 U8195 ( .B1(n9607), .B2(n9606), .A(n9604), .ZN(n7490) );
  OR2_X1 U8196 ( .A1(n7205), .A2(n12926), .ZN(n6913) );
  INV_X1 U8197 ( .A(n12929), .ZN(n7230) );
  INV_X1 U8198 ( .A(n12930), .ZN(n7229) );
  NAND2_X1 U8199 ( .A1(n7489), .A2(n7488), .ZN(n9609) );
  AND2_X1 U8200 ( .A1(n9610), .A2(n6570), .ZN(n7488) );
  NAND2_X1 U8201 ( .A1(n7489), .A2(n6570), .ZN(n9612) );
  NAND2_X1 U8202 ( .A1(n6745), .A2(n7218), .ZN(n12943) );
  OR2_X1 U8203 ( .A1(n7219), .A2(n12940), .ZN(n7218) );
  INV_X1 U8204 ( .A(n12939), .ZN(n7219) );
  AND2_X1 U8205 ( .A1(n12944), .A2(n6912), .ZN(n6911) );
  INV_X1 U8206 ( .A(n12942), .ZN(n6912) );
  NAND2_X1 U8207 ( .A1(n12945), .A2(n12942), .ZN(n6910) );
  OAI21_X1 U8208 ( .B1(n6673), .B2(n6671), .A(n7484), .ZN(n9623) );
  NAND2_X1 U8209 ( .A1(n9618), .A2(n9620), .ZN(n7484) );
  AOI21_X1 U8210 ( .B1(n9616), .B2(n6672), .A(n9615), .ZN(n6673) );
  OAI21_X1 U8211 ( .B1(n9616), .B2(n6672), .A(n6491), .ZN(n6671) );
  AOI22_X1 U8212 ( .A1(n12344), .A2(n9471), .B1(n9470), .B2(n12523), .ZN(n9476) );
  OAI21_X1 U8213 ( .B1(n11089), .B2(n7122), .A(n14965), .ZN(n7121) );
  NAND2_X1 U8214 ( .A1(n15036), .A2(n9188), .ZN(n9373) );
  AOI21_X1 U8215 ( .B1(n6923), .B2(n7231), .A(n6480), .ZN(n6922) );
  NAND2_X1 U8216 ( .A1(n12806), .A2(n12805), .ZN(n6691) );
  INV_X1 U8217 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7614) );
  INV_X1 U8218 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7615) );
  INV_X1 U8219 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6654) );
  NAND2_X1 U8220 ( .A1(n9629), .A2(n9631), .ZN(n7481) );
  INV_X1 U8221 ( .A(n8011), .ZN(n6694) );
  OAI21_X1 U8222 ( .B1(n7533), .B2(n7419), .A(n7536), .ZN(n7414) );
  NOR2_X1 U8223 ( .A1(n7419), .A2(n7417), .ZN(n7416) );
  INV_X1 U8224 ( .A(n7532), .ZN(n7417) );
  OAI21_X1 U8225 ( .B1(n9926), .B2(n9934), .A(n6729), .ZN(n7531) );
  NAND2_X1 U8226 ( .A1(n9926), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6729) );
  INV_X1 U8227 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6893) );
  NAND2_X1 U8228 ( .A1(n14183), .A2(n14184), .ZN(n14185) );
  NOR2_X1 U8229 ( .A1(n6815), .A2(n9797), .ZN(n6814) );
  INV_X1 U8230 ( .A(n7519), .ZN(n6815) );
  NAND2_X1 U8231 ( .A1(n6802), .A2(n6800), .ZN(n9816) );
  AOI21_X1 U8232 ( .B1(n6803), .B2(n6808), .A(n6801), .ZN(n6800) );
  NOR2_X1 U8233 ( .A1(n7342), .A2(n6804), .ZN(n6803) );
  OR2_X1 U8234 ( .A1(n9790), .A2(n12140), .ZN(n9791) );
  INV_X1 U8235 ( .A(n10743), .ZN(n6788) );
  NAND2_X1 U8236 ( .A1(n9335), .A2(n11952), .ZN(n7326) );
  INV_X1 U8237 ( .A(n9485), .ZN(n9316) );
  NOR2_X1 U8238 ( .A1(n6485), .A2(n10526), .ZN(n7059) );
  INV_X1 U8239 ( .A(n7058), .ZN(n7057) );
  OAI21_X1 U8240 ( .B1(n10715), .B2(n6485), .A(n10526), .ZN(n7058) );
  OAI21_X1 U8241 ( .B1(n10639), .B2(n6562), .A(n6987), .ZN(n10512) );
  AND2_X1 U8242 ( .A1(n11531), .A2(n11530), .ZN(n11609) );
  NAND2_X1 U8243 ( .A1(n7048), .A2(n12235), .ZN(n12259) );
  OR2_X1 U8244 ( .A1(n12281), .A2(n12303), .ZN(n6984) );
  INV_X1 U8245 ( .A(n12250), .ZN(n6981) );
  INV_X1 U8246 ( .A(n12263), .ZN(n7069) );
  INV_X1 U8247 ( .A(n12417), .ZN(n9215) );
  NAND2_X1 U8248 ( .A1(n9401), .A2(n9402), .ZN(n7141) );
  INV_X1 U8249 ( .A(n9406), .ZN(n7137) );
  INV_X1 U8250 ( .A(n9402), .ZN(n7138) );
  NAND2_X1 U8251 ( .A1(n6629), .A2(n9353), .ZN(n12394) );
  INV_X1 U8252 ( .A(n12639), .ZN(n10284) );
  NAND2_X1 U8253 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n11814), .ZN(n8739) );
  INV_X1 U8254 ( .A(n9054), .ZN(n7312) );
  INV_X1 U8255 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7125) );
  INV_X1 U8256 ( .A(n8971), .ZN(n7124) );
  NOR2_X1 U8257 ( .A1(n8018), .A2(n8017), .ZN(n8016) );
  AND2_X1 U8258 ( .A1(n7909), .A2(n7688), .ZN(n7948) );
  AND2_X1 U8259 ( .A1(n7897), .A2(n10921), .ZN(n7247) );
  AND2_X1 U8260 ( .A1(n8016), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8032) );
  NOR2_X1 U8261 ( .A1(n6742), .A2(n12791), .ZN(n12978) );
  NAND2_X1 U8262 ( .A1(n6733), .A2(n6732), .ZN(n12803) );
  INV_X1 U8263 ( .A(n13152), .ZN(n7157) );
  NOR2_X1 U8264 ( .A1(n12946), .A2(n7046), .ZN(n7045) );
  INV_X1 U8265 ( .A(n7047), .ZN(n7046) );
  INV_X1 U8266 ( .A(n11896), .ZN(n7168) );
  NOR2_X1 U8267 ( .A1(n13179), .A2(n7167), .ZN(n7166) );
  NOR2_X1 U8268 ( .A1(n13201), .A2(n7168), .ZN(n7167) );
  NOR2_X1 U8269 ( .A1(n13182), .A2(n13194), .ZN(n7047) );
  AOI21_X1 U8270 ( .B1(n11919), .B2(n11920), .A(n7094), .ZN(n7093) );
  INV_X1 U8271 ( .A(n12989), .ZN(n7094) );
  INV_X1 U8272 ( .A(n11920), .ZN(n7091) );
  NAND2_X1 U8273 ( .A1(n6639), .A2(n6637), .ZN(n6641) );
  AND2_X1 U8274 ( .A1(n6589), .A2(n6638), .ZN(n6637) );
  OR2_X1 U8275 ( .A1(n13002), .A2(n7151), .ZN(n7150) );
  INV_X1 U8276 ( .A(n10968), .ZN(n7151) );
  INV_X1 U8277 ( .A(n10957), .ZN(n7087) );
  NAND2_X1 U8278 ( .A1(n11179), .A2(n11363), .ZN(n11300) );
  NOR2_X1 U8279 ( .A1(n11037), .A2(n14892), .ZN(n11179) );
  NOR2_X1 U8280 ( .A1(n7678), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6646) );
  NOR2_X1 U8281 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7758) );
  INV_X1 U8282 ( .A(n13502), .ZN(n7389) );
  NOR2_X1 U8283 ( .A1(n9703), .A2(n7455), .ZN(n7454) );
  NAND2_X1 U8284 ( .A1(n13879), .A2(n7456), .ZN(n7455) );
  AND2_X1 U8285 ( .A1(n9702), .A2(n13907), .ZN(n7456) );
  XNOR2_X1 U8286 ( .A(n13870), .B(n13753), .ZN(n7453) );
  NAND2_X1 U8287 ( .A1(n7478), .A2(n7474), .ZN(n7473) );
  INV_X1 U8288 ( .A(n7477), .ZN(n7474) );
  AND2_X1 U8289 ( .A1(n9643), .A2(n7479), .ZN(n7477) );
  AOI21_X1 U8290 ( .B1(n13849), .B2(P1_REG1_REG_17__SCAN_IN), .A(n14562), .ZN(
        n13851) );
  NOR2_X1 U8291 ( .A1(n14087), .A2(n6952), .ZN(n6951) );
  INV_X1 U8292 ( .A(n6953), .ZN(n6952) );
  NOR2_X1 U8293 ( .A1(n14093), .A2(n6828), .ZN(n6953) );
  AOI21_X1 U8294 ( .B1(n11472), .B2(n7258), .A(n7257), .ZN(n7256) );
  INV_X1 U8295 ( .A(n8676), .ZN(n7257) );
  INV_X1 U8296 ( .A(n8675), .ZN(n7258) );
  NOR2_X1 U8297 ( .A1(n14453), .A2(n11381), .ZN(n6962) );
  INV_X1 U8298 ( .A(n8384), .ZN(n7173) );
  AND2_X1 U8299 ( .A1(n9521), .A2(n8278), .ZN(n7177) );
  NAND2_X1 U8300 ( .A1(n9686), .A2(n9521), .ZN(n7175) );
  INV_X1 U8301 ( .A(n6950), .ZN(n14022) );
  NAND2_X1 U8302 ( .A1(n8239), .A2(n7487), .ZN(n7486) );
  XNOR2_X1 U8303 ( .A(n9650), .B(SI_29_), .ZN(n9648) );
  INV_X1 U8304 ( .A(n6706), .ZN(n6705) );
  OAI21_X1 U8305 ( .B1(n7597), .B2(n6609), .A(n7602), .ZN(n6706) );
  NAND2_X1 U8306 ( .A1(n8158), .A2(n7597), .ZN(n8161) );
  NAND2_X1 U8307 ( .A1(n6757), .A2(n7588), .ZN(n6765) );
  NAND2_X1 U8308 ( .A1(n8106), .A2(n7587), .ZN(n6757) );
  OR2_X1 U8309 ( .A1(n7580), .A2(n7579), .ZN(n7581) );
  AND2_X1 U8310 ( .A1(n8507), .A2(n8509), .ZN(n7501) );
  AOI21_X1 U8311 ( .B1(n6888), .B2(n6890), .A(n6885), .ZN(n6884) );
  INV_X1 U8312 ( .A(n7564), .ZN(n6885) );
  AOI21_X1 U8313 ( .B1(n7900), .B2(n7428), .A(n6565), .ZN(n7427) );
  INV_X1 U8314 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8332) );
  XNOR2_X1 U8315 ( .A(n7541), .B(SI_6_), .ZN(n7822) );
  NAND2_X1 U8316 ( .A1(n6772), .A2(n6731), .ZN(n7523) );
  OR2_X1 U8317 ( .A1(n7522), .A2(n9898), .ZN(n6772) );
  XNOR2_X1 U8318 ( .A(n14181), .B(n7029), .ZN(n14240) );
  INV_X1 U8319 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7029) );
  XNOR2_X1 U8320 ( .A(n14185), .B(n7000), .ZN(n14228) );
  INV_X1 U8321 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7000) );
  AOI21_X1 U8322 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14199), .A(n14198), .ZN(
        n14200) );
  AND2_X1 U8323 ( .A1(n14267), .A2(n14266), .ZN(n14198) );
  NOR2_X1 U8324 ( .A1(n6478), .A2(n14478), .ZN(n7006) );
  NAND2_X1 U8325 ( .A1(n9821), .A2(n9820), .ZN(n7339) );
  NAND2_X1 U8326 ( .A1(n9788), .A2(n11312), .ZN(n7355) );
  OR2_X1 U8327 ( .A1(n8822), .A2(n8798), .ZN(n8799) );
  INV_X1 U8328 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8910) );
  AND2_X1 U8329 ( .A1(n12074), .A2(n9827), .ZN(n12101) );
  NAND2_X1 U8330 ( .A1(n9823), .A2(n9822), .ZN(n12100) );
  NOR2_X1 U8331 ( .A1(n9132), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U8332 ( .A1(n9777), .A2(n12190), .ZN(n7362) );
  INV_X1 U8333 ( .A(n12043), .ZN(n6808) );
  NAND2_X1 U8334 ( .A1(n11662), .A2(n9791), .ZN(n12059) );
  AND2_X1 U8335 ( .A1(n9860), .A2(n9859), .ZN(n12170) );
  OR2_X1 U8336 ( .A1(n10446), .A2(n15082), .ZN(n10448) );
  OR2_X1 U8337 ( .A1(n10442), .A2(n15049), .ZN(n10443) );
  NAND2_X1 U8338 ( .A1(n10443), .A2(n10406), .ZN(n10407) );
  NAND2_X1 U8339 ( .A1(n10398), .A2(n10397), .ZN(n10521) );
  OR2_X1 U8340 ( .A1(n10641), .A2(n15085), .ZN(n10717) );
  NAND2_X1 U8341 ( .A1(n10524), .A2(n10715), .ZN(n10719) );
  OR2_X1 U8342 ( .A1(n10524), .A2(n7056), .ZN(n7052) );
  INV_X1 U8343 ( .A(n7059), .ZN(n7056) );
  AOI22_X1 U8344 ( .A1(n7057), .A2(n6485), .B1(n7059), .B2(n7055), .ZN(n7054)
         );
  OR2_X1 U8345 ( .A1(n8857), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U8346 ( .A1(n7053), .A2(n7057), .ZN(n10529) );
  OR2_X1 U8347 ( .A1(n10524), .A2(n6485), .ZN(n7053) );
  OR2_X1 U8348 ( .A1(n10625), .A2(n14997), .ZN(n10623) );
  NAND2_X1 U8349 ( .A1(n6996), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6995) );
  NAND2_X1 U8350 ( .A1(n6997), .A2(n11059), .ZN(n6996) );
  INV_X1 U8351 ( .A(n10664), .ZN(n6997) );
  AND2_X1 U8352 ( .A1(n6995), .A2(n6994), .ZN(n14933) );
  NOR2_X1 U8353 ( .A1(n14932), .A2(n14933), .ZN(n14931) );
  AND2_X1 U8354 ( .A1(n7077), .A2(n7078), .ZN(n14936) );
  AND2_X1 U8355 ( .A1(n11518), .A2(n11517), .ZN(n11603) );
  XNOR2_X1 U8356 ( .A(n11609), .B(n11610), .ZN(n11532) );
  OAI21_X1 U8357 ( .B1(n11789), .B2(n11790), .A(n11791), .ZN(n11792) );
  NOR2_X1 U8358 ( .A1(n11792), .A2(n11793), .ZN(n12200) );
  AND2_X1 U8359 ( .A1(n11780), .A2(n11779), .ZN(n12192) );
  NAND2_X1 U8360 ( .A1(n6763), .A2(n6507), .ZN(n7050) );
  NOR2_X1 U8361 ( .A1(n12575), .A2(n12236), .ZN(n12261) );
  OR2_X1 U8362 ( .A1(n7069), .A2(n7067), .ZN(n7062) );
  OR2_X1 U8363 ( .A1(n12271), .A2(n12303), .ZN(n7068) );
  OAI21_X1 U8364 ( .B1(n6874), .B2(n6876), .A(n6873), .ZN(n12277) );
  NAND2_X1 U8365 ( .A1(n6618), .A2(n12230), .ZN(n6876) );
  NOR2_X1 U8366 ( .A1(n12305), .A2(n12304), .ZN(n12308) );
  XNOR2_X1 U8367 ( .A(n6881), .B(n12322), .ZN(n6880) );
  INV_X1 U8368 ( .A(n12323), .ZN(n6881) );
  NOR2_X1 U8369 ( .A1(n11247), .A2(n10459), .ZN(n6882) );
  INV_X1 U8370 ( .A(n9745), .ZN(n9752) );
  NOR2_X1 U8371 ( .A1(n7132), .A2(n7129), .ZN(n7128) );
  OAI21_X1 U8372 ( .B1(n7130), .B2(n7129), .A(n9342), .ZN(n7127) );
  INV_X1 U8373 ( .A(n9343), .ZN(n7129) );
  OR2_X1 U8374 ( .A1(n9161), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U8375 ( .A1(n9112), .A2(n9111), .ZN(n9121) );
  NOR2_X1 U8376 ( .A1(n9091), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9102) );
  NAND2_X1 U8377 ( .A1(n6747), .A2(n7448), .ZN(n12438) );
  AOI21_X1 U8378 ( .B1(n6475), .B2(n12470), .A(n6554), .ZN(n7448) );
  NAND2_X1 U8379 ( .A1(n6748), .A2(n6475), .ZN(n6747) );
  AND2_X1 U8380 ( .A1(n9048), .A2(n9047), .ZN(n9063) );
  NAND2_X1 U8381 ( .A1(n9063), .A2(n9062), .ZN(n9079) );
  AOI21_X1 U8382 ( .B1(n7110), .B2(n9430), .A(n6547), .ZN(n7108) );
  INV_X1 U8383 ( .A(n7111), .ZN(n7110) );
  NAND2_X1 U8384 ( .A1(n6749), .A2(n9209), .ZN(n12477) );
  OR2_X1 U8385 ( .A1(n9015), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9035) );
  CLKBUF_X1 U8386 ( .A(n12494), .Z(n6749) );
  AOI21_X1 U8387 ( .B1(n7115), .B2(n7117), .A(n7113), .ZN(n7112) );
  INV_X1 U8388 ( .A(n9417), .ZN(n7113) );
  OR2_X1 U8389 ( .A1(n8979), .A2(n8765), .ZN(n8988) );
  OAI21_X1 U8390 ( .B1(n11455), .B2(n7139), .A(n7136), .ZN(n11509) );
  INV_X1 U8391 ( .A(n7140), .ZN(n7139) );
  AOI21_X1 U8392 ( .B1(n7140), .B2(n7138), .A(n7137), .ZN(n7136) );
  AND2_X1 U8393 ( .A1(n9325), .A2(n7141), .ZN(n7140) );
  AND2_X1 U8394 ( .A1(n8911), .A2(n8910), .ZN(n8929) );
  NAND2_X1 U8395 ( .A1(n9199), .A2(n9198), .ZN(n11199) );
  NOR2_X1 U8396 ( .A1(n8894), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8911) );
  NAND2_X1 U8397 ( .A1(n11092), .A2(n9391), .ZN(n14964) );
  NAND2_X1 U8398 ( .A1(n11090), .A2(n11089), .ZN(n11092) );
  INV_X1 U8399 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n10626) );
  AND4_X1 U8400 ( .A1(n8884), .A2(n8883), .A3(n8882), .A4(n8881), .ZN(n14987)
         );
  CLKBUF_X1 U8401 ( .A(n14979), .Z(n15003) );
  INV_X1 U8402 ( .A(n9366), .ZN(n15015) );
  NAND2_X1 U8403 ( .A1(n9288), .A2(n9287), .ZN(n9313) );
  NAND2_X1 U8404 ( .A1(n7126), .A2(n7130), .ZN(n9289) );
  NAND2_X1 U8405 ( .A1(n12354), .A2(n7133), .ZN(n7126) );
  NAND2_X1 U8406 ( .A1(n12443), .A2(n9449), .ZN(n12430) );
  NAND2_X1 U8407 ( .A1(n9014), .A2(n9013), .ZN(n12166) );
  NAND2_X1 U8408 ( .A1(n15043), .A2(n15052), .ZN(n14362) );
  AND3_X1 U8409 ( .A1(n10284), .A2(n9770), .A3(n9758), .ZN(n9854) );
  INV_X1 U8410 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8767) );
  AND2_X1 U8411 ( .A1(n14164), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7319) );
  NAND2_X1 U8412 ( .A1(n6751), .A2(n8762), .ZN(n6856) );
  NAND2_X1 U8413 ( .A1(n7124), .A2(n6859), .ZN(n6858) );
  NOR2_X1 U8414 ( .A1(n7123), .A2(n8762), .ZN(n6859) );
  INV_X1 U8415 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7460) );
  AND2_X1 U8416 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n6860) );
  NAND2_X1 U8417 ( .A1(n9241), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9246) );
  XNOR2_X1 U8418 ( .A(n9257), .B(n9256), .ZN(n10388) );
  OAI21_X1 U8419 ( .B1(n9255), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9257) );
  OR2_X1 U8420 ( .A1(n9175), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n9177) );
  NAND2_X1 U8421 ( .A1(n9171), .A2(n9170), .ZN(n9255) );
  INV_X1 U8422 ( .A(n9177), .ZN(n9171) );
  INV_X1 U8423 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7364) );
  NAND2_X1 U8424 ( .A1(n9026), .A2(n7365), .ZN(n9056) );
  INV_X1 U8425 ( .A(n7298), .ZN(n7297) );
  AND2_X1 U8426 ( .A1(n8995), .A2(n9010), .ZN(n9026) );
  NAND2_X1 U8427 ( .A1(n7124), .A2(n8751), .ZN(n8973) );
  NOR2_X1 U8428 ( .A1(n7288), .A2(n6564), .ZN(n7287) );
  OR2_X1 U8429 ( .A1(n8919), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8920) );
  NOR2_X1 U8430 ( .A1(n8920), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8950) );
  XNOR2_X1 U8431 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8854) );
  INV_X1 U8432 ( .A(n13065), .ZN(n10800) );
  OR2_X1 U8433 ( .A1(n7845), .A2(n7844), .ZN(n7867) );
  OR2_X1 U8434 ( .A1(n7867), .A2(n13073), .ZN(n7886) );
  OR2_X1 U8435 ( .A1(n8074), .A2(n8073), .ZN(n8095) );
  NAND2_X1 U8436 ( .A1(n10052), .A2(n10058), .ZN(n12773) );
  INV_X1 U8437 ( .A(n7898), .ZN(n6936) );
  OR2_X1 U8438 ( .A1(n7917), .A2(n7916), .ZN(n6939) );
  INV_X1 U8439 ( .A(n7247), .ZN(n6934) );
  AND2_X1 U8440 ( .A1(n8067), .A2(n8043), .ZN(n7249) );
  CLKBUF_X1 U8441 ( .A(n10795), .Z(n10796) );
  OR2_X1 U8442 ( .A1(n7983), .A2(n7982), .ZN(n8000) );
  AND3_X1 U8443 ( .A1(n8004), .A2(n8003), .A3(n8002), .ZN(n12887) );
  NAND2_X1 U8444 ( .A1(n12786), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7084) );
  AND4_X1 U8445 ( .A1(n6652), .A2(n7763), .A3(n7762), .A4(n6651), .ZN(n10575)
         );
  NAND2_X1 U8446 ( .A1(n7745), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6652) );
  AND2_X1 U8447 ( .A1(n11929), .A2(n13449), .ZN(n7746) );
  NAND2_X1 U8448 ( .A1(n14754), .A2(n10081), .ZN(n10135) );
  NAND2_X1 U8449 ( .A1(n10135), .A2(n10136), .ZN(n10134) );
  NAND2_X1 U8450 ( .A1(n10540), .A2(n10539), .ZN(n10541) );
  NOR2_X1 U8451 ( .A1(n10541), .A2(n10542), .ZN(n11107) );
  INV_X1 U8452 ( .A(n13308), .ZN(n12796) );
  AND2_X1 U8453 ( .A1(n8209), .A2(n8208), .ZN(n12957) );
  AND2_X1 U8454 ( .A1(n13112), .A2(n13101), .ZN(n7161) );
  AND2_X1 U8455 ( .A1(n7153), .A2(n6503), .ZN(n13116) );
  AND2_X1 U8456 ( .A1(n7720), .A2(n7719), .ZN(n13135) );
  NAND2_X1 U8457 ( .A1(n13211), .A2(n7045), .ZN(n13168) );
  NAND2_X1 U8458 ( .A1(n13164), .A2(n13163), .ZN(n13162) );
  NAND2_X1 U8459 ( .A1(n7103), .A2(n11924), .ZN(n6898) );
  NAND2_X1 U8460 ( .A1(n13200), .A2(n13201), .ZN(n13199) );
  NAND2_X1 U8461 ( .A1(n13211), .A2(n13416), .ZN(n13191) );
  NOR2_X1 U8462 ( .A1(n13269), .A2(n7040), .ZN(n7038) );
  NAND2_X1 U8463 ( .A1(n11654), .A2(n6482), .ZN(n13286) );
  NAND2_X1 U8464 ( .A1(n6476), .A2(n13013), .ZN(n11889) );
  AOI21_X1 U8465 ( .B1(n7144), .B2(n7146), .A(n6513), .ZN(n7142) );
  INV_X1 U8466 ( .A(n7144), .ZN(n7143) );
  NAND2_X1 U8467 ( .A1(n6736), .A2(n13007), .ZN(n11293) );
  NAND2_X1 U8468 ( .A1(n6661), .A2(n11178), .ZN(n11298) );
  NAND2_X1 U8469 ( .A1(n11177), .A2(n11176), .ZN(n6661) );
  INV_X1 U8470 ( .A(n13005), .ZN(n11176) );
  NAND2_X1 U8471 ( .A1(n7037), .A2(n7036), .ZN(n11037) );
  OAI21_X1 U8472 ( .B1(n10956), .B2(n7085), .A(n6663), .ZN(n11133) );
  INV_X1 U8473 ( .A(n7086), .ZN(n7085) );
  AOI21_X1 U8474 ( .B1(n6462), .B2(n7086), .A(n6518), .ZN(n6663) );
  NOR2_X1 U8475 ( .A1(n10958), .A2(n7087), .ZN(n7086) );
  NOR2_X1 U8476 ( .A1(n10606), .A2(n12849), .ZN(n11283) );
  OR2_X1 U8477 ( .A1(n10771), .A2(n12841), .ZN(n10606) );
  OAI21_X1 U8478 ( .B1(n6636), .B2(n12996), .A(n6633), .ZN(n10592) );
  AOI21_X1 U8479 ( .B1(n10765), .B2(n6634), .A(n6552), .ZN(n6633) );
  INV_X1 U8480 ( .A(n10567), .ZN(n6634) );
  NAND2_X1 U8481 ( .A1(n10772), .A2(n14860), .ZN(n10771) );
  INV_X1 U8482 ( .A(n12992), .ZN(n10837) );
  NAND2_X1 U8483 ( .A1(n7760), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7035) );
  NAND2_X1 U8484 ( .A1(n8070), .A2(n10078), .ZN(n7034) );
  AND2_X1 U8485 ( .A1(n10355), .A2(n7033), .ZN(n10840) );
  NAND2_X1 U8486 ( .A1(n12991), .A2(n10348), .ZN(n10574) );
  CLKBUF_X1 U8487 ( .A(n12991), .Z(n6735) );
  INV_X1 U8488 ( .A(n13198), .ZN(n13281) );
  NAND2_X1 U8489 ( .A1(n13441), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6653) );
  AND2_X1 U8490 ( .A1(n8013), .A2(n8028), .ZN(n11739) );
  OR2_X1 U8491 ( .A1(n7978), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7996) );
  AND2_X1 U8492 ( .A1(n7920), .A2(n7906), .ZN(n10237) );
  INV_X1 U8493 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n7824) );
  AND2_X1 U8494 ( .A1(n7789), .A2(n7788), .ZN(n10086) );
  OR2_X1 U8495 ( .A1(n8447), .A2(n8252), .ZN(n8461) );
  INV_X1 U8496 ( .A(n13491), .ZN(n7393) );
  NAND2_X1 U8497 ( .A1(n13487), .A2(n13486), .ZN(n7394) );
  AND2_X1 U8498 ( .A1(n8695), .A2(n8599), .ZN(n13633) );
  NAND2_X1 U8499 ( .A1(n13693), .A2(n13692), .ZN(n7401) );
  NOR2_X1 U8500 ( .A1(n8403), .A2(n8402), .ZN(n8418) );
  NOR2_X1 U8501 ( .A1(n8461), .A2(n15104), .ZN(n8475) );
  NAND2_X1 U8502 ( .A1(n7408), .A2(n7407), .ZN(n13674) );
  INV_X1 U8503 ( .A(n13663), .ZN(n7407) );
  INV_X1 U8504 ( .A(n13662), .ZN(n7408) );
  AND2_X1 U8505 ( .A1(n8475), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8492) );
  NAND2_X1 U8506 ( .A1(n8290), .A2(n9890), .ZN(n7262) );
  OR2_X1 U8507 ( .A1(n8378), .A2(n8377), .ZN(n8390) );
  OAI21_X1 U8508 ( .B1(n13693), .B2(n7399), .A(n7395), .ZN(n6690) );
  AOI21_X1 U8509 ( .B1(n7398), .B2(n7397), .A(n7396), .ZN(n7395) );
  INV_X1 U8510 ( .A(n13692), .ZN(n7397) );
  OR2_X1 U8511 ( .A1(n10014), .A2(n13783), .ZN(n14385) );
  INV_X1 U8512 ( .A(n7409), .ZN(n7406) );
  AOI21_X1 U8513 ( .B1(n7409), .B2(n7405), .A(n7404), .ZN(n7403) );
  INV_X1 U8514 ( .A(n13528), .ZN(n7404) );
  INV_X1 U8515 ( .A(n10894), .ZN(n7366) );
  INV_X1 U8516 ( .A(n9727), .ZN(n9728) );
  OR2_X1 U8517 ( .A1(n9641), .A2(n6526), .ZN(n6664) );
  OR2_X1 U8518 ( .A1(n9642), .A2(n6526), .ZN(n6665) );
  NAND2_X1 U8519 ( .A1(n9637), .A2(n9638), .ZN(n9636) );
  NAND2_X1 U8520 ( .A1(n7180), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8499) );
  INV_X1 U8521 ( .A(n8606), .ZN(n8530) );
  NAND2_X1 U8522 ( .A1(n7180), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8356) );
  AND2_X1 U8523 ( .A1(n6969), .A2(n6968), .ZN(n13815) );
  NAND2_X1 U8524 ( .A1(n13805), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6968) );
  INV_X1 U8525 ( .A(n6720), .ZN(n13784) );
  NOR2_X1 U8526 ( .A1(n10435), .A2(n10434), .ZN(n10733) );
  AND2_X1 U8527 ( .A1(n11430), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6973) );
  NAND2_X1 U8528 ( .A1(n11421), .A2(n11422), .ZN(n11857) );
  AND2_X1 U8529 ( .A1(n11865), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6976) );
  AOI21_X1 U8530 ( .B1(n11865), .B2(P1_REG1_REG_13__SCAN_IN), .A(n14510), .ZN(
        n14532) );
  AND2_X1 U8531 ( .A1(n13828), .A2(n13829), .ZN(n7503) );
  AND2_X1 U8532 ( .A1(n6958), .A2(n6956), .ZN(n6955) );
  NAND2_X1 U8533 ( .A1(n6843), .A2(n6846), .ZN(n13922) );
  NAND3_X1 U8534 ( .A1(n6951), .A2(n13988), .A3(n13660), .ZN(n13929) );
  NAND2_X1 U8535 ( .A1(n6951), .A2(n13988), .ZN(n13946) );
  NAND2_X1 U8536 ( .A1(n13988), .A2(n14101), .ZN(n13974) );
  NAND2_X1 U8537 ( .A1(n6950), .A2(n6949), .ZN(n14009) );
  INV_X1 U8538 ( .A(n14113), .ZN(n6949) );
  NAND2_X1 U8539 ( .A1(n6824), .A2(n9600), .ZN(n14001) );
  NOR2_X1 U8540 ( .A1(n14019), .A2(n6826), .ZN(n6825) );
  INV_X1 U8541 ( .A(n9595), .ZN(n6826) );
  OR2_X1 U8542 ( .A1(n14439), .A2(n14416), .ZN(n11772) );
  OAI21_X1 U8543 ( .B1(n11342), .B2(n9694), .A(n7256), .ZN(n14402) );
  AND2_X1 U8544 ( .A1(n6487), .A2(n11001), .ZN(n11475) );
  NAND2_X1 U8545 ( .A1(n11001), .A2(n6962), .ZN(n11351) );
  NAND2_X1 U8546 ( .A1(n10999), .A2(n8671), .ZN(n11215) );
  NAND2_X1 U8547 ( .A1(n11215), .A2(n11214), .ZN(n11213) );
  NAND2_X1 U8548 ( .A1(n11001), .A2(n14718), .ZN(n11219) );
  NOR2_X1 U8549 ( .A1(n10854), .A2(n10901), .ZN(n14600) );
  CLKBUF_X1 U8550 ( .A(n10817), .Z(n10818) );
  NAND2_X1 U8551 ( .A1(n8291), .A2(n6724), .ZN(n10476) );
  AND2_X1 U8552 ( .A1(n8292), .A2(n6517), .ZN(n6724) );
  NAND2_X1 U8553 ( .A1(n6821), .A2(n8655), .ZN(n10374) );
  NAND2_X1 U8554 ( .A1(n14606), .A2(n9686), .ZN(n6821) );
  NAND2_X1 U8555 ( .A1(n9512), .A2(n9510), .ZN(n14606) );
  INV_X1 U8556 ( .A(n9686), .ZN(n14605) );
  INV_X1 U8557 ( .A(n14385), .ZN(n13732) );
  AND2_X1 U8558 ( .A1(n13888), .A2(n6522), .ZN(n14060) );
  INV_X1 U8559 ( .A(n14675), .ZN(n14617) );
  NAND2_X1 U8560 ( .A1(n14406), .A2(n9575), .ZN(n11754) );
  INV_X1 U8561 ( .A(n14717), .ZN(n14706) );
  NAND2_X1 U8562 ( .A1(n7283), .A2(n8666), .ZN(n10692) );
  OR2_X1 U8563 ( .A1(n10201), .A2(n13858), .ZN(n14709) );
  INV_X1 U8564 ( .A(n10876), .ZN(n14670) );
  INV_X1 U8565 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8240) );
  INV_X1 U8566 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n6822) );
  INV_X1 U8567 ( .A(n7486), .ZN(n6686) );
  XNOR2_X1 U8568 ( .A(n6699), .B(n9673), .ZN(n13440) );
  NAND2_X1 U8569 ( .A1(n7433), .A2(n7431), .ZN(n9671) );
  XNOR2_X1 U8570 ( .A(n9649), .B(n9648), .ZN(n13447) );
  AND2_X1 U8571 ( .A1(n8611), .A2(n7612), .ZN(n8609) );
  INV_X1 U8572 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8232) );
  XNOR2_X1 U8573 ( .A(n8636), .B(n8635), .ZN(n9922) );
  INV_X1 U8574 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8635) );
  OAI21_X1 U8575 ( .B1(n8634), .B2(P1_IR_REG_22__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U8576 ( .A1(n7570), .A2(n10421), .ZN(n7571) );
  NAND2_X1 U8577 ( .A1(n7571), .A2(n7573), .ZN(n8046) );
  NAND2_X1 U8578 ( .A1(n6700), .A2(SI_18_), .ZN(n7573) );
  INV_X1 U8579 ( .A(n7570), .ZN(n6700) );
  OAI21_X1 U8580 ( .B1(n7899), .B2(n7900), .A(n7553), .ZN(n7919) );
  NAND2_X1 U8581 ( .A1(n7451), .A2(n7549), .ZN(n7879) );
  NAND2_X1 U8582 ( .A1(n7418), .A2(n7535), .ZN(n7804) );
  NAND2_X1 U8583 ( .A1(n7783), .A2(n7533), .ZN(n7418) );
  XNOR2_X1 U8584 ( .A(n14228), .B(n14229), .ZN(n14245) );
  NOR2_X1 U8585 ( .A1(n14252), .A2(n14253), .ZN(n14256) );
  AOI21_X1 U8586 ( .B1(n14952), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n14197), .ZN(
        n14267) );
  AND2_X1 U8587 ( .A1(n14226), .A2(n14227), .ZN(n14197) );
  AOI21_X1 U8588 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14507), .A(n14204), .ZN(
        n14224) );
  AND3_X1 U8589 ( .A1(n8908), .A2(n8907), .A3(n8906), .ZN(n11151) );
  INV_X1 U8590 ( .A(n6798), .ZN(n6792) );
  NAND2_X1 U8591 ( .A1(n6794), .A2(n6797), .ZN(n6793) );
  OR2_X1 U8592 ( .A1(n9836), .A2(n9835), .ZN(n6797) );
  NOR2_X1 U8593 ( .A1(n12024), .A2(n12025), .ZN(n12168) );
  AND2_X1 U8594 ( .A1(n7356), .A2(n7355), .ZN(n11664) );
  NAND2_X1 U8595 ( .A1(n10363), .A2(n7363), .ZN(n10650) );
  AND3_X1 U8596 ( .A1(n8845), .A2(n8844), .A3(n8843), .ZN(n10655) );
  OR2_X1 U8597 ( .A1(n10391), .A2(n10647), .ZN(n8843) );
  NAND2_X1 U8598 ( .A1(n9807), .A2(n6809), .ZN(n12044) );
  AND2_X1 U8599 ( .A1(n11960), .A2(n7338), .ZN(n7337) );
  AND2_X1 U8600 ( .A1(n11955), .A2(n14914), .ZN(n7338) );
  NAND2_X1 U8601 ( .A1(n11146), .A2(n9783), .ZN(n11310) );
  NOR2_X1 U8602 ( .A1(n9773), .A2(n7331), .ZN(n10318) );
  AND2_X1 U8603 ( .A1(n7333), .A2(n7332), .ZN(n7331) );
  NAND2_X1 U8604 ( .A1(n7344), .A2(n7343), .ZN(n12051) );
  NAND2_X1 U8605 ( .A1(n12111), .A2(n12110), .ZN(n7344) );
  NAND2_X1 U8606 ( .A1(n7347), .A2(n7349), .ZN(n12085) );
  NAND2_X1 U8607 ( .A1(n10741), .A2(n6790), .ZN(n10914) );
  NAND2_X1 U8608 ( .A1(n10742), .A2(n10743), .ZN(n10741) );
  NAND2_X1 U8609 ( .A1(n11308), .A2(n9786), .ZN(n11484) );
  OAI211_X1 U8610 ( .C1(n10391), .C2(n15207), .A(n7411), .B(n8820), .ZN(n14917) );
  NAND2_X1 U8611 ( .A1(n10391), .A2(n7412), .ZN(n7411) );
  INV_X1 U8612 ( .A(n9882), .ZN(n7412) );
  NAND2_X1 U8613 ( .A1(n6805), .A2(n6806), .ZN(n12111) );
  OR2_X1 U8614 ( .A1(n9807), .A2(n6808), .ZN(n6805) );
  NAND2_X1 U8615 ( .A1(n11662), .A2(n6817), .ZN(n6816) );
  AND3_X1 U8616 ( .A1(n9106), .A2(n9105), .A3(n9104), .ZN(n12428) );
  XNOR2_X1 U8617 ( .A(n9775), .B(n15036), .ZN(n10365) );
  NAND2_X1 U8618 ( .A1(n10364), .A2(n10365), .ZN(n10363) );
  OR2_X1 U8619 ( .A1(n9804), .A2(n12088), .ZN(n9805) );
  NAND2_X1 U8620 ( .A1(n6783), .A2(n6785), .ZN(n6781) );
  NAND2_X1 U8621 ( .A1(n6780), .A2(n6783), .ZN(n10948) );
  OR2_X1 U8622 ( .A1(n10742), .A2(n6785), .ZN(n6780) );
  AND2_X1 U8623 ( .A1(n9860), .A2(n9845), .ZN(n14916) );
  AND2_X1 U8624 ( .A1(n10319), .A2(n11320), .ZN(n12161) );
  AND2_X1 U8625 ( .A1(n9844), .A2(n15012), .ZN(n12177) );
  NAND2_X1 U8626 ( .A1(n12024), .A2(n9799), .ZN(n7348) );
  INV_X1 U8627 ( .A(n12161), .ZN(n12174) );
  NOR2_X1 U8628 ( .A1(n10276), .A2(n10387), .ZN(n9855) );
  NAND2_X1 U8629 ( .A1(n9493), .A2(n9492), .ZN(n9494) );
  NAND2_X1 U8630 ( .A1(n7321), .A2(n7334), .ZN(n9339) );
  XNOR2_X1 U8631 ( .A(n7322), .B(n9767), .ZN(n7321) );
  INV_X1 U8632 ( .A(n12353), .ZN(n12179) );
  INV_X1 U8633 ( .A(n12367), .ZN(n12340) );
  NAND2_X1 U8634 ( .A1(n9153), .A2(n9152), .ZN(n12379) );
  INV_X1 U8635 ( .A(n12428), .ZN(n12181) );
  INV_X1 U8636 ( .A(n12440), .ZN(n12466) );
  INV_X1 U8637 ( .A(n14347), .ZN(n12184) );
  INV_X1 U8638 ( .A(n12140), .ZN(n12185) );
  NAND2_X1 U8639 ( .A1(n8824), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8825) );
  OAI21_X1 U8640 ( .B1(n10502), .B2(n10501), .A(n6556), .ZN(n10637) );
  NAND2_X1 U8641 ( .A1(n6990), .A2(n10709), .ZN(n10714) );
  NAND2_X1 U8642 ( .A1(n10712), .A2(n10710), .ZN(n6990) );
  AOI21_X1 U8643 ( .B1(n10621), .B2(n10622), .A(n6861), .ZN(n10668) );
  AND2_X1 U8644 ( .A1(n10507), .A2(n10634), .ZN(n6861) );
  NAND2_X1 U8645 ( .A1(n7079), .A2(n7078), .ZN(n10680) );
  NOR2_X1 U8646 ( .A1(n7077), .A2(n11076), .ZN(n11075) );
  NOR2_X1 U8647 ( .A1(n6995), .A2(n11056), .ZN(n11055) );
  NAND2_X1 U8648 ( .A1(n6996), .A2(n6994), .ZN(n10665) );
  NAND2_X1 U8649 ( .A1(n11070), .A2(n11069), .ZN(n11242) );
  XNOR2_X1 U8650 ( .A(n11603), .B(n11610), .ZN(n11519) );
  NOR2_X1 U8651 ( .A1(n11519), .A2(n11521), .ZN(n11604) );
  AND2_X1 U8652 ( .A1(n6867), .A2(n6866), .ZN(n11523) );
  INV_X1 U8653 ( .A(n6991), .ZN(n11607) );
  INV_X1 U8654 ( .A(n6763), .ZN(n12211) );
  NOR2_X1 U8655 ( .A1(n12247), .A2(n12246), .ZN(n12249) );
  NOR2_X1 U8656 ( .A1(n12283), .A2(n12284), .ZN(n12304) );
  AOI21_X1 U8657 ( .B1(n12272), .B2(n12271), .A(n12303), .ZN(n12290) );
  NOR2_X1 U8658 ( .A1(n8785), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n14333) );
  NOR2_X1 U8659 ( .A1(n9237), .A2(n7509), .ZN(n9238) );
  NAND2_X1 U8660 ( .A1(n7135), .A2(n7133), .ZN(n12343) );
  AND2_X1 U8661 ( .A1(n9120), .A2(n9119), .ZN(n12542) );
  NAND2_X1 U8662 ( .A1(n7447), .A2(n7444), .ZN(n12391) );
  NAND2_X1 U8663 ( .A1(n7442), .A2(n9214), .ZN(n12414) );
  NAND2_X1 U8664 ( .A1(n12463), .A2(n6475), .ZN(n12451) );
  NAND2_X1 U8665 ( .A1(n12488), .A2(n9434), .ZN(n12471) );
  NAND2_X1 U8666 ( .A1(n14341), .A2(n9205), .ZN(n12510) );
  NAND2_X1 U8667 ( .A1(n11511), .A2(n9409), .ZN(n14340) );
  OAI21_X1 U8668 ( .B1(n11455), .B2(n9401), .A(n9402), .ZN(n11411) );
  NAND2_X1 U8669 ( .A1(n7436), .A2(n7437), .ZN(n11457) );
  NOR2_X1 U8670 ( .A1(n10287), .A2(n10286), .ZN(n15000) );
  NAND2_X1 U8671 ( .A1(n15000), .A2(n15023), .ZN(n14958) );
  INV_X1 U8672 ( .A(n9313), .ZN(n12020) );
  INV_X1 U8673 ( .A(n11963), .ZN(n12589) );
  INV_X1 U8674 ( .A(n12072), .ZN(n12598) );
  INV_X1 U8675 ( .A(n12050), .ZN(n12610) );
  INV_X1 U8676 ( .A(n12115), .ZN(n12614) );
  NAND2_X1 U8677 ( .A1(n9078), .A2(n9077), .ZN(n12618) );
  INV_X1 U8678 ( .A(n12166), .ZN(n12629) );
  AND2_X1 U8679 ( .A1(n10388), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12640) );
  XNOR2_X1 U8680 ( .A(n6722), .B(n6721), .ZN(n12647) );
  INV_X1 U8681 ( .A(n9294), .ZN(n6721) );
  CLKBUF_X1 U8682 ( .A(n8772), .Z(n12644) );
  XNOR2_X1 U8683 ( .A(n9303), .B(n7327), .ZN(n11883) );
  INV_X1 U8684 ( .A(n9302), .ZN(n7327) );
  INV_X1 U8685 ( .A(n7320), .ZN(n9142) );
  NAND2_X1 U8686 ( .A1(n9242), .A2(n9241), .ZN(n11764) );
  NAND2_X1 U8687 ( .A1(n9245), .A2(n6500), .ZN(n11702) );
  AOI21_X1 U8688 ( .B1(n8734), .B2(n7306), .A(n6497), .ZN(n9108) );
  NAND2_X1 U8689 ( .A1(n8734), .A2(n7308), .ZN(n9099) );
  INV_X1 U8690 ( .A(n9338), .ZN(n10661) );
  INV_X1 U8691 ( .A(SI_19_), .ZN(n10457) );
  NAND2_X1 U8692 ( .A1(n7310), .A2(n8730), .ZN(n9055) );
  OR2_X1 U8693 ( .A1(n9042), .A2(n6601), .ZN(n7310) );
  INV_X1 U8694 ( .A(SI_17_), .ZN(n10327) );
  INV_X1 U8695 ( .A(SI_16_), .ZN(n10246) );
  INV_X1 U8696 ( .A(SI_14_), .ZN(n10099) );
  NAND2_X1 U8697 ( .A1(n7302), .A2(n8723), .ZN(n8994) );
  NAND2_X1 U8698 ( .A1(n8985), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7302) );
  INV_X1 U8699 ( .A(SI_13_), .ZN(n9969) );
  INV_X1 U8700 ( .A(SI_12_), .ZN(n9959) );
  NAND2_X1 U8701 ( .A1(n7289), .A2(n7290), .ZN(n8948) );
  INV_X1 U8702 ( .A(SI_9_), .ZN(n9892) );
  NAND2_X1 U8703 ( .A1(n7293), .A2(n8715), .ZN(n8936) );
  NAND2_X1 U8704 ( .A1(n7295), .A2(n7294), .ZN(n7293) );
  NAND2_X1 U8705 ( .A1(n7314), .A2(n8709), .ZN(n8886) );
  OAI21_X1 U8706 ( .B1(n8812), .B2(n8811), .A(n7075), .ZN(n7074) );
  NAND2_X1 U8707 ( .A1(n12769), .A2(n7242), .ZN(n12650) );
  INV_X1 U8708 ( .A(n12892), .ZN(n14380) );
  INV_X1 U8709 ( .A(n8156), .ZN(n6925) );
  NAND2_X1 U8710 ( .A1(n11187), .A2(n7898), .ZN(n11273) );
  AOI21_X1 U8711 ( .B1(n12799), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n6519), .ZN(
        n7082) );
  NAND2_X1 U8712 ( .A1(n8072), .A2(n8071), .ZN(n13251) );
  NAND2_X1 U8713 ( .A1(n6947), .A2(n7238), .ZN(n6942) );
  NAND2_X1 U8714 ( .A1(n6941), .A2(n7238), .ZN(n6940) );
  INV_X1 U8715 ( .A(n6944), .ZN(n6941) );
  NAND2_X1 U8716 ( .A1(n6516), .A2(n7241), .ZN(n7240) );
  NAND2_X1 U8717 ( .A1(n13072), .A2(n10484), .ZN(n11942) );
  INV_X1 U8718 ( .A(n12671), .ZN(n8123) );
  NAND2_X1 U8719 ( .A1(n12734), .A2(n8105), .ZN(n12672) );
  INV_X1 U8720 ( .A(n6616), .ZN(n7816) );
  CLKBUF_X1 U8721 ( .A(n12713), .Z(n12725) );
  CLKBUF_X1 U8722 ( .A(n12689), .Z(n12690) );
  NAND2_X1 U8723 ( .A1(n7248), .A2(n10921), .ZN(n11189) );
  NAND2_X1 U8724 ( .A1(n6927), .A2(n6539), .ZN(n11690) );
  OR2_X1 U8725 ( .A1(n8215), .A2(n12982), .ZN(n12751) );
  OAI211_X1 U8726 ( .C1(n7248), .C2(n6933), .A(n6939), .B(n6932), .ZN(n11541)
         );
  NAND2_X1 U8727 ( .A1(n6934), .A2(n6935), .ZN(n6932) );
  INV_X1 U8728 ( .A(n6933), .ZN(n6935) );
  NAND2_X1 U8729 ( .A1(n12725), .A2(n8043), .ZN(n12761) );
  NAND2_X1 U8730 ( .A1(n7836), .A2(n7837), .ZN(n10910) );
  NAND2_X1 U8731 ( .A1(n12700), .A2(n7821), .ZN(n10909) );
  OR2_X2 U8732 ( .A1(n8215), .A2(n8214), .ZN(n12759) );
  CLKBUF_X1 U8733 ( .A(n11834), .Z(n11835) );
  INV_X1 U8734 ( .A(n12759), .ZN(n14376) );
  XNOR2_X1 U8735 ( .A(n13027), .B(n13026), .ZN(n13028) );
  NOR2_X1 U8736 ( .A1(n13021), .A2(n13020), .ZN(n13024) );
  INV_X1 U8737 ( .A(n6742), .ZN(n13038) );
  INV_X1 U8738 ( .A(n12956), .ZN(n13045) );
  INV_X1 U8739 ( .A(n10575), .ZN(n13069) );
  NAND2_X1 U8740 ( .A1(n10112), .A2(n10111), .ZN(n10113) );
  NAND2_X1 U8741 ( .A1(n10113), .A2(n10114), .ZN(n10128) );
  NAND2_X1 U8742 ( .A1(n10210), .A2(n10209), .ZN(n13077) );
  NAND2_X1 U8743 ( .A1(n13077), .A2(n13078), .ZN(n13076) );
  AND2_X1 U8744 ( .A1(n6622), .A2(n6571), .ZN(n11439) );
  NOR2_X1 U8745 ( .A1(n14814), .A2(n12008), .ZN(n12009) );
  XNOR2_X1 U8746 ( .A(n13088), .B(n13095), .ZN(n13090) );
  INV_X1 U8747 ( .A(n7097), .ZN(n13139) );
  INV_X1 U8748 ( .A(n13322), .ZN(n13137) );
  INV_X1 U8749 ( .A(n7162), .ZN(n7152) );
  NAND2_X1 U8750 ( .A1(n7104), .A2(n7102), .ZN(n13188) );
  AND2_X1 U8751 ( .A1(n7104), .A2(n6512), .ZN(n13189) );
  INV_X1 U8752 ( .A(n7103), .ZN(n7102) );
  AND2_X1 U8753 ( .A1(n11923), .A2(n11922), .ZN(n13209) );
  NAND2_X1 U8754 ( .A1(n8093), .A2(n8092), .ZN(n13353) );
  NAND2_X1 U8755 ( .A1(n13265), .A2(n11920), .ZN(n13239) );
  NAND2_X1 U8756 ( .A1(n11917), .A2(n11916), .ZN(n13284) );
  AND2_X1 U8757 ( .A1(n7999), .A2(n7998), .ZN(n12886) );
  NAND2_X1 U8758 ( .A1(n11560), .A2(n11559), .ZN(n11648) );
  NAND2_X1 U8759 ( .A1(n11134), .A2(n10968), .ZN(n11039) );
  NAND2_X1 U8760 ( .A1(n7088), .A2(n10957), .ZN(n11281) );
  NAND2_X1 U8761 ( .A1(n10956), .A2(n12998), .ZN(n7088) );
  NAND2_X1 U8762 ( .A1(n6636), .A2(n10567), .ZN(n10764) );
  INV_X1 U8763 ( .A(n13238), .ZN(n13295) );
  INV_X1 U8764 ( .A(n10355), .ZN(n12815) );
  AND2_X2 U8765 ( .A1(n11048), .A2(n10346), .ZN(n14912) );
  NAND2_X1 U8766 ( .A1(n6726), .A2(n6479), .ZN(n13398) );
  INV_X1 U8767 ( .A(n6774), .ZN(n6726) );
  AOI21_X1 U8768 ( .B1(n13318), .B2(n14880), .A(n13317), .ZN(n6753) );
  INV_X1 U8769 ( .A(n13182), .ZN(n13412) );
  INV_X1 U8770 ( .A(n13212), .ZN(n13420) );
  NAND2_X1 U8771 ( .A1(n7944), .A2(n7943), .ZN(n12883) );
  AND2_X2 U8772 ( .A1(n11048), .A2(n11047), .ZN(n15282) );
  AND2_X1 U8773 ( .A1(n10057), .A2(n9868), .ZN(n14835) );
  INV_X1 U8774 ( .A(n7693), .ZN(n11929) );
  NAND2_X1 U8775 ( .A1(n7685), .A2(n7628), .ZN(n7632) );
  XNOR2_X1 U8776 ( .A(n7640), .B(P2_IR_REG_25__SCAN_IN), .ZN(n13461) );
  INV_X1 U8777 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11845) );
  NAND2_X1 U8778 ( .A1(n7643), .A2(n7645), .ZN(n11846) );
  INV_X1 U8779 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n15219) );
  INV_X1 U8780 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10558) );
  INV_X1 U8781 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10184) );
  INV_X1 U8782 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10037) );
  INV_X1 U8783 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9965) );
  INV_X1 U8784 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9954) );
  INV_X1 U8785 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9941) );
  INV_X1 U8786 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9920) );
  NAND2_X1 U8787 ( .A1(n7394), .A2(n13491), .ZN(n14392) );
  NAND2_X1 U8788 ( .A1(n7394), .A2(n7392), .ZN(n14394) );
  AOI21_X1 U8789 ( .B1(n7375), .B2(n7378), .A(n6527), .ZN(n7373) );
  NOR2_X1 U8790 ( .A1(n7384), .A2(n13632), .ZN(n7382) );
  OAI22_X1 U8791 ( .A1(n7385), .A2(n7384), .B1(n13632), .B2(n7387), .ZN(n7383)
         );
  NAND2_X1 U8792 ( .A1(n13597), .A2(n13632), .ZN(n7386) );
  AND2_X1 U8793 ( .A1(n7380), .A2(n6524), .ZN(n11263) );
  INV_X1 U8794 ( .A(n7371), .ZN(n10163) );
  NAND2_X1 U8795 ( .A1(n8271), .A2(n6682), .ZN(n10167) );
  NAND2_X1 U8796 ( .A1(n7401), .A2(n13550), .ZN(n13641) );
  NAND2_X1 U8797 ( .A1(n11681), .A2(n11680), .ZN(n11724) );
  NAND2_X1 U8798 ( .A1(n7367), .A2(n10891), .ZN(n10893) );
  NAND2_X1 U8799 ( .A1(n7402), .A2(n7409), .ZN(n13676) );
  NAND2_X1 U8800 ( .A1(n13662), .A2(n13673), .ZN(n7402) );
  INV_X1 U8801 ( .A(n13683), .ZN(n13577) );
  NAND2_X1 U8802 ( .A1(n7372), .A2(n7375), .ZN(n11370) );
  OR2_X1 U8803 ( .A1(n11262), .A2(n7378), .ZN(n7372) );
  NAND2_X1 U8804 ( .A1(n11637), .A2(n11636), .ZN(n11640) );
  NAND2_X1 U8805 ( .A1(n10010), .A2(n14612), .ZN(n14398) );
  NAND2_X1 U8806 ( .A1(n10016), .A2(n10015), .ZN(n13751) );
  NAND2_X1 U8807 ( .A1(n7180), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9660) );
  NAND2_X1 U8808 ( .A1(n7180), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8581) );
  NAND2_X1 U8809 ( .A1(n7180), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8423) );
  NAND2_X1 U8810 ( .A1(n8295), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8342) );
  AND2_X1 U8811 ( .A1(n6850), .A2(n6849), .ZN(n6853) );
  NAND2_X1 U8812 ( .A1(n8294), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8276) );
  NAND2_X1 U8813 ( .A1(n8295), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6852) );
  INV_X1 U8814 ( .A(n6969), .ZN(n13799) );
  INV_X1 U8815 ( .A(n6972), .ZN(n10038) );
  NOR2_X1 U8816 ( .A1(n10041), .A2(n10040), .ZN(n10248) );
  AND2_X1 U8817 ( .A1(n6972), .A2(n6971), .ZN(n10041) );
  NAND2_X1 U8818 ( .A1(n10044), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6971) );
  NOR2_X1 U8819 ( .A1(n10250), .A2(n10249), .ZN(n10431) );
  AOI21_X1 U8820 ( .B1(n10252), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10251), .ZN(
        n10255) );
  NAND2_X1 U8821 ( .A1(n10728), .A2(n6770), .ZN(n10729) );
  OR2_X1 U8822 ( .A1(n10734), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6770) );
  NAND2_X1 U8823 ( .A1(n10729), .A2(n10730), .ZN(n10986) );
  NOR2_X1 U8824 ( .A1(n10984), .A2(n10983), .ZN(n11419) );
  AOI21_X1 U8825 ( .B1(n11428), .B2(P1_REG1_REG_10__SCAN_IN), .A(n11427), .ZN(
        n14497) );
  AND2_X1 U8826 ( .A1(n13842), .A2(n13841), .ZN(n14546) );
  AND2_X1 U8827 ( .A1(n14560), .A2(n14559), .ZN(n14562) );
  NAND2_X1 U8828 ( .A1(n6963), .A2(n6964), .ZN(n14573) );
  NOR2_X1 U8829 ( .A1(n6965), .A2(n6967), .ZN(n14571) );
  INV_X1 U8830 ( .A(n13837), .ZN(n6963) );
  XNOR2_X1 U8831 ( .A(n8615), .B(n9703), .ZN(n14059) );
  OR2_X1 U8832 ( .A1(n6960), .A2(n13628), .ZN(n7511) );
  AND2_X1 U8833 ( .A1(n7190), .A2(n7189), .ZN(n13884) );
  NAND2_X1 U8834 ( .A1(n13911), .A2(n7512), .ZN(n13906) );
  INV_X1 U8835 ( .A(n14066), .ZN(n13904) );
  INV_X1 U8836 ( .A(n13915), .ZN(n14070) );
  AND2_X1 U8837 ( .A1(n7191), .A2(n6521), .ZN(n13928) );
  NAND2_X1 U8838 ( .A1(n13944), .A2(n8685), .ZN(n13926) );
  NAND2_X1 U8839 ( .A1(n14095), .A2(n8566), .ZN(n13952) );
  NAND2_X1 U8840 ( .A1(n13956), .A2(n8682), .ZN(n13941) );
  INV_X1 U8841 ( .A(n14108), .ZN(n13992) );
  NAND2_X1 U8842 ( .A1(n14003), .A2(n8680), .ZN(n13986) );
  NAND2_X1 U8843 ( .A1(n13999), .A2(n8531), .ZN(n13984) );
  NAND2_X1 U8844 ( .A1(n8521), .A2(n8520), .ZN(n13997) );
  NAND2_X1 U8845 ( .A1(n8512), .A2(n8511), .ZN(n14027) );
  NAND2_X1 U8846 ( .A1(n8679), .A2(n9595), .ZN(n14018) );
  AND2_X1 U8847 ( .A1(n8498), .A2(n8497), .ZN(n14044) );
  OAI21_X1 U8848 ( .B1(n11822), .B2(n7280), .A(n7278), .ZN(n14035) );
  NAND2_X1 U8849 ( .A1(n8491), .A2(n8490), .ZN(n14423) );
  NAND2_X1 U8850 ( .A1(n11752), .A2(n9582), .ZN(n11768) );
  NAND2_X1 U8851 ( .A1(n8474), .A2(n8473), .ZN(n14430) );
  NAND2_X1 U8852 ( .A1(n14410), .A2(n8454), .ZN(n11751) );
  NAND2_X1 U8853 ( .A1(n8438), .A2(n8437), .ZN(n14412) );
  NAND2_X1 U8854 ( .A1(n11473), .A2(n11472), .ZN(n11471) );
  NAND2_X1 U8855 ( .A1(n11342), .A2(n8675), .ZN(n11473) );
  CLKBUF_X1 U8856 ( .A(n11348), .Z(n11350) );
  CLKBUF_X1 U8857 ( .A(n11210), .Z(n11212) );
  NAND2_X1 U8858 ( .A1(n10933), .A2(n10937), .ZN(n7174) );
  NAND2_X1 U8859 ( .A1(n10934), .A2(n8670), .ZN(n10997) );
  NAND2_X1 U8860 ( .A1(n10696), .A2(n8668), .ZN(n10936) );
  CLKBUF_X1 U8861 ( .A(n10687), .Z(n10688) );
  CLKBUF_X1 U8862 ( .A(n10750), .Z(n10752) );
  CLKBUF_X1 U8863 ( .A(n14587), .Z(n14588) );
  CLKBUF_X1 U8864 ( .A(n10850), .Z(n10852) );
  OR2_X1 U8865 ( .A1(n14648), .A2(n10200), .ZN(n14016) );
  OR2_X1 U8866 ( .A1(n14648), .A2(n10008), .ZN(n14640) );
  NAND2_X1 U8867 ( .A1(n10191), .A2(n10006), .ZN(n14612) );
  NAND2_X1 U8868 ( .A1(n14052), .A2(n14051), .ZN(n14136) );
  OAI21_X1 U8869 ( .B1(n6956), .B2(n14717), .A(n14049), .ZN(n14050) );
  NOR2_X1 U8870 ( .A1(n11847), .A2(n14162), .ZN(n9938) );
  AND2_X1 U8871 ( .A1(n9922), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9937) );
  INV_X1 U8872 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8248) );
  INV_X1 U8873 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14157) );
  INV_X1 U8874 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14164) );
  XNOR2_X1 U8875 ( .A(n8629), .B(P1_IR_REG_26__SCAN_IN), .ZN(n14162) );
  NAND2_X1 U8876 ( .A1(n8628), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8629) );
  XNOR2_X1 U8877 ( .A(n8627), .B(P1_IR_REG_25__SCAN_IN), .ZN(n14168) );
  AND2_X1 U8878 ( .A1(n8143), .A2(n8145), .ZN(n11816) );
  NAND2_X1 U8879 ( .A1(n8634), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8619) );
  INV_X1 U8880 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11556) );
  NAND2_X1 U8881 ( .A1(n8112), .A2(n8111), .ZN(n11557) );
  OAI21_X1 U8882 ( .B1(n8616), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8621) );
  INV_X1 U8883 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10559) );
  INV_X1 U8884 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10441) );
  INV_X1 U8885 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10589) );
  INV_X1 U8886 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10274) );
  INV_X1 U8887 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9955) );
  INV_X1 U8888 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9945) );
  INV_X1 U8889 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9932) );
  AND2_X1 U8890 ( .A1(n8317), .A2(n8331), .ZN(n13823) );
  INV_X1 U8891 ( .A(n7526), .ZN(n7756) );
  MUX2_X1 U8892 ( .A(n8241), .B(n8285), .S(P1_IR_REG_2__SCAN_IN), .Z(n8286) );
  NAND2_X1 U8893 ( .A1(n8269), .A2(n8268), .ZN(n9985) );
  CLKBUF_X1 U8894 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n6720) );
  INV_X1 U8895 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14232) );
  XNOR2_X1 U8896 ( .A(n14245), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15285) );
  XNOR2_X1 U8897 ( .A(n14256), .B(n7003), .ZN(n14295) );
  XNOR2_X1 U8898 ( .A(n14259), .B(n14258), .ZN(n15290) );
  INV_X1 U8899 ( .A(n7001), .ZN(n14299) );
  OAI21_X1 U8900 ( .B1(n14296), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6523), .ZN(
        n7001) );
  INV_X1 U8901 ( .A(n14302), .ZN(n7025) );
  AND2_X1 U8902 ( .A1(n7024), .A2(n7022), .ZN(n14272) );
  NOR2_X1 U8903 ( .A1(n14485), .A2(n14286), .ZN(n14314) );
  NAND2_X1 U8904 ( .A1(n14314), .A2(n14315), .ZN(n14313) );
  XNOR2_X1 U8905 ( .A(n14318), .B(n14319), .ZN(n14317) );
  INV_X1 U8906 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n11994) );
  NOR2_X1 U8907 ( .A1(n14317), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n14321) );
  INV_X1 U8908 ( .A(n6986), .ZN(n11231) );
  INV_X1 U8909 ( .A(n6993), .ZN(n12221) );
  AOI21_X1 U8910 ( .B1(n6741), .B2(n14924), .A(n6740), .ZN(n6739) );
  INV_X1 U8911 ( .A(n9868), .ZN(n9869) );
  NAND2_X1 U8912 ( .A1(n6759), .A2(n7106), .ZN(n6758) );
  OAI21_X1 U8913 ( .B1(n13115), .B2(n13298), .A(n6658), .ZN(P2_U3237) );
  AND2_X1 U8914 ( .A1(n6660), .A2(n6659), .ZN(n6658) );
  AOI21_X1 U8915 ( .B1(n13313), .B2(n13288), .A(n13114), .ZN(n6659) );
  INV_X1 U8916 ( .A(n6905), .ZN(n6904) );
  OAI22_X1 U8917 ( .A1(n6742), .A2(P2_U3088), .B1(n11992), .B2(n13464), .ZN(
        n6905) );
  MUX2_X1 U8918 ( .A(n13860), .B(n13859), .S(n13858), .Z(n13862) );
  OR2_X1 U8919 ( .A1(n14740), .A2(n7265), .ZN(n7264) );
  INV_X1 U8920 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7265) );
  OR2_X1 U8921 ( .A1(n14724), .A2(n7182), .ZN(n7181) );
  INV_X1 U8922 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7182) );
  INV_X1 U8923 ( .A(n7013), .ZN(n14477) );
  INV_X1 U8924 ( .A(n14482), .ZN(n7010) );
  AND2_X1 U8925 ( .A1(n12457), .A2(n9212), .ZN(n6475) );
  INV_X2 U8926 ( .A(n12814), .ZN(n12872) );
  INV_X1 U8927 ( .A(n9617), .ZN(n6672) );
  INV_X1 U8928 ( .A(n10315), .ZN(n11951) );
  INV_X1 U8929 ( .A(n14101), .ZN(n6828) );
  AND2_X1 U8930 ( .A1(n13914), .A2(n6958), .ZN(n6477) );
  AND2_X1 U8931 ( .A1(n14481), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n6478) );
  AND2_X1 U8932 ( .A1(n6776), .A2(n13109), .ZN(n6479) );
  AND2_X1 U8933 ( .A1(n7232), .A2(n12954), .ZN(n6480) );
  XNOR2_X1 U8934 ( .A(n10315), .B(n15024), .ZN(n9775) );
  AND2_X1 U8935 ( .A1(n13211), .A2(n7047), .ZN(n6481) );
  AND2_X1 U8936 ( .A1(n12886), .A2(n7042), .ZN(n6482) );
  AND2_X1 U8937 ( .A1(n7150), .A2(n10969), .ZN(n6483) );
  XNOR2_X1 U8938 ( .A(n13124), .B(n13045), .ZN(n13120) );
  OR2_X1 U8939 ( .A1(n6831), .A2(n14608), .ZN(n6484) );
  INV_X1 U8940 ( .A(n13985), .ZN(n7273) );
  AND2_X1 U8941 ( .A1(n10525), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6485) );
  AND2_X1 U8942 ( .A1(n7054), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n6486) );
  AND2_X1 U8943 ( .A1(n6962), .A2(n6961), .ZN(n6487) );
  AND2_X1 U8944 ( .A1(n9353), .A2(n9352), .ZN(n12401) );
  NAND2_X1 U8945 ( .A1(n7573), .A2(n6545), .ZN(n8044) );
  INV_X1 U8946 ( .A(n13269), .ZN(n13429) );
  NAND2_X1 U8947 ( .A1(n8054), .A2(n8053), .ZN(n13269) );
  AND2_X1 U8948 ( .A1(n7351), .A2(n6810), .ZN(n6488) );
  AND2_X1 U8949 ( .A1(n9511), .A2(n9510), .ZN(n6489) );
  INV_X1 U8950 ( .A(n13327), .ZN(n7044) );
  INV_X1 U8951 ( .A(n14301), .ZN(n7028) );
  NAND2_X1 U8952 ( .A1(n14061), .A2(n13628), .ZN(n8687) );
  INV_X1 U8953 ( .A(n8687), .ZN(n6831) );
  NOR2_X1 U8954 ( .A1(n6478), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U8955 ( .A1(n9619), .A2(n7485), .ZN(n6491) );
  AND2_X1 U8956 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n7296), .ZN(n6492) );
  NAND2_X1 U8957 ( .A1(n9582), .A2(n9695), .ZN(n6493) );
  XOR2_X1 U8958 ( .A(n13754), .B(n9645), .Z(n9703) );
  INV_X1 U8959 ( .A(n9551), .ZN(n7468) );
  AND3_X1 U8960 ( .A1(n8617), .A2(n7501), .A3(n8618), .ZN(n6494) );
  INV_X1 U8961 ( .A(n7238), .ZN(n7237) );
  NOR2_X1 U8962 ( .A1(n12649), .A2(n7239), .ZN(n7238) );
  AND2_X1 U8963 ( .A1(n7517), .A2(n8700), .ZN(n6495) );
  AND2_X1 U8964 ( .A1(n8123), .A2(n8105), .ZN(n6496) );
  AND2_X1 U8965 ( .A1(n11932), .A2(n8251), .ZN(n8353) );
  AND2_X1 U8966 ( .A1(n11556), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6497) );
  MUX2_X1 U8967 ( .A(n10394), .B(P3_U3897), .S(n10393), .Z(n14948) );
  INV_X1 U8968 ( .A(n9799), .ZN(n7350) );
  AND2_X1 U8969 ( .A1(n7306), .A2(n7305), .ZN(n6498) );
  INV_X1 U8970 ( .A(n9141), .ZN(n6764) );
  NAND3_X1 U8971 ( .A1(n8276), .A2(n6853), .A3(n6852), .ZN(n10017) );
  OR2_X1 U8972 ( .A1(n9810), .A2(n12441), .ZN(n6499) );
  INV_X1 U8973 ( .A(n8819), .ZN(n9305) );
  AND2_X2 U8974 ( .A1(n8817), .A2(n9925), .ZN(n8819) );
  NAND2_X1 U8975 ( .A1(n8995), .A2(n6752), .ZN(n6500) );
  OR3_X1 U8976 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        n10395), .ZN(n6501) );
  AND3_X1 U8977 ( .A1(n6820), .A2(n6819), .A3(n8840), .ZN(n8995) );
  NAND2_X2 U8978 ( .A1(n11876), .A2(n12198), .ZN(n8817) );
  XNOR2_X1 U8979 ( .A(n8619), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9504) );
  NAND2_X1 U8980 ( .A1(n7758), .A2(n6917), .ZN(n7620) );
  NAND2_X1 U8981 ( .A1(n7524), .A2(SI_0_), .ZN(n9882) );
  AND2_X1 U8982 ( .A1(n7401), .A2(n7398), .ZN(n6502) );
  INV_X1 U8983 ( .A(n8304), .ZN(n8692) );
  AND2_X1 U8984 ( .A1(n12877), .A2(n12876), .ZN(n6504) );
  AND2_X1 U8985 ( .A1(n12843), .A2(n12842), .ZN(n6505) );
  AND2_X1 U8986 ( .A1(n13210), .A2(n11922), .ZN(n6506) );
  OR2_X1 U8987 ( .A1(n12210), .A2(n12209), .ZN(n6507) );
  OR2_X1 U8988 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n8741), .ZN(n6508) );
  AND2_X1 U8989 ( .A1(n8157), .A2(n8156), .ZN(n6509) );
  AND2_X1 U8990 ( .A1(n9647), .A2(n7475), .ZN(n6510) );
  AND2_X1 U8991 ( .A1(n12924), .A2(n12923), .ZN(n6511) );
  INV_X1 U8992 ( .A(n9697), .ZN(n11753) );
  INV_X1 U8993 ( .A(n10484), .ZN(n7033) );
  INV_X1 U8994 ( .A(n7900), .ZN(n7430) );
  XNOR2_X1 U8995 ( .A(n7523), .B(SI_1_), .ZN(n7740) );
  OR2_X1 U8996 ( .A1(n13212), .A2(n13051), .ZN(n6512) );
  AND2_X1 U8997 ( .A1(n12892), .A2(n13057), .ZN(n6513) );
  OR2_X1 U8998 ( .A1(n9598), .A2(n14034), .ZN(n6514) );
  NOR2_X1 U8999 ( .A1(n13308), .A2(n13314), .ZN(n6515) );
  XOR2_X1 U9000 ( .A(n13111), .B(n8212), .Z(n6516) );
  OR2_X1 U9001 ( .A1(n8546), .A2(n9994), .ZN(n6517) );
  INV_X1 U9002 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13442) );
  NAND2_X1 U9003 ( .A1(n8575), .A2(n8574), .ZN(n14082) );
  AND2_X1 U9004 ( .A1(n12853), .A2(n13064), .ZN(n6518) );
  AND2_X1 U9005 ( .A1(n8070), .A2(n10083), .ZN(n6519) );
  NAND2_X1 U9006 ( .A1(n7582), .A2(n7581), .ZN(n7591) );
  AND2_X1 U9007 ( .A1(n14034), .A2(n7277), .ZN(n6520) );
  NAND2_X1 U9008 ( .A1(n9505), .A2(n7462), .ZN(n9506) );
  INV_X1 U9009 ( .A(n14478), .ZN(n7009) );
  NAND2_X1 U9010 ( .A1(n13950), .A2(n8684), .ZN(n6521) );
  NAND2_X1 U9011 ( .A1(n7339), .A2(n12100), .ZN(n12034) );
  NOR2_X1 U9012 ( .A1(n8237), .A2(n8483), .ZN(n8625) );
  NAND2_X1 U9013 ( .A1(n13914), .A2(n6957), .ZN(n6522) );
  OR2_X1 U9014 ( .A1(n14265), .A2(n14264), .ZN(n6523) );
  NAND2_X1 U9015 ( .A1(n11260), .A2(n11259), .ZN(n6524) );
  AND2_X1 U9016 ( .A1(n9252), .A2(n9247), .ZN(n6525) );
  NAND4_X1 U9017 ( .A1(n7613), .A2(n6917), .A3(n6916), .A4(n6915), .ZN(n7784)
         );
  NOR2_X1 U9018 ( .A1(n7470), .A2(n6510), .ZN(n6526) );
  INV_X1 U9019 ( .A(n7133), .ZN(n7132) );
  NOR2_X1 U9020 ( .A1(n12339), .A2(n7134), .ZN(n7133) );
  NAND2_X1 U9021 ( .A1(n8568), .A2(n8567), .ZN(n14087) );
  AND2_X1 U9022 ( .A1(n11369), .A2(n11368), .ZN(n6527) );
  NOR2_X1 U9023 ( .A1(n12892), .A2(n13057), .ZN(n6528) );
  AND2_X1 U9024 ( .A1(n9418), .A2(n9205), .ZN(n6529) );
  AND2_X1 U9025 ( .A1(n9809), .A2(n12452), .ZN(n6530) );
  AND2_X1 U9026 ( .A1(n7045), .A2(n7044), .ZN(n6531) );
  INV_X1 U9027 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7805) );
  INV_X1 U9028 ( .A(n12953), .ZN(n6923) );
  NAND2_X1 U9029 ( .A1(n10156), .A2(n10157), .ZN(n10265) );
  OR2_X1 U9030 ( .A1(n9493), .A2(n15044), .ZN(n6532) );
  INV_X1 U9031 ( .A(n12949), .ZN(n6908) );
  NAND2_X1 U9032 ( .A1(n6887), .A2(n7558), .ZN(n7975) );
  NAND2_X1 U9033 ( .A1(n8614), .A2(n8613), .ZN(n9645) );
  NAND2_X1 U9034 ( .A1(n13988), .A2(n6953), .ZN(n6954) );
  AND2_X1 U9035 ( .A1(n9140), .A2(n9351), .ZN(n6533) );
  INV_X1 U9036 ( .A(n13194), .ZN(n13416) );
  NAND2_X1 U9037 ( .A1(n6897), .A2(n8132), .ZN(n13194) );
  AND2_X1 U9038 ( .A1(n9210), .A2(n9209), .ZN(n6534) );
  NOR2_X1 U9039 ( .A1(n9710), .A2(n9726), .ZN(n6535) );
  INV_X1 U9040 ( .A(n8714), .ZN(n7294) );
  AND2_X1 U9041 ( .A1(n12282), .A2(n12281), .ZN(n6536) );
  XOR2_X1 U9042 ( .A(P3_IR_REG_27__SCAN_IN), .B(n8841), .Z(n6537) );
  AND2_X1 U9043 ( .A1(n14000), .A2(n8680), .ZN(n6538) );
  AND2_X1 U9044 ( .A1(n11691), .A2(n6926), .ZN(n6539) );
  AND2_X1 U9045 ( .A1(n11638), .A2(n11636), .ZN(n6540) );
  AND2_X1 U9046 ( .A1(n9697), .A2(n8454), .ZN(n6541) );
  AND2_X1 U9047 ( .A1(n6691), .A2(n13025), .ZN(n6542) );
  AND2_X1 U9048 ( .A1(n7119), .A2(n9393), .ZN(n6543) );
  AND2_X1 U9049 ( .A1(n13992), .A2(n13762), .ZN(n6544) );
  NOR2_X1 U9050 ( .A1(n7333), .A2(n7330), .ZN(n9773) );
  AND2_X1 U9051 ( .A1(n7571), .A2(n7572), .ZN(n6545) );
  INV_X1 U9052 ( .A(n12954), .ZN(n7234) );
  AND2_X1 U9053 ( .A1(n9317), .A2(n9319), .ZN(n6546) );
  INV_X1 U9054 ( .A(n6840), .ZN(n13921) );
  NAND2_X1 U9055 ( .A1(n13922), .A2(n13923), .ZN(n6840) );
  AND2_X1 U9056 ( .A1(n12095), .A2(n12088), .ZN(n6547) );
  AND2_X1 U9057 ( .A1(n9819), .A2(n12378), .ZN(n6548) );
  AND2_X1 U9058 ( .A1(n11292), .A2(n11165), .ZN(n13007) );
  AND2_X1 U9059 ( .A1(n8240), .A2(n6822), .ZN(n6549) );
  NAND2_X1 U9060 ( .A1(n7233), .A2(n6923), .ZN(n6550) );
  NOR2_X1 U9061 ( .A1(n11381), .A2(n13772), .ZN(n6551) );
  NOR2_X1 U9062 ( .A1(n12836), .A2(n13067), .ZN(n6552) );
  NOR2_X1 U9063 ( .A1(n12865), .A2(n10970), .ZN(n6553) );
  NOR2_X1 U9064 ( .A1(n12559), .A2(n12466), .ZN(n6554) );
  AND2_X1 U9065 ( .A1(n7490), .A2(n6514), .ZN(n6555) );
  OR2_X1 U9066 ( .A1(n10500), .A2(n10519), .ZN(n6556) );
  INV_X1 U9067 ( .A(n6847), .ZN(n6846) );
  NOR2_X1 U9068 ( .A1(n13660), .A2(n13758), .ZN(n6847) );
  AND2_X1 U9069 ( .A1(n7010), .A2(n7012), .ZN(n6557) );
  INV_X1 U9070 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8762) );
  AND2_X1 U9071 ( .A1(n7466), .A2(n6756), .ZN(n6558) );
  OR2_X1 U9072 ( .A1(n13137), .A2(n12654), .ZN(n6559) );
  OR2_X1 U9073 ( .A1(n13088), .A2(n12804), .ZN(n6560) );
  AND2_X1 U9074 ( .A1(n6901), .A2(n12866), .ZN(n6561) );
  INV_X1 U9075 ( .A(n7040), .ZN(n7039) );
  NAND2_X1 U9076 ( .A1(n6482), .A2(n7041), .ZN(n7040) );
  OR2_X1 U9077 ( .A1(n10711), .A2(n10640), .ZN(n6562) );
  INV_X1 U9078 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7676) );
  AND2_X1 U9079 ( .A1(n7556), .A2(n9959), .ZN(n6563) );
  AND2_X1 U9080 ( .A1(n9967), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6564) );
  AND2_X1 U9081 ( .A1(n7555), .A2(n9952), .ZN(n6565) );
  INV_X1 U9082 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9934) );
  INV_X1 U9083 ( .A(n7399), .ZN(n7398) );
  NAND2_X1 U9084 ( .A1(n7400), .A2(n13550), .ZN(n7399) );
  INV_X1 U9085 ( .A(n7445), .ZN(n7444) );
  NAND2_X1 U9086 ( .A1(n7446), .A2(n9217), .ZN(n7445) );
  NAND2_X1 U9087 ( .A1(n6577), .A2(n7457), .ZN(n7123) );
  INV_X1 U9088 ( .A(n7123), .ZN(n6751) );
  AND2_X1 U9089 ( .A1(n9394), .A2(n11198), .ZN(n6566) );
  AND2_X1 U9090 ( .A1(n10891), .A2(n7366), .ZN(n6568) );
  NAND2_X1 U9091 ( .A1(n8594), .A2(n8593), .ZN(n14061) );
  INV_X1 U9092 ( .A(n14061), .ZN(n6960) );
  INV_X1 U9093 ( .A(n9337), .ZN(n9481) );
  NAND2_X1 U9094 ( .A1(n12020), .A2(n12178), .ZN(n9337) );
  AND2_X1 U9095 ( .A1(n9515), .A2(n9514), .ZN(n6569) );
  INV_X1 U9096 ( .A(n6947), .ZN(n6946) );
  AND2_X1 U9097 ( .A1(n12681), .A2(n6948), .ZN(n6947) );
  AND2_X1 U9098 ( .A1(n12167), .A2(n7352), .ZN(n7351) );
  NAND2_X1 U9099 ( .A1(n9778), .A2(n14988), .ZN(n6790) );
  INV_X1 U9100 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9963) );
  INV_X1 U9101 ( .A(n12835), .ZN(n7226) );
  INV_X1 U9102 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14180) );
  NAND2_X1 U9103 ( .A1(n8757), .A2(n7460), .ZN(n7459) );
  INV_X1 U9104 ( .A(n7459), .ZN(n6752) );
  NAND2_X1 U9105 ( .A1(n9255), .A2(n9173), .ZN(n10881) );
  INV_X1 U9106 ( .A(n9695), .ZN(n7275) );
  OR2_X1 U9107 ( .A1(n9607), .A2(n9606), .ZN(n6570) );
  OR2_X1 U9108 ( .A1(n11437), .A2(n11436), .ZN(n6571) );
  NAND2_X1 U9109 ( .A1(n9658), .A2(n9657), .ZN(n13870) );
  INV_X1 U9110 ( .A(n13870), .ZN(n6956) );
  AND3_X1 U9111 ( .A1(n7775), .A2(n7774), .A3(n7083), .ZN(n6572) );
  OAI22_X1 U9112 ( .A1(n7252), .A2(n7740), .B1(n9914), .B2(n7251), .ZN(n7526)
         );
  AND2_X1 U9113 ( .A1(n7156), .A2(n13120), .ZN(n6573) );
  AND2_X1 U9114 ( .A1(n6794), .A2(n6792), .ZN(n6574) );
  AND2_X1 U9115 ( .A1(n7469), .A2(n6535), .ZN(n6575) );
  AND2_X1 U9116 ( .A1(n13823), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6576) );
  AND2_X1 U9117 ( .A1(n8751), .A2(n7125), .ZN(n6577) );
  AND2_X1 U9118 ( .A1(n12395), .A2(n9351), .ZN(n6578) );
  AND2_X1 U9119 ( .A1(n9478), .A2(n9477), .ZN(n6579) );
  AND2_X1 U9120 ( .A1(n9520), .A2(n9519), .ZN(n6580) );
  AND2_X1 U9121 ( .A1(n9096), .A2(n9449), .ZN(n6581) );
  AND2_X1 U9122 ( .A1(n13199), .A2(n11896), .ZN(n6582) );
  AND2_X1 U9123 ( .A1(n9225), .A2(n9224), .ZN(n6583) );
  NOR2_X1 U9124 ( .A1(n8716), .A2(n7292), .ZN(n7291) );
  AND2_X1 U9125 ( .A1(n13124), .A2(n13045), .ZN(n6584) );
  AND2_X1 U9126 ( .A1(n6506), .A2(n11924), .ZN(n6585) );
  AND2_X1 U9127 ( .A1(n12339), .A2(n9224), .ZN(n6586) );
  OR2_X1 U9128 ( .A1(n12941), .A2(n12939), .ZN(n6587) );
  AND2_X1 U9129 ( .A1(n13022), .A2(n6515), .ZN(n6588) );
  INV_X1 U9130 ( .A(n9643), .ZN(n7476) );
  AND2_X1 U9131 ( .A1(n7096), .A2(n13277), .ZN(n6589) );
  OR2_X1 U9132 ( .A1(n7240), .A2(n7236), .ZN(n6590) );
  NAND2_X1 U9133 ( .A1(n7230), .A2(n12930), .ZN(n6591) );
  AND2_X1 U9134 ( .A1(n8617), .A2(n7501), .ZN(n6592) );
  INV_X1 U9135 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8509) );
  OR2_X1 U9136 ( .A1(n9539), .A2(n7500), .ZN(n6593) );
  NAND2_X1 U9137 ( .A1(n9630), .A2(n7483), .ZN(n6594) );
  INV_X1 U9138 ( .A(n13766), .ZN(n7279) );
  INV_X1 U9139 ( .A(n8290), .ZN(n8312) );
  OR2_X1 U9140 ( .A1(n9589), .A2(n9590), .ZN(n6595) );
  INV_X1 U9141 ( .A(n13699), .ZN(n7396) );
  NAND2_X1 U9142 ( .A1(n11835), .A2(n8009), .ZN(n12688) );
  AND2_X1 U9143 ( .A1(n9026), .A2(n9025), .ZN(n9030) );
  NAND2_X1 U9144 ( .A1(n11690), .A2(n7246), .ZN(n14372) );
  NAND2_X1 U9145 ( .A1(n11690), .A2(n7974), .ZN(n14373) );
  NAND2_X1 U9146 ( .A1(n6641), .A2(n11918), .ZN(n13264) );
  INV_X1 U9147 ( .A(n13264), .ZN(n7095) );
  NOR2_X1 U9148 ( .A1(n7354), .A2(n11485), .ZN(n6596) );
  AND4_X1 U9149 ( .A1(n8993), .A2(n8992), .A3(n8991), .A4(n8990), .ZN(n12029)
         );
  INV_X1 U9150 ( .A(n12029), .ZN(n14344) );
  NAND2_X1 U9151 ( .A1(n11654), .A2(n7039), .ZN(n7043) );
  INV_X1 U9152 ( .A(n6871), .ZN(n6870) );
  NAND2_X1 U9153 ( .A1(n6872), .A2(n11069), .ZN(n6871) );
  INV_X1 U9154 ( .A(n12416), .ZN(n12180) );
  AND3_X1 U9155 ( .A1(n9116), .A2(n9115), .A3(n9114), .ZN(n12416) );
  OR2_X1 U9156 ( .A1(n11611), .A2(n11612), .ZN(n7081) );
  OR2_X1 U9157 ( .A1(n11108), .A2(n11109), .ZN(n6622) );
  INV_X1 U9158 ( .A(n8045), .ZN(n7572) );
  AND2_X1 U9159 ( .A1(n7025), .A2(n7028), .ZN(n6597) );
  AND2_X1 U9160 ( .A1(n9800), .A2(n9801), .ZN(n6598) );
  AND2_X1 U9161 ( .A1(n12119), .A2(n14344), .ZN(n6599) );
  AND2_X1 U9162 ( .A1(n7575), .A2(n10457), .ZN(n6600) );
  NOR2_X1 U9163 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n15219), .ZN(n6601) );
  INV_X1 U9164 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7301) );
  AND2_X1 U9165 ( .A1(n6878), .A2(n6877), .ZN(n6602) );
  OR2_X1 U9166 ( .A1(n13251), .A2(n12756), .ZN(n6603) );
  NAND2_X1 U9167 ( .A1(n11237), .A2(n11529), .ZN(n6604) );
  AND2_X1 U9168 ( .A1(n12463), .A2(n9212), .ZN(n6605) );
  INV_X1 U9169 ( .A(n11391), .ZN(n11393) );
  AND2_X1 U9170 ( .A1(n7365), .A2(n7364), .ZN(n6606) );
  AND2_X1 U9171 ( .A1(n7344), .A2(n6499), .ZN(n6607) );
  NAND2_X1 U9172 ( .A1(n13755), .A2(n14387), .ZN(n6608) );
  OR2_X1 U9173 ( .A1(n11272), .A2(n6936), .ZN(n6933) );
  NAND2_X1 U9174 ( .A1(n10331), .A2(n13226), .ZN(n13248) );
  INV_X2 U9175 ( .A(n15080), .ZN(n15081) );
  NAND2_X1 U9176 ( .A1(n11308), .A2(n6596), .ZN(n7356) );
  INV_X1 U9177 ( .A(SI_18_), .ZN(n10421) );
  NAND2_X1 U9178 ( .A1(n7598), .A2(n7599), .ZN(n6609) );
  INV_X1 U9179 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11453) );
  NAND2_X1 U9180 ( .A1(n8373), .A2(n8372), .ZN(n10933) );
  OR2_X1 U9181 ( .A1(n15096), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n6610) );
  XOR2_X1 U9182 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .Z(n6611) );
  NAND2_X1 U9183 ( .A1(n7174), .A2(n8384), .ZN(n10995) );
  NAND2_X1 U9184 ( .A1(n6816), .A2(n7519), .ZN(n12118) );
  NAND2_X1 U9185 ( .A1(n9250), .A2(n9249), .ZN(n9770) );
  INV_X1 U9186 ( .A(n9770), .ZN(n7335) );
  AND2_X1 U9187 ( .A1(n6777), .A2(n9252), .ZN(n6612) );
  NAND2_X1 U9188 ( .A1(n7248), .A2(n7247), .ZN(n11187) );
  XNOR2_X1 U9189 ( .A(n9246), .B(P3_IR_REG_26__SCAN_IN), .ZN(n9252) );
  NOR2_X1 U9190 ( .A1(n12324), .A2(n6882), .ZN(n6613) );
  INV_X1 U9191 ( .A(n7037), .ZN(n11139) );
  AND2_X1 U9192 ( .A1(n7348), .A2(n7351), .ZN(n6614) );
  AND2_X1 U9193 ( .A1(n6867), .A2(n6868), .ZN(n6615) );
  OR2_X1 U9194 ( .A1(n11234), .A2(n11235), .ZN(n7072) );
  INV_X1 U9195 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n15251) );
  INV_X1 U9196 ( .A(n7067), .ZN(n7066) );
  NAND2_X1 U9197 ( .A1(n12271), .A2(n12303), .ZN(n7067) );
  INV_X1 U9198 ( .A(n12865), .ZN(n7036) );
  NAND2_X1 U9199 ( .A1(n8031), .A2(n8030), .ZN(n13287) );
  INV_X1 U9200 ( .A(n13287), .ZN(n7041) );
  INV_X1 U9201 ( .A(n12303), .ZN(n12296) );
  NAND2_X1 U9202 ( .A1(n8416), .A2(n8415), .ZN(n11678) );
  INV_X1 U9203 ( .A(n11678), .ZN(n6961) );
  NAND2_X1 U9204 ( .A1(n6928), .A2(n7826), .ZN(n12849) );
  INV_X1 U9205 ( .A(n12849), .ZN(n6657) );
  NAND2_X1 U9206 ( .A1(n8690), .A2(n8689), .ZN(n14630) );
  AND2_X1 U9207 ( .A1(n8696), .A2(n14612), .ZN(n14648) );
  INV_X1 U9208 ( .A(n14648), .ZN(n14008) );
  AND2_X2 U9209 ( .A1(n11588), .A2(n11587), .ZN(n14740) );
  INV_X1 U9210 ( .A(n9107), .ZN(n7305) );
  INV_X1 U9211 ( .A(n11241), .ZN(n6869) );
  INV_X1 U9212 ( .A(n13091), .ZN(n12804) );
  NAND2_X1 U9213 ( .A1(n8015), .A2(n8014), .ZN(n13372) );
  INV_X1 U9214 ( .A(n13372), .ZN(n7042) );
  XOR2_X1 U9215 ( .A(n7818), .B(n7819), .Z(n6616) );
  INV_X1 U9216 ( .A(n11236), .ZN(n7071) );
  AND2_X1 U9217 ( .A1(n12006), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6617) );
  NAND2_X1 U9218 ( .A1(n12254), .A2(n12280), .ZN(n6618) );
  AND2_X1 U9219 ( .A1(n10363), .A2(n7361), .ZN(n6619) );
  AND2_X1 U9220 ( .A1(n10664), .A2(n10678), .ZN(n11056) );
  AND2_X1 U9221 ( .A1(n7069), .A2(n12296), .ZN(n6620) );
  INV_X1 U9222 ( .A(n9322), .ZN(n15038) );
  INV_X1 U9223 ( .A(n7461), .ZN(n9663) );
  OAI21_X1 U9224 ( .B1(n9506), .B2(n10011), .A(n10019), .ZN(n7461) );
  AND2_X1 U9225 ( .A1(n14169), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6621) );
  INV_X1 U9226 ( .A(n6983), .ZN(n6982) );
  NAND2_X1 U9227 ( .A1(n12281), .A2(n12303), .ZN(n6983) );
  INV_X1 U9228 ( .A(n10305), .ZN(n6624) );
  INV_X1 U9229 ( .A(n9769), .ZN(n7334) );
  INV_X1 U9230 ( .A(n6989), .ZN(n10712) );
  NOR2_X1 U9231 ( .A1(n10639), .A2(n10640), .ZN(n6989) );
  INV_X1 U9232 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7014) );
  INV_X1 U9233 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7031) );
  INV_X1 U9234 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6773) );
  INV_X1 U9235 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7296) );
  INV_X1 U9236 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6915) );
  INV_X1 U9237 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7003) );
  OAI222_X1 U9238 ( .A1(n14163), .A2(n9932), .B1(n14166), .B2(n9931), .C1(
        n10003), .C2(P1_U3086), .ZN(P1_U3350) );
  OAI222_X1 U9239 ( .A1(n14163), .A2(n9934), .B1(n14166), .B2(n9933), .C1(
        n9994), .C2(P1_U3086), .ZN(P1_U3352) );
  OAI222_X1 U9240 ( .A1(n14163), .A2(n9967), .B1(n14171), .B2(n9966), .C1(
        P1_U3086), .C2(n10991), .ZN(P1_U3345) );
  OAI222_X1 U9241 ( .A1(n14163), .A2(n10186), .B1(n14171), .B2(n10185), .C1(
        P1_U3086), .C2(n11426), .ZN(P1_U3343) );
  NAND2_X2 U9242 ( .A1(n7524), .A2(P1_U3086), .ZN(n14163) );
  XNOR2_X1 U9243 ( .A(n12192), .B(n12210), .ZN(n11781) );
  XNOR2_X1 U9244 ( .A(n11437), .B(n11436), .ZN(n11108) );
  NAND2_X1 U9245 ( .A1(n11197), .A2(n11198), .ZN(n6623) );
  NAND2_X1 U9246 ( .A1(n14766), .A2(n10087), .ZN(n10090) );
  NAND2_X1 U9247 ( .A1(n13076), .A2(n10212), .ZN(n14781) );
  NAND2_X1 U9248 ( .A1(n14741), .A2(n10079), .ZN(n14755) );
  NOR2_X2 U9249 ( .A1(n8759), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n8768) );
  NAND4_X2 U9250 ( .A1(n8840), .A2(n8750), .A3(n8749), .A4(n8748), .ZN(n8971)
         );
  NAND2_X1 U9251 ( .A1(n12405), .A2(n9352), .ZN(n6629) );
  NAND2_X1 U9252 ( .A1(n12418), .A2(n9354), .ZN(n6630) );
  NAND2_X1 U9253 ( .A1(n7107), .A2(n9366), .ZN(n8830) );
  AND2_X2 U9254 ( .A1(n9373), .A2(n9368), .ZN(n9366) );
  INV_X1 U9255 ( .A(n10765), .ZN(n12996) );
  NOR2_X2 U9256 ( .A1(n7938), .A2(n7618), .ZN(n6647) );
  NAND3_X1 U9257 ( .A1(n7204), .A2(n7202), .A3(n6645), .ZN(n7633) );
  AND2_X1 U9258 ( .A1(n6647), .A2(n7626), .ZN(n6645) );
  NAND2_X1 U9259 ( .A1(n7786), .A2(n6647), .ZN(n7678) );
  AOI21_X2 U9260 ( .B1(n11653), .B2(n11652), .A(n11651), .ZN(n11713) );
  NAND2_X1 U9261 ( .A1(n6727), .A2(n7901), .ZN(n6650) );
  NAND2_X2 U9262 ( .A1(n13449), .A2(n7693), .ZN(n12790) );
  XNOR2_X1 U9263 ( .A(n13113), .B(n13112), .ZN(n13315) );
  OAI22_X1 U9264 ( .A1(n11298), .A2(n11297), .B1(n13060), .B2(n12875), .ZN(
        n11401) );
  NAND3_X1 U9265 ( .A1(n6665), .A2(n7469), .A3(n6664), .ZN(n9733) );
  NAND3_X1 U9266 ( .A1(n6665), .A2(n6575), .A3(n6664), .ZN(n9735) );
  NOR2_X4 U9267 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n8267) );
  NAND3_X1 U9268 ( .A1(n9523), .A2(n9518), .A3(n6668), .ZN(n6670) );
  NAND3_X1 U9269 ( .A1(n6670), .A2(n9526), .A3(n6669), .ZN(n9529) );
  NAND2_X1 U9270 ( .A1(n9523), .A2(n6580), .ZN(n6669) );
  OAI22_X1 U9271 ( .A1(n9561), .A2(n6674), .B1(n6675), .B2(n9562), .ZN(n9565)
         );
  NAND3_X1 U9272 ( .A1(n6680), .A2(n6593), .A3(n6679), .ZN(n6678) );
  OR2_X1 U9273 ( .A1(n9537), .A2(n9538), .ZN(n6679) );
  NAND2_X1 U9274 ( .A1(n6681), .A2(n9536), .ZN(n6680) );
  NAND2_X1 U9275 ( .A1(n9537), .A2(n9538), .ZN(n6681) );
  INV_X2 U9276 ( .A(n10167), .ZN(n14652) );
  NOR2_X1 U9277 ( .A1(n8270), .A2(n6683), .ZN(n6682) );
  NOR2_X2 U9278 ( .A1(n8628), .A2(n7486), .ZN(n8242) );
  INV_X1 U9279 ( .A(n6684), .ZN(n6823) );
  NOR2_X1 U9280 ( .A1(n8628), .A2(n6685), .ZN(n6684) );
  XNOR2_X2 U9281 ( .A(n6687), .B(n8248), .ZN(n11932) );
  NAND2_X1 U9282 ( .A1(n10160), .A2(n10265), .ZN(n10162) );
  NAND2_X1 U9283 ( .A1(n10887), .A2(n10886), .ZN(n7367) );
  NAND2_X2 U9284 ( .A1(n13729), .A2(n13730), .ZN(n13728) );
  NAND2_X1 U9285 ( .A1(n13604), .A2(n13605), .ZN(n13570) );
  NAND2_X1 U9286 ( .A1(n6690), .A2(n13700), .ZN(n13604) );
  OAI21_X2 U9287 ( .B1(n13662), .B2(n7406), .A(n7403), .ZN(n13708) );
  XNOR2_X2 U9288 ( .A(n13508), .B(n13507), .ZN(n13744) );
  OAI21_X2 U9289 ( .B1(n6886), .B2(n6694), .A(n6692), .ZN(n8025) );
  OAI21_X1 U9290 ( .B1(n9649), .B2(n6698), .A(n6695), .ZN(n6699) );
  NAND2_X1 U9291 ( .A1(n6702), .A2(n7546), .ZN(n7857) );
  NAND2_X1 U9292 ( .A1(n7839), .A2(n7544), .ZN(n6702) );
  NAND2_X1 U9293 ( .A1(n7838), .A2(n7546), .ZN(n6703) );
  INV_X1 U9294 ( .A(n7546), .ZN(n6704) );
  NAND2_X1 U9295 ( .A1(n7543), .A2(n7542), .ZN(n7839) );
  NAND2_X1 U9296 ( .A1(n6707), .A2(n7416), .ZN(n7415) );
  NAND2_X1 U9297 ( .A1(n6707), .A2(n7532), .ZN(n7783) );
  NAND2_X1 U9298 ( .A1(n7770), .A2(n7530), .ZN(n6707) );
  NAND2_X1 U9299 ( .A1(n6708), .A2(n7591), .ZN(n7592) );
  NAND3_X1 U9300 ( .A1(n7591), .A2(n7590), .A3(n8130), .ZN(n6708) );
  OAI21_X1 U9301 ( .B1(n8129), .B2(n8130), .A(n6708), .ZN(n11993) );
  INV_X1 U9302 ( .A(n10715), .ZN(n7055) );
  NOR2_X1 U9303 ( .A1(n11532), .A2(n11520), .ZN(n11611) );
  INV_X1 U9304 ( .A(n11076), .ZN(n7078) );
  NOR2_X1 U9305 ( .A1(n11078), .A2(n11465), .ZN(n11234) );
  INV_X1 U9306 ( .A(n7070), .ZN(n12264) );
  NAND2_X1 U9307 ( .A1(n12330), .A2(n6739), .ZN(P3_U3201) );
  XOR2_X1 U9308 ( .A(n6762), .B(n6761), .Z(n6741) );
  NAND2_X1 U9309 ( .A1(n7529), .A2(n7528), .ZN(n7770) );
  NAND2_X1 U9310 ( .A1(n6713), .A2(n6712), .ZN(n12802) );
  NAND2_X1 U9311 ( .A1(n6560), .A2(n6461), .ZN(n6712) );
  OR2_X1 U9312 ( .A1(n12801), .A2(n6461), .ZN(n6713) );
  OR2_X1 U9313 ( .A1(n8781), .A2(n8779), .ZN(n7318) );
  OAI21_X1 U9314 ( .B1(n9396), .B2(n9395), .A(n6566), .ZN(n9400) );
  NAND2_X1 U9315 ( .A1(n6719), .A2(n12355), .ZN(n9468) );
  NAND2_X1 U9316 ( .A1(n9466), .A2(n9467), .ZN(n6719) );
  NAND2_X2 U9317 ( .A1(n11884), .A2(n11879), .ZN(n8822) );
  NAND2_X1 U9318 ( .A1(n8729), .A2(n8728), .ZN(n9042) );
  OR3_X1 U9319 ( .A1(n9420), .A2(n9419), .A3(n9418), .ZN(n9425) );
  NOR2_X1 U9320 ( .A1(n9284), .A2(n9283), .ZN(n9285) );
  NOR2_X1 U9321 ( .A1(n9156), .A2(n9154), .ZN(n8742) );
  NOR2_X1 U9322 ( .A1(n13632), .A2(n13597), .ZN(n7385) );
  NAND2_X1 U9323 ( .A1(n7503), .A2(n14543), .ZN(n14542) );
  NAND2_X1 U9324 ( .A1(n7266), .A2(n14740), .ZN(n7263) );
  NAND2_X1 U9325 ( .A1(n7186), .A2(n14714), .ZN(n7185) );
  NOR2_X1 U9326 ( .A1(n14528), .A2(n6975), .ZN(n13827) );
  NOR2_X1 U9327 ( .A1(n14499), .A2(n6973), .ZN(n11421) );
  NOR2_X1 U9328 ( .A1(n13813), .A2(n6576), .ZN(n9997) );
  AOI21_X1 U9329 ( .B1(n7320), .B2(n6764), .A(n6621), .ZN(n9156) );
  AOI21_X1 U9330 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n14157), .A(n9285), .ZN(
        n9291) );
  NAND2_X1 U9331 ( .A1(n6883), .A2(n7551), .ZN(n7899) );
  NAND2_X1 U9332 ( .A1(n10577), .A2(n10576), .ZN(n10613) );
  AOI21_X1 U9333 ( .B1(n13116), .B2(n13101), .A(n13112), .ZN(n13103) );
  INV_X1 U9334 ( .A(n13312), .ZN(n6776) );
  XNOR2_X1 U9335 ( .A(n11903), .B(n13020), .ZN(n11912) );
  OAI21_X1 U9336 ( .B1(n9529), .B2(n9528), .A(n9527), .ZN(n9531) );
  OAI22_X1 U9337 ( .A1(n9535), .A2(n7480), .B1(n9534), .B2(n9533), .ZN(n9537)
         );
  NAND2_X1 U9338 ( .A1(n9549), .A2(n9548), .ZN(n9552) );
  AOI21_X1 U9339 ( .B1(n9522), .B2(n9521), .A(n10372), .ZN(n9523) );
  XNOR2_X1 U9340 ( .A(n13827), .B(n8458), .ZN(n11860) );
  NOR2_X1 U9341 ( .A1(n9980), .A2(n13782), .ZN(n9992) );
  NOR2_X1 U9342 ( .A1(n14526), .A2(n14527), .ZN(n14528) );
  NOR2_X1 U9343 ( .A1(n14500), .A2(n14501), .ZN(n14499) );
  NAND2_X1 U9344 ( .A1(n13447), .A2(n12782), .ZN(n11902) );
  NAND2_X1 U9345 ( .A1(n7589), .A2(n6765), .ZN(n7590) );
  AND2_X2 U9346 ( .A1(n10053), .A2(n9926), .ZN(n7901) );
  AOI21_X1 U9347 ( .B1(n13121), .B2(n7155), .A(n6584), .ZN(n13113) );
  XNOR2_X1 U9348 ( .A(n11926), .B(n13020), .ZN(n13311) );
  XNOR2_X1 U9349 ( .A(n8157), .B(n6925), .ZN(n11972) );
  NAND2_X1 U9350 ( .A1(n8101), .A2(n12738), .ZN(n12734) );
  NAND2_X2 U9351 ( .A1(n10801), .A2(n7855), .ZN(n10923) );
  NAND2_X1 U9352 ( .A1(n14372), .A2(n7989), .ZN(n8008) );
  NAND2_X1 U9353 ( .A1(n7901), .A2(n9897), .ZN(n7743) );
  NAND2_X1 U9354 ( .A1(n12673), .A2(n8128), .ZN(n8141) );
  NAND2_X1 U9355 ( .A1(n6943), .A2(n6947), .ZN(n12682) );
  NAND2_X1 U9356 ( .A1(n12700), .A2(n7244), .ZN(n10795) );
  NAND2_X1 U9357 ( .A1(n8039), .A2(n12718), .ZN(n12713) );
  NAND2_X1 U9358 ( .A1(n10489), .A2(n7768), .ZN(n9875) );
  NAND2_X1 U9359 ( .A1(n7781), .A2(n7780), .ZN(n9873) );
  NAND2_X1 U9360 ( .A1(n11834), .A2(n6929), .ZN(n12689) );
  NAND2_X2 U9361 ( .A1(n6728), .A2(n6743), .ZN(n10495) );
  INV_X1 U9362 ( .A(n11949), .ZN(n6728) );
  XNOR2_X1 U9363 ( .A(n7752), .B(n7754), .ZN(n11949) );
  INV_X1 U9364 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n6894) );
  INV_X1 U9365 ( .A(P1_RD_REG_SCAN_IN), .ZN(n6896) );
  NAND2_X1 U9366 ( .A1(n8195), .A2(n7609), .ZN(n8610) );
  NAND2_X1 U9367 ( .A1(n7451), .A2(n7450), .ZN(n6883) );
  NAND2_X1 U9368 ( .A1(n7522), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6731) );
  OAI21_X1 U9369 ( .B1(n10017), .B2(n10203), .A(n9509), .ZN(n9685) );
  INV_X1 U9370 ( .A(n11171), .ZN(n6736) );
  NAND2_X1 U9371 ( .A1(n7154), .A2(n7158), .ZN(n13117) );
  NAND2_X1 U9372 ( .A1(n13119), .A2(n13198), .ZN(n6755) );
  NAND3_X1 U9373 ( .A1(n10265), .A2(n10150), .A3(n10149), .ZN(n7368) );
  INV_X4 U9374 ( .A(n13629), .ZN(n13587) );
  NAND2_X1 U9375 ( .A1(n7433), .A2(n9651), .ZN(n9654) );
  INV_X1 U9376 ( .A(n6967), .ZN(n6964) );
  NOR2_X1 U9377 ( .A1(n13789), .A2(n6970), .ZN(n13801) );
  NOR2_X1 U9378 ( .A1(n11419), .A2(n6974), .ZN(n14501) );
  NOR2_X1 U9379 ( .A1(n14515), .A2(n6976), .ZN(n14526) );
  OAI21_X1 U9380 ( .B1(n9591), .B2(n7496), .A(n6595), .ZN(n9594) );
  AOI21_X1 U9381 ( .B1(n9552), .B2(n7466), .A(n7464), .ZN(n7463) );
  OAI21_X1 U9382 ( .B1(n6769), .B2(n6768), .A(n14413), .ZN(n9580) );
  NAND2_X1 U9383 ( .A1(n6738), .A2(n8302), .ZN(n10850) );
  NAND3_X1 U9384 ( .A1(n7176), .A2(n7175), .A3(n10372), .ZN(n6738) );
  OAI21_X2 U9385 ( .B1(n13487), .B2(n7391), .A(n7388), .ZN(n13508) );
  NAND2_X1 U9386 ( .A1(n8508), .A2(n6592), .ZN(n8622) );
  NAND2_X1 U9387 ( .A1(n13882), .A2(n7511), .ZN(n8615) );
  OAI21_X1 U9388 ( .B1(n14058), .B2(n14638), .A(n6495), .ZN(P1_U3356) );
  NAND3_X1 U9389 ( .A1(n7369), .A2(n10268), .A3(n7368), .ZN(n10468) );
  XNOR2_X1 U9390 ( .A(n8610), .B(n8609), .ZN(n14156) );
  INV_X1 U9391 ( .A(n14059), .ZN(n7186) );
  NAND2_X1 U9392 ( .A1(n7183), .A2(n7181), .ZN(P1_U3525) );
  NAND3_X1 U9393 ( .A1(n13883), .A2(n7190), .A3(n7189), .ZN(n13882) );
  NAND2_X1 U9394 ( .A1(n6991), .A2(n11602), .ZN(n11780) );
  INV_X1 U9395 ( .A(n7074), .ZN(n7073) );
  NAND2_X1 U9396 ( .A1(n7817), .A2(n7816), .ZN(n12700) );
  NOR2_X4 U9397 ( .A1(n11978), .A2(n6509), .ZN(n12728) );
  NAND2_X1 U9398 ( .A1(n6938), .A2(n6937), .ZN(n11538) );
  BUF_X4 U9399 ( .A(n8817), .Z(n10391) );
  NAND2_X1 U9400 ( .A1(n9228), .A2(n9227), .ZN(n9744) );
  NAND2_X1 U9401 ( .A1(n10785), .A2(n10784), .ZN(n10783) );
  NAND2_X1 U9402 ( .A1(n12350), .A2(n9221), .ZN(n9225) );
  NAND2_X2 U9403 ( .A1(n14341), .A2(n6529), .ZN(n12508) );
  NAND2_X1 U9404 ( .A1(n12496), .A2(n12495), .ZN(n12494) );
  OAI21_X2 U9405 ( .B1(n12402), .B2(n7445), .A(n7443), .ZN(n12377) );
  NAND2_X1 U9406 ( .A1(n12424), .A2(n12429), .ZN(n7442) );
  NAND3_X1 U9407 ( .A1(n12968), .A2(n12967), .A3(n12969), .ZN(n6744) );
  NAND2_X1 U9408 ( .A1(n7958), .A2(n7959), .ZN(n6887) );
  OAI21_X2 U9409 ( .B1(n6511), .B2(n7227), .A(n7228), .ZN(n12933) );
  NAND3_X1 U9410 ( .A1(n12938), .A2(n12937), .A3(n6587), .ZN(n6745) );
  OR3_X1 U9411 ( .A1(n6914), .A2(n7206), .A3(n7205), .ZN(n12925) );
  NAND2_X1 U9412 ( .A1(n7421), .A2(n7420), .ZN(n7958) );
  NAND2_X1 U9413 ( .A1(n11293), .A2(n11292), .ZN(n11386) );
  NOR2_X2 U9414 ( .A1(n9168), .A2(n8756), .ZN(n8757) );
  NAND2_X1 U9415 ( .A1(n8161), .A2(n7598), .ZN(n8175) );
  OAI21_X2 U9416 ( .B1(n13264), .B2(n7092), .A(n7089), .ZN(n13219) );
  OAI21_X1 U9417 ( .B1(n13315), .B2(n14851), .A(n6775), .ZN(n6774) );
  NAND2_X1 U9418 ( .A1(n10838), .A2(n10837), .ZN(n10565) );
  AOI21_X1 U9419 ( .B1(n6760), .B2(n13248), .A(n6758), .ZN(n7105) );
  INV_X1 U9420 ( .A(n13310), .ZN(n6760) );
  NAND3_X1 U9421 ( .A1(n7317), .A2(n7315), .A3(n8703), .ZN(n8838) );
  NAND2_X1 U9422 ( .A1(n9898), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8701) );
  NAND2_X1 U9423 ( .A1(n6532), .A2(n9494), .ZN(n9497) );
  NAND2_X1 U9424 ( .A1(n8865), .A2(n8864), .ZN(n7314) );
  NAND2_X1 U9425 ( .A1(n8740), .A2(n8739), .ZN(n8741) );
  AND2_X2 U9426 ( .A1(n9745), .A2(n6579), .ZN(n9482) );
  XNOR2_X1 U9427 ( .A(n11232), .B(n11233), .ZN(n11078) );
  NAND2_X1 U9428 ( .A1(n7169), .A2(n6603), .ZN(n13240) );
  NAND2_X1 U9429 ( .A1(n10833), .A2(n12992), .ZN(n10577) );
  NAND2_X1 U9430 ( .A1(n7633), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7634) );
  NAND2_X1 U9431 ( .A1(n7592), .A2(n7593), .ZN(n7595) );
  NAND2_X1 U9432 ( .A1(n13877), .A2(n6829), .ZN(n6830) );
  NAND4_X1 U9433 ( .A1(n6894), .A2(n6893), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6766) );
  NAND2_X2 U9434 ( .A1(n14168), .A2(n6767), .ZN(n10023) );
  NAND2_X1 U9435 ( .A1(n8612), .A2(n8611), .ZN(n9649) );
  NAND2_X1 U9436 ( .A1(n7594), .A2(SI_23_), .ZN(n8143) );
  NAND2_X2 U9437 ( .A1(n11724), .A2(n11723), .ZN(n13487) );
  NAND2_X2 U9438 ( .A1(n13718), .A2(n11019), .ZN(n11262) );
  NAND2_X1 U9439 ( .A1(n6993), .A2(n6992), .ZN(n12222) );
  XNOR2_X1 U9440 ( .A(n11226), .B(n11233), .ZN(n11057) );
  NAND2_X1 U9441 ( .A1(n12803), .A2(n12802), .ZN(n12969) );
  NAND2_X1 U9442 ( .A1(n9613), .A2(n9614), .ZN(n9616) );
  NOR2_X1 U9443 ( .A1(n9572), .A2(n9573), .ZN(n6768) );
  NAND2_X1 U9444 ( .A1(n7482), .A2(n7481), .ZN(n9633) );
  INV_X4 U9445 ( .A(n8279), .ZN(n9659) );
  AND2_X2 U9446 ( .A1(n11972), .A2(n6924), .ZN(n11978) );
  NOR2_X1 U9447 ( .A1(n7160), .A2(n7159), .ZN(n7158) );
  INV_X1 U9448 ( .A(n7741), .ZN(n7252) );
  OAI21_X1 U9449 ( .B1(n13311), .B2(n13238), .A(n7105), .ZN(P2_U3236) );
  INV_X1 U9450 ( .A(n13241), .ZN(n7169) );
  NAND2_X1 U9451 ( .A1(n7514), .A2(n7165), .ZN(n7164) );
  AOI21_X1 U9452 ( .B1(n13200), .B2(n7166), .A(n7164), .ZN(n7163) );
  NAND3_X1 U9453 ( .A1(n9817), .A2(n12416), .A3(n9818), .ZN(n12129) );
  NAND2_X1 U9454 ( .A1(n9817), .A2(n9818), .ZN(n12128) );
  NAND2_X1 U9455 ( .A1(n6783), .A2(n10742), .ZN(n6782) );
  NAND3_X1 U9456 ( .A1(n6782), .A2(n10947), .A3(n6781), .ZN(n10946) );
  NAND2_X1 U9457 ( .A1(n12156), .A2(n6574), .ZN(n6791) );
  OAI211_X1 U9458 ( .C1(n12156), .C2(n6793), .A(n6791), .B(n14914), .ZN(n9867)
         );
  NAND2_X1 U9459 ( .A1(n12156), .A2(n12158), .ZN(n12157) );
  OAI21_X1 U9460 ( .B1(n12156), .B2(n9835), .A(n6798), .ZN(n11966) );
  NAND2_X1 U9461 ( .A1(n9807), .A2(n6803), .ZN(n6802) );
  OR2_X1 U9462 ( .A1(n9808), .A2(n12440), .ZN(n6809) );
  AND2_X1 U9463 ( .A1(n8750), .A2(n8748), .ZN(n6819) );
  NAND2_X1 U9464 ( .A1(n8995), .A2(n8757), .ZN(n9243) );
  NAND2_X2 U9465 ( .A1(n14659), .A2(n10164), .ZN(n9521) );
  NAND2_X1 U9466 ( .A1(n8242), .A2(n8240), .ZN(n8247) );
  NAND2_X1 U9467 ( .A1(n8679), .A2(n6825), .ZN(n6824) );
  NAND3_X1 U9468 ( .A1(n8688), .A2(n14630), .A3(n6831), .ZN(n6833) );
  NAND2_X1 U9469 ( .A1(n7255), .A2(n6837), .ZN(n6835) );
  NAND2_X1 U9470 ( .A1(n6835), .A2(n6836), .ZN(n11766) );
  NAND2_X1 U9471 ( .A1(n13944), .A2(n6844), .ZN(n6843) );
  NAND3_X1 U9472 ( .A1(n11932), .A2(n8251), .A3(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6849) );
  NAND2_X2 U9473 ( .A1(n8255), .A2(n14155), .ZN(n8279) );
  AND2_X2 U9474 ( .A1(n11932), .A2(n14155), .ZN(n8295) );
  NOR2_X1 U9475 ( .A1(n6856), .A2(n8971), .ZN(n6854) );
  NAND2_X1 U9476 ( .A1(n6752), .A2(n6854), .ZN(n6855) );
  NAND2_X4 U9477 ( .A1(n6857), .A2(n6855), .ZN(n12198) );
  AOI22_X2 U9478 ( .A1(n7459), .A2(n6860), .B1(n6858), .B2(n6537), .ZN(n6857)
         );
  INV_X1 U9479 ( .A(n11240), .ZN(n6872) );
  NOR2_X1 U9480 ( .A1(n12277), .A2(n12276), .ZN(n12295) );
  AOI21_X1 U9481 ( .B1(n12251), .B2(n6618), .A(n6875), .ZN(n6873) );
  INV_X1 U9482 ( .A(n12229), .ZN(n6874) );
  INV_X1 U9483 ( .A(n12251), .ZN(n6877) );
  NAND2_X1 U9484 ( .A1(n12229), .A2(n12230), .ZN(n6878) );
  NAND2_X1 U9485 ( .A1(n7958), .A2(n6888), .ZN(n6886) );
  NAND2_X1 U9486 ( .A1(n8086), .A2(n6891), .ZN(n7582) );
  MUX2_X1 U9487 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n9925), .Z(n7541) );
  NAND4_X1 U9488 ( .A1(n7520), .A2(n11994), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n6896), .ZN(n6895) );
  NAND2_X1 U9489 ( .A1(n12844), .A2(n12845), .ZN(n12843) );
  NAND3_X1 U9490 ( .A1(n12861), .A2(n7216), .A3(n12860), .ZN(n6903) );
  OAI21_X1 U9491 ( .B1(n11993), .B2(n13459), .A(n6904), .ZN(P2_U3305) );
  OR2_X1 U9492 ( .A1(n12943), .A2(n6911), .ZN(n6906) );
  NAND2_X1 U9493 ( .A1(n12943), .A2(n6910), .ZN(n6909) );
  OR3_X1 U9494 ( .A1(n6914), .A2(n7206), .A3(n6913), .ZN(n12927) );
  NAND2_X1 U9495 ( .A1(n6919), .A2(n6922), .ZN(n12960) );
  NAND3_X1 U9496 ( .A1(n12951), .A2(n12950), .A3(n6920), .ZN(n6919) );
  MUX2_X1 U9497 ( .A(n13068), .B(n12833), .S(n12872), .Z(n12835) );
  OAI21_X1 U9498 ( .B1(n11579), .B2(n11575), .A(n11576), .ZN(n11692) );
  NAND2_X1 U9499 ( .A1(n11575), .A2(n11576), .ZN(n6926) );
  NAND2_X1 U9500 ( .A1(n11574), .A2(n11576), .ZN(n6927) );
  XNOR2_X1 U9501 ( .A(n7823), .B(n7822), .ZN(n9918) );
  NAND2_X1 U9502 ( .A1(n11833), .A2(n8005), .ZN(n11834) );
  NAND2_X1 U9503 ( .A1(n7248), .A2(n6939), .ZN(n6931) );
  OAI21_X1 U9504 ( .B1(n6931), .B2(n6934), .A(n6930), .ZN(n6938) );
  MUX2_X1 U9505 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n7522), .Z(n7534) );
  NAND2_X1 U9506 ( .A1(n12728), .A2(n8174), .ZN(n6943) );
  NOR2_X1 U9507 ( .A1(n12728), .A2(n12727), .ZN(n12726) );
  OAI21_X1 U9508 ( .B1(n12728), .B2(n6946), .A(n6944), .ZN(n12769) );
  OAI21_X1 U9509 ( .B1(n12728), .B2(n6942), .A(n6940), .ZN(n12651) );
  INV_X1 U9510 ( .A(n6954), .ZN(n13959) );
  NAND2_X1 U9511 ( .A1(n13914), .A2(n13904), .ZN(n13899) );
  NAND3_X1 U9512 ( .A1(n6487), .A2(n11591), .A3(n11001), .ZN(n14415) );
  INV_X1 U9513 ( .A(n13836), .ZN(n6966) );
  NAND2_X1 U9514 ( .A1(n12249), .A2(n6982), .ZN(n6977) );
  OAI21_X1 U9515 ( .B1(n6981), .B2(n6983), .A(n6984), .ZN(n6979) );
  INV_X1 U9516 ( .A(n6988), .ZN(n6987) );
  OAI21_X1 U9517 ( .B1(n10710), .B2(n10711), .A(n10511), .ZN(n6988) );
  INV_X1 U9518 ( .A(n11056), .ZN(n6994) );
  NAND2_X1 U9519 ( .A1(n7002), .A2(n14257), .ZN(n14259) );
  NAND3_X1 U9520 ( .A1(n7005), .A2(n7004), .A3(n7011), .ZN(n14285) );
  INV_X1 U9521 ( .A(n14479), .ZN(n7007) );
  NAND2_X1 U9522 ( .A1(n14473), .A2(n14474), .ZN(n14472) );
  NAND2_X1 U9523 ( .A1(n14473), .A2(n7017), .ZN(n7016) );
  OR2_X1 U9524 ( .A1(n14474), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n7017) );
  XNOR2_X1 U9525 ( .A(n14274), .B(n14273), .ZN(n14476) );
  NAND2_X1 U9526 ( .A1(n7024), .A2(n7026), .ZN(n14469) );
  NAND2_X1 U9527 ( .A1(n7019), .A2(n7018), .ZN(n7024) );
  INV_X1 U9528 ( .A(n14297), .ZN(n7018) );
  NOR2_X1 U9529 ( .A1(n14297), .A2(n7020), .ZN(n14302) );
  INV_X1 U9530 ( .A(n7021), .ZN(n7020) );
  AND2_X1 U9531 ( .A1(n7021), .A2(n7027), .ZN(n7019) );
  NOR2_X1 U9532 ( .A1(n7023), .A2(n14470), .ZN(n7022) );
  MUX2_X1 U9533 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13465), .S(n10053), .Z(n10484)
         );
  NOR2_X2 U9534 ( .A1(n10839), .A2(n12833), .ZN(n10772) );
  NOR2_X2 U9535 ( .A1(n11282), .A2(n14885), .ZN(n7037) );
  AND2_X1 U9536 ( .A1(n13122), .A2(n6515), .ZN(n13096) );
  NAND2_X1 U9537 ( .A1(n13122), .A2(n6588), .ZN(n13095) );
  AND2_X1 U9538 ( .A1(n13122), .A2(n13111), .ZN(n13108) );
  NAND2_X1 U9539 ( .A1(n11654), .A2(n7038), .ZN(n13267) );
  INV_X1 U9540 ( .A(n7043), .ZN(n13285) );
  NAND2_X1 U9541 ( .A1(n10524), .A2(n7057), .ZN(n7051) );
  NAND3_X1 U9542 ( .A1(n7052), .A2(n7051), .A3(n7054), .ZN(n10627) );
  AOI21_X1 U9543 ( .B1(n12264), .B2(n7066), .A(n7061), .ZN(n7060) );
  NAND2_X1 U9544 ( .A1(n12272), .A2(n7066), .ZN(n7065) );
  NAND3_X1 U9545 ( .A1(n7065), .A2(n7068), .A3(n7064), .ZN(n12273) );
  INV_X2 U9546 ( .A(n10566), .ZN(n12833) );
  XNOR2_X1 U9547 ( .A(n11983), .B(n10566), .ZN(n10611) );
  NAND2_X1 U9548 ( .A1(n11923), .A2(n6585), .ZN(n7101) );
  NAND2_X1 U9549 ( .A1(n9771), .A2(n9184), .ZN(n7107) );
  XNOR2_X1 U9550 ( .A(n15015), .B(n7107), .ZN(n15056) );
  NAND2_X1 U9551 ( .A1(n12486), .A2(n7110), .ZN(n7109) );
  NAND2_X1 U9552 ( .A1(n8968), .A2(n7115), .ZN(n7114) );
  NAND2_X1 U9553 ( .A1(n11090), .A2(n7120), .ZN(n7118) );
  INV_X1 U9554 ( .A(n7121), .ZN(n7120) );
  AOI21_X1 U9555 ( .B1(n12354), .B2(n7128), .A(n7127), .ZN(n9751) );
  NAND2_X1 U9556 ( .A1(n12443), .A2(n6581), .ZN(n12432) );
  AND4_X2 U9557 ( .A1(n8800), .A2(n8801), .A3(n8802), .A4(n8799), .ZN(n10786)
         );
  INV_X1 U9558 ( .A(n10611), .ZN(n12994) );
  NAND2_X1 U9559 ( .A1(n12394), .A2(n12393), .ZN(n12395) );
  NAND2_X1 U9560 ( .A1(n12190), .A2(n10791), .ZN(n9372) );
  NAND2_X1 U9561 ( .A1(n11135), .A2(n6483), .ZN(n7148) );
  NAND2_X1 U9562 ( .A1(n7148), .A2(n7149), .ZN(n11166) );
  AOI21_X1 U9563 ( .B1(n6483), .B2(n7151), .A(n6553), .ZN(n7149) );
  NAND2_X1 U9564 ( .A1(n13143), .A2(n7156), .ZN(n7154) );
  AOI21_X1 U9565 ( .B1(n13143), .B2(n13152), .A(n7152), .ZN(n13131) );
  INV_X1 U9566 ( .A(n7163), .ZN(n13157) );
  INV_X1 U9567 ( .A(n7620), .ZN(n7204) );
  NAND2_X1 U9568 ( .A1(n10933), .A2(n7170), .ZN(n7172) );
  NOR2_X1 U9569 ( .A1(n10932), .A2(n9692), .ZN(n7170) );
  NAND2_X1 U9570 ( .A1(n7172), .A2(n7171), .ZN(n11210) );
  NAND2_X1 U9571 ( .A1(n7178), .A2(n7177), .ZN(n7176) );
  OR2_X2 U9572 ( .A1(n14624), .A2(n14623), .ZN(n7178) );
  NAND2_X1 U9573 ( .A1(n7178), .A2(n8278), .ZN(n14604) );
  NAND2_X1 U9574 ( .A1(n7179), .A2(n9521), .ZN(n10371) );
  NAND2_X1 U9575 ( .A1(n14604), .A2(n14605), .ZN(n7179) );
  CLKBUF_X1 U9576 ( .A(n8295), .Z(n7180) );
  NAND2_X1 U9577 ( .A1(n13911), .A2(n7187), .ZN(n7190) );
  INV_X1 U9578 ( .A(n7190), .ZN(n13905) );
  CLKBUF_X1 U9579 ( .A(n7195), .Z(n7191) );
  INV_X1 U9580 ( .A(n7191), .ZN(n13951) );
  AND2_X1 U9581 ( .A1(n7626), .A2(n7203), .ZN(n7201) );
  OAI22_X2 U9582 ( .A1(n7210), .A2(n6504), .B1(n7212), .B2(n12885), .ZN(n12899) );
  INV_X1 U9583 ( .A(n12884), .ZN(n7212) );
  OAI22_X2 U9584 ( .A1(n7213), .A2(n6505), .B1(n7215), .B2(n12851), .ZN(n12856) );
  INV_X1 U9585 ( .A(n12850), .ZN(n7215) );
  INV_X1 U9586 ( .A(n12862), .ZN(n7217) );
  NAND2_X1 U9587 ( .A1(n12871), .A2(n7221), .ZN(n7220) );
  OAI22_X2 U9588 ( .A1(n6561), .A2(n7220), .B1(n12874), .B2(n7222), .ZN(n12878) );
  INV_X1 U9589 ( .A(n12873), .ZN(n7222) );
  NAND2_X1 U9590 ( .A1(n7223), .A2(n7225), .ZN(n12838) );
  NAND3_X1 U9591 ( .A1(n12832), .A2(n12831), .A3(n7224), .ZN(n7223) );
  OR2_X1 U9592 ( .A1(n7226), .A2(n12834), .ZN(n7224) );
  NAND2_X1 U9593 ( .A1(n12927), .A2(n6591), .ZN(n7227) );
  INV_X1 U9594 ( .A(n12682), .ZN(n7235) );
  AOI21_X1 U9595 ( .B1(n7235), .B2(n7238), .A(n6590), .ZN(n8217) );
  NAND2_X1 U9596 ( .A1(n12734), .A2(n6496), .ZN(n12673) );
  NAND2_X2 U9597 ( .A1(n10923), .A2(n10922), .ZN(n7248) );
  NAND2_X1 U9598 ( .A1(n12713), .A2(n7249), .ZN(n12659) );
  NAND2_X2 U9599 ( .A1(n7790), .A2(n7250), .ZN(n12836) );
  XNOR2_X1 U9600 ( .A(n7783), .B(n7782), .ZN(n9890) );
  NAND2_X1 U9601 ( .A1(n11342), .A2(n7256), .ZN(n7255) );
  AND2_X4 U9602 ( .A1(n8546), .A2(n9926), .ZN(n9674) );
  OAI211_X1 U9603 ( .C1(n14058), .C2(n14738), .A(n7263), .B(n7264), .ZN(
        P1_U3557) );
  NAND2_X1 U9604 ( .A1(n13956), .A2(n7267), .ZN(n13944) );
  NAND2_X1 U9605 ( .A1(n7276), .A2(n6520), .ZN(n8679) );
  NAND2_X1 U9606 ( .A1(n11822), .A2(n7278), .ZN(n7276) );
  NAND2_X1 U9607 ( .A1(n8918), .A2(n7291), .ZN(n7289) );
  NAND2_X1 U9608 ( .A1(n7289), .A2(n7287), .ZN(n8718) );
  NAND2_X1 U9609 ( .A1(n7299), .A2(n7297), .ZN(n9009) );
  OAI21_X1 U9610 ( .B1(n8723), .B2(n6611), .A(n8725), .ZN(n7298) );
  NAND2_X1 U9611 ( .A1(n8985), .A2(n7300), .ZN(n7299) );
  NAND2_X1 U9612 ( .A1(n7303), .A2(n7304), .ZN(n8738) );
  NAND2_X1 U9613 ( .A1(n8734), .A2(n6498), .ZN(n7303) );
  NAND2_X1 U9614 ( .A1(n9042), .A2(n8730), .ZN(n7309) );
  NAND2_X1 U9615 ( .A1(n7309), .A2(n7311), .ZN(n8731) );
  NAND2_X1 U9616 ( .A1(n7316), .A2(n8702), .ZN(n7315) );
  INV_X1 U9617 ( .A(n8701), .ZN(n7316) );
  NAND3_X1 U9618 ( .A1(n8809), .A2(n8810), .A3(n8702), .ZN(n7317) );
  NAND2_X1 U9619 ( .A1(n8808), .A2(n8701), .ZN(n8793) );
  NAND2_X1 U9620 ( .A1(n8809), .A2(n8810), .ZN(n8808) );
  NOR2_X1 U9621 ( .A1(n15031), .A2(n10315), .ZN(n7332) );
  NAND2_X1 U9622 ( .A1(n11966), .A2(n7337), .ZN(n11965) );
  NAND3_X1 U9623 ( .A1(n7339), .A2(n12100), .A3(n9824), .ZN(n12035) );
  INV_X1 U9624 ( .A(n9816), .ZN(n9814) );
  INV_X1 U9625 ( .A(n7356), .ZN(n11483) );
  OAI21_X1 U9626 ( .B1(n7361), .B2(n7360), .A(n7357), .ZN(n10742) );
  NAND2_X1 U9627 ( .A1(n10364), .A2(n7358), .ZN(n7357) );
  NAND2_X1 U9628 ( .A1(n9026), .A2(n6606), .ZN(n9074) );
  NAND2_X1 U9629 ( .A1(n10149), .A2(n10150), .ZN(n7371) );
  INV_X1 U9630 ( .A(n10162), .ZN(n7370) );
  NAND2_X1 U9631 ( .A1(n10265), .A2(n10162), .ZN(n7369) );
  NAND2_X1 U9632 ( .A1(n10266), .A2(n10265), .ZN(n10267) );
  NAND2_X1 U9633 ( .A1(n7370), .A2(n7371), .ZN(n10266) );
  NAND2_X1 U9634 ( .A1(n11262), .A2(n7375), .ZN(n7374) );
  NAND2_X1 U9635 ( .A1(n13728), .A2(n7382), .ZN(n7381) );
  OAI211_X1 U9636 ( .C1(n13728), .C2(n7386), .A(n7383), .B(n7381), .ZN(n13639)
         );
  NAND2_X2 U9637 ( .A1(n10023), .A2(n10019), .ZN(n13629) );
  AND2_X1 U9638 ( .A1(n15033), .A2(n14917), .ZN(n15037) );
  NAND2_X1 U9639 ( .A1(n7415), .A2(n7413), .ZN(n7539) );
  INV_X1 U9640 ( .A(n7414), .ZN(n7413) );
  NAND2_X1 U9641 ( .A1(n7899), .A2(n7423), .ZN(n7421) );
  NAND2_X1 U9642 ( .A1(n7436), .A2(n7434), .ZN(n11460) );
  NAND2_X1 U9643 ( .A1(n9225), .A2(n6586), .ZN(n12338) );
  INV_X1 U9644 ( .A(n8196), .ZN(n7608) );
  NAND2_X2 U9645 ( .A1(n14343), .A2(n14342), .ZN(n14341) );
  NAND3_X1 U9646 ( .A1(n9709), .A2(n7454), .A3(n7453), .ZN(n7452) );
  NAND3_X1 U9647 ( .A1(n6752), .A2(n8995), .A3(n8758), .ZN(n9241) );
  INV_X1 U9648 ( .A(n9644), .ZN(n7479) );
  NAND3_X1 U9649 ( .A1(n9628), .A2(n9627), .A3(n6594), .ZN(n7482) );
  INV_X1 U9650 ( .A(n9629), .ZN(n7483) );
  INV_X1 U9651 ( .A(n9618), .ZN(n7485) );
  INV_X1 U9652 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7487) );
  NAND2_X1 U9653 ( .A1(n8508), .A2(n8507), .ZN(n8616) );
  NAND2_X1 U9654 ( .A1(n8508), .A2(n6494), .ZN(n8634) );
  CLKBUF_X1 U9655 ( .A(n11979), .Z(n12708) );
  AOI21_X2 U9656 ( .B1(n11286), .B2(n10966), .A(n10965), .ZN(n11135) );
  INV_X1 U9657 ( .A(n8204), .ZN(n8167) );
  CLKBUF_X1 U9658 ( .A(n11574), .Z(n11579) );
  NAND2_X1 U9659 ( .A1(n7773), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U9660 ( .A1(n9239), .A2(n9238), .ZN(n12336) );
  INV_X1 U9661 ( .A(n12651), .ZN(n12652) );
  OAI21_X1 U9662 ( .B1(n9341), .B2(n9340), .A(n9339), .ZN(n9498) );
  XNOR2_X1 U9663 ( .A(n9318), .B(n10459), .ZN(n9341) );
  AOI21_X1 U9664 ( .B1(n12650), .B2(n12649), .A(n12759), .ZN(n12653) );
  INV_X1 U9665 ( .A(n13088), .ZN(n13393) );
  AND4_X4 U9666 ( .A1(n8836), .A2(n8835), .A3(n8834), .A4(n8833), .ZN(n15018)
         );
  NAND2_X1 U9667 ( .A1(n9184), .A2(n9361), .ZN(n9322) );
  AND4_X2 U9668 ( .A1(n8807), .A2(n8806), .A3(n8805), .A4(n8804), .ZN(n8829)
         );
  BUF_X4 U9669 ( .A(n8822), .Z(n9309) );
  INV_X1 U9670 ( .A(n8506), .ZN(n8508) );
  OR2_X1 U9671 ( .A1(n8550), .A2(n8280), .ZN(n8281) );
  NAND4_X2 U9672 ( .A1(n8876), .A2(n8875), .A3(n8874), .A4(n8873), .ZN(n12188)
         );
  NAND2_X1 U9673 ( .A1(n8817), .A2(n9926), .ZN(n8839) );
  INV_X1 U9674 ( .A(n11932), .ZN(n8255) );
  NAND2_X1 U9675 ( .A1(n8829), .A2(n10320), .ZN(n9184) );
  NOR2_X1 U9676 ( .A1(n9926), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12646) );
  CLKBUF_X1 U9677 ( .A(n12424), .Z(n12425) );
  INV_X1 U9678 ( .A(n11190), .ZN(n7897) );
  OR2_X1 U9679 ( .A1(n12020), .A2(n12638), .ZN(n7504) );
  OR2_X1 U9680 ( .A1(n12020), .A2(n12585), .ZN(n7505) );
  AND3_X2 U9681 ( .A1(n10283), .A2(n9278), .A3(n9277), .ZN(n15096) );
  AND2_X1 U9682 ( .A1(n9729), .A2(n9728), .ZN(n7506) );
  XNOR2_X1 U9683 ( .A(n13042), .B(n13023), .ZN(n7507) );
  INV_X1 U9684 ( .A(SI_26_), .ZN(n11852) );
  INV_X1 U9685 ( .A(n9692), .ZN(n10996) );
  AND2_X1 U9686 ( .A1(n12981), .A2(n12980), .ZN(n7508) );
  AND2_X1 U9687 ( .A1(n12178), .A2(n15035), .ZN(n7509) );
  OR2_X1 U9688 ( .A1(n7550), .A2(n9892), .ZN(n7510) );
  NAND2_X1 U9689 ( .A1(n7608), .A2(n7607), .ZN(n8195) );
  AND2_X1 U9690 ( .A1(n13159), .A2(n13156), .ZN(n7514) );
  INV_X1 U9691 ( .A(SI_20_), .ZN(n10659) );
  INV_X1 U9692 ( .A(n7746), .ZN(n7791) );
  INV_X1 U9693 ( .A(n11817), .ZN(n9737) );
  AND2_X1 U9694 ( .A1(n12799), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n7515) );
  INV_X1 U9695 ( .A(SI_23_), .ZN(n11322) );
  INV_X1 U9696 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11086) );
  INV_X1 U9697 ( .A(n9098), .ZN(n8735) );
  AND2_X1 U9698 ( .A1(n9926), .A2(P2_U3088), .ZN(n13450) );
  INV_X1 U9699 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n15119) );
  INV_X1 U9700 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7844) );
  INV_X1 U9701 ( .A(n9418), .ZN(n12515) );
  AND2_X1 U9702 ( .A1(n8261), .A2(n8260), .ZN(n7516) );
  INV_X1 U9703 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11087) );
  INV_X1 U9704 ( .A(n12904), .ZN(n13013) );
  NAND2_X1 U9705 ( .A1(n12659), .A2(n8082), .ZN(n12666) );
  AND2_X1 U9706 ( .A1(n9795), .A2(n9794), .ZN(n7519) );
  MUX2_X1 U9707 ( .A(n12808), .B(n12807), .S(n12814), .Z(n12810) );
  INV_X1 U9708 ( .A(n9532), .ZN(n9533) );
  NAND2_X1 U9709 ( .A1(n12847), .A2(n12846), .ZN(n12848) );
  NAND2_X1 U9710 ( .A1(n12870), .A2(n12869), .ZN(n12871) );
  INV_X1 U9711 ( .A(n9578), .ZN(n9579) );
  INV_X1 U9712 ( .A(n9585), .ZN(n9586) );
  OR4_X1 U9713 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n8646) );
  INV_X1 U9714 ( .A(n14980), .ZN(n9193) );
  INV_X1 U9715 ( .A(n13072), .ZN(n10347) );
  INV_X1 U9716 ( .A(n12378), .ZN(n9824) );
  INV_X1 U9717 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n9111) );
  NOR2_X1 U9718 ( .A1(n14981), .A2(n9193), .ZN(n14982) );
  INV_X1 U9719 ( .A(n7922), .ZN(n7760) );
  INV_X1 U9720 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8239) );
  INV_X1 U9721 ( .A(n8197), .ZN(n7607) );
  INV_X1 U9722 ( .A(n12482), .ZN(n9801) );
  NAND2_X1 U9723 ( .A1(n9814), .A2(n9813), .ZN(n9817) );
  INV_X1 U9724 ( .A(n12457), .ZN(n9070) );
  INV_X1 U9725 ( .A(n12429), .ZN(n9096) );
  INV_X1 U9726 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8758) );
  INV_X1 U9727 ( .A(n7737), .ZN(n12984) );
  INV_X1 U9728 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8094) );
  INV_X1 U9729 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15221) );
  NAND2_X1 U9730 ( .A1(n10613), .A2(n10611), .ZN(n10579) );
  NOR2_X1 U9731 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7639) );
  INV_X1 U9732 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n15104) );
  NOR2_X1 U9733 ( .A1(n14627), .A2(n10264), .ZN(n14616) );
  INV_X1 U9734 ( .A(P1_B_REG_SCAN_IN), .ZN(n8637) );
  INV_X1 U9735 ( .A(n9784), .ZN(n9785) );
  INV_X1 U9736 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n9062) );
  AND2_X1 U9737 ( .A1(n10459), .A2(n10661), .ZN(n9492) );
  OR2_X1 U9738 ( .A1(n9121), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9132) );
  INV_X1 U9739 ( .A(n11879), .ZN(n8774) );
  OR2_X1 U9740 ( .A1(n9159), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9161) );
  INV_X1 U9741 ( .A(n12376), .ZN(n9140) );
  NAND2_X2 U9742 ( .A1(n11033), .A2(n9230), .ZN(n9499) );
  INV_X1 U9743 ( .A(n11508), .ZN(n8967) );
  OR2_X1 U9744 ( .A1(n9492), .A2(n9499), .ZN(n9848) );
  OR2_X1 U9745 ( .A1(n9295), .A2(n11971), .ZN(n8782) );
  NAND2_X1 U9746 ( .A1(n10782), .A2(n9376), .ZN(n15002) );
  NAND2_X1 U9747 ( .A1(n14160), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8743) );
  AND2_X1 U9748 ( .A1(n7884), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7909) );
  NOR2_X1 U9749 ( .A1(n11942), .A2(n13106), .ZN(n7751) );
  INV_X1 U9750 ( .A(n9874), .ZN(n7780) );
  NOR2_X1 U9751 ( .A1(n8116), .A2(n12675), .ZN(n8115) );
  OR2_X1 U9752 ( .A1(n12975), .A2(n12974), .ZN(n12976) );
  OR2_X1 U9753 ( .A1(n8179), .A2(n7690), .ZN(n7719) );
  OR2_X1 U9754 ( .A1(n8095), .A2(n8094), .ZN(n8116) );
  NAND2_X1 U9755 ( .A1(n8032), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8074) );
  INV_X1 U9756 ( .A(n7734), .ZN(n7727) );
  INV_X1 U9757 ( .A(n13283), .ZN(n13277) );
  AND2_X1 U9758 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7679) );
  INV_X1 U9759 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8389) );
  INV_X1 U9760 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n8377) );
  INV_X1 U9761 ( .A(n11641), .ZN(n11638) );
  OR2_X1 U9762 ( .A1(n8515), .A2(n8253), .ZN(n8524) );
  INV_X1 U9763 ( .A(n8353), .ZN(n8304) );
  INV_X1 U9764 ( .A(n9645), .ZN(n14054) );
  INV_X1 U9765 ( .A(n14633), .ZN(n14387) );
  INV_X1 U9766 ( .A(n10476), .ZN(n8301) );
  NAND2_X1 U9767 ( .A1(n8277), .A2(n10167), .ZN(n9510) );
  INV_X1 U9768 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8617) );
  OR2_X1 U9769 ( .A1(n8385), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n8398) );
  INV_X1 U9770 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8227) );
  INV_X1 U9771 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14210) );
  OR2_X1 U9772 ( .A1(n9079), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9091) );
  OR2_X1 U9773 ( .A1(n11147), .A2(n11311), .ZN(n9783) );
  NOR2_X1 U9774 ( .A1(n9035), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U9775 ( .A1(n14968), .A2(n9785), .ZN(n9786) );
  OR2_X1 U9776 ( .A1(n8940), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8979) );
  INV_X1 U9777 ( .A(n14916), .ZN(n12172) );
  OR2_X1 U9778 ( .A1(n8766), .A2(n14333), .ZN(n12332) );
  INV_X1 U9779 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14191) );
  OR2_X1 U9780 ( .A1(n10392), .A2(n10400), .ZN(n10403) );
  INV_X1 U9781 ( .A(n12401), .ZN(n12404) );
  INV_X1 U9782 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8928) );
  NAND2_X1 U9783 ( .A1(n12640), .A2(n9870), .ZN(n10387) );
  INV_X1 U9784 ( .A(n10881), .ZN(n9230) );
  OR2_X1 U9785 ( .A1(n9295), .A2(n11875), .ZN(n8763) );
  OR2_X1 U9786 ( .A1(n9088), .A2(n7584), .ZN(n9109) );
  AND3_X1 U9787 ( .A1(n7335), .A2(n9758), .A3(n12639), .ZN(n9850) );
  INV_X1 U9788 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n12701) );
  AND2_X1 U9789 ( .A1(n11986), .A2(n7798), .ZN(n7799) );
  OR2_X1 U9790 ( .A1(n13126), .A2(n8167), .ZN(n7699) );
  AND2_X1 U9791 ( .A1(n8056), .A2(n8035), .ZN(n13290) );
  INV_X1 U9792 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n13073) );
  INV_X1 U9793 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11836) );
  INV_X1 U9794 ( .A(n13106), .ZN(n13089) );
  INV_X1 U9795 ( .A(n13036), .ZN(n12771) );
  AND2_X1 U9796 ( .A1(n12990), .A2(n12989), .ZN(n13242) );
  INV_X1 U9797 ( .A(n13010), .ZN(n11392) );
  OR2_X1 U9798 ( .A1(n10334), .A2(n11417), .ZN(n10569) );
  INV_X1 U9799 ( .A(n12824), .ZN(n14844) );
  INV_X1 U9800 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n7666) );
  OR2_X1 U9801 ( .A1(n8028), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n8050) );
  OR2_X1 U9802 ( .A1(n8390), .A2(n8389), .ZN(n8403) );
  NOR2_X1 U9803 ( .A1(n15248), .A2(n8569), .ZN(n8576) );
  INV_X1 U9804 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13694) );
  INV_X1 U9805 ( .A(n8561), .ZN(n8547) );
  INV_X1 U9806 ( .A(n14397), .ZN(n13737) );
  NOR2_X1 U9807 ( .A1(n8524), .A2(n13694), .ZN(n8534) );
  NAND2_X1 U9808 ( .A1(n8492), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8515) );
  INV_X1 U9809 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14182) );
  INV_X1 U9810 ( .A(n13942), .ZN(n8683) );
  INV_X1 U9811 ( .A(n14017), .ZN(n14019) );
  OR2_X1 U9812 ( .A1(n10014), .A2(n14159), .ZN(n14633) );
  INV_X1 U9813 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14229) );
  AOI22_X1 U9814 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14193), .B1(n14255), .B2(
        n14192), .ZN(n14194) );
  AND2_X1 U9815 ( .A1(n9841), .A2(n9840), .ZN(n14914) );
  AND2_X1 U9816 ( .A1(n9312), .A2(n9236), .ZN(n11958) );
  AND4_X1 U9817 ( .A1(n9040), .A2(n9039), .A3(n9038), .A4(n9037), .ZN(n12500)
         );
  INV_X1 U9818 ( .A(n14943), .ZN(n14922) );
  NOR2_X1 U9819 ( .A1(n10403), .A2(n10402), .ZN(n14923) );
  INV_X1 U9820 ( .A(n15019), .ZN(n15034) );
  AND2_X1 U9821 ( .A1(n15050), .A2(n14953), .ZN(n12520) );
  OR2_X1 U9822 ( .A1(n10387), .A2(n15030), .ZN(n9843) );
  NAND2_X1 U9823 ( .A1(n9767), .A2(n10661), .ZN(n15044) );
  OR2_X1 U9824 ( .A1(n9275), .A2(n12639), .ZN(n9278) );
  OR2_X1 U9825 ( .A1(n9295), .A2(n11701), .ZN(n9130) );
  INV_X1 U9826 ( .A(n15023), .ZN(n15030) );
  INV_X1 U9827 ( .A(n15052), .ZN(n15079) );
  INV_X1 U9828 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9010) );
  INV_X1 U9829 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8903) );
  NAND2_X1 U9830 ( .A1(n7851), .A2(n10797), .ZN(n10801) );
  INV_X1 U9831 ( .A(n13049), .ZN(n12730) );
  INV_X1 U9832 ( .A(n12751), .ZN(n14378) );
  NAND2_X1 U9833 ( .A1(n7687), .A2(n13226), .ZN(n14381) );
  INV_X1 U9834 ( .A(n14384), .ZN(n12770) );
  AND2_X1 U9835 ( .A1(n10089), .A2(n10088), .ZN(n14784) );
  INV_X1 U9836 ( .A(n14784), .ZN(n14813) );
  OAI21_X1 U9837 ( .B1(n10057), .B2(n10056), .A(n10055), .ZN(n10089) );
  INV_X1 U9838 ( .A(n11910), .ZN(n11911) );
  AND2_X1 U9839 ( .A1(n8150), .A2(n8165), .ZN(n13177) );
  INV_X1 U9840 ( .A(n13226), .ZN(n13289) );
  NAND2_X1 U9841 ( .A1(n10569), .A2(n8213), .ZN(n14891) );
  INV_X1 U9842 ( .A(n14851), .ZN(n14880) );
  NOR2_X1 U9843 ( .A1(n11046), .A2(n14832), .ZN(n11047) );
  OR2_X1 U9844 ( .A1(n7648), .A2(n13458), .ZN(n14828) );
  XNOR2_X1 U9845 ( .A(n7667), .B(n7666), .ZN(n11812) );
  AND2_X1 U9846 ( .A1(n7942), .A2(n7978), .ZN(n10538) );
  INV_X1 U9847 ( .A(n13464), .ZN(n9894) );
  AND4_X1 U9848 ( .A1(n8555), .A2(n8554), .A3(n8553), .A4(n8552), .ZN(n13642)
         );
  AND4_X1 U9849 ( .A1(n8466), .A2(n8465), .A3(n8464), .A4(n8463), .ZN(n14386)
         );
  NAND3_X2 U9850 ( .A1(n8263), .A2(n8262), .A3(n7516), .ZN(n10028) );
  INV_X1 U9851 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14193) );
  OR2_X1 U9852 ( .A1(n14493), .A2(n9975), .ZN(n14576) );
  OR3_X1 U9853 ( .A1(n14493), .A2(n6459), .A3(n14159), .ZN(n14572) );
  INV_X1 U9854 ( .A(n14572), .ZN(n14554) );
  INV_X1 U9855 ( .A(n14566), .ZN(n14582) );
  NAND2_X1 U9856 ( .A1(n14078), .A2(n7513), .ZN(n13913) );
  INV_X1 U9857 ( .A(n14640), .ZN(n14409) );
  INV_X1 U9858 ( .A(n14011), .ZN(n14644) );
  AOI21_X1 U9859 ( .B1(n10196), .B2(n9939), .A(n9938), .ZN(n11587) );
  AND2_X1 U9860 ( .A1(n14690), .A2(n14709), .ZN(n14442) );
  INV_X1 U9861 ( .A(n14630), .ZN(n14608) );
  INV_X1 U9862 ( .A(n14690), .ZN(n14712) );
  INV_X1 U9863 ( .A(n14442), .ZN(n14714) );
  OR2_X1 U9864 ( .A1(n14168), .A2(n14162), .ZN(n9936) );
  AND2_X1 U9865 ( .A1(n10400), .A2(n10399), .ZN(n14921) );
  INV_X1 U9866 ( .A(n9789), .ZN(n11671) );
  INV_X1 U9867 ( .A(n14914), .ZN(n12153) );
  AND2_X1 U9868 ( .A1(n9312), .A2(n9301), .ZN(n14332) );
  NAND2_X1 U9869 ( .A1(n9128), .A2(n9127), .ZN(n12378) );
  INV_X1 U9870 ( .A(n12514), .ZN(n12497) );
  INV_X1 U9871 ( .A(n11311), .ZN(n12187) );
  INV_X1 U9872 ( .A(n14921), .ZN(n14951) );
  INV_X1 U9873 ( .A(n14923), .ZN(n14940) );
  AND2_X1 U9874 ( .A1(n12484), .A2(n12483), .ZN(n12570) );
  OR2_X1 U9875 ( .A1(n9843), .A2(n15044), .ZN(n15012) );
  NAND2_X1 U9876 ( .A1(n10287), .A2(n15012), .ZN(n15050) );
  INV_X1 U9877 ( .A(n9280), .ZN(n9281) );
  NAND2_X1 U9878 ( .A1(n15096), .A2(n15023), .ZN(n12585) );
  INV_X1 U9879 ( .A(n15096), .ZN(n15094) );
  INV_X1 U9880 ( .A(n12155), .ZN(n12594) );
  INV_X1 U9881 ( .A(n12095), .ZN(n12623) );
  AND2_X1 U9882 ( .A1(n14365), .A2(n14364), .ZN(n14371) );
  AND2_X1 U9883 ( .A1(n9760), .A2(n9759), .ZN(n15080) );
  NAND2_X1 U9884 ( .A1(n9948), .A2(n12640), .ZN(n9957) );
  INV_X1 U9885 ( .A(n8775), .ZN(n11884) );
  INV_X1 U9886 ( .A(SI_25_), .ZN(n15233) );
  INV_X1 U9887 ( .A(SI_15_), .ZN(n10172) );
  INV_X1 U9888 ( .A(SI_11_), .ZN(n9952) );
  NAND2_X1 U9889 ( .A1(n12653), .A2(n12652), .ZN(n12658) );
  OR2_X1 U9890 ( .A1(n8222), .A2(n6516), .ZN(n8223) );
  INV_X1 U9891 ( .A(n12957), .ZN(n13044) );
  INV_X1 U9892 ( .A(n12887), .ZN(n13056) );
  OR2_X1 U9893 ( .A1(n14772), .A2(P2_U3088), .ZN(n14827) );
  OR2_X1 U9894 ( .A1(n10089), .A2(P2_U3088), .ZN(n14811) );
  NAND2_X1 U9895 ( .A1(n13248), .A2(n10562), .ZN(n13238) );
  NAND2_X1 U9896 ( .A1(n14912), .A2(n14891), .ZN(n13370) );
  INV_X1 U9897 ( .A(n14912), .ZN(n14910) );
  INV_X1 U9898 ( .A(n15282), .ZN(n14899) );
  NAND2_X1 U9899 ( .A1(n14835), .A2(n14828), .ZN(n14829) );
  INV_X1 U9900 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13448) );
  INV_X1 U9901 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11814) );
  INV_X1 U9902 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U9903 ( .A1(n10475), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14401) );
  INV_X1 U9904 ( .A(n14087), .ZN(n13950) );
  INV_X1 U9905 ( .A(n13635), .ZN(n13754) );
  OAI21_X1 U9906 ( .B1(n14006), .B2(n8530), .A(n8529), .ZN(n13763) );
  OR2_X1 U9907 ( .A1(n14493), .A2(n13783), .ZN(n14566) );
  INV_X1 U9908 ( .A(n14491), .ZN(n14585) );
  OR2_X1 U9909 ( .A1(n8696), .A2(n14023), .ZN(n14011) );
  OR2_X1 U9910 ( .A1(n14648), .A2(n14608), .ZN(n14032) );
  INV_X1 U9911 ( .A(n14740), .ZN(n14738) );
  INV_X1 U9912 ( .A(n14724), .ZN(n14722) );
  AND2_X2 U9913 ( .A1(n11588), .A2(n10199), .ZN(n14724) );
  INV_X1 U9914 ( .A(n9936), .ZN(n10194) );
  INV_X1 U9915 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11819) );
  INV_X1 U9916 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10777) );
  INV_X1 U9917 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10186) );
  NAND2_X1 U9918 ( .A1(n9925), .A2(P1_U3086), .ZN(n14171) );
  AND2_X2 U9919 ( .A1(n12640), .A2(n9871), .ZN(P3_U3897) );
  NOR2_X1 U9920 ( .A1(n10057), .A2(n9869), .ZN(P2_U3947) );
  AND2_X2 U9921 ( .A1(n9937), .A2(n10018), .ZN(P1_U4016) );
  MUX2_X1 U9922 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n7524), .Z(n7593) );
  AND2_X1 U9923 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n7521) );
  NAND2_X1 U9924 ( .A1(n7522), .A2(n7521), .ZN(n8275) );
  INV_X1 U9925 ( .A(SI_1_), .ZN(n9914) );
  INV_X1 U9926 ( .A(n7757), .ZN(n7525) );
  NAND2_X1 U9927 ( .A1(n7526), .A2(n7525), .ZN(n7529) );
  NAND2_X1 U9928 ( .A1(n7527), .A2(SI_2_), .ZN(n7528) );
  XNOR2_X1 U9929 ( .A(n7531), .B(SI_3_), .ZN(n7769) );
  INV_X1 U9930 ( .A(n7769), .ZN(n7530) );
  NAND2_X1 U9931 ( .A1(n7531), .A2(SI_3_), .ZN(n7532) );
  NAND2_X1 U9932 ( .A1(n7534), .A2(SI_4_), .ZN(n7535) );
  MUX2_X1 U9933 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9926), .Z(n7537) );
  INV_X1 U9934 ( .A(n7803), .ZN(n7536) );
  NAND2_X1 U9935 ( .A1(n7537), .A2(SI_5_), .ZN(n7538) );
  NAND2_X1 U9936 ( .A1(n7823), .A2(n7540), .ZN(n7543) );
  NAND2_X1 U9937 ( .A1(n7541), .A2(SI_6_), .ZN(n7542) );
  MUX2_X1 U9938 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9926), .Z(n7545) );
  XNOR2_X1 U9939 ( .A(n7545), .B(SI_7_), .ZN(n7838) );
  INV_X1 U9940 ( .A(n7838), .ZN(n7544) );
  NAND2_X1 U9941 ( .A1(n7545), .A2(SI_7_), .ZN(n7546) );
  MUX2_X1 U9942 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9926), .Z(n7548) );
  XNOR2_X1 U9943 ( .A(n7548), .B(SI_8_), .ZN(n7856) );
  INV_X1 U9944 ( .A(n7856), .ZN(n7547) );
  NAND2_X1 U9945 ( .A1(n7548), .A2(SI_8_), .ZN(n7549) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9926), .Z(n7877) );
  INV_X1 U9947 ( .A(n7877), .ZN(n7550) );
  NAND2_X1 U9948 ( .A1(n7550), .A2(n9892), .ZN(n7551) );
  NAND2_X1 U9949 ( .A1(n7552), .A2(SI_10_), .ZN(n7553) );
  OAI21_X1 U9950 ( .B1(n7552), .B2(SI_10_), .A(n7553), .ZN(n7900) );
  MUX2_X1 U9951 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9926), .Z(n7554) );
  XNOR2_X1 U9952 ( .A(n7554), .B(SI_11_), .ZN(n7918) );
  INV_X1 U9953 ( .A(n7554), .ZN(n7555) );
  MUX2_X1 U9954 ( .A(n10186), .B(n10184), .S(n9926), .Z(n7556) );
  XNOR2_X1 U9955 ( .A(n7556), .B(SI_12_), .ZN(n7936) );
  MUX2_X1 U9956 ( .A(n10274), .B(n7301), .S(n9926), .Z(n7557) );
  XNOR2_X1 U9957 ( .A(n7557), .B(SI_13_), .ZN(n7959) );
  NAND2_X1 U9958 ( .A1(n7557), .A2(n9969), .ZN(n7558) );
  MUX2_X1 U9959 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9926), .Z(n7991) );
  INV_X1 U9960 ( .A(n7991), .ZN(n7976) );
  MUX2_X1 U9961 ( .A(n10589), .B(n10558), .S(n9926), .Z(n7993) );
  INV_X1 U9962 ( .A(n7993), .ZN(n7559) );
  NAND2_X1 U9963 ( .A1(n7559), .A2(SI_15_), .ZN(n7562) );
  OAI21_X1 U9964 ( .B1(n10099), .B2(n7976), .A(n7562), .ZN(n7560) );
  INV_X1 U9965 ( .A(n7560), .ZN(n7561) );
  NOR2_X1 U9966 ( .A1(n7991), .A2(SI_14_), .ZN(n7563) );
  AOI22_X1 U9967 ( .A1(n7563), .A2(n7562), .B1(n10172), .B2(n7993), .ZN(n7564)
         );
  MUX2_X1 U9968 ( .A(n10441), .B(n10461), .S(n9926), .Z(n7565) );
  NAND2_X1 U9969 ( .A1(n7565), .A2(n10246), .ZN(n7566) );
  MUX2_X1 U9970 ( .A(n10559), .B(n15219), .S(n9926), .Z(n7567) );
  NAND2_X1 U9971 ( .A1(n7567), .A2(n10327), .ZN(n7568) );
  INV_X1 U9972 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10749) );
  MUX2_X1 U9973 ( .A(n10777), .B(n10749), .S(n9926), .Z(n8045) );
  MUX2_X1 U9974 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9926), .Z(n7574) );
  XNOR2_X1 U9975 ( .A(n7574), .B(SI_19_), .ZN(n8068) );
  INV_X1 U9976 ( .A(n7574), .ZN(n7575) );
  MUX2_X1 U9977 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n9926), .Z(n8088) );
  MUX2_X1 U9978 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n7524), .Z(n7578) );
  INV_X1 U9979 ( .A(n7577), .ZN(n7580) );
  OAI21_X1 U9980 ( .B1(SI_21_), .B2(n7578), .A(n7583), .ZN(n8107) );
  INV_X1 U9981 ( .A(n8107), .ZN(n8109) );
  AND2_X1 U9982 ( .A1(n8109), .A2(SI_22_), .ZN(n7579) );
  INV_X1 U9983 ( .A(SI_22_), .ZN(n7584) );
  INV_X1 U9984 ( .A(n7587), .ZN(n7585) );
  OR2_X1 U9985 ( .A1(n7585), .A2(n8109), .ZN(n7588) );
  AND2_X1 U9986 ( .A1(n8088), .A2(n7588), .ZN(n7586) );
  NAND2_X1 U9987 ( .A1(n8087), .A2(n7586), .ZN(n7589) );
  MUX2_X1 U9988 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9926), .Z(n8130) );
  OAI21_X1 U9989 ( .B1(n7593), .B2(n7592), .A(n7595), .ZN(n8144) );
  INV_X1 U9990 ( .A(n8144), .ZN(n7594) );
  NAND2_X1 U9991 ( .A1(n8143), .A2(n7595), .ZN(n8158) );
  MUX2_X1 U9992 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9926), .Z(n7596) );
  NAND2_X1 U9993 ( .A1(n7596), .A2(SI_24_), .ZN(n7598) );
  OAI21_X1 U9994 ( .B1(SI_24_), .B2(n7596), .A(n7598), .ZN(n8159) );
  INV_X1 U9995 ( .A(n8159), .ZN(n7597) );
  MUX2_X1 U9996 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9926), .Z(n7600) );
  XNOR2_X1 U9997 ( .A(n7600), .B(SI_25_), .ZN(n8176) );
  INV_X1 U9998 ( .A(n8176), .ZN(n7599) );
  INV_X1 U9999 ( .A(n7600), .ZN(n7601) );
  NAND2_X1 U10000 ( .A1(n7601), .A2(n15233), .ZN(n7602) );
  INV_X1 U10001 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13457) );
  MUX2_X1 U10002 ( .A(n14164), .B(n13457), .S(n9926), .Z(n7730) );
  INV_X1 U10003 ( .A(n7730), .ZN(n7603) );
  INV_X1 U10004 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14160) );
  INV_X1 U10005 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13455) );
  MUX2_X1 U10006 ( .A(n14160), .B(n13455), .S(n9926), .Z(n7604) );
  INV_X1 U10007 ( .A(SI_27_), .ZN(n11971) );
  NAND2_X1 U10008 ( .A1(n7604), .A2(n11971), .ZN(n7609) );
  INV_X1 U10009 ( .A(n7604), .ZN(n7605) );
  NAND2_X1 U10010 ( .A1(n7605), .A2(SI_27_), .ZN(n7606) );
  NAND2_X1 U10011 ( .A1(n7609), .A2(n7606), .ZN(n8197) );
  INV_X1 U10012 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13453) );
  MUX2_X1 U10013 ( .A(n14157), .B(n13453), .S(n9926), .Z(n7610) );
  INV_X1 U10014 ( .A(SI_28_), .ZN(n11875) );
  NAND2_X1 U10015 ( .A1(n7610), .A2(n11875), .ZN(n8611) );
  INV_X1 U10016 ( .A(n7610), .ZN(n7611) );
  NAND2_X1 U10017 ( .A1(n7611), .A2(SI_28_), .ZN(n7612) );
  NAND4_X1 U10018 ( .A1(n7617), .A2(n7616), .A3(n7615), .A4(n7614), .ZN(n7618)
         );
  NAND2_X1 U10019 ( .A1(n7680), .A2(n7619), .ZN(n7625) );
  NOR2_X1 U10020 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n7624) );
  NOR2_X1 U10021 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n7623) );
  INV_X1 U10022 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7621) );
  NAND4_X1 U10023 ( .A1(n7624), .A2(n7623), .A3(n7622), .A4(n7621), .ZN(n7629)
         );
  NOR3_X1 U10024 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n7626) );
  NOR2_X1 U10025 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n7627) );
  AOI21_X1 U10026 ( .B1(n7629), .B2(n7628), .A(n7627), .ZN(n7630) );
  AND2_X1 U10027 ( .A1(n7633), .A2(n7630), .ZN(n7631) );
  INV_X1 U10028 ( .A(n7692), .ZN(n7636) );
  NAND2_X1 U10029 ( .A1(n14156), .A2(n12782), .ZN(n7638) );
  INV_X4 U10030 ( .A(n7922), .ZN(n12799) );
  NAND2_X1 U10031 ( .A1(n12799), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7637) );
  NAND2_X1 U10032 ( .A1(n7669), .A2(n7639), .ZN(n7665) );
  NAND2_X1 U10033 ( .A1(n7645), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7640) );
  NAND2_X1 U10034 ( .A1(n7641), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7642) );
  MUX2_X1 U10035 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7642), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n7643) );
  XOR2_X1 U10036 ( .A(P2_B_REG_SCAN_IN), .B(n11846), .Z(n7644) );
  NOR2_X1 U10037 ( .A1(n13461), .A2(n7644), .ZN(n7648) );
  NAND2_X1 U10038 ( .A1(n13458), .A2(n11846), .ZN(n7649) );
  INV_X1 U10039 ( .A(n14831), .ZN(n7661) );
  NOR4_X1 U10040 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n7653) );
  NOR4_X1 U10041 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n7652) );
  NOR4_X1 U10042 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n7651) );
  NOR4_X1 U10043 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n7650) );
  NAND4_X1 U10044 ( .A1(n7653), .A2(n7652), .A3(n7651), .A4(n7650), .ZN(n7660)
         );
  NOR2_X1 U10045 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .ZN(
        n7657) );
  NOR4_X1 U10046 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n7656) );
  NOR4_X1 U10047 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n7655) );
  NOR4_X1 U10048 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n7654) );
  NAND4_X1 U10049 ( .A1(n7657), .A2(n7656), .A3(n7655), .A4(n7654), .ZN(n7659)
         );
  INV_X1 U10050 ( .A(n14828), .ZN(n7658) );
  OAI21_X1 U10051 ( .B1(n7660), .B2(n7659), .A(n7658), .ZN(n10344) );
  NAND2_X1 U10052 ( .A1(n7661), .A2(n10344), .ZN(n7711) );
  INV_X1 U10053 ( .A(n7711), .ZN(n7668) );
  INV_X1 U10054 ( .A(n13458), .ZN(n7662) );
  INV_X1 U10055 ( .A(n11846), .ZN(n7663) );
  NAND2_X1 U10056 ( .A1(n7663), .A2(n13461), .ZN(n7664) );
  NAND2_X1 U10057 ( .A1(n7665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7667) );
  INV_X1 U10058 ( .A(n14835), .ZN(n14832) );
  NOR2_X1 U10059 ( .A1(n14834), .A2(n14832), .ZN(n10330) );
  NAND2_X1 U10060 ( .A1(n7668), .A2(n10330), .ZN(n8215) );
  XNOR2_X2 U10061 ( .A(n7671), .B(n7670), .ZN(n7735) );
  INV_X1 U10062 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7672) );
  NAND2_X1 U10063 ( .A1(n7735), .A2(n11515), .ZN(n10334) );
  XNOR2_X2 U10064 ( .A(n7677), .B(n7676), .ZN(n11417) );
  OR2_X1 U10065 ( .A1(n8215), .A2(n10569), .ZN(n7687) );
  NAND2_X1 U10066 ( .A1(n8028), .A2(n7679), .ZN(n7684) );
  NAND2_X1 U10067 ( .A1(n7680), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n7682) );
  XNOR2_X1 U10068 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_19__SCAN_IN), .ZN(
        n7681) );
  NAND2_X1 U10069 ( .A1(n7682), .A2(n7681), .ZN(n7683) );
  AND3_X2 U10070 ( .A1(n7685), .A2(n7684), .A3(n7683), .ZN(n12979) );
  NAND2_X1 U10071 ( .A1(n11417), .A2(n12979), .ZN(n12791) );
  INV_X1 U10072 ( .A(n12791), .ZN(n13030) );
  OR2_X1 U10073 ( .A1(n14895), .A2(n13029), .ZN(n10343) );
  INV_X1 U10074 ( .A(n10343), .ZN(n7686) );
  NAND2_X1 U10075 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7810) );
  NOR2_X1 U10076 ( .A1(n7810), .A2(n12701), .ZN(n7809) );
  NAND2_X1 U10077 ( .A1(n7809), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7845) );
  INV_X1 U10078 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7885) );
  NOR2_X1 U10079 ( .A1(n7886), .A2(n7885), .ZN(n7884) );
  AND2_X1 U10080 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n7688) );
  NAND2_X1 U10081 ( .A1(n7948), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7983) );
  INV_X1 U10082 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7982) );
  INV_X1 U10083 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8017) );
  INV_X1 U10084 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8073) );
  INV_X1 U10085 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12675) );
  AND2_X1 U10086 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n7689) );
  NAND2_X1 U10087 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n7690) );
  INV_X1 U10088 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12655) );
  NOR2_X1 U10089 ( .A1(n7719), .A2(n12655), .ZN(n7700) );
  INV_X1 U10090 ( .A(n7700), .ZN(n7708) );
  NAND2_X1 U10091 ( .A1(n7719), .A2(n12655), .ZN(n7691) );
  NAND2_X1 U10092 ( .A1(n7708), .A2(n7691), .ZN(n13126) );
  NAND2_X1 U10093 ( .A1(n7692), .A2(n6469), .ZN(n13441) );
  AND2_X4 U10094 ( .A1(n7693), .A2(n7694), .ZN(n8204) );
  INV_X1 U10095 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13125) );
  INV_X2 U10096 ( .A(n7791), .ZN(n12786) );
  NAND2_X1 U10097 ( .A1(n12786), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7696) );
  NAND2_X1 U10098 ( .A1(n7773), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7695) );
  OAI211_X1 U10099 ( .C1(n12790), .C2(n13125), .A(n7696), .B(n7695), .ZN(n7697) );
  INV_X1 U10100 ( .A(n7697), .ZN(n7698) );
  INV_X1 U10101 ( .A(n10058), .ZN(n10059) );
  NAND2_X1 U10102 ( .A1(n13045), .A2(n13036), .ZN(n7706) );
  AND2_X1 U10103 ( .A1(n7700), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n11914) );
  INV_X1 U10104 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U10105 ( .A1(n12786), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n7702) );
  NAND2_X1 U10106 ( .A1(n12785), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7701) );
  OAI211_X1 U10107 ( .C1(n7703), .C2(n12790), .A(n7702), .B(n7701), .ZN(n7704)
         );
  AOI21_X1 U10108 ( .B1(n11914), .B2(n8204), .A(n7704), .ZN(n12795) );
  OR2_X1 U10109 ( .A1(n12795), .A2(n12773), .ZN(n7705) );
  AND2_X1 U10110 ( .A1(n7706), .A2(n7705), .ZN(n13102) );
  NAND2_X1 U10111 ( .A1(n11417), .A2(n13026), .ZN(n12982) );
  INV_X1 U10112 ( .A(n11914), .ZN(n7710) );
  INV_X1 U10113 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U10114 ( .A1(n7708), .A2(n7707), .ZN(n7709) );
  OAI21_X1 U10115 ( .B1(n7711), .B2(n14834), .A(n10343), .ZN(n7715) );
  INV_X1 U10116 ( .A(n10052), .ZN(n7713) );
  INV_X1 U10117 ( .A(n12982), .ZN(n7712) );
  OR2_X1 U10118 ( .A1(n7713), .A2(n7712), .ZN(n13034) );
  AND3_X1 U10119 ( .A1(n10057), .A2(n11812), .A3(n13034), .ZN(n7714) );
  NAND2_X1 U10120 ( .A1(n7715), .A2(n7714), .ZN(n10482) );
  NAND2_X1 U10121 ( .A1(n10482), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14384) );
  AOI22_X1 U10122 ( .A1(n13105), .A2(n12770), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n7716) );
  OAI21_X1 U10123 ( .B1(n13102), .B2(n12751), .A(n7716), .ZN(n8218) );
  INV_X1 U10124 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n7718) );
  INV_X1 U10125 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7717) );
  OAI21_X1 U10126 ( .B1(n8179), .B2(n7718), .A(n7717), .ZN(n7720) );
  NAND2_X1 U10127 ( .A1(n13135), .A2(n8204), .ZN(n7726) );
  INV_X1 U10128 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n7723) );
  NAND2_X1 U10129 ( .A1(n7773), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7722) );
  NAND2_X1 U10130 ( .A1(n12786), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7721) );
  OAI211_X1 U10131 ( .C1(n7723), .C2(n12790), .A(n7722), .B(n7721), .ZN(n7724)
         );
  INV_X1 U10132 ( .A(n7724), .ZN(n7725) );
  NAND2_X1 U10133 ( .A1(n7726), .A2(n7725), .ZN(n13046) );
  INV_X2 U10134 ( .A(n10334), .ZN(n7728) );
  NAND2_X4 U10135 ( .A1(n7728), .A2(n7727), .ZN(n13231) );
  NAND2_X1 U10136 ( .A1(n13046), .A2(n13089), .ZN(n8191) );
  INV_X1 U10137 ( .A(n8191), .ZN(n8194) );
  XNOR2_X1 U10138 ( .A(n7730), .B(SI_26_), .ZN(n7731) );
  XNOR2_X1 U10139 ( .A(n7729), .B(n7731), .ZN(n13456) );
  NAND2_X1 U10140 ( .A1(n13456), .A2(n12782), .ZN(n7733) );
  NAND2_X1 U10141 ( .A1(n12799), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n7732) );
  XNOR2_X1 U10142 ( .A(n7735), .B(n7737), .ZN(n7736) );
  NAND2_X1 U10143 ( .A1(n7736), .A2(n13026), .ZN(n10335) );
  XNOR2_X1 U10144 ( .A(n13322), .B(n8210), .ZN(n8193) );
  NAND2_X1 U10145 ( .A1(n7746), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7739) );
  INV_X1 U10146 ( .A(n12790), .ZN(n7745) );
  NAND2_X1 U10147 ( .A1(n13231), .A2(n13070), .ZN(n7754) );
  XNOR2_X1 U10148 ( .A(n7741), .B(n7740), .ZN(n9897) );
  INV_X2 U10149 ( .A(n10053), .ZN(n8070) );
  NAND2_X1 U10150 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7742) );
  XNOR2_X1 U10151 ( .A(n7742), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10078) );
  INV_X1 U10152 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9898) );
  XNOR2_X1 U10153 ( .A(n7744), .B(n10355), .ZN(n7752) );
  NAND2_X1 U10154 ( .A1(n7773), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U10155 ( .A1(n8204), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U10156 ( .A1(n7745), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7748) );
  NAND2_X1 U10157 ( .A1(n7746), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7747) );
  XNOR2_X1 U10158 ( .A(n9882), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13465) );
  NOR2_X1 U10159 ( .A1(n7744), .A2(n10484), .ZN(n11940) );
  CLKBUF_X1 U10160 ( .A(n7752), .Z(n7753) );
  NAND2_X1 U10161 ( .A1(n7753), .A2(n7754), .ZN(n7755) );
  NAND2_X1 U10162 ( .A1(n10495), .A2(n7755), .ZN(n7764) );
  XNOR2_X1 U10163 ( .A(n7757), .B(n7756), .ZN(n9943) );
  OR2_X1 U10164 ( .A1(n7758), .A2(n7805), .ZN(n7759) );
  XNOR2_X1 U10165 ( .A(n7759), .B(P2_IR_REG_2__SCAN_IN), .ZN(n10080) );
  AOI22_X1 U10166 ( .A1(n7760), .A2(P1_DATAO_REG_2__SCAN_IN), .B1(n8070), .B2(
        n10080), .ZN(n7761) );
  XNOR2_X1 U10167 ( .A(n7744), .B(n12824), .ZN(n7765) );
  NAND2_X1 U10168 ( .A1(n7746), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7763) );
  NAND2_X1 U10169 ( .A1(n7773), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7762) );
  INV_X4 U10170 ( .A(n12790), .ZN(n11906) );
  NAND2_X1 U10171 ( .A1(n13231), .A2(n13069), .ZN(n7766) );
  XNOR2_X1 U10172 ( .A(n7765), .B(n7766), .ZN(n10494) );
  NAND2_X1 U10173 ( .A1(n7764), .A2(n10494), .ZN(n10489) );
  INV_X1 U10174 ( .A(n7765), .ZN(n7767) );
  NAND2_X1 U10175 ( .A1(n7767), .A2(n7766), .ZN(n7768) );
  INV_X1 U10176 ( .A(n9875), .ZN(n7781) );
  XNOR2_X1 U10177 ( .A(n7770), .B(n7769), .ZN(n9895) );
  NAND2_X1 U10178 ( .A1(n9895), .A2(n7901), .ZN(n7772) );
  NAND2_X1 U10179 ( .A1(n7620), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7771) );
  XNOR2_X1 U10180 ( .A(n7771), .B(P2_IR_REG_3__SCAN_IN), .ZN(n10083) );
  XNOR2_X1 U10181 ( .A(n7744), .B(n12833), .ZN(n7778) );
  INV_X1 U10182 ( .A(n7778), .ZN(n11982) );
  NAND2_X1 U10183 ( .A1(n7773), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7775) );
  INV_X1 U10184 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U10185 ( .A1(n8204), .A2(n10616), .ZN(n7774) );
  AND2_X1 U10186 ( .A1(n13231), .A2(n13068), .ZN(n7777) );
  INV_X1 U10187 ( .A(n7777), .ZN(n7776) );
  NAND2_X1 U10188 ( .A1(n11982), .A2(n7776), .ZN(n7779) );
  NAND2_X1 U10189 ( .A1(n7778), .A2(n7777), .ZN(n7798) );
  NAND2_X1 U10190 ( .A1(n7779), .A2(n7798), .ZN(n9874) );
  NAND2_X1 U10191 ( .A1(n7784), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7785) );
  MUX2_X1 U10192 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7785), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n7789) );
  INV_X1 U10193 ( .A(n7787), .ZN(n7788) );
  AOI22_X1 U10194 ( .A1(n12799), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8070), 
        .B2(n10086), .ZN(n7790) );
  XNOR2_X1 U10195 ( .A(n7744), .B(n12836), .ZN(n12705) );
  NAND2_X1 U10196 ( .A1(n7773), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7797) );
  NAND2_X1 U10197 ( .A1(n7746), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7796) );
  INV_X1 U10198 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n7792) );
  NAND2_X1 U10199 ( .A1(n10616), .A2(n7792), .ZN(n7793) );
  AND2_X1 U10200 ( .A1(n7793), .A2(n7810), .ZN(n11990) );
  NAND2_X1 U10201 ( .A1(n8204), .A2(n11990), .ZN(n7795) );
  NAND2_X1 U10202 ( .A1(n11906), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7794) );
  NAND4_X1 U10203 ( .A1(n7797), .A2(n7796), .A3(n7795), .A4(n7794), .ZN(n13067) );
  NAND2_X1 U10204 ( .A1(n13231), .A2(n13067), .ZN(n7800) );
  XNOR2_X1 U10205 ( .A(n12705), .B(n7800), .ZN(n11986) );
  NAND2_X1 U10206 ( .A1(n9873), .A2(n7799), .ZN(n11979) );
  INV_X1 U10207 ( .A(n7800), .ZN(n7801) );
  OR2_X1 U10208 ( .A1(n12705), .A2(n7801), .ZN(n7802) );
  NAND2_X1 U10209 ( .A1(n11979), .A2(n7802), .ZN(n7817) );
  XNOR2_X1 U10210 ( .A(n7804), .B(n7803), .ZN(n9899) );
  NAND2_X1 U10211 ( .A1(n9899), .A2(n7901), .ZN(n7808) );
  OR2_X1 U10212 ( .A1(n7787), .A2(n7805), .ZN(n7806) );
  XNOR2_X1 U10213 ( .A(n7806), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U10214 ( .A1(n12799), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8070), 
        .B2(n10110), .ZN(n7807) );
  NAND2_X1 U10215 ( .A1(n7808), .A2(n7807), .ZN(n12841) );
  XNOR2_X1 U10216 ( .A(n12841), .B(n8210), .ZN(n7818) );
  NAND2_X1 U10217 ( .A1(n12785), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7815) );
  NAND2_X1 U10218 ( .A1(n12786), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7814) );
  INV_X1 U10219 ( .A(n7809), .ZN(n7828) );
  NAND2_X1 U10220 ( .A1(n7810), .A2(n12701), .ZN(n7811) );
  AND2_X1 U10221 ( .A1(n7828), .A2(n7811), .ZN(n12704) );
  NAND2_X1 U10222 ( .A1(n8204), .A2(n12704), .ZN(n7813) );
  NAND2_X1 U10223 ( .A1(n11906), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7812) );
  NAND4_X1 U10224 ( .A1(n7815), .A2(n7814), .A3(n7813), .A4(n7812), .ZN(n13066) );
  NAND2_X1 U10225 ( .A1(n13231), .A2(n13066), .ZN(n7819) );
  INV_X1 U10226 ( .A(n7818), .ZN(n7820) );
  NAND2_X1 U10227 ( .A1(n7820), .A2(n7819), .ZN(n7821) );
  NAND2_X1 U10228 ( .A1(n7787), .A2(n7824), .ZN(n7840) );
  NAND2_X1 U10229 ( .A1(n7840), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7825) );
  XNOR2_X1 U10230 ( .A(n7825), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U10231 ( .A1(n12799), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8070), 
        .B2(n10126), .ZN(n7826) );
  NAND2_X1 U10232 ( .A1(n12786), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7832) );
  INV_X1 U10233 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U10234 ( .A1(n7828), .A2(n7827), .ZN(n7829) );
  AND2_X1 U10235 ( .A1(n7845), .A2(n7829), .ZN(n10904) );
  NAND2_X1 U10236 ( .A1(n8204), .A2(n10904), .ZN(n7831) );
  NAND2_X1 U10237 ( .A1(n11906), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7830) );
  AND2_X1 U10238 ( .A1(n13231), .A2(n13065), .ZN(n7834) );
  NAND2_X1 U10239 ( .A1(n7833), .A2(n7834), .ZN(n7837) );
  INV_X1 U10240 ( .A(n7833), .ZN(n10799) );
  INV_X1 U10241 ( .A(n7834), .ZN(n7835) );
  NAND2_X1 U10242 ( .A1(n10799), .A2(n7835), .ZN(n7836) );
  NAND2_X1 U10243 ( .A1(n10795), .A2(n7837), .ZN(n7851) );
  XNOR2_X1 U10244 ( .A(n7839), .B(n7838), .ZN(n9929) );
  NAND2_X1 U10245 ( .A1(n9929), .A2(n7901), .ZN(n7843) );
  NAND2_X1 U10246 ( .A1(n7858), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7841) );
  XNOR2_X1 U10247 ( .A(n7841), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U10248 ( .A1(n12799), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n8070), 
        .B2(n10216), .ZN(n7842) );
  NAND2_X1 U10249 ( .A1(n7843), .A2(n7842), .ZN(n12853) );
  XNOR2_X1 U10250 ( .A(n12853), .B(n8210), .ZN(n7854) );
  NAND2_X1 U10251 ( .A1(n12786), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7850) );
  NAND2_X1 U10252 ( .A1(n12785), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U10253 ( .A1(n7845), .A2(n7844), .ZN(n7846) );
  AND2_X1 U10254 ( .A1(n7867), .A2(n7846), .ZN(n11284) );
  NAND2_X1 U10255 ( .A1(n8204), .A2(n11284), .ZN(n7848) );
  NAND2_X1 U10256 ( .A1(n11906), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7847) );
  NAND4_X1 U10257 ( .A1(n7850), .A2(n7849), .A3(n7848), .A4(n7847), .ZN(n13064) );
  NAND2_X1 U10258 ( .A1(n13231), .A2(n13064), .ZN(n7852) );
  XNOR2_X1 U10259 ( .A(n7854), .B(n7852), .ZN(n10797) );
  INV_X1 U10260 ( .A(n7852), .ZN(n7853) );
  NAND2_X1 U10261 ( .A1(n7854), .A2(n7853), .ZN(n7855) );
  XNOR2_X1 U10262 ( .A(n7857), .B(n7856), .ZN(n9953) );
  NAND2_X1 U10263 ( .A1(n9953), .A2(n7901), .ZN(n7866) );
  NOR2_X1 U10264 ( .A1(n7858), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n7862) );
  INV_X1 U10265 ( .A(n7862), .ZN(n7859) );
  NAND2_X1 U10266 ( .A1(n7859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7860) );
  MUX2_X1 U10267 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7860), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n7863) );
  INV_X1 U10268 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U10269 ( .A1(n7862), .A2(n7861), .ZN(n7902) );
  NAND2_X1 U10270 ( .A1(n7863), .A2(n7902), .ZN(n13079) );
  OAI22_X1 U10271 ( .A1(n13079), .A2(n10053), .B1(n7922), .B2(n9954), .ZN(
        n7864) );
  INV_X1 U10272 ( .A(n7864), .ZN(n7865) );
  NAND2_X1 U10273 ( .A1(n7866), .A2(n7865), .ZN(n14885) );
  XNOR2_X1 U10274 ( .A(n14885), .B(n8201), .ZN(n7873) );
  NAND2_X1 U10275 ( .A1(n7773), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U10276 ( .A1(n12786), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7871) );
  NAND2_X1 U10277 ( .A1(n7867), .A2(n13073), .ZN(n7868) );
  NAND2_X1 U10278 ( .A1(n7886), .A2(n7868), .ZN(n10928) );
  INV_X1 U10279 ( .A(n10928), .ZN(n11140) );
  NAND2_X1 U10280 ( .A1(n8204), .A2(n11140), .ZN(n7870) );
  NAND2_X1 U10281 ( .A1(n11906), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7869) );
  NAND4_X1 U10282 ( .A1(n7872), .A2(n7871), .A3(n7870), .A4(n7869), .ZN(n13063) );
  NAND2_X1 U10283 ( .A1(n13231), .A2(n13063), .ZN(n7874) );
  NAND2_X1 U10284 ( .A1(n7873), .A2(n7874), .ZN(n10922) );
  INV_X1 U10285 ( .A(n7873), .ZN(n7876) );
  INV_X1 U10286 ( .A(n7874), .ZN(n7875) );
  NAND2_X1 U10287 ( .A1(n7876), .A2(n7875), .ZN(n10921) );
  XNOR2_X1 U10288 ( .A(n7877), .B(SI_9_), .ZN(n7878) );
  XNOR2_X1 U10289 ( .A(n7879), .B(n7878), .ZN(n9961) );
  NAND2_X1 U10290 ( .A1(n9961), .A2(n7901), .ZN(n7883) );
  NAND2_X1 U10291 ( .A1(n7902), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7880) );
  XNOR2_X1 U10292 ( .A(n7880), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U10293 ( .A1(n7922), .A2(n9963), .ZN(n7881) );
  AOI21_X1 U10294 ( .B1(n10222), .B2(n8070), .A(n7881), .ZN(n7882) );
  NAND2_X1 U10295 ( .A1(n7883), .A2(n7882), .ZN(n12865) );
  XNOR2_X1 U10296 ( .A(n12865), .B(n8201), .ZN(n7892) );
  NAND2_X1 U10297 ( .A1(n12785), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U10298 ( .A1(n12786), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7890) );
  INV_X1 U10299 ( .A(n7884), .ZN(n7910) );
  NAND2_X1 U10300 ( .A1(n7886), .A2(n7885), .ZN(n7887) );
  AND2_X1 U10301 ( .A1(n7910), .A2(n7887), .ZN(n11194) );
  NAND2_X1 U10302 ( .A1(n8204), .A2(n11194), .ZN(n7889) );
  NAND2_X1 U10303 ( .A1(n11906), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7888) );
  NAND4_X1 U10304 ( .A1(n7891), .A2(n7890), .A3(n7889), .A4(n7888), .ZN(n13062) );
  NAND2_X1 U10305 ( .A1(n13231), .A2(n13062), .ZN(n7893) );
  NAND2_X1 U10306 ( .A1(n7892), .A2(n7893), .ZN(n7898) );
  INV_X1 U10307 ( .A(n7892), .ZN(n7895) );
  INV_X1 U10308 ( .A(n7893), .ZN(n7894) );
  NAND2_X1 U10309 ( .A1(n7895), .A2(n7894), .ZN(n7896) );
  NAND2_X1 U10310 ( .A1(n7898), .A2(n7896), .ZN(n11190) );
  XNOR2_X1 U10311 ( .A(n7899), .B(n7430), .ZN(n9964) );
  NAND2_X1 U10312 ( .A1(n9964), .A2(n7901), .ZN(n7908) );
  OR2_X1 U10313 ( .A1(n7902), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7903) );
  NAND2_X1 U10314 ( .A1(n7903), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7905) );
  INV_X1 U10315 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U10316 ( .A1(n7905), .A2(n7904), .ZN(n7920) );
  OR2_X1 U10317 ( .A1(n7905), .A2(n7904), .ZN(n7906) );
  AOI22_X1 U10318 ( .A1(n10237), .A2(n8070), .B1(n12799), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n7907) );
  XNOR2_X1 U10319 ( .A(n14892), .B(n8201), .ZN(n7917) );
  NAND2_X1 U10320 ( .A1(n12785), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7915) );
  NAND2_X1 U10321 ( .A1(n12786), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7914) );
  INV_X1 U10322 ( .A(n7909), .ZN(n7947) );
  INV_X1 U10323 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n15103) );
  NAND2_X1 U10324 ( .A1(n7910), .A2(n15103), .ZN(n7911) );
  AND2_X1 U10325 ( .A1(n7947), .A2(n7911), .ZN(n11277) );
  NAND2_X1 U10326 ( .A1(n8204), .A2(n11277), .ZN(n7913) );
  NAND2_X1 U10327 ( .A1(n11906), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7912) );
  NAND4_X1 U10328 ( .A1(n7915), .A2(n7914), .A3(n7913), .A4(n7912), .ZN(n13061) );
  NAND2_X1 U10329 ( .A1(n13231), .A2(n13061), .ZN(n7916) );
  XNOR2_X1 U10330 ( .A(n7917), .B(n7916), .ZN(n11272) );
  XNOR2_X1 U10331 ( .A(n7919), .B(n7918), .ZN(n10035) );
  NAND2_X1 U10332 ( .A1(n10035), .A2(n12782), .ZN(n7925) );
  NAND2_X1 U10333 ( .A1(n7920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7921) );
  XNOR2_X1 U10334 ( .A(n7921), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10304) );
  NOR2_X1 U10335 ( .A1(n7922), .A2(n10037), .ZN(n7923) );
  AOI21_X1 U10336 ( .B1(n10304), .B2(n8070), .A(n7923), .ZN(n7924) );
  XNOR2_X1 U10337 ( .A(n12875), .B(n8201), .ZN(n7930) );
  NAND2_X1 U10338 ( .A1(n12785), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7929) );
  NAND2_X1 U10339 ( .A1(n12786), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7928) );
  XNOR2_X1 U10340 ( .A(n7947), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n11542) );
  NAND2_X1 U10341 ( .A1(n8204), .A2(n11542), .ZN(n7927) );
  NAND2_X1 U10342 ( .A1(n11906), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7926) );
  NAND4_X1 U10343 ( .A1(n7929), .A2(n7928), .A3(n7927), .A4(n7926), .ZN(n13060) );
  NAND2_X1 U10344 ( .A1(n13231), .A2(n13060), .ZN(n7931) );
  NAND2_X1 U10345 ( .A1(n7930), .A2(n7931), .ZN(n7935) );
  INV_X1 U10346 ( .A(n7930), .ZN(n7933) );
  INV_X1 U10347 ( .A(n7931), .ZN(n7932) );
  NAND2_X1 U10348 ( .A1(n7933), .A2(n7932), .ZN(n7934) );
  NAND2_X1 U10349 ( .A1(n7935), .A2(n7934), .ZN(n11540) );
  NAND2_X1 U10350 ( .A1(n11538), .A2(n7935), .ZN(n11574) );
  XNOR2_X1 U10351 ( .A(n7937), .B(n7936), .ZN(n10183) );
  NAND2_X1 U10352 ( .A1(n10183), .A2(n12782), .ZN(n7944) );
  INV_X1 U10353 ( .A(n7938), .ZN(n7939) );
  NAND2_X1 U10354 ( .A1(n7787), .A2(n7939), .ZN(n7941) );
  NAND2_X1 U10355 ( .A1(n7941), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7940) );
  MUX2_X1 U10356 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7940), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n7942) );
  AOI22_X1 U10357 ( .A1(n12799), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8070), 
        .B2(n10538), .ZN(n7943) );
  XNOR2_X1 U10358 ( .A(n12883), .B(n8201), .ZN(n7954) );
  NAND2_X1 U10359 ( .A1(n12785), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7953) );
  NAND2_X1 U10360 ( .A1(n12786), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7952) );
  INV_X1 U10361 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7946) );
  INV_X1 U10362 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7945) );
  OAI21_X1 U10363 ( .B1(n7947), .B2(n7946), .A(n7945), .ZN(n7949) );
  INV_X1 U10364 ( .A(n7948), .ZN(n7963) );
  AND2_X1 U10365 ( .A1(n7949), .A2(n7963), .ZN(n11580) );
  NAND2_X1 U10366 ( .A1(n8204), .A2(n11580), .ZN(n7951) );
  NAND2_X1 U10367 ( .A1(n11906), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7950) );
  NAND4_X1 U10368 ( .A1(n7953), .A2(n7952), .A3(n7951), .A4(n7950), .ZN(n13059) );
  NAND2_X1 U10369 ( .A1(n13231), .A2(n13059), .ZN(n7955) );
  AND2_X1 U10370 ( .A1(n7954), .A2(n7955), .ZN(n11575) );
  INV_X1 U10371 ( .A(n7954), .ZN(n7957) );
  INV_X1 U10372 ( .A(n7955), .ZN(n7956) );
  NAND2_X1 U10373 ( .A1(n7957), .A2(n7956), .ZN(n11576) );
  XNOR2_X1 U10374 ( .A(n7958), .B(n7959), .ZN(n10260) );
  NAND2_X1 U10375 ( .A1(n10260), .A2(n12782), .ZN(n7962) );
  NAND2_X1 U10376 ( .A1(n7978), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7960) );
  XNOR2_X1 U10377 ( .A(n7960), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11111) );
  AOI22_X1 U10378 ( .A1(n12799), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n11111), 
        .B2(n8070), .ZN(n7961) );
  XNOR2_X1 U10379 ( .A(n13386), .B(n8210), .ZN(n7969) );
  INV_X1 U10380 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11693) );
  NAND2_X1 U10381 ( .A1(n7963), .A2(n11693), .ZN(n7964) );
  AND2_X1 U10382 ( .A1(n7983), .A2(n7964), .ZN(n11696) );
  NAND2_X1 U10383 ( .A1(n11696), .A2(n8204), .ZN(n7968) );
  NAND2_X1 U10384 ( .A1(n12786), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7967) );
  NAND2_X1 U10385 ( .A1(n11906), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7966) );
  NAND2_X1 U10386 ( .A1(n12785), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7965) );
  NAND4_X1 U10387 ( .A1(n7968), .A2(n7967), .A3(n7966), .A4(n7965), .ZN(n13058) );
  AND2_X1 U10388 ( .A1(n13231), .A2(n13058), .ZN(n7970) );
  NAND2_X1 U10389 ( .A1(n7969), .A2(n7970), .ZN(n7974) );
  INV_X1 U10390 ( .A(n7969), .ZN(n7972) );
  INV_X1 U10391 ( .A(n7970), .ZN(n7971) );
  NAND2_X1 U10392 ( .A1(n7972), .A2(n7971), .ZN(n7973) );
  AND2_X1 U10393 ( .A1(n7974), .A2(n7973), .ZN(n11691) );
  XNOR2_X1 U10394 ( .A(n7975), .B(n10099), .ZN(n7992) );
  INV_X1 U10395 ( .A(n7992), .ZN(n7977) );
  XNOR2_X1 U10396 ( .A(n7977), .B(n7976), .ZN(n10423) );
  NAND2_X1 U10397 ( .A1(n10423), .A2(n12782), .ZN(n7981) );
  NAND2_X1 U10398 ( .A1(n7996), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7979) );
  XNOR2_X1 U10399 ( .A(n7979), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14803) );
  AOI22_X1 U10400 ( .A1(n12799), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n14803), 
        .B2(n8070), .ZN(n7980) );
  XNOR2_X1 U10401 ( .A(n12892), .B(n8210), .ZN(n7988) );
  NAND2_X1 U10402 ( .A1(n7983), .A2(n7982), .ZN(n7984) );
  NAND2_X1 U10403 ( .A1(n8000), .A2(n7984), .ZN(n14383) );
  AOI22_X1 U10404 ( .A1(n11906), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n12785), 
        .B2(P2_REG1_REG_14__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U10405 ( .A1(n12786), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7985) );
  OAI211_X1 U10406 ( .C1(n14383), .C2(n8167), .A(n7986), .B(n7985), .ZN(n13057) );
  NAND2_X1 U10407 ( .A1(n13231), .A2(n13057), .ZN(n7987) );
  XNOR2_X1 U10408 ( .A(n7988), .B(n7987), .ZN(n14374) );
  NAND2_X1 U10409 ( .A1(n7988), .A2(n7987), .ZN(n7989) );
  INV_X1 U10410 ( .A(n7975), .ZN(n7990) );
  OAI22_X1 U10411 ( .A1(n7992), .A2(n7991), .B1(n7990), .B2(SI_14_), .ZN(n7995) );
  XNOR2_X1 U10412 ( .A(n7993), .B(SI_15_), .ZN(n7994) );
  XNOR2_X1 U10413 ( .A(n7995), .B(n7994), .ZN(n10557) );
  NAND2_X1 U10414 ( .A1(n10557), .A2(n12782), .ZN(n7999) );
  OAI21_X1 U10415 ( .B1(n7996), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7997) );
  XNOR2_X1 U10416 ( .A(n7997), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U10417 ( .A1(n11441), .A2(n8070), .B1(n12799), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n7998) );
  XNOR2_X1 U10418 ( .A(n12886), .B(n8201), .ZN(n8006) );
  XNOR2_X1 U10419 ( .A(n8008), .B(n8006), .ZN(n11833) );
  NAND2_X1 U10420 ( .A1(n8000), .A2(n11836), .ZN(n8001) );
  AND2_X1 U10421 ( .A1(n8018), .A2(n8001), .ZN(n11840) );
  NAND2_X1 U10422 ( .A1(n11840), .A2(n8204), .ZN(n8004) );
  AOI22_X1 U10423 ( .A1(n12786), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n12785), 
        .B2(P2_REG1_REG_15__SCAN_IN), .ZN(n8003) );
  NAND2_X1 U10424 ( .A1(n11906), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8002) );
  NOR2_X1 U10425 ( .A1(n12887), .A2(n13106), .ZN(n8005) );
  INV_X1 U10426 ( .A(n8006), .ZN(n8007) );
  OR2_X1 U10427 ( .A1(n8008), .A2(n8007), .ZN(n8009) );
  XNOR2_X1 U10428 ( .A(n8010), .B(n8011), .ZN(n10440) );
  NAND2_X1 U10429 ( .A1(n10440), .A2(n12782), .ZN(n8015) );
  NAND2_X1 U10430 ( .A1(n7678), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8012) );
  MUX2_X1 U10431 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8012), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8013) );
  AOI22_X1 U10432 ( .A1(n12799), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8070), 
        .B2(n11739), .ZN(n8014) );
  XNOR2_X1 U10433 ( .A(n13372), .B(n8201), .ZN(n12720) );
  INV_X1 U10434 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11444) );
  INV_X1 U10435 ( .A(n8016), .ZN(n8034) );
  NAND2_X1 U10436 ( .A1(n8018), .A2(n8017), .ZN(n8019) );
  NAND2_X1 U10437 ( .A1(n8034), .A2(n8019), .ZN(n12696) );
  OR2_X1 U10438 ( .A1(n12696), .A2(n8167), .ZN(n8021) );
  AOI22_X1 U10439 ( .A1(n12786), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n12785), 
        .B2(P2_REG1_REG_16__SCAN_IN), .ZN(n8020) );
  OAI211_X1 U10440 ( .C1(n12790), .C2(n11444), .A(n8021), .B(n8020), .ZN(
        n13055) );
  NAND2_X1 U10441 ( .A1(n13055), .A2(n13089), .ZN(n8023) );
  XNOR2_X1 U10442 ( .A(n12720), .B(n8023), .ZN(n12692) );
  INV_X1 U10443 ( .A(n12692), .ZN(n8022) );
  NAND2_X1 U10444 ( .A1(n12720), .A2(n8023), .ZN(n8024) );
  NAND2_X1 U10445 ( .A1(n12689), .A2(n8024), .ZN(n8039) );
  XNOR2_X1 U10446 ( .A(n8025), .B(n8026), .ZN(n10556) );
  NAND2_X1 U10447 ( .A1(n10556), .A2(n12782), .ZN(n8031) );
  NAND2_X1 U10448 ( .A1(n8028), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8027) );
  MUX2_X1 U10449 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8027), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n8029) );
  AND2_X1 U10450 ( .A1(n8029), .A2(n8050), .ZN(n12006) );
  AOI22_X1 U10451 ( .A1(n12799), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n12006), 
        .B2(n8070), .ZN(n8030) );
  XNOR2_X1 U10452 ( .A(n13287), .B(n8201), .ZN(n8042) );
  INV_X1 U10453 ( .A(n8032), .ZN(n8056) );
  INV_X1 U10454 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U10455 ( .A1(n8034), .A2(n8033), .ZN(n8035) );
  INV_X1 U10456 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n15133) );
  NAND2_X1 U10457 ( .A1(n12785), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U10458 ( .A1(n11906), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8036) );
  OAI211_X1 U10459 ( .C1(n7791), .C2(n15133), .A(n8037), .B(n8036), .ZN(n8038)
         );
  AOI21_X1 U10460 ( .B1(n13290), .B2(n8204), .A(n8038), .ZN(n12755) );
  NOR2_X1 U10461 ( .A1(n12755), .A2(n13106), .ZN(n8040) );
  XNOR2_X1 U10462 ( .A(n8042), .B(n8040), .ZN(n12718) );
  INV_X1 U10463 ( .A(n8040), .ZN(n8041) );
  NAND2_X1 U10464 ( .A1(n8042), .A2(n8041), .ZN(n8043) );
  NAND2_X1 U10465 ( .A1(n8046), .A2(n8045), .ZN(n8047) );
  NAND2_X1 U10466 ( .A1(n8044), .A2(n8047), .ZN(n10778) );
  OR2_X1 U10467 ( .A1(n10778), .A2(n8131), .ZN(n8054) );
  NAND2_X1 U10468 ( .A1(n8050), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8048) );
  MUX2_X1 U10469 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8048), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n8049) );
  INV_X1 U10470 ( .A(n8049), .ZN(n8052) );
  NOR2_X1 U10471 ( .A1(n8050), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n8051) );
  NOR2_X1 U10472 ( .A1(n8052), .A2(n8051), .ZN(n12002) );
  AOI22_X1 U10473 ( .A1(n12002), .A2(n8070), .B1(n12799), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n8053) );
  XNOR2_X1 U10474 ( .A(n13269), .B(n8210), .ZN(n8063) );
  INV_X1 U10475 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8055) );
  NAND2_X1 U10476 ( .A1(n8056), .A2(n8055), .ZN(n8057) );
  NAND2_X1 U10477 ( .A1(n8074), .A2(n8057), .ZN(n13270) );
  OR2_X1 U10478 ( .A1(n13270), .A2(n8167), .ZN(n8062) );
  INV_X1 U10479 ( .A(n12785), .ZN(n8182) );
  INV_X1 U10480 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n14815) );
  NAND2_X1 U10481 ( .A1(n11906), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8059) );
  NAND2_X1 U10482 ( .A1(n12786), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8058) );
  OAI211_X1 U10483 ( .C1(n8182), .C2(n14815), .A(n8059), .B(n8058), .ZN(n8060)
         );
  INV_X1 U10484 ( .A(n8060), .ZN(n8061) );
  NAND2_X1 U10485 ( .A1(n8062), .A2(n8061), .ZN(n13053) );
  AND2_X1 U10486 ( .A1(n13053), .A2(n13231), .ZN(n8064) );
  NAND2_X1 U10487 ( .A1(n8063), .A2(n8064), .ZN(n8081) );
  INV_X1 U10488 ( .A(n8063), .ZN(n12660) );
  INV_X1 U10489 ( .A(n8064), .ZN(n8065) );
  NAND2_X1 U10490 ( .A1(n12660), .A2(n8065), .ZN(n8066) );
  NAND2_X1 U10491 ( .A1(n8081), .A2(n8066), .ZN(n12760) );
  INV_X1 U10492 ( .A(n12760), .ZN(n8067) );
  XNOR2_X1 U10493 ( .A(n8069), .B(n8068), .ZN(n11085) );
  NAND2_X1 U10494 ( .A1(n11085), .A2(n12782), .ZN(n8072) );
  AOI22_X1 U10495 ( .A1(n12799), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n12979), 
        .B2(n8070), .ZN(n8071) );
  XNOR2_X1 U10496 ( .A(n13251), .B(n8210), .ZN(n12737) );
  NAND2_X1 U10497 ( .A1(n8074), .A2(n8073), .ZN(n8075) );
  NAND2_X1 U10498 ( .A1(n8095), .A2(n8075), .ZN(n13252) );
  OR2_X1 U10499 ( .A1(n13252), .A2(n8167), .ZN(n8080) );
  INV_X1 U10500 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n15252) );
  NAND2_X1 U10501 ( .A1(n11906), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8077) );
  NAND2_X1 U10502 ( .A1(n12786), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8076) );
  OAI211_X1 U10503 ( .C1(n8182), .C2(n15252), .A(n8077), .B(n8076), .ZN(n8078)
         );
  INV_X1 U10504 ( .A(n8078), .ZN(n8079) );
  NAND2_X1 U10505 ( .A1(n8080), .A2(n8079), .ZN(n13052) );
  NAND2_X1 U10506 ( .A1(n13052), .A2(n13089), .ZN(n8083) );
  XNOR2_X1 U10507 ( .A(n12737), .B(n8083), .ZN(n12669) );
  AND2_X1 U10508 ( .A1(n12669), .A2(n8081), .ZN(n8082) );
  INV_X1 U10509 ( .A(n12737), .ZN(n8084) );
  NAND2_X1 U10510 ( .A1(n8084), .A2(n8083), .ZN(n8085) );
  NAND2_X1 U10511 ( .A1(n12666), .A2(n8085), .ZN(n8101) );
  INV_X1 U10512 ( .A(n8087), .ZN(n8090) );
  INV_X1 U10513 ( .A(n8088), .ZN(n8089) );
  NAND2_X1 U10514 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  NAND2_X1 U10515 ( .A1(n11416), .A2(n12782), .ZN(n8093) );
  NAND2_X1 U10516 ( .A1(n12799), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8092) );
  XNOR2_X1 U10517 ( .A(n13353), .B(n8210), .ZN(n8102) );
  NAND2_X1 U10518 ( .A1(n8095), .A2(n8094), .ZN(n8096) );
  NAND2_X1 U10519 ( .A1(n8116), .A2(n8096), .ZN(n13227) );
  INV_X1 U10520 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n13228) );
  NAND2_X1 U10521 ( .A1(n12785), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8098) );
  NAND2_X1 U10522 ( .A1(n12786), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8097) );
  OAI211_X1 U10523 ( .C1(n13228), .C2(n12790), .A(n8098), .B(n8097), .ZN(n8099) );
  INV_X1 U10524 ( .A(n8099), .ZN(n8100) );
  NAND2_X1 U10525 ( .A1(n12928), .A2(n13089), .ZN(n8103) );
  XNOR2_X1 U10526 ( .A(n8102), .B(n8103), .ZN(n12738) );
  INV_X1 U10527 ( .A(n8102), .ZN(n8104) );
  NAND2_X1 U10528 ( .A1(n8104), .A2(n8103), .ZN(n8105) );
  AND2_X1 U10529 ( .A1(n8086), .A2(n8106), .ZN(n8108) );
  NAND2_X1 U10530 ( .A1(n8108), .A2(n8107), .ZN(n8112) );
  INV_X1 U10531 ( .A(n8108), .ZN(n8110) );
  NAND2_X1 U10532 ( .A1(n8110), .A2(n8109), .ZN(n8111) );
  NAND2_X1 U10533 ( .A1(n12799), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8113) );
  XNOR2_X1 U10534 ( .A(n13212), .B(n8201), .ZN(n8124) );
  INV_X1 U10535 ( .A(n8115), .ZN(n8148) );
  NAND2_X1 U10536 ( .A1(n8116), .A2(n12675), .ZN(n8117) );
  AND2_X1 U10537 ( .A1(n8148), .A2(n8117), .ZN(n13213) );
  NAND2_X1 U10538 ( .A1(n13213), .A2(n8204), .ZN(n8122) );
  INV_X1 U10539 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n15128) );
  NAND2_X1 U10540 ( .A1(n12786), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8119) );
  NAND2_X1 U10541 ( .A1(n11906), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8118) );
  OAI211_X1 U10542 ( .C1(n8182), .C2(n15128), .A(n8119), .B(n8118), .ZN(n8120)
         );
  INV_X1 U10543 ( .A(n8120), .ZN(n8121) );
  NAND2_X1 U10544 ( .A1(n8122), .A2(n8121), .ZN(n13051) );
  NAND2_X1 U10545 ( .A1(n13051), .A2(n13089), .ZN(n8125) );
  XNOR2_X1 U10546 ( .A(n8124), .B(n8125), .ZN(n12671) );
  INV_X1 U10547 ( .A(n8124), .ZN(n8127) );
  INV_X1 U10548 ( .A(n8125), .ZN(n8126) );
  NAND2_X1 U10549 ( .A1(n8127), .A2(n8126), .ZN(n8128) );
  NAND2_X1 U10550 ( .A1(n12799), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8132) );
  XNOR2_X1 U10551 ( .A(n13194), .B(n8201), .ZN(n8139) );
  XNOR2_X1 U10552 ( .A(n8141), .B(n8139), .ZN(n12746) );
  XNOR2_X1 U10553 ( .A(n8148), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n13195) );
  NAND2_X1 U10554 ( .A1(n13195), .A2(n8204), .ZN(n8138) );
  INV_X1 U10555 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8135) );
  NAND2_X1 U10556 ( .A1(n12786), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8134) );
  NAND2_X1 U10557 ( .A1(n7773), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n8133) );
  OAI211_X1 U10558 ( .C1(n8135), .C2(n12790), .A(n8134), .B(n8133), .ZN(n8136)
         );
  INV_X1 U10559 ( .A(n8136), .ZN(n8137) );
  NAND2_X1 U10560 ( .A1(n8138), .A2(n8137), .ZN(n13050) );
  NAND2_X1 U10561 ( .A1(n13050), .A2(n13089), .ZN(n12745) );
  INV_X1 U10562 ( .A(n8139), .ZN(n8140) );
  NOR2_X1 U10563 ( .A1(n8141), .A2(n8140), .ZN(n8142) );
  NAND2_X1 U10564 ( .A1(n8144), .A2(n11322), .ZN(n8145) );
  NAND2_X1 U10565 ( .A1(n11816), .A2(n12782), .ZN(n8147) );
  NAND2_X1 U10566 ( .A1(n12799), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8146) );
  XNOR2_X1 U10567 ( .A(n13182), .B(n8210), .ZN(n8156) );
  INV_X1 U10568 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12750) );
  INV_X1 U10569 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n11973) );
  OAI21_X1 U10570 ( .B1(n8148), .B2(n12750), .A(n11973), .ZN(n8150) );
  INV_X1 U10571 ( .A(n8149), .ZN(n8165) );
  NAND2_X1 U10572 ( .A1(n13177), .A2(n8204), .ZN(n8155) );
  INV_X1 U10573 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n15246) );
  NAND2_X1 U10574 ( .A1(n12785), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8152) );
  NAND2_X1 U10575 ( .A1(n11906), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8151) );
  OAI211_X1 U10576 ( .C1(n7791), .C2(n15246), .A(n8152), .B(n8151), .ZN(n8153)
         );
  INV_X1 U10577 ( .A(n8153), .ZN(n8154) );
  NAND2_X1 U10578 ( .A1(n8155), .A2(n8154), .ZN(n13049) );
  INV_X1 U10579 ( .A(n8158), .ZN(n8160) );
  NAND2_X1 U10580 ( .A1(n8160), .A2(n8159), .ZN(n8162) );
  NAND2_X1 U10581 ( .A1(n11844), .A2(n12782), .ZN(n8164) );
  NAND2_X1 U10582 ( .A1(n12799), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8163) );
  XNOR2_X1 U10583 ( .A(n12946), .B(n8210), .ZN(n12680) );
  INV_X1 U10584 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n15225) );
  NAND2_X1 U10585 ( .A1(n8165), .A2(n15225), .ZN(n8166) );
  NAND2_X1 U10586 ( .A1(n8179), .A2(n8166), .ZN(n13165) );
  OR2_X1 U10587 ( .A1(n13165), .A2(n8167), .ZN(n8172) );
  INV_X1 U10588 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n15208) );
  NAND2_X1 U10589 ( .A1(n11906), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8169) );
  NAND2_X1 U10590 ( .A1(n12786), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8168) );
  OAI211_X1 U10591 ( .C1(n8182), .C2(n15208), .A(n8169), .B(n8168), .ZN(n8170)
         );
  INV_X1 U10592 ( .A(n8170), .ZN(n8171) );
  NAND2_X1 U10593 ( .A1(n8172), .A2(n8171), .ZN(n13048) );
  AND2_X1 U10594 ( .A1(n13048), .A2(n13231), .ZN(n8173) );
  NAND2_X1 U10595 ( .A1(n12680), .A2(n8173), .ZN(n8174) );
  OAI21_X1 U10596 ( .B1(n12680), .B2(n8173), .A(n8174), .ZN(n12727) );
  INV_X1 U10597 ( .A(n8174), .ZN(n8190) );
  XNOR2_X1 U10598 ( .A(n8175), .B(n8176), .ZN(n13460) );
  NAND2_X1 U10599 ( .A1(n13460), .A2(n12782), .ZN(n8178) );
  NAND2_X1 U10600 ( .A1(n12799), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8177) );
  XNOR2_X1 U10601 ( .A(n13327), .B(n8210), .ZN(n8186) );
  XNOR2_X1 U10602 ( .A(n8179), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n13149) );
  NAND2_X1 U10603 ( .A1(n13149), .A2(n8204), .ZN(n8185) );
  INV_X1 U10604 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n15249) );
  NAND2_X1 U10605 ( .A1(n12786), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8181) );
  NAND2_X1 U10606 ( .A1(n11906), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8180) );
  OAI211_X1 U10607 ( .C1(n15249), .C2(n8182), .A(n8181), .B(n8180), .ZN(n8183)
         );
  INV_X1 U10608 ( .A(n8183), .ZN(n8184) );
  NAND2_X1 U10609 ( .A1(n8185), .A2(n8184), .ZN(n13047) );
  AND2_X1 U10610 ( .A1(n13047), .A2(n13231), .ZN(n8187) );
  NAND2_X1 U10611 ( .A1(n8186), .A2(n8187), .ZN(n8192) );
  INV_X1 U10612 ( .A(n8186), .ZN(n12766) );
  INV_X1 U10613 ( .A(n8187), .ZN(n8188) );
  NAND2_X1 U10614 ( .A1(n12766), .A2(n8188), .ZN(n8189) );
  AND2_X1 U10615 ( .A1(n8192), .A2(n8189), .ZN(n12681) );
  XNOR2_X1 U10616 ( .A(n8193), .B(n8191), .ZN(n12780) );
  NAND2_X1 U10617 ( .A1(n8196), .A2(n8197), .ZN(n8198) );
  NAND2_X1 U10618 ( .A1(n8195), .A2(n8198), .ZN(n8225) );
  NAND2_X1 U10619 ( .A1(n8225), .A2(n12782), .ZN(n8200) );
  NAND2_X1 U10620 ( .A1(n12799), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8199) );
  XNOR2_X1 U10621 ( .A(n13402), .B(n8201), .ZN(n8219) );
  NOR2_X1 U10622 ( .A1(n12956), .A2(n13106), .ZN(n8202) );
  NAND2_X1 U10623 ( .A1(n8219), .A2(n8202), .ZN(n8203) );
  OAI21_X1 U10624 ( .B1(n8219), .B2(n8202), .A(n8203), .ZN(n12649) );
  INV_X1 U10625 ( .A(n8203), .ZN(n8216) );
  NAND2_X1 U10626 ( .A1(n13105), .A2(n8204), .ZN(n8209) );
  INV_X1 U10627 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n13110) );
  NAND2_X1 U10628 ( .A1(n7773), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U10629 ( .A1(n12786), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8205) );
  OAI211_X1 U10630 ( .C1(n13110), .C2(n12790), .A(n8206), .B(n8205), .ZN(n8207) );
  INV_X1 U10631 ( .A(n8207), .ZN(n8208) );
  OR2_X1 U10632 ( .A1(n12957), .A2(n13106), .ZN(n8211) );
  XNOR2_X1 U10633 ( .A(n8211), .B(n8210), .ZN(n8212) );
  OR2_X1 U10634 ( .A1(n10334), .A2(n13026), .ZN(n8213) );
  OR2_X1 U10635 ( .A1(n14891), .A2(n10052), .ZN(n8214) );
  INV_X1 U10636 ( .A(n8219), .ZN(n8220) );
  NAND2_X1 U10637 ( .A1(n14376), .A2(n13089), .ZN(n12765) );
  NOR3_X1 U10638 ( .A1(n8220), .A2(n12956), .A3(n12765), .ZN(n8221) );
  AOI21_X1 U10639 ( .B1(n12651), .B2(n14376), .A(n8221), .ZN(n8222) );
  NAND2_X1 U10640 ( .A1(n8224), .A2(n8223), .ZN(P2_U3192) );
  NOR2_X1 U10641 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8230) );
  NAND4_X1 U10642 ( .A1(n8230), .A2(n8229), .A3(n8228), .A4(n8412), .ZN(n8484)
         );
  NAND2_X1 U10643 ( .A1(n8232), .A2(n8231), .ZN(n8233) );
  NOR2_X1 U10644 ( .A1(n8484), .A2(n8233), .ZN(n8238) );
  NOR2_X1 U10645 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), 
        .ZN(n8235) );
  NOR2_X1 U10646 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8234) );
  NAND4_X1 U10647 ( .A1(n8235), .A2(n8234), .A3(n8509), .A4(n8617), .ZN(n8237)
         );
  NAND3_X1 U10648 ( .A1(n8456), .A2(n8470), .A3(n8236), .ZN(n8483) );
  NAND3_X1 U10649 ( .A1(n8486), .A2(n8238), .A3(n8625), .ZN(n8628) );
  OR2_X1 U10650 ( .A1(n8242), .A2(n8241), .ZN(n8243) );
  NAND2_X1 U10651 ( .A1(n8225), .A2(n9656), .ZN(n8246) );
  NAND2_X1 U10652 ( .A1(n9674), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U10653 ( .A1(n8247), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8249) );
  NAND2_X1 U10654 ( .A1(n8692), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8258) );
  INV_X1 U10655 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n15248) );
  AND3_X1 U10656 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U10657 ( .A1(n8337), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8351) );
  INV_X1 U10658 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8350) );
  NOR2_X1 U10659 ( .A1(n8351), .A2(n8350), .ZN(n8366) );
  NAND2_X1 U10660 ( .A1(n8366), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8378) );
  INV_X1 U10661 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10662 ( .A1(n8418), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U10663 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n8252) );
  NAND2_X1 U10664 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n8253) );
  NAND2_X1 U10665 ( .A1(n8534), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8548) );
  INV_X1 U10666 ( .A(n8548), .ZN(n8254) );
  NAND2_X1 U10667 ( .A1(n8254), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U10668 ( .A1(n8547), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8569) );
  NAND2_X1 U10669 ( .A1(n8576), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8587) );
  INV_X1 U10670 ( .A(n8587), .ZN(n8577) );
  NAND2_X1 U10671 ( .A1(n8577), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8586) );
  XNOR2_X1 U10672 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n8586), .ZN(n13902) );
  NAND2_X1 U10673 ( .A1(n8606), .A2(n13902), .ZN(n8257) );
  NAND2_X1 U10674 ( .A1(n9659), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8256) );
  NAND4_X1 U10675 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n13756) );
  INV_X1 U10676 ( .A(n13756), .ZN(n13634) );
  NAND2_X1 U10677 ( .A1(n8295), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10678 ( .A1(n9659), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U10679 ( .A1(n8353), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U10680 ( .A1(n8294), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8260) );
  INV_X1 U10681 ( .A(n10028), .ZN(n8277) );
  NAND2_X1 U10682 ( .A1(n8290), .A2(n9897), .ZN(n8271) );
  NAND2_X1 U10683 ( .A1(n9926), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8265) );
  AOI21_X1 U10684 ( .B1(n14159), .B2(n6459), .A(n8265), .ZN(n8270) );
  NAND2_X1 U10685 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8266) );
  MUX2_X1 U10686 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8266), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8269) );
  INV_X1 U10687 ( .A(n8267), .ZN(n8268) );
  INV_X1 U10688 ( .A(n9985), .ZN(n9993) );
  INV_X1 U10689 ( .A(SI_0_), .ZN(n8273) );
  INV_X1 U10690 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8272) );
  OAI21_X1 U10691 ( .B1(n9926), .B2(n8273), .A(n8272), .ZN(n8274) );
  NAND2_X1 U10692 ( .A1(n8275), .A2(n8274), .ZN(n14175) );
  INV_X1 U10693 ( .A(n14628), .ZN(n10203) );
  NAND2_X1 U10694 ( .A1(n10203), .A2(n10017), .ZN(n9509) );
  INV_X1 U10695 ( .A(n9509), .ZN(n14623) );
  NAND2_X1 U10696 ( .A1(n8277), .A2(n14652), .ZN(n8278) );
  NAND2_X1 U10697 ( .A1(n8294), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8283) );
  NAND2_X1 U10698 ( .A1(n8353), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n8282) );
  INV_X1 U10699 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8280) );
  NAND4_X2 U10700 ( .A1(n8284), .A2(n8283), .A3(n8282), .A4(n8281), .ZN(n13780) );
  NAND2_X1 U10701 ( .A1(n9674), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8288) );
  NOR2_X1 U10702 ( .A1(n8267), .A2(n8241), .ZN(n8285) );
  NAND2_X1 U10703 ( .A1(n9921), .A2(n13788), .ZN(n8287) );
  OAI211_X2 U10704 ( .C1(n8312), .C2(n9943), .A(n8288), .B(n8287), .ZN(n10264)
         );
  NAND2_X1 U10705 ( .A1(n13780), .A2(n10264), .ZN(n9519) );
  OR2_X1 U10706 ( .A1(n8314), .A2(n8241), .ZN(n8289) );
  XNOR2_X1 U10707 ( .A(n8289), .B(n8313), .ZN(n9994) );
  NAND2_X1 U10708 ( .A1(n9895), .A2(n8290), .ZN(n8292) );
  NAND2_X1 U10709 ( .A1(n9674), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8291) );
  INV_X1 U10710 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8293) );
  NAND2_X1 U10711 ( .A1(n8294), .A2(n8293), .ZN(n8300) );
  NAND2_X1 U10712 ( .A1(n8353), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8299) );
  INV_X1 U10713 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n8296) );
  INV_X1 U10714 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9995) );
  OR2_X1 U10715 ( .A1(n8279), .A2(n9995), .ZN(n8297) );
  INV_X1 U10716 ( .A(n10847), .ZN(n13779) );
  NAND2_X1 U10717 ( .A1(n9525), .A2(n9524), .ZN(n10372) );
  NAND2_X1 U10718 ( .A1(n10847), .A2(n8301), .ZN(n8302) );
  INV_X1 U10719 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8303) );
  XNOR2_X1 U10720 ( .A(n8303), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n10861) );
  NAND2_X1 U10721 ( .A1(n8606), .A2(n10861), .ZN(n8311) );
  INV_X1 U10722 ( .A(n8304), .ZN(n8339) );
  NAND2_X1 U10723 ( .A1(n8339), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8310) );
  INV_X1 U10724 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n8306) );
  OR2_X1 U10725 ( .A1(n8305), .A2(n8306), .ZN(n8309) );
  INV_X1 U10726 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n8307) );
  OR2_X1 U10727 ( .A1(n8550), .A2(n8307), .ZN(n8308) );
  AND4_X2 U10728 ( .A1(n8311), .A2(n8310), .A3(n8309), .A4(n8308), .ZN(n10871)
         );
  NAND2_X1 U10729 ( .A1(n6725), .A2(n8313), .ZN(n8316) );
  NAND2_X1 U10730 ( .A1(n8316), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8315) );
  MUX2_X1 U10731 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8315), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n8317) );
  XNOR2_X1 U10732 ( .A(n10871), .B(n10876), .ZN(n10851) );
  NAND2_X1 U10733 ( .A1(n10850), .A2(n10851), .ZN(n8319) );
  NAND2_X1 U10734 ( .A1(n14670), .A2(n10871), .ZN(n8318) );
  NAND2_X1 U10735 ( .A1(n8319), .A2(n8318), .ZN(n10817) );
  NAND2_X1 U10736 ( .A1(n9899), .A2(n9656), .ZN(n8322) );
  NAND2_X1 U10737 ( .A1(n8331), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8320) );
  XNOR2_X1 U10738 ( .A(n8320), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10044) );
  AOI22_X1 U10739 ( .A1(n9674), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n9921), .B2(
        n10044), .ZN(n8321) );
  NAND2_X1 U10740 ( .A1(n8322), .A2(n8321), .ZN(n10901) );
  NAND2_X1 U10741 ( .A1(n9659), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U10742 ( .A1(n8295), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8326) );
  AOI21_X1 U10743 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8323) );
  NOR2_X1 U10744 ( .A1(n8323), .A2(n8337), .ZN(n10895) );
  NAND2_X1 U10745 ( .A1(n8606), .A2(n10895), .ZN(n8325) );
  NAND2_X1 U10746 ( .A1(n8339), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8324) );
  XNOR2_X1 U10747 ( .A(n10901), .B(n13777), .ZN(n10819) );
  INV_X1 U10748 ( .A(n10819), .ZN(n8328) );
  NAND2_X1 U10749 ( .A1(n10817), .A2(n8328), .ZN(n8330) );
  OR2_X1 U10750 ( .A1(n10901), .A2(n13777), .ZN(n8329) );
  NAND2_X1 U10751 ( .A1(n8330), .A2(n8329), .ZN(n14587) );
  NAND2_X1 U10752 ( .A1(n9918), .A2(n9656), .ZN(n8336) );
  INV_X1 U10753 ( .A(n8331), .ZN(n8333) );
  NAND2_X1 U10754 ( .A1(n8333), .A2(n8332), .ZN(n8346) );
  NAND2_X1 U10755 ( .A1(n8346), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8334) );
  XNOR2_X1 U10756 ( .A(n8334), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U10757 ( .A1(n9674), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n9921), .B2(
        n10252), .ZN(n8335) );
  NAND2_X1 U10758 ( .A1(n8336), .A2(n8335), .ZN(n13723) );
  NAND2_X1 U10759 ( .A1(n9659), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8343) );
  OAI21_X1 U10760 ( .B1(n8337), .B2(P1_REG3_REG_6__SCAN_IN), .A(n8351), .ZN(
        n14594) );
  INV_X1 U10761 ( .A(n14594), .ZN(n8338) );
  NAND2_X1 U10762 ( .A1(n8606), .A2(n8338), .ZN(n8341) );
  NAND2_X1 U10763 ( .A1(n8339), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8340) );
  NAND4_X1 U10764 ( .A1(n8343), .A2(n8342), .A3(n8341), .A4(n8340), .ZN(n13776) );
  XNOR2_X1 U10765 ( .A(n13723), .B(n13776), .ZN(n9688) );
  INV_X1 U10766 ( .A(n9688), .ZN(n14589) );
  NAND2_X1 U10767 ( .A1(n14587), .A2(n14589), .ZN(n8345) );
  OR2_X1 U10768 ( .A1(n13723), .A2(n13776), .ZN(n8344) );
  NAND2_X1 U10769 ( .A1(n8345), .A2(n8344), .ZN(n10750) );
  NAND2_X1 U10770 ( .A1(n9929), .A2(n9656), .ZN(n8349) );
  OAI21_X1 U10771 ( .B1(n8346), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8347) );
  XNOR2_X1 U10772 ( .A(n8347), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U10773 ( .A1(n9674), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n9921), .B2(
        n10432), .ZN(n8348) );
  NAND2_X1 U10774 ( .A1(n8349), .A2(n8348), .ZN(n11029) );
  NAND2_X1 U10775 ( .A1(n9659), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8357) );
  AND2_X1 U10776 ( .A1(n8351), .A2(n8350), .ZN(n8352) );
  NOR2_X1 U10777 ( .A1(n8366), .A2(n8352), .ZN(n11024) );
  NAND2_X1 U10778 ( .A1(n8606), .A2(n11024), .ZN(n8355) );
  NAND2_X1 U10779 ( .A1(n8339), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8354) );
  NAND4_X1 U10780 ( .A1(n8357), .A2(n8356), .A3(n8355), .A4(n8354), .ZN(n13775) );
  XNOR2_X1 U10781 ( .A(n11029), .B(n13775), .ZN(n10751) );
  INV_X1 U10782 ( .A(n10751), .ZN(n10753) );
  NAND2_X1 U10783 ( .A1(n10750), .A2(n10753), .ZN(n8359) );
  OR2_X1 U10784 ( .A1(n11029), .A2(n13775), .ZN(n8358) );
  NAND2_X1 U10785 ( .A1(n8359), .A2(n8358), .ZN(n10687) );
  NAND2_X1 U10786 ( .A1(n9953), .A2(n9656), .ZN(n8365) );
  NOR2_X1 U10787 ( .A1(n8486), .A2(n8241), .ZN(n8360) );
  MUX2_X1 U10788 ( .A(n8241), .B(n8360), .S(P1_IR_REG_8__SCAN_IN), .Z(n8363)
         );
  INV_X1 U10789 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8361) );
  NAND2_X1 U10790 ( .A1(n8486), .A2(n8361), .ZN(n8385) );
  INV_X1 U10791 ( .A(n8385), .ZN(n8362) );
  NOR2_X1 U10792 ( .A1(n8363), .A2(n8362), .ZN(n10734) );
  AOI22_X1 U10793 ( .A1(n9674), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9921), .B2(
        n10734), .ZN(n8364) );
  NAND2_X1 U10794 ( .A1(n8365), .A2(n8364), .ZN(n11257) );
  NAND2_X1 U10795 ( .A1(n9659), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8371) );
  OR2_X1 U10796 ( .A1(n8366), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8367) );
  AND2_X1 U10797 ( .A1(n8378), .A2(n8367), .ZN(n11269) );
  NAND2_X1 U10798 ( .A1(n8606), .A2(n11269), .ZN(n8369) );
  NAND2_X1 U10799 ( .A1(n8692), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8368) );
  NAND4_X1 U10800 ( .A1(n8371), .A2(n8370), .A3(n8369), .A4(n8368), .ZN(n13774) );
  INV_X1 U10801 ( .A(n13774), .ZN(n8667) );
  XNOR2_X1 U10802 ( .A(n11257), .B(n8667), .ZN(n10691) );
  NAND2_X1 U10803 ( .A1(n10687), .A2(n10691), .ZN(n8373) );
  OR2_X1 U10804 ( .A1(n11257), .A2(n13774), .ZN(n8372) );
  NAND2_X1 U10805 ( .A1(n9961), .A2(n9656), .ZN(n8376) );
  NAND2_X1 U10806 ( .A1(n8385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8374) );
  XNOR2_X1 U10807 ( .A(n8374), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U10808 ( .A1(n9674), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9921), .B2(
        n10987), .ZN(n8375) );
  NAND2_X1 U10809 ( .A1(n8376), .A2(n8375), .ZN(n14705) );
  NAND2_X1 U10810 ( .A1(n9659), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8383) );
  NAND2_X1 U10811 ( .A1(n8295), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U10812 ( .A1(n8378), .A2(n8377), .ZN(n8379) );
  AND2_X1 U10813 ( .A1(n8390), .A2(n8379), .ZN(n11338) );
  NAND2_X1 U10814 ( .A1(n8606), .A2(n11338), .ZN(n8381) );
  NAND2_X1 U10815 ( .A1(n8692), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8380) );
  NAND4_X1 U10816 ( .A1(n8383), .A2(n8382), .A3(n8381), .A4(n8380), .ZN(n13773) );
  XNOR2_X1 U10817 ( .A(n14705), .B(n13773), .ZN(n10932) );
  INV_X1 U10818 ( .A(n10932), .ZN(n10937) );
  OR2_X1 U10819 ( .A1(n14705), .A2(n13773), .ZN(n8384) );
  NAND2_X1 U10820 ( .A1(n9964), .A2(n9656), .ZN(n8388) );
  NAND2_X1 U10821 ( .A1(n8398), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8386) );
  XNOR2_X1 U10822 ( .A(n8386), .B(P1_IR_REG_10__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U10823 ( .A1(n9674), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n9921), 
        .B2(n11428), .ZN(n8387) );
  NAND2_X1 U10824 ( .A1(n8295), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10825 ( .A1(n9659), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10826 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  AND2_X1 U10827 ( .A1(n8403), .A2(n8391), .ZN(n11380) );
  NAND2_X1 U10828 ( .A1(n8606), .A2(n11380), .ZN(n8393) );
  NAND2_X1 U10829 ( .A1(n8339), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8392) );
  NAND4_X1 U10830 ( .A1(n8395), .A2(n8394), .A3(n8393), .A4(n8392), .ZN(n13772) );
  INV_X1 U10831 ( .A(n13772), .ZN(n8396) );
  OR2_X1 U10832 ( .A1(n11381), .A2(n8396), .ZN(n8671) );
  NAND2_X1 U10833 ( .A1(n11381), .A2(n8396), .ZN(n8397) );
  AND2_X1 U10834 ( .A1(n8671), .A2(n8397), .ZN(n9692) );
  NAND2_X1 U10835 ( .A1(n10035), .A2(n9656), .ZN(n8401) );
  NOR2_X1 U10836 ( .A1(n8398), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n8413) );
  OR2_X1 U10837 ( .A1(n8413), .A2(n8241), .ZN(n8399) );
  XNOR2_X1 U10838 ( .A(n8399), .B(P1_IR_REG_11__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U10839 ( .A1(n9674), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9921), 
        .B2(n11430), .ZN(n8400) );
  NAND2_X1 U10840 ( .A1(n8295), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8409) );
  AND2_X1 U10841 ( .A1(n8403), .A2(n8402), .ZN(n8404) );
  NOR2_X1 U10842 ( .A1(n8418), .A2(n8404), .ZN(n11642) );
  NAND2_X1 U10843 ( .A1(n8606), .A2(n11642), .ZN(n8408) );
  INV_X1 U10844 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8405) );
  OR2_X1 U10845 ( .A1(n8550), .A2(n8405), .ZN(n8407) );
  NAND2_X1 U10846 ( .A1(n8692), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8406) );
  NAND4_X1 U10847 ( .A1(n8409), .A2(n8408), .A3(n8407), .A4(n8406), .ZN(n13771) );
  XNOR2_X1 U10848 ( .A(n14453), .B(n13771), .ZN(n11214) );
  INV_X1 U10849 ( .A(n11214), .ZN(n11211) );
  NAND2_X1 U10850 ( .A1(n11210), .A2(n11211), .ZN(n8411) );
  OR2_X1 U10851 ( .A1(n14453), .A2(n13771), .ZN(n8410) );
  NAND2_X1 U10852 ( .A1(n8411), .A2(n8410), .ZN(n11348) );
  NAND2_X1 U10853 ( .A1(n10183), .A2(n9656), .ZN(n8416) );
  NAND2_X1 U10854 ( .A1(n8413), .A2(n8412), .ZN(n8414) );
  NAND2_X1 U10855 ( .A1(n8414), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8427) );
  XNOR2_X1 U10856 ( .A(n8427), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U10857 ( .A1(n9674), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9921), 
        .B2(n11862), .ZN(n8415) );
  NAND2_X1 U10858 ( .A1(n8692), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8422) );
  INV_X1 U10859 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8417) );
  OR2_X1 U10860 ( .A1(n8550), .A2(n8417), .ZN(n8421) );
  OR2_X1 U10861 ( .A1(n8418), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n8419) );
  AND2_X1 U10862 ( .A1(n8419), .A2(n8447), .ZN(n11687) );
  NAND2_X1 U10863 ( .A1(n8606), .A2(n11687), .ZN(n8420) );
  NAND4_X1 U10864 ( .A1(n8423), .A2(n8422), .A3(n8421), .A4(n8420), .ZN(n13770) );
  INV_X1 U10865 ( .A(n13770), .ZN(n8674) );
  XNOR2_X1 U10866 ( .A(n11678), .B(n8674), .ZN(n11349) );
  NAND2_X1 U10867 ( .A1(n11348), .A2(n11349), .ZN(n8425) );
  OR2_X1 U10868 ( .A1(n11678), .A2(n13770), .ZN(n8424) );
  NAND2_X1 U10869 ( .A1(n8425), .A2(n8424), .ZN(n11469) );
  NAND2_X1 U10870 ( .A1(n10260), .A2(n9656), .ZN(n8430) );
  INV_X1 U10871 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U10872 ( .A1(n8427), .A2(n8426), .ZN(n8428) );
  NAND2_X1 U10873 ( .A1(n8428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8440) );
  XNOR2_X1 U10874 ( .A(n8440), .B(P1_IR_REG_13__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U10875 ( .A1(n9674), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n11865), 
        .B2(n9921), .ZN(n8429) );
  NAND2_X1 U10876 ( .A1(n8295), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U10877 ( .A1(n8692), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8433) );
  XNOR2_X1 U10878 ( .A(n8447), .B(P1_REG3_REG_13__SCAN_IN), .ZN(n11477) );
  NAND2_X1 U10879 ( .A1(n8606), .A2(n11477), .ZN(n8432) );
  NAND2_X1 U10880 ( .A1(n9659), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8431) );
  NAND4_X1 U10881 ( .A1(n8434), .A2(n8433), .A3(n8432), .A4(n8431), .ZN(n14388) );
  INV_X1 U10882 ( .A(n14388), .ZN(n8435) );
  OR2_X1 U10883 ( .A1(n11733), .A2(n8435), .ZN(n8676) );
  NAND2_X1 U10884 ( .A1(n11733), .A2(n8435), .ZN(n8436) );
  NAND2_X1 U10885 ( .A1(n8676), .A2(n8436), .ZN(n9694) );
  NAND2_X1 U10886 ( .A1(n11469), .A2(n9694), .ZN(n8438) );
  OR2_X1 U10887 ( .A1(n11733), .A2(n14388), .ZN(n8437) );
  NAND2_X1 U10888 ( .A1(n10423), .A2(n9656), .ZN(n8444) );
  INV_X1 U10889 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8439) );
  NAND2_X1 U10890 ( .A1(n8440), .A2(n8439), .ZN(n8441) );
  NAND2_X1 U10891 ( .A1(n8441), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8442) );
  XNOR2_X1 U10892 ( .A(n8442), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14525) );
  AOI22_X1 U10893 ( .A1(n14525), .A2(n9921), .B1(n9674), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8443) );
  INV_X1 U10894 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8446) );
  INV_X1 U10895 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8445) );
  OAI21_X1 U10896 ( .B1(n8447), .B2(n8446), .A(n8445), .ZN(n8448) );
  NAND2_X1 U10897 ( .A1(n8448), .A2(n8461), .ZN(n14400) );
  INV_X1 U10898 ( .A(n14400), .ZN(n14408) );
  NAND2_X1 U10899 ( .A1(n8606), .A2(n14408), .ZN(n8453) );
  NAND2_X1 U10900 ( .A1(n8692), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n8452) );
  INV_X1 U10901 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8449) );
  OR2_X1 U10902 ( .A1(n8305), .A2(n8449), .ZN(n8451) );
  INV_X1 U10903 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11858) );
  OR2_X1 U10904 ( .A1(n8550), .A2(n11858), .ZN(n8450) );
  NAND2_X1 U10905 ( .A1(n14414), .A2(n13495), .ZN(n9574) );
  INV_X1 U10906 ( .A(n13495), .ZN(n13769) );
  NAND2_X1 U10907 ( .A1(n14414), .A2(n13769), .ZN(n8454) );
  NAND2_X1 U10908 ( .A1(n10557), .A2(n9656), .ZN(n8460) );
  INV_X1 U10909 ( .A(n8484), .ZN(n8455) );
  NAND2_X1 U10910 ( .A1(n8486), .A2(n8455), .ZN(n8624) );
  NAND2_X1 U10911 ( .A1(n8624), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8457) );
  XNOR2_X1 U10912 ( .A(n8457), .B(n8456), .ZN(n13840) );
  INV_X1 U10913 ( .A(n13840), .ZN(n8458) );
  AOI22_X1 U10914 ( .A1(n9674), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9921), 
        .B2(n8458), .ZN(n8459) );
  AND2_X1 U10915 ( .A1(n8461), .A2(n15104), .ZN(n8462) );
  NOR2_X1 U10916 ( .A1(n8475), .A2(n8462), .ZN(n13745) );
  NAND2_X1 U10917 ( .A1(n13745), .A2(n8606), .ZN(n8466) );
  NAND2_X1 U10918 ( .A1(n9659), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8465) );
  NAND2_X1 U10919 ( .A1(n8692), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U10920 ( .A1(n14439), .A2(n14386), .ZN(n9581) );
  NAND2_X1 U10921 ( .A1(n9582), .A2(n9581), .ZN(n9697) );
  INV_X1 U10922 ( .A(n14386), .ZN(n13768) );
  OR2_X1 U10923 ( .A1(n14439), .A2(n13768), .ZN(n8467) );
  NAND2_X1 U10924 ( .A1(n10440), .A2(n9656), .ZN(n8474) );
  OR2_X1 U10925 ( .A1(n8624), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U10926 ( .A1(n8469), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8468) );
  MUX2_X1 U10927 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8468), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n8472) );
  INV_X1 U10928 ( .A(n8469), .ZN(n8471) );
  NAND2_X1 U10929 ( .A1(n8471), .A2(n8470), .ZN(n8487) );
  NAND2_X1 U10930 ( .A1(n8472), .A2(n8487), .ZN(n14549) );
  INV_X1 U10931 ( .A(n14549), .ZN(n13844) );
  AOI22_X1 U10932 ( .A1(n9674), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9921), 
        .B2(n13844), .ZN(n8473) );
  NOR2_X1 U10933 ( .A1(n8475), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8476) );
  OR2_X1 U10934 ( .A1(n8492), .A2(n8476), .ZN(n13665) );
  NAND2_X1 U10935 ( .A1(n9659), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10936 ( .A1(n8295), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8477) );
  AND2_X1 U10937 ( .A1(n8478), .A2(n8477), .ZN(n8480) );
  NAND2_X1 U10938 ( .A1(n8692), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8479) );
  OAI211_X1 U10939 ( .C1(n13665), .C2(n8530), .A(n8480), .B(n8479), .ZN(n13767) );
  XNOR2_X1 U10940 ( .A(n14430), .B(n13767), .ZN(n9695) );
  NAND2_X1 U10941 ( .A1(n11776), .A2(n7275), .ZN(n8482) );
  OR2_X1 U10942 ( .A1(n14430), .A2(n13767), .ZN(n8481) );
  NAND2_X1 U10943 ( .A1(n10556), .A2(n9656), .ZN(n8491) );
  NOR2_X1 U10944 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  NAND2_X1 U10945 ( .A1(n8486), .A2(n8485), .ZN(n8506) );
  NAND2_X1 U10946 ( .A1(n8487), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8488) );
  MUX2_X1 U10947 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8488), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n8489) );
  AND2_X1 U10948 ( .A1(n8506), .A2(n8489), .ZN(n13849) );
  AOI22_X1 U10949 ( .A1(n9674), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9921), 
        .B2(n13849), .ZN(n8490) );
  OR2_X1 U10950 ( .A1(n8492), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U10951 ( .A1(n8515), .A2(n8493), .ZN(n13670) );
  NAND2_X1 U10952 ( .A1(n8692), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8494) );
  OAI211_X1 U10953 ( .C1(n13670), .C2(n8530), .A(n8495), .B(n8494), .ZN(n13766) );
  NOR2_X1 U10954 ( .A1(n14423), .A2(n13766), .ZN(n9682) );
  NAND2_X1 U10955 ( .A1(n14423), .A2(n13766), .ZN(n9683) );
  OR2_X1 U10956 ( .A1(n10778), .A2(n8312), .ZN(n8498) );
  NAND2_X1 U10957 ( .A1(n8506), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8496) );
  XNOR2_X1 U10958 ( .A(n8496), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14581) );
  AOI22_X1 U10959 ( .A1(n9674), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9921), 
        .B2(n14581), .ZN(n8497) );
  XNOR2_X1 U10960 ( .A(n8515), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n14041) );
  NAND2_X1 U10961 ( .A1(n14041), .A2(n8606), .ZN(n8504) );
  INV_X1 U10962 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U10963 ( .A1(n8692), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8500) );
  OAI211_X1 U10964 ( .C1(n8550), .C2(n8501), .A(n8500), .B(n8499), .ZN(n8502)
         );
  INV_X1 U10965 ( .A(n8502), .ZN(n8503) );
  NAND2_X1 U10966 ( .A1(n8504), .A2(n8503), .ZN(n13765) );
  INV_X1 U10967 ( .A(n13765), .ZN(n13530) );
  NOR2_X1 U10968 ( .A1(n14044), .A2(n13530), .ZN(n8505) );
  NAND2_X1 U10969 ( .A1(n11085), .A2(n9656), .ZN(n8512) );
  AOI22_X1 U10970 ( .A1(n9674), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14023), 
        .B2(n9921), .ZN(n8511) );
  INV_X1 U10971 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8514) );
  INV_X1 U10972 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8513) );
  OAI21_X1 U10973 ( .B1(n8515), .B2(n8514), .A(n8513), .ZN(n8516) );
  NAND2_X1 U10974 ( .A1(n8516), .A2(n8524), .ZN(n13620) );
  OR2_X1 U10975 ( .A1(n13620), .A2(n8530), .ZN(n8519) );
  AOI22_X1 U10976 ( .A1(n9659), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n8295), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U10977 ( .A1(n8692), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8517) );
  AND3_X1 U10978 ( .A1(n8519), .A2(n8518), .A3(n8517), .ZN(n13711) );
  NAND2_X1 U10979 ( .A1(n14027), .A2(n13711), .ZN(n9600) );
  NAND2_X1 U10980 ( .A1(n14020), .A2(n14019), .ZN(n8521) );
  INV_X1 U10981 ( .A(n13711), .ZN(n13764) );
  OR2_X1 U10982 ( .A1(n14027), .A2(n13764), .ZN(n8520) );
  NAND2_X1 U10983 ( .A1(n11416), .A2(n9656), .ZN(n8523) );
  NAND2_X1 U10984 ( .A1(n9674), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8522) );
  AND2_X1 U10985 ( .A1(n8524), .A2(n13694), .ZN(n8525) );
  OR2_X1 U10986 ( .A1(n8525), .A2(n8534), .ZN(n14006) );
  INV_X1 U10987 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n14119) );
  NAND2_X1 U10988 ( .A1(n8295), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8527) );
  NAND2_X1 U10989 ( .A1(n9659), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8526) );
  OAI211_X1 U10990 ( .C1(n8304), .C2(n14119), .A(n8527), .B(n8526), .ZN(n8528)
         );
  INV_X1 U10991 ( .A(n8528), .ZN(n8529) );
  XNOR2_X1 U10992 ( .A(n14113), .B(n13763), .ZN(n13996) );
  NAND2_X1 U10993 ( .A1(n14113), .A2(n13763), .ZN(n8531) );
  NAND2_X1 U10994 ( .A1(n9674), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8532) );
  OR2_X1 U10995 ( .A1(n8534), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8535) );
  AND2_X1 U10996 ( .A1(n8535), .A2(n8548), .ZN(n13989) );
  NAND2_X1 U10997 ( .A1(n13989), .A2(n8606), .ZN(n8541) );
  INV_X1 U10998 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U10999 ( .A1(n8692), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U11000 ( .A1(n9659), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8536) );
  OAI211_X1 U11001 ( .C1(n8305), .C2(n8538), .A(n8537), .B(n8536), .ZN(n8539)
         );
  INV_X1 U11002 ( .A(n8539), .ZN(n8540) );
  NAND2_X1 U11003 ( .A1(n8541), .A2(n8540), .ZN(n13762) );
  INV_X1 U11004 ( .A(n13762), .ZN(n8542) );
  NAND2_X1 U11005 ( .A1(n13992), .A2(n8542), .ZN(n8544) );
  NAND2_X1 U11006 ( .A1(n14108), .A2(n13762), .ZN(n8543) );
  NAND2_X1 U11007 ( .A1(n8544), .A2(n8543), .ZN(n13985) );
  NAND2_X1 U11008 ( .A1(n8129), .A2(n9925), .ZN(n8545) );
  XNOR2_X1 U11009 ( .A(n8545), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14174) );
  NAND2_X1 U11010 ( .A1(n14174), .A2(n8546), .ZN(n14101) );
  INV_X1 U11011 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13703) );
  AOI21_X1 U11012 ( .B1(n13703), .B2(n8548), .A(n8547), .ZN(n13975) );
  NAND2_X1 U11013 ( .A1(n8606), .A2(n13975), .ZN(n8555) );
  NAND2_X1 U11014 ( .A1(n8692), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8554) );
  INV_X1 U11015 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8549) );
  OR2_X1 U11016 ( .A1(n8550), .A2(n8549), .ZN(n8553) );
  INV_X1 U11017 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8551) );
  OR2_X1 U11018 ( .A1(n8305), .A2(n8551), .ZN(n8552) );
  XNOR2_X1 U11019 ( .A(n14101), .B(n13642), .ZN(n13970) );
  INV_X1 U11020 ( .A(n13970), .ZN(n13972) );
  NAND2_X1 U11021 ( .A1(n13973), .A2(n13972), .ZN(n8557) );
  NAND2_X1 U11022 ( .A1(n14101), .A2(n13642), .ZN(n8556) );
  NAND2_X1 U11023 ( .A1(n8557), .A2(n8556), .ZN(n13966) );
  NAND2_X1 U11024 ( .A1(n11816), .A2(n9656), .ZN(n8559) );
  NAND2_X1 U11025 ( .A1(n9674), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U11026 ( .A1(n9659), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8565) );
  INV_X1 U11027 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13612) );
  INV_X1 U11028 ( .A(n8569), .ZN(n8560) );
  AOI21_X1 U11029 ( .B1(n13612), .B2(n8561), .A(n8560), .ZN(n13961) );
  NAND2_X1 U11030 ( .A1(n8606), .A2(n13961), .ZN(n8563) );
  NAND2_X1 U11031 ( .A1(n8692), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8562) );
  NAND4_X1 U11032 ( .A1(n8565), .A2(n8564), .A3(n8563), .A4(n8562), .ZN(n13760) );
  XNOR2_X1 U11033 ( .A(n14093), .B(n13760), .ZN(n13967) );
  OR2_X2 U11034 ( .A1(n13966), .A2(n13967), .ZN(n14095) );
  NAND2_X1 U11035 ( .A1(n14093), .A2(n13760), .ZN(n8566) );
  NAND2_X1 U11036 ( .A1(n11844), .A2(n9656), .ZN(n8568) );
  NAND2_X1 U11037 ( .A1(n9674), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8567) );
  NAND2_X1 U11038 ( .A1(n9659), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11039 ( .A1(n8295), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8572) );
  AOI21_X1 U11040 ( .B1(n15248), .B2(n8569), .A(n8576), .ZN(n13948) );
  NAND2_X1 U11041 ( .A1(n8606), .A2(n13948), .ZN(n8571) );
  NAND2_X1 U11042 ( .A1(n8692), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8570) );
  NAND4_X1 U11043 ( .A1(n8573), .A2(n8572), .A3(n8571), .A4(n8570), .ZN(n13759) );
  INV_X1 U11044 ( .A(n13759), .ZN(n8684) );
  XNOR2_X1 U11045 ( .A(n14087), .B(n8684), .ZN(n13942) );
  NAND2_X1 U11046 ( .A1(n13460), .A2(n9656), .ZN(n8575) );
  NAND2_X1 U11047 ( .A1(n9674), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8574) );
  NAND2_X1 U11048 ( .A1(n9659), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8582) );
  INV_X1 U11049 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13656) );
  INV_X1 U11050 ( .A(n8576), .ZN(n8578) );
  AOI21_X1 U11051 ( .B1(n13656), .B2(n8578), .A(n8577), .ZN(n13931) );
  NAND2_X1 U11052 ( .A1(n8606), .A2(n13931), .ZN(n8580) );
  NAND2_X1 U11053 ( .A1(n8692), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8579) );
  NAND4_X1 U11054 ( .A1(n8582), .A2(n8581), .A3(n8580), .A4(n8579), .ZN(n13758) );
  INV_X1 U11055 ( .A(n13758), .ZN(n8583) );
  XNOR2_X1 U11056 ( .A(n14082), .B(n8583), .ZN(n13927) );
  INV_X1 U11057 ( .A(n14082), .ZN(n13660) );
  NAND2_X1 U11058 ( .A1(n13456), .A2(n9656), .ZN(n8585) );
  NAND2_X1 U11059 ( .A1(n9674), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U11060 ( .A1(n8295), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U11061 ( .A1(n9659), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8590) );
  INV_X1 U11062 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13735) );
  INV_X1 U11063 ( .A(n8586), .ZN(n8595) );
  AOI21_X1 U11064 ( .B1(n13735), .B2(n8587), .A(n8595), .ZN(n13916) );
  NAND2_X1 U11065 ( .A1(n8606), .A2(n13916), .ZN(n8589) );
  NAND2_X1 U11066 ( .A1(n8692), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8588) );
  NAND4_X1 U11067 ( .A1(n8591), .A2(n8590), .A3(n8589), .A4(n8588), .ZN(n13757) );
  NAND2_X1 U11068 ( .A1(n13915), .A2(n13599), .ZN(n13893) );
  OR2_X1 U11069 ( .A1(n13915), .A2(n13599), .ZN(n8592) );
  NAND2_X1 U11070 ( .A1(n13893), .A2(n8592), .ZN(n13912) );
  XNOR2_X1 U11071 ( .A(n14066), .B(n13756), .ZN(n13907) );
  NAND2_X1 U11072 ( .A1(n14156), .A2(n9656), .ZN(n8594) );
  NAND2_X1 U11073 ( .A1(n9674), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8593) );
  NAND2_X1 U11074 ( .A1(n9659), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8603) );
  NAND2_X1 U11075 ( .A1(n8295), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U11076 ( .A1(n8596), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8695) );
  INV_X1 U11077 ( .A(n8596), .ZN(n8598) );
  INV_X1 U11078 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11079 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  NAND2_X1 U11080 ( .A1(n8606), .A2(n13633), .ZN(n8601) );
  NAND2_X1 U11081 ( .A1(n8692), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8600) );
  NAND4_X1 U11082 ( .A1(n8603), .A2(n8602), .A3(n8601), .A4(n8600), .ZN(n13755) );
  OR2_X1 U11083 ( .A1(n14061), .A2(n13628), .ZN(n8604) );
  AOI22_X1 U11084 ( .A1(n9659), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8295), .B2(
        P1_REG0_REG_29__SCAN_IN), .ZN(n8608) );
  INV_X1 U11085 ( .A(n8695), .ZN(n8605) );
  AOI22_X1 U11086 ( .A1(n8692), .A2(P1_REG1_REG_29__SCAN_IN), .B1(n8606), .B2(
        n8605), .ZN(n8607) );
  AND2_X1 U11087 ( .A1(n8608), .A2(n8607), .ZN(n13635) );
  NAND2_X1 U11088 ( .A1(n8610), .A2(n8609), .ZN(n8612) );
  INV_X1 U11089 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15205) );
  MUX2_X1 U11090 ( .A(n15205), .B(n13448), .S(n9926), .Z(n9650) );
  NAND2_X1 U11091 ( .A1(n13447), .A2(n9656), .ZN(n8614) );
  NAND2_X1 U11092 ( .A1(n9674), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8613) );
  XNOR2_X2 U11093 ( .A(n8620), .B(P1_IR_REG_21__SCAN_IN), .ZN(n10011) );
  NAND2_X1 U11094 ( .A1(n9504), .A2(n10011), .ZN(n10014) );
  MUX2_X1 U11095 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8621), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n8623) );
  AND2_X1 U11096 ( .A1(n11454), .A2(n13858), .ZN(n10012) );
  INV_X1 U11097 ( .A(n8624), .ZN(n8626) );
  NAND2_X1 U11098 ( .A1(n8626), .A2(n8625), .ZN(n8630) );
  OR2_X2 U11099 ( .A1(n8630), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n8632) );
  NAND2_X1 U11100 ( .A1(n8632), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11101 ( .A1(n8630), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8631) );
  MUX2_X1 U11102 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8631), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8633) );
  AND2_X2 U11103 ( .A1(n8633), .A2(n8632), .ZN(n11847) );
  OAI211_X1 U11104 ( .C1(n10014), .C2(n10012), .A(n10023), .B(n9922), .ZN(
        n10472) );
  INV_X4 U11105 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OR2_X1 U11106 ( .A1(n10472), .A2(P1_U3086), .ZN(n10193) );
  NOR2_X1 U11107 ( .A1(n14168), .A2(n8637), .ZN(n8638) );
  MUX2_X1 U11108 ( .A(n8638), .B(n8637), .S(n11847), .Z(n8639) );
  INV_X1 U11109 ( .A(n8639), .ZN(n8640) );
  NAND2_X1 U11110 ( .A1(n8640), .A2(n14162), .ZN(n10190) );
  NOR4_X1 U11111 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n8649) );
  NOR4_X1 U11112 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n8648) );
  NOR4_X1 U11113 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n8644) );
  NOR4_X1 U11114 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n8643) );
  NOR4_X1 U11115 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n8642) );
  NOR4_X1 U11116 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n8641) );
  NAND4_X1 U11117 ( .A1(n8644), .A2(n8643), .A3(n8642), .A4(n8641), .ZN(n8645)
         );
  NOR4_X1 U11118 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n8646), .A4(n8645), .ZN(n8647) );
  NAND3_X1 U11119 ( .A1(n8649), .A2(n8648), .A3(n8647), .ZN(n10188) );
  INV_X1 U11120 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10195) );
  NOR2_X1 U11121 ( .A1(n10188), .A2(n10195), .ZN(n8650) );
  OR2_X1 U11122 ( .A1(n10190), .A2(n8650), .ZN(n8651) );
  NAND2_X1 U11123 ( .A1(n8651), .A2(n9936), .ZN(n10004) );
  NOR2_X1 U11124 ( .A1(n10193), .A2(n10004), .ZN(n8652) );
  INV_X1 U11125 ( .A(n10190), .ZN(n10196) );
  INV_X1 U11126 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9939) );
  INV_X1 U11127 ( .A(n11587), .ZN(n10199) );
  NAND2_X1 U11128 ( .A1(n8652), .A2(n10199), .ZN(n8696) );
  OR2_X4 U11129 ( .A1(n10201), .A2(n10011), .ZN(n14675) );
  AND2_X1 U11130 ( .A1(n9937), .A2(n10023), .ZN(n10006) );
  NAND2_X2 U11131 ( .A1(n9505), .A2(n10019), .ZN(n13625) );
  OR2_X1 U11132 ( .A1(n9505), .A2(n10019), .ZN(n8653) );
  NAND2_X1 U11133 ( .A1(n13625), .A2(n8653), .ZN(n10200) );
  NAND2_X1 U11134 ( .A1(n9513), .A2(n8654), .ZN(n9512) );
  NAND2_X1 U11135 ( .A1(n10164), .A2(n10264), .ZN(n8655) );
  INV_X1 U11136 ( .A(n10372), .ZN(n10375) );
  NAND2_X1 U11137 ( .A1(n10374), .A2(n10375), .ZN(n10373) );
  NAND2_X1 U11138 ( .A1(n10373), .A2(n9524), .ZN(n10845) );
  INV_X1 U11139 ( .A(n10851), .ZN(n8656) );
  NAND2_X1 U11140 ( .A1(n10845), .A2(n8656), .ZN(n8658) );
  NAND2_X1 U11141 ( .A1(n10876), .A2(n10871), .ZN(n8657) );
  NAND2_X1 U11142 ( .A1(n8658), .A2(n8657), .ZN(n10820) );
  NAND2_X1 U11143 ( .A1(n10820), .A2(n10819), .ZN(n8661) );
  INV_X1 U11144 ( .A(n13777), .ZN(n8659) );
  NAND2_X1 U11145 ( .A1(n10901), .A2(n8659), .ZN(n8660) );
  NAND2_X1 U11146 ( .A1(n8661), .A2(n8660), .ZN(n14590) );
  NAND2_X1 U11147 ( .A1(n14590), .A2(n9688), .ZN(n8664) );
  INV_X1 U11148 ( .A(n13776), .ZN(n8662) );
  NAND2_X1 U11149 ( .A1(n13723), .A2(n8662), .ZN(n8663) );
  NAND2_X1 U11150 ( .A1(n8664), .A2(n8663), .ZN(n10754) );
  INV_X1 U11151 ( .A(n13775), .ZN(n8665) );
  NAND2_X1 U11152 ( .A1(n11029), .A2(n8665), .ZN(n8666) );
  OR2_X1 U11153 ( .A1(n11257), .A2(n8667), .ZN(n8668) );
  INV_X1 U11154 ( .A(n13773), .ZN(n8669) );
  NAND2_X1 U11155 ( .A1(n14705), .A2(n8669), .ZN(n8670) );
  INV_X1 U11156 ( .A(n13771), .ZN(n8672) );
  OR2_X1 U11157 ( .A1(n14453), .A2(n8672), .ZN(n8673) );
  INV_X1 U11158 ( .A(n11349), .ZN(n11343) );
  OR2_X1 U11159 ( .A1(n11678), .A2(n8674), .ZN(n8675) );
  INV_X1 U11160 ( .A(n9694), .ZN(n11472) );
  INV_X1 U11161 ( .A(n13767), .ZN(n11823) );
  NAND2_X1 U11162 ( .A1(n14430), .A2(n11823), .ZN(n8677) );
  NAND2_X1 U11163 ( .A1(n11766), .A2(n8677), .ZN(n11822) );
  INV_X1 U11164 ( .A(n14423), .ZN(n8678) );
  XNOR2_X1 U11165 ( .A(n14130), .B(n13765), .ZN(n14034) );
  NAND2_X1 U11166 ( .A1(n14044), .A2(n13765), .ZN(n9595) );
  INV_X1 U11167 ( .A(n13996), .ZN(n14000) );
  INV_X1 U11168 ( .A(n13763), .ZN(n13643) );
  OR2_X1 U11169 ( .A1(n14113), .A2(n13643), .ZN(n8680) );
  INV_X1 U11170 ( .A(n13642), .ZN(n13761) );
  NAND2_X1 U11171 ( .A1(n13967), .A2(n13957), .ZN(n13956) );
  INV_X1 U11172 ( .A(n13760), .ZN(n8681) );
  NAND2_X1 U11173 ( .A1(n14093), .A2(n8681), .ZN(n8682) );
  OR2_X1 U11174 ( .A1(n14087), .A2(n8684), .ZN(n8685) );
  INV_X1 U11175 ( .A(n13912), .ZN(n13923) );
  INV_X1 U11176 ( .A(n13893), .ZN(n8686) );
  OAI21_X1 U11177 ( .B1(n13904), .B2(n13756), .A(n13895), .ZN(n13878) );
  NAND2_X1 U11178 ( .A1(n13878), .A2(n13879), .ZN(n13877) );
  INV_X1 U11179 ( .A(n9703), .ZN(n8688) );
  NAND2_X1 U11180 ( .A1(n9504), .A2(n14023), .ZN(n8690) );
  INV_X1 U11181 ( .A(n11454), .ZN(n9507) );
  NAND2_X1 U11182 ( .A1(n10011), .A2(n9507), .ZN(n8689) );
  INV_X1 U11183 ( .A(n11733), .ZN(n11591) );
  NAND2_X1 U11184 ( .A1(n14652), .A2(n14628), .ZN(n14627) );
  NAND2_X1 U11185 ( .A1(n14616), .A2(n8301), .ZN(n10853) );
  OR2_X1 U11186 ( .A1(n10853), .A2(n10876), .ZN(n10854) );
  INV_X1 U11187 ( .A(n13723), .ZN(n14682) );
  AND2_X1 U11188 ( .A1(n14600), .A2(n14682), .ZN(n14598) );
  INV_X1 U11189 ( .A(n11029), .ZN(n14692) );
  NAND2_X1 U11190 ( .A1(n14598), .A2(n14692), .ZN(n10689) );
  OR2_X1 U11191 ( .A1(n10689), .A2(n11257), .ZN(n10939) );
  INV_X1 U11192 ( .A(n11381), .ZN(n14718) );
  OR2_X1 U11193 ( .A1(n14414), .A2(n14415), .ZN(n14416) );
  OR2_X1 U11194 ( .A1(n11772), .A2(n14430), .ZN(n11827) );
  NOR2_X2 U11195 ( .A1(n14108), .A2(n14009), .ZN(n13988) );
  NOR2_X2 U11196 ( .A1(n13915), .A2(n13929), .ZN(n13914) );
  AOI21_X1 U11197 ( .B1(n9645), .B2(n6522), .A(n6477), .ZN(n14056) );
  NOR2_X1 U11198 ( .A1(n14011), .A2(n14675), .ZN(n13920) );
  INV_X1 U11199 ( .A(n10011), .ZN(n11558) );
  NAND2_X1 U11200 ( .A1(n11558), .A2(n9507), .ZN(n9704) );
  OR2_X1 U11201 ( .A1(n9704), .A2(n9504), .ZN(n10008) );
  INV_X1 U11202 ( .A(n14159), .ZN(n13783) );
  NOR2_X1 U11203 ( .A1(n6459), .A2(n8637), .ZN(n8691) );
  NOR2_X1 U11204 ( .A1(n14385), .A2(n8691), .ZN(n13865) );
  INV_X1 U11205 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n15130) );
  NAND2_X1 U11206 ( .A1(n9659), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U11207 ( .A1(n8692), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8693) );
  OAI211_X1 U11208 ( .C1(n8305), .C2(n15130), .A(n8694), .B(n8693), .ZN(n13753) );
  NAND2_X1 U11209 ( .A1(n13865), .A2(n13753), .ZN(n14053) );
  OAI22_X1 U11210 ( .A1(n8696), .A2(n14053), .B1(n8695), .B2(n14612), .ZN(
        n8697) );
  AOI21_X1 U11211 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n14648), .A(n8697), .ZN(
        n8698) );
  OAI21_X1 U11212 ( .B1(n14054), .B2(n14640), .A(n8698), .ZN(n8699) );
  AOI21_X1 U11213 ( .B1(n14056), .B2(n13920), .A(n8699), .ZN(n8700) );
  INV_X1 U11214 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9942) );
  NAND2_X1 U11215 ( .A1(n9942), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8702) );
  INV_X1 U11216 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9901) );
  NAND2_X1 U11217 ( .A1(n9901), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8703) );
  INV_X1 U11218 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9896) );
  AND2_X1 U11219 ( .A1(n9896), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U11220 ( .A1(n9934), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U11221 ( .A1(n8853), .A2(n8854), .ZN(n8708) );
  INV_X1 U11222 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n8706) );
  NAND2_X1 U11223 ( .A1(n8706), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8707) );
  NAND2_X1 U11224 ( .A1(n9932), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U11225 ( .A1(n9920), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U11226 ( .A1(n9945), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U11227 ( .A1(n8712), .A2(n8710), .ZN(n8885) );
  INV_X1 U11228 ( .A(n8885), .ZN(n8711) );
  NAND2_X1 U11229 ( .A1(n8888), .A2(n8712), .ZN(n8902) );
  XNOR2_X1 U11230 ( .A(n8713), .B(P1_DATAO_REG_7__SCAN_IN), .ZN(n8901) );
  OAI22_X2 U11231 ( .A1(n8902), .A2(n8901), .B1(P2_DATAO_REG_7__SCAN_IN), .B2(
        n9941), .ZN(n8918) );
  AND2_X1 U11232 ( .A1(n9955), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11233 ( .A1(n9954), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8715) );
  AND2_X1 U11234 ( .A1(n9963), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8716) );
  INV_X1 U11235 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U11236 ( .A1(n9965), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8717) );
  NAND2_X1 U11237 ( .A1(n8718), .A2(n8717), .ZN(n8961) );
  XNOR2_X1 U11238 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8969) );
  NAND2_X1 U11239 ( .A1(n8970), .A2(n8969), .ZN(n8721) );
  NAND2_X1 U11240 ( .A1(n10186), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U11241 ( .A1(n8722), .A2(n10274), .ZN(n8723) );
  INV_X1 U11242 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U11243 ( .A1(n8724), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8725) );
  XNOR2_X1 U11244 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n9007) );
  NAND2_X1 U11245 ( .A1(n9009), .A2(n9007), .ZN(n8727) );
  NAND2_X1 U11246 ( .A1(n10589), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8726) );
  NAND2_X1 U11247 ( .A1(n8727), .A2(n8726), .ZN(n9024) );
  XNOR2_X1 U11248 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n9022) );
  NAND2_X1 U11249 ( .A1(n9024), .A2(n9022), .ZN(n8729) );
  NAND2_X1 U11250 ( .A1(n10441), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U11251 ( .A1(n15219), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8730) );
  XNOR2_X1 U11252 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .ZN(n9054) );
  AOI22_X1 U11253 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n11086), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n11087), .ZN(n9071) );
  AOI22_X1 U11254 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n11453), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n15251), .ZN(n9086) );
  INV_X1 U11255 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11514) );
  AOI22_X1 U11256 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(
        P1_DATAO_REG_21__SCAN_IN), .B1(n11514), .B2(n11556), .ZN(n9098) );
  INV_X1 U11257 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11992) );
  INV_X1 U11258 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8736) );
  AOI22_X1 U11259 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n11992), .B2(n8736), .ZN(n9107) );
  AOI22_X1 U11260 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n11814), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n11819), .ZN(n9118) );
  NAND2_X1 U11261 ( .A1(n9117), .A2(n9118), .ZN(n8740) );
  INV_X1 U11262 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13463) );
  INV_X1 U11263 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14169) );
  AOI22_X1 U11264 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n13463), .B2(n14169), .ZN(n9141) );
  AOI22_X1 U11265 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n13457), .B2(n14164), .ZN(n9154) );
  AOI22_X1 U11266 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13455), .B2(n14160), .ZN(n8779) );
  AOI22_X1 U11267 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(
        P1_DATAO_REG_28__SCAN_IN), .B1(n13453), .B2(n14157), .ZN(n9283) );
  INV_X1 U11268 ( .A(n9283), .ZN(n8744) );
  XNOR2_X1 U11269 ( .A(n9284), .B(n8744), .ZN(n11873) );
  INV_X1 U11270 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8745) );
  AND2_X2 U11271 ( .A1(n10404), .A2(n8745), .ZN(n8840) );
  NOR2_X1 U11272 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n8747) );
  NOR2_X1 U11273 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8746) );
  AND2_X1 U11274 ( .A1(n8747), .A2(n8746), .ZN(n8750) );
  NOR2_X1 U11275 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n8749) );
  NOR3_X2 U11276 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .A3(
        P3_IR_REG_4__SCAN_IN), .ZN(n8748) );
  INV_X1 U11277 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8751) );
  NOR2_X1 U11278 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n8753) );
  NAND4_X1 U11279 ( .A1(n8753), .A2(n8752), .A3(n9057), .A4(n9010), .ZN(n9168)
         );
  NAND4_X1 U11280 ( .A1(n8755), .A2(n9170), .A3(n8754), .A4(n9256), .ZN(n8756)
         );
  INV_X1 U11281 ( .A(n8768), .ZN(n8770) );
  NAND2_X1 U11282 ( .A1(n8759), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8760) );
  MUX2_X1 U11283 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8760), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n8761) );
  NAND2_X1 U11284 ( .A1(n11873), .A2(n8819), .ZN(n8764) );
  NOR2_X1 U11286 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8871) );
  NAND2_X1 U11287 ( .A1(n8871), .A2(n10626), .ZN(n8878) );
  NAND2_X1 U11288 ( .A1(n8929), .A2(n8928), .ZN(n8940) );
  NAND2_X1 U11289 ( .A1(n11525), .A2(n11619), .ZN(n8765) );
  NAND2_X1 U11290 ( .A1(n9001), .A2(n15221), .ZN(n9015) );
  INV_X1 U11291 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9047) );
  INV_X1 U11292 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n12054) );
  INV_X1 U11293 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U11294 ( .A1(n9147), .A2(n9146), .ZN(n9159) );
  AND2_X1 U11295 ( .A1(n8785), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U11296 ( .A1(n8768), .A2(n8767), .ZN(n8772) );
  XNOR2_X2 U11297 ( .A(n8769), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8775) );
  NAND2_X1 U11298 ( .A1(n8770), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8771) );
  INV_X1 U11299 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12587) );
  NAND2_X1 U11300 ( .A1(n8893), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8777) );
  AND2_X2 U11301 ( .A1(n8775), .A2(n11879), .ZN(n9000) );
  NAND2_X1 U11302 ( .A1(n9306), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8776) );
  OAI211_X1 U11303 ( .C1(n12587), .C2(n9309), .A(n8777), .B(n8776), .ZN(n8778)
         );
  AOI21_X1 U11304 ( .B1(n12332), .B2(n9231), .A(n8778), .ZN(n9748) );
  NAND2_X1 U11305 ( .A1(n11963), .A2(n9748), .ZN(n9342) );
  INV_X1 U11306 ( .A(n8779), .ZN(n8780) );
  XNOR2_X1 U11307 ( .A(n8781), .B(n8780), .ZN(n11968) );
  NAND2_X1 U11308 ( .A1(n11968), .A2(n9143), .ZN(n8783) );
  NAND2_X1 U11309 ( .A1(n9161), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8784) );
  NAND2_X1 U11310 ( .A1(n8785), .A2(n8784), .ZN(n12345) );
  NAND2_X1 U11311 ( .A1(n12345), .A2(n9231), .ZN(n8791) );
  INV_X1 U11312 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n8788) );
  NAND2_X1 U11313 ( .A1(n8893), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U11314 ( .A1(n9306), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8786) );
  OAI211_X1 U11315 ( .C1(n8788), .C2(n9309), .A(n8787), .B(n8786), .ZN(n8789)
         );
  INV_X1 U11316 ( .A(n8789), .ZN(n8790) );
  NAND2_X1 U11317 ( .A1(n12523), .A2(n12353), .ZN(n9167) );
  NAND2_X1 U11318 ( .A1(n9473), .A2(n9167), .ZN(n12339) );
  XNOR2_X1 U11319 ( .A(n9901), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n8792) );
  XNOR2_X1 U11320 ( .A(n8793), .B(n8792), .ZN(n9886) );
  NAND2_X1 U11321 ( .A1(n8819), .A2(n9886), .ZN(n8797) );
  OR2_X1 U11322 ( .A1(n8839), .A2(SI_2_), .ZN(n8796) );
  OR2_X1 U11323 ( .A1(n10391), .A2(n10416), .ZN(n8795) );
  AND3_X2 U11324 ( .A1(n8797), .A2(n8796), .A3(n8795), .ZN(n15024) );
  INV_X1 U11325 ( .A(n15024), .ZN(n9188) );
  NAND2_X1 U11326 ( .A1(n9000), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8802) );
  NAND2_X1 U11327 ( .A1(n8823), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8801) );
  NAND2_X1 U11328 ( .A1(n8824), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8800) );
  INV_X1 U11329 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8798) );
  INV_X1 U11330 ( .A(n10786), .ZN(n15036) );
  NAND2_X1 U11331 ( .A1(n10786), .A2(n15024), .ZN(n9368) );
  NAND2_X1 U11332 ( .A1(n9000), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8807) );
  INV_X1 U11333 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U11334 ( .A1(n8823), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8804) );
  OAI21_X1 U11335 ( .B1(n8810), .B2(n8809), .A(n8808), .ZN(n9913) );
  NAND2_X1 U11336 ( .A1(n8819), .A2(n9913), .ZN(n8816) );
  NAND2_X1 U11337 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8812) );
  OR2_X1 U11338 ( .A1(n8817), .A2(n10456), .ZN(n8815) );
  NAND2_X1 U11339 ( .A1(n7333), .A2(n15031), .ZN(n9361) );
  INV_X1 U11340 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n15207) );
  XNOR2_X1 U11341 ( .A(n8818), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U11342 ( .A1(n8819), .A2(n9881), .ZN(n8820) );
  INV_X1 U11343 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8821) );
  OR2_X1 U11344 ( .A1(n8822), .A2(n8821), .ZN(n8828) );
  NAND2_X1 U11345 ( .A1(n9000), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U11346 ( .A1(n8823), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8826) );
  NOR2_X2 U11347 ( .A1(n10311), .A2(n15033), .ZN(n9359) );
  NAND2_X1 U11348 ( .A1(n9361), .A2(n9359), .ZN(n9771) );
  INV_X1 U11349 ( .A(n15031), .ZN(n10320) );
  NAND2_X1 U11350 ( .A1(n8830), .A2(n9368), .ZN(n10780) );
  NAND2_X1 U11351 ( .A1(n9000), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8836) );
  INV_X1 U11352 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U11353 ( .A1(n9134), .A2(n8831), .ZN(n8835) );
  NAND2_X1 U11354 ( .A1(n8893), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8834) );
  INV_X1 U11355 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8832) );
  XNOR2_X1 U11356 ( .A(n9896), .B(P2_DATAO_REG_3__SCAN_IN), .ZN(n8837) );
  XNOR2_X1 U11357 ( .A(n8838), .B(n8837), .ZN(n9909) );
  NAND2_X1 U11358 ( .A1(n8819), .A2(n9909), .ZN(n8845) );
  OR2_X1 U11359 ( .A1(n8839), .A2(SI_3_), .ZN(n8844) );
  OR2_X1 U11360 ( .A1(n8840), .A2(n8841), .ZN(n8842) );
  XNOR2_X1 U11361 ( .A(n8842), .B(P3_IR_REG_3__SCAN_IN), .ZN(n10647) );
  NAND2_X1 U11362 ( .A1(n15018), .A2(n10655), .ZN(n9376) );
  INV_X2 U11363 ( .A(n15018), .ZN(n12190) );
  INV_X1 U11364 ( .A(n10655), .ZN(n10791) );
  AND2_X1 U11365 ( .A1(n9376), .A2(n9372), .ZN(n10779) );
  NAND2_X1 U11366 ( .A1(n10780), .A2(n10779), .ZN(n10782) );
  AND2_X1 U11367 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8846) );
  NOR2_X1 U11368 ( .A1(n8871), .A2(n8846), .ZN(n15013) );
  INV_X1 U11369 ( .A(n15013), .ZN(n8847) );
  NAND2_X1 U11370 ( .A1(n9134), .A2(n8847), .ZN(n8852) );
  NAND2_X1 U11371 ( .A1(n8893), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U11372 ( .A1(n9000), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8850) );
  INV_X1 U11373 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8848) );
  OR2_X1 U11374 ( .A1(n9309), .A2(n8848), .ZN(n8849) );
  AND4_X2 U11375 ( .A1(n8852), .A2(n8851), .A3(n8850), .A4(n8849), .ZN(n14988)
         );
  XNOR2_X1 U11376 ( .A(n8853), .B(n8854), .ZN(n9903) );
  NAND2_X1 U11377 ( .A1(n8819), .A2(n9903), .ZN(n8861) );
  OR2_X1 U11378 ( .A1(n9088), .A2(SI_4_), .ZN(n8860) );
  INV_X1 U11379 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8855) );
  NAND2_X1 U11380 ( .A1(n8840), .A2(n8855), .ZN(n8857) );
  NAND2_X1 U11381 ( .A1(n8857), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8856) );
  MUX2_X1 U11382 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8856), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8858) );
  OR2_X1 U11383 ( .A1(n10391), .A2(n10724), .ZN(n8859) );
  NAND2_X1 U11384 ( .A1(n14988), .A2(n14999), .ZN(n9377) );
  INV_X1 U11385 ( .A(n14988), .ZN(n12189) );
  INV_X1 U11386 ( .A(n14999), .ZN(n8862) );
  NAND2_X1 U11387 ( .A1(n12189), .A2(n8862), .ZN(n9378) );
  NAND2_X1 U11388 ( .A1(n15002), .A2(n15004), .ZN(n8863) );
  NAND2_X1 U11389 ( .A1(n8863), .A2(n9377), .ZN(n14978) );
  XNOR2_X1 U11390 ( .A(n8865), .B(n8864), .ZN(n9906) );
  NAND2_X1 U11391 ( .A1(n8819), .A2(n9906), .ZN(n8869) );
  OR2_X1 U11392 ( .A1(n9088), .A2(SI_5_), .ZN(n8868) );
  NAND2_X1 U11393 ( .A1(n8889), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8866) );
  XNOR2_X1 U11394 ( .A(n8866), .B(P3_IR_REG_5__SCAN_IN), .ZN(n10634) );
  OR2_X1 U11395 ( .A1(n10391), .A2(n10634), .ZN(n8867) );
  INV_X1 U11396 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8870) );
  OR2_X1 U11397 ( .A1(n9309), .A2(n8870), .ZN(n8876) );
  NAND2_X1 U11398 ( .A1(n8893), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U11399 ( .A1(n9000), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8874) );
  OR2_X1 U11400 ( .A1(n8871), .A2(n10626), .ZN(n8872) );
  NAND2_X1 U11401 ( .A1(n8878), .A2(n8872), .ZN(n14995) );
  NAND2_X1 U11402 ( .A1(n9134), .A2(n14995), .ZN(n8873) );
  XNOR2_X2 U11403 ( .A(n14994), .B(n12188), .ZN(n14981) );
  NAND2_X1 U11404 ( .A1(n14978), .A2(n14981), .ZN(n8877) );
  INV_X1 U11405 ( .A(n12188), .ZN(n15005) );
  NAND2_X1 U11406 ( .A1(n15005), .A2(n14994), .ZN(n9382) );
  NAND2_X1 U11407 ( .A1(n8877), .A2(n9382), .ZN(n11090) );
  NAND2_X1 U11408 ( .A1(n6463), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8884) );
  NAND2_X1 U11409 ( .A1(n9306), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8883) );
  NAND2_X1 U11410 ( .A1(n8878), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8879) );
  NAND2_X1 U11411 ( .A1(n8894), .A2(n8879), .ZN(n11103) );
  NAND2_X1 U11412 ( .A1(n9134), .A2(n11103), .ZN(n8882) );
  INV_X1 U11413 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8880) );
  OR2_X1 U11414 ( .A1(n9309), .A2(n8880), .ZN(n8881) );
  INV_X1 U11415 ( .A(SI_6_), .ZN(n9911) );
  INV_X2 U11416 ( .A(n9305), .ZN(n9143) );
  NAND2_X1 U11417 ( .A1(n8886), .A2(n8885), .ZN(n8887) );
  NAND2_X1 U11418 ( .A1(n8888), .A2(n8887), .ZN(n9910) );
  NAND2_X1 U11419 ( .A1(n9143), .A2(n9910), .ZN(n8892) );
  NOR2_X1 U11420 ( .A1(n8889), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8904) );
  OR2_X1 U11421 ( .A1(n8904), .A2(n8841), .ZN(n8890) );
  XNOR2_X1 U11422 ( .A(n8890), .B(n8903), .ZN(n10675) );
  OR2_X1 U11423 ( .A1(n10391), .A2(n10675), .ZN(n8891) );
  OAI211_X1 U11424 ( .C1(n9088), .C2(n9911), .A(n8892), .B(n8891), .ZN(n10952)
         );
  NAND2_X1 U11425 ( .A1(n14987), .A2(n10952), .ZN(n9391) );
  INV_X1 U11426 ( .A(n10952), .ZN(n11102) );
  NAND2_X1 U11427 ( .A1(n14969), .A2(n11102), .ZN(n9389) );
  NAND2_X1 U11428 ( .A1(n9306), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U11429 ( .A1(n6463), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8899) );
  AND2_X1 U11430 ( .A1(n8894), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8895) );
  OR2_X1 U11431 ( .A1(n8895), .A2(n8911), .ZN(n14974) );
  NAND2_X1 U11432 ( .A1(n9231), .A2(n14974), .ZN(n8898) );
  INV_X1 U11433 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8896) );
  OR2_X1 U11434 ( .A1(n9309), .A2(n8896), .ZN(n8897) );
  XNOR2_X1 U11435 ( .A(n8902), .B(n8901), .ZN(n9917) );
  NAND2_X1 U11436 ( .A1(n9143), .A2(n9917), .ZN(n8908) );
  OR2_X1 U11437 ( .A1(n9088), .A2(SI_7_), .ZN(n8907) );
  NAND2_X1 U11438 ( .A1(n8904), .A2(n8903), .ZN(n8919) );
  NAND2_X1 U11439 ( .A1(n8919), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8905) );
  XNOR2_X1 U11440 ( .A(n8905), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11059) );
  OR2_X1 U11441 ( .A1(n10391), .A2(n11059), .ZN(n8906) );
  NAND2_X1 U11442 ( .A1(n11311), .A2(n11151), .ZN(n9393) );
  INV_X1 U11443 ( .A(n11151), .ZN(n14973) );
  NAND2_X1 U11444 ( .A1(n12187), .A2(n14973), .ZN(n9392) );
  INV_X1 U11445 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8909) );
  OR2_X1 U11446 ( .A1(n9309), .A2(n8909), .ZN(n8916) );
  NAND2_X1 U11447 ( .A1(n9000), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U11448 ( .A1(n6463), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8914) );
  NOR2_X1 U11449 ( .A1(n8911), .A2(n8910), .ZN(n8912) );
  OR2_X1 U11450 ( .A1(n8929), .A2(n8912), .ZN(n11307) );
  NAND2_X1 U11451 ( .A1(n9231), .A2(n11307), .ZN(n8913) );
  NAND4_X1 U11452 ( .A1(n8916), .A2(n8915), .A3(n8914), .A4(n8913), .ZN(n14968) );
  INV_X1 U11453 ( .A(SI_8_), .ZN(n9888) );
  XNOR2_X1 U11454 ( .A(n9954), .B(P2_DATAO_REG_8__SCAN_IN), .ZN(n8917) );
  XNOR2_X1 U11455 ( .A(n8918), .B(n8917), .ZN(n9887) );
  NAND2_X1 U11456 ( .A1(n9143), .A2(n9887), .ZN(n8925) );
  INV_X1 U11457 ( .A(n8950), .ZN(n8923) );
  NAND2_X1 U11458 ( .A1(n8920), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8921) );
  MUX2_X1 U11459 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8921), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8922) );
  NAND2_X1 U11460 ( .A1(n8923), .A2(n8922), .ZN(n11077) );
  OR2_X1 U11461 ( .A1(n10391), .A2(n11077), .ZN(n8924) );
  OAI211_X1 U11462 ( .C1(n9088), .C2(n9888), .A(n8925), .B(n8924), .ZN(n11315)
         );
  XNOR2_X1 U11463 ( .A(n14968), .B(n11315), .ZN(n11198) );
  INV_X1 U11464 ( .A(n14968), .ZN(n11458) );
  NAND2_X1 U11465 ( .A1(n11458), .A2(n11315), .ZN(n8926) );
  INV_X1 U11466 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n8927) );
  OR2_X1 U11467 ( .A1(n9309), .A2(n8927), .ZN(n8934) );
  OR2_X1 U11468 ( .A1(n8929), .A2(n8928), .ZN(n8930) );
  AND2_X1 U11469 ( .A1(n8940), .A2(n8930), .ZN(n14962) );
  INV_X1 U11470 ( .A(n14962), .ZN(n11490) );
  NAND2_X1 U11471 ( .A1(n9231), .A2(n11490), .ZN(n8933) );
  NAND2_X1 U11472 ( .A1(n6463), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U11473 ( .A1(n9306), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8931) );
  NAND4_X1 U11474 ( .A1(n8934), .A2(n8933), .A3(n8932), .A4(n8931), .ZN(n12186) );
  XNOR2_X1 U11475 ( .A(n9963), .B(P2_DATAO_REG_9__SCAN_IN), .ZN(n8935) );
  XNOR2_X1 U11476 ( .A(n8936), .B(n8935), .ZN(n9893) );
  NAND2_X1 U11477 ( .A1(n9143), .A2(n9893), .ZN(n8939) );
  OR2_X1 U11478 ( .A1(n8950), .A2(n8841), .ZN(n8937) );
  XNOR2_X1 U11479 ( .A(n8937), .B(P3_IR_REG_9__SCAN_IN), .ZN(n11233) );
  OR2_X1 U11480 ( .A1(n10391), .A2(n11233), .ZN(n8938) );
  OAI211_X1 U11481 ( .C1(n9088), .C2(SI_9_), .A(n8939), .B(n8938), .ZN(n14957)
         );
  NOR2_X1 U11482 ( .A1(n12186), .A2(n14957), .ZN(n9401) );
  NAND2_X1 U11483 ( .A1(n12186), .A2(n14957), .ZN(n9402) );
  NAND2_X1 U11484 ( .A1(n6463), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8946) );
  NAND2_X1 U11485 ( .A1(n9000), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8945) );
  NAND2_X1 U11486 ( .A1(n8940), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U11487 ( .A1(n8979), .A2(n8941), .ZN(n11668) );
  NAND2_X1 U11488 ( .A1(n9134), .A2(n11668), .ZN(n8944) );
  INV_X1 U11489 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8942) );
  OR2_X1 U11490 ( .A1(n9309), .A2(n8942), .ZN(n8943) );
  XNOR2_X1 U11491 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8947) );
  XNOR2_X1 U11492 ( .A(n8948), .B(n8947), .ZN(n9905) );
  NAND2_X1 U11493 ( .A1(n9905), .A2(n9143), .ZN(n8954) );
  INV_X1 U11494 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U11495 ( .A1(n8950), .A2(n8949), .ZN(n8962) );
  NAND2_X1 U11496 ( .A1(n8962), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8951) );
  XNOR2_X1 U11497 ( .A(n8951), .B(P3_IR_REG_10__SCAN_IN), .ZN(n11529) );
  OAI22_X1 U11498 ( .A1(n9295), .A2(SI_10_), .B1(n11529), .B2(n10391), .ZN(
        n8952) );
  INV_X1 U11499 ( .A(n8952), .ZN(n8953) );
  NAND2_X1 U11500 ( .A1(n12140), .A2(n9789), .ZN(n9407) );
  NAND2_X1 U11501 ( .A1(n12185), .A2(n11671), .ZN(n9406) );
  INV_X1 U11502 ( .A(n11509), .ZN(n8968) );
  NAND2_X1 U11503 ( .A1(n6463), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U11504 ( .A1(n9306), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8958) );
  XNOR2_X1 U11505 ( .A(n8979), .B(P3_REG3_REG_11__SCAN_IN), .ZN(n12144) );
  NAND2_X1 U11506 ( .A1(n9231), .A2(n12144), .ZN(n8957) );
  INV_X1 U11507 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n8955) );
  OR2_X1 U11508 ( .A1(n9309), .A2(n8955), .ZN(n8956) );
  XNOR2_X1 U11509 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8960) );
  XNOR2_X1 U11510 ( .A(n8961), .B(n8960), .ZN(n9949) );
  NAND2_X1 U11511 ( .A1(n9949), .A2(n9143), .ZN(n8966) );
  OAI21_X1 U11512 ( .B1(n8962), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8963) );
  XNOR2_X1 U11513 ( .A(n8963), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11610) );
  INV_X1 U11514 ( .A(n11610), .ZN(n9950) );
  OAI22_X1 U11515 ( .A1(n9295), .A2(n9952), .B1(n10391), .B2(n9950), .ZN(n8964) );
  INV_X1 U11516 ( .A(n8964), .ZN(n8965) );
  NAND2_X1 U11517 ( .A1(n8966), .A2(n8965), .ZN(n11505) );
  NAND2_X1 U11518 ( .A1(n14347), .A2(n11505), .ZN(n9409) );
  INV_X1 U11519 ( .A(n11505), .ZN(n12137) );
  NAND2_X1 U11520 ( .A1(n12137), .A2(n12184), .ZN(n9413) );
  NAND2_X1 U11521 ( .A1(n9409), .A2(n9413), .ZN(n11508) );
  XNOR2_X1 U11522 ( .A(n8970), .B(n8969), .ZN(n9960) );
  NAND2_X1 U11523 ( .A1(n9960), .A2(n9143), .ZN(n8977) );
  NAND2_X1 U11524 ( .A1(n8971), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8972) );
  MUX2_X1 U11525 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8972), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8974) );
  AND2_X1 U11526 ( .A1(n8974), .A2(n8973), .ZN(n11618) );
  OAI22_X1 U11527 ( .A1(n9295), .A2(SI_12_), .B1(n11618), .B2(n10391), .ZN(
        n8975) );
  INV_X1 U11528 ( .A(n8975), .ZN(n8976) );
  NAND2_X1 U11529 ( .A1(n8977), .A2(n8976), .ZN(n14348) );
  INV_X1 U11530 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8978) );
  OR2_X1 U11531 ( .A1(n9309), .A2(n8978), .ZN(n8984) );
  NAND2_X1 U11532 ( .A1(n6463), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8983) );
  NAND2_X1 U11533 ( .A1(n9306), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8982) );
  OAI21_X1 U11534 ( .B1(n8979), .B2(P3_REG3_REG_11__SCAN_IN), .A(
        P3_REG3_REG_12__SCAN_IN), .ZN(n8980) );
  NAND2_X1 U11535 ( .A1(n8980), .A2(n8988), .ZN(n14349) );
  NAND2_X1 U11536 ( .A1(n9134), .A2(n14349), .ZN(n8981) );
  NAND4_X1 U11537 ( .A1(n8984), .A2(n8983), .A3(n8982), .A4(n8981), .ZN(n12183) );
  OR2_X1 U11538 ( .A1(n14348), .A2(n12183), .ZN(n9417) );
  NAND2_X1 U11539 ( .A1(n14348), .A2(n12183), .ZN(n9415) );
  XNOR2_X1 U11540 ( .A(n8985), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9970) );
  NAND2_X1 U11541 ( .A1(n8973), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8986) );
  XNOR2_X1 U11542 ( .A(n8986), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12210) );
  OAI22_X1 U11543 ( .A1(n9088), .A2(SI_13_), .B1(n12210), .B2(n10391), .ZN(
        n8987) );
  AOI21_X1 U11544 ( .B1(n9970), .B2(n9143), .A(n8987), .ZN(n12125) );
  NAND2_X1 U11545 ( .A1(n6463), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U11546 ( .A1(n9306), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8992) );
  AND2_X1 U11547 ( .A1(n8988), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8989) );
  OR2_X1 U11548 ( .A1(n8989), .A2(n9001), .ZN(n12517) );
  NAND2_X1 U11549 ( .A1(n9231), .A2(n12517), .ZN(n8991) );
  INV_X1 U11550 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12635) );
  OR2_X1 U11551 ( .A1(n9309), .A2(n12635), .ZN(n8990) );
  AND2_X1 U11552 ( .A1(n12125), .A2(n12029), .ZN(n9206) );
  INV_X1 U11553 ( .A(n12125), .ZN(n12637) );
  NAND2_X1 U11554 ( .A1(n12637), .A2(n14344), .ZN(n9422) );
  XNOR2_X1 U11555 ( .A(n8994), .B(n6611), .ZN(n10098) );
  NAND2_X1 U11556 ( .A1(n10098), .A2(n9143), .ZN(n8999) );
  OR2_X1 U11557 ( .A1(n8995), .A2(n8841), .ZN(n8996) );
  XNOR2_X1 U11558 ( .A(n8996), .B(n9010), .ZN(n12197) );
  OAI22_X1 U11559 ( .A1(n9295), .A2(n10099), .B1(n10391), .B2(n12197), .ZN(
        n8997) );
  INV_X1 U11560 ( .A(n8997), .ZN(n8998) );
  NAND2_X1 U11561 ( .A1(n8999), .A2(n8998), .ZN(n12031) );
  NAND2_X1 U11562 ( .A1(n6463), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9006) );
  NAND2_X1 U11563 ( .A1(n9000), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9005) );
  OR2_X1 U11564 ( .A1(n9001), .A2(n15221), .ZN(n9002) );
  NAND2_X1 U11565 ( .A1(n9015), .A2(n9002), .ZN(n12026) );
  NAND2_X1 U11566 ( .A1(n9231), .A2(n12026), .ZN(n9004) );
  INV_X1 U11567 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12631) );
  OR2_X1 U11568 ( .A1(n9309), .A2(n12631), .ZN(n9003) );
  OR2_X1 U11569 ( .A1(n12031), .A2(n12514), .ZN(n9426) );
  NAND2_X1 U11570 ( .A1(n12031), .A2(n12514), .ZN(n9435) );
  NAND2_X1 U11571 ( .A1(n9426), .A2(n9435), .ZN(n11806) );
  INV_X1 U11572 ( .A(n9007), .ZN(n9008) );
  XNOR2_X1 U11573 ( .A(n9009), .B(n9008), .ZN(n10171) );
  NAND2_X1 U11574 ( .A1(n10171), .A2(n9143), .ZN(n9014) );
  OR2_X1 U11575 ( .A1(n9026), .A2(n8841), .ZN(n9011) );
  XNOR2_X1 U11576 ( .A(n9011), .B(n9025), .ZN(n12260) );
  OAI22_X1 U11577 ( .A1(n9295), .A2(n10172), .B1(n10391), .B2(n12260), .ZN(
        n9012) );
  INV_X1 U11578 ( .A(n9012), .ZN(n9013) );
  INV_X1 U11579 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12627) );
  OR2_X1 U11580 ( .A1(n9309), .A2(n12627), .ZN(n9020) );
  NAND2_X1 U11581 ( .A1(n6463), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U11582 ( .A1(n9306), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n9018) );
  NAND2_X1 U11583 ( .A1(n9015), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9016) );
  NAND2_X1 U11584 ( .A1(n9035), .A2(n9016), .ZN(n12503) );
  NAND2_X1 U11585 ( .A1(n9134), .A2(n12503), .ZN(n9017) );
  NAND4_X1 U11586 ( .A1(n9020), .A2(n9019), .A3(n9018), .A4(n9017), .ZN(n12482) );
  XNOR2_X1 U11587 ( .A(n12166), .B(n12482), .ZN(n12501) );
  NAND2_X1 U11588 ( .A1(n12502), .A2(n12501), .ZN(n9021) );
  NAND2_X1 U11589 ( .A1(n12166), .A2(n9801), .ZN(n9433) );
  NAND2_X1 U11590 ( .A1(n9021), .A2(n9433), .ZN(n12486) );
  INV_X1 U11591 ( .A(n9022), .ZN(n9023) );
  XNOR2_X1 U11592 ( .A(n9024), .B(n9023), .ZN(n10245) );
  NAND2_X1 U11593 ( .A1(n10245), .A2(n9143), .ZN(n9034) );
  NOR2_X1 U11594 ( .A1(n9030), .A2(n8841), .ZN(n9027) );
  MUX2_X1 U11595 ( .A(n8841), .B(n9027), .S(P3_IR_REG_16__SCAN_IN), .Z(n9028)
         );
  INV_X1 U11596 ( .A(n9028), .ZN(n9031) );
  NAND2_X1 U11597 ( .A1(n9031), .A2(n9056), .ZN(n12280) );
  OAI22_X1 U11598 ( .A1(n9088), .A2(n10246), .B1(n10391), .B2(n12280), .ZN(
        n9032) );
  INV_X1 U11599 ( .A(n9032), .ZN(n9033) );
  NAND2_X1 U11600 ( .A1(n9034), .A2(n9033), .ZN(n12567) );
  NAND2_X1 U11601 ( .A1(n6463), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n9040) );
  NAND2_X1 U11602 ( .A1(n9306), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n9039) );
  AND2_X1 U11603 ( .A1(n9035), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9036) );
  OR2_X1 U11604 ( .A1(n9036), .A2(n9048), .ZN(n12489) );
  NAND2_X1 U11605 ( .A1(n9231), .A2(n12489), .ZN(n9038) );
  INV_X1 U11606 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n15131) );
  OR2_X1 U11607 ( .A1(n9309), .A2(n15131), .ZN(n9037) );
  OR2_X1 U11608 ( .A1(n12567), .A2(n12500), .ZN(n9437) );
  NAND2_X1 U11609 ( .A1(n12567), .A2(n12500), .ZN(n9434) );
  XNOR2_X1 U11610 ( .A(n15219), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n9041) );
  XNOR2_X1 U11611 ( .A(n9042), .B(n9041), .ZN(n10326) );
  NAND2_X1 U11612 ( .A1(n10326), .A2(n9143), .ZN(n9046) );
  NAND2_X1 U11613 ( .A1(n9056), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9043) );
  XNOR2_X1 U11614 ( .A(n9043), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12303) );
  OAI22_X1 U11615 ( .A1(n9295), .A2(n10327), .B1(n10391), .B2(n12296), .ZN(
        n9044) );
  INV_X1 U11616 ( .A(n9044), .ZN(n9045) );
  INV_X1 U11617 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12621) );
  OR2_X1 U11618 ( .A1(n9309), .A2(n12621), .ZN(n9053) );
  NAND2_X1 U11619 ( .A1(n6463), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U11620 ( .A1(n9306), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9051) );
  NOR2_X1 U11621 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  OR2_X1 U11622 ( .A1(n9063), .A2(n9049), .ZN(n12472) );
  NAND2_X1 U11623 ( .A1(n9231), .A2(n12472), .ZN(n9050) );
  NAND4_X1 U11624 ( .A1(n9053), .A2(n9052), .A3(n9051), .A4(n9050), .ZN(n12481) );
  XNOR2_X1 U11625 ( .A(n12095), .B(n12481), .ZN(n12470) );
  INV_X1 U11626 ( .A(n12481), .ZN(n12088) );
  XNOR2_X1 U11627 ( .A(n9055), .B(n9054), .ZN(n10420) );
  NAND2_X1 U11628 ( .A1(n10420), .A2(n9143), .ZN(n9061) );
  NAND2_X1 U11629 ( .A1(n9074), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9058) );
  XNOR2_X1 U11630 ( .A(n9058), .B(n9057), .ZN(n12306) );
  OAI22_X1 U11631 ( .A1(n9088), .A2(n10421), .B1(n10391), .B2(n12306), .ZN(
        n9059) );
  INV_X1 U11632 ( .A(n9059), .ZN(n9060) );
  NAND2_X1 U11633 ( .A1(n9061), .A2(n9060), .ZN(n12559) );
  NAND2_X1 U11634 ( .A1(n9306), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9069) );
  OR2_X1 U11635 ( .A1(n9063), .A2(n9062), .ZN(n9064) );
  NAND2_X1 U11636 ( .A1(n9079), .A2(n9064), .ZN(n12458) );
  NAND2_X1 U11637 ( .A1(n9134), .A2(n12458), .ZN(n9068) );
  NAND2_X1 U11638 ( .A1(n6463), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9067) );
  INV_X1 U11639 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n9065) );
  OR2_X1 U11640 ( .A1(n9309), .A2(n9065), .ZN(n9066) );
  OR2_X1 U11641 ( .A1(n12559), .A2(n12440), .ZN(n12442) );
  NAND2_X1 U11642 ( .A1(n12559), .A2(n12440), .ZN(n9443) );
  NAND2_X1 U11643 ( .A1(n12442), .A2(n9443), .ZN(n12457) );
  INV_X1 U11644 ( .A(n9071), .ZN(n9072) );
  XNOR2_X1 U11645 ( .A(n9073), .B(n9072), .ZN(n10458) );
  NAND2_X1 U11646 ( .A1(n10458), .A2(n9143), .ZN(n9078) );
  OAI22_X1 U11647 ( .A1(n9295), .A2(SI_19_), .B1(n9767), .B2(n10391), .ZN(
        n9076) );
  INV_X1 U11648 ( .A(n9076), .ZN(n9077) );
  NAND2_X1 U11649 ( .A1(n6463), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U11650 ( .A1(n9306), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U11651 ( .A1(n9079), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9080) );
  NAND2_X1 U11652 ( .A1(n9091), .A2(n9080), .ZN(n12446) );
  NAND2_X1 U11653 ( .A1(n9231), .A2(n12446), .ZN(n9082) );
  INV_X1 U11654 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12616) );
  OR2_X1 U11655 ( .A1(n9309), .A2(n12616), .ZN(n9081) );
  XNOR2_X1 U11656 ( .A(n12618), .B(n12427), .ZN(n12444) );
  AND2_X1 U11657 ( .A1(n12444), .A2(n12442), .ZN(n9085) );
  OR2_X1 U11658 ( .A1(n12618), .A2(n12452), .ZN(n9449) );
  XNOR2_X1 U11659 ( .A(n9087), .B(n9086), .ZN(n10658) );
  NAND2_X1 U11660 ( .A1(n10658), .A2(n9143), .ZN(n9090) );
  AND2_X1 U11661 ( .A1(n9091), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9092) );
  OR2_X1 U11662 ( .A1(n9092), .A2(n9102), .ZN(n12433) );
  NAND2_X1 U11663 ( .A1(n12433), .A2(n9231), .ZN(n9095) );
  AOI22_X1 U11664 ( .A1(n6463), .A2(P3_REG1_REG_20__SCAN_IN), .B1(n9306), .B2(
        P3_REG2_REG_20__SCAN_IN), .ZN(n9094) );
  INV_X1 U11665 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12612) );
  OR2_X1 U11666 ( .A1(n9309), .A2(n12612), .ZN(n9093) );
  NAND2_X1 U11667 ( .A1(n12614), .A2(n12182), .ZN(n9097) );
  NAND2_X1 U11668 ( .A1(n12432), .A2(n9097), .ZN(n12418) );
  XNOR2_X1 U11669 ( .A(n9099), .B(n8735), .ZN(n10878) );
  NAND2_X1 U11670 ( .A1(n10878), .A2(n9143), .ZN(n9101) );
  INV_X1 U11671 ( .A(SI_21_), .ZN(n10880) );
  NOR2_X1 U11672 ( .A1(n9102), .A2(n12054), .ZN(n9103) );
  OR2_X1 U11673 ( .A1(n9112), .A2(n9103), .ZN(n12419) );
  NAND2_X1 U11674 ( .A1(n12419), .A2(n9134), .ZN(n9106) );
  AOI22_X1 U11675 ( .A1(n6463), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n9306), .B2(
        P3_REG2_REG_21__SCAN_IN), .ZN(n9105) );
  INV_X1 U11676 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12608) );
  OR2_X1 U11677 ( .A1(n9309), .A2(n12608), .ZN(n9104) );
  NAND2_X1 U11678 ( .A1(n12050), .A2(n12428), .ZN(n9354) );
  XNOR2_X1 U11679 ( .A(n9108), .B(n7305), .ZN(n11032) );
  NAND2_X1 U11680 ( .A1(n11032), .A2(n9143), .ZN(n9110) );
  OR2_X1 U11681 ( .A1(n9112), .A2(n9111), .ZN(n9113) );
  NAND2_X1 U11682 ( .A1(n9121), .A2(n9113), .ZN(n12407) );
  NAND2_X1 U11683 ( .A1(n12407), .A2(n9231), .ZN(n9116) );
  AOI22_X1 U11684 ( .A1(n8893), .A2(P3_REG1_REG_22__SCAN_IN), .B1(n9306), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n9115) );
  INV_X1 U11685 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n15236) );
  OR2_X1 U11686 ( .A1(n9309), .A2(n15236), .ZN(n9114) );
  NAND2_X1 U11687 ( .A1(n12406), .A2(n12416), .ZN(n9352) );
  XNOR2_X1 U11688 ( .A(n9118), .B(n9117), .ZN(n11319) );
  NAND2_X1 U11689 ( .A1(n11319), .A2(n9143), .ZN(n9120) );
  OR2_X1 U11690 ( .A1(n9295), .A2(n11322), .ZN(n9119) );
  NAND2_X1 U11691 ( .A1(n9121), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9122) );
  NAND2_X1 U11692 ( .A1(n9132), .A2(n9122), .ZN(n12396) );
  NAND2_X1 U11693 ( .A1(n12396), .A2(n9231), .ZN(n9128) );
  INV_X1 U11694 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n9125) );
  NAND2_X1 U11695 ( .A1(n9306), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9124) );
  NAND2_X1 U11696 ( .A1(n8893), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9123) );
  OAI211_X1 U11697 ( .C1(n9309), .C2(n9125), .A(n9124), .B(n9123), .ZN(n9126)
         );
  INV_X1 U11698 ( .A(n9126), .ZN(n9127) );
  NAND2_X1 U11699 ( .A1(n12542), .A2(n12378), .ZN(n9351) );
  NAND2_X1 U11700 ( .A1(n9819), .A2(n9824), .ZN(n9350) );
  XNOR2_X1 U11701 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9129), .ZN(n11699) );
  NAND2_X1 U11702 ( .A1(n11699), .A2(n9143), .ZN(n9131) );
  INV_X1 U11703 ( .A(SI_24_), .ZN(n11701) );
  AND2_X1 U11704 ( .A1(n9132), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9133) );
  OR2_X1 U11705 ( .A1(n9133), .A2(n9147), .ZN(n12383) );
  NAND2_X1 U11706 ( .A1(n12383), .A2(n9134), .ZN(n9139) );
  INV_X1 U11707 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12600) );
  NAND2_X1 U11708 ( .A1(n9306), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9136) );
  NAND2_X1 U11709 ( .A1(n8893), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9135) );
  OAI211_X1 U11710 ( .C1(n12600), .C2(n9309), .A(n9136), .B(n9135), .ZN(n9137)
         );
  INV_X1 U11711 ( .A(n9137), .ZN(n9138) );
  NAND2_X1 U11712 ( .A1(n12602), .A2(n12364), .ZN(n9349) );
  INV_X1 U11713 ( .A(n12602), .ZN(n9218) );
  NAND2_X1 U11714 ( .A1(n9218), .A2(n12389), .ZN(n9348) );
  NAND2_X1 U11715 ( .A1(n9349), .A2(n9348), .ZN(n12376) );
  XNOR2_X1 U11716 ( .A(n9142), .B(n6764), .ZN(n11763) );
  NAND2_X1 U11717 ( .A1(n11763), .A2(n9143), .ZN(n9145) );
  OR2_X1 U11718 ( .A1(n9147), .A2(n9146), .ZN(n9148) );
  NAND2_X1 U11719 ( .A1(n9159), .A2(n9148), .ZN(n12370) );
  NAND2_X1 U11720 ( .A1(n12370), .A2(n9231), .ZN(n9153) );
  INV_X1 U11721 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12596) );
  NAND2_X1 U11722 ( .A1(n9306), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9150) );
  NAND2_X1 U11723 ( .A1(n8893), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9149) );
  OAI211_X1 U11724 ( .C1(n9309), .C2(n12596), .A(n9150), .B(n9149), .ZN(n9151)
         );
  INV_X1 U11725 ( .A(n9151), .ZN(n9152) );
  XNOR2_X1 U11726 ( .A(n12072), .B(n12379), .ZN(n12368) );
  NAND2_X1 U11727 ( .A1(n12072), .A2(n12352), .ZN(n9344) );
  INV_X1 U11728 ( .A(n9154), .ZN(n9155) );
  XNOR2_X1 U11729 ( .A(n9156), .B(n9155), .ZN(n11850) );
  NAND2_X1 U11730 ( .A1(n11850), .A2(n9143), .ZN(n9158) );
  NAND2_X1 U11731 ( .A1(n9159), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9160) );
  NAND2_X1 U11732 ( .A1(n9161), .A2(n9160), .ZN(n12356) );
  NAND2_X1 U11733 ( .A1(n12356), .A2(n9231), .ZN(n9166) );
  INV_X1 U11734 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12592) );
  NAND2_X1 U11735 ( .A1(n8893), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9163) );
  NAND2_X1 U11736 ( .A1(n9306), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9162) );
  OAI211_X1 U11737 ( .C1(n12592), .C2(n9309), .A(n9163), .B(n9162), .ZN(n9164)
         );
  INV_X1 U11738 ( .A(n9164), .ZN(n9165) );
  NAND2_X1 U11739 ( .A1(n12155), .A2(n12367), .ZN(n9222) );
  INV_X1 U11740 ( .A(n9222), .ZN(n9472) );
  XNOR2_X1 U11741 ( .A(n11952), .B(n9289), .ZN(n12331) );
  INV_X1 U11742 ( .A(n9168), .ZN(n9169) );
  NAND2_X1 U11743 ( .A1(n8995), .A2(n9169), .ZN(n9175) );
  NAND2_X1 U11744 ( .A1(n9177), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9172) );
  MUX2_X1 U11745 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9172), .S(
        P3_IR_REG_21__SCAN_IN), .Z(n9173) );
  OR2_X1 U11746 ( .A1(n9767), .A2(n9230), .ZN(n9181) );
  NAND2_X1 U11747 ( .A1(n9255), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9174) );
  NAND2_X1 U11748 ( .A1(n9175), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9176) );
  MUX2_X1 U11749 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9176), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n9178) );
  NAND2_X1 U11750 ( .A1(n10881), .A2(n10661), .ZN(n9179) );
  XNOR2_X1 U11751 ( .A(n11033), .B(n9179), .ZN(n9180) );
  NAND2_X1 U11752 ( .A1(n9181), .A2(n9180), .ZN(n9847) );
  INV_X1 U11753 ( .A(n9767), .ZN(n10459) );
  NAND3_X1 U11754 ( .A1(n9847), .A2(n9492), .A3(n15030), .ZN(n9183) );
  NAND2_X1 U11755 ( .A1(n11033), .A2(n9338), .ZN(n9182) );
  OR2_X1 U11756 ( .A1(n9767), .A2(n9182), .ZN(n9276) );
  AND2_X1 U11757 ( .A1(n9183), .A2(n9276), .ZN(n15043) );
  OR2_X1 U11758 ( .A1(n15044), .A2(n11033), .ZN(n15052) );
  INV_X1 U11759 ( .A(n15037), .ZN(n9185) );
  NAND2_X1 U11760 ( .A1(n9322), .A2(n9185), .ZN(n9187) );
  NAND2_X1 U11761 ( .A1(n8829), .A2(n15031), .ZN(n9186) );
  NAND2_X1 U11762 ( .A1(n9187), .A2(n9186), .ZN(n15016) );
  NAND2_X1 U11763 ( .A1(n15015), .A2(n15016), .ZN(n15014) );
  NAND2_X1 U11764 ( .A1(n10786), .A2(n9188), .ZN(n9189) );
  AND2_X2 U11765 ( .A1(n15014), .A2(n9189), .ZN(n10785) );
  INV_X1 U11766 ( .A(n10779), .ZN(n10784) );
  NAND2_X1 U11767 ( .A1(n12190), .A2(n10655), .ZN(n9190) );
  NAND2_X1 U11768 ( .A1(n10783), .A2(n9190), .ZN(n14979) );
  INV_X1 U11769 ( .A(n15004), .ZN(n15001) );
  INV_X1 U11770 ( .A(n14994), .ZN(n9386) );
  NAND2_X1 U11771 ( .A1(n15005), .A2(n9386), .ZN(n9192) );
  AND2_X1 U11772 ( .A1(n15001), .A2(n9192), .ZN(n9191) );
  NAND2_X1 U11773 ( .A1(n14979), .A2(n9191), .ZN(n9196) );
  INV_X1 U11774 ( .A(n9192), .ZN(n9194) );
  NAND2_X1 U11775 ( .A1(n12189), .A2(n14999), .ZN(n14980) );
  OR2_X1 U11776 ( .A1(n9194), .A2(n14982), .ZN(n9195) );
  NAND2_X1 U11777 ( .A1(n9196), .A2(n9195), .ZN(n11095) );
  INV_X1 U11778 ( .A(n11089), .ZN(n11094) );
  NAND2_X1 U11779 ( .A1(n11095), .A2(n11094), .ZN(n11093) );
  NAND2_X1 U11780 ( .A1(n14969), .A2(n10952), .ZN(n9197) );
  NAND2_X1 U11781 ( .A1(n11093), .A2(n9197), .ZN(n14966) );
  INV_X1 U11782 ( .A(n14965), .ZN(n14963) );
  NAND2_X1 U11783 ( .A1(n14966), .A2(n14963), .ZN(n9199) );
  NAND2_X1 U11784 ( .A1(n12187), .A2(n11151), .ZN(n9198) );
  AND2_X1 U11785 ( .A1(n14968), .A2(n11315), .ZN(n9200) );
  INV_X1 U11786 ( .A(n14957), .ZN(n9201) );
  XNOR2_X1 U11787 ( .A(n12186), .B(n9201), .ZN(n11456) );
  NAND2_X1 U11788 ( .A1(n12186), .A2(n9201), .ZN(n9202) );
  NAND2_X1 U11789 ( .A1(n11460), .A2(n9202), .ZN(n11407) );
  NAND2_X1 U11790 ( .A1(n11407), .A2(n11410), .ZN(n11406) );
  NAND2_X1 U11791 ( .A1(n12185), .A2(n9789), .ZN(n9203) );
  NAND2_X1 U11792 ( .A1(n11406), .A2(n9203), .ZN(n11502) );
  NAND2_X1 U11793 ( .A1(n11502), .A2(n11508), .ZN(n11501) );
  NAND2_X1 U11794 ( .A1(n12184), .A2(n11505), .ZN(n9204) );
  NAND2_X1 U11795 ( .A1(n11501), .A2(n9204), .ZN(n14343) );
  INV_X1 U11796 ( .A(n14339), .ZN(n14342) );
  INV_X1 U11797 ( .A(n12183), .ZN(n12513) );
  OR2_X1 U11798 ( .A1(n14348), .A2(n12513), .ZN(n9205) );
  INV_X1 U11799 ( .A(n9206), .ZN(n9421) );
  NAND2_X1 U11800 ( .A1(n9421), .A2(n9422), .ZN(n9418) );
  OR2_X1 U11801 ( .A1(n12125), .A2(n14344), .ZN(n11802) );
  AND2_X1 U11802 ( .A1(n11806), .A2(n11802), .ZN(n9207) );
  NAND2_X1 U11803 ( .A1(n12508), .A2(n9207), .ZN(n11801) );
  NAND2_X1 U11804 ( .A1(n12031), .A2(n12497), .ZN(n9208) );
  NAND2_X1 U11805 ( .A1(n11801), .A2(n9208), .ZN(n12496) );
  INV_X1 U11806 ( .A(n12501), .ZN(n12495) );
  NAND2_X1 U11807 ( .A1(n12166), .A2(n12482), .ZN(n9209) );
  INV_X1 U11808 ( .A(n12500), .ZN(n12467) );
  OR2_X1 U11809 ( .A1(n12567), .A2(n12467), .ZN(n9211) );
  NAND2_X1 U11810 ( .A1(n12095), .A2(n12481), .ZN(n9212) );
  AND2_X1 U11811 ( .A1(n12618), .A2(n12427), .ZN(n9213) );
  OAI22_X1 U11812 ( .A1(n12438), .A2(n9213), .B1(n12427), .B2(n12618), .ZN(
        n12424) );
  NAND2_X1 U11813 ( .A1(n12115), .A2(n12182), .ZN(n9214) );
  OR2_X1 U11814 ( .A1(n12050), .A2(n12181), .ZN(n9216) );
  OR2_X1 U11815 ( .A1(n12406), .A2(n12180), .ZN(n9217) );
  NAND2_X1 U11816 ( .A1(n12377), .A2(n12376), .ZN(n12375) );
  NAND2_X1 U11817 ( .A1(n9218), .A2(n12364), .ZN(n9219) );
  NAND2_X1 U11818 ( .A1(n12375), .A2(n9219), .ZN(n12363) );
  INV_X1 U11819 ( .A(n12368), .ZN(n12362) );
  NAND2_X1 U11820 ( .A1(n12363), .A2(n12362), .ZN(n12361) );
  NAND2_X1 U11821 ( .A1(n12072), .A2(n12379), .ZN(n9220) );
  NAND2_X1 U11822 ( .A1(n12361), .A2(n9220), .ZN(n12350) );
  OR2_X1 U11823 ( .A1(n12155), .A2(n12340), .ZN(n9221) );
  NAND2_X1 U11824 ( .A1(n12355), .A2(n12155), .ZN(n9224) );
  INV_X1 U11825 ( .A(n12339), .ZN(n12344) );
  OR2_X1 U11826 ( .A1(n12523), .A2(n12179), .ZN(n9226) );
  INV_X1 U11827 ( .A(n11952), .ZN(n9227) );
  NAND2_X1 U11828 ( .A1(n9767), .A2(n11033), .ZN(n9754) );
  NAND2_X1 U11829 ( .A1(n9230), .A2(n9338), .ZN(n9340) );
  NAND3_X1 U11830 ( .A1(n9744), .A2(n9229), .A3(n15039), .ZN(n9239) );
  OR2_X1 U11831 ( .A1(n11876), .A2(n12198), .ZN(n10402) );
  NAND2_X1 U11832 ( .A1(n10402), .A2(n10391), .ZN(n9845) );
  INV_X1 U11833 ( .A(n9845), .ZN(n9859) );
  NOR2_X1 U11834 ( .A1(n12353), .A2(n15019), .ZN(n9237) );
  NAND2_X1 U11835 ( .A1(n14333), .A2(n9231), .ZN(n9312) );
  INV_X1 U11836 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U11837 ( .A1(n9306), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9233) );
  NAND2_X1 U11838 ( .A1(n8893), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9232) );
  OAI211_X1 U11839 ( .C1(n9309), .C2(n9234), .A(n9233), .B(n9232), .ZN(n9235)
         );
  INV_X1 U11840 ( .A(n9235), .ZN(n9236) );
  INV_X1 U11841 ( .A(n11958), .ZN(n12178) );
  AOI21_X1 U11842 ( .B1(n12331), .B2(n14362), .A(n12336), .ZN(n12586) );
  NAND2_X1 U11843 ( .A1(n6500), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9240) );
  MUX2_X1 U11844 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9240), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n9242) );
  NAND2_X1 U11845 ( .A1(n9243), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9244) );
  MUX2_X1 U11846 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9244), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n9245) );
  INV_X1 U11847 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9247) );
  INV_X1 U11848 ( .A(n11702), .ZN(n9248) );
  OR2_X1 U11849 ( .A1(n9252), .A2(n9248), .ZN(n9249) );
  INV_X1 U11850 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9251) );
  NAND2_X1 U11851 ( .A1(n6612), .A2(n9251), .ZN(n9254) );
  INV_X1 U11852 ( .A(n9252), .ZN(n11853) );
  NAND2_X1 U11853 ( .A1(n11853), .A2(n11764), .ZN(n9253) );
  XNOR2_X1 U11854 ( .A(n9770), .B(n12639), .ZN(n9271) );
  NOR2_X1 U11855 ( .A1(n11764), .A2(n11702), .ZN(n9258) );
  NAND2_X1 U11856 ( .A1(n9252), .A2(n9258), .ZN(n9870) );
  INV_X1 U11857 ( .A(n6612), .ZN(n9948) );
  NOR2_X1 U11858 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_24__SCAN_IN), .ZN(
        n9262) );
  NOR4_X1 U11859 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n9261) );
  NOR4_X1 U11860 ( .A1(P3_D_REG_27__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n9260) );
  NOR4_X1 U11861 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_20__SCAN_IN), .A3(
        P3_D_REG_19__SCAN_IN), .A4(P3_D_REG_18__SCAN_IN), .ZN(n9259) );
  NAND4_X1 U11862 ( .A1(n9262), .A2(n9261), .A3(n9260), .A4(n9259), .ZN(n9268)
         );
  NOR4_X1 U11863 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9266) );
  NOR4_X1 U11864 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9265) );
  NOR4_X1 U11865 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9264) );
  NOR4_X1 U11866 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9263) );
  NAND4_X1 U11867 ( .A1(n9266), .A2(n9265), .A3(n9264), .A4(n9263), .ZN(n9267)
         );
  NOR2_X1 U11868 ( .A1(n9268), .A2(n9267), .ZN(n9269) );
  NOR2_X1 U11869 ( .A1(n9948), .A2(n9269), .ZN(n9756) );
  NOR2_X1 U11870 ( .A1(n10387), .A2(n9756), .ZN(n9270) );
  INV_X1 U11871 ( .A(n9492), .ZN(n9500) );
  INV_X1 U11872 ( .A(n11033), .ZN(n9273) );
  NAND2_X1 U11873 ( .A1(n15023), .A2(n10661), .ZN(n9272) );
  OAI21_X1 U11874 ( .B1(n9767), .B2(n9273), .A(n9272), .ZN(n9274) );
  AOI21_X1 U11875 ( .B1(n9500), .B2(n9274), .A(n10389), .ZN(n9275) );
  NAND2_X1 U11876 ( .A1(n9276), .A2(n9499), .ZN(n10280) );
  NAND2_X1 U11877 ( .A1(n9848), .A2(n10280), .ZN(n10281) );
  NAND2_X1 U11878 ( .A1(n10281), .A2(n12639), .ZN(n9277) );
  OR2_X1 U11879 ( .A1(n12586), .A2(n15094), .ZN(n9282) );
  INV_X1 U11880 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9279) );
  OAI22_X1 U11881 ( .A1(n12589), .A2(n12585), .B1(n15096), .B2(n9279), .ZN(
        n9280) );
  NAND2_X1 U11882 ( .A1(n9282), .A2(n9281), .ZN(P3_U3487) );
  OAI22_X1 U11883 ( .A1(n15205), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n13448), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9290) );
  INV_X1 U11884 ( .A(n9290), .ZN(n9286) );
  XNOR2_X1 U11885 ( .A(n9291), .B(n9286), .ZN(n11877) );
  NAND2_X1 U11886 ( .A1(n11877), .A2(n9143), .ZN(n9288) );
  INV_X1 U11887 ( .A(SI_29_), .ZN(n11878) );
  OR2_X1 U11888 ( .A1(n9295), .A2(n11878), .ZN(n9287) );
  INV_X1 U11889 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11928) );
  INV_X1 U11890 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n11930) );
  NOR2_X1 U11891 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n11930), .ZN(n9292) );
  INV_X1 U11892 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13443) );
  INV_X1 U11893 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9293) );
  AOI22_X1 U11894 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n13443), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n9293), .ZN(n9294) );
  NAND2_X1 U11895 ( .A1(n12647), .A2(n9143), .ZN(n9297) );
  INV_X1 U11896 ( .A(SI_31_), .ZN(n12642) );
  OR2_X1 U11897 ( .A1(n9295), .A2(n12642), .ZN(n9296) );
  INV_X1 U11898 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14366) );
  NAND2_X1 U11899 ( .A1(n8893), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U11900 ( .A1(n9306), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n9298) );
  OAI211_X1 U11901 ( .C1(n14366), .C2(n9309), .A(n9299), .B(n9298), .ZN(n9300)
         );
  INV_X1 U11902 ( .A(n9300), .ZN(n9301) );
  NOR2_X1 U11903 ( .A1(n9315), .A2(n14332), .ZN(n9488) );
  AOI22_X1 U11904 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n11928), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n11930), .ZN(n9302) );
  INV_X1 U11905 ( .A(SI_30_), .ZN(n11882) );
  OR2_X1 U11906 ( .A1(n9295), .A2(n11882), .ZN(n9304) );
  INV_X1 U11907 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14368) );
  NAND2_X1 U11908 ( .A1(n8893), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n9308) );
  NAND2_X1 U11909 ( .A1(n9306), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n9307) );
  OAI211_X1 U11910 ( .C1(n14368), .C2(n9309), .A(n9308), .B(n9307), .ZN(n9310)
         );
  INV_X1 U11911 ( .A(n9310), .ZN(n9311) );
  AND2_X1 U11912 ( .A1(n9312), .A2(n9311), .ZN(n10705) );
  AND2_X1 U11913 ( .A1(n14355), .A2(n10705), .ZN(n9486) );
  AOI21_X1 U11914 ( .B1(n14355), .B2(n14332), .A(n9336), .ZN(n9314) );
  NAND2_X1 U11915 ( .A1(n9315), .A2(n14332), .ZN(n9319) );
  OR2_X1 U11916 ( .A1(n14355), .A2(n10705), .ZN(n9485) );
  INV_X1 U11917 ( .A(n9319), .ZN(n9489) );
  INV_X1 U11918 ( .A(n12444), .ZN(n9332) );
  INV_X1 U11919 ( .A(n12470), .ZN(n12464) );
  INV_X1 U11920 ( .A(n11806), .ZN(n9424) );
  NAND2_X1 U11921 ( .A1(n15033), .A2(n10311), .ZN(n9364) );
  INV_X1 U11922 ( .A(n9364), .ZN(n9321) );
  NOR2_X1 U11923 ( .A1(n9359), .A2(n9321), .ZN(n14913) );
  NAND3_X1 U11924 ( .A1(n14913), .A2(n9366), .A3(n15004), .ZN(n9324) );
  NAND4_X1 U11925 ( .A1(n15038), .A2(n10779), .A3(n11089), .A4(n14965), .ZN(
        n9323) );
  NOR2_X1 U11926 ( .A1(n9324), .A2(n9323), .ZN(n9326) );
  AND4_X1 U11927 ( .A1(n9326), .A2(n14981), .A3(n9325), .A4(n11198), .ZN(n9327) );
  NAND4_X1 U11928 ( .A1(n9327), .A2(n11456), .A3(n8967), .A4(n14339), .ZN(
        n9328) );
  NOR2_X1 U11929 ( .A1(n9328), .A2(n9418), .ZN(n9329) );
  NAND4_X1 U11930 ( .A1(n12485), .A2(n9424), .A3(n9329), .A4(n12501), .ZN(
        n9330) );
  OR3_X1 U11931 ( .A1(n12457), .A2(n12464), .A3(n9330), .ZN(n9331) );
  NOR4_X1 U11932 ( .A1(n12429), .A2(n9215), .A3(n9332), .A4(n9331), .ZN(n9333)
         );
  NAND4_X1 U11933 ( .A1(n12393), .A2(n12355), .A3(n12401), .A4(n9333), .ZN(
        n9334) );
  NOR4_X1 U11934 ( .A1(n12339), .A2(n12362), .A3(n9334), .A4(n12376), .ZN(
        n9335) );
  INV_X1 U11935 ( .A(n9336), .ZN(n9479) );
  NAND2_X1 U11936 ( .A1(n10881), .A2(n9338), .ZN(n9769) );
  MUX2_X1 U11937 ( .A(n9343), .B(n9342), .S(n9499), .Z(n9478) );
  NAND2_X1 U11938 ( .A1(n12340), .A2(n9499), .ZN(n9469) );
  INV_X1 U11939 ( .A(n9344), .ZN(n9346) );
  NOR2_X1 U11940 ( .A1(n12072), .A2(n12352), .ZN(n9345) );
  MUX2_X1 U11941 ( .A(n9346), .B(n9345), .S(n9499), .Z(n9347) );
  INV_X1 U11942 ( .A(n9347), .ZN(n9467) );
  MUX2_X1 U11943 ( .A(n9349), .B(n9348), .S(n9499), .Z(n9465) );
  MUX2_X1 U11944 ( .A(n9351), .B(n9350), .S(n10389), .Z(n9463) );
  MUX2_X1 U11945 ( .A(n9353), .B(n9352), .S(n9499), .Z(n9461) );
  INV_X1 U11946 ( .A(n9354), .ZN(n9357) );
  INV_X1 U11947 ( .A(n9355), .ZN(n9356) );
  MUX2_X1 U11948 ( .A(n9357), .B(n9356), .S(n9499), .Z(n9358) );
  INV_X1 U11949 ( .A(n9358), .ZN(n9459) );
  INV_X1 U11950 ( .A(n9359), .ZN(n15032) );
  NAND2_X1 U11951 ( .A1(n9360), .A2(n9364), .ZN(n9363) );
  INV_X1 U11952 ( .A(n9361), .ZN(n9362) );
  NAND3_X1 U11953 ( .A1(n15038), .A2(n10389), .A3(n9364), .ZN(n9365) );
  NAND3_X1 U11954 ( .A1(n9367), .A2(n9366), .A3(n9365), .ZN(n9371) );
  NAND2_X1 U11955 ( .A1(n9376), .A2(n9368), .ZN(n9369) );
  NAND2_X1 U11956 ( .A1(n9369), .A2(n9499), .ZN(n9370) );
  NAND2_X1 U11957 ( .A1(n9371), .A2(n9370), .ZN(n9375) );
  AOI21_X1 U11958 ( .B1(n9372), .B2(n9373), .A(n9499), .ZN(n9374) );
  AOI21_X1 U11959 ( .B1(n9375), .B2(n9372), .A(n9374), .ZN(n9381) );
  OAI21_X1 U11960 ( .B1(n9499), .B2(n9376), .A(n15004), .ZN(n9380) );
  MUX2_X1 U11961 ( .A(n9378), .B(n9377), .S(n9499), .Z(n9379) );
  OAI211_X1 U11962 ( .C1(n9381), .C2(n9380), .A(n14981), .B(n9379), .ZN(n9385)
         );
  NAND2_X1 U11963 ( .A1(n9391), .A2(n9382), .ZN(n9383) );
  NAND2_X1 U11964 ( .A1(n9383), .A2(n10389), .ZN(n9384) );
  NAND2_X1 U11965 ( .A1(n9385), .A2(n9384), .ZN(n9390) );
  NAND2_X1 U11966 ( .A1(n12188), .A2(n9386), .ZN(n9387) );
  AOI21_X1 U11967 ( .B1(n9389), .B2(n9387), .A(n10389), .ZN(n9388) );
  AOI21_X1 U11968 ( .B1(n9390), .B2(n9389), .A(n9388), .ZN(n9396) );
  OAI21_X1 U11969 ( .B1(n10389), .B2(n9391), .A(n14965), .ZN(n9395) );
  MUX2_X1 U11970 ( .A(n9393), .B(n9392), .S(n9499), .Z(n9394) );
  NAND2_X1 U11971 ( .A1(n11315), .A2(n9499), .ZN(n9398) );
  OR2_X1 U11972 ( .A1(n11315), .A2(n9499), .ZN(n9397) );
  MUX2_X1 U11973 ( .A(n9398), .B(n9397), .S(n14968), .Z(n9399) );
  NAND3_X1 U11974 ( .A1(n9400), .A2(n11456), .A3(n9399), .ZN(n9405) );
  INV_X1 U11975 ( .A(n9401), .ZN(n9403) );
  MUX2_X1 U11976 ( .A(n9403), .B(n9402), .S(n9499), .Z(n9404) );
  AOI21_X1 U11977 ( .B1(n9405), .B2(n9404), .A(n11410), .ZN(n9412) );
  MUX2_X1 U11978 ( .A(n9407), .B(n9406), .S(n9499), .Z(n9408) );
  NAND2_X1 U11979 ( .A1(n9408), .A2(n8967), .ZN(n9411) );
  AND2_X1 U11980 ( .A1(n9417), .A2(n9409), .ZN(n9410) );
  AOI21_X1 U11981 ( .B1(n9415), .B2(n9413), .A(n9499), .ZN(n9414) );
  AOI21_X1 U11982 ( .B1(n9416), .B2(n9415), .A(n9414), .ZN(n9420) );
  NOR2_X1 U11983 ( .A1(n9417), .A2(n9499), .ZN(n9419) );
  MUX2_X1 U11984 ( .A(n9422), .B(n9421), .S(n9499), .Z(n9423) );
  NAND4_X1 U11985 ( .A1(n9425), .A2(n9424), .A3(n12501), .A4(n9423), .ZN(n9432) );
  INV_X1 U11986 ( .A(n9426), .ZN(n9427) );
  NAND2_X1 U11987 ( .A1(n12501), .A2(n9427), .ZN(n9428) );
  OAI211_X1 U11988 ( .C1(n9801), .C2(n12166), .A(n9428), .B(n9437), .ZN(n9429)
         );
  NAND2_X1 U11989 ( .A1(n9429), .A2(n9499), .ZN(n9431) );
  INV_X1 U11990 ( .A(n9434), .ZN(n9430) );
  AOI21_X1 U11991 ( .B1(n9432), .B2(n9431), .A(n9430), .ZN(n9439) );
  OAI211_X1 U11992 ( .C1(n12495), .C2(n9435), .A(n9434), .B(n9433), .ZN(n9436)
         );
  AND2_X1 U11993 ( .A1(n9436), .A2(n10389), .ZN(n9438) );
  OAI22_X1 U11994 ( .A1(n9439), .A2(n9438), .B1(n9499), .B2(n9437), .ZN(n9442)
         );
  NAND2_X1 U11995 ( .A1(n12618), .A2(n12452), .ZN(n9448) );
  OAI21_X1 U11996 ( .B1(n12088), .B2(n12095), .A(n12442), .ZN(n9440) );
  NAND2_X1 U11997 ( .A1(n9440), .A2(n9443), .ZN(n9441) );
  NAND3_X1 U11998 ( .A1(n9448), .A2(n10389), .A3(n9441), .ZN(n9445) );
  AOI22_X1 U11999 ( .A1(n9442), .A2(n12470), .B1(n9445), .B2(n6547), .ZN(n9447) );
  NAND3_X1 U12000 ( .A1(n9449), .A2(n9499), .A3(n9443), .ZN(n9444) );
  NAND2_X1 U12001 ( .A1(n9445), .A2(n9444), .ZN(n9446) );
  OAI21_X1 U12002 ( .B1(n9447), .B2(n12457), .A(n9446), .ZN(n9454) );
  INV_X1 U12003 ( .A(n9448), .ZN(n9451) );
  INV_X1 U12004 ( .A(n9449), .ZN(n9450) );
  MUX2_X1 U12005 ( .A(n9451), .B(n9450), .S(n10389), .Z(n9452) );
  INV_X1 U12006 ( .A(n9452), .ZN(n9453) );
  NAND3_X1 U12007 ( .A1(n9454), .A2(n9096), .A3(n9453), .ZN(n9457) );
  NAND3_X1 U12008 ( .A1(n12115), .A2(n12441), .A3(n9499), .ZN(n9456) );
  NAND3_X1 U12009 ( .A1(n12614), .A2(n10389), .A3(n12182), .ZN(n9455) );
  NAND4_X1 U12010 ( .A1(n12417), .A2(n9457), .A3(n9456), .A4(n9455), .ZN(n9458) );
  NAND3_X1 U12011 ( .A1(n12401), .A2(n9459), .A3(n9458), .ZN(n9460) );
  NAND3_X1 U12012 ( .A1(n9461), .A2(n9460), .A3(n12393), .ZN(n9462) );
  NAND3_X1 U12013 ( .A1(n9140), .A2(n9463), .A3(n9462), .ZN(n9464) );
  NAND3_X1 U12014 ( .A1(n12368), .A2(n9465), .A3(n9464), .ZN(n9466) );
  OAI21_X1 U12015 ( .B1(n9469), .B2(n12155), .A(n9468), .ZN(n9471) );
  NOR2_X1 U12016 ( .A1(n12179), .A2(n9499), .ZN(n9470) );
  NAND2_X1 U12017 ( .A1(n9473), .A2(n9472), .ZN(n9474) );
  MUX2_X1 U12018 ( .A(n9474), .B(n9473), .S(n9499), .Z(n9475) );
  NAND3_X1 U12019 ( .A1(n11952), .A2(n9476), .A3(n9475), .ZN(n9477) );
  INV_X1 U12020 ( .A(n9482), .ZN(n9480) );
  NAND2_X1 U12021 ( .A1(n9480), .A2(n9479), .ZN(n9484) );
  NOR2_X1 U12022 ( .A1(n9482), .A2(n9481), .ZN(n9483) );
  OAI21_X1 U12023 ( .B1(n9487), .B2(n9486), .A(n9485), .ZN(n9491) );
  INV_X1 U12024 ( .A(n9488), .ZN(n9490) );
  AOI21_X1 U12025 ( .B1(n9491), .B2(n9490), .A(n9489), .ZN(n9493) );
  INV_X1 U12026 ( .A(n10388), .ZN(n9495) );
  NAND2_X1 U12027 ( .A1(n9495), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11320) );
  INV_X1 U12028 ( .A(n11320), .ZN(n9496) );
  OAI21_X1 U12029 ( .B1(n9498), .B2(n9497), .A(n9496), .ZN(n9503) );
  OR2_X1 U12030 ( .A1(n9500), .A2(n9499), .ZN(n10276) );
  INV_X1 U12031 ( .A(n11876), .ZN(n10393) );
  NAND3_X1 U12032 ( .A1(n9855), .A2(n10393), .A3(n12198), .ZN(n9501) );
  OAI211_X1 U12033 ( .C1(n11033), .C2(n11320), .A(n9501), .B(P3_B_REG_SCAN_IN), 
        .ZN(n9502) );
  NAND2_X1 U12034 ( .A1(n9503), .A2(n9502), .ZN(P3_U3296) );
  NAND2_X1 U12035 ( .A1(n9506), .A2(n9507), .ZN(n9508) );
  AND2_X2 U12036 ( .A1(n9663), .A2(n9508), .ZN(n9541) );
  INV_X4 U12037 ( .A(n9541), .ZN(n9680) );
  MUX2_X1 U12038 ( .A(n14388), .B(n11733), .S(n9680), .Z(n9573) );
  INV_X1 U12039 ( .A(n10019), .ZN(n9677) );
  NAND2_X1 U12040 ( .A1(n9685), .A2(n9677), .ZN(n9511) );
  NAND2_X1 U12041 ( .A1(n9512), .A2(n9541), .ZN(n9515) );
  NAND2_X1 U12042 ( .A1(n9680), .A2(n9513), .ZN(n9514) );
  NAND2_X1 U12043 ( .A1(n9541), .A2(n10167), .ZN(n9517) );
  NAND2_X1 U12044 ( .A1(n9680), .A2(n14652), .ZN(n9516) );
  INV_X1 U12045 ( .A(n9520), .ZN(n9522) );
  MUX2_X1 U12046 ( .A(n9525), .B(n9524), .S(n9680), .Z(n9526) );
  MUX2_X1 U12047 ( .A(n14670), .B(n10871), .S(n9680), .Z(n9528) );
  INV_X1 U12048 ( .A(n10871), .ZN(n13778) );
  MUX2_X1 U12049 ( .A(n13778), .B(n10876), .S(n9680), .Z(n9527) );
  NAND2_X1 U12050 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  NAND2_X1 U12051 ( .A1(n9531), .A2(n9530), .ZN(n9535) );
  MUX2_X1 U12052 ( .A(n13777), .B(n10901), .S(n9680), .Z(n9534) );
  MUX2_X1 U12053 ( .A(n10901), .B(n13777), .S(n9680), .Z(n9532) );
  INV_X1 U12054 ( .A(n9680), .ZN(n9555) );
  MUX2_X1 U12055 ( .A(n13776), .B(n13723), .S(n9555), .Z(n9538) );
  MUX2_X1 U12056 ( .A(n13776), .B(n13723), .S(n9680), .Z(n9536) );
  MUX2_X1 U12057 ( .A(n13775), .B(n11029), .S(n9680), .Z(n9540) );
  MUX2_X1 U12058 ( .A(n13775), .B(n11029), .S(n9541), .Z(n9539) );
  MUX2_X1 U12059 ( .A(n13774), .B(n11257), .S(n9541), .Z(n9545) );
  NAND2_X1 U12060 ( .A1(n9544), .A2(n9545), .ZN(n9543) );
  MUX2_X1 U12061 ( .A(n13774), .B(n11257), .S(n9680), .Z(n9542) );
  NAND2_X1 U12062 ( .A1(n9543), .A2(n9542), .ZN(n9549) );
  INV_X1 U12063 ( .A(n9544), .ZN(n9547) );
  INV_X1 U12064 ( .A(n9545), .ZN(n9546) );
  NAND2_X1 U12065 ( .A1(n9547), .A2(n9546), .ZN(n9548) );
  MUX2_X1 U12066 ( .A(n13773), .B(n14705), .S(n9680), .Z(n9553) );
  INV_X1 U12067 ( .A(n9680), .ZN(n9550) );
  MUX2_X1 U12068 ( .A(n13773), .B(n14705), .S(n9550), .Z(n9551) );
  INV_X1 U12069 ( .A(n9553), .ZN(n9554) );
  MUX2_X1 U12070 ( .A(n13772), .B(n11381), .S(n9555), .Z(n9557) );
  MUX2_X1 U12071 ( .A(n13772), .B(n11381), .S(n9680), .Z(n9556) );
  NAND2_X1 U12072 ( .A1(n9559), .A2(n9558), .ZN(n9561) );
  MUX2_X1 U12073 ( .A(n13771), .B(n14453), .S(n9680), .Z(n9562) );
  MUX2_X1 U12074 ( .A(n13771), .B(n14453), .S(n9550), .Z(n9560) );
  MUX2_X1 U12075 ( .A(n13770), .B(n11678), .S(n9550), .Z(n9566) );
  MUX2_X1 U12076 ( .A(n13770), .B(n11678), .S(n9680), .Z(n9563) );
  NAND2_X1 U12077 ( .A1(n9564), .A2(n9563), .ZN(n9570) );
  INV_X1 U12078 ( .A(n9565), .ZN(n9568) );
  INV_X1 U12079 ( .A(n9566), .ZN(n9567) );
  NAND2_X1 U12080 ( .A1(n9568), .A2(n9567), .ZN(n9569) );
  NAND2_X1 U12081 ( .A1(n9570), .A2(n9569), .ZN(n9572) );
  MUX2_X1 U12082 ( .A(n14388), .B(n11733), .S(n9550), .Z(n9571) );
  NAND2_X1 U12083 ( .A1(n9581), .A2(n9574), .ZN(n9577) );
  NAND2_X1 U12084 ( .A1(n9582), .A2(n9575), .ZN(n9576) );
  MUX2_X1 U12085 ( .A(n9577), .B(n9576), .S(n9680), .Z(n9578) );
  NAND2_X1 U12086 ( .A1(n9580), .A2(n9579), .ZN(n9587) );
  INV_X1 U12087 ( .A(n9581), .ZN(n9584) );
  INV_X1 U12088 ( .A(n9582), .ZN(n9583) );
  MUX2_X1 U12089 ( .A(n9584), .B(n9583), .S(n9550), .Z(n9585) );
  NAND2_X1 U12090 ( .A1(n9587), .A2(n9586), .ZN(n9591) );
  MUX2_X1 U12091 ( .A(n13767), .B(n14430), .S(n9680), .Z(n9590) );
  INV_X1 U12092 ( .A(n14430), .ZN(n9588) );
  MUX2_X1 U12093 ( .A(n11823), .B(n9588), .S(n9550), .Z(n9589) );
  MUX2_X1 U12094 ( .A(n7279), .B(n8678), .S(n9550), .Z(n9592) );
  OAI21_X1 U12095 ( .B1(n9594), .B2(n9683), .A(n9593), .ZN(n9599) );
  OAI21_X1 U12096 ( .B1(n14044), .B2(n13765), .A(n9600), .ZN(n9597) );
  NAND2_X1 U12097 ( .A1(n9601), .A2(n9595), .ZN(n9596) );
  MUX2_X1 U12098 ( .A(n9597), .B(n9596), .S(n9550), .Z(n9598) );
  INV_X1 U12099 ( .A(n9600), .ZN(n9603) );
  INV_X1 U12100 ( .A(n9601), .ZN(n9602) );
  MUX2_X1 U12101 ( .A(n9603), .B(n9602), .S(n9680), .Z(n9604) );
  MUX2_X1 U12102 ( .A(n14113), .B(n13763), .S(n9550), .Z(n9605) );
  INV_X1 U12103 ( .A(n9605), .ZN(n9607) );
  MUX2_X1 U12104 ( .A(n14113), .B(n13763), .S(n9680), .Z(n9606) );
  MUX2_X1 U12105 ( .A(n13762), .B(n14108), .S(n9550), .Z(n9610) );
  MUX2_X1 U12106 ( .A(n14108), .B(n13762), .S(n9550), .Z(n9608) );
  NAND2_X1 U12107 ( .A1(n9609), .A2(n9608), .ZN(n9614) );
  INV_X1 U12108 ( .A(n9610), .ZN(n9611) );
  NAND2_X1 U12109 ( .A1(n9612), .A2(n9611), .ZN(n9613) );
  MUX2_X1 U12110 ( .A(n14101), .B(n13642), .S(n9550), .Z(n9617) );
  MUX2_X1 U12111 ( .A(n13642), .B(n14101), .S(n9550), .Z(n9615) );
  MUX2_X1 U12112 ( .A(n13760), .B(n14093), .S(n9550), .Z(n9619) );
  MUX2_X1 U12113 ( .A(n14093), .B(n13760), .S(n9550), .Z(n9618) );
  INV_X1 U12114 ( .A(n9619), .ZN(n9620) );
  MUX2_X1 U12115 ( .A(n14087), .B(n13759), .S(n9555), .Z(n9624) );
  NAND2_X1 U12116 ( .A1(n9623), .A2(n9624), .ZN(n9622) );
  MUX2_X1 U12117 ( .A(n13759), .B(n14087), .S(n9550), .Z(n9621) );
  NAND2_X1 U12118 ( .A1(n9622), .A2(n9621), .ZN(n9628) );
  INV_X1 U12119 ( .A(n9623), .ZN(n9626) );
  INV_X1 U12120 ( .A(n9624), .ZN(n9625) );
  NAND2_X1 U12121 ( .A1(n9626), .A2(n9625), .ZN(n9627) );
  MUX2_X1 U12122 ( .A(n13758), .B(n14082), .S(n9550), .Z(n9630) );
  MUX2_X1 U12123 ( .A(n13758), .B(n14082), .S(n9680), .Z(n9629) );
  INV_X1 U12124 ( .A(n9630), .ZN(n9631) );
  MUX2_X1 U12125 ( .A(n13757), .B(n13915), .S(n9680), .Z(n9634) );
  MUX2_X1 U12126 ( .A(n13757), .B(n13915), .S(n9555), .Z(n9632) );
  MUX2_X1 U12127 ( .A(n14066), .B(n13756), .S(n9680), .Z(n9638) );
  MUX2_X1 U12128 ( .A(n14066), .B(n13756), .S(n9550), .Z(n9635) );
  NAND2_X1 U12129 ( .A1(n9636), .A2(n9635), .ZN(n9642) );
  INV_X1 U12130 ( .A(n9637), .ZN(n9640) );
  INV_X1 U12131 ( .A(n9638), .ZN(n9639) );
  NAND2_X1 U12132 ( .A1(n9640), .A2(n9639), .ZN(n9641) );
  MUX2_X1 U12133 ( .A(n13755), .B(n14061), .S(n9680), .Z(n9643) );
  MUX2_X1 U12134 ( .A(n13755), .B(n14061), .S(n9550), .Z(n9644) );
  MUX2_X1 U12135 ( .A(n13635), .B(n14054), .S(n9555), .Z(n9647) );
  MUX2_X1 U12136 ( .A(n9645), .B(n13754), .S(n9550), .Z(n9646) );
  NAND2_X1 U12137 ( .A1(n9650), .A2(n11878), .ZN(n9651) );
  MUX2_X1 U12138 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7524), .Z(n9652) );
  NAND2_X1 U12139 ( .A1(n9652), .A2(SI_30_), .ZN(n9670) );
  OAI21_X1 U12140 ( .B1(n9652), .B2(SI_30_), .A(n9670), .ZN(n9653) );
  NAND2_X1 U12141 ( .A1(n9654), .A2(n9653), .ZN(n9655) );
  NAND2_X1 U12142 ( .A1(n12783), .A2(n9656), .ZN(n9658) );
  NAND2_X1 U12143 ( .A1(n9674), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9657) );
  INV_X1 U12144 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9662) );
  NAND2_X1 U12145 ( .A1(n9659), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9661) );
  OAI211_X1 U12146 ( .C1(n8304), .C2(n9662), .A(n9661), .B(n9660), .ZN(n13864)
         );
  OAI21_X1 U12147 ( .B1(n13864), .B2(n7461), .A(n13753), .ZN(n9664) );
  INV_X1 U12148 ( .A(n9664), .ZN(n9665) );
  MUX2_X1 U12149 ( .A(n13870), .B(n9665), .S(n9680), .Z(n9708) );
  INV_X1 U12150 ( .A(n13864), .ZN(n9667) );
  INV_X1 U12151 ( .A(n9506), .ZN(n9666) );
  OAI22_X1 U12152 ( .A1(n9680), .A2(n9667), .B1(n10011), .B2(n9666), .ZN(n9668) );
  AND2_X1 U12153 ( .A1(n9668), .A2(n13753), .ZN(n9669) );
  AOI21_X1 U12154 ( .B1(n13870), .B2(n9680), .A(n9669), .ZN(n9707) );
  NOR2_X1 U12155 ( .A1(n9708), .A2(n9707), .ZN(n9710) );
  MUX2_X1 U12156 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9926), .Z(n9672) );
  XNOR2_X1 U12157 ( .A(n9672), .B(SI_31_), .ZN(n9673) );
  NAND2_X1 U12158 ( .A1(n13440), .A2(n9656), .ZN(n9676) );
  NAND2_X1 U12159 ( .A1(n9674), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9675) );
  NAND2_X1 U12160 ( .A1(n9680), .A2(n13864), .ZN(n9712) );
  NAND2_X1 U12161 ( .A1(n10014), .A2(n10201), .ZN(n9678) );
  NAND2_X1 U12162 ( .A1(n9677), .A2(n14023), .ZN(n10825) );
  AND2_X1 U12163 ( .A1(n9678), .A2(n10825), .ZN(n9719) );
  INV_X1 U12164 ( .A(n9719), .ZN(n9679) );
  AND2_X1 U12165 ( .A1(n9679), .A2(n9704), .ZN(n9715) );
  NOR2_X1 U12166 ( .A1(n9680), .A2(n13864), .ZN(n9714) );
  NAND2_X1 U12167 ( .A1(n13866), .A2(n9714), .ZN(n9681) );
  OAI211_X1 U12168 ( .C1(n13866), .C2(n9712), .A(n9715), .B(n9681), .ZN(n9726)
         );
  INV_X1 U12169 ( .A(n9682), .ZN(n9684) );
  NAND2_X1 U12170 ( .A1(n9684), .A2(n9683), .ZN(n11821) );
  NAND4_X1 U12171 ( .A1(n10375), .A2(n14624), .A3(n9685), .A4(n9686), .ZN(
        n9687) );
  NOR2_X1 U12172 ( .A1(n9687), .A2(n10851), .ZN(n9689) );
  NAND4_X1 U12173 ( .A1(n10751), .A2(n9689), .A3(n9688), .A4(n10819), .ZN(
        n9690) );
  NOR2_X1 U12174 ( .A1(n10691), .A2(n9690), .ZN(n9691) );
  NAND4_X1 U12175 ( .A1(n11214), .A2(n9692), .A3(n9691), .A4(n10932), .ZN(
        n9693) );
  NOR3_X1 U12176 ( .A1(n9694), .A2(n11349), .A3(n9693), .ZN(n9696) );
  NAND4_X1 U12177 ( .A1(n11821), .A2(n9696), .A3(n14413), .A4(n9695), .ZN(
        n9698) );
  NOR2_X1 U12178 ( .A1(n9698), .A2(n9697), .ZN(n9699) );
  AND4_X1 U12179 ( .A1(n13985), .A2(n14017), .A3(n9699), .A4(n14034), .ZN(
        n9700) );
  NAND4_X1 U12180 ( .A1(n13967), .A2(n13970), .A3(n9700), .A4(n13996), .ZN(
        n9701) );
  NOR4_X1 U12181 ( .A1(n13912), .A2(n13927), .A3(n13942), .A4(n9701), .ZN(
        n9702) );
  INV_X1 U12182 ( .A(n9704), .ZN(n9705) );
  NAND2_X1 U12183 ( .A1(n9706), .A2(n9705), .ZN(n9729) );
  AND2_X1 U12184 ( .A1(n9708), .A2(n9707), .ZN(n9730) );
  INV_X1 U12185 ( .A(n9730), .ZN(n9725) );
  NAND2_X1 U12186 ( .A1(n9709), .A2(n9719), .ZN(n9731) );
  INV_X1 U12187 ( .A(n9731), .ZN(n9711) );
  NAND2_X1 U12188 ( .A1(n9711), .A2(n9710), .ZN(n9724) );
  AND2_X1 U12189 ( .A1(n9715), .A2(n13864), .ZN(n9713) );
  MUX2_X1 U12190 ( .A(n9719), .B(n9713), .S(n9712), .Z(n9722) );
  INV_X1 U12191 ( .A(n9714), .ZN(n9718) );
  INV_X1 U12192 ( .A(n9715), .ZN(n9716) );
  OAI21_X1 U12193 ( .B1(n13864), .B2(n9716), .A(n9718), .ZN(n9717) );
  OAI21_X1 U12194 ( .B1(n9719), .B2(n9718), .A(n9717), .ZN(n9720) );
  NAND2_X1 U12195 ( .A1(n13866), .A2(n9720), .ZN(n9721) );
  OAI21_X1 U12196 ( .B1(n13866), .B2(n9722), .A(n9721), .ZN(n9723) );
  OAI211_X1 U12197 ( .C1(n9726), .C2(n9725), .A(n9724), .B(n9723), .ZN(n9727)
         );
  NOR2_X1 U12198 ( .A1(n9731), .A2(n9730), .ZN(n9732) );
  NAND2_X1 U12199 ( .A1(n9733), .A2(n9732), .ZN(n9734) );
  NAND3_X1 U12200 ( .A1(n9735), .A2(n7506), .A3(n9734), .ZN(n9738) );
  INV_X1 U12201 ( .A(n9922), .ZN(n9736) );
  NAND2_X1 U12202 ( .A1(n9736), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11817) );
  NAND2_X1 U12203 ( .A1(n9738), .A2(n9737), .ZN(n9742) );
  NOR3_X1 U12204 ( .A1(n10193), .A2(n6459), .A3(n14633), .ZN(n9740) );
  OAI21_X1 U12205 ( .B1(n11817), .B2(n9504), .A(P1_B_REG_SCAN_IN), .ZN(n9739)
         );
  OR2_X1 U12206 ( .A1(n9740), .A2(n9739), .ZN(n9741) );
  NAND2_X1 U12207 ( .A1(n9742), .A2(n9741), .ZN(P1_U3242) );
  INV_X1 U12208 ( .A(n9748), .ZN(n12341) );
  NAND2_X1 U12209 ( .A1(n11963), .A2(n12341), .ZN(n9743) );
  NAND2_X1 U12210 ( .A1(n9744), .A2(n9743), .ZN(n9746) );
  XNOR2_X1 U12211 ( .A(n9746), .B(n9745), .ZN(n9750) );
  NAND2_X1 U12212 ( .A1(n10393), .A2(P3_B_REG_SCAN_IN), .ZN(n9747) );
  NAND2_X1 U12213 ( .A1(n15035), .A2(n9747), .ZN(n14331) );
  OAI22_X1 U12214 ( .A1(n9748), .A2(n15019), .B1(n10705), .B2(n14331), .ZN(
        n9749) );
  AOI21_X2 U12215 ( .B1(n9750), .B2(n15039), .A(n9749), .ZN(n12018) );
  XNOR2_X1 U12216 ( .A(n9752), .B(n9751), .ZN(n12022) );
  NAND2_X1 U12217 ( .A1(n12022), .A2(n14362), .ZN(n9753) );
  NAND2_X1 U12218 ( .A1(n12018), .A2(n9753), .ZN(n9764) );
  OR2_X1 U12219 ( .A1(n9754), .A2(n9769), .ZN(n9846) );
  NOR2_X1 U12220 ( .A1(n9846), .A2(n10387), .ZN(n9755) );
  OR2_X1 U12221 ( .A1(n9855), .A2(n9755), .ZN(n9757) );
  INV_X1 U12222 ( .A(n9756), .ZN(n9758) );
  NAND2_X1 U12223 ( .A1(n9757), .A2(n9850), .ZN(n9760) );
  INV_X1 U12224 ( .A(n10387), .ZN(n9840) );
  NAND3_X1 U12225 ( .A1(n9854), .A2(n9840), .A3(n9847), .ZN(n9759) );
  OR2_X1 U12226 ( .A1(n9764), .A2(n15080), .ZN(n9762) );
  NAND2_X1 U12227 ( .A1(n15080), .A2(n9234), .ZN(n9761) );
  NAND2_X1 U12228 ( .A1(n9762), .A2(n9761), .ZN(n9763) );
  OR2_X1 U12229 ( .A1(n15080), .A2(n15030), .ZN(n12638) );
  NAND2_X1 U12230 ( .A1(n9763), .A2(n7504), .ZN(P3_U3456) );
  OR2_X1 U12231 ( .A1(n9764), .A2(n15094), .ZN(n9765) );
  NAND2_X1 U12232 ( .A1(n9765), .A2(n6610), .ZN(n9766) );
  NAND2_X1 U12233 ( .A1(n9766), .A2(n7505), .ZN(P3_U3488) );
  NAND2_X1 U12234 ( .A1(n9767), .A2(n10881), .ZN(n9768) );
  XNOR2_X1 U12235 ( .A(n12523), .B(n11951), .ZN(n11959) );
  NOR2_X1 U12236 ( .A1(n11959), .A2(n12179), .ZN(n11954) );
  XNOR2_X1 U12237 ( .A(n12559), .B(n10315), .ZN(n9808) );
  XNOR2_X1 U12238 ( .A(n14957), .B(n10315), .ZN(n9787) );
  INV_X1 U12239 ( .A(n9787), .ZN(n9788) );
  INV_X1 U12240 ( .A(n12186), .ZN(n11312) );
  XNOR2_X1 U12241 ( .A(n14999), .B(n10315), .ZN(n9778) );
  XNOR2_X1 U12242 ( .A(n10655), .B(n10315), .ZN(n9776) );
  INV_X1 U12243 ( .A(n9776), .ZN(n9777) );
  OAI21_X1 U12244 ( .B1(n15037), .B2(n10315), .A(n9771), .ZN(n9772) );
  NAND2_X1 U12245 ( .A1(n9772), .A2(n10318), .ZN(n10317) );
  INV_X1 U12246 ( .A(n9773), .ZN(n9774) );
  NAND2_X1 U12247 ( .A1(n10317), .A2(n9774), .ZN(n10364) );
  XNOR2_X1 U12248 ( .A(n9776), .B(n15018), .ZN(n10651) );
  XNOR2_X1 U12249 ( .A(n12189), .B(n9778), .ZN(n10743) );
  XNOR2_X1 U12250 ( .A(n14994), .B(n10315), .ZN(n9779) );
  XNOR2_X1 U12251 ( .A(n9779), .B(n12188), .ZN(n10915) );
  XNOR2_X1 U12252 ( .A(n10952), .B(n10315), .ZN(n9780) );
  XNOR2_X1 U12253 ( .A(n14969), .B(n9780), .ZN(n10947) );
  INV_X1 U12254 ( .A(n9780), .ZN(n9781) );
  NAND2_X1 U12255 ( .A1(n9781), .A2(n14969), .ZN(n9782) );
  NAND2_X1 U12256 ( .A1(n10946), .A2(n9782), .ZN(n11148) );
  XNOR2_X1 U12257 ( .A(n14965), .B(n10315), .ZN(n11147) );
  XNOR2_X1 U12258 ( .A(n11315), .B(n10315), .ZN(n9784) );
  XNOR2_X1 U12259 ( .A(n9784), .B(n14968), .ZN(n11309) );
  XNOR2_X1 U12260 ( .A(n9787), .B(n12186), .ZN(n11485) );
  XNOR2_X1 U12261 ( .A(n9789), .B(n10315), .ZN(n9790) );
  XNOR2_X1 U12262 ( .A(n12185), .B(n9790), .ZN(n11663) );
  XOR2_X1 U12263 ( .A(n10315), .B(n14348), .Z(n12061) );
  XNOR2_X1 U12264 ( .A(n11505), .B(n10315), .ZN(n9793) );
  OAI22_X1 U12265 ( .A1(n12061), .A2(n12513), .B1(n14347), .B2(n9793), .ZN(
        n9796) );
  INV_X1 U12266 ( .A(n9793), .ZN(n12060) );
  OAI21_X1 U12267 ( .B1(n12060), .B2(n12184), .A(n12183), .ZN(n9792) );
  NAND2_X1 U12268 ( .A1(n12061), .A2(n9792), .ZN(n9795) );
  NAND3_X1 U12269 ( .A1(n9793), .A2(n12513), .A3(n14347), .ZN(n9794) );
  XNOR2_X1 U12270 ( .A(n12125), .B(n11951), .ZN(n12119) );
  NOR2_X1 U12271 ( .A1(n12119), .A2(n14344), .ZN(n9797) );
  XNOR2_X1 U12272 ( .A(n12031), .B(n10315), .ZN(n9798) );
  NAND2_X1 U12273 ( .A1(n9798), .A2(n12514), .ZN(n9799) );
  OAI21_X1 U12274 ( .B1(n9798), .B2(n12514), .A(n9799), .ZN(n12025) );
  XNOR2_X1 U12275 ( .A(n12166), .B(n10315), .ZN(n9800) );
  XNOR2_X1 U12276 ( .A(n9800), .B(n12482), .ZN(n12167) );
  XNOR2_X1 U12277 ( .A(n12567), .B(n10315), .ZN(n9802) );
  XNOR2_X1 U12278 ( .A(n9802), .B(n12500), .ZN(n12084) );
  NAND2_X1 U12279 ( .A1(n7502), .A2(n9803), .ZN(n12092) );
  XNOR2_X1 U12280 ( .A(n12095), .B(n10315), .ZN(n9804) );
  XNOR2_X1 U12281 ( .A(n9804), .B(n12481), .ZN(n12093) );
  NAND2_X1 U12282 ( .A1(n12092), .A2(n12093), .ZN(n9806) );
  NAND2_X1 U12283 ( .A1(n9806), .A2(n9805), .ZN(n12147) );
  XNOR2_X1 U12284 ( .A(n9808), .B(n12466), .ZN(n12148) );
  NAND2_X1 U12285 ( .A1(n12147), .A2(n12148), .ZN(n9807) );
  XNOR2_X1 U12286 ( .A(n12618), .B(n10315), .ZN(n9809) );
  XNOR2_X1 U12287 ( .A(n9809), .B(n12427), .ZN(n12043) );
  XNOR2_X1 U12288 ( .A(n12115), .B(n10315), .ZN(n9810) );
  XNOR2_X1 U12289 ( .A(n9810), .B(n12182), .ZN(n12110) );
  XNOR2_X1 U12290 ( .A(n12050), .B(n11951), .ZN(n9811) );
  NOR2_X1 U12291 ( .A1(n9811), .A2(n12181), .ZN(n9812) );
  AOI21_X1 U12292 ( .B1(n9811), .B2(n12181), .A(n9812), .ZN(n12052) );
  XNOR2_X1 U12293 ( .A(n12406), .B(n10315), .ZN(n9815) );
  INV_X1 U12294 ( .A(n9815), .ZN(n9813) );
  NAND2_X1 U12295 ( .A1(n9816), .A2(n9815), .ZN(n9818) );
  INV_X1 U12296 ( .A(n9823), .ZN(n9821) );
  XNOR2_X1 U12297 ( .A(n9819), .B(n10315), .ZN(n9822) );
  INV_X1 U12298 ( .A(n9822), .ZN(n9820) );
  NAND2_X1 U12299 ( .A1(n12035), .A2(n12100), .ZN(n9828) );
  XNOR2_X1 U12300 ( .A(n12602), .B(n11951), .ZN(n9825) );
  NAND2_X1 U12301 ( .A1(n9825), .A2(n12389), .ZN(n12074) );
  INV_X1 U12302 ( .A(n9825), .ZN(n9826) );
  NAND2_X1 U12303 ( .A1(n9826), .A2(n12364), .ZN(n9827) );
  NAND2_X1 U12304 ( .A1(n9828), .A2(n12101), .ZN(n12073) );
  NAND2_X1 U12305 ( .A1(n12073), .A2(n12074), .ZN(n9832) );
  XNOR2_X1 U12306 ( .A(n12072), .B(n10315), .ZN(n9829) );
  NAND2_X1 U12307 ( .A1(n9829), .A2(n12352), .ZN(n9833) );
  INV_X1 U12308 ( .A(n9829), .ZN(n9830) );
  NAND2_X1 U12309 ( .A1(n9830), .A2(n12379), .ZN(n9831) );
  NAND2_X1 U12310 ( .A1(n9832), .A2(n12075), .ZN(n12077) );
  NAND2_X1 U12311 ( .A1(n12077), .A2(n9833), .ZN(n12156) );
  XNOR2_X1 U12312 ( .A(n12155), .B(n11951), .ZN(n9834) );
  NOR2_X1 U12313 ( .A1(n9834), .A2(n12340), .ZN(n9835) );
  AOI21_X1 U12314 ( .B1(n9834), .B2(n12340), .A(n9835), .ZN(n12158) );
  INV_X1 U12315 ( .A(n9846), .ZN(n9837) );
  NAND2_X1 U12316 ( .A1(n9854), .A2(n9837), .ZN(n9839) );
  NAND3_X1 U12317 ( .A1(n9850), .A2(n9847), .A3(n15030), .ZN(n9838) );
  NAND2_X1 U12318 ( .A1(n9839), .A2(n9838), .ZN(n9841) );
  INV_X1 U12319 ( .A(n12523), .ZN(n12347) );
  INV_X1 U12320 ( .A(n9843), .ZN(n9842) );
  NAND2_X1 U12321 ( .A1(n9850), .A2(n9842), .ZN(n9844) );
  AND2_X1 U12322 ( .A1(n9854), .A2(n9855), .ZN(n9860) );
  INV_X1 U12323 ( .A(n12345), .ZN(n9862) );
  NOR2_X1 U12324 ( .A1(n9854), .A2(n9846), .ZN(n9852) );
  INV_X1 U12325 ( .A(n9847), .ZN(n9849) );
  OAI211_X1 U12326 ( .C1(n9850), .C2(n9849), .A(n9870), .B(n9848), .ZN(n9851)
         );
  OR2_X1 U12327 ( .A1(n9852), .A2(n9851), .ZN(n9853) );
  NAND2_X1 U12328 ( .A1(n9853), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9858) );
  INV_X1 U12329 ( .A(n9854), .ZN(n9856) );
  NAND2_X1 U12330 ( .A1(n9856), .A2(n9855), .ZN(n9857) );
  AND2_X1 U12331 ( .A1(n9858), .A2(n9857), .ZN(n10319) );
  AOI22_X1 U12332 ( .A1(n12340), .A2(n12170), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9861) );
  OAI21_X1 U12333 ( .B1(n9862), .B2(n12161), .A(n9861), .ZN(n9863) );
  AOI21_X1 U12334 ( .B1(n12341), .B2(n14916), .A(n9863), .ZN(n9864) );
  OAI21_X1 U12335 ( .B1(n12347), .B2(n12177), .A(n9864), .ZN(n9865) );
  INV_X1 U12336 ( .A(n9865), .ZN(n9866) );
  NAND2_X1 U12337 ( .A1(n9867), .A2(n9866), .ZN(P3_U3154) );
  INV_X1 U12338 ( .A(n9870), .ZN(n9871) );
  INV_X1 U12339 ( .A(n10023), .ZN(n10018) );
  INV_X1 U12340 ( .A(n9873), .ZN(n11985) );
  AOI211_X1 U12341 ( .C1(n9875), .C2(n9874), .A(n12759), .B(n11985), .ZN(n9880) );
  MUX2_X1 U12342 ( .A(P2_U3088), .B(n12770), .S(n10616), .Z(n9879) );
  INV_X1 U12343 ( .A(n14381), .ZN(n12776) );
  OR2_X1 U12344 ( .A1(n12773), .A2(n6635), .ZN(n9877) );
  NAND2_X1 U12345 ( .A1(n13036), .A2(n13069), .ZN(n9876) );
  AND2_X1 U12346 ( .A1(n9877), .A2(n9876), .ZN(n14853) );
  OAI22_X1 U12347 ( .A1(n12776), .A2(n10566), .B1(n14853), .B2(n12751), .ZN(
        n9878) );
  OR3_X1 U12348 ( .A1(n9880), .A2(n9879), .A3(n9878), .ZN(P2_U3190) );
  INV_X2 U12349 ( .A(n12646), .ZN(n11970) );
  INV_X1 U12350 ( .A(n9881), .ZN(n9884) );
  MUX2_X1 U12351 ( .A(n9882), .B(n15207), .S(P3_STATE_REG_SCAN_IN), .Z(n9883)
         );
  OAI21_X1 U12352 ( .B1(n11970), .B2(n9884), .A(n9883), .ZN(P3_U3295) );
  INV_X1 U12353 ( .A(n10416), .ZN(n10519) );
  INV_X1 U12354 ( .A(SI_2_), .ZN(n9885) );
  NAND2_X2 U12355 ( .A1(n9926), .A2(P3_U3151), .ZN(n11881) );
  OAI222_X1 U12356 ( .A1(n10519), .A2(P3_U3151), .B1(n11970), .B2(n9886), .C1(
        n9885), .C2(n11881), .ZN(P3_U3293) );
  INV_X1 U12357 ( .A(n9887), .ZN(n9889) );
  OAI222_X1 U12358 ( .A1(n11970), .A2(n9889), .B1(n11881), .B2(n9888), .C1(
        n11077), .C2(P3_U3151), .ZN(P3_U3287) );
  INV_X1 U12359 ( .A(n9890), .ZN(n9928) );
  INV_X2 U12360 ( .A(n13450), .ZN(n13459) );
  NAND2_X2 U12361 ( .A1(n9925), .A2(P2_U3088), .ZN(n13464) );
  NAND2_X1 U12362 ( .A1(n9894), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9891) );
  NAND2_X1 U12363 ( .A1(n10086), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14771) );
  OAI211_X1 U12364 ( .C1(n9928), .C2(n13459), .A(n9891), .B(n14771), .ZN(
        P2_U3323) );
  INV_X1 U12365 ( .A(n11233), .ZN(n11073) );
  OAI222_X1 U12366 ( .A1(n11073), .A2(P3_U3151), .B1(n11970), .B2(n9893), .C1(
        n9892), .C2(n11881), .ZN(P3_U3286) );
  INV_X1 U12367 ( .A(n9895), .ZN(n9933) );
  INV_X1 U12368 ( .A(n10083), .ZN(n10146) );
  OAI222_X1 U12369 ( .A1(n13464), .A2(n9896), .B1(n13459), .B2(n9933), .C1(
        P2_U3088), .C2(n10146), .ZN(P2_U3324) );
  INV_X1 U12370 ( .A(n9897), .ZN(n9935) );
  INV_X1 U12371 ( .A(n10078), .ZN(n14745) );
  OAI222_X1 U12372 ( .A1(n13464), .A2(n9898), .B1(n13459), .B2(n9935), .C1(
        P2_U3088), .C2(n14745), .ZN(P2_U3326) );
  INV_X1 U12373 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9900) );
  INV_X1 U12374 ( .A(n9899), .ZN(n9931) );
  INV_X1 U12375 ( .A(n10110), .ZN(n10097) );
  OAI222_X1 U12376 ( .A1(n13464), .A2(n9900), .B1(n13459), .B2(n9931), .C1(
        P2_U3088), .C2(n10097), .ZN(P2_U3322) );
  INV_X1 U12377 ( .A(n10080), .ZN(n14758) );
  OAI222_X1 U12378 ( .A1(n13464), .A2(n9901), .B1(n13459), .B2(n9943), .C1(
        P2_U3088), .C2(n14758), .ZN(P2_U3325) );
  INV_X1 U12379 ( .A(SI_4_), .ZN(n9902) );
  INV_X1 U12380 ( .A(n10724), .ZN(n10525) );
  OAI222_X1 U12381 ( .A1(n11970), .A2(n9903), .B1(n11881), .B2(n9902), .C1(
        n10525), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12382 ( .A(SI_10_), .ZN(n9904) );
  INV_X1 U12383 ( .A(n11529), .ZN(n11246) );
  OAI222_X1 U12384 ( .A1(n11970), .A2(n9905), .B1(n11881), .B2(n9904), .C1(
        n11246), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12385 ( .A(n10634), .ZN(n10526) );
  INV_X1 U12386 ( .A(SI_5_), .ZN(n9907) );
  OAI222_X1 U12387 ( .A1(P3_U3151), .A2(n10526), .B1(n11881), .B2(n9907), .C1(
        n11970), .C2(n9906), .ZN(P3_U3290) );
  INV_X1 U12388 ( .A(n10647), .ZN(n10522) );
  INV_X1 U12389 ( .A(SI_3_), .ZN(n9908) );
  OAI222_X1 U12390 ( .A1(n10522), .A2(P3_U3151), .B1(n11970), .B2(n9909), .C1(
        n9908), .C2(n11881), .ZN(P3_U3292) );
  INV_X1 U12391 ( .A(n9910), .ZN(n9912) );
  OAI222_X1 U12392 ( .A1(n10675), .A2(P3_U3151), .B1(n11970), .B2(n9912), .C1(
        n9911), .C2(n11881), .ZN(P3_U3289) );
  INV_X1 U12393 ( .A(n9913), .ZN(n9915) );
  OAI222_X1 U12394 ( .A1(n10456), .A2(P3_U3151), .B1(n11970), .B2(n9915), .C1(
        n9914), .C2(n11881), .ZN(P3_U3294) );
  INV_X1 U12395 ( .A(n11059), .ZN(n10678) );
  INV_X1 U12396 ( .A(SI_7_), .ZN(n9916) );
  OAI222_X1 U12397 ( .A1(n10678), .A2(P3_U3151), .B1(n11970), .B2(n9917), .C1(
        n9916), .C2(n11881), .ZN(P3_U3288) );
  INV_X1 U12398 ( .A(n9918), .ZN(n9946) );
  INV_X1 U12399 ( .A(n10126), .ZN(n9919) );
  OAI222_X1 U12400 ( .A1(n13464), .A2(n9920), .B1(n13459), .B2(n9946), .C1(
        P2_U3088), .C2(n9919), .ZN(P2_U3321) );
  OR2_X1 U12401 ( .A1(n10006), .A2(n9737), .ZN(n9972) );
  INV_X1 U12402 ( .A(n10014), .ZN(n9923) );
  AOI21_X1 U12403 ( .B1(n9923), .B2(n9922), .A(n9921), .ZN(n9971) );
  INV_X1 U12404 ( .A(n9971), .ZN(n9924) );
  AND2_X1 U12405 ( .A1(n9972), .A2(n9924), .ZN(n14491) );
  NOR2_X1 U12406 ( .A1(n14491), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U12407 ( .A(n14171), .ZN(n11815) );
  INV_X1 U12408 ( .A(n11815), .ZN(n14166) );
  INV_X1 U12409 ( .A(n14163), .ZN(n14151) );
  AOI22_X1 U12410 ( .A1(n13823), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n14151), .ZN(n9927) );
  OAI21_X1 U12411 ( .B1(n9928), .B2(n14166), .A(n9927), .ZN(P1_U3351) );
  INV_X1 U12412 ( .A(n9929), .ZN(n9940) );
  AOI22_X1 U12413 ( .A1(n10432), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n14151), .ZN(n9930) );
  OAI21_X1 U12414 ( .B1(n9940), .B2(n14171), .A(n9930), .ZN(P1_U3348) );
  INV_X1 U12415 ( .A(n10044), .ZN(n10003) );
  OAI222_X1 U12416 ( .A1(n9985), .A2(P1_U3086), .B1(n14166), .B2(n9935), .C1(
        n6773), .C2(n14163), .ZN(P1_U3354) );
  AOI22_X1 U12417 ( .A1(n14650), .A2(n10195), .B1(n10194), .B2(n9937), .ZN(
        P1_U3446) );
  AOI22_X1 U12418 ( .A1(n14650), .A2(n9939), .B1(n9938), .B2(n9937), .ZN(
        P1_U3445) );
  INV_X1 U12419 ( .A(n10216), .ZN(n10133) );
  OAI222_X1 U12420 ( .A1(n13464), .A2(n9941), .B1(n13459), .B2(n9940), .C1(
        P2_U3088), .C2(n10133), .ZN(P2_U3320) );
  INV_X1 U12421 ( .A(n13788), .ZN(n9944) );
  OAI222_X1 U12422 ( .A1(n9944), .A2(P1_U3086), .B1(n14166), .B2(n9943), .C1(
        n9942), .C2(n14163), .ZN(P1_U3353) );
  INV_X1 U12423 ( .A(n10252), .ZN(n9947) );
  OAI222_X1 U12424 ( .A1(n9947), .A2(P1_U3086), .B1(n14166), .B2(n9946), .C1(
        n9945), .C2(n14163), .ZN(P1_U3349) );
  AND2_X1 U12425 ( .A1(n9957), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12426 ( .A1(n9957), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12427 ( .A1(n9957), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12428 ( .A1(n9957), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12429 ( .A1(n9957), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12430 ( .A1(n9957), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12431 ( .A1(n9957), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12432 ( .A1(n9957), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12433 ( .A1(n9957), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12434 ( .A1(n9957), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12435 ( .A1(n9957), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12436 ( .A1(n9957), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12437 ( .A1(n9957), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12438 ( .A1(n9957), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12439 ( .A1(n9957), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12440 ( .A1(n9957), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12441 ( .A1(n9957), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12442 ( .A1(n9957), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12443 ( .A1(n9957), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12444 ( .A1(n9957), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12445 ( .A1(n9957), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12446 ( .A1(n9957), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12447 ( .A1(n9957), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12448 ( .A1(n9957), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12449 ( .A1(n9957), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12450 ( .A1(n9957), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12451 ( .A1(n9957), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12452 ( .A1(n9957), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  INV_X1 U12453 ( .A(n9949), .ZN(n9951) );
  OAI222_X1 U12454 ( .A1(n11881), .A2(n9952), .B1(n11970), .B2(n9951), .C1(
        P3_U3151), .C2(n9950), .ZN(P3_U3284) );
  INV_X1 U12455 ( .A(n9953), .ZN(n9956) );
  OAI222_X1 U12456 ( .A1(n13464), .A2(n9954), .B1(n13459), .B2(n9956), .C1(
        P2_U3088), .C2(n13079), .ZN(P2_U3319) );
  INV_X1 U12457 ( .A(n10734), .ZN(n10430) );
  OAI222_X1 U12458 ( .A1(n10430), .A2(P1_U3086), .B1(n14171), .B2(n9956), .C1(
        n9955), .C2(n14163), .ZN(P1_U3347) );
  INV_X1 U12459 ( .A(n9957), .ZN(n9958) );
  INV_X1 U12460 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n15245) );
  NOR2_X1 U12461 ( .A1(n9958), .A2(n15245), .ZN(P3_U3241) );
  INV_X1 U12462 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n15218) );
  NOR2_X1 U12463 ( .A1(n9958), .A2(n15218), .ZN(P3_U3244) );
  INV_X1 U12464 ( .A(n11618), .ZN(n11787) );
  OAI222_X1 U12465 ( .A1(n11970), .A2(n9960), .B1(n11881), .B2(n9959), .C1(
        n11787), .C2(P3_U3151), .ZN(P3_U3283) );
  INV_X1 U12466 ( .A(n10987), .ZN(n10732) );
  INV_X1 U12467 ( .A(n9961), .ZN(n9962) );
  OAI222_X1 U12468 ( .A1(n10732), .A2(P1_U3086), .B1(n14171), .B2(n9962), .C1(
        n7296), .C2(n14163), .ZN(P1_U3346) );
  INV_X1 U12469 ( .A(n10222), .ZN(n14792) );
  OAI222_X1 U12470 ( .A1(n13464), .A2(n9963), .B1(n13459), .B2(n9962), .C1(
        P2_U3088), .C2(n14792), .ZN(P2_U3318) );
  INV_X1 U12471 ( .A(n9964), .ZN(n9966) );
  INV_X1 U12472 ( .A(n10237), .ZN(n10227) );
  OAI222_X1 U12473 ( .A1(n13459), .A2(n9966), .B1(n10227), .B2(P2_U3088), .C1(
        n9965), .C2(n13464), .ZN(P2_U3317) );
  INV_X1 U12474 ( .A(n11428), .ZN(n10991) );
  INV_X1 U12475 ( .A(n12210), .ZN(n9968) );
  OAI222_X1 U12476 ( .A1(n11970), .A2(n9970), .B1(n11881), .B2(n9969), .C1(
        n9968), .C2(P3_U3151), .ZN(P3_U3282) );
  NAND2_X1 U12477 ( .A1(n9972), .A2(n9971), .ZN(n14493) );
  NAND2_X1 U12478 ( .A1(n6720), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9978) );
  INV_X1 U12479 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n14725) );
  MUX2_X1 U12480 ( .A(n14725), .B(P1_REG1_REG_1__SCAN_IN), .S(n9985), .Z(n9974) );
  INV_X1 U12481 ( .A(n9974), .ZN(n9977) );
  AND2_X1 U12482 ( .A1(n6720), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9973) );
  NAND2_X1 U12483 ( .A1(n9974), .A2(n9973), .ZN(n9987) );
  INV_X1 U12484 ( .A(n9987), .ZN(n9976) );
  INV_X1 U12485 ( .A(n6459), .ZN(n9975) );
  AOI211_X1 U12486 ( .C1(n9978), .C2(n9977), .A(n9976), .B(n14576), .ZN(n9982)
         );
  INV_X1 U12487 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9979) );
  MUX2_X1 U12488 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9979), .S(n9985), .Z(n9980)
         );
  NAND2_X1 U12489 ( .A1(n6720), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13782) );
  AOI211_X1 U12490 ( .C1(n9980), .C2(n13782), .A(n9992), .B(n14572), .ZN(n9981) );
  NOR2_X1 U12491 ( .A1(n9982), .A2(n9981), .ZN(n9984) );
  AOI22_X1 U12492 ( .A1(n14491), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9983) );
  OAI211_X1 U12493 ( .C1(n9985), .C2(n14566), .A(n9984), .B(n9983), .ZN(
        P1_U3244) );
  XOR2_X1 U12494 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n10044), .Z(n9991) );
  INV_X1 U12495 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n14727) );
  MUX2_X1 U12496 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n14727), .S(n13788), .Z(
        n13795) );
  NAND2_X1 U12497 ( .A1(n9993), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U12498 ( .A1(n9987), .A2(n9986), .ZN(n13794) );
  NAND2_X1 U12499 ( .A1(n13795), .A2(n13794), .ZN(n13793) );
  NAND2_X1 U12500 ( .A1(n13788), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U12501 ( .A1(n13793), .A2(n9988), .ZN(n13807) );
  XNOR2_X1 U12502 ( .A(n9994), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n13808) );
  NAND2_X1 U12503 ( .A1(n13807), .A2(n13808), .ZN(n13806) );
  INV_X1 U12504 ( .A(n9994), .ZN(n13805) );
  NAND2_X1 U12505 ( .A1(n13805), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9989) );
  NAND2_X1 U12506 ( .A1(n13806), .A2(n9989), .ZN(n13819) );
  INV_X1 U12507 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15265) );
  MUX2_X1 U12508 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n15265), .S(n13823), .Z(
        n13818) );
  AND2_X1 U12509 ( .A1(n13819), .A2(n13818), .ZN(n13821) );
  NAND2_X1 U12510 ( .A1(n9990), .A2(n9991), .ZN(n10043) );
  OAI21_X1 U12511 ( .B1(n9991), .B2(n9990), .A(n10043), .ZN(n9999) );
  AOI21_X1 U12512 ( .B1(n9993), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9992), .ZN(
        n13791) );
  MUX2_X1 U12513 ( .A(n8280), .B(P1_REG2_REG_2__SCAN_IN), .S(n13788), .Z(
        n13790) );
  MUX2_X1 U12514 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9995), .S(n9994), .Z(n13800) );
  XNOR2_X1 U12515 ( .A(n13823), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n13814) );
  NOR2_X1 U12516 ( .A1(n13815), .A2(n13814), .ZN(n13813) );
  XNOR2_X1 U12517 ( .A(n10044), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9996) );
  AOI211_X1 U12518 ( .C1(n9997), .C2(n9996), .A(n14572), .B(n10038), .ZN(n9998) );
  AOI21_X1 U12519 ( .B1(n14558), .B2(n9999), .A(n9998), .ZN(n10002) );
  NAND2_X1 U12520 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10898) );
  INV_X1 U12521 ( .A(n10898), .ZN(n10000) );
  AOI21_X1 U12522 ( .B1(n14491), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n10000), .ZN(
        n10001) );
  OAI211_X1 U12523 ( .C1(n10003), .C2(n14566), .A(n10002), .B(n10001), .ZN(
        P1_U3248) );
  INV_X1 U12524 ( .A(n10004), .ZN(n10005) );
  NAND2_X1 U12525 ( .A1(n11587), .A2(n10005), .ZN(n10030) );
  INV_X1 U12526 ( .A(n10030), .ZN(n10007) );
  AND2_X1 U12527 ( .A1(n10007), .A2(n10006), .ZN(n10016) );
  INV_X1 U12528 ( .A(n10008), .ZN(n10009) );
  NAND2_X1 U12529 ( .A1(n10016), .A2(n10009), .ZN(n10010) );
  INV_X1 U12530 ( .A(n14398), .ZN(n13742) );
  NOR2_X1 U12531 ( .A1(n10012), .A2(n10011), .ZN(n10013) );
  AND2_X1 U12532 ( .A1(n14717), .A2(n10014), .ZN(n10015) );
  AND2_X2 U12533 ( .A1(n14675), .A2(n13587), .ZN(n10463) );
  NAND2_X1 U12534 ( .A1(n10017), .A2(n10463), .ZN(n10022) );
  OR2_X2 U12535 ( .A1(n10019), .A2(n10018), .ZN(n13627) );
  OAI22_X1 U12536 ( .A1(n14628), .A2(n13627), .B1(n10023), .B2(n13784), .ZN(
        n10020) );
  INV_X1 U12537 ( .A(n10020), .ZN(n10021) );
  AND2_X1 U12538 ( .A1(n10022), .A2(n10021), .ZN(n10027) );
  INV_X2 U12539 ( .A(n13627), .ZN(n10153) );
  NAND2_X1 U12540 ( .A1(n10017), .A2(n6460), .ZN(n10026) );
  INV_X1 U12541 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14488) );
  OAI22_X1 U12542 ( .A1(n14628), .A2(n13629), .B1(n10023), .B2(n14488), .ZN(
        n10024) );
  INV_X1 U12543 ( .A(n10024), .ZN(n10025) );
  NAND2_X1 U12544 ( .A1(n10026), .A2(n10025), .ZN(n10147) );
  NAND2_X1 U12545 ( .A1(n10027), .A2(n10147), .ZN(n10150) );
  OAI21_X1 U12546 ( .B1(n10027), .B2(n10147), .A(n10150), .ZN(n13781) );
  NOR2_X2 U12547 ( .A1(n10030), .A2(n10193), .ZN(n14397) );
  NAND2_X1 U12548 ( .A1(n14629), .A2(n13732), .ZN(n11934) );
  INV_X1 U12549 ( .A(n10191), .ZN(n10029) );
  NAND2_X1 U12550 ( .A1(n10030), .A2(n10029), .ZN(n10474) );
  INV_X1 U12551 ( .A(n10193), .ZN(n10031) );
  NAND2_X1 U12552 ( .A1(n10474), .A2(n10031), .ZN(n10270) );
  INV_X1 U12553 ( .A(n10270), .ZN(n10032) );
  INV_X1 U12554 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11933) );
  OAI22_X1 U12555 ( .A1(n13737), .A2(n11934), .B1(n10032), .B2(n11933), .ZN(
        n10033) );
  AOI21_X1 U12556 ( .B1(n14395), .B2(n13781), .A(n10033), .ZN(n10034) );
  OAI21_X1 U12557 ( .B1(n13742), .B2(n14628), .A(n10034), .ZN(P1_U3232) );
  INV_X1 U12558 ( .A(n11430), .ZN(n14498) );
  INV_X1 U12559 ( .A(n10035), .ZN(n10036) );
  INV_X1 U12560 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n15224) );
  OAI222_X1 U12561 ( .A1(n14498), .A2(P1_U3086), .B1(n14171), .B2(n10036), 
        .C1(n15224), .C2(n14163), .ZN(P1_U3344) );
  INV_X1 U12562 ( .A(n10304), .ZN(n10296) );
  OAI222_X1 U12563 ( .A1(n13464), .A2(n10037), .B1(n13459), .B2(n10036), .C1(
        P2_U3088), .C2(n10296), .ZN(P2_U3316) );
  INV_X1 U12564 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10039) );
  MUX2_X1 U12565 ( .A(n10039), .B(P1_REG2_REG_6__SCAN_IN), .S(n10252), .Z(
        n10040) );
  AOI211_X1 U12566 ( .C1(n10041), .C2(n10040), .A(n14572), .B(n10248), .ZN(
        n10051) );
  INV_X1 U12567 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10042) );
  MUX2_X1 U12568 ( .A(n10042), .B(P1_REG1_REG_6__SCAN_IN), .S(n10252), .Z(
        n10046) );
  OAI21_X1 U12569 ( .B1(n10044), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10043), .ZN(
        n10045) );
  NOR2_X1 U12570 ( .A1(n10045), .A2(n10046), .ZN(n10251) );
  AOI211_X1 U12571 ( .C1(n10046), .C2(n10045), .A(n14576), .B(n10251), .ZN(
        n10050) );
  NAND2_X1 U12572 ( .A1(n14582), .A2(n10252), .ZN(n10048) );
  NAND2_X1 U12573 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10047) );
  OAI211_X1 U12574 ( .C1(n14193), .C2(n14585), .A(n10048), .B(n10047), .ZN(
        n10049) );
  OR3_X1 U12575 ( .A1(n10051), .A2(n10050), .A3(n10049), .ZN(P1_U3249) );
  INV_X1 U12576 ( .A(n11812), .ZN(n10056) );
  NAND2_X1 U12577 ( .A1(n10052), .A2(n11812), .ZN(n10054) );
  NAND2_X1 U12578 ( .A1(n10054), .A2(n10053), .ZN(n10055) );
  NAND2_X1 U12579 ( .A1(n10089), .A2(n10058), .ZN(n14772) );
  INV_X1 U12580 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10074) );
  NAND2_X1 U12581 ( .A1(n10059), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13451) );
  NOR2_X1 U12582 ( .A1(n13451), .A2(n13454), .ZN(n10060) );
  INV_X1 U12583 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10061) );
  MUX2_X1 U12584 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10061), .S(n10086), .Z(
        n14775) );
  INV_X1 U12585 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10062) );
  XNOR2_X1 U12586 ( .A(n10080), .B(n10062), .ZN(n14760) );
  NAND2_X1 U12587 ( .A1(n10078), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10064) );
  OAI21_X1 U12588 ( .B1(n10078), .B2(P2_REG2_REG_1__SCAN_IN), .A(n10064), .ZN(
        n14747) );
  NAND2_X1 U12589 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10063) );
  OR2_X1 U12590 ( .A1(n14747), .A2(n10063), .ZN(n14750) );
  NAND2_X1 U12591 ( .A1(n14750), .A2(n10064), .ZN(n14761) );
  NAND2_X1 U12592 ( .A1(n14760), .A2(n14761), .ZN(n10066) );
  NAND2_X1 U12593 ( .A1(n10080), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10065) );
  NAND2_X1 U12594 ( .A1(n10066), .A2(n10065), .ZN(n10139) );
  INV_X1 U12595 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10618) );
  MUX2_X1 U12596 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10618), .S(n10083), .Z(
        n10140) );
  NAND2_X1 U12597 ( .A1(n10139), .A2(n10140), .ZN(n10138) );
  NAND2_X1 U12598 ( .A1(n10083), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10067) );
  NAND2_X1 U12599 ( .A1(n10138), .A2(n10067), .ZN(n14776) );
  NAND2_X1 U12600 ( .A1(n14775), .A2(n14776), .ZN(n14774) );
  NAND2_X1 U12601 ( .A1(n10086), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10071) );
  NAND2_X1 U12602 ( .A1(n14774), .A2(n10071), .ZN(n10069) );
  INV_X1 U12603 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10586) );
  MUX2_X1 U12604 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10586), .S(n10110), .Z(
        n10068) );
  NAND2_X1 U12605 ( .A1(n10069), .A2(n10068), .ZN(n10106) );
  MUX2_X1 U12606 ( .A(n10586), .B(P2_REG2_REG_5__SCAN_IN), .S(n10110), .Z(
        n10070) );
  NAND3_X1 U12607 ( .A1(n14774), .A2(n10071), .A3(n10070), .ZN(n10072) );
  NAND3_X1 U12608 ( .A1(n14805), .A2(n10106), .A3(n10072), .ZN(n10073) );
  OAI21_X1 U12609 ( .B1(n10074), .B2(n14811), .A(n10073), .ZN(n10095) );
  INV_X1 U12610 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10075) );
  XNOR2_X1 U12611 ( .A(n10110), .B(n10075), .ZN(n10091) );
  INV_X1 U12612 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10076) );
  XNOR2_X1 U12613 ( .A(n10080), .B(n10076), .ZN(n14756) );
  INV_X1 U12614 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10077) );
  XNOR2_X1 U12615 ( .A(n10078), .B(n10077), .ZN(n14743) );
  AND2_X1 U12616 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14742) );
  NAND2_X1 U12617 ( .A1(n14743), .A2(n14742), .ZN(n14741) );
  NAND2_X1 U12618 ( .A1(n10078), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10079) );
  NAND2_X1 U12619 ( .A1(n10080), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10081) );
  INV_X1 U12620 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10082) );
  XNOR2_X1 U12621 ( .A(n10083), .B(n10082), .ZN(n10136) );
  NAND2_X1 U12622 ( .A1(n10083), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10084) );
  NAND2_X1 U12623 ( .A1(n10134), .A2(n10084), .ZN(n14767) );
  INV_X1 U12624 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10085) );
  XNOR2_X1 U12625 ( .A(n10086), .B(n10085), .ZN(n14768) );
  NAND2_X1 U12626 ( .A1(n14767), .A2(n14768), .ZN(n14766) );
  NAND2_X1 U12627 ( .A1(n10086), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10087) );
  INV_X1 U12628 ( .A(n13454), .ZN(n13035) );
  NOR2_X1 U12629 ( .A1(n13451), .A2(n13035), .ZN(n10088) );
  OAI211_X1 U12630 ( .C1(n10091), .C2(n10090), .A(n14784), .B(n10112), .ZN(
        n10092) );
  INV_X1 U12631 ( .A(n10092), .ZN(n10094) );
  AND2_X1 U12632 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10093) );
  NOR3_X1 U12633 ( .A1(n10095), .A2(n10094), .A3(n10093), .ZN(n10096) );
  OAI21_X1 U12634 ( .B1(n10097), .B2(n14827), .A(n10096), .ZN(P2_U3219) );
  INV_X1 U12635 ( .A(n10098), .ZN(n10100) );
  OAI222_X1 U12636 ( .A1(n11970), .A2(n10100), .B1(n11881), .B2(n10099), .C1(
        n12197), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12637 ( .A(n14827), .ZN(n14804) );
  NAND2_X1 U12638 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10906) );
  INV_X1 U12639 ( .A(n10906), .ZN(n10109) );
  NAND2_X1 U12640 ( .A1(n10110), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10105) );
  NAND2_X1 U12641 ( .A1(n10106), .A2(n10105), .ZN(n10103) );
  INV_X1 U12642 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10101) );
  MUX2_X1 U12643 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10101), .S(n10126), .Z(
        n10102) );
  NAND2_X1 U12644 ( .A1(n10103), .A2(n10102), .ZN(n10122) );
  MUX2_X1 U12645 ( .A(n10101), .B(P2_REG2_REG_6__SCAN_IN), .S(n10126), .Z(
        n10104) );
  NAND3_X1 U12646 ( .A1(n10106), .A2(n10105), .A3(n10104), .ZN(n10107) );
  AND3_X1 U12647 ( .A1(n14805), .A2(n10122), .A3(n10107), .ZN(n10108) );
  AOI211_X1 U12648 ( .C1(n14804), .C2(n10126), .A(n10109), .B(n10108), .ZN(
        n10116) );
  INV_X1 U12649 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10610) );
  MUX2_X1 U12650 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10610), .S(n10126), .Z(
        n10114) );
  NAND2_X1 U12651 ( .A1(n10110), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10111) );
  OAI211_X1 U12652 ( .C1(n10114), .C2(n10113), .A(n14784), .B(n10128), .ZN(
        n10115) );
  OAI211_X1 U12653 ( .C1(n7003), .C2(n14811), .A(n10116), .B(n10115), .ZN(
        P2_U3220) );
  INV_X1 U12654 ( .A(n14811), .ZN(n14819) );
  NOR2_X1 U12655 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7844), .ZN(n10125) );
  NAND2_X1 U12656 ( .A1(n10126), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10121) );
  NAND2_X1 U12657 ( .A1(n10122), .A2(n10121), .ZN(n10119) );
  INV_X1 U12658 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10117) );
  MUX2_X1 U12659 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10117), .S(n10216), .Z(
        n10118) );
  NAND2_X1 U12660 ( .A1(n10119), .A2(n10118), .ZN(n13082) );
  MUX2_X1 U12661 ( .A(n10117), .B(P2_REG2_REG_7__SCAN_IN), .S(n10216), .Z(
        n10120) );
  NAND3_X1 U12662 ( .A1(n10122), .A2(n10121), .A3(n10120), .ZN(n10123) );
  AND3_X1 U12663 ( .A1(n14805), .A2(n13082), .A3(n10123), .ZN(n10124) );
  AOI211_X1 U12664 ( .C1(n14819), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n10125), .B(
        n10124), .ZN(n10132) );
  INV_X1 U12665 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n14906) );
  MUX2_X1 U12666 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n14906), .S(n10216), .Z(
        n10130) );
  NAND2_X1 U12667 ( .A1(n10126), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10127) );
  NAND2_X1 U12668 ( .A1(n10128), .A2(n10127), .ZN(n10129) );
  OAI211_X1 U12669 ( .C1(n10130), .C2(n10129), .A(n14784), .B(n10210), .ZN(
        n10131) );
  OAI211_X1 U12670 ( .C1(n14827), .C2(n10133), .A(n10132), .B(n10131), .ZN(
        P2_U3221) );
  OAI211_X1 U12671 ( .C1(n10136), .C2(n10135), .A(n14784), .B(n10134), .ZN(
        n10137) );
  INV_X1 U12672 ( .A(n10137), .ZN(n10144) );
  INV_X1 U12673 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10142) );
  OAI211_X1 U12674 ( .C1(n10140), .C2(n10139), .A(n14805), .B(n10138), .ZN(
        n10141) );
  OAI21_X1 U12675 ( .B1(n10142), .B2(n14811), .A(n10141), .ZN(n10143) );
  AOI211_X1 U12676 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(P2_U3088), .A(n10144), 
        .B(n10143), .ZN(n10145) );
  OAI21_X1 U12677 ( .B1(n10146), .B2(n14827), .A(n10145), .ZN(P2_U3217) );
  INV_X1 U12678 ( .A(n10147), .ZN(n10148) );
  NAND2_X1 U12679 ( .A1(n10148), .A2(n13625), .ZN(n10149) );
  NAND2_X1 U12680 ( .A1(n14629), .A2(n10153), .ZN(n10152) );
  NAND2_X1 U12681 ( .A1(n10167), .A2(n13587), .ZN(n10151) );
  NAND2_X1 U12682 ( .A1(n14629), .A2(n10463), .ZN(n10155) );
  NAND2_X1 U12683 ( .A1(n10167), .A2(n10153), .ZN(n10154) );
  AND2_X1 U12684 ( .A1(n10155), .A2(n10154), .ZN(n10157) );
  INV_X1 U12685 ( .A(n10156), .ZN(n10159) );
  INV_X1 U12686 ( .A(n10157), .ZN(n10158) );
  NAND2_X1 U12687 ( .A1(n10159), .A2(n10158), .ZN(n10160) );
  INV_X1 U12688 ( .A(n10266), .ZN(n10161) );
  AOI21_X1 U12689 ( .B1(n10163), .B2(n10162), .A(n10161), .ZN(n10170) );
  INV_X1 U12690 ( .A(n10017), .ZN(n14625) );
  NOR2_X1 U12691 ( .A1(n10164), .A2(n14385), .ZN(n14636) );
  INV_X1 U12692 ( .A(n14636), .ZN(n10165) );
  OAI21_X1 U12693 ( .B1(n14625), .B2(n14633), .A(n10165), .ZN(n10166) );
  AOI22_X1 U12694 ( .A1(n10166), .A2(n14397), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10270), .ZN(n10169) );
  NAND2_X1 U12695 ( .A1(n14398), .A2(n10167), .ZN(n10168) );
  OAI211_X1 U12696 ( .C1(n10170), .C2(n13751), .A(n10169), .B(n10168), .ZN(
        P1_U3222) );
  INV_X1 U12697 ( .A(n10171), .ZN(n10173) );
  OAI222_X1 U12698 ( .A1(n11970), .A2(n10173), .B1(n11881), .B2(n10172), .C1(
        n12260), .C2(P3_U3151), .ZN(P3_U3280) );
  AOI22_X1 U12699 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n14805), .B1(n14784), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10178) );
  INV_X1 U12700 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10174) );
  NAND2_X1 U12701 ( .A1(n14784), .A2(n10174), .ZN(n10176) );
  INV_X1 U12702 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n14748) );
  NAND2_X1 U12703 ( .A1(n14805), .A2(n14748), .ZN(n10175) );
  AND3_X1 U12704 ( .A1(n14827), .A2(n10176), .A3(n10175), .ZN(n10177) );
  MUX2_X1 U12705 ( .A(n10178), .B(n10177), .S(P2_IR_REG_0__SCAN_IN), .Z(n10182) );
  INV_X1 U12706 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10179) );
  INV_X1 U12707 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10488) );
  OAI22_X1 U12708 ( .A1(n14811), .A2(n10179), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10488), .ZN(n10180) );
  INV_X1 U12709 ( .A(n10180), .ZN(n10181) );
  NAND2_X1 U12710 ( .A1(n10182), .A2(n10181), .ZN(P2_U3214) );
  INV_X1 U12711 ( .A(n10183), .ZN(n10185) );
  INV_X1 U12712 ( .A(n10538), .ZN(n10545) );
  OAI222_X1 U12713 ( .A1(n13459), .A2(n10185), .B1(n10545), .B2(P2_U3088), 
        .C1(n10184), .C2(n13464), .ZN(P2_U3315) );
  INV_X1 U12714 ( .A(n11862), .ZN(n11426) );
  NAND2_X1 U12715 ( .A1(n12928), .A2(n13071), .ZN(n10187) );
  OAI21_X1 U12716 ( .B1(n11453), .B2(n13071), .A(n10187), .ZN(P2_U3551) );
  INV_X1 U12717 ( .A(n10188), .ZN(n10189) );
  NOR2_X1 U12718 ( .A1(n10190), .A2(n10189), .ZN(n10192) );
  OR3_X1 U12719 ( .A1(n10193), .A2(n10192), .A3(n10191), .ZN(n10198) );
  AOI21_X1 U12720 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(n10197) );
  NOR2_X1 U12721 ( .A1(n10198), .A2(n10197), .ZN(n11588) );
  INV_X1 U12722 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10207) );
  OR2_X1 U12723 ( .A1(n10200), .A2(n14023), .ZN(n14690) );
  NOR2_X1 U12724 ( .A1(n14714), .A2(n14630), .ZN(n10205) );
  NAND3_X1 U12725 ( .A1(n10203), .A2(n10202), .A3(n11558), .ZN(n10204) );
  OAI211_X1 U12726 ( .C1(n10205), .C2(n9685), .A(n11934), .B(n10204), .ZN(
        n14134) );
  NAND2_X1 U12727 ( .A1(n14134), .A2(n14724), .ZN(n10206) );
  OAI21_X1 U12728 ( .B1(n14724), .B2(n10207), .A(n10206), .ZN(P1_U3459) );
  INV_X1 U12729 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10208) );
  MUX2_X1 U12730 ( .A(n10208), .B(P2_REG1_REG_10__SCAN_IN), .S(n10237), .Z(
        n10215) );
  NAND2_X1 U12731 ( .A1(n10216), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10209) );
  INV_X1 U12732 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14908) );
  MUX2_X1 U12733 ( .A(n14908), .B(P2_REG1_REG_8__SCAN_IN), .S(n13079), .Z(
        n13078) );
  INV_X1 U12734 ( .A(n13079), .ZN(n10211) );
  NAND2_X1 U12735 ( .A1(n10211), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10212) );
  INV_X1 U12736 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10213) );
  MUX2_X1 U12737 ( .A(n10213), .B(P2_REG1_REG_9__SCAN_IN), .S(n10222), .Z(
        n14780) );
  OR2_X1 U12738 ( .A1(n14781), .A2(n14780), .ZN(n14783) );
  OAI21_X1 U12739 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n10222), .A(n14783), .ZN(
        n10214) );
  NOR2_X1 U12740 ( .A1(n10214), .A2(n10215), .ZN(n10236) );
  AOI211_X1 U12741 ( .C1(n10215), .C2(n10214), .A(n14813), .B(n10236), .ZN(
        n10230) );
  NAND2_X1 U12742 ( .A1(n10216), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n13081) );
  NAND2_X1 U12743 ( .A1(n13082), .A2(n13081), .ZN(n10219) );
  INV_X1 U12744 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10217) );
  MUX2_X1 U12745 ( .A(n10217), .B(P2_REG2_REG_8__SCAN_IN), .S(n13079), .Z(
        n10218) );
  NAND2_X1 U12746 ( .A1(n10219), .A2(n10218), .ZN(n13084) );
  OR2_X1 U12747 ( .A1(n13079), .A2(n10217), .ZN(n10220) );
  AND2_X1 U12748 ( .A1(n13084), .A2(n10220), .ZN(n14788) );
  INV_X1 U12749 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10221) );
  MUX2_X1 U12750 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10221), .S(n10222), .Z(
        n14787) );
  NAND2_X1 U12751 ( .A1(n14788), .A2(n14787), .ZN(n14786) );
  OAI21_X1 U12752 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n10222), .A(n14786), .ZN(
        n10225) );
  INV_X1 U12753 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10223) );
  MUX2_X1 U12754 ( .A(n10223), .B(P2_REG2_REG_10__SCAN_IN), .S(n10237), .Z(
        n10224) );
  INV_X1 U12755 ( .A(n14805), .ZN(n14823) );
  NOR2_X1 U12756 ( .A1(n10225), .A2(n10224), .ZN(n10231) );
  AOI211_X1 U12757 ( .C1(n10225), .C2(n10224), .A(n14823), .B(n10231), .ZN(
        n10229) );
  NOR2_X1 U12758 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n15103), .ZN(n11276) );
  AOI21_X1 U12759 ( .B1(n14819), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n11276), 
        .ZN(n10226) );
  OAI21_X1 U12760 ( .B1(n10227), .B2(n14827), .A(n10226), .ZN(n10228) );
  OR3_X1 U12761 ( .A1(n10230), .A2(n10229), .A3(n10228), .ZN(P2_U3224) );
  AOI21_X1 U12762 ( .B1(n10237), .B2(P2_REG2_REG_10__SCAN_IN), .A(n10231), 
        .ZN(n10234) );
  INV_X1 U12763 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10297) );
  MUX2_X1 U12764 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10297), .S(n10304), .Z(
        n10233) );
  AND2_X1 U12765 ( .A1(n10234), .A2(n10233), .ZN(n10295) );
  INV_X1 U12766 ( .A(n10295), .ZN(n10232) );
  OAI21_X1 U12767 ( .B1(n10234), .B2(n10233), .A(n10232), .ZN(n10243) );
  NAND2_X1 U12768 ( .A1(n14819), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n10235) );
  NAND2_X1 U12769 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11543)
         );
  OAI211_X1 U12770 ( .C1(n14827), .C2(n10296), .A(n10235), .B(n11543), .ZN(
        n10242) );
  AOI21_X1 U12771 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n10237), .A(n10236), 
        .ZN(n10240) );
  INV_X1 U12772 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10238) );
  MUX2_X1 U12773 ( .A(n10238), .B(P2_REG1_REG_11__SCAN_IN), .S(n10304), .Z(
        n10239) );
  NOR2_X1 U12774 ( .A1(n10240), .A2(n10239), .ZN(n10303) );
  AOI211_X1 U12775 ( .C1(n10240), .C2(n10239), .A(n14813), .B(n10303), .ZN(
        n10241) );
  AOI211_X1 U12776 ( .C1(n14805), .C2(n10243), .A(n10242), .B(n10241), .ZN(
        n10244) );
  INV_X1 U12777 ( .A(n10244), .ZN(P2_U3225) );
  INV_X1 U12778 ( .A(n10245), .ZN(n10247) );
  OAI222_X1 U12779 ( .A1(n11970), .A2(n10247), .B1(n12280), .B2(P3_U3151), 
        .C1(n10246), .C2(n11881), .ZN(P3_U3279) );
  AOI21_X1 U12780 ( .B1(n10252), .B2(P1_REG2_REG_6__SCAN_IN), .A(n10248), .ZN(
        n10250) );
  XNOR2_X1 U12781 ( .A(n10432), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n10249) );
  AOI211_X1 U12782 ( .C1(n10250), .C2(n10249), .A(n14572), .B(n10431), .ZN(
        n10259) );
  INV_X1 U12783 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10253) );
  MUX2_X1 U12784 ( .A(n10253), .B(P1_REG1_REG_7__SCAN_IN), .S(n10432), .Z(
        n10254) );
  NOR2_X1 U12785 ( .A1(n10255), .A2(n10254), .ZN(n10425) );
  AOI211_X1 U12786 ( .C1(n10255), .C2(n10254), .A(n14576), .B(n10425), .ZN(
        n10258) );
  INV_X1 U12787 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14261) );
  NAND2_X1 U12788 ( .A1(n14582), .A2(n10432), .ZN(n10256) );
  NAND2_X1 U12789 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11025) );
  OAI211_X1 U12790 ( .C1(n14261), .C2(n14585), .A(n10256), .B(n11025), .ZN(
        n10257) );
  OR3_X1 U12791 ( .A1(n10259), .A2(n10258), .A3(n10257), .ZN(P1_U3250) );
  INV_X1 U12792 ( .A(n10260), .ZN(n10275) );
  INV_X1 U12793 ( .A(n11111), .ZN(n10552) );
  OAI222_X1 U12794 ( .A1(n13459), .A2(n10275), .B1(n10552), .B2(P2_U3088), 
        .C1(n7301), .C2(n13464), .ZN(P2_U3314) );
  NAND2_X1 U12795 ( .A1(n13780), .A2(n10153), .ZN(n10262) );
  NAND2_X1 U12796 ( .A1(n10264), .A2(n13587), .ZN(n10261) );
  NAND2_X1 U12797 ( .A1(n10262), .A2(n10261), .ZN(n10263) );
  XNOR2_X1 U12798 ( .A(n10263), .B(n13625), .ZN(n10464) );
  INV_X1 U12799 ( .A(n10463), .ZN(n11011) );
  AOI22_X1 U12800 ( .A1(n13780), .A2(n10463), .B1(n13555), .B2(n10264), .ZN(
        n10465) );
  XNOR2_X1 U12801 ( .A(n10464), .B(n10465), .ZN(n10268) );
  OAI21_X1 U12802 ( .B1(n10268), .B2(n10267), .A(n10468), .ZN(n10269) );
  NAND2_X1 U12803 ( .A1(n10269), .A2(n14395), .ZN(n10273) );
  AOI22_X1 U12804 ( .A1(n13779), .A2(n13732), .B1(n14387), .B2(n14629), .ZN(
        n14607) );
  INV_X1 U12805 ( .A(n14607), .ZN(n10271) );
  AOI22_X1 U12806 ( .A1(n10271), .A2(n14397), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10270), .ZN(n10272) );
  OAI211_X1 U12807 ( .C1(n14659), .C2(n13742), .A(n10273), .B(n10272), .ZN(
        P1_U3237) );
  INV_X1 U12808 ( .A(n11865), .ZN(n14520) );
  OAI222_X1 U12809 ( .A1(P1_U3086), .A2(n14520), .B1(n14171), .B2(n10275), 
        .C1(n10274), .C2(n14163), .ZN(P1_U3342) );
  NAND2_X1 U12810 ( .A1(n10276), .A2(n15030), .ZN(n10277) );
  OAI22_X1 U12811 ( .A1(n14913), .A2(n10277), .B1(n8829), .B2(n15017), .ZN(
        n10313) );
  INV_X1 U12812 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10395) );
  OAI22_X1 U12813 ( .A1(n12585), .A2(n10311), .B1(n15096), .B2(n10395), .ZN(
        n10278) );
  AOI21_X1 U12814 ( .B1(n10313), .B2(n15096), .A(n10278), .ZN(n10279) );
  INV_X1 U12815 ( .A(n10279), .ZN(P3_U3459) );
  INV_X1 U12816 ( .A(n10280), .ZN(n10285) );
  NAND2_X1 U12817 ( .A1(n10281), .A2(n10284), .ZN(n10282) );
  INV_X1 U12818 ( .A(n15044), .ZN(n10286) );
  INV_X1 U12819 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10289) );
  INV_X1 U12820 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10288) );
  OAI22_X1 U12821 ( .A1(n15050), .A2(n10289), .B1(n10288), .B2(n15012), .ZN(
        n10290) );
  AOI21_X1 U12822 ( .B1(n10313), .B2(n15050), .A(n10290), .ZN(n10291) );
  OAI21_X1 U12823 ( .B1(n10311), .B2(n14958), .A(n10291), .ZN(P3_U3233) );
  INV_X1 U12824 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10292) );
  OR2_X1 U12825 ( .A1(n10538), .A2(n10292), .ZN(n10294) );
  NAND2_X1 U12826 ( .A1(n10538), .A2(n10292), .ZN(n10293) );
  NAND2_X1 U12827 ( .A1(n10294), .A2(n10293), .ZN(n10300) );
  AOI21_X1 U12828 ( .B1(n10297), .B2(n10296), .A(n10295), .ZN(n10298) );
  INV_X1 U12829 ( .A(n10298), .ZN(n10299) );
  NAND2_X1 U12830 ( .A1(n10300), .A2(n10299), .ZN(n10547) );
  OAI21_X1 U12831 ( .B1(n10300), .B2(n10299), .A(n10547), .ZN(n10301) );
  AOI22_X1 U12832 ( .A1(n14819), .A2(P2_ADDR_REG_12__SCAN_IN), .B1(n14805), 
        .B2(n10301), .ZN(n10310) );
  NAND2_X1 U12833 ( .A1(n10538), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10302) );
  OAI21_X1 U12834 ( .B1(n10538), .B2(P2_REG1_REG_12__SCAN_IN), .A(n10302), 
        .ZN(n10305) );
  AOI21_X1 U12835 ( .B1(n10304), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10303), 
        .ZN(n10306) );
  OAI21_X1 U12836 ( .B1(n6624), .B2(n10306), .A(n10540), .ZN(n10308) );
  NAND2_X1 U12837 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n11581)
         );
  INV_X1 U12838 ( .A(n11581), .ZN(n10307) );
  AOI21_X1 U12839 ( .B1(n14784), .B2(n10308), .A(n10307), .ZN(n10309) );
  OAI211_X1 U12840 ( .C1(n10545), .C2(n14827), .A(n10310), .B(n10309), .ZN(
        P2_U3226) );
  OAI22_X1 U12841 ( .A1(n10311), .A2(n12638), .B1(n15081), .B2(n8821), .ZN(
        n10312) );
  AOI21_X1 U12842 ( .B1(n10313), .B2(n15081), .A(n10312), .ZN(n10314) );
  INV_X1 U12843 ( .A(n10314), .ZN(P3_U3390) );
  NAND3_X1 U12844 ( .A1(n9322), .A2(n15032), .A3(n10315), .ZN(n10316) );
  OAI211_X1 U12845 ( .C1(n10318), .C2(n9185), .A(n10317), .B(n10316), .ZN(
        n10324) );
  AND2_X1 U12846 ( .A1(n10319), .A2(n12640), .ZN(n14920) );
  INV_X1 U12847 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10445) );
  INV_X1 U12848 ( .A(n12177), .ZN(n14918) );
  AOI22_X1 U12849 ( .A1(n15036), .A2(n14916), .B1(n10320), .B2(n14918), .ZN(
        n10322) );
  NAND2_X1 U12850 ( .A1(n12170), .A2(n15033), .ZN(n10321) );
  OAI211_X1 U12851 ( .C1(n14920), .C2(n10445), .A(n10322), .B(n10321), .ZN(
        n10323) );
  AOI21_X1 U12852 ( .B1(n10324), .B2(n14914), .A(n10323), .ZN(n10325) );
  INV_X1 U12853 ( .A(n10325), .ZN(P3_U3162) );
  INV_X1 U12854 ( .A(n10326), .ZN(n10328) );
  OAI222_X1 U12855 ( .A1(n11970), .A2(n10328), .B1(n12296), .B2(P3_U3151), 
        .C1(n10327), .C2(n11881), .ZN(P3_U3278) );
  NAND2_X1 U12856 ( .A1(n14831), .A2(n13034), .ZN(n11046) );
  INV_X1 U12857 ( .A(n11046), .ZN(n10329) );
  NAND3_X1 U12858 ( .A1(n10330), .A2(n10329), .A3(n10344), .ZN(n10331) );
  NOR2_X1 U12859 ( .A1(n11515), .A2(n12791), .ZN(n12784) );
  NAND2_X1 U12860 ( .A1(n13248), .A2(n12784), .ZN(n13258) );
  INV_X1 U12861 ( .A(n13258), .ZN(n10333) );
  OAI21_X1 U12862 ( .B1(n13072), .B2(n10484), .A(n11942), .ZN(n14838) );
  INV_X1 U12863 ( .A(n14838), .ZN(n10332) );
  NAND2_X1 U12864 ( .A1(n10333), .A2(n10332), .ZN(n10342) );
  NAND2_X1 U12865 ( .A1(n7728), .A2(n10484), .ZN(n14836) );
  NAND2_X1 U12866 ( .A1(n13029), .A2(n7734), .ZN(n10337) );
  AOI21_X1 U12867 ( .B1(n10336), .B2(n13281), .A(n14838), .ZN(n10339) );
  NOR2_X1 U12868 ( .A1(n12773), .A2(n7147), .ZN(n10483) );
  NOR2_X1 U12869 ( .A1(n10339), .A2(n10483), .ZN(n14837) );
  OAI21_X1 U12870 ( .B1(n13030), .B2(n14836), .A(n14837), .ZN(n10340) );
  AOI22_X1 U12871 ( .A1(n13248), .A2(n10340), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13289), .ZN(n10341) );
  OAI211_X1 U12872 ( .C1(n14748), .C2(n13248), .A(n10342), .B(n10341), .ZN(
        P2_U3265) );
  AND3_X1 U12873 ( .A1(n10344), .A2(n14834), .A3(n10343), .ZN(n11048) );
  NAND2_X1 U12874 ( .A1(n14835), .A2(n13034), .ZN(n10345) );
  NOR2_X1 U12875 ( .A1(n14831), .A2(n10345), .ZN(n10346) );
  NAND2_X1 U12876 ( .A1(n10347), .A2(n10484), .ZN(n12807) );
  INV_X1 U12877 ( .A(n12807), .ZN(n10348) );
  OAI21_X1 U12878 ( .B1(n10348), .B2(n6735), .A(n10574), .ZN(n10349) );
  NAND2_X1 U12879 ( .A1(n10349), .A2(n13198), .ZN(n10353) );
  NAND2_X1 U12880 ( .A1(n13036), .A2(n13072), .ZN(n10351) );
  OR2_X1 U12881 ( .A1(n12773), .A2(n10575), .ZN(n10350) );
  NAND2_X1 U12882 ( .A1(n10351), .A2(n10350), .ZN(n11943) );
  INV_X1 U12883 ( .A(n11943), .ZN(n10352) );
  NAND2_X1 U12884 ( .A1(n10353), .A2(n10352), .ZN(n10814) );
  INV_X1 U12885 ( .A(n10840), .ZN(n10354) );
  OAI211_X1 U12886 ( .C1(n10355), .C2(n7033), .A(n13106), .B(n10354), .ZN(
        n10812) );
  NAND2_X1 U12887 ( .A1(n14891), .A2(n12815), .ZN(n10356) );
  NAND2_X1 U12888 ( .A1(n10812), .A2(n10356), .ZN(n10357) );
  NOR2_X1 U12889 ( .A1(n10814), .A2(n10357), .ZN(n10361) );
  XNOR2_X1 U12890 ( .A(n11942), .B(n6735), .ZN(n10816) );
  INV_X1 U12891 ( .A(n10816), .ZN(n10358) );
  INV_X1 U12892 ( .A(n10336), .ZN(n14890) );
  NAND2_X1 U12893 ( .A1(n10358), .A2(n14890), .ZN(n10360) );
  INV_X1 U12894 ( .A(n14895), .ZN(n14873) );
  NAND2_X1 U12895 ( .A1(n10358), .A2(n14873), .ZN(n10359) );
  AND3_X1 U12896 ( .A1(n10361), .A2(n10360), .A3(n10359), .ZN(n14842) );
  NAND2_X1 U12897 ( .A1(n14910), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10362) );
  OAI21_X1 U12898 ( .B1(n14910), .B2(n14842), .A(n10362), .ZN(P2_U3500) );
  OAI21_X1 U12899 ( .B1(n10365), .B2(n10364), .A(n10363), .ZN(n10369) );
  INV_X1 U12900 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10401) );
  AOI22_X1 U12901 ( .A1(n12190), .A2(n14916), .B1(n15024), .B2(n14918), .ZN(
        n10367) );
  NAND2_X1 U12902 ( .A1(n12170), .A2(n7333), .ZN(n10366) );
  OAI211_X1 U12903 ( .C1(n14920), .C2(n10401), .A(n10367), .B(n10366), .ZN(
        n10368) );
  AOI21_X1 U12904 ( .B1(n10369), .B2(n14914), .A(n10368), .ZN(n10370) );
  INV_X1 U12905 ( .A(n10370), .ZN(P3_U3177) );
  XNOR2_X1 U12906 ( .A(n10371), .B(n10372), .ZN(n14668) );
  INV_X1 U12907 ( .A(n14668), .ZN(n10386) );
  OAI21_X1 U12908 ( .B1(n10375), .B2(n10374), .A(n10373), .ZN(n10377) );
  NAND2_X1 U12909 ( .A1(n13780), .A2(n14387), .ZN(n10376) );
  OAI21_X1 U12910 ( .B1(n10871), .B2(n14385), .A(n10376), .ZN(n10477) );
  AOI21_X1 U12911 ( .B1(n10377), .B2(n14630), .A(n10477), .ZN(n10378) );
  INV_X1 U12912 ( .A(n10378), .ZN(n14666) );
  OR2_X1 U12913 ( .A1(n14616), .A2(n8301), .ZN(n10379) );
  NAND2_X1 U12914 ( .A1(n10853), .A2(n10379), .ZN(n14665) );
  INV_X1 U12915 ( .A(n14665), .ZN(n10380) );
  NAND2_X1 U12916 ( .A1(n13920), .A2(n10380), .ZN(n10383) );
  NOR2_X1 U12917 ( .A1(n14612), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10381) );
  AOI21_X1 U12918 ( .B1(n14648), .B2(P1_REG2_REG_3__SCAN_IN), .A(n10381), .ZN(
        n10382) );
  OAI211_X1 U12919 ( .C1(n8301), .C2(n14640), .A(n10383), .B(n10382), .ZN(
        n10384) );
  AOI21_X1 U12920 ( .B1(n14666), .B2(n14008), .A(n10384), .ZN(n10385) );
  OAI21_X1 U12921 ( .B1(n10386), .B2(n14016), .A(n10385), .ZN(P1_U3290) );
  NAND2_X1 U12922 ( .A1(n10387), .A2(n11320), .ZN(n10399) );
  INV_X1 U12923 ( .A(n10399), .ZN(n10392) );
  NAND2_X1 U12924 ( .A1(n10389), .A2(n10388), .ZN(n10390) );
  NAND2_X1 U12925 ( .A1(n10391), .A2(n10390), .ZN(n10400) );
  INV_X1 U12926 ( .A(n10403), .ZN(n10394) );
  INV_X1 U12927 ( .A(n14948), .ZN(n11247) );
  NAND2_X1 U12928 ( .A1(n10394), .A2(n12198), .ZN(n14937) );
  INV_X1 U12929 ( .A(n14937), .ZN(n14924) );
  INV_X1 U12930 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15261) );
  MUX2_X1 U12931 ( .A(n15261), .B(P3_REG1_REG_2__SCAN_IN), .S(n10416), .Z(
        n10398) );
  NOR2_X1 U12932 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10395), .ZN(n10396) );
  INV_X1 U12933 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15082) );
  NAND2_X1 U12934 ( .A1(n10448), .A2(n6501), .ZN(n10397) );
  OAI21_X1 U12935 ( .B1(n10398), .B2(n10397), .A(n10521), .ZN(n10412) );
  OAI22_X1 U12936 ( .A1(n14951), .A2(n14180), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10401), .ZN(n10411) );
  INV_X1 U12937 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n15029) );
  MUX2_X1 U12938 ( .A(n15029), .B(P3_REG2_REG_2__SCAN_IN), .S(n10416), .Z(
        n10408) );
  AND2_X1 U12939 ( .A1(n15207), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10405) );
  NAND2_X1 U12940 ( .A1(n10404), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10406) );
  OAI21_X1 U12941 ( .B1(n10456), .B2(n10405), .A(n10406), .ZN(n10442) );
  INV_X1 U12942 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15049) );
  NAND2_X1 U12943 ( .A1(n10407), .A2(n10408), .ZN(n10509) );
  OAI21_X1 U12944 ( .B1(n10408), .B2(n10407), .A(n10509), .ZN(n10409) );
  AND2_X1 U12945 ( .A1(n14923), .A2(n10409), .ZN(n10410) );
  AOI211_X1 U12946 ( .C1(n14924), .C2(n10412), .A(n10411), .B(n10410), .ZN(
        n10419) );
  MUX2_X1 U12947 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n12198), .Z(n10413) );
  XOR2_X1 U12948 ( .A(n10456), .B(n10413), .Z(n10452) );
  MUX2_X1 U12949 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n12198), .Z(n14926) );
  NOR2_X1 U12950 ( .A1(n14926), .A2(n15207), .ZN(n14925) );
  INV_X1 U12951 ( .A(n10456), .ZN(n10415) );
  INV_X1 U12952 ( .A(n10413), .ZN(n10414) );
  AOI22_X1 U12953 ( .A1(n10452), .A2(n14925), .B1(n10415), .B2(n10414), .ZN(
        n10502) );
  MUX2_X1 U12954 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12198), .Z(n10500) );
  XOR2_X1 U12955 ( .A(n10416), .B(n10500), .Z(n10501) );
  XNOR2_X1 U12956 ( .A(n10502), .B(n10501), .ZN(n10417) );
  NAND2_X1 U12957 ( .A1(P3_U3897), .A2(n11876), .ZN(n14943) );
  NAND2_X1 U12958 ( .A1(n10417), .A2(n14922), .ZN(n10418) );
  OAI211_X1 U12959 ( .C1(n11247), .C2(n10519), .A(n10419), .B(n10418), .ZN(
        P3_U3184) );
  INV_X1 U12960 ( .A(n10420), .ZN(n10422) );
  OAI222_X1 U12961 ( .A1(n12306), .A2(P3_U3151), .B1(n11970), .B2(n10422), 
        .C1(n10421), .C2(n11881), .ZN(P3_U3277) );
  INV_X1 U12962 ( .A(n10423), .ZN(n10553) );
  AOI22_X1 U12963 ( .A1(n14525), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n14151), .ZN(n10424) );
  OAI21_X1 U12964 ( .B1(n10553), .B2(n14171), .A(n10424), .ZN(P1_U3341) );
  AOI21_X1 U12965 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n10432), .A(n10425), .ZN(
        n10428) );
  INV_X1 U12966 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10426) );
  MUX2_X1 U12967 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10426), .S(n10734), .Z(
        n10427) );
  NAND2_X1 U12968 ( .A1(n10428), .A2(n10427), .ZN(n10728) );
  OAI21_X1 U12969 ( .B1(n10428), .B2(n10427), .A(n10728), .ZN(n10438) );
  AND2_X1 U12970 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n11268) );
  AOI21_X1 U12971 ( .B1(n14491), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n11268), .ZN(
        n10429) );
  OAI21_X1 U12972 ( .B1(n14566), .B2(n10430), .A(n10429), .ZN(n10437) );
  AOI21_X1 U12973 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n10432), .A(n10431), .ZN(
        n10435) );
  INV_X1 U12974 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10433) );
  MUX2_X1 U12975 ( .A(n10433), .B(P1_REG2_REG_8__SCAN_IN), .S(n10734), .Z(
        n10434) );
  AOI211_X1 U12976 ( .C1(n10435), .C2(n10434), .A(n14572), .B(n10733), .ZN(
        n10436) );
  AOI211_X1 U12977 ( .C1(n14558), .C2(n10438), .A(n10437), .B(n10436), .ZN(
        n10439) );
  INV_X1 U12978 ( .A(n10439), .ZN(P1_U3251) );
  INV_X1 U12979 ( .A(n10440), .ZN(n10460) );
  OAI222_X1 U12980 ( .A1(P1_U3086), .A2(n14549), .B1(n14171), .B2(n10460), 
        .C1(n10441), .C2(n14163), .ZN(P1_U3339) );
  INV_X1 U12981 ( .A(n10442), .ZN(n10444) );
  OAI21_X1 U12982 ( .B1(n10444), .B2(P3_REG2_REG_1__SCAN_IN), .A(n10443), .ZN(
        n10451) );
  OAI22_X1 U12983 ( .A1(n14951), .A2(n14179), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10445), .ZN(n10450) );
  NAND2_X1 U12984 ( .A1(n10446), .A2(n15082), .ZN(n10447) );
  AOI21_X1 U12985 ( .B1(n10448), .B2(n10447), .A(n14937), .ZN(n10449) );
  AOI211_X1 U12986 ( .C1(n14923), .C2(n10451), .A(n10450), .B(n10449), .ZN(
        n10455) );
  XNOR2_X1 U12987 ( .A(n10452), .B(n14925), .ZN(n10453) );
  NAND2_X1 U12988 ( .A1(n10453), .A2(n14922), .ZN(n10454) );
  OAI211_X1 U12989 ( .C1(n11247), .C2(n10456), .A(n10455), .B(n10454), .ZN(
        P3_U3183) );
  OAI222_X1 U12990 ( .A1(n10459), .A2(P3_U3151), .B1(n11970), .B2(n10458), 
        .C1(n10457), .C2(n11881), .ZN(P3_U3276) );
  INV_X1 U12991 ( .A(n11739), .ZN(n11737) );
  OAI222_X1 U12992 ( .A1(n13464), .A2(n10461), .B1(n11737), .B2(P2_U3088), 
        .C1(n13459), .C2(n10460), .ZN(P2_U3311) );
  OAI22_X1 U12993 ( .A1(n10847), .A2(n13627), .B1(n8301), .B2(n13629), .ZN(
        n10462) );
  XNOR2_X1 U12994 ( .A(n10462), .B(n13625), .ZN(n10866) );
  OAI22_X1 U12995 ( .A1(n10847), .A2(n11011), .B1(n8301), .B2(n13627), .ZN(
        n10865) );
  XNOR2_X1 U12996 ( .A(n10866), .B(n10865), .ZN(n10471) );
  INV_X1 U12997 ( .A(n10464), .ZN(n10466) );
  NAND2_X1 U12998 ( .A1(n10466), .A2(n10465), .ZN(n10467) );
  NAND2_X1 U12999 ( .A1(n10468), .A2(n10467), .ZN(n10470) );
  OR2_X1 U13000 ( .A1(n10470), .A2(n10471), .ZN(n10868) );
  INV_X1 U13001 ( .A(n10868), .ZN(n10469) );
  AOI211_X1 U13002 ( .C1(n10471), .C2(n10470), .A(n13751), .B(n10469), .ZN(
        n10481) );
  INV_X1 U13003 ( .A(n10472), .ZN(n10473) );
  NAND2_X1 U13004 ( .A1(n10474), .A2(n10473), .ZN(n10475) );
  NAND2_X1 U13005 ( .A1(n14398), .A2(n10476), .ZN(n10479) );
  AOI22_X1 U13006 ( .A1(n14397), .A2(n10477), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10478) );
  OAI211_X1 U13007 ( .C1(n14401), .C2(P1_REG3_REG_3__SCAN_IN), .A(n10479), .B(
        n10478), .ZN(n10480) );
  OR2_X1 U13008 ( .A1(n10481), .A2(n10480), .ZN(P1_U3218) );
  NOR2_X1 U13009 ( .A1(n10482), .A2(P2_U3088), .ZN(n11946) );
  INV_X1 U13010 ( .A(n12765), .ZN(n12744) );
  NAND2_X1 U13011 ( .A1(n13072), .A2(n7033), .ZN(n12808) );
  INV_X1 U13012 ( .A(n12808), .ZN(n12811) );
  AOI22_X1 U13013 ( .A1(n12744), .A2(n12811), .B1(n14378), .B2(n10483), .ZN(
        n10487) );
  AOI21_X1 U13014 ( .B1(n13072), .B2(n13089), .A(n12759), .ZN(n10485) );
  OAI21_X1 U13015 ( .B1(n10485), .B2(n14381), .A(n10484), .ZN(n10486) );
  OAI211_X1 U13016 ( .C1(n11946), .C2(n10488), .A(n10487), .B(n10486), .ZN(
        P2_U3204) );
  INV_X1 U13017 ( .A(n11946), .ZN(n10493) );
  OR2_X1 U13018 ( .A1(n12773), .A2(n11983), .ZN(n10491) );
  NAND2_X1 U13019 ( .A1(n13036), .A2(n13070), .ZN(n10490) );
  AND2_X1 U13020 ( .A1(n10491), .A2(n10490), .ZN(n10834) );
  OAI22_X1 U13021 ( .A1(n12776), .A2(n14844), .B1(n10834), .B2(n12751), .ZN(
        n10492) );
  AOI21_X1 U13022 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n10493), .A(n10492), .ZN(
        n10499) );
  OAI22_X1 U13023 ( .A1(n12765), .A2(n7147), .B1(n7753), .B2(n12759), .ZN(
        n10497) );
  INV_X1 U13024 ( .A(n10494), .ZN(n10496) );
  NAND3_X1 U13025 ( .A1(n10497), .A2(n10496), .A3(n10495), .ZN(n10498) );
  OAI211_X1 U13026 ( .C1(n10489), .C2(n12759), .A(n10499), .B(n10498), .ZN(
        P2_U3209) );
  MUX2_X1 U13027 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12198), .Z(n10666) );
  XNOR2_X1 U13028 ( .A(n10666), .B(n10675), .ZN(n10667) );
  MUX2_X1 U13029 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12198), .Z(n10503) );
  XNOR2_X1 U13030 ( .A(n10503), .B(n10647), .ZN(n10638) );
  INV_X1 U13031 ( .A(n10503), .ZN(n10504) );
  MUX2_X1 U13032 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12198), .Z(n10505) );
  XOR2_X1 U13033 ( .A(n10724), .B(n10505), .Z(n10708) );
  MUX2_X1 U13034 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12198), .Z(n10506) );
  XNOR2_X1 U13035 ( .A(n10506), .B(n10634), .ZN(n10622) );
  INV_X1 U13036 ( .A(n10506), .ZN(n10507) );
  XOR2_X1 U13037 ( .A(n10667), .B(n10668), .Z(n10537) );
  NOR2_X1 U13038 ( .A1(n11247), .A2(n10675), .ZN(n10535) );
  NAND2_X1 U13039 ( .A1(n10519), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U13040 ( .A1(n10509), .A2(n10508), .ZN(n10510) );
  NAND2_X1 U13041 ( .A1(n10510), .A2(n10522), .ZN(n10710) );
  OAI21_X1 U13042 ( .B1(n10510), .B2(n10522), .A(n10710), .ZN(n10639) );
  INV_X1 U13043 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10640) );
  XNOR2_X1 U13044 ( .A(n10724), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n10709) );
  NAND2_X1 U13045 ( .A1(n10525), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10511) );
  NAND2_X1 U13046 ( .A1(n10512), .A2(n10526), .ZN(n10516) );
  OAI21_X1 U13047 ( .B1(n10512), .B2(n10526), .A(n10516), .ZN(n10625) );
  INV_X1 U13048 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n14997) );
  NAND2_X1 U13049 ( .A1(n10623), .A2(n10516), .ZN(n10514) );
  INV_X1 U13050 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10513) );
  MUX2_X1 U13051 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n10513), .S(n10675), .Z(
        n10515) );
  NAND2_X1 U13052 ( .A1(n10514), .A2(n10515), .ZN(n10663) );
  INV_X1 U13053 ( .A(n10515), .ZN(n10517) );
  NAND3_X1 U13054 ( .A1(n10623), .A2(n10517), .A3(n10516), .ZN(n10518) );
  AOI21_X1 U13055 ( .B1(n10663), .B2(n10518), .A(n14940), .ZN(n10534) );
  NAND2_X1 U13056 ( .A1(n10519), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10520) );
  NAND2_X1 U13057 ( .A1(n10521), .A2(n10520), .ZN(n10523) );
  NAND2_X1 U13058 ( .A1(n10523), .A2(n10522), .ZN(n10716) );
  OAI21_X1 U13059 ( .B1(n10523), .B2(n10522), .A(n10716), .ZN(n10641) );
  INV_X1 U13060 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15085) );
  NAND2_X1 U13061 ( .A1(n10717), .A2(n10716), .ZN(n10524) );
  XNOR2_X1 U13062 ( .A(n10724), .B(P3_REG1_REG_4__SCAN_IN), .ZN(n10715) );
  INV_X1 U13063 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15089) );
  NAND2_X1 U13064 ( .A1(n10629), .A2(n10529), .ZN(n10527) );
  INV_X1 U13065 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15091) );
  MUX2_X1 U13066 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n15091), .S(n10675), .Z(
        n10528) );
  NAND2_X1 U13067 ( .A1(n10527), .A2(n10528), .ZN(n10677) );
  INV_X1 U13068 ( .A(n10528), .ZN(n10530) );
  NAND3_X1 U13069 ( .A1(n10629), .A2(n10530), .A3(n10529), .ZN(n10531) );
  AOI21_X1 U13070 ( .B1(n10677), .B2(n10531), .A(n14937), .ZN(n10533) );
  NAND2_X1 U13071 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n10949) );
  OAI21_X1 U13072 ( .B1(n14951), .B2(n14191), .A(n10949), .ZN(n10532) );
  NOR4_X1 U13073 ( .A1(n10535), .A2(n10534), .A3(n10533), .A4(n10532), .ZN(
        n10536) );
  OAI21_X1 U13074 ( .B1(n10537), .B2(n14943), .A(n10536), .ZN(P3_U3188) );
  XNOR2_X1 U13075 ( .A(n11111), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n10542) );
  OR2_X1 U13076 ( .A1(n10538), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10539) );
  AOI211_X1 U13077 ( .C1(n10542), .C2(n10541), .A(n11107), .B(n14813), .ZN(
        n10544) );
  NOR2_X1 U13078 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11693), .ZN(n10543) );
  NOR2_X1 U13079 ( .A1(n10544), .A2(n10543), .ZN(n10551) );
  NAND2_X1 U13080 ( .A1(n10545), .A2(n10292), .ZN(n10546) );
  NAND2_X1 U13081 ( .A1(n10547), .A2(n10546), .ZN(n11113) );
  INV_X1 U13082 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10548) );
  MUX2_X1 U13083 ( .A(n10548), .B(P2_REG2_REG_13__SCAN_IN), .S(n11111), .Z(
        n11112) );
  XOR2_X1 U13084 ( .A(n11113), .B(n11112), .Z(n10549) );
  AOI22_X1 U13085 ( .A1(n14819), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(n14805), 
        .B2(n10549), .ZN(n10550) );
  OAI211_X1 U13086 ( .C1(n10552), .C2(n14827), .A(n10551), .B(n10550), .ZN(
        P2_U3227) );
  INV_X1 U13087 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10555) );
  INV_X1 U13088 ( .A(n14803), .ZN(n10554) );
  OAI222_X1 U13089 ( .A1(n13464), .A2(n10555), .B1(n10554), .B2(P2_U3088), 
        .C1(n13459), .C2(n10553), .ZN(P2_U3313) );
  INV_X1 U13090 ( .A(n10556), .ZN(n10560) );
  INV_X1 U13091 ( .A(n12006), .ZN(n11999) );
  OAI222_X1 U13092 ( .A1(n13459), .A2(n10560), .B1(n11999), .B2(P2_U3088), 
        .C1(n15219), .C2(n13464), .ZN(P2_U3310) );
  INV_X1 U13093 ( .A(n10557), .ZN(n10590) );
  INV_X1 U13094 ( .A(n11441), .ZN(n11436) );
  OAI222_X1 U13095 ( .A1(n13459), .A2(n10590), .B1(n11436), .B2(P2_U3088), 
        .C1(n10558), .C2(n13464), .ZN(P2_U3312) );
  INV_X1 U13096 ( .A(n13849), .ZN(n14565) );
  OAI222_X1 U13097 ( .A1(P1_U3086), .A2(n14565), .B1(n14171), .B2(n10560), 
        .C1(n10559), .C2(n14163), .ZN(P1_U3338) );
  INV_X1 U13098 ( .A(n12784), .ZN(n10561) );
  NAND2_X1 U13099 ( .A1(n10336), .A2(n10561), .ZN(n10562) );
  INV_X1 U13100 ( .A(n11942), .ZN(n10563) );
  OAI22_X1 U13101 ( .A1(n12991), .A2(n10563), .B1(n13070), .B2(n12815), .ZN(
        n10838) );
  NAND2_X1 U13102 ( .A1(n14844), .A2(n10575), .ZN(n10564) );
  NAND2_X1 U13103 ( .A1(n10565), .A2(n10564), .ZN(n10612) );
  OR2_X1 U13104 ( .A1(n12833), .A2(n13068), .ZN(n10567) );
  XNOR2_X1 U13105 ( .A(n12841), .B(n13066), .ZN(n12999) );
  XNOR2_X1 U13106 ( .A(n10592), .B(n12999), .ZN(n14866) );
  INV_X1 U13107 ( .A(n12836), .ZN(n14860) );
  NAND2_X1 U13108 ( .A1(n14844), .A2(n10840), .ZN(n10839) );
  INV_X1 U13109 ( .A(n10606), .ZN(n10568) );
  AOI211_X1 U13110 ( .C1(n12841), .C2(n10771), .A(n13089), .B(n10568), .ZN(
        n14867) );
  INV_X1 U13111 ( .A(n10569), .ZN(n10570) );
  INV_X1 U13112 ( .A(n12841), .ZN(n14869) );
  INV_X1 U13113 ( .A(n12704), .ZN(n10571) );
  OAI22_X1 U13114 ( .A1(n13293), .A2(n14869), .B1(n10571), .B2(n13226), .ZN(
        n10572) );
  AOI21_X1 U13115 ( .B1(n13288), .B2(n14867), .A(n10572), .ZN(n10588) );
  NAND2_X1 U13116 ( .A1(n7147), .A2(n12815), .ZN(n10573) );
  NAND2_X1 U13117 ( .A1(n10575), .A2(n12824), .ZN(n10576) );
  NAND2_X1 U13118 ( .A1(n12833), .A2(n11983), .ZN(n10578) );
  NAND2_X1 U13119 ( .A1(n10579), .A2(n10578), .ZN(n10766) );
  NAND2_X1 U13120 ( .A1(n10766), .A2(n12996), .ZN(n10581) );
  NAND2_X1 U13121 ( .A1(n12836), .A2(n6635), .ZN(n10580) );
  XNOR2_X1 U13122 ( .A(n10597), .B(n12999), .ZN(n10585) );
  OR2_X1 U13123 ( .A1(n12773), .A2(n10800), .ZN(n10583) );
  NAND2_X1 U13124 ( .A1(n13036), .A2(n13067), .ZN(n10582) );
  AND2_X1 U13125 ( .A1(n10583), .A2(n10582), .ZN(n12702) );
  INV_X1 U13126 ( .A(n12702), .ZN(n10584) );
  AOI21_X1 U13127 ( .B1(n10585), .B2(n13198), .A(n10584), .ZN(n14865) );
  MUX2_X1 U13128 ( .A(n10586), .B(n14865), .S(n13248), .Z(n10587) );
  OAI211_X1 U13129 ( .C1(n13238), .C2(n14866), .A(n10588), .B(n10587), .ZN(
        P2_U3260) );
  OAI222_X1 U13130 ( .A1(P1_U3086), .A2(n13840), .B1(n14171), .B2(n10590), 
        .C1(n10589), .C2(n14163), .ZN(P1_U3340) );
  INV_X1 U13131 ( .A(n12999), .ZN(n10591) );
  NAND2_X1 U13132 ( .A1(n10592), .A2(n10591), .ZN(n10594) );
  OR2_X1 U13133 ( .A1(n12841), .A2(n13066), .ZN(n10593) );
  NAND2_X1 U13134 ( .A1(n12849), .A2(n10800), .ZN(n10962) );
  NAND2_X1 U13135 ( .A1(n10962), .A2(n10595), .ZN(n12998) );
  XNOR2_X1 U13136 ( .A(n10956), .B(n12998), .ZN(n11155) );
  INV_X1 U13137 ( .A(n13066), .ZN(n10767) );
  AND2_X1 U13138 ( .A1(n12841), .A2(n10767), .ZN(n10596) );
  OR2_X1 U13139 ( .A1(n12841), .A2(n10767), .ZN(n10598) );
  NAND2_X1 U13140 ( .A1(n10599), .A2(n12998), .ZN(n10600) );
  NAND2_X1 U13141 ( .A1(n10963), .A2(n10600), .ZN(n10603) );
  NAND2_X1 U13142 ( .A1(n13036), .A2(n13066), .ZN(n10602) );
  INV_X1 U13143 ( .A(n13064), .ZN(n10964) );
  OR2_X1 U13144 ( .A1(n12773), .A2(n10964), .ZN(n10601) );
  NAND2_X1 U13145 ( .A1(n10602), .A2(n10601), .ZN(n10905) );
  AOI21_X1 U13146 ( .B1(n10603), .B2(n13198), .A(n10905), .ZN(n10605) );
  NAND2_X1 U13147 ( .A1(n11155), .A2(n14890), .ZN(n10604) );
  NAND2_X1 U13148 ( .A1(n10605), .A2(n10604), .ZN(n11156) );
  INV_X1 U13149 ( .A(n14891), .ZN(n14876) );
  AOI211_X1 U13150 ( .C1(n12849), .C2(n10606), .A(n13089), .B(n11283), .ZN(
        n11160) );
  INV_X1 U13151 ( .A(n11160), .ZN(n10607) );
  OAI21_X1 U13152 ( .B1(n6657), .B2(n14876), .A(n10607), .ZN(n10608) );
  AOI211_X1 U13153 ( .C1(n14873), .C2(n11155), .A(n11156), .B(n10608), .ZN(
        n15280) );
  OR2_X1 U13154 ( .A1(n15280), .A2(n14910), .ZN(n10609) );
  OAI21_X1 U13155 ( .B1(n14912), .B2(n10610), .A(n10609), .ZN(P2_U3505) );
  XNOR2_X1 U13156 ( .A(n10612), .B(n10611), .ZN(n14852) );
  INV_X1 U13157 ( .A(n13293), .ZN(n13230) );
  AOI211_X1 U13158 ( .C1(n12833), .C2(n10839), .A(n13231), .B(n10772), .ZN(
        n14855) );
  AOI22_X1 U13159 ( .A1(n13230), .A2(n12833), .B1(n13288), .B2(n14855), .ZN(
        n10620) );
  INV_X1 U13160 ( .A(n14853), .ZN(n10615) );
  XNOR2_X1 U13161 ( .A(n10613), .B(n12994), .ZN(n10614) );
  NOR2_X1 U13162 ( .A1(n10614), .A2(n13281), .ZN(n14857) );
  AOI211_X1 U13163 ( .C1(n13289), .C2(n10616), .A(n10615), .B(n14857), .ZN(
        n10617) );
  MUX2_X1 U13164 ( .A(n10618), .B(n10617), .S(n13248), .Z(n10619) );
  OAI211_X1 U13165 ( .C1(n13238), .C2(n14852), .A(n10620), .B(n10619), .ZN(
        P2_U3262) );
  XOR2_X1 U13166 ( .A(n10622), .B(n10621), .Z(n10636) );
  INV_X1 U13167 ( .A(n10623), .ZN(n10624) );
  AOI21_X1 U13168 ( .B1(n14997), .B2(n10625), .A(n10624), .ZN(n10632) );
  NOR2_X1 U13169 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10626), .ZN(n10917) );
  NAND2_X1 U13170 ( .A1(n10627), .A2(n15089), .ZN(n10628) );
  AOI21_X1 U13171 ( .B1(n10629), .B2(n10628), .A(n14937), .ZN(n10630) );
  AOI211_X1 U13172 ( .C1(n14921), .C2(P3_ADDR_REG_5__SCAN_IN), .A(n10917), .B(
        n10630), .ZN(n10631) );
  OAI21_X1 U13173 ( .B1(n10632), .B2(n14940), .A(n10631), .ZN(n10633) );
  AOI21_X1 U13174 ( .B1(n10634), .B2(n14948), .A(n10633), .ZN(n10635) );
  OAI21_X1 U13175 ( .B1(n10636), .B2(n14943), .A(n10635), .ZN(P3_U3187) );
  XOR2_X1 U13176 ( .A(n10638), .B(n10637), .Z(n10649) );
  AOI21_X1 U13177 ( .B1(n10640), .B2(n10639), .A(n6989), .ZN(n10645) );
  NOR2_X1 U13178 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n8831), .ZN(n10654) );
  NAND2_X1 U13179 ( .A1(n10641), .A2(n15085), .ZN(n10642) );
  AOI21_X1 U13180 ( .B1(n10717), .B2(n10642), .A(n14937), .ZN(n10643) );
  AOI211_X1 U13181 ( .C1(n14921), .C2(P3_ADDR_REG_3__SCAN_IN), .A(n10654), .B(
        n10643), .ZN(n10644) );
  OAI21_X1 U13182 ( .B1(n10645), .B2(n14940), .A(n10644), .ZN(n10646) );
  AOI21_X1 U13183 ( .B1(n10647), .B2(n14948), .A(n10646), .ZN(n10648) );
  OAI21_X1 U13184 ( .B1(n10649), .B2(n14943), .A(n10648), .ZN(P3_U3185) );
  AOI211_X1 U13185 ( .C1(n10651), .C2(n10650), .A(n12153), .B(n6619), .ZN(
        n10652) );
  INV_X1 U13186 ( .A(n10652), .ZN(n10657) );
  INV_X1 U13187 ( .A(n12170), .ZN(n12141) );
  OAI22_X1 U13188 ( .A1(n14988), .A2(n12172), .B1(n12141), .B2(n10786), .ZN(
        n10653) );
  AOI211_X1 U13189 ( .C1(n10655), .C2(n14918), .A(n10654), .B(n10653), .ZN(
        n10656) );
  OAI211_X1 U13190 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12161), .A(n10657), .B(
        n10656), .ZN(P3_U3158) );
  INV_X1 U13191 ( .A(n10658), .ZN(n10660) );
  OAI222_X1 U13192 ( .A1(n10661), .A2(P3_U3151), .B1(n11970), .B2(n10660), 
        .C1(n10659), .C2(n11881), .ZN(P3_U3275) );
  NAND2_X1 U13193 ( .A1(n10675), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10662) );
  NAND2_X1 U13194 ( .A1(n10663), .A2(n10662), .ZN(n10664) );
  INV_X1 U13195 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n14976) );
  AOI21_X1 U13196 ( .B1(n10665), .B2(n14976), .A(n11055), .ZN(n10686) );
  OAI22_X1 U13197 ( .A1(n10668), .A2(n10667), .B1(n10666), .B2(n10675), .ZN(
        n10670) );
  MUX2_X1 U13198 ( .A(n14976), .B(n15098), .S(n12198), .Z(n11060) );
  XOR2_X1 U13199 ( .A(n11059), .B(n11060), .Z(n10669) );
  NAND2_X1 U13200 ( .A1(n10669), .A2(n10670), .ZN(n11061) );
  OAI21_X1 U13201 ( .B1(n10670), .B2(n10669), .A(n11061), .ZN(n10671) );
  NAND2_X1 U13202 ( .A1(n10671), .A2(n14922), .ZN(n10685) );
  INV_X1 U13203 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n10674) );
  INV_X1 U13204 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n10672) );
  NOR2_X1 U13205 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10672), .ZN(n11150) );
  INV_X1 U13206 ( .A(n11150), .ZN(n10673) );
  OAI21_X1 U13207 ( .B1(n14951), .B2(n10674), .A(n10673), .ZN(n10683) );
  NAND2_X1 U13208 ( .A1(n10675), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10676) );
  NAND2_X1 U13209 ( .A1(n10677), .A2(n10676), .ZN(n10679) );
  AND2_X1 U13210 ( .A1(n10679), .A2(n10678), .ZN(n11076) );
  INV_X1 U13211 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15098) );
  AOI21_X1 U13212 ( .B1(n10680), .B2(n15098), .A(n11075), .ZN(n10681) );
  NOR2_X1 U13213 ( .A1(n10681), .A2(n14937), .ZN(n10682) );
  AOI211_X1 U13214 ( .C1(n14948), .C2(n11059), .A(n10683), .B(n10682), .ZN(
        n10684) );
  OAI211_X1 U13215 ( .C1(n10686), .C2(n14940), .A(n10685), .B(n10684), .ZN(
        P3_U3189) );
  XNOR2_X1 U13216 ( .A(n10688), .B(n10691), .ZN(n14701) );
  INV_X1 U13217 ( .A(n14701), .ZN(n10703) );
  INV_X1 U13218 ( .A(n10689), .ZN(n10690) );
  INV_X1 U13219 ( .A(n11257), .ZN(n14699) );
  OAI211_X1 U13220 ( .C1(n10690), .C2(n14699), .A(n14617), .B(n10939), .ZN(
        n14697) );
  AOI21_X1 U13221 ( .B1(n10692), .B2(n10691), .A(n14608), .ZN(n10697) );
  NAND2_X1 U13222 ( .A1(n13775), .A2(n14387), .ZN(n10694) );
  NAND2_X1 U13223 ( .A1(n13773), .A2(n13732), .ZN(n10693) );
  AND2_X1 U13224 ( .A1(n10694), .A2(n10693), .ZN(n11266) );
  INV_X1 U13225 ( .A(n11266), .ZN(n10695) );
  AOI21_X1 U13226 ( .B1(n10697), .B2(n10696), .A(n10695), .ZN(n14698) );
  OAI21_X1 U13227 ( .B1(n14023), .B2(n14697), .A(n14698), .ZN(n10698) );
  NAND2_X1 U13228 ( .A1(n10698), .A2(n14008), .ZN(n10702) );
  INV_X1 U13229 ( .A(n11269), .ZN(n10699) );
  OAI22_X1 U13230 ( .A1(n14008), .A2(n10433), .B1(n10699), .B2(n14612), .ZN(
        n10700) );
  AOI21_X1 U13231 ( .B1(n14409), .B2(n11257), .A(n10700), .ZN(n10701) );
  OAI211_X1 U13232 ( .C1(n14016), .C2(n10703), .A(n10702), .B(n10701), .ZN(
        P1_U3285) );
  INV_X1 U13233 ( .A(P3_U3897), .ZN(n12191) );
  NAND2_X1 U13234 ( .A1(n12191), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10704) );
  OAI21_X1 U13235 ( .B1(n10705), .B2(n12191), .A(n10704), .ZN(P3_U3521) );
  NAND2_X1 U13236 ( .A1(n12191), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(n10706) );
  OAI21_X1 U13237 ( .B1(n14332), .B2(n12191), .A(n10706), .ZN(P3_U3522) );
  XOR2_X1 U13238 ( .A(n10708), .B(n10707), .Z(n10726) );
  INV_X1 U13239 ( .A(n10709), .ZN(n10711) );
  NAND3_X1 U13240 ( .A1(n10712), .A2(n10711), .A3(n10710), .ZN(n10713) );
  AOI21_X1 U13241 ( .B1(n10714), .B2(n10713), .A(n14940), .ZN(n10723) );
  AND2_X1 U13242 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10746) );
  NAND3_X1 U13243 ( .A1(n10717), .A2(n7055), .A3(n10716), .ZN(n10718) );
  AOI21_X1 U13244 ( .B1(n10719), .B2(n10718), .A(n14937), .ZN(n10720) );
  AOI211_X1 U13245 ( .C1(n14921), .C2(P3_ADDR_REG_4__SCAN_IN), .A(n10746), .B(
        n10720), .ZN(n10721) );
  INV_X1 U13246 ( .A(n10721), .ZN(n10722) );
  AOI211_X1 U13247 ( .C1(n14948), .C2(n10724), .A(n10723), .B(n10722), .ZN(
        n10725) );
  OAI21_X1 U13248 ( .B1(n10726), .B2(n14943), .A(n10725), .ZN(P3_U3186) );
  INV_X1 U13249 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10727) );
  MUX2_X1 U13250 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10727), .S(n10987), .Z(
        n10730) );
  OAI21_X1 U13251 ( .B1(n10730), .B2(n10729), .A(n10986), .ZN(n10739) );
  NAND2_X1 U13252 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11335) );
  NAND2_X1 U13253 ( .A1(n14491), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n10731) );
  OAI211_X1 U13254 ( .C1(n14566), .C2(n10732), .A(n11335), .B(n10731), .ZN(
        n10738) );
  AOI21_X1 U13255 ( .B1(n10734), .B2(P1_REG2_REG_8__SCAN_IN), .A(n10733), .ZN(
        n10736) );
  XNOR2_X1 U13256 ( .A(n10987), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n10735) );
  NOR2_X1 U13257 ( .A1(n10736), .A2(n10735), .ZN(n10982) );
  AOI211_X1 U13258 ( .C1(n10736), .C2(n10735), .A(n14572), .B(n10982), .ZN(
        n10737) );
  AOI211_X1 U13259 ( .C1(n14558), .C2(n10739), .A(n10738), .B(n10737), .ZN(
        n10740) );
  INV_X1 U13260 ( .A(n10740), .ZN(P1_U3252) );
  OAI21_X1 U13261 ( .B1(n10743), .B2(n10742), .A(n10741), .ZN(n10744) );
  NAND2_X1 U13262 ( .A1(n10744), .A2(n14914), .ZN(n10748) );
  OAI22_X1 U13263 ( .A1(n15005), .A2(n12172), .B1(n12141), .B2(n15018), .ZN(
        n10745) );
  AOI211_X1 U13264 ( .C1(n14999), .C2(n14918), .A(n10746), .B(n10745), .ZN(
        n10747) );
  OAI211_X1 U13265 ( .C1(n15013), .C2(n12161), .A(n10748), .B(n10747), .ZN(
        P3_U3170) );
  INV_X1 U13266 ( .A(n12002), .ZN(n14826) );
  OAI222_X1 U13267 ( .A1(n13459), .A2(n10778), .B1(n14826), .B2(P2_U3088), 
        .C1(n10749), .C2(n13464), .ZN(P2_U3309) );
  XNOR2_X1 U13268 ( .A(n10752), .B(n10751), .ZN(n14689) );
  XNOR2_X1 U13269 ( .A(n10754), .B(n10753), .ZN(n10757) );
  NAND2_X1 U13270 ( .A1(n13776), .A2(n14387), .ZN(n10756) );
  NAND2_X1 U13271 ( .A1(n13774), .A2(n13732), .ZN(n10755) );
  AND2_X1 U13272 ( .A1(n10756), .A2(n10755), .ZN(n11027) );
  OAI21_X1 U13273 ( .B1(n10757), .B2(n14608), .A(n11027), .ZN(n14694) );
  NAND2_X1 U13274 ( .A1(n14694), .A2(n14008), .ZN(n10763) );
  XNOR2_X1 U13275 ( .A(n14598), .B(n11029), .ZN(n10758) );
  NAND2_X1 U13276 ( .A1(n10758), .A2(n14617), .ZN(n14691) );
  INV_X1 U13277 ( .A(n14691), .ZN(n10761) );
  INV_X2 U13278 ( .A(n14008), .ZN(n14638) );
  INV_X1 U13279 ( .A(n14612), .ZN(n14637) );
  AOI22_X1 U13280 ( .A1(n14638), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n11024), 
        .B2(n14637), .ZN(n10759) );
  OAI21_X1 U13281 ( .B1(n14692), .B2(n14640), .A(n10759), .ZN(n10760) );
  AOI21_X1 U13282 ( .B1(n10761), .B2(n14644), .A(n10760), .ZN(n10762) );
  OAI211_X1 U13283 ( .C1(n14016), .C2(n14689), .A(n10763), .B(n10762), .ZN(
        P1_U3286) );
  XNOR2_X1 U13284 ( .A(n10764), .B(n10765), .ZN(n14863) );
  XNOR2_X1 U13285 ( .A(n10766), .B(n10765), .ZN(n10770) );
  OR2_X1 U13286 ( .A1(n12773), .A2(n10767), .ZN(n10769) );
  NAND2_X1 U13287 ( .A1(n13036), .A2(n13068), .ZN(n10768) );
  AND2_X1 U13288 ( .A1(n10769), .A2(n10768), .ZN(n11981) );
  OAI21_X1 U13289 ( .B1(n10770), .B2(n13281), .A(n11981), .ZN(n14862) );
  MUX2_X1 U13290 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n14862), .S(n13248), .Z(
        n10775) );
  INV_X1 U13291 ( .A(n13288), .ZN(n13184) );
  OAI211_X1 U13292 ( .C1(n14860), .C2(n10772), .A(n13106), .B(n10771), .ZN(
        n14858) );
  AOI22_X1 U13293 ( .A1(n13230), .A2(n12836), .B1(n13289), .B2(n11990), .ZN(
        n10773) );
  OAI21_X1 U13294 ( .B1(n13184), .B2(n14858), .A(n10773), .ZN(n10774) );
  AOI211_X1 U13295 ( .C1(n14863), .C2(n13295), .A(n10775), .B(n10774), .ZN(
        n10776) );
  INV_X1 U13296 ( .A(n10776), .ZN(P2_U3261) );
  INV_X1 U13297 ( .A(n14581), .ZN(n13850) );
  OAI222_X1 U13298 ( .A1(P1_U3086), .A2(n13850), .B1(n14166), .B2(n10778), 
        .C1(n10777), .C2(n14163), .ZN(P1_U3337) );
  OR2_X1 U13299 ( .A1(n10780), .A2(n10779), .ZN(n10781) );
  NAND2_X1 U13300 ( .A1(n10782), .A2(n10781), .ZN(n15062) );
  INV_X1 U13301 ( .A(n15062), .ZN(n10794) );
  OR2_X1 U13302 ( .A1(n15044), .A2(n10881), .ZN(n15026) );
  INV_X1 U13303 ( .A(n15026), .ZN(n14993) );
  NAND2_X1 U13304 ( .A1(n15050), .A2(n14993), .ZN(n11204) );
  OAI211_X1 U13305 ( .C1(n10785), .C2(n10784), .A(n10783), .B(n15039), .ZN(
        n10789) );
  INV_X1 U13306 ( .A(n15043), .ZN(n11098) );
  OAI22_X1 U13307 ( .A1(n14988), .A2(n15017), .B1(n10786), .B2(n15019), .ZN(
        n10787) );
  AOI21_X1 U13308 ( .B1(n15062), .B2(n11098), .A(n10787), .ZN(n10788) );
  NAND2_X1 U13309 ( .A1(n10789), .A2(n10788), .ZN(n15060) );
  MUX2_X1 U13310 ( .A(n15060), .B(P3_REG2_REG_3__SCAN_IN), .S(n14334), .Z(
        n10790) );
  INV_X1 U13311 ( .A(n10790), .ZN(n10793) );
  NOR2_X1 U13312 ( .A1(n10791), .A2(n15030), .ZN(n15061) );
  INV_X2 U13313 ( .A(n15012), .ZN(n15046) );
  AOI22_X1 U13314 ( .A1(n15061), .A2(n15000), .B1(n15046), .B2(n8831), .ZN(
        n10792) );
  OAI211_X1 U13315 ( .C1(n10794), .C2(n11204), .A(n10793), .B(n10792), .ZN(
        P3_U3230) );
  INV_X1 U13316 ( .A(n12853), .ZN(n14877) );
  INV_X1 U13317 ( .A(n10797), .ZN(n10798) );
  AOI21_X1 U13318 ( .B1(n10796), .B2(n10798), .A(n12759), .ZN(n10803) );
  NOR3_X1 U13319 ( .A1(n12765), .A2(n10800), .A3(n10799), .ZN(n10802) );
  OAI21_X1 U13320 ( .B1(n10803), .B2(n10802), .A(n10801), .ZN(n10808) );
  INV_X1 U13321 ( .A(n13063), .ZN(n10967) );
  OR2_X1 U13322 ( .A1(n12773), .A2(n10967), .ZN(n10805) );
  NAND2_X1 U13323 ( .A1(n13036), .A2(n13065), .ZN(n10804) );
  AND2_X1 U13324 ( .A1(n10805), .A2(n10804), .ZN(n11287) );
  OAI22_X1 U13325 ( .A1(n12751), .A2(n11287), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7844), .ZN(n10806) );
  AOI21_X1 U13326 ( .B1(n11284), .B2(n12770), .A(n10806), .ZN(n10807) );
  OAI211_X1 U13327 ( .C1(n14877), .C2(n12776), .A(n10808), .B(n10807), .ZN(
        P2_U3185) );
  INV_X1 U13328 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10809) );
  INV_X1 U13329 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11945) );
  OAI22_X1 U13330 ( .A1(n13248), .A2(n10809), .B1(n11945), .B2(n13226), .ZN(
        n10810) );
  AOI21_X1 U13331 ( .B1(n13230), .B2(n12815), .A(n10810), .ZN(n10811) );
  OAI21_X1 U13332 ( .B1(n13184), .B2(n10812), .A(n10811), .ZN(n10813) );
  AOI21_X1 U13333 ( .B1(n13248), .B2(n10814), .A(n10813), .ZN(n10815) );
  OAI21_X1 U13334 ( .B1(n13238), .B2(n10816), .A(n10815), .ZN(P2_U3264) );
  XNOR2_X1 U13335 ( .A(n10818), .B(n10819), .ZN(n10824) );
  XNOR2_X1 U13336 ( .A(n10820), .B(n10819), .ZN(n10822) );
  NAND2_X1 U13337 ( .A1(n13776), .A2(n13732), .ZN(n10821) );
  OAI21_X1 U13338 ( .B1(n10871), .B2(n14633), .A(n10821), .ZN(n10896) );
  AOI21_X1 U13339 ( .B1(n10822), .B2(n14630), .A(n10896), .ZN(n10823) );
  OAI21_X1 U13340 ( .B1(n10824), .B2(n14690), .A(n10823), .ZN(n14677) );
  INV_X1 U13341 ( .A(n14677), .ZN(n10832) );
  INV_X1 U13342 ( .A(n10824), .ZN(n14679) );
  NOR2_X1 U13343 ( .A1(n14638), .A2(n10825), .ZN(n14645) );
  INV_X1 U13344 ( .A(n10901), .ZN(n14674) );
  INV_X1 U13345 ( .A(n10854), .ZN(n10827) );
  INV_X1 U13346 ( .A(n14600), .ZN(n10826) );
  OAI21_X1 U13347 ( .B1(n14674), .B2(n10827), .A(n10826), .ZN(n14676) );
  INV_X1 U13348 ( .A(n13920), .ZN(n11935) );
  AOI22_X1 U13349 ( .A1(n14638), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n10895), 
        .B2(n14637), .ZN(n10829) );
  NAND2_X1 U13350 ( .A1(n14409), .A2(n10901), .ZN(n10828) );
  OAI211_X1 U13351 ( .C1(n14676), .C2(n11935), .A(n10829), .B(n10828), .ZN(
        n10830) );
  AOI21_X1 U13352 ( .B1(n14679), .B2(n14645), .A(n10830), .ZN(n10831) );
  OAI21_X1 U13353 ( .B1(n10832), .B2(n14638), .A(n10831), .ZN(P1_U3288) );
  XNOR2_X1 U13354 ( .A(n12992), .B(n10833), .ZN(n10836) );
  INV_X1 U13355 ( .A(n10834), .ZN(n10835) );
  AOI21_X1 U13356 ( .B1(n10836), .B2(n13198), .A(n10835), .ZN(n14845) );
  XNOR2_X1 U13357 ( .A(n10837), .B(n10838), .ZN(n14849) );
  OAI211_X1 U13358 ( .C1(n14844), .C2(n10840), .A(n13106), .B(n10839), .ZN(
        n14843) );
  AOI22_X1 U13359 ( .A1(n13298), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n13289), .ZN(n10842) );
  NAND2_X1 U13360 ( .A1(n13230), .A2(n12824), .ZN(n10841) );
  OAI211_X1 U13361 ( .C1(n13184), .C2(n14843), .A(n10842), .B(n10841), .ZN(
        n10843) );
  AOI21_X1 U13362 ( .B1(n13295), .B2(n14849), .A(n10843), .ZN(n10844) );
  OAI21_X1 U13363 ( .B1(n13298), .B2(n14845), .A(n10844), .ZN(P2_U3263) );
  XNOR2_X1 U13364 ( .A(n10845), .B(n10851), .ZN(n10849) );
  NAND2_X1 U13365 ( .A1(n13777), .A2(n13732), .ZN(n10846) );
  OAI21_X1 U13366 ( .B1(n10847), .B2(n14633), .A(n10846), .ZN(n10862) );
  INV_X1 U13367 ( .A(n10862), .ZN(n10848) );
  OAI21_X1 U13368 ( .B1(n10849), .B2(n14608), .A(n10848), .ZN(n14671) );
  INV_X1 U13369 ( .A(n14671), .ZN(n10860) );
  XNOR2_X1 U13370 ( .A(n10852), .B(n10851), .ZN(n14673) );
  INV_X1 U13371 ( .A(n14016), .ZN(n14419) );
  INV_X1 U13372 ( .A(n10853), .ZN(n10855) );
  OAI211_X1 U13373 ( .C1(n10855), .C2(n14670), .A(n14617), .B(n10854), .ZN(
        n14669) );
  NAND2_X1 U13374 ( .A1(n14409), .A2(n10876), .ZN(n10857) );
  AOI22_X1 U13375 ( .A1(n14638), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n10861), 
        .B2(n14637), .ZN(n10856) );
  OAI211_X1 U13376 ( .C1(n14669), .C2(n14011), .A(n10857), .B(n10856), .ZN(
        n10858) );
  AOI21_X1 U13377 ( .B1(n14673), .B2(n14419), .A(n10858), .ZN(n10859) );
  OAI21_X1 U13378 ( .B1(n10860), .B2(n14638), .A(n10859), .ZN(P1_U3289) );
  INV_X1 U13379 ( .A(n10861), .ZN(n10864) );
  NAND2_X1 U13380 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13812) );
  NAND2_X1 U13381 ( .A1(n14397), .A2(n10862), .ZN(n10863) );
  OAI211_X1 U13382 ( .C1(n14401), .C2(n10864), .A(n13812), .B(n10863), .ZN(
        n10875) );
  NAND2_X1 U13383 ( .A1(n10866), .A2(n10865), .ZN(n10867) );
  NAND2_X1 U13384 ( .A1(n13778), .A2(n10463), .ZN(n10870) );
  OR2_X1 U13385 ( .A1(n14670), .A2(n13627), .ZN(n10869) );
  AND2_X1 U13386 ( .A1(n10870), .A2(n10869), .ZN(n10888) );
  OAI22_X1 U13387 ( .A1(n14670), .A2(n13629), .B1(n10871), .B2(n13627), .ZN(
        n10872) );
  XNOR2_X1 U13388 ( .A(n10872), .B(n13625), .ZN(n10886) );
  XNOR2_X1 U13389 ( .A(n10887), .B(n10886), .ZN(n10873) );
  NOR2_X1 U13390 ( .A1(n10873), .A2(n13751), .ZN(n10874) );
  AOI211_X1 U13391 ( .C1(n10876), .C2(n14398), .A(n10875), .B(n10874), .ZN(
        n10877) );
  INV_X1 U13392 ( .A(n10877), .ZN(P1_U3230) );
  INV_X1 U13393 ( .A(n10878), .ZN(n10879) );
  OAI222_X1 U13394 ( .A1(P3_U3151), .A2(n10881), .B1(n11881), .B2(n10880), 
        .C1(n11970), .C2(n10879), .ZN(P3_U3274) );
  NAND2_X1 U13395 ( .A1(n10901), .A2(n13587), .ZN(n10883) );
  NAND2_X1 U13396 ( .A1(n13777), .A2(n6460), .ZN(n10882) );
  NAND2_X1 U13397 ( .A1(n10883), .A2(n10882), .ZN(n10884) );
  XNOR2_X1 U13398 ( .A(n10884), .B(n13561), .ZN(n11014) );
  AND2_X1 U13399 ( .A1(n13777), .A2(n10463), .ZN(n10885) );
  AOI21_X1 U13400 ( .B1(n10901), .B2(n13555), .A(n10885), .ZN(n11013) );
  XNOR2_X1 U13401 ( .A(n11014), .B(n11013), .ZN(n10894) );
  INV_X1 U13402 ( .A(n10888), .ZN(n10889) );
  NAND2_X1 U13403 ( .A1(n10890), .A2(n10889), .ZN(n10891) );
  INV_X1 U13404 ( .A(n13717), .ZN(n10892) );
  AOI21_X1 U13405 ( .B1(n10894), .B2(n10893), .A(n10892), .ZN(n10903) );
  INV_X1 U13406 ( .A(n10895), .ZN(n10899) );
  NAND2_X1 U13407 ( .A1(n14397), .A2(n10896), .ZN(n10897) );
  OAI211_X1 U13408 ( .C1(n14401), .C2(n10899), .A(n10898), .B(n10897), .ZN(
        n10900) );
  AOI21_X1 U13409 ( .B1(n10901), .B2(n14398), .A(n10900), .ZN(n10902) );
  OAI21_X1 U13410 ( .B1(n10903), .B2(n13751), .A(n10902), .ZN(P1_U3227) );
  INV_X1 U13411 ( .A(n10904), .ZN(n11158) );
  NAND2_X1 U13412 ( .A1(n14378), .A2(n10905), .ZN(n10907) );
  OAI211_X1 U13413 ( .C1(n14384), .C2(n11158), .A(n10907), .B(n10906), .ZN(
        n10912) );
  INV_X1 U13414 ( .A(n10796), .ZN(n10908) );
  AOI211_X1 U13415 ( .C1(n10910), .C2(n10909), .A(n12759), .B(n10908), .ZN(
        n10911) );
  AOI211_X1 U13416 ( .C1(n12849), .C2(n14381), .A(n10912), .B(n10911), .ZN(
        n10913) );
  INV_X1 U13417 ( .A(n10913), .ZN(P2_U3211) );
  XOR2_X1 U13418 ( .A(n10915), .B(n10914), .Z(n10920) );
  OAI22_X1 U13419 ( .A1(n14988), .A2(n12141), .B1(n12172), .B2(n14987), .ZN(
        n10916) );
  AOI211_X1 U13420 ( .C1(n14994), .C2(n14918), .A(n10917), .B(n10916), .ZN(
        n10919) );
  NAND2_X1 U13421 ( .A1(n12174), .A2(n14995), .ZN(n10918) );
  OAI211_X1 U13422 ( .C1(n10920), .C2(n12153), .A(n10919), .B(n10918), .ZN(
        P3_U3167) );
  NAND2_X1 U13423 ( .A1(n10922), .A2(n10921), .ZN(n10924) );
  XOR2_X1 U13424 ( .A(n10924), .B(n10923), .Z(n10931) );
  NAND2_X1 U13425 ( .A1(n13036), .A2(n13064), .ZN(n10926) );
  INV_X1 U13426 ( .A(n13062), .ZN(n10970) );
  OR2_X1 U13427 ( .A1(n12773), .A2(n10970), .ZN(n10925) );
  NAND2_X1 U13428 ( .A1(n10926), .A2(n10925), .ZN(n11136) );
  AOI22_X1 U13429 ( .A1(n14378), .A2(n11136), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10927) );
  OAI21_X1 U13430 ( .B1(n10928), .B2(n14384), .A(n10927), .ZN(n10929) );
  AOI21_X1 U13431 ( .B1(n14885), .B2(n14381), .A(n10929), .ZN(n10930) );
  OAI21_X1 U13432 ( .B1(n10931), .B2(n12759), .A(n10930), .ZN(P2_U3193) );
  XNOR2_X1 U13433 ( .A(n10933), .B(n10932), .ZN(n14708) );
  INV_X1 U13434 ( .A(n10934), .ZN(n10935) );
  AOI21_X1 U13435 ( .B1(n10937), .B2(n10936), .A(n10935), .ZN(n10938) );
  AOI22_X1 U13436 ( .A1(n14387), .A2(n13774), .B1(n13772), .B2(n13732), .ZN(
        n11336) );
  OAI21_X1 U13437 ( .B1(n10938), .B2(n14608), .A(n11336), .ZN(n14703) );
  INV_X1 U13438 ( .A(n14705), .ZN(n11341) );
  NAND2_X1 U13439 ( .A1(n10939), .A2(n14705), .ZN(n10940) );
  NAND2_X1 U13440 ( .A1(n10940), .A2(n14617), .ZN(n10941) );
  NOR2_X1 U13441 ( .A1(n11001), .A2(n10941), .ZN(n14704) );
  NAND2_X1 U13442 ( .A1(n14704), .A2(n14644), .ZN(n10943) );
  AOI22_X1 U13443 ( .A1(n14638), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11338), 
        .B2(n14637), .ZN(n10942) );
  OAI211_X1 U13444 ( .C1(n11341), .C2(n14640), .A(n10943), .B(n10942), .ZN(
        n10944) );
  AOI21_X1 U13445 ( .B1(n14703), .B2(n14008), .A(n10944), .ZN(n10945) );
  OAI21_X1 U13446 ( .B1(n14016), .B2(n14708), .A(n10945), .ZN(P1_U3284) );
  INV_X1 U13447 ( .A(n11103), .ZN(n10955) );
  OAI211_X1 U13448 ( .C1(n10948), .C2(n10947), .A(n10946), .B(n14914), .ZN(
        n10954) );
  INV_X1 U13449 ( .A(n10949), .ZN(n10951) );
  OAI22_X1 U13450 ( .A1(n15005), .A2(n12141), .B1(n12172), .B2(n11311), .ZN(
        n10950) );
  AOI211_X1 U13451 ( .C1(n10952), .C2(n14918), .A(n10951), .B(n10950), .ZN(
        n10953) );
  OAI211_X1 U13452 ( .C1(n10955), .C2(n12161), .A(n10954), .B(n10953), .ZN(
        P3_U3179) );
  OR2_X1 U13453 ( .A1(n12849), .A2(n13065), .ZN(n10957) );
  NOR2_X1 U13454 ( .A1(n12853), .A2(n13064), .ZN(n10958) );
  XNOR2_X1 U13455 ( .A(n14885), .B(n13063), .ZN(n13002) );
  INV_X1 U13456 ( .A(n13002), .ZN(n11132) );
  NAND2_X1 U13457 ( .A1(n14885), .A2(n13063), .ZN(n10959) );
  XNOR2_X1 U13458 ( .A(n12865), .B(n10970), .ZN(n13004) );
  NAND2_X1 U13459 ( .A1(n11036), .A2(n13004), .ZN(n10961) );
  NAND2_X1 U13460 ( .A1(n12865), .A2(n13062), .ZN(n10960) );
  NAND2_X1 U13461 ( .A1(n10961), .A2(n10960), .ZN(n11177) );
  XNOR2_X1 U13462 ( .A(n14892), .B(n13061), .ZN(n13005) );
  XNOR2_X1 U13463 ( .A(n11177), .B(n11176), .ZN(n14896) );
  OR2_X1 U13464 ( .A1(n12853), .A2(n10964), .ZN(n10966) );
  AND2_X1 U13465 ( .A1(n12853), .A2(n10964), .ZN(n10965) );
  OR2_X1 U13466 ( .A1(n14885), .A2(n10967), .ZN(n10968) );
  NAND2_X1 U13467 ( .A1(n12865), .A2(n10970), .ZN(n10969) );
  XNOR2_X1 U13468 ( .A(n11166), .B(n11176), .ZN(n10971) );
  NAND2_X1 U13469 ( .A1(n10971), .A2(n13198), .ZN(n10974) );
  INV_X1 U13470 ( .A(n13060), .ZN(n11164) );
  OR2_X1 U13471 ( .A1(n12773), .A2(n11164), .ZN(n10973) );
  NAND2_X1 U13472 ( .A1(n13036), .A2(n13062), .ZN(n10972) );
  AND2_X1 U13473 ( .A1(n10973), .A2(n10972), .ZN(n11274) );
  OAI211_X1 U13474 ( .C1(n14896), .C2(n10336), .A(n10974), .B(n11274), .ZN(
        n14898) );
  NAND2_X1 U13475 ( .A1(n14898), .A2(n13248), .ZN(n10981) );
  INV_X1 U13476 ( .A(n11277), .ZN(n10975) );
  OAI22_X1 U13477 ( .A1(n13248), .A2(n10223), .B1(n10975), .B2(n13226), .ZN(
        n10979) );
  NAND2_X1 U13478 ( .A1(n14877), .A2(n11283), .ZN(n11282) );
  NAND2_X1 U13479 ( .A1(n14892), .A2(n11037), .ZN(n10976) );
  NAND2_X1 U13480 ( .A1(n10976), .A2(n13106), .ZN(n10977) );
  OR2_X1 U13481 ( .A1(n11179), .A2(n10977), .ZN(n14894) );
  NOR2_X1 U13482 ( .A1(n14894), .A2(n13184), .ZN(n10978) );
  AOI211_X1 U13483 ( .C1(n13230), .C2(n14892), .A(n10979), .B(n10978), .ZN(
        n10980) );
  OAI211_X1 U13484 ( .C1(n14896), .C2(n13258), .A(n10981), .B(n10980), .ZN(
        P2_U3255) );
  AOI21_X1 U13485 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n10987), .A(n10982), .ZN(
        n10984) );
  XNOR2_X1 U13486 ( .A(n11428), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n10983) );
  AOI211_X1 U13487 ( .C1(n10984), .C2(n10983), .A(n14572), .B(n11419), .ZN(
        n10994) );
  INV_X1 U13488 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10985) );
  MUX2_X1 U13489 ( .A(n10985), .B(P1_REG1_REG_10__SCAN_IN), .S(n11428), .Z(
        n10989) );
  OAI21_X1 U13490 ( .B1(n10987), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10986), .ZN(
        n10988) );
  NOR2_X1 U13491 ( .A1(n10988), .A2(n10989), .ZN(n11427) );
  AOI211_X1 U13492 ( .C1(n10989), .C2(n10988), .A(n14576), .B(n11427), .ZN(
        n10993) );
  NAND2_X1 U13493 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11375)
         );
  NAND2_X1 U13494 ( .A1(n14491), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n10990) );
  OAI211_X1 U13495 ( .C1(n14566), .C2(n10991), .A(n11375), .B(n10990), .ZN(
        n10992) );
  OR3_X1 U13496 ( .A1(n10994), .A2(n10993), .A3(n10992), .ZN(P1_U3253) );
  XNOR2_X1 U13497 ( .A(n10995), .B(n10996), .ZN(n14715) );
  INV_X1 U13498 ( .A(n14715), .ZN(n11007) );
  NAND2_X1 U13499 ( .A1(n10997), .A2(n10996), .ZN(n10998) );
  NAND3_X1 U13500 ( .A1(n10999), .A2(n14630), .A3(n10998), .ZN(n11000) );
  NAND2_X1 U13501 ( .A1(n13773), .A2(n14387), .ZN(n11376) );
  NAND2_X1 U13502 ( .A1(n11000), .A2(n11376), .ZN(n14720) );
  OAI211_X1 U13503 ( .C1(n14718), .C2(n11001), .A(n11219), .B(n14617), .ZN(
        n11002) );
  NAND2_X1 U13504 ( .A1(n13771), .A2(n13732), .ZN(n11377) );
  AND2_X1 U13505 ( .A1(n11002), .A2(n11377), .ZN(n14716) );
  AOI22_X1 U13506 ( .A1(n14648), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11380), 
        .B2(n14637), .ZN(n11004) );
  NAND2_X1 U13507 ( .A1(n11381), .A2(n14409), .ZN(n11003) );
  OAI211_X1 U13508 ( .C1(n14716), .C2(n14011), .A(n11004), .B(n11003), .ZN(
        n11005) );
  AOI21_X1 U13509 ( .B1(n14720), .B2(n14008), .A(n11005), .ZN(n11006) );
  OAI21_X1 U13510 ( .B1(n11007), .B2(n14016), .A(n11006), .ZN(P1_U3283) );
  NAND2_X1 U13511 ( .A1(n13723), .A2(n13587), .ZN(n11009) );
  NAND2_X1 U13512 ( .A1(n13776), .A2(n13555), .ZN(n11008) );
  NAND2_X1 U13513 ( .A1(n11009), .A2(n11008), .ZN(n11010) );
  XNOR2_X1 U13514 ( .A(n11010), .B(n13625), .ZN(n11018) );
  AND2_X1 U13515 ( .A1(n13776), .A2(n10463), .ZN(n11012) );
  AOI21_X1 U13516 ( .B1(n13723), .B2(n13555), .A(n11012), .ZN(n11016) );
  XNOR2_X1 U13517 ( .A(n11018), .B(n11016), .ZN(n13719) );
  NAND2_X1 U13518 ( .A1(n11014), .A2(n11013), .ZN(n13716) );
  AND2_X1 U13519 ( .A1(n13719), .A2(n13716), .ZN(n11015) );
  INV_X1 U13520 ( .A(n11016), .ZN(n11017) );
  NAND2_X1 U13521 ( .A1(n11018), .A2(n11017), .ZN(n11019) );
  NAND2_X1 U13522 ( .A1(n11029), .A2(n13587), .ZN(n11021) );
  NAND2_X1 U13523 ( .A1(n13775), .A2(n13555), .ZN(n11020) );
  NAND2_X1 U13524 ( .A1(n11021), .A2(n11020), .ZN(n11022) );
  XNOR2_X1 U13525 ( .A(n11022), .B(n13625), .ZN(n11260) );
  AND2_X1 U13526 ( .A1(n13775), .A2(n10463), .ZN(n11023) );
  AOI21_X1 U13527 ( .B1(n11029), .B2(n6460), .A(n11023), .ZN(n11258) );
  XNOR2_X1 U13528 ( .A(n11260), .B(n11258), .ZN(n11261) );
  XNOR2_X1 U13529 ( .A(n11262), .B(n11261), .ZN(n11031) );
  INV_X1 U13530 ( .A(n14401), .ZN(n13739) );
  NAND2_X1 U13531 ( .A1(n13739), .A2(n11024), .ZN(n11026) );
  OAI211_X1 U13532 ( .C1(n11027), .C2(n13737), .A(n11026), .B(n11025), .ZN(
        n11028) );
  AOI21_X1 U13533 ( .B1(n11029), .B2(n14398), .A(n11028), .ZN(n11030) );
  OAI21_X1 U13534 ( .B1(n11031), .B2(n13751), .A(n11030), .ZN(P1_U3213) );
  INV_X1 U13535 ( .A(n11032), .ZN(n11035) );
  OAI22_X1 U13536 ( .A1(n11033), .A2(P3_U3151), .B1(SI_22_), .B2(n11881), .ZN(
        n11034) );
  AOI21_X1 U13537 ( .B1(n11035), .B2(n12646), .A(n11034), .ZN(P3_U3273) );
  XNOR2_X1 U13538 ( .A(n11036), .B(n13004), .ZN(n11131) );
  INV_X1 U13539 ( .A(n11131), .ZN(n11044) );
  INV_X1 U13540 ( .A(n11037), .ZN(n11038) );
  AOI211_X1 U13541 ( .C1(n12865), .C2(n11139), .A(n13231), .B(n11038), .ZN(
        n11128) );
  XNOR2_X1 U13542 ( .A(n11039), .B(n13004), .ZN(n11040) );
  NAND2_X1 U13543 ( .A1(n11040), .A2(n13198), .ZN(n11043) );
  INV_X1 U13544 ( .A(n13061), .ZN(n11167) );
  OR2_X1 U13545 ( .A1(n12773), .A2(n11167), .ZN(n11042) );
  NAND2_X1 U13546 ( .A1(n13036), .A2(n13063), .ZN(n11041) );
  AND2_X1 U13547 ( .A1(n11042), .A2(n11041), .ZN(n11191) );
  OAI211_X1 U13548 ( .C1(n11131), .C2(n10336), .A(n11043), .B(n11191), .ZN(
        n11125) );
  AOI211_X1 U13549 ( .C1(n14873), .C2(n11044), .A(n11128), .B(n11125), .ZN(
        n11052) );
  INV_X1 U13550 ( .A(n13370), .ZN(n13379) );
  AOI22_X1 U13551 ( .A1(n13379), .A2(n12865), .B1(n14910), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11045) );
  OAI21_X1 U13552 ( .B1(n11052), .B2(n14910), .A(n11045), .ZN(P2_U3508) );
  NAND2_X1 U13553 ( .A1(n15282), .A2(n14891), .ZN(n13432) );
  INV_X1 U13554 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n11049) );
  OAI22_X1 U13555 ( .A1(n7036), .A2(n13432), .B1(n15282), .B2(n11049), .ZN(
        n11050) );
  INV_X1 U13556 ( .A(n11050), .ZN(n11051) );
  OAI21_X1 U13557 ( .B1(n11052), .B2(n14899), .A(n11051), .ZN(P2_U3457) );
  INV_X1 U13558 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11058) );
  INV_X1 U13559 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11053) );
  MUX2_X1 U13560 ( .A(P3_REG2_REG_8__SCAN_IN), .B(n11053), .S(n11077), .Z(
        n11054) );
  INV_X1 U13561 ( .A(n11054), .ZN(n14932) );
  AOI21_X1 U13562 ( .B1(n11058), .B2(n11057), .A(n11227), .ZN(n11084) );
  MUX2_X1 U13563 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12198), .Z(n11063) );
  INV_X1 U13564 ( .A(n11077), .ZN(n14947) );
  XNOR2_X1 U13565 ( .A(n11063), .B(n14947), .ZN(n14941) );
  NAND2_X1 U13566 ( .A1(n11060), .A2(n11059), .ZN(n11062) );
  NAND2_X1 U13567 ( .A1(n11062), .A2(n11061), .ZN(n14942) );
  NAND2_X1 U13568 ( .A1(n14941), .A2(n14942), .ZN(n11066) );
  INV_X1 U13569 ( .A(n11063), .ZN(n11064) );
  NAND2_X1 U13570 ( .A1(n11064), .A2(n14947), .ZN(n11065) );
  NAND2_X1 U13571 ( .A1(n11066), .A2(n11065), .ZN(n11070) );
  MUX2_X1 U13572 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12198), .Z(n11067) );
  NAND2_X1 U13573 ( .A1(n11067), .A2(n11073), .ZN(n11069) );
  INV_X1 U13574 ( .A(n11067), .ZN(n11068) );
  NAND2_X1 U13575 ( .A1(n11068), .A2(n11233), .ZN(n11241) );
  AND2_X1 U13576 ( .A1(n11241), .A2(n11069), .ZN(n11071) );
  OAI22_X1 U13577 ( .A1(n11242), .A2(n6869), .B1(n11071), .B2(n11070), .ZN(
        n11082) );
  AND2_X1 U13578 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11487) );
  AOI21_X1 U13579 ( .B1(n14921), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11487), .ZN(
        n11072) );
  OAI21_X1 U13580 ( .B1(n11247), .B2(n11073), .A(n11072), .ZN(n11081) );
  INV_X1 U13581 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11465) );
  INV_X1 U13582 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11074) );
  MUX2_X1 U13583 ( .A(n11074), .B(P3_REG1_REG_8__SCAN_IN), .S(n11077), .Z(
        n14935) );
  NOR2_X1 U13584 ( .A1(n14935), .A2(n14936), .ZN(n14934) );
  AOI21_X1 U13585 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n11077), .A(n14934), .ZN(
        n11232) );
  AOI21_X1 U13586 ( .B1(n11465), .B2(n11078), .A(n11234), .ZN(n11079) );
  NOR2_X1 U13587 ( .A1(n11079), .A2(n14937), .ZN(n11080) );
  AOI211_X1 U13588 ( .C1(n14922), .C2(n11082), .A(n11081), .B(n11080), .ZN(
        n11083) );
  OAI21_X1 U13589 ( .B1(n11084), .B2(n14940), .A(n11083), .ZN(P3_U3191) );
  INV_X1 U13590 ( .A(n11085), .ZN(n11088) );
  OAI222_X1 U13591 ( .A1(n13464), .A2(n11086), .B1(n13459), .B2(n11088), .C1(
        P2_U3088), .C2(n13026), .ZN(P2_U3308) );
  OAI222_X1 U13592 ( .A1(n13858), .A2(P1_U3086), .B1(n14166), .B2(n11088), 
        .C1(n11087), .C2(n14163), .ZN(P1_U3336) );
  OR2_X1 U13593 ( .A1(n11090), .A2(n11089), .ZN(n11091) );
  NAND2_X1 U13594 ( .A1(n11092), .A2(n11091), .ZN(n15072) );
  INV_X1 U13595 ( .A(n15072), .ZN(n11106) );
  OAI211_X1 U13596 ( .C1(n11095), .C2(n11094), .A(n11093), .B(n15039), .ZN(
        n11100) );
  NAND2_X1 U13597 ( .A1(n12188), .A2(n15034), .ZN(n11096) );
  OAI21_X1 U13598 ( .B1(n11311), .B2(n15017), .A(n11096), .ZN(n11097) );
  AOI21_X1 U13599 ( .B1(n15072), .B2(n11098), .A(n11097), .ZN(n11099) );
  NAND2_X1 U13600 ( .A1(n11100), .A2(n11099), .ZN(n15070) );
  MUX2_X1 U13601 ( .A(n15070), .B(P3_REG2_REG_6__SCAN_IN), .S(n14334), .Z(
        n11101) );
  INV_X1 U13602 ( .A(n11101), .ZN(n11105) );
  NOR2_X1 U13603 ( .A1(n11102), .A2(n15030), .ZN(n15071) );
  AOI22_X1 U13604 ( .A1(n15071), .A2(n15000), .B1(n15046), .B2(n11103), .ZN(
        n11104) );
  OAI211_X1 U13605 ( .C1(n11106), .C2(n11204), .A(n11105), .B(n11104), .ZN(
        P3_U3227) );
  AOI21_X1 U13606 ( .B1(n11111), .B2(P2_REG1_REG_13__SCAN_IN), .A(n11107), 
        .ZN(n14800) );
  XNOR2_X1 U13607 ( .A(n14803), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14799) );
  NOR2_X1 U13608 ( .A1(n14800), .A2(n14799), .ZN(n14798) );
  AOI21_X1 U13609 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n14803), .A(n14798), 
        .ZN(n11437) );
  INV_X1 U13610 ( .A(n11108), .ZN(n11110) );
  INV_X1 U13611 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11109) );
  OAI211_X1 U13612 ( .C1(n11110), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14784), 
        .B(n6622), .ZN(n11124) );
  NOR2_X1 U13613 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11836), .ZN(n11122) );
  NAND2_X1 U13614 ( .A1(n11111), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11115) );
  OR2_X1 U13615 ( .A1(n11113), .A2(n11112), .ZN(n11114) );
  NAND2_X1 U13616 ( .A1(n11115), .A2(n11114), .ZN(n11116) );
  NAND2_X1 U13617 ( .A1(n14803), .A2(n11116), .ZN(n11117) );
  XOR2_X1 U13618 ( .A(n14803), .B(n11116), .Z(n14807) );
  NAND2_X1 U13619 ( .A1(n14807), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n14806) );
  NAND2_X1 U13620 ( .A1(n11117), .A2(n14806), .ZN(n11440) );
  INV_X1 U13621 ( .A(n11440), .ZN(n11118) );
  XNOR2_X1 U13622 ( .A(n11441), .B(n11118), .ZN(n11119) );
  NAND2_X1 U13623 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n11119), .ZN(n11442) );
  OAI211_X1 U13624 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n11119), .A(n14805), 
        .B(n11442), .ZN(n11120) );
  INV_X1 U13625 ( .A(n11120), .ZN(n11121) );
  AOI211_X1 U13626 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n14819), .A(n11122), 
        .B(n11121), .ZN(n11123) );
  OAI211_X1 U13627 ( .C1(n14827), .C2(n11436), .A(n11124), .B(n11123), .ZN(
        P2_U3229) );
  NAND2_X1 U13628 ( .A1(n11125), .A2(n13248), .ZN(n11130) );
  AOI22_X1 U13629 ( .A1(n13298), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11194), 
        .B2(n13289), .ZN(n11126) );
  OAI21_X1 U13630 ( .B1(n7036), .B2(n13293), .A(n11126), .ZN(n11127) );
  AOI21_X1 U13631 ( .B1(n11128), .B2(n13288), .A(n11127), .ZN(n11129) );
  OAI211_X1 U13632 ( .C1(n11131), .C2(n13258), .A(n11130), .B(n11129), .ZN(
        P2_U3256) );
  XNOR2_X1 U13633 ( .A(n11133), .B(n11132), .ZN(n14887) );
  OAI211_X1 U13634 ( .C1(n11135), .C2(n13002), .A(n11134), .B(n13198), .ZN(
        n11138) );
  INV_X1 U13635 ( .A(n11136), .ZN(n11137) );
  NAND2_X1 U13636 ( .A1(n11138), .A2(n11137), .ZN(n14883) );
  INV_X1 U13637 ( .A(n14885), .ZN(n11143) );
  AOI211_X1 U13638 ( .C1(n14885), .C2(n11282), .A(n13089), .B(n7037), .ZN(
        n14884) );
  NAND2_X1 U13639 ( .A1(n14884), .A2(n13288), .ZN(n11142) );
  AOI22_X1 U13640 ( .A1(n13298), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n11140), 
        .B2(n13289), .ZN(n11141) );
  OAI211_X1 U13641 ( .C1(n11143), .C2(n13293), .A(n11142), .B(n11141), .ZN(
        n11144) );
  AOI21_X1 U13642 ( .B1(n13248), .B2(n14883), .A(n11144), .ZN(n11145) );
  OAI21_X1 U13643 ( .B1(n14887), .B2(n13238), .A(n11145), .ZN(P2_U3257) );
  INV_X1 U13644 ( .A(n14974), .ZN(n11154) );
  OAI211_X1 U13645 ( .C1(n11148), .C2(n11147), .A(n11146), .B(n14914), .ZN(
        n11153) );
  OAI22_X1 U13646 ( .A1(n11458), .A2(n12172), .B1(n12141), .B2(n14987), .ZN(
        n11149) );
  AOI211_X1 U13647 ( .C1(n11151), .C2(n14918), .A(n11150), .B(n11149), .ZN(
        n11152) );
  OAI211_X1 U13648 ( .C1(n11154), .C2(n12161), .A(n11153), .B(n11152), .ZN(
        P3_U3153) );
  INV_X1 U13649 ( .A(n11155), .ZN(n11163) );
  MUX2_X1 U13650 ( .A(n11156), .B(P2_REG2_REG_6__SCAN_IN), .S(n13298), .Z(
        n11157) );
  INV_X1 U13651 ( .A(n11157), .ZN(n11162) );
  OAI22_X1 U13652 ( .A1(n13293), .A2(n6657), .B1(n13226), .B2(n11158), .ZN(
        n11159) );
  AOI21_X1 U13653 ( .B1(n11160), .B2(n13288), .A(n11159), .ZN(n11161) );
  OAI211_X1 U13654 ( .C1(n11163), .C2(n13258), .A(n11162), .B(n11161), .ZN(
        P2_U3259) );
  NAND2_X1 U13655 ( .A1(n12875), .A2(n11164), .ZN(n11292) );
  OR2_X1 U13656 ( .A1(n12875), .A2(n11164), .ZN(n11165) );
  INV_X1 U13657 ( .A(n13007), .ZN(n11172) );
  NAND2_X1 U13658 ( .A1(n11166), .A2(n13005), .ZN(n11169) );
  OR2_X1 U13659 ( .A1(n14892), .A2(n11167), .ZN(n11168) );
  NAND2_X1 U13660 ( .A1(n11169), .A2(n11168), .ZN(n11171) );
  INV_X1 U13661 ( .A(n11293), .ZN(n11170) );
  AOI21_X1 U13662 ( .B1(n11172), .B2(n11171), .A(n11170), .ZN(n11175) );
  INV_X1 U13663 ( .A(n13059), .ZN(n11387) );
  OR2_X1 U13664 ( .A1(n12773), .A2(n11387), .ZN(n11174) );
  NAND2_X1 U13665 ( .A1(n13036), .A2(n13061), .ZN(n11173) );
  AND2_X1 U13666 ( .A1(n11174), .A2(n11173), .ZN(n11545) );
  OAI21_X1 U13667 ( .B1(n11175), .B2(n13281), .A(n11545), .ZN(n11358) );
  INV_X1 U13668 ( .A(n11358), .ZN(n11186) );
  NAND2_X1 U13669 ( .A1(n14892), .A2(n13061), .ZN(n11178) );
  XNOR2_X1 U13670 ( .A(n11298), .B(n13007), .ZN(n11360) );
  INV_X1 U13671 ( .A(n12875), .ZN(n11363) );
  INV_X1 U13672 ( .A(n11179), .ZN(n11181) );
  INV_X1 U13673 ( .A(n11300), .ZN(n11180) );
  AOI211_X1 U13674 ( .C1(n12875), .C2(n11181), .A(n13089), .B(n11180), .ZN(
        n11359) );
  NAND2_X1 U13675 ( .A1(n11359), .A2(n13288), .ZN(n11183) );
  AOI22_X1 U13676 ( .A1(n13298), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n11542), 
        .B2(n13289), .ZN(n11182) );
  OAI211_X1 U13677 ( .C1(n11363), .C2(n13293), .A(n11183), .B(n11182), .ZN(
        n11184) );
  AOI21_X1 U13678 ( .B1(n13295), .B2(n11360), .A(n11184), .ZN(n11185) );
  OAI21_X1 U13679 ( .B1(n11186), .B2(n13298), .A(n11185), .ZN(P2_U3254) );
  INV_X1 U13680 ( .A(n11187), .ZN(n11188) );
  AOI21_X1 U13681 ( .B1(n11190), .B2(n11189), .A(n11188), .ZN(n11196) );
  NAND2_X1 U13682 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n14794) );
  OAI21_X1 U13683 ( .B1(n12751), .B2(n11191), .A(n14794), .ZN(n11193) );
  NOR2_X1 U13684 ( .A1(n7036), .A2(n12776), .ZN(n11192) );
  AOI211_X1 U13685 ( .C1(n12770), .C2(n11194), .A(n11193), .B(n11192), .ZN(
        n11195) );
  OAI21_X1 U13686 ( .B1(n11196), .B2(n12759), .A(n11195), .ZN(P2_U3203) );
  XOR2_X1 U13687 ( .A(n11198), .B(n11197), .Z(n11203) );
  XNOR2_X1 U13688 ( .A(n11199), .B(n11198), .ZN(n11200) );
  NAND2_X1 U13689 ( .A1(n11200), .A2(n15039), .ZN(n11202) );
  AOI22_X1 U13690 ( .A1(n12187), .A2(n15034), .B1(n15035), .B2(n12186), .ZN(
        n11201) );
  OAI211_X1 U13691 ( .C1(n11203), .C2(n15043), .A(n11202), .B(n11201), .ZN(
        n15076) );
  INV_X1 U13692 ( .A(n15076), .ZN(n11209) );
  INV_X1 U13693 ( .A(n11203), .ZN(n15078) );
  INV_X1 U13694 ( .A(n11204), .ZN(n15047) );
  INV_X1 U13695 ( .A(n11315), .ZN(n11205) );
  NOR2_X1 U13696 ( .A1(n11205), .A2(n15030), .ZN(n15077) );
  AOI22_X1 U13697 ( .A1(n15077), .A2(n15000), .B1(n15046), .B2(n11307), .ZN(
        n11206) );
  OAI21_X1 U13698 ( .B1(n11053), .B2(n15050), .A(n11206), .ZN(n11207) );
  AOI21_X1 U13699 ( .B1(n15078), .B2(n15047), .A(n11207), .ZN(n11208) );
  OAI21_X1 U13700 ( .B1(n11209), .B2(n14334), .A(n11208), .ZN(P3_U3225) );
  XNOR2_X1 U13701 ( .A(n11212), .B(n11211), .ZN(n14452) );
  INV_X1 U13702 ( .A(n14452), .ZN(n11225) );
  OAI211_X1 U13703 ( .C1(n11215), .C2(n11214), .A(n11213), .B(n14630), .ZN(
        n11218) );
  NAND2_X1 U13704 ( .A1(n13772), .A2(n14387), .ZN(n11217) );
  NAND2_X1 U13705 ( .A1(n13770), .A2(n13732), .ZN(n11216) );
  AND2_X1 U13706 ( .A1(n11217), .A2(n11216), .ZN(n11644) );
  NAND2_X1 U13707 ( .A1(n11218), .A2(n11644), .ZN(n14457) );
  AOI21_X1 U13708 ( .B1(n11219), .B2(n14453), .A(n14675), .ZN(n11220) );
  NAND2_X1 U13709 ( .A1(n11220), .A2(n11351), .ZN(n14455) );
  AOI22_X1 U13710 ( .A1(n14638), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11642), 
        .B2(n14637), .ZN(n11222) );
  NAND2_X1 U13711 ( .A1(n14453), .A2(n14409), .ZN(n11221) );
  OAI211_X1 U13712 ( .C1(n14455), .C2(n14011), .A(n11222), .B(n11221), .ZN(
        n11223) );
  AOI21_X1 U13713 ( .B1(n14457), .B2(n14008), .A(n11223), .ZN(n11224) );
  OAI21_X1 U13714 ( .B1(n14016), .B2(n11225), .A(n11224), .ZN(P1_U3282) );
  NOR2_X1 U13715 ( .A1(n11233), .A2(n11226), .ZN(n11228) );
  INV_X1 U13716 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11516) );
  MUX2_X1 U13717 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n11516), .S(n11529), .Z(
        n11230) );
  INV_X1 U13718 ( .A(n11518), .ZN(n11229) );
  AOI21_X1 U13719 ( .B1(n11231), .B2(n11230), .A(n11229), .ZN(n11252) );
  NOR2_X1 U13720 ( .A1(n11233), .A2(n11232), .ZN(n11235) );
  INV_X1 U13721 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11528) );
  MUX2_X1 U13722 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n11528), .S(n11529), .Z(
        n11236) );
  OAI21_X1 U13723 ( .B1(n7072), .B2(n7071), .A(n11531), .ZN(n11250) );
  MUX2_X1 U13724 ( .A(n11516), .B(n11528), .S(n12198), .Z(n11237) );
  INV_X1 U13725 ( .A(n11237), .ZN(n11238) );
  NAND2_X1 U13726 ( .A1(n11238), .A2(n11246), .ZN(n11239) );
  NAND2_X1 U13727 ( .A1(n6604), .A2(n11239), .ZN(n11240) );
  NAND3_X1 U13728 ( .A1(n11242), .A2(n11241), .A3(n11240), .ZN(n11243) );
  AOI21_X1 U13729 ( .B1(n6615), .B2(n11243), .A(n14943), .ZN(n11249) );
  NAND2_X1 U13730 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(P3_U3151), .ZN(n11666)
         );
  INV_X1 U13731 ( .A(n11666), .ZN(n11244) );
  AOI21_X1 U13732 ( .B1(n14921), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11244), 
        .ZN(n11245) );
  OAI21_X1 U13733 ( .B1(n11247), .B2(n11246), .A(n11245), .ZN(n11248) );
  AOI211_X1 U13734 ( .C1(n11250), .C2(n14924), .A(n11249), .B(n11248), .ZN(
        n11251) );
  OAI21_X1 U13735 ( .B1(n11252), .B2(n14940), .A(n11251), .ZN(P3_U3192) );
  NAND2_X1 U13736 ( .A1(n11257), .A2(n13587), .ZN(n11254) );
  NAND2_X1 U13737 ( .A1(n13774), .A2(n13555), .ZN(n11253) );
  NAND2_X1 U13738 ( .A1(n11254), .A2(n11253), .ZN(n11255) );
  XNOR2_X1 U13739 ( .A(n11255), .B(n13625), .ZN(n11323) );
  AND2_X1 U13740 ( .A1(n13774), .A2(n10463), .ZN(n11256) );
  AOI21_X1 U13741 ( .B1(n11257), .B2(n6460), .A(n11256), .ZN(n11324) );
  XNOR2_X1 U13742 ( .A(n11323), .B(n11324), .ZN(n11264) );
  INV_X1 U13743 ( .A(n11258), .ZN(n11259) );
  OAI21_X1 U13744 ( .B1(n11264), .B2(n11263), .A(n11332), .ZN(n11265) );
  NAND2_X1 U13745 ( .A1(n11265), .A2(n14395), .ZN(n11271) );
  NOR2_X1 U13746 ( .A1(n13737), .A2(n11266), .ZN(n11267) );
  AOI211_X1 U13747 ( .C1(n13739), .C2(n11269), .A(n11268), .B(n11267), .ZN(
        n11270) );
  OAI211_X1 U13748 ( .C1(n14699), .C2(n13742), .A(n11271), .B(n11270), .ZN(
        P1_U3221) );
  XNOR2_X1 U13749 ( .A(n11273), .B(n11272), .ZN(n11280) );
  NOR2_X1 U13750 ( .A1(n12751), .A2(n11274), .ZN(n11275) );
  AOI211_X1 U13751 ( .C1(n12770), .C2(n11277), .A(n11276), .B(n11275), .ZN(
        n11279) );
  NAND2_X1 U13752 ( .A1(n14892), .A2(n14381), .ZN(n11278) );
  OAI211_X1 U13753 ( .C1(n11280), .C2(n12759), .A(n11279), .B(n11278), .ZN(
        P2_U3189) );
  XNOR2_X1 U13754 ( .A(n12853), .B(n13064), .ZN(n13000) );
  XOR2_X1 U13755 ( .A(n13000), .B(n11281), .Z(n14881) );
  OAI211_X1 U13756 ( .C1(n14877), .C2(n11283), .A(n13106), .B(n11282), .ZN(
        n14875) );
  AOI22_X1 U13757 ( .A1(n13230), .A2(n12853), .B1(n11284), .B2(n13289), .ZN(
        n11285) );
  OAI21_X1 U13758 ( .B1(n13184), .B2(n14875), .A(n11285), .ZN(n11290) );
  XOR2_X1 U13759 ( .A(n11286), .B(n13000), .Z(n11288) );
  OAI21_X1 U13760 ( .B1(n11288), .B2(n13281), .A(n11287), .ZN(n14878) );
  MUX2_X1 U13761 ( .A(n14878), .B(P2_REG2_REG_7__SCAN_IN), .S(n13298), .Z(
        n11289) );
  AOI211_X1 U13762 ( .C1(n13295), .C2(n14881), .A(n11290), .B(n11289), .ZN(
        n11291) );
  INV_X1 U13763 ( .A(n11291), .ZN(P2_U3258) );
  OR2_X1 U13764 ( .A1(n12883), .A2(n13059), .ZN(n11402) );
  NAND2_X1 U13765 ( .A1(n12883), .A2(n13059), .ZN(n11400) );
  NAND2_X1 U13766 ( .A1(n11402), .A2(n11400), .ZN(n13008) );
  XOR2_X1 U13767 ( .A(n11386), .B(n13008), .Z(n11296) );
  INV_X1 U13768 ( .A(n13058), .ZN(n12896) );
  OR2_X1 U13769 ( .A1(n12773), .A2(n12896), .ZN(n11295) );
  NAND2_X1 U13770 ( .A1(n13036), .A2(n13060), .ZN(n11294) );
  AND2_X1 U13771 ( .A1(n11295), .A2(n11294), .ZN(n11583) );
  OAI21_X1 U13772 ( .B1(n11296), .B2(n13281), .A(n11583), .ZN(n11493) );
  INV_X1 U13773 ( .A(n11493), .ZN(n11306) );
  AND2_X1 U13774 ( .A1(n12875), .A2(n13060), .ZN(n11297) );
  XOR2_X1 U13775 ( .A(n11401), .B(n13008), .Z(n11495) );
  INV_X1 U13776 ( .A(n12883), .ZN(n11303) );
  OR2_X1 U13777 ( .A1(n11300), .A2(n12883), .ZN(n11398) );
  INV_X1 U13778 ( .A(n11398), .ZN(n11299) );
  AOI211_X1 U13779 ( .C1(n12883), .C2(n11300), .A(n13231), .B(n11299), .ZN(
        n11494) );
  NAND2_X1 U13780 ( .A1(n11494), .A2(n13288), .ZN(n11302) );
  AOI22_X1 U13781 ( .A1(n13298), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11580), 
        .B2(n13289), .ZN(n11301) );
  OAI211_X1 U13782 ( .C1(n11303), .C2(n13293), .A(n11302), .B(n11301), .ZN(
        n11304) );
  AOI21_X1 U13783 ( .B1(n13295), .B2(n11495), .A(n11304), .ZN(n11305) );
  OAI21_X1 U13784 ( .B1(n11306), .B2(n13298), .A(n11305), .ZN(P2_U3253) );
  INV_X1 U13785 ( .A(n11307), .ZN(n11318) );
  OAI211_X1 U13786 ( .C1(n11310), .C2(n11309), .A(n11308), .B(n14914), .ZN(
        n11317) );
  NAND2_X1 U13787 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n14949) );
  INV_X1 U13788 ( .A(n14949), .ZN(n11314) );
  OAI22_X1 U13789 ( .A1(n11312), .A2(n12172), .B1(n12141), .B2(n11311), .ZN(
        n11313) );
  AOI211_X1 U13790 ( .C1(n11315), .C2(n14918), .A(n11314), .B(n11313), .ZN(
        n11316) );
  OAI211_X1 U13791 ( .C1(n11318), .C2(n12161), .A(n11317), .B(n11316), .ZN(
        P3_U3161) );
  NAND2_X1 U13792 ( .A1(n11319), .A2(n12646), .ZN(n11321) );
  OAI211_X1 U13793 ( .C1(n11322), .C2(n11881), .A(n11321), .B(n11320), .ZN(
        P3_U3272) );
  INV_X1 U13794 ( .A(n11323), .ZN(n11325) );
  NAND2_X1 U13795 ( .A1(n11325), .A2(n11324), .ZN(n11330) );
  AND2_X1 U13796 ( .A1(n11332), .A2(n11330), .ZN(n11334) );
  NAND2_X1 U13797 ( .A1(n14705), .A2(n13587), .ZN(n11327) );
  NAND2_X1 U13798 ( .A1(n13773), .A2(n13555), .ZN(n11326) );
  NAND2_X1 U13799 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  XNOR2_X1 U13800 ( .A(n11328), .B(n13625), .ZN(n11369) );
  AND2_X1 U13801 ( .A1(n13773), .A2(n10463), .ZN(n11329) );
  AOI21_X1 U13802 ( .B1(n14705), .B2(n6460), .A(n11329), .ZN(n11367) );
  XNOR2_X1 U13803 ( .A(n11369), .B(n11367), .ZN(n11333) );
  AND2_X1 U13804 ( .A1(n11333), .A2(n11330), .ZN(n11331) );
  OAI211_X1 U13805 ( .C1(n11334), .C2(n11333), .A(n14395), .B(n11370), .ZN(
        n11340) );
  OAI21_X1 U13806 ( .B1(n13737), .B2(n11336), .A(n11335), .ZN(n11337) );
  AOI21_X1 U13807 ( .B1(n11338), .B2(n13739), .A(n11337), .ZN(n11339) );
  OAI211_X1 U13808 ( .C1(n11341), .C2(n13742), .A(n11340), .B(n11339), .ZN(
        P1_U3231) );
  OAI211_X1 U13809 ( .C1(n11344), .C2(n11343), .A(n11342), .B(n14630), .ZN(
        n11347) );
  NAND2_X1 U13810 ( .A1(n13771), .A2(n14387), .ZN(n11346) );
  NAND2_X1 U13811 ( .A1(n14388), .A2(n13732), .ZN(n11345) );
  AND2_X1 U13812 ( .A1(n11346), .A2(n11345), .ZN(n11685) );
  NAND2_X1 U13813 ( .A1(n11347), .A2(n11685), .ZN(n14309) );
  INV_X1 U13814 ( .A(n14309), .ZN(n11357) );
  XNOR2_X1 U13815 ( .A(n11350), .B(n11349), .ZN(n14305) );
  AND2_X1 U13816 ( .A1(n11678), .A2(n11351), .ZN(n11352) );
  OR2_X1 U13817 ( .A1(n11475), .A2(n11352), .ZN(n14306) );
  AOI22_X1 U13818 ( .A1(n14638), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11687), 
        .B2(n14637), .ZN(n11354) );
  NAND2_X1 U13819 ( .A1(n11678), .A2(n14409), .ZN(n11353) );
  OAI211_X1 U13820 ( .C1(n14306), .C2(n11935), .A(n11354), .B(n11353), .ZN(
        n11355) );
  AOI21_X1 U13821 ( .B1(n14305), .B2(n14419), .A(n11355), .ZN(n11356) );
  OAI21_X1 U13822 ( .B1(n11357), .B2(n14638), .A(n11356), .ZN(P1_U3281) );
  AOI211_X1 U13823 ( .C1(n11360), .C2(n14880), .A(n11359), .B(n11358), .ZN(
        n11366) );
  AOI22_X1 U13824 ( .A1(n12875), .A2(n13379), .B1(n14910), .B2(
        P2_REG1_REG_11__SCAN_IN), .ZN(n11361) );
  OAI21_X1 U13825 ( .B1(n11366), .B2(n14910), .A(n11361), .ZN(P2_U3510) );
  INV_X1 U13826 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11362) );
  OAI22_X1 U13827 ( .A1(n11363), .A2(n13432), .B1(n15282), .B2(n11362), .ZN(
        n11364) );
  INV_X1 U13828 ( .A(n11364), .ZN(n11365) );
  OAI21_X1 U13829 ( .B1(n11366), .B2(n14899), .A(n11365), .ZN(P2_U3463) );
  INV_X1 U13830 ( .A(n11367), .ZN(n11368) );
  NAND2_X1 U13831 ( .A1(n11381), .A2(n13587), .ZN(n11372) );
  NAND2_X1 U13832 ( .A1(n13772), .A2(n13555), .ZN(n11371) );
  NAND2_X1 U13833 ( .A1(n11372), .A2(n11371), .ZN(n11373) );
  XNOR2_X1 U13834 ( .A(n11373), .B(n13625), .ZN(n11635) );
  AND2_X1 U13835 ( .A1(n13772), .A2(n10463), .ZN(n11374) );
  AOI21_X1 U13836 ( .B1(n11381), .B2(n6460), .A(n11374), .ZN(n11633) );
  XNOR2_X1 U13837 ( .A(n11635), .B(n11633), .ZN(n11631) );
  XNOR2_X1 U13838 ( .A(n11632), .B(n11631), .ZN(n11384) );
  INV_X1 U13839 ( .A(n11375), .ZN(n11379) );
  AOI21_X1 U13840 ( .B1(n11377), .B2(n11376), .A(n13737), .ZN(n11378) );
  AOI211_X1 U13841 ( .C1(n13739), .C2(n11380), .A(n11379), .B(n11378), .ZN(
        n11383) );
  NAND2_X1 U13842 ( .A1(n11381), .A2(n14398), .ZN(n11382) );
  OAI211_X1 U13843 ( .C1(n11384), .C2(n13751), .A(n11383), .B(n11382), .ZN(
        P1_U3217) );
  OR2_X1 U13844 ( .A1(n12883), .A2(n11387), .ZN(n11385) );
  NAND2_X1 U13845 ( .A1(n11386), .A2(n11385), .ZN(n11389) );
  NAND2_X1 U13846 ( .A1(n12883), .A2(n11387), .ZN(n11388) );
  OR2_X1 U13847 ( .A1(n13386), .A2(n12896), .ZN(n11559) );
  NAND2_X1 U13848 ( .A1(n13386), .A2(n12896), .ZN(n11390) );
  NAND2_X1 U13849 ( .A1(n11559), .A2(n11390), .ZN(n13010) );
  AOI21_X1 U13850 ( .B1(n11391), .B2(n13010), .A(n13281), .ZN(n11397) );
  NAND2_X1 U13851 ( .A1(n13036), .A2(n13059), .ZN(n11395) );
  INV_X1 U13852 ( .A(n13057), .ZN(n12893) );
  OR2_X1 U13853 ( .A1(n12773), .A2(n12893), .ZN(n11394) );
  AND2_X1 U13854 ( .A1(n11395), .A2(n11394), .ZN(n11694) );
  INV_X1 U13855 ( .A(n11694), .ZN(n11396) );
  AOI21_X1 U13856 ( .B1(n11397), .B2(n11560), .A(n11396), .ZN(n13388) );
  AOI211_X1 U13857 ( .C1(n13386), .C2(n11398), .A(n13089), .B(n11564), .ZN(
        n13385) );
  INV_X1 U13858 ( .A(n13386), .ZN(n12895) );
  AOI22_X1 U13859 ( .A1(n13298), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11696), 
        .B2(n13289), .ZN(n11399) );
  OAI21_X1 U13860 ( .B1(n12895), .B2(n13293), .A(n11399), .ZN(n11404) );
  XOR2_X1 U13861 ( .A(n13010), .B(n11570), .Z(n13389) );
  NOR2_X1 U13862 ( .A1(n13389), .A2(n13238), .ZN(n11403) );
  AOI211_X1 U13863 ( .C1(n13385), .C2(n13288), .A(n11404), .B(n11403), .ZN(
        n11405) );
  OAI21_X1 U13864 ( .B1(n13298), .B2(n13388), .A(n11405), .ZN(P2_U3252) );
  OAI211_X1 U13865 ( .C1(n11407), .C2(n11410), .A(n11406), .B(n15039), .ZN(
        n11409) );
  AOI22_X1 U13866 ( .A1(n12184), .A2(n15035), .B1(n15034), .B2(n12186), .ZN(
        n11408) );
  NAND2_X1 U13867 ( .A1(n11409), .A2(n11408), .ZN(n11549) );
  INV_X1 U13868 ( .A(n11549), .ZN(n11415) );
  XNOR2_X1 U13869 ( .A(n11411), .B(n11410), .ZN(n11550) );
  NAND2_X1 U13870 ( .A1(n15043), .A2(n15026), .ZN(n14953) );
  AOI22_X1 U13871 ( .A1(n14334), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n15046), 
        .B2(n11668), .ZN(n11412) );
  OAI21_X1 U13872 ( .B1(n14958), .B2(n11671), .A(n11412), .ZN(n11413) );
  AOI21_X1 U13873 ( .B1(n11550), .B2(n12520), .A(n11413), .ZN(n11414) );
  OAI21_X1 U13874 ( .B1(n11415), .B2(n14334), .A(n11414), .ZN(P3_U3223) );
  INV_X1 U13875 ( .A(n11416), .ZN(n11452) );
  OAI222_X1 U13876 ( .A1(n13459), .A2(n11452), .B1(n11417), .B2(P2_U3088), 
        .C1(n15251), .C2(n13464), .ZN(P2_U3307) );
  NOR2_X1 U13877 ( .A1(n11862), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11418) );
  AOI21_X1 U13878 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n11862), .A(n11418), 
        .ZN(n11422) );
  MUX2_X1 U13879 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n8405), .S(n11430), .Z(
        n11420) );
  INV_X1 U13880 ( .A(n11420), .ZN(n14500) );
  OAI21_X1 U13881 ( .B1(n11422), .B2(n11421), .A(n11857), .ZN(n11425) );
  NAND2_X1 U13882 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11684)
         );
  NAND2_X1 U13883 ( .A1(n14491), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n11423) );
  OAI211_X1 U13884 ( .C1(n14566), .C2(n11426), .A(n11684), .B(n11423), .ZN(
        n11424) );
  AOI21_X1 U13885 ( .B1(n11425), .B2(n14554), .A(n11424), .ZN(n11435) );
  INV_X1 U13886 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14311) );
  AOI22_X1 U13887 ( .A1(n11862), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n14311), 
        .B2(n11426), .ZN(n11432) );
  INV_X1 U13888 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11429) );
  MUX2_X1 U13889 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n11429), .S(n11430), .Z(
        n14496) );
  NAND2_X1 U13890 ( .A1(n14497), .A2(n14496), .ZN(n14495) );
  OAI21_X1 U13891 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n11430), .A(n14495), 
        .ZN(n11431) );
  NAND2_X1 U13892 ( .A1(n11432), .A2(n11431), .ZN(n11864) );
  OAI21_X1 U13893 ( .B1(n11432), .B2(n11431), .A(n11864), .ZN(n11433) );
  NAND2_X1 U13894 ( .A1(n11433), .A2(n14558), .ZN(n11434) );
  NAND2_X1 U13895 ( .A1(n11435), .A2(n11434), .ZN(P1_U3255) );
  XNOR2_X1 U13896 ( .A(n11739), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n11438) );
  AOI211_X1 U13897 ( .C1(n11439), .C2(n11438), .A(n14813), .B(n11738), .ZN(
        n11451) );
  NAND2_X1 U13898 ( .A1(n11441), .A2(n11440), .ZN(n11443) );
  NAND2_X1 U13899 ( .A1(n11443), .A2(n11442), .ZN(n11446) );
  MUX2_X1 U13900 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n11444), .S(n11739), .Z(
        n11445) );
  NAND2_X1 U13901 ( .A1(n11446), .A2(n11445), .ZN(n11736) );
  OAI211_X1 U13902 ( .C1(n11446), .C2(n11445), .A(n11736), .B(n14805), .ZN(
        n11447) );
  INV_X1 U13903 ( .A(n11447), .ZN(n11450) );
  NAND2_X1 U13904 ( .A1(n14819), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n11448) );
  NAND2_X1 U13905 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n12694)
         );
  OAI211_X1 U13906 ( .C1(n14827), .C2(n11737), .A(n11448), .B(n12694), .ZN(
        n11449) );
  OR3_X1 U13907 ( .A1(n11451), .A2(n11450), .A3(n11449), .ZN(P2_U3230) );
  OAI222_X1 U13908 ( .A1(n11454), .A2(P1_U3086), .B1(n14163), .B2(n11453), 
        .C1(n11452), .C2(n14166), .ZN(P1_U3335) );
  INV_X1 U13909 ( .A(n14362), .ZN(n11462) );
  XOR2_X1 U13910 ( .A(n11455), .B(n11456), .Z(n14955) );
  AOI21_X1 U13911 ( .B1(n11457), .B2(n11456), .A(n12512), .ZN(n11461) );
  OAI22_X1 U13912 ( .A1(n11458), .A2(n15019), .B1(n12140), .B2(n15017), .ZN(
        n11459) );
  AOI21_X1 U13913 ( .B1(n11461), .B2(n11460), .A(n11459), .ZN(n14954) );
  OAI21_X1 U13914 ( .B1(n11462), .B2(n14955), .A(n14954), .ZN(n11467) );
  OAI22_X1 U13915 ( .A1(n14957), .A2(n12638), .B1(n15081), .B2(n8927), .ZN(
        n11463) );
  AOI21_X1 U13916 ( .B1(n11467), .B2(n15081), .A(n11463), .ZN(n11464) );
  INV_X1 U13917 ( .A(n11464), .ZN(P3_U3417) );
  OAI22_X1 U13918 ( .A1(n12585), .A2(n14957), .B1(n15096), .B2(n11465), .ZN(
        n11466) );
  AOI21_X1 U13919 ( .B1(n11467), .B2(n15096), .A(n11466), .ZN(n11468) );
  INV_X1 U13920 ( .A(n11468), .ZN(P3_U3468) );
  CLKBUF_X1 U13921 ( .A(n11469), .Z(n11470) );
  XNOR2_X1 U13922 ( .A(n11470), .B(n11472), .ZN(n11595) );
  OAI21_X1 U13923 ( .B1(n11473), .B2(n11472), .A(n11471), .ZN(n11474) );
  INV_X1 U13924 ( .A(n11474), .ZN(n11593) );
  INV_X1 U13925 ( .A(n14032), .ZN(n13987) );
  OAI211_X1 U13926 ( .C1(n11591), .C2(n11475), .A(n14617), .B(n14415), .ZN(
        n11590) );
  NAND2_X1 U13927 ( .A1(n13770), .A2(n14387), .ZN(n11476) );
  OAI21_X1 U13928 ( .B1(n13495), .B2(n14385), .A(n11476), .ZN(n11729) );
  INV_X1 U13929 ( .A(n11729), .ZN(n11589) );
  INV_X1 U13930 ( .A(n11477), .ZN(n11731) );
  OAI22_X1 U13931 ( .A1(n14638), .A2(n11589), .B1(n11731), .B2(n14612), .ZN(
        n11479) );
  NOR2_X1 U13932 ( .A1(n11591), .A2(n14640), .ZN(n11478) );
  AOI211_X1 U13933 ( .C1(n14648), .C2(P1_REG2_REG_13__SCAN_IN), .A(n11479), 
        .B(n11478), .ZN(n11480) );
  OAI21_X1 U13934 ( .B1(n14011), .B2(n11590), .A(n11480), .ZN(n11481) );
  AOI21_X1 U13935 ( .B1(n11593), .B2(n13987), .A(n11481), .ZN(n11482) );
  OAI21_X1 U13936 ( .B1(n11595), .B2(n14016), .A(n11482), .ZN(P1_U3280) );
  AOI21_X1 U13937 ( .B1(n11485), .B2(n11484), .A(n11483), .ZN(n11492) );
  NOR2_X1 U13938 ( .A1(n12172), .A2(n12140), .ZN(n11486) );
  AOI211_X1 U13939 ( .C1(n12170), .C2(n14968), .A(n11487), .B(n11486), .ZN(
        n11488) );
  OAI21_X1 U13940 ( .B1(n12177), .B2(n14957), .A(n11488), .ZN(n11489) );
  AOI21_X1 U13941 ( .B1(n11490), .B2(n12174), .A(n11489), .ZN(n11491) );
  OAI21_X1 U13942 ( .B1(n11492), .B2(n12153), .A(n11491), .ZN(P3_U3171) );
  AOI211_X1 U13943 ( .C1(n11495), .C2(n14880), .A(n11494), .B(n11493), .ZN(
        n11500) );
  INV_X1 U13944 ( .A(n13432), .ZN(n13434) );
  INV_X1 U13945 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11496) );
  NOR2_X1 U13946 ( .A1(n15282), .A2(n11496), .ZN(n11497) );
  AOI21_X1 U13947 ( .B1(n12883), .B2(n13434), .A(n11497), .ZN(n11498) );
  OAI21_X1 U13948 ( .B1(n11500), .B2(n14899), .A(n11498), .ZN(P2_U3466) );
  AOI22_X1 U13949 ( .A1(n12883), .A2(n13379), .B1(n14910), .B2(
        P2_REG1_REG_12__SCAN_IN), .ZN(n11499) );
  OAI21_X1 U13950 ( .B1(n11500), .B2(n14910), .A(n11499), .ZN(P2_U3511) );
  OAI211_X1 U13951 ( .C1(n11508), .C2(n11502), .A(n11501), .B(n15039), .ZN(
        n11504) );
  AOI22_X1 U13952 ( .A1(n12185), .A2(n15034), .B1(n15035), .B2(n12183), .ZN(
        n11503) );
  AND2_X1 U13953 ( .A1(n11504), .A2(n11503), .ZN(n14365) );
  AND2_X1 U13954 ( .A1(n11505), .A2(n15023), .ZN(n14361) );
  INV_X1 U13955 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11521) );
  INV_X1 U13956 ( .A(n12144), .ZN(n11506) );
  OAI22_X1 U13957 ( .A1(n15050), .A2(n11521), .B1(n11506), .B2(n15012), .ZN(
        n11507) );
  AOI21_X1 U13958 ( .B1(n15000), .B2(n14361), .A(n11507), .ZN(n11513) );
  NAND2_X1 U13959 ( .A1(n11509), .A2(n11508), .ZN(n11510) );
  NAND2_X1 U13960 ( .A1(n11511), .A2(n11510), .ZN(n14363) );
  NAND2_X1 U13961 ( .A1(n14363), .A2(n12520), .ZN(n11512) );
  OAI211_X1 U13962 ( .C1(n14365), .C2(n14334), .A(n11513), .B(n11512), .ZN(
        P3_U3222) );
  OAI222_X1 U13963 ( .A1(n13459), .A2(n11557), .B1(n11515), .B2(P2_U3088), 
        .C1(n11514), .C2(n13464), .ZN(P2_U3306) );
  OR2_X1 U13964 ( .A1(n11529), .A2(n11516), .ZN(n11517) );
  AOI21_X1 U13965 ( .B1(n11521), .B2(n11519), .A(n11604), .ZN(n11537) );
  INV_X1 U13966 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11520) );
  MUX2_X1 U13967 ( .A(n11521), .B(n11520), .S(n12198), .Z(n11522) );
  NAND2_X1 U13968 ( .A1(n11522), .A2(n11610), .ZN(n11617) );
  OAI21_X1 U13969 ( .B1(n11522), .B2(n11610), .A(n11617), .ZN(n11524) );
  AOI21_X1 U13970 ( .B1(n11524), .B2(n11523), .A(n11615), .ZN(n11527) );
  NOR2_X1 U13971 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11525), .ZN(n12138) );
  AOI21_X1 U13972 ( .B1(n14921), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n12138), 
        .ZN(n11526) );
  OAI21_X1 U13973 ( .B1(n11527), .B2(n14943), .A(n11526), .ZN(n11535) );
  OR2_X1 U13974 ( .A1(n11529), .A2(n11528), .ZN(n11530) );
  AOI21_X1 U13975 ( .B1(n11520), .B2(n11532), .A(n11611), .ZN(n11533) );
  NOR2_X1 U13976 ( .A1(n11533), .A2(n14937), .ZN(n11534) );
  AOI211_X1 U13977 ( .C1(n14948), .C2(n11610), .A(n11535), .B(n11534), .ZN(
        n11536) );
  OAI21_X1 U13978 ( .B1(n11537), .B2(n14940), .A(n11536), .ZN(P3_U3193) );
  INV_X1 U13979 ( .A(n11538), .ZN(n11539) );
  AOI21_X1 U13980 ( .B1(n11541), .B2(n11540), .A(n11539), .ZN(n11548) );
  NAND2_X1 U13981 ( .A1(n12770), .A2(n11542), .ZN(n11544) );
  OAI211_X1 U13982 ( .C1(n11545), .C2(n12751), .A(n11544), .B(n11543), .ZN(
        n11546) );
  AOI21_X1 U13983 ( .B1(n12875), .B2(n14381), .A(n11546), .ZN(n11547) );
  OAI21_X1 U13984 ( .B1(n11548), .B2(n12759), .A(n11547), .ZN(P2_U3208) );
  AOI21_X1 U13985 ( .B1(n14362), .B2(n11550), .A(n11549), .ZN(n11555) );
  OAI22_X1 U13986 ( .A1(n12585), .A2(n11671), .B1(n15096), .B2(n11528), .ZN(
        n11551) );
  INV_X1 U13987 ( .A(n11551), .ZN(n11552) );
  OAI21_X1 U13988 ( .B1(n11555), .B2(n15094), .A(n11552), .ZN(P3_U3469) );
  OAI22_X1 U13989 ( .A1(n11671), .A2(n12638), .B1(n15081), .B2(n8942), .ZN(
        n11553) );
  INV_X1 U13990 ( .A(n11553), .ZN(n11554) );
  OAI21_X1 U13991 ( .B1(n11555), .B2(n15080), .A(n11554), .ZN(P3_U3420) );
  OAI222_X1 U13992 ( .A1(P1_U3086), .A2(n11558), .B1(n14166), .B2(n11557), 
        .C1(n11556), .C2(n14163), .ZN(P1_U3334) );
  OR2_X1 U13993 ( .A1(n14380), .A2(n13057), .ZN(n11652) );
  NAND2_X1 U13994 ( .A1(n14380), .A2(n13057), .ZN(n11650) );
  NAND2_X1 U13995 ( .A1(n11652), .A2(n11650), .ZN(n13011) );
  XOR2_X1 U13996 ( .A(n13011), .B(n11648), .Z(n11563) );
  OR2_X1 U13997 ( .A1(n12887), .A2(n12773), .ZN(n11562) );
  NAND2_X1 U13998 ( .A1(n13036), .A2(n13058), .ZN(n11561) );
  NAND2_X1 U13999 ( .A1(n11562), .A2(n11561), .ZN(n14379) );
  AOI21_X1 U14000 ( .B1(n11563), .B2(n13198), .A(n14379), .ZN(n13382) );
  INV_X1 U14001 ( .A(n11564), .ZN(n11565) );
  AND2_X1 U14002 ( .A1(n12892), .A2(n11564), .ZN(n11654) );
  AOI211_X1 U14003 ( .C1(n14380), .C2(n11565), .A(n13231), .B(n11654), .ZN(
        n13381) );
  INV_X1 U14004 ( .A(n14383), .ZN(n11566) );
  AOI22_X1 U14005 ( .A1(n13298), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11566), 
        .B2(n13289), .ZN(n11567) );
  OAI21_X1 U14006 ( .B1(n12892), .B2(n13293), .A(n11567), .ZN(n11572) );
  NAND2_X1 U14007 ( .A1(n13386), .A2(n13058), .ZN(n11569) );
  NOR2_X1 U14008 ( .A1(n13386), .A2(n13058), .ZN(n11568) );
  XOR2_X1 U14009 ( .A(n13011), .B(n11653), .Z(n13384) );
  NOR2_X1 U14010 ( .A1(n13384), .A2(n13238), .ZN(n11571) );
  AOI211_X1 U14011 ( .C1(n13381), .C2(n13288), .A(n11572), .B(n11571), .ZN(
        n11573) );
  OAI21_X1 U14012 ( .B1(n13298), .B2(n13382), .A(n11573), .ZN(P2_U3251) );
  INV_X1 U14013 ( .A(n11575), .ZN(n11577) );
  NAND2_X1 U14014 ( .A1(n11577), .A2(n11576), .ZN(n11578) );
  XNOR2_X1 U14015 ( .A(n11579), .B(n11578), .ZN(n11586) );
  NAND2_X1 U14016 ( .A1(n12770), .A2(n11580), .ZN(n11582) );
  OAI211_X1 U14017 ( .C1(n11583), .C2(n12751), .A(n11582), .B(n11581), .ZN(
        n11584) );
  AOI21_X1 U14018 ( .B1(n12883), .B2(n14381), .A(n11584), .ZN(n11585) );
  OAI21_X1 U14019 ( .B1(n11586), .B2(n12759), .A(n11585), .ZN(P2_U3196) );
  INV_X1 U14020 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11597) );
  OAI211_X1 U14021 ( .C1(n11591), .C2(n14717), .A(n11590), .B(n11589), .ZN(
        n11592) );
  AOI21_X1 U14022 ( .B1(n11593), .B2(n14630), .A(n11592), .ZN(n11594) );
  OAI21_X1 U14023 ( .B1(n14442), .B2(n11595), .A(n11594), .ZN(n11598) );
  NAND2_X1 U14024 ( .A1(n11598), .A2(n14740), .ZN(n11596) );
  OAI21_X1 U14025 ( .B1(n14740), .B2(n11597), .A(n11596), .ZN(P1_U3541) );
  INV_X1 U14026 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11600) );
  NAND2_X1 U14027 ( .A1(n11598), .A2(n14724), .ZN(n11599) );
  OAI21_X1 U14028 ( .B1(n14724), .B2(n11600), .A(n11599), .ZN(P1_U3498) );
  NAND2_X1 U14029 ( .A1(n11618), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n11601) );
  OAI21_X1 U14030 ( .B1(n11618), .B2(P3_REG2_REG_12__SCAN_IN), .A(n11601), 
        .ZN(n11602) );
  INV_X1 U14031 ( .A(n11602), .ZN(n11608) );
  NOR2_X1 U14032 ( .A1(n11610), .A2(n11603), .ZN(n11605) );
  INV_X1 U14033 ( .A(n11780), .ZN(n11606) );
  AOI21_X1 U14034 ( .B1(n11608), .B2(n11607), .A(n11606), .ZN(n11626) );
  NOR2_X1 U14035 ( .A1(n11610), .A2(n11609), .ZN(n11612) );
  NAND2_X1 U14036 ( .A1(n11618), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n11613) );
  OAI21_X1 U14037 ( .B1(n11618), .B2(P3_REG1_REG_12__SCAN_IN), .A(n11613), 
        .ZN(n11614) );
  OAI21_X1 U14038 ( .B1(n7081), .B2(n11614), .A(n11784), .ZN(n11624) );
  MUX2_X1 U14039 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12198), .Z(n11788) );
  XNOR2_X1 U14040 ( .A(n11788), .B(n11787), .ZN(n11790) );
  INV_X1 U14041 ( .A(n11615), .ZN(n11616) );
  XNOR2_X1 U14042 ( .A(n11790), .B(n11789), .ZN(n11622) );
  NAND2_X1 U14043 ( .A1(n14948), .A2(n11618), .ZN(n11621) );
  NOR2_X1 U14044 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11619), .ZN(n12064) );
  AOI21_X1 U14045 ( .B1(n14921), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12064), 
        .ZN(n11620) );
  OAI211_X1 U14046 ( .C1(n11622), .C2(n14943), .A(n11621), .B(n11620), .ZN(
        n11623) );
  AOI21_X1 U14047 ( .B1(n11624), .B2(n14924), .A(n11623), .ZN(n11625) );
  OAI21_X1 U14048 ( .B1(n11626), .B2(n14940), .A(n11625), .ZN(P3_U3194) );
  NAND2_X1 U14049 ( .A1(n14453), .A2(n13587), .ZN(n11628) );
  NAND2_X1 U14050 ( .A1(n13771), .A2(n13555), .ZN(n11627) );
  NAND2_X1 U14051 ( .A1(n11628), .A2(n11627), .ZN(n11629) );
  XNOR2_X1 U14052 ( .A(n11629), .B(n13561), .ZN(n11673) );
  AND2_X1 U14053 ( .A1(n13771), .A2(n10463), .ZN(n11630) );
  AOI21_X1 U14054 ( .B1(n14453), .B2(n6460), .A(n11630), .ZN(n11672) );
  XNOR2_X1 U14055 ( .A(n11673), .B(n11672), .ZN(n11641) );
  INV_X1 U14056 ( .A(n11633), .ZN(n11634) );
  NAND2_X1 U14057 ( .A1(n11635), .A2(n11634), .ZN(n11636) );
  INV_X1 U14058 ( .A(n11681), .ZN(n11639) );
  AOI21_X1 U14059 ( .B1(n11641), .B2(n11640), .A(n11639), .ZN(n11647) );
  NAND2_X1 U14060 ( .A1(n13739), .A2(n11642), .ZN(n11643) );
  NAND2_X1 U14061 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14505)
         );
  OAI211_X1 U14062 ( .C1(n11644), .C2(n13737), .A(n11643), .B(n14505), .ZN(
        n11645) );
  AOI21_X1 U14063 ( .B1(n14453), .B2(n14398), .A(n11645), .ZN(n11646) );
  OAI21_X1 U14064 ( .B1(n11647), .B2(n13751), .A(n11646), .ZN(P1_U3236) );
  XNOR2_X1 U14065 ( .A(n13435), .B(n12887), .ZN(n13015) );
  INV_X1 U14066 ( .A(n13015), .ZN(n11703) );
  XNOR2_X1 U14067 ( .A(n11704), .B(n11703), .ZN(n11649) );
  INV_X1 U14068 ( .A(n12773), .ZN(n12749) );
  AOI22_X1 U14069 ( .A1(n13055), .A2(n12749), .B1(n13036), .B2(n13057), .ZN(
        n11837) );
  OAI21_X1 U14070 ( .B1(n11649), .B2(n13281), .A(n11837), .ZN(n13376) );
  INV_X1 U14071 ( .A(n13376), .ZN(n11661) );
  INV_X1 U14072 ( .A(n11650), .ZN(n11651) );
  XNOR2_X1 U14073 ( .A(n11713), .B(n13015), .ZN(n13378) );
  INV_X1 U14074 ( .A(n11654), .ZN(n11656) );
  INV_X1 U14075 ( .A(n11710), .ZN(n11655) );
  AOI211_X1 U14076 ( .C1(n13435), .C2(n11656), .A(n13231), .B(n11655), .ZN(
        n13377) );
  NAND2_X1 U14077 ( .A1(n13377), .A2(n13288), .ZN(n11658) );
  AOI22_X1 U14078 ( .A1(n13298), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11840), 
        .B2(n13289), .ZN(n11657) );
  OAI211_X1 U14079 ( .C1(n12886), .C2(n13293), .A(n11658), .B(n11657), .ZN(
        n11659) );
  AOI21_X1 U14080 ( .B1(n13295), .B2(n13378), .A(n11659), .ZN(n11660) );
  OAI21_X1 U14081 ( .B1(n13298), .B2(n11661), .A(n11660), .ZN(P2_U3250) );
  OAI211_X1 U14082 ( .C1(n11664), .C2(n11663), .A(n11662), .B(n14914), .ZN(
        n11670) );
  NAND2_X1 U14083 ( .A1(n12170), .A2(n12186), .ZN(n11665) );
  OAI211_X1 U14084 ( .C1(n12172), .C2(n14347), .A(n11666), .B(n11665), .ZN(
        n11667) );
  AOI21_X1 U14085 ( .B1(n12174), .B2(n11668), .A(n11667), .ZN(n11669) );
  OAI211_X1 U14086 ( .C1(n12177), .C2(n11671), .A(n11670), .B(n11669), .ZN(
        P3_U3157) );
  NAND2_X1 U14087 ( .A1(n11673), .A2(n11672), .ZN(n11679) );
  AND2_X1 U14088 ( .A1(n11681), .A2(n11679), .ZN(n11683) );
  NAND2_X1 U14089 ( .A1(n11678), .A2(n13587), .ZN(n11675) );
  NAND2_X1 U14090 ( .A1(n13770), .A2(n13555), .ZN(n11674) );
  NAND2_X1 U14091 ( .A1(n11675), .A2(n11674), .ZN(n11676) );
  XNOR2_X1 U14092 ( .A(n11676), .B(n13625), .ZN(n11722) );
  AND2_X1 U14093 ( .A1(n13770), .A2(n10463), .ZN(n11677) );
  AOI21_X1 U14094 ( .B1(n11678), .B2(n6460), .A(n11677), .ZN(n11720) );
  XNOR2_X1 U14095 ( .A(n11722), .B(n11720), .ZN(n11682) );
  AND2_X1 U14096 ( .A1(n11682), .A2(n11679), .ZN(n11680) );
  OAI211_X1 U14097 ( .C1(n11683), .C2(n11682), .A(n14395), .B(n11724), .ZN(
        n11689) );
  OAI21_X1 U14098 ( .B1(n13737), .B2(n11685), .A(n11684), .ZN(n11686) );
  AOI21_X1 U14099 ( .B1(n11687), .B2(n13739), .A(n11686), .ZN(n11688) );
  OAI211_X1 U14100 ( .C1(n6961), .C2(n13742), .A(n11689), .B(n11688), .ZN(
        P1_U3224) );
  OAI211_X1 U14101 ( .C1(n11692), .C2(n11691), .A(n11690), .B(n14376), .ZN(
        n11698) );
  OAI22_X1 U14102 ( .A1(n12751), .A2(n11694), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11693), .ZN(n11695) );
  AOI21_X1 U14103 ( .B1(n11696), .B2(n12770), .A(n11695), .ZN(n11697) );
  OAI211_X1 U14104 ( .C1(n12895), .C2(n12776), .A(n11698), .B(n11697), .ZN(
        P2_U3206) );
  INV_X1 U14105 ( .A(n11699), .ZN(n11700) );
  OAI222_X1 U14106 ( .A1(n11702), .A2(P3_U3151), .B1(n11881), .B2(n11701), 
        .C1(n11970), .C2(n11700), .ZN(P3_U3271) );
  INV_X1 U14107 ( .A(n13055), .ZN(n12719) );
  XNOR2_X1 U14108 ( .A(n13372), .B(n12719), .ZN(n12904) );
  OAI21_X1 U14109 ( .B1(n6476), .B2(n13013), .A(n11889), .ZN(n11708) );
  OR2_X1 U14110 ( .A1(n12755), .A2(n12773), .ZN(n11707) );
  NAND2_X1 U14111 ( .A1(n13056), .A2(n13036), .ZN(n11706) );
  NAND2_X1 U14112 ( .A1(n11707), .A2(n11706), .ZN(n12693) );
  AOI21_X1 U14113 ( .B1(n11708), .B2(n13198), .A(n12693), .ZN(n13373) );
  INV_X1 U14114 ( .A(n13286), .ZN(n11709) );
  AOI211_X1 U14115 ( .C1(n13372), .C2(n11710), .A(n13231), .B(n11709), .ZN(
        n13371) );
  INV_X1 U14116 ( .A(n12696), .ZN(n11711) );
  AOI22_X1 U14117 ( .A1(n13298), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n11711), 
        .B2(n13289), .ZN(n11712) );
  OAI21_X1 U14118 ( .B1(n7042), .B2(n13293), .A(n11712), .ZN(n11718) );
  NAND2_X1 U14119 ( .A1(n12886), .A2(n12887), .ZN(n11714) );
  NAND2_X1 U14120 ( .A1(n11715), .A2(n13013), .ZN(n11716) );
  NAND2_X1 U14121 ( .A1(n11917), .A2(n11716), .ZN(n13375) );
  NOR2_X1 U14122 ( .A1(n13375), .A2(n13238), .ZN(n11717) );
  AOI211_X1 U14123 ( .C1(n13371), .C2(n13288), .A(n11718), .B(n11717), .ZN(
        n11719) );
  OAI21_X1 U14124 ( .B1(n13298), .B2(n13373), .A(n11719), .ZN(P2_U3249) );
  INV_X1 U14125 ( .A(n11720), .ZN(n11721) );
  NAND2_X1 U14126 ( .A1(n11722), .A2(n11721), .ZN(n11723) );
  NAND2_X1 U14127 ( .A1(n11733), .A2(n13587), .ZN(n11726) );
  NAND2_X1 U14128 ( .A1(n14388), .A2(n13555), .ZN(n11725) );
  NAND2_X1 U14129 ( .A1(n11726), .A2(n11725), .ZN(n11727) );
  XNOR2_X1 U14130 ( .A(n11727), .B(n13625), .ZN(n13490) );
  AND2_X1 U14131 ( .A1(n14388), .A2(n10463), .ZN(n11728) );
  AOI21_X1 U14132 ( .B1(n11733), .B2(n6460), .A(n11728), .ZN(n13488) );
  XNOR2_X1 U14133 ( .A(n13490), .B(n13488), .ZN(n13486) );
  XNOR2_X1 U14134 ( .A(n13487), .B(n13486), .ZN(n11735) );
  NAND2_X1 U14135 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14522)
         );
  NAND2_X1 U14136 ( .A1(n14397), .A2(n11729), .ZN(n11730) );
  OAI211_X1 U14137 ( .C1(n14401), .C2(n11731), .A(n14522), .B(n11730), .ZN(
        n11732) );
  AOI21_X1 U14138 ( .B1(n11733), .B2(n14398), .A(n11732), .ZN(n11734) );
  OAI21_X1 U14139 ( .B1(n11735), .B2(n13751), .A(n11734), .ZN(P1_U3234) );
  INV_X1 U14140 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12000) );
  MUX2_X1 U14141 ( .A(n12000), .B(P2_REG2_REG_17__SCAN_IN), .S(n12006), .Z(
        n11995) );
  OAI21_X1 U14142 ( .B1(n11444), .B2(n11737), .A(n11736), .ZN(n11996) );
  XOR2_X1 U14143 ( .A(n11995), .B(n11996), .Z(n11748) );
  AOI21_X1 U14144 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n11739), .A(n11738), 
        .ZN(n11741) );
  XNOR2_X1 U14145 ( .A(n12006), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n11740) );
  NOR2_X1 U14146 ( .A1(n11741), .A2(n11740), .ZN(n12005) );
  AOI211_X1 U14147 ( .C1(n11741), .C2(n11740), .A(n14813), .B(n12005), .ZN(
        n11746) );
  NOR2_X1 U14148 ( .A1(n14827), .A2(n11999), .ZN(n11745) );
  AND2_X1 U14149 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n11744) );
  INV_X1 U14150 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n11742) );
  NOR2_X1 U14151 ( .A1(n14811), .A2(n11742), .ZN(n11743) );
  NOR4_X1 U14152 ( .A1(n11746), .A2(n11745), .A3(n11744), .A4(n11743), .ZN(
        n11747) );
  OAI21_X1 U14153 ( .B1(n14823), .B2(n11748), .A(n11747), .ZN(P2_U3231) );
  INV_X1 U14154 ( .A(n11749), .ZN(n11750) );
  AOI21_X1 U14155 ( .B1(n11753), .B2(n11751), .A(n11750), .ZN(n14443) );
  OAI211_X1 U14156 ( .C1(n11754), .C2(n11753), .A(n11752), .B(n14630), .ZN(
        n14440) );
  INV_X1 U14157 ( .A(n14440), .ZN(n11756) );
  NAND2_X1 U14158 ( .A1(n13767), .A2(n13732), .ZN(n11755) );
  OAI21_X1 U14159 ( .B1(n13495), .B2(n14633), .A(n11755), .ZN(n14438) );
  OAI21_X1 U14160 ( .B1(n11756), .B2(n14438), .A(n14008), .ZN(n11762) );
  INV_X1 U14161 ( .A(n11772), .ZN(n11757) );
  AOI211_X1 U14162 ( .C1(n14439), .C2(n14416), .A(n14675), .B(n11757), .ZN(
        n14437) );
  INV_X1 U14163 ( .A(n14439), .ZN(n11759) );
  AOI22_X1 U14164 ( .A1(n14638), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13745), 
        .B2(n14637), .ZN(n11758) );
  OAI21_X1 U14165 ( .B1(n11759), .B2(n14640), .A(n11758), .ZN(n11760) );
  AOI21_X1 U14166 ( .B1(n14437), .B2(n14644), .A(n11760), .ZN(n11761) );
  OAI211_X1 U14167 ( .C1(n14443), .C2(n14016), .A(n11762), .B(n11761), .ZN(
        P1_U3278) );
  INV_X1 U14168 ( .A(n11763), .ZN(n11765) );
  OAI222_X1 U14169 ( .A1(n11970), .A2(n11765), .B1(P3_U3151), .B2(n11764), 
        .C1(n15233), .C2(n11881), .ZN(P3_U3270) );
  INV_X1 U14170 ( .A(n11766), .ZN(n11767) );
  AOI21_X1 U14171 ( .B1(n7275), .B2(n11768), .A(n11767), .ZN(n14433) );
  INV_X1 U14172 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11771) );
  OAI22_X1 U14173 ( .A1(n7279), .A2(n14385), .B1(n14386), .B2(n14633), .ZN(
        n14429) );
  INV_X1 U14174 ( .A(n13665), .ZN(n11769) );
  AOI22_X1 U14175 ( .A1(n14008), .A2(n14429), .B1(n11769), .B2(n14637), .ZN(
        n11770) );
  OAI21_X1 U14176 ( .B1(n11771), .B2(n14008), .A(n11770), .ZN(n11775) );
  AOI21_X1 U14177 ( .B1(n11772), .B2(n14430), .A(n14675), .ZN(n11773) );
  NAND2_X1 U14178 ( .A1(n11773), .A2(n11827), .ZN(n14431) );
  NOR2_X1 U14179 ( .A1(n14431), .A2(n14011), .ZN(n11774) );
  AOI211_X1 U14180 ( .C1(n14409), .C2(n14430), .A(n11775), .B(n11774), .ZN(
        n11778) );
  XNOR2_X1 U14181 ( .A(n11776), .B(n7275), .ZN(n14435) );
  NAND2_X1 U14182 ( .A1(n14435), .A2(n14419), .ZN(n11777) );
  OAI211_X1 U14183 ( .C1(n14433), .C2(n14032), .A(n11778), .B(n11777), .ZN(
        P1_U3277) );
  INV_X1 U14184 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11782) );
  NAND2_X1 U14185 ( .A1(n11787), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n11779) );
  AOI21_X1 U14186 ( .B1(n11782), .B2(n11781), .A(n12193), .ZN(n11800) );
  INV_X1 U14187 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12583) );
  NAND2_X1 U14188 ( .A1(n11787), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n11783) );
  XNOR2_X1 U14189 ( .A(n12210), .B(n12209), .ZN(n11785) );
  AOI21_X1 U14190 ( .B1(n12583), .B2(n11785), .A(n12211), .ZN(n11786) );
  NOR2_X1 U14191 ( .A1(n11786), .A2(n14937), .ZN(n11798) );
  MUX2_X1 U14192 ( .A(n11782), .B(n12583), .S(n12198), .Z(n12195) );
  XNOR2_X1 U14193 ( .A(n12195), .B(n12210), .ZN(n11793) );
  NAND2_X1 U14194 ( .A1(n11788), .A2(n11787), .ZN(n11791) );
  AOI21_X1 U14195 ( .B1(n11793), .B2(n11792), .A(n12200), .ZN(n11796) );
  NAND2_X1 U14196 ( .A1(n14948), .A2(n12210), .ZN(n11795) );
  AND2_X1 U14197 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12121) );
  AOI21_X1 U14198 ( .B1(n14921), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12121), 
        .ZN(n11794) );
  OAI211_X1 U14199 ( .C1(n11796), .C2(n14943), .A(n11795), .B(n11794), .ZN(
        n11797) );
  NOR2_X1 U14200 ( .A1(n11798), .A2(n11797), .ZN(n11799) );
  OAI21_X1 U14201 ( .B1(n11800), .B2(n14940), .A(n11799), .ZN(P3_U3195) );
  NAND2_X1 U14202 ( .A1(n11801), .A2(n15039), .ZN(n11805) );
  AOI21_X1 U14203 ( .B1(n12508), .B2(n11802), .A(n11806), .ZN(n11804) );
  AOI22_X1 U14204 ( .A1(n14344), .A2(n15034), .B1(n15035), .B2(n12482), .ZN(
        n11803) );
  OAI21_X1 U14205 ( .B1(n11805), .B2(n11804), .A(n11803), .ZN(n12577) );
  INV_X1 U14206 ( .A(n12577), .ZN(n11811) );
  XNOR2_X1 U14207 ( .A(n11807), .B(n11806), .ZN(n12578) );
  INV_X1 U14208 ( .A(n12031), .ZN(n12633) );
  AOI22_X1 U14209 ( .A1(n14334), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15046), 
        .B2(n12026), .ZN(n11808) );
  OAI21_X1 U14210 ( .B1(n12633), .B2(n14958), .A(n11808), .ZN(n11809) );
  AOI21_X1 U14211 ( .B1(n12578), .B2(n12520), .A(n11809), .ZN(n11810) );
  OAI21_X1 U14212 ( .B1(n11811), .B2(n14334), .A(n11810), .ZN(P3_U3219) );
  NAND2_X1 U14213 ( .A1(n11816), .A2(n13450), .ZN(n11813) );
  OR2_X1 U14214 ( .A1(n11812), .A2(P2_U3088), .ZN(n13040) );
  OAI211_X1 U14215 ( .C1(n11814), .C2(n13464), .A(n11813), .B(n13040), .ZN(
        P2_U3304) );
  NAND2_X1 U14216 ( .A1(n11816), .A2(n11815), .ZN(n11818) );
  OAI211_X1 U14217 ( .C1(n11819), .C2(n14163), .A(n11818), .B(n11817), .ZN(
        P1_U3332) );
  XNOR2_X1 U14218 ( .A(n11820), .B(n11821), .ZN(n14426) );
  XNOR2_X1 U14219 ( .A(n11822), .B(n11821), .ZN(n14428) );
  NAND2_X1 U14220 ( .A1(n14428), .A2(n13987), .ZN(n11832) );
  INV_X1 U14221 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13832) );
  OAI22_X1 U14222 ( .A1(n13530), .A2(n14385), .B1(n11823), .B2(n14633), .ZN(
        n14422) );
  INV_X1 U14223 ( .A(n13670), .ZN(n11824) );
  AOI22_X1 U14224 ( .A1(n14422), .A2(n14008), .B1(n11824), .B2(n14637), .ZN(
        n11825) );
  OAI21_X1 U14225 ( .B1(n13832), .B2(n14008), .A(n11825), .ZN(n11830) );
  INV_X1 U14226 ( .A(n11826), .ZN(n14040) );
  AOI21_X1 U14227 ( .B1(n11827), .B2(n14423), .A(n14675), .ZN(n11828) );
  NAND2_X1 U14228 ( .A1(n14040), .A2(n11828), .ZN(n14424) );
  NOR2_X1 U14229 ( .A1(n14424), .A2(n14011), .ZN(n11829) );
  AOI211_X1 U14230 ( .C1(n14409), .C2(n14423), .A(n11830), .B(n11829), .ZN(
        n11831) );
  OAI211_X1 U14231 ( .C1(n14426), .C2(n14016), .A(n11832), .B(n11831), .ZN(
        P1_U3276) );
  AOI22_X1 U14232 ( .A1(n11833), .A2(n14376), .B1(n12744), .B2(n13056), .ZN(
        n11843) );
  INV_X1 U14233 ( .A(n11835), .ZN(n11842) );
  OAI22_X1 U14234 ( .A1(n12751), .A2(n11837), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11836), .ZN(n11839) );
  NOR2_X1 U14235 ( .A1(n12886), .A2(n12776), .ZN(n11838) );
  AOI211_X1 U14236 ( .C1(n12770), .C2(n11840), .A(n11839), .B(n11838), .ZN(
        n11841) );
  OAI21_X1 U14237 ( .B1(n11843), .B2(n11842), .A(n11841), .ZN(P2_U3213) );
  INV_X1 U14238 ( .A(n11844), .ZN(n11848) );
  OAI222_X1 U14239 ( .A1(n13459), .A2(n11848), .B1(P2_U3088), .B2(n11846), 
        .C1(n11845), .C2(n13464), .ZN(P2_U3303) );
  INV_X1 U14240 ( .A(n11847), .ZN(n11849) );
  OAI222_X1 U14241 ( .A1(P1_U3086), .A2(n11849), .B1(n14166), .B2(n11848), 
        .C1(n15119), .C2(n14163), .ZN(P1_U3331) );
  INV_X1 U14242 ( .A(n11850), .ZN(n11851) );
  OAI222_X1 U14243 ( .A1(n11853), .A2(P3_U3151), .B1(n11881), .B2(n11852), 
        .C1(n11970), .C2(n11851), .ZN(P3_U3269) );
  OR2_X1 U14244 ( .A1(n11865), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11855) );
  NAND2_X1 U14245 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n11865), .ZN(n11854) );
  NAND2_X1 U14246 ( .A1(n11855), .A2(n11854), .ZN(n14513) );
  OR2_X1 U14247 ( .A1(n11862), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11856) );
  NAND2_X1 U14248 ( .A1(n11857), .A2(n11856), .ZN(n14514) );
  MUX2_X1 U14249 ( .A(n11858), .B(P1_REG2_REG_14__SCAN_IN), .S(n14525), .Z(
        n14527) );
  INV_X1 U14250 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11859) );
  NAND2_X1 U14251 ( .A1(n11860), .A2(n11859), .ZN(n13828) );
  OAI21_X1 U14252 ( .B1(n11860), .B2(n11859), .A(n13828), .ZN(n11871) );
  INV_X1 U14253 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11861) );
  MUX2_X1 U14254 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n11861), .S(n14525), .Z(
        n14533) );
  OR2_X1 U14255 ( .A1(n11862), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11863) );
  NAND2_X1 U14256 ( .A1(n11864), .A2(n11863), .ZN(n14509) );
  MUX2_X1 U14257 ( .A(n11597), .B(P1_REG1_REG_13__SCAN_IN), .S(n11865), .Z(
        n14508) );
  NOR2_X1 U14258 ( .A1(n14509), .A2(n14508), .ZN(n14510) );
  NAND2_X1 U14259 ( .A1(n14533), .A2(n14532), .ZN(n14531) );
  OAI21_X1 U14260 ( .B1(n14525), .B2(P1_REG1_REG_14__SCAN_IN), .A(n14531), 
        .ZN(n13839) );
  INV_X1 U14261 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14445) );
  OAI21_X1 U14262 ( .B1(n11866), .B2(n14445), .A(n13841), .ZN(n11867) );
  NAND2_X1 U14263 ( .A1(n11867), .A2(n14558), .ZN(n11869) );
  NOR2_X1 U14264 ( .A1(n15104), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13746) );
  AOI21_X1 U14265 ( .B1(n14491), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n13746), 
        .ZN(n11868) );
  OAI211_X1 U14266 ( .C1(n14566), .C2(n13840), .A(n11869), .B(n11868), .ZN(
        n11870) );
  AOI21_X1 U14267 ( .B1(n14554), .B2(n11871), .A(n11870), .ZN(n11872) );
  INV_X1 U14268 ( .A(n11872), .ZN(P1_U3258) );
  INV_X1 U14269 ( .A(n11873), .ZN(n11874) );
  OAI222_X1 U14270 ( .A1(P3_U3151), .A2(n11876), .B1(n11881), .B2(n11875), 
        .C1(n11970), .C2(n11874), .ZN(P3_U3267) );
  INV_X1 U14271 ( .A(n11877), .ZN(n11880) );
  OAI222_X1 U14272 ( .A1(n11970), .A2(n11880), .B1(n11879), .B2(P3_U3151), 
        .C1(n11878), .C2(n11881), .ZN(P3_U3266) );
  OAI222_X1 U14273 ( .A1(n11884), .A2(P3_U3151), .B1(n11970), .B2(n11883), 
        .C1(n11882), .C2(n11881), .ZN(P3_U3265) );
  NAND2_X1 U14274 ( .A1(n13314), .A2(n12957), .ZN(n11885) );
  NAND2_X1 U14275 ( .A1(n13416), .A2(n13050), .ZN(n11896) );
  INV_X1 U14276 ( .A(n13050), .ZN(n11886) );
  NAND2_X1 U14277 ( .A1(n13194), .A2(n11886), .ZN(n11887) );
  NAND2_X1 U14278 ( .A1(n13372), .A2(n12719), .ZN(n11888) );
  OR2_X1 U14279 ( .A1(n13287), .A2(n12755), .ZN(n12912) );
  NAND2_X1 U14280 ( .A1(n13287), .A2(n12755), .ZN(n12913) );
  INV_X1 U14281 ( .A(n13053), .ZN(n12714) );
  AND2_X1 U14282 ( .A1(n13269), .A2(n12714), .ZN(n11890) );
  NAND2_X1 U14283 ( .A1(n13429), .A2(n13053), .ZN(n11891) );
  INV_X1 U14284 ( .A(n13052), .ZN(n12756) );
  NAND2_X1 U14285 ( .A1(n13251), .A2(n12756), .ZN(n13243) );
  XNOR2_X1 U14286 ( .A(n13353), .B(n12928), .ZN(n13220) );
  INV_X1 U14287 ( .A(n12928), .ZN(n11892) );
  NAND2_X1 U14288 ( .A1(n13353), .A2(n11892), .ZN(n11893) );
  NAND2_X1 U14289 ( .A1(n13420), .A2(n13051), .ZN(n11895) );
  INV_X1 U14290 ( .A(n13051), .ZN(n12735) );
  AND2_X1 U14291 ( .A1(n13212), .A2(n12735), .ZN(n11894) );
  XNOR2_X1 U14292 ( .A(n13182), .B(n12730), .ZN(n13179) );
  NAND2_X1 U14293 ( .A1(n13408), .A2(n13048), .ZN(n11897) );
  INV_X1 U14294 ( .A(n13048), .ZN(n11925) );
  NAND2_X1 U14295 ( .A1(n12946), .A2(n11925), .ZN(n11898) );
  NAND2_X1 U14296 ( .A1(n11897), .A2(n11898), .ZN(n13163) );
  INV_X1 U14297 ( .A(n13163), .ZN(n13159) );
  NAND2_X1 U14298 ( .A1(n13412), .A2(n13049), .ZN(n13156) );
  XNOR2_X1 U14299 ( .A(n13327), .B(n13047), .ZN(n13152) );
  INV_X1 U14300 ( .A(n13047), .ZN(n12772) );
  NAND2_X1 U14301 ( .A1(n13137), .A2(n13046), .ZN(n12988) );
  INV_X1 U14302 ( .A(n12988), .ZN(n11899) );
  INV_X1 U14303 ( .A(n13046), .ZN(n12654) );
  NAND2_X1 U14304 ( .A1(n13322), .A2(n12654), .ZN(n12987) );
  NAND2_X1 U14305 ( .A1(n13124), .A2(n12956), .ZN(n13101) );
  NAND2_X1 U14306 ( .A1(n12799), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11901) );
  XNOR2_X1 U14307 ( .A(n13308), .B(n12795), .ZN(n13020) );
  INV_X1 U14308 ( .A(P2_B_REG_SCAN_IN), .ZN(n11904) );
  NOR2_X1 U14309 ( .A1(n13454), .A2(n11904), .ZN(n11905) );
  NOR2_X1 U14310 ( .A1(n12773), .A2(n11905), .ZN(n13092) );
  NAND2_X1 U14311 ( .A1(n12785), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n11909) );
  NAND2_X1 U14312 ( .A1(n11906), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n11908) );
  NAND2_X1 U14313 ( .A1(n12786), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n11907) );
  AND3_X1 U14314 ( .A1(n11909), .A2(n11908), .A3(n11907), .ZN(n12794) );
  INV_X1 U14315 ( .A(n12794), .ZN(n13042) );
  AOI22_X1 U14316 ( .A1(n13044), .A2(n13036), .B1(n13092), .B2(n13042), .ZN(
        n11910) );
  AOI21_X2 U14317 ( .B1(n11912), .B2(n13198), .A(n11911), .ZN(n13310) );
  OR2_X1 U14318 ( .A1(n13353), .A2(n13249), .ZN(n13232) );
  NOR2_X2 U14319 ( .A1(n13212), .A2(n13232), .ZN(n13211) );
  NOR2_X2 U14320 ( .A1(n13322), .A2(n13147), .ZN(n13134) );
  AND2_X1 U14321 ( .A1(n13402), .A2(n13134), .ZN(n13122) );
  INV_X1 U14322 ( .A(n13108), .ZN(n11913) );
  AOI211_X1 U14323 ( .C1(n13308), .C2(n11913), .A(n13089), .B(n13096), .ZN(
        n13307) );
  AOI22_X1 U14324 ( .A1(n11914), .A2(n13289), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13298), .ZN(n11915) );
  OAI21_X1 U14325 ( .B1(n12796), .B2(n13293), .A(n11915), .ZN(n11927) );
  INV_X1 U14326 ( .A(n13201), .ZN(n13190) );
  XNOR2_X1 U14327 ( .A(n13212), .B(n13051), .ZN(n13016) );
  NAND2_X1 U14328 ( .A1(n13372), .A2(n13055), .ZN(n11916) );
  INV_X1 U14329 ( .A(n12755), .ZN(n13054) );
  NAND2_X1 U14330 ( .A1(n13287), .A2(n13054), .ZN(n11918) );
  XNOR2_X1 U14331 ( .A(n13269), .B(n12714), .ZN(n13266) );
  INV_X1 U14332 ( .A(n13266), .ZN(n11919) );
  NAND2_X1 U14333 ( .A1(n13429), .A2(n12714), .ZN(n11920) );
  NAND2_X1 U14334 ( .A1(n13251), .A2(n13052), .ZN(n12989) );
  OR2_X1 U14335 ( .A1(n13251), .A2(n13052), .ZN(n12990) );
  NOR2_X1 U14336 ( .A1(n13353), .A2(n12928), .ZN(n11921) );
  NAND2_X1 U14337 ( .A1(n13353), .A2(n12928), .ZN(n11922) );
  NAND2_X1 U14338 ( .A1(n13194), .A2(n13050), .ZN(n11924) );
  OAI22_X1 U14339 ( .A1(n13113), .A2(n13112), .B1(n13111), .B2(n12957), .ZN(
        n11926) );
  INV_X1 U14340 ( .A(n12783), .ZN(n11931) );
  OAI222_X1 U14341 ( .A1(n13459), .A2(n11931), .B1(n11929), .B2(P2_U3088), 
        .C1(n11928), .C2(n13464), .ZN(P2_U3297) );
  OAI222_X1 U14342 ( .A1(P1_U3086), .A2(n11932), .B1(n14171), .B2(n11931), 
        .C1(n11930), .C2(n14163), .ZN(P1_U3325) );
  NOR2_X1 U14343 ( .A1(n14419), .A2(n13987), .ZN(n11939) );
  OAI22_X1 U14344 ( .A1(n14648), .A2(n11934), .B1(n11933), .B2(n14612), .ZN(
        n11937) );
  AOI21_X1 U14345 ( .B1(n11935), .B2(n14640), .A(n14628), .ZN(n11936) );
  AOI211_X1 U14346 ( .C1(n14648), .C2(P1_REG2_REG_0__SCAN_IN), .A(n11937), .B(
        n11936), .ZN(n11938) );
  OAI21_X1 U14347 ( .B1(n11939), .B2(n9685), .A(n11938), .ZN(P1_U3293) );
  INV_X1 U14348 ( .A(n11940), .ZN(n11941) );
  OAI22_X1 U14349 ( .A1(n12765), .A2(n11942), .B1(n12759), .B2(n11941), .ZN(
        n11948) );
  AOI22_X1 U14350 ( .A1(n14378), .A2(n11943), .B1(n14381), .B2(n12815), .ZN(
        n11944) );
  OAI21_X1 U14351 ( .B1(n11946), .B2(n11945), .A(n11944), .ZN(n11947) );
  AOI21_X1 U14352 ( .B1(n11949), .B2(n11948), .A(n11947), .ZN(n11950) );
  OAI21_X1 U14353 ( .B1(n12759), .B2(n10495), .A(n11950), .ZN(P2_U3194) );
  XNOR2_X1 U14354 ( .A(n11952), .B(n11951), .ZN(n11960) );
  INV_X1 U14355 ( .A(n11960), .ZN(n11953) );
  NAND2_X1 U14356 ( .A1(n11953), .A2(n14914), .ZN(n11967) );
  INV_X1 U14357 ( .A(n11954), .ZN(n11955) );
  AOI22_X1 U14358 ( .A1(n12332), .A2(n12174), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11957) );
  NAND2_X1 U14359 ( .A1(n12179), .A2(n12170), .ZN(n11956) );
  OAI211_X1 U14360 ( .C1(n11958), .C2(n12172), .A(n11957), .B(n11956), .ZN(
        n11962) );
  NOR4_X1 U14361 ( .A1(n11960), .A2(n11959), .A3(n12153), .A4(n12179), .ZN(
        n11961) );
  AOI211_X1 U14362 ( .C1(n11963), .C2(n14918), .A(n11962), .B(n11961), .ZN(
        n11964) );
  OAI211_X1 U14363 ( .C1(n11967), .C2(n11966), .A(n11965), .B(n11964), .ZN(
        P3_U3160) );
  INV_X1 U14364 ( .A(n11968), .ZN(n11969) );
  OAI222_X1 U14365 ( .A1(P3_U3151), .A2(n12198), .B1(n11881), .B2(n11971), 
        .C1(n11970), .C2(n11969), .ZN(P3_U3268) );
  AOI22_X1 U14366 ( .A1(n11972), .A2(n14376), .B1(n12744), .B2(n13049), .ZN(
        n11977) );
  AOI22_X1 U14367 ( .A1(n13048), .A2(n12749), .B1(n13036), .B2(n13050), .ZN(
        n13173) );
  OAI22_X1 U14368 ( .A1(n13173), .A2(n12751), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11973), .ZN(n11975) );
  NOR2_X1 U14369 ( .A1(n13412), .A2(n12776), .ZN(n11974) );
  AOI211_X1 U14370 ( .C1(n12770), .C2(n13177), .A(n11975), .B(n11974), .ZN(
        n11976) );
  OAI21_X1 U14371 ( .B1(n11978), .B2(n11977), .A(n11976), .ZN(P2_U3188) );
  NAND2_X1 U14372 ( .A1(n14381), .A2(n12836), .ZN(n11980) );
  NAND2_X1 U14373 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n14769) );
  OAI211_X1 U14374 ( .C1(n11981), .C2(n12751), .A(n11980), .B(n14769), .ZN(
        n11989) );
  NOR3_X1 U14375 ( .A1(n12765), .A2(n11983), .A3(n11982), .ZN(n11984) );
  AOI21_X1 U14376 ( .B1(n11985), .B2(n14376), .A(n11984), .ZN(n11987) );
  NOR2_X1 U14377 ( .A1(n11987), .A2(n11986), .ZN(n11988) );
  AOI211_X1 U14378 ( .C1(n12770), .C2(n11990), .A(n11989), .B(n11988), .ZN(
        n11991) );
  OAI21_X1 U14379 ( .B1(n12759), .B2(n12708), .A(n11991), .ZN(P2_U3202) );
  INV_X1 U14380 ( .A(n11995), .ZN(n11997) );
  NAND2_X1 U14381 ( .A1(n11997), .A2(n11996), .ZN(n11998) );
  OAI21_X1 U14382 ( .B1(n12000), .B2(n11999), .A(n11998), .ZN(n12001) );
  NOR2_X1 U14383 ( .A1(n12002), .A2(n12001), .ZN(n12003) );
  XNOR2_X1 U14384 ( .A(n12002), .B(n12001), .ZN(n14821) );
  NOR2_X1 U14385 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14821), .ZN(n14820) );
  NOR2_X1 U14386 ( .A1(n12003), .A2(n14820), .ZN(n12004) );
  XOR2_X1 U14387 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n12004), .Z(n12010) );
  NOR2_X1 U14388 ( .A1(n12007), .A2(n14826), .ZN(n12008) );
  XNOR2_X1 U14389 ( .A(n12009), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U14390 ( .A1(n12010), .A2(n14805), .B1(n14784), .B2(n12013), .ZN(
        n12016) );
  INV_X1 U14391 ( .A(n12010), .ZN(n12011) );
  NAND2_X1 U14392 ( .A1(n14805), .A2(n12011), .ZN(n12012) );
  OAI211_X1 U14393 ( .C1(n12013), .C2(n14813), .A(n14827), .B(n12012), .ZN(
        n12014) );
  INV_X1 U14394 ( .A(n12014), .ZN(n12015) );
  MUX2_X1 U14395 ( .A(n12016), .B(n12015), .S(n12979), .Z(n12017) );
  NAND2_X1 U14396 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12663)
         );
  OAI211_X1 U14397 ( .C1(n11994), .C2(n14811), .A(n12017), .B(n12663), .ZN(
        P2_U3233) );
  AOI22_X1 U14398 ( .A1(n14333), .A2(n15046), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n14334), .ZN(n12019) );
  OAI21_X1 U14399 ( .B1(n12020), .B2(n14958), .A(n12019), .ZN(n12021) );
  AOI21_X1 U14400 ( .B1(n12022), .B2(n12520), .A(n12021), .ZN(n12023) );
  OAI21_X1 U14401 ( .B1(n12018), .B2(n14334), .A(n12023), .ZN(P3_U3204) );
  AOI21_X1 U14402 ( .B1(n12025), .B2(n12024), .A(n12168), .ZN(n12033) );
  NAND2_X1 U14403 ( .A1(n12174), .A2(n12026), .ZN(n12028) );
  NOR2_X1 U14404 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15221), .ZN(n12205) );
  AOI21_X1 U14405 ( .B1(n14916), .B2(n12482), .A(n12205), .ZN(n12027) );
  OAI211_X1 U14406 ( .C1(n12029), .C2(n12141), .A(n12028), .B(n12027), .ZN(
        n12030) );
  AOI21_X1 U14407 ( .B1(n12031), .B2(n14918), .A(n12030), .ZN(n12032) );
  OAI21_X1 U14408 ( .B1(n12033), .B2(n12153), .A(n12032), .ZN(P3_U3155) );
  INV_X1 U14409 ( .A(n12035), .ZN(n12103) );
  AOI21_X1 U14410 ( .B1(n12378), .B2(n12034), .A(n12103), .ZN(n12042) );
  INV_X1 U14411 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12036) );
  OAI22_X1 U14412 ( .A1(n12416), .A2(n12141), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12036), .ZN(n12037) );
  AOI21_X1 U14413 ( .B1(n12364), .B2(n14916), .A(n12037), .ZN(n12039) );
  NAND2_X1 U14414 ( .A1(n12174), .A2(n12396), .ZN(n12038) );
  OAI211_X1 U14415 ( .C1(n12542), .C2(n12177), .A(n12039), .B(n12038), .ZN(
        n12040) );
  INV_X1 U14416 ( .A(n12040), .ZN(n12041) );
  OAI21_X1 U14417 ( .B1(n12042), .B2(n12153), .A(n12041), .ZN(P3_U3156) );
  XNOR2_X1 U14418 ( .A(n12044), .B(n12043), .ZN(n12049) );
  NAND2_X1 U14419 ( .A1(n12466), .A2(n12170), .ZN(n12045) );
  NAND2_X1 U14420 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12316)
         );
  OAI211_X1 U14421 ( .C1(n12441), .C2(n12172), .A(n12045), .B(n12316), .ZN(
        n12047) );
  NOR2_X1 U14422 ( .A1(n12618), .A2(n12177), .ZN(n12046) );
  AOI211_X1 U14423 ( .C1(n12446), .C2(n12174), .A(n12047), .B(n12046), .ZN(
        n12048) );
  OAI21_X1 U14424 ( .B1(n12049), .B2(n12153), .A(n12048), .ZN(P3_U3159) );
  OAI21_X1 U14425 ( .B1(n12052), .B2(n6607), .A(n12051), .ZN(n12053) );
  NAND2_X1 U14426 ( .A1(n12053), .A2(n14914), .ZN(n12058) );
  NOR2_X1 U14427 ( .A1(n12441), .A2(n12141), .ZN(n12056) );
  OAI22_X1 U14428 ( .A1(n12416), .A2(n12172), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12054), .ZN(n12055) );
  AOI211_X1 U14429 ( .C1(n12419), .C2(n12174), .A(n12056), .B(n12055), .ZN(
        n12057) );
  OAI211_X1 U14430 ( .C1(n12610), .C2(n12177), .A(n12058), .B(n12057), .ZN(
        P3_U3163) );
  XNOR2_X1 U14431 ( .A(n12059), .B(n12060), .ZN(n12136) );
  OAI22_X1 U14432 ( .A1(n12136), .A2(n12184), .B1(n12060), .B2(n12059), .ZN(
        n12063) );
  XNOR2_X1 U14433 ( .A(n12061), .B(n12183), .ZN(n12062) );
  XNOR2_X1 U14434 ( .A(n12063), .B(n12062), .ZN(n12070) );
  NOR2_X1 U14435 ( .A1(n14348), .A2(n12177), .ZN(n12069) );
  INV_X1 U14436 ( .A(n14349), .ZN(n12067) );
  AOI21_X1 U14437 ( .B1(n14344), .B2(n14916), .A(n12064), .ZN(n12066) );
  NAND2_X1 U14438 ( .A1(n12184), .A2(n12170), .ZN(n12065) );
  OAI211_X1 U14439 ( .C1(n12161), .C2(n12067), .A(n12066), .B(n12065), .ZN(
        n12068) );
  AOI211_X1 U14440 ( .C1(n12070), .C2(n14914), .A(n12069), .B(n12068), .ZN(
        n12071) );
  INV_X1 U14441 ( .A(n12071), .ZN(P3_U3164) );
  INV_X1 U14442 ( .A(n12073), .ZN(n12104) );
  INV_X1 U14443 ( .A(n12074), .ZN(n12076) );
  NOR3_X1 U14444 ( .A1(n12104), .A2(n12076), .A3(n12075), .ZN(n12079) );
  INV_X1 U14445 ( .A(n12077), .ZN(n12078) );
  OAI21_X1 U14446 ( .B1(n12079), .B2(n12078), .A(n14914), .ZN(n12083) );
  AOI22_X1 U14447 ( .A1(n12364), .A2(n12170), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12080) );
  OAI21_X1 U14448 ( .B1(n12367), .B2(n12172), .A(n12080), .ZN(n12081) );
  AOI21_X1 U14449 ( .B1(n12370), .B2(n12174), .A(n12081), .ZN(n12082) );
  OAI211_X1 U14450 ( .C1(n12598), .C2(n12177), .A(n12083), .B(n12082), .ZN(
        P3_U3165) );
  INV_X1 U14451 ( .A(n12567), .ZN(n12491) );
  AOI21_X1 U14452 ( .B1(n12085), .B2(n12084), .A(n12153), .ZN(n12086) );
  NAND2_X1 U14453 ( .A1(n12086), .A2(n7502), .ZN(n12091) );
  NAND2_X1 U14454 ( .A1(n12170), .A2(n12482), .ZN(n12087) );
  NAND2_X1 U14455 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12257)
         );
  OAI211_X1 U14456 ( .C1(n12172), .C2(n12088), .A(n12087), .B(n12257), .ZN(
        n12089) );
  AOI21_X1 U14457 ( .B1(n12174), .B2(n12489), .A(n12089), .ZN(n12090) );
  OAI211_X1 U14458 ( .C1(n12491), .C2(n12177), .A(n12091), .B(n12090), .ZN(
        P3_U3166) );
  XNOR2_X1 U14459 ( .A(n12092), .B(n12093), .ZN(n12099) );
  NAND2_X1 U14460 ( .A1(n12467), .A2(n12170), .ZN(n12094) );
  NAND2_X1 U14461 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12274)
         );
  OAI211_X1 U14462 ( .C1(n12440), .C2(n12172), .A(n12094), .B(n12274), .ZN(
        n12097) );
  NOR2_X1 U14463 ( .A1(n12623), .A2(n12177), .ZN(n12096) );
  AOI211_X1 U14464 ( .C1(n12472), .C2(n12174), .A(n12097), .B(n12096), .ZN(
        n12098) );
  OAI21_X1 U14465 ( .B1(n12099), .B2(n12153), .A(n12098), .ZN(P3_U3168) );
  INV_X1 U14466 ( .A(n12100), .ZN(n12102) );
  NOR3_X1 U14467 ( .A1(n12103), .A2(n12102), .A3(n12101), .ZN(n12105) );
  OAI21_X1 U14468 ( .B1(n12105), .B2(n12104), .A(n14914), .ZN(n12109) );
  AOI22_X1 U14469 ( .A1(n12378), .A2(n12170), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12106) );
  OAI21_X1 U14470 ( .B1(n12352), .B2(n12172), .A(n12106), .ZN(n12107) );
  AOI21_X1 U14471 ( .B1(n12383), .B2(n12174), .A(n12107), .ZN(n12108) );
  OAI211_X1 U14472 ( .C1(n12602), .C2(n12177), .A(n12109), .B(n12108), .ZN(
        P3_U3169) );
  XNOR2_X1 U14473 ( .A(n12111), .B(n12110), .ZN(n12117) );
  AOI22_X1 U14474 ( .A1(n12181), .A2(n14916), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12113) );
  NAND2_X1 U14475 ( .A1(n12174), .A2(n12433), .ZN(n12112) );
  OAI211_X1 U14476 ( .C1(n12427), .C2(n12141), .A(n12113), .B(n12112), .ZN(
        n12114) );
  AOI21_X1 U14477 ( .B1(n12115), .B2(n14918), .A(n12114), .ZN(n12116) );
  OAI21_X1 U14478 ( .B1(n12117), .B2(n12153), .A(n12116), .ZN(P3_U3173) );
  XNOR2_X1 U14479 ( .A(n12119), .B(n14344), .ZN(n12120) );
  XNOR2_X1 U14480 ( .A(n12118), .B(n12120), .ZN(n12127) );
  NAND2_X1 U14481 ( .A1(n12174), .A2(n12517), .ZN(n12123) );
  AOI21_X1 U14482 ( .B1(n12497), .B2(n14916), .A(n12121), .ZN(n12122) );
  OAI211_X1 U14483 ( .C1(n12513), .C2(n12141), .A(n12123), .B(n12122), .ZN(
        n12124) );
  AOI21_X1 U14484 ( .B1(n12125), .B2(n14918), .A(n12124), .ZN(n12126) );
  OAI21_X1 U14485 ( .B1(n12127), .B2(n12153), .A(n12126), .ZN(P3_U3174) );
  INV_X1 U14486 ( .A(n12129), .ZN(n12130) );
  AOI21_X1 U14487 ( .B1(n12180), .B2(n12128), .A(n12130), .ZN(n12135) );
  AOI22_X1 U14488 ( .A1(n12378), .A2(n14916), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12132) );
  NAND2_X1 U14489 ( .A1(n12174), .A2(n12407), .ZN(n12131) );
  OAI211_X1 U14490 ( .C1(n12428), .C2(n12141), .A(n12132), .B(n12131), .ZN(
        n12133) );
  AOI21_X1 U14491 ( .B1(n12406), .B2(n14918), .A(n12133), .ZN(n12134) );
  OAI21_X1 U14492 ( .B1(n12135), .B2(n12153), .A(n12134), .ZN(P3_U3175) );
  XNOR2_X1 U14493 ( .A(n12136), .B(n14347), .ZN(n12146) );
  NOR2_X1 U14494 ( .A1(n12137), .A2(n12177), .ZN(n12143) );
  AOI21_X1 U14495 ( .B1(n14916), .B2(n12183), .A(n12138), .ZN(n12139) );
  OAI21_X1 U14496 ( .B1(n12141), .B2(n12140), .A(n12139), .ZN(n12142) );
  AOI211_X1 U14497 ( .C1(n12144), .C2(n12174), .A(n12143), .B(n12142), .ZN(
        n12145) );
  OAI21_X1 U14498 ( .B1(n12146), .B2(n12153), .A(n12145), .ZN(P3_U3176) );
  XNOR2_X1 U14499 ( .A(n12147), .B(n12148), .ZN(n12154) );
  NAND2_X1 U14500 ( .A1(n12170), .A2(n12481), .ZN(n12149) );
  NAND2_X1 U14501 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12294)
         );
  OAI211_X1 U14502 ( .C1(n12172), .C2(n12427), .A(n12149), .B(n12294), .ZN(
        n12151) );
  INV_X1 U14503 ( .A(n12559), .ZN(n12460) );
  NOR2_X1 U14504 ( .A1(n12460), .A2(n12177), .ZN(n12150) );
  AOI211_X1 U14505 ( .C1(n12458), .C2(n12174), .A(n12151), .B(n12150), .ZN(
        n12152) );
  OAI21_X1 U14506 ( .B1(n12154), .B2(n12153), .A(n12152), .ZN(P3_U3178) );
  OAI21_X1 U14507 ( .B1(n12158), .B2(n12156), .A(n12157), .ZN(n12159) );
  NAND2_X1 U14508 ( .A1(n12159), .A2(n14914), .ZN(n12165) );
  INV_X1 U14509 ( .A(n12356), .ZN(n12162) );
  AOI22_X1 U14510 ( .A1(n12379), .A2(n12170), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12160) );
  OAI21_X1 U14511 ( .B1(n12162), .B2(n12161), .A(n12160), .ZN(n12163) );
  AOI21_X1 U14512 ( .B1(n12179), .B2(n14916), .A(n12163), .ZN(n12164) );
  OAI211_X1 U14513 ( .C1(n12594), .C2(n12177), .A(n12165), .B(n12164), .ZN(
        P3_U3180) );
  NOR3_X1 U14514 ( .A1(n12168), .A2(n7350), .A3(n12167), .ZN(n12169) );
  OAI21_X1 U14515 ( .B1(n6614), .B2(n12169), .A(n14914), .ZN(n12176) );
  NAND2_X1 U14516 ( .A1(n12497), .A2(n12170), .ZN(n12171) );
  NAND2_X1 U14517 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12232)
         );
  OAI211_X1 U14518 ( .C1(n12500), .C2(n12172), .A(n12171), .B(n12232), .ZN(
        n12173) );
  AOI21_X1 U14519 ( .B1(n12503), .B2(n12174), .A(n12173), .ZN(n12175) );
  OAI211_X1 U14520 ( .C1(n12629), .C2(n12177), .A(n12176), .B(n12175), .ZN(
        P3_U3181) );
  MUX2_X1 U14521 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12178), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14522 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12341), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14523 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12179), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14524 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12340), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14525 ( .A(n12379), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12191), .Z(
        P3_U3516) );
  MUX2_X1 U14526 ( .A(n12364), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12191), .Z(
        P3_U3515) );
  MUX2_X1 U14527 ( .A(n12378), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12191), .Z(
        P3_U3514) );
  MUX2_X1 U14528 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12180), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14529 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12181), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14530 ( .A(n12182), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12191), .Z(
        P3_U3511) );
  MUX2_X1 U14531 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12452), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14532 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12466), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14533 ( .A(n12481), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12191), .Z(
        P3_U3508) );
  MUX2_X1 U14534 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12467), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14535 ( .A(n12482), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12191), .Z(
        P3_U3506) );
  MUX2_X1 U14536 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12497), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14537 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n14344), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14538 ( .A(n12183), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12191), .Z(
        P3_U3503) );
  MUX2_X1 U14539 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12184), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14540 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12185), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14541 ( .A(n12186), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12191), .Z(
        P3_U3500) );
  MUX2_X1 U14542 ( .A(n14968), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12191), .Z(
        P3_U3499) );
  MUX2_X1 U14543 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12187), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14544 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n14969), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14545 ( .A(n12188), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12191), .Z(
        P3_U3496) );
  MUX2_X1 U14546 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12189), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14547 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12190), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14548 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n15036), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14549 ( .A(n7333), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12191), .Z(
        P3_U3492) );
  MUX2_X1 U14550 ( .A(n15033), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12191), .Z(
        P3_U3491) );
  NAND2_X1 U14551 ( .A1(n12197), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12225) );
  OAI21_X1 U14552 ( .B1(n12197), .B2(P3_REG2_REG_14__SCAN_IN), .A(n12225), 
        .ZN(n12220) );
  NOR2_X1 U14553 ( .A1(n12210), .A2(n12192), .ZN(n12194) );
  XOR2_X1 U14554 ( .A(n12220), .B(n12221), .Z(n12219) );
  INV_X1 U14555 ( .A(n12197), .ZN(n12217) );
  NAND2_X1 U14556 ( .A1(n12195), .A2(n12210), .ZN(n12203) );
  INV_X1 U14557 ( .A(n12200), .ZN(n12196) );
  NAND2_X1 U14558 ( .A1(n12203), .A2(n12196), .ZN(n12199) );
  NAND2_X1 U14559 ( .A1(n12197), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12235) );
  OAI21_X1 U14560 ( .B1(n12197), .B2(P3_REG1_REG_14__SCAN_IN), .A(n12235), 
        .ZN(n12212) );
  MUX2_X1 U14561 ( .A(n12220), .B(n12212), .S(n12198), .Z(n12201) );
  NAND2_X1 U14562 ( .A1(n12199), .A2(n12201), .ZN(n12204) );
  NOR2_X1 U14563 ( .A1(n12201), .A2(n12200), .ZN(n12202) );
  NAND2_X1 U14564 ( .A1(n12203), .A2(n12202), .ZN(n12227) );
  NAND3_X1 U14565 ( .A1(n12204), .A2(n14922), .A3(n12227), .ZN(n12208) );
  NAND2_X1 U14566 ( .A1(n14921), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n12207) );
  INV_X1 U14567 ( .A(n12205), .ZN(n12206) );
  NAND3_X1 U14568 ( .A1(n12208), .A2(n12207), .A3(n12206), .ZN(n12216) );
  AOI21_X1 U14569 ( .B1(n12213), .B2(n12212), .A(n12234), .ZN(n12214) );
  NOR2_X1 U14570 ( .A1(n12214), .A2(n14937), .ZN(n12215) );
  AOI211_X1 U14571 ( .C1(n14948), .C2(n12217), .A(n12216), .B(n12215), .ZN(
        n12218) );
  OAI21_X1 U14572 ( .B1(n14940), .B2(n12219), .A(n12218), .ZN(P3_U3196) );
  INV_X1 U14573 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12224) );
  NAND2_X1 U14574 ( .A1(n12225), .A2(n12222), .ZN(n12245) );
  AOI21_X1 U14575 ( .B1(n12224), .B2(n12223), .A(n12246), .ZN(n12242) );
  INV_X1 U14576 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12575) );
  MUX2_X1 U14577 ( .A(n12224), .B(n12575), .S(n12198), .Z(n12230) );
  MUX2_X1 U14578 ( .A(n12225), .B(n12235), .S(n12198), .Z(n12226) );
  NAND2_X1 U14579 ( .A1(n12227), .A2(n12226), .ZN(n12228) );
  NOR2_X1 U14580 ( .A1(n12228), .A2(n12260), .ZN(n12251) );
  AOI21_X1 U14581 ( .B1(n12260), .B2(n12228), .A(n12251), .ZN(n12229) );
  OAI21_X1 U14582 ( .B1(n12230), .B2(n12229), .A(n6878), .ZN(n12240) );
  INV_X1 U14583 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14211) );
  INV_X1 U14584 ( .A(n12260), .ZN(n12231) );
  NAND2_X1 U14585 ( .A1(n14948), .A2(n12231), .ZN(n12233) );
  OAI211_X1 U14586 ( .C1(n14211), .C2(n14951), .A(n12233), .B(n12232), .ZN(
        n12239) );
  XNOR2_X1 U14587 ( .A(n12260), .B(n12259), .ZN(n12236) );
  AOI21_X1 U14588 ( .B1(n12575), .B2(n12236), .A(n12261), .ZN(n12237) );
  NOR2_X1 U14589 ( .A1(n12237), .A2(n14937), .ZN(n12238) );
  AOI211_X1 U14590 ( .C1(n14922), .C2(n12240), .A(n12239), .B(n12238), .ZN(
        n12241) );
  OAI21_X1 U14591 ( .B1(n12242), .B2(n14940), .A(n12241), .ZN(P3_U3197) );
  INV_X1 U14592 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12252) );
  OR2_X1 U14593 ( .A1(n12280), .A2(n12252), .ZN(n12244) );
  NAND2_X1 U14594 ( .A1(n12280), .A2(n12252), .ZN(n12243) );
  AND2_X1 U14595 ( .A1(n12244), .A2(n12243), .ZN(n12250) );
  AND2_X1 U14596 ( .A1(n12260), .A2(n12245), .ZN(n12247) );
  INV_X1 U14597 ( .A(n12282), .ZN(n12248) );
  AOI21_X1 U14598 ( .B1(n12250), .B2(n12249), .A(n12248), .ZN(n12270) );
  INV_X1 U14599 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12571) );
  MUX2_X1 U14600 ( .A(n12252), .B(n12571), .S(n12198), .Z(n12253) );
  INV_X1 U14601 ( .A(n12280), .ZN(n12256) );
  NAND2_X1 U14602 ( .A1(n12253), .A2(n12256), .ZN(n12275) );
  MUX2_X1 U14603 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n12198), .Z(n12254) );
  NAND2_X1 U14604 ( .A1(n12275), .A2(n6618), .ZN(n12255) );
  XNOR2_X1 U14605 ( .A(n6602), .B(n12255), .ZN(n12268) );
  INV_X1 U14606 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14281) );
  NAND2_X1 U14607 ( .A1(n14948), .A2(n12256), .ZN(n12258) );
  OAI211_X1 U14608 ( .C1(n14281), .C2(n14951), .A(n12258), .B(n12257), .ZN(
        n12267) );
  AND2_X1 U14609 ( .A1(n12260), .A2(n12259), .ZN(n12262) );
  NAND2_X1 U14610 ( .A1(n12280), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n12271) );
  OAI21_X1 U14611 ( .B1(n12280), .B2(P3_REG1_REG_16__SCAN_IN), .A(n12271), 
        .ZN(n12263) );
  NAND2_X1 U14612 ( .A1(n12264), .A2(n12263), .ZN(n12265) );
  AOI21_X1 U14613 ( .B1(n12272), .B2(n12265), .A(n14937), .ZN(n12266) );
  AOI211_X1 U14614 ( .C1(n14922), .C2(n12268), .A(n12267), .B(n12266), .ZN(
        n12269) );
  OAI21_X1 U14615 ( .B1(n12270), .B2(n14940), .A(n12269), .ZN(P3_U3198) );
  INV_X1 U14616 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12565) );
  AOI21_X1 U14617 ( .B1(n12565), .B2(n12273), .A(n12289), .ZN(n12288) );
  INV_X1 U14618 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15260) );
  OAI21_X1 U14619 ( .B1(n14951), .B2(n15260), .A(n12274), .ZN(n12279) );
  MUX2_X1 U14620 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12198), .Z(n12297) );
  XNOR2_X1 U14621 ( .A(n12297), .B(n12296), .ZN(n12276) );
  AOI211_X1 U14622 ( .C1(n12277), .C2(n12276), .A(n12295), .B(n14943), .ZN(
        n12278) );
  AOI211_X1 U14623 ( .C1(n14948), .C2(n12303), .A(n12279), .B(n12278), .ZN(
        n12287) );
  NAND2_X1 U14624 ( .A1(n12280), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12281) );
  INV_X1 U14625 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12284) );
  AND2_X1 U14626 ( .A1(n12283), .A2(n12284), .ZN(n12285) );
  OAI21_X1 U14627 ( .B1(n12285), .B2(n12304), .A(n14923), .ZN(n12286) );
  OAI211_X1 U14628 ( .C1(n12288), .C2(n14937), .A(n12287), .B(n12286), .ZN(
        P3_U3199) );
  NOR2_X1 U14629 ( .A1(n12290), .A2(n12289), .ZN(n12293) );
  NAND2_X1 U14630 ( .A1(n12306), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n12314) );
  OAI21_X1 U14631 ( .B1(n12306), .B2(P3_REG1_REG_18__SCAN_IN), .A(n12314), 
        .ZN(n12292) );
  INV_X1 U14632 ( .A(n12315), .ZN(n12291) );
  AOI21_X1 U14633 ( .B1(n12293), .B2(n12292), .A(n12291), .ZN(n12313) );
  INV_X1 U14634 ( .A(n12306), .ZN(n12318) );
  INV_X1 U14635 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n14325) );
  OAI21_X1 U14636 ( .B1(n14951), .B2(n14325), .A(n12294), .ZN(n12302) );
  MUX2_X1 U14637 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12198), .Z(n12299) );
  AOI21_X1 U14638 ( .B1(n12297), .B2(n12296), .A(n12295), .ZN(n12319) );
  XOR2_X1 U14639 ( .A(n12306), .B(n12319), .Z(n12298) );
  NOR2_X1 U14640 ( .A1(n12298), .A2(n12299), .ZN(n12317) );
  AOI21_X1 U14641 ( .B1(n12299), .B2(n12298), .A(n12317), .ZN(n12300) );
  NOR2_X1 U14642 ( .A1(n12300), .A2(n14943), .ZN(n12301) );
  AOI211_X1 U14643 ( .C1(n14948), .C2(n12318), .A(n12302), .B(n12301), .ZN(
        n12312) );
  NOR2_X1 U14644 ( .A1(n12303), .A2(n6536), .ZN(n12305) );
  NAND2_X1 U14645 ( .A1(n12306), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12325) );
  OAI21_X1 U14646 ( .B1(n12306), .B2(P3_REG2_REG_18__SCAN_IN), .A(n12325), 
        .ZN(n12307) );
  INV_X1 U14647 ( .A(n12326), .ZN(n12310) );
  AND2_X1 U14648 ( .A1(n12308), .A2(n12307), .ZN(n12309) );
  OAI21_X1 U14649 ( .B1(n12310), .B2(n12309), .A(n14923), .ZN(n12311) );
  OAI211_X1 U14650 ( .C1(n12313), .C2(n14937), .A(n12312), .B(n12311), .ZN(
        P3_U3200) );
  XNOR2_X1 U14651 ( .A(n9767), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12321) );
  OAI21_X1 U14652 ( .B1(n14951), .B2(n6894), .A(n12316), .ZN(n12324) );
  AOI21_X1 U14653 ( .B1(n12319), .B2(n12318), .A(n12317), .ZN(n12323) );
  INV_X1 U14654 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12320) );
  MUX2_X1 U14655 ( .A(n12320), .B(P3_REG2_REG_19__SCAN_IN), .S(n9767), .Z(
        n12327) );
  MUX2_X1 U14656 ( .A(n12327), .B(n12321), .S(n12198), .Z(n12322) );
  NAND2_X1 U14657 ( .A1(n12326), .A2(n12325), .ZN(n12328) );
  XNOR2_X1 U14658 ( .A(n12328), .B(n12327), .ZN(n12329) );
  NAND2_X1 U14659 ( .A1(n12329), .A2(n14923), .ZN(n12330) );
  NAND2_X1 U14660 ( .A1(n12331), .A2(n12520), .ZN(n12334) );
  AOI22_X1 U14661 ( .A1(n12332), .A2(n15046), .B1(n14334), .B2(
        P3_REG2_REG_28__SCAN_IN), .ZN(n12333) );
  OAI211_X1 U14662 ( .C1(n12589), .C2(n14958), .A(n12334), .B(n12333), .ZN(
        n12335) );
  AOI21_X1 U14663 ( .B1(n12336), .B2(n15050), .A(n12335), .ZN(n12337) );
  INV_X1 U14664 ( .A(n12337), .ZN(P3_U3205) );
  OAI21_X1 U14665 ( .B1(n6583), .B2(n12339), .A(n12338), .ZN(n12342) );
  AOI222_X1 U14666 ( .A1(n15039), .A2(n12342), .B1(n12341), .B2(n15035), .C1(
        n12340), .C2(n15034), .ZN(n12526) );
  OAI21_X1 U14667 ( .B1(n12344), .B2(n6567), .A(n12343), .ZN(n12524) );
  AOI22_X1 U14668 ( .A1(n12345), .A2(n15046), .B1(n14334), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12346) );
  OAI21_X1 U14669 ( .B1(n12347), .B2(n14958), .A(n12346), .ZN(n12348) );
  AOI21_X1 U14670 ( .B1(n12524), .B2(n12520), .A(n12348), .ZN(n12349) );
  OAI21_X1 U14671 ( .B1(n12526), .B2(n14334), .A(n12349), .ZN(P3_U3206) );
  XOR2_X1 U14672 ( .A(n12350), .B(n12355), .Z(n12351) );
  OAI222_X1 U14673 ( .A1(n15017), .A2(n12353), .B1(n15019), .B2(n12352), .C1(
        n12351), .C2(n12512), .ZN(n12527) );
  INV_X1 U14674 ( .A(n12527), .ZN(n12360) );
  XNOR2_X1 U14675 ( .A(n12355), .B(n12354), .ZN(n12528) );
  AOI22_X1 U14676 ( .A1(n12356), .A2(n15046), .B1(n14334), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12357) );
  OAI21_X1 U14677 ( .B1(n12594), .B2(n14958), .A(n12357), .ZN(n12358) );
  AOI21_X1 U14678 ( .B1(n12528), .B2(n12520), .A(n12358), .ZN(n12359) );
  OAI21_X1 U14679 ( .B1(n12360), .B2(n14334), .A(n12359), .ZN(P3_U3207) );
  OAI211_X1 U14680 ( .C1(n12363), .C2(n12362), .A(n12361), .B(n15039), .ZN(
        n12366) );
  NAND2_X1 U14681 ( .A1(n12364), .A2(n15034), .ZN(n12365) );
  OAI211_X1 U14682 ( .C1(n12367), .C2(n15017), .A(n12366), .B(n12365), .ZN(
        n12531) );
  INV_X1 U14683 ( .A(n12531), .ZN(n12374) );
  XNOR2_X1 U14684 ( .A(n12369), .B(n12368), .ZN(n12532) );
  AOI22_X1 U14685 ( .A1(n12370), .A2(n15046), .B1(n14334), .B2(
        P3_REG2_REG_25__SCAN_IN), .ZN(n12371) );
  OAI21_X1 U14686 ( .B1(n12598), .B2(n14958), .A(n12371), .ZN(n12372) );
  AOI21_X1 U14687 ( .B1(n12532), .B2(n12520), .A(n12372), .ZN(n12373) );
  OAI21_X1 U14688 ( .B1(n12374), .B2(n14334), .A(n12373), .ZN(P3_U3208) );
  OAI211_X1 U14689 ( .C1(n12377), .C2(n12376), .A(n12375), .B(n15039), .ZN(
        n12381) );
  AOI22_X1 U14690 ( .A1(n12379), .A2(n15035), .B1(n15034), .B2(n12378), .ZN(
        n12380) );
  NAND2_X1 U14691 ( .A1(n12381), .A2(n12380), .ZN(n12535) );
  INV_X1 U14692 ( .A(n12535), .ZN(n12387) );
  OAI21_X1 U14693 ( .B1(n6578), .B2(n9140), .A(n12382), .ZN(n12536) );
  AOI22_X1 U14694 ( .A1(n12383), .A2(n15046), .B1(n14334), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n12384) );
  OAI21_X1 U14695 ( .B1(n12602), .B2(n14958), .A(n12384), .ZN(n12385) );
  AOI21_X1 U14696 ( .B1(n12536), .B2(n12520), .A(n12385), .ZN(n12386) );
  OAI21_X1 U14697 ( .B1(n12387), .B2(n14334), .A(n12386), .ZN(P3_U3209) );
  AOI21_X1 U14698 ( .B1(n12388), .B2(n12393), .A(n12512), .ZN(n12392) );
  OAI22_X1 U14699 ( .A1(n12389), .A2(n15017), .B1(n12416), .B2(n15019), .ZN(
        n12390) );
  AOI21_X1 U14700 ( .B1(n12392), .B2(n12391), .A(n12390), .ZN(n12541) );
  OR2_X1 U14701 ( .A1(n12394), .A2(n12393), .ZN(n12539) );
  NAND3_X1 U14702 ( .A1(n12539), .A2(n12395), .A3(n12520), .ZN(n12398) );
  AOI22_X1 U14703 ( .A1(n12396), .A2(n15046), .B1(n14334), .B2(
        P3_REG2_REG_23__SCAN_IN), .ZN(n12397) );
  OAI211_X1 U14704 ( .C1(n12542), .C2(n14958), .A(n12398), .B(n12397), .ZN(
        n12399) );
  INV_X1 U14705 ( .A(n12399), .ZN(n12400) );
  OAI21_X1 U14706 ( .B1(n12541), .B2(n14334), .A(n12400), .ZN(P3_U3210) );
  XNOR2_X1 U14707 ( .A(n12402), .B(n12401), .ZN(n12403) );
  OAI222_X1 U14708 ( .A1(n15017), .A2(n9824), .B1(n15019), .B2(n12428), .C1(
        n12512), .C2(n12403), .ZN(n12543) );
  INV_X1 U14709 ( .A(n12543), .ZN(n12411) );
  XNOR2_X1 U14710 ( .A(n12405), .B(n12404), .ZN(n12544) );
  INV_X1 U14711 ( .A(n12406), .ZN(n12606) );
  AOI22_X1 U14712 ( .A1(n12407), .A2(n15046), .B1(n14334), .B2(
        P3_REG2_REG_22__SCAN_IN), .ZN(n12408) );
  OAI21_X1 U14713 ( .B1(n12606), .B2(n14958), .A(n12408), .ZN(n12409) );
  AOI21_X1 U14714 ( .B1(n12544), .B2(n12520), .A(n12409), .ZN(n12410) );
  OAI21_X1 U14715 ( .B1(n12411), .B2(n14334), .A(n12410), .ZN(P3_U3211) );
  INV_X1 U14716 ( .A(n12412), .ZN(n12413) );
  AOI21_X1 U14717 ( .B1(n12417), .B2(n12414), .A(n12413), .ZN(n12415) );
  OAI222_X1 U14718 ( .A1(n15017), .A2(n12416), .B1(n15019), .B2(n12441), .C1(
        n12512), .C2(n12415), .ZN(n12547) );
  INV_X1 U14719 ( .A(n12547), .ZN(n12423) );
  XOR2_X1 U14720 ( .A(n12418), .B(n12417), .Z(n12548) );
  AOI22_X1 U14721 ( .A1(P3_REG2_REG_21__SCAN_IN), .A2(n14334), .B1(n12419), 
        .B2(n15046), .ZN(n12420) );
  OAI21_X1 U14722 ( .B1(n12610), .B2(n14958), .A(n12420), .ZN(n12421) );
  AOI21_X1 U14723 ( .B1(n12548), .B2(n12520), .A(n12421), .ZN(n12422) );
  OAI21_X1 U14724 ( .B1(n12423), .B2(n14334), .A(n12422), .ZN(P3_U3212) );
  XNOR2_X1 U14725 ( .A(n12425), .B(n12429), .ZN(n12426) );
  OAI222_X1 U14726 ( .A1(n15017), .A2(n12428), .B1(n15019), .B2(n12427), .C1(
        n12512), .C2(n12426), .ZN(n12551) );
  NAND2_X1 U14727 ( .A1(n12430), .A2(n12429), .ZN(n12431) );
  AND2_X1 U14728 ( .A1(n12432), .A2(n12431), .ZN(n12552) );
  NAND2_X1 U14729 ( .A1(n12552), .A2(n12520), .ZN(n12435) );
  AOI22_X1 U14730 ( .A1(n14334), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n15046), 
        .B2(n12433), .ZN(n12434) );
  OAI211_X1 U14731 ( .C1(n12614), .C2(n14958), .A(n12435), .B(n12434), .ZN(
        n12436) );
  AOI21_X1 U14732 ( .B1(n12551), .B2(n15050), .A(n12436), .ZN(n12437) );
  INV_X1 U14733 ( .A(n12437), .ZN(P3_U3213) );
  XNOR2_X1 U14734 ( .A(n12438), .B(n12444), .ZN(n12439) );
  OAI222_X1 U14735 ( .A1(n15017), .A2(n12441), .B1(n15019), .B2(n12440), .C1(
        n12512), .C2(n12439), .ZN(n12555) );
  INV_X1 U14736 ( .A(n12555), .ZN(n12450) );
  AND2_X1 U14737 ( .A1(n12454), .A2(n12442), .ZN(n12445) );
  OAI21_X1 U14738 ( .B1(n12445), .B2(n12444), .A(n12443), .ZN(n12556) );
  AOI22_X1 U14739 ( .A1(n14334), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n15046), 
        .B2(n12446), .ZN(n12447) );
  OAI21_X1 U14740 ( .B1(n12618), .B2(n14958), .A(n12447), .ZN(n12448) );
  AOI21_X1 U14741 ( .B1(n12556), .B2(n12520), .A(n12448), .ZN(n12449) );
  OAI21_X1 U14742 ( .B1(n12450), .B2(n14334), .A(n12449), .ZN(P3_U3214) );
  OAI21_X1 U14743 ( .B1(n6605), .B2(n12457), .A(n12451), .ZN(n12453) );
  AOI222_X1 U14744 ( .A1(n15039), .A2(n12453), .B1(n12452), .B2(n15035), .C1(
        n12481), .C2(n15034), .ZN(n12562) );
  INV_X1 U14745 ( .A(n12454), .ZN(n12455) );
  AOI21_X1 U14746 ( .B1(n12457), .B2(n12456), .A(n12455), .ZN(n12560) );
  AOI22_X1 U14747 ( .A1(n14334), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15046), 
        .B2(n12458), .ZN(n12459) );
  OAI21_X1 U14748 ( .B1(n12460), .B2(n14958), .A(n12459), .ZN(n12461) );
  AOI21_X1 U14749 ( .B1(n12560), .B2(n12520), .A(n12461), .ZN(n12462) );
  OAI21_X1 U14750 ( .B1(n12562), .B2(n14334), .A(n12462), .ZN(P3_U3215) );
  OAI211_X1 U14751 ( .C1(n12465), .C2(n12464), .A(n12463), .B(n15039), .ZN(
        n12469) );
  AOI22_X1 U14752 ( .A1(n15034), .A2(n12467), .B1(n12466), .B2(n15035), .ZN(
        n12468) );
  NAND2_X1 U14753 ( .A1(n12469), .A2(n12468), .ZN(n12563) );
  INV_X1 U14754 ( .A(n12563), .ZN(n12476) );
  XNOR2_X1 U14755 ( .A(n12471), .B(n12470), .ZN(n12564) );
  AOI22_X1 U14756 ( .A1(n14334), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15046), 
        .B2(n12472), .ZN(n12473) );
  OAI21_X1 U14757 ( .B1(n12623), .B2(n14958), .A(n12473), .ZN(n12474) );
  AOI21_X1 U14758 ( .B1(n12564), .B2(n12520), .A(n12474), .ZN(n12475) );
  OAI21_X1 U14759 ( .B1(n12476), .B2(n14334), .A(n12475), .ZN(P3_U3216) );
  NAND2_X1 U14760 ( .A1(n12477), .A2(n12485), .ZN(n12478) );
  NAND2_X1 U14761 ( .A1(n12479), .A2(n12478), .ZN(n12480) );
  NAND2_X1 U14762 ( .A1(n12480), .A2(n15039), .ZN(n12484) );
  AOI22_X1 U14763 ( .A1(n15034), .A2(n12482), .B1(n12481), .B2(n15035), .ZN(
        n12483) );
  OR2_X1 U14764 ( .A1(n12486), .A2(n12485), .ZN(n12487) );
  NAND2_X1 U14765 ( .A1(n12488), .A2(n12487), .ZN(n12568) );
  AOI22_X1 U14766 ( .A1(n14334), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15046), 
        .B2(n12489), .ZN(n12490) );
  OAI21_X1 U14767 ( .B1(n12491), .B2(n14958), .A(n12490), .ZN(n12492) );
  AOI21_X1 U14768 ( .B1(n12568), .B2(n12520), .A(n12492), .ZN(n12493) );
  OAI21_X1 U14769 ( .B1(n12570), .B2(n14334), .A(n12493), .ZN(P3_U3217) );
  OAI211_X1 U14770 ( .C1(n12496), .C2(n12495), .A(n6749), .B(n15039), .ZN(
        n12499) );
  NAND2_X1 U14771 ( .A1(n12497), .A2(n15034), .ZN(n12498) );
  OAI211_X1 U14772 ( .C1(n12500), .C2(n15017), .A(n12499), .B(n12498), .ZN(
        n12573) );
  INV_X1 U14773 ( .A(n12573), .ZN(n12507) );
  XNOR2_X1 U14774 ( .A(n12502), .B(n12501), .ZN(n12574) );
  AOI22_X1 U14775 ( .A1(n14334), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15046), 
        .B2(n12503), .ZN(n12504) );
  OAI21_X1 U14776 ( .B1(n12629), .B2(n14958), .A(n12504), .ZN(n12505) );
  AOI21_X1 U14777 ( .B1(n12574), .B2(n12520), .A(n12505), .ZN(n12506) );
  OAI21_X1 U14778 ( .B1(n12507), .B2(n14334), .A(n12506), .ZN(P3_U3218) );
  INV_X1 U14779 ( .A(n12508), .ZN(n12509) );
  AOI21_X1 U14780 ( .B1(n12515), .B2(n12510), .A(n12509), .ZN(n12511) );
  OAI222_X1 U14781 ( .A1(n15017), .A2(n12514), .B1(n15019), .B2(n12513), .C1(
        n12512), .C2(n12511), .ZN(n12581) );
  INV_X1 U14782 ( .A(n12581), .ZN(n12522) );
  XNOR2_X1 U14783 ( .A(n12516), .B(n12515), .ZN(n12582) );
  AOI22_X1 U14784 ( .A1(n14334), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n15046), 
        .B2(n12517), .ZN(n12518) );
  OAI21_X1 U14785 ( .B1(n12637), .B2(n14958), .A(n12518), .ZN(n12519) );
  AOI21_X1 U14786 ( .B1(n12582), .B2(n12520), .A(n12519), .ZN(n12521) );
  OAI21_X1 U14787 ( .B1(n12522), .B2(n14334), .A(n12521), .ZN(P3_U3220) );
  AOI22_X1 U14788 ( .A1(n12524), .A2(n14362), .B1(n15023), .B2(n12523), .ZN(
        n12525) );
  NAND2_X1 U14789 ( .A1(n12526), .A2(n12525), .ZN(n12590) );
  MUX2_X1 U14790 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12590), .S(n15096), .Z(
        P3_U3486) );
  INV_X1 U14791 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12529) );
  AOI21_X1 U14792 ( .B1(n12528), .B2(n14362), .A(n12527), .ZN(n12591) );
  MUX2_X1 U14793 ( .A(n12529), .B(n12591), .S(n15096), .Z(n12530) );
  OAI21_X1 U14794 ( .B1(n12594), .B2(n12585), .A(n12530), .ZN(P3_U3485) );
  INV_X1 U14795 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12533) );
  AOI21_X1 U14796 ( .B1(n14362), .B2(n12532), .A(n12531), .ZN(n12595) );
  MUX2_X1 U14797 ( .A(n12533), .B(n12595), .S(n15096), .Z(n12534) );
  OAI21_X1 U14798 ( .B1(n12598), .B2(n12585), .A(n12534), .ZN(P3_U3484) );
  INV_X1 U14799 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12537) );
  AOI21_X1 U14800 ( .B1(n14362), .B2(n12536), .A(n12535), .ZN(n12599) );
  MUX2_X1 U14801 ( .A(n12537), .B(n12599), .S(n15096), .Z(n12538) );
  OAI21_X1 U14802 ( .B1(n12602), .B2(n12585), .A(n12538), .ZN(P3_U3483) );
  NAND3_X1 U14803 ( .A1(n12539), .A2(n12395), .A3(n14362), .ZN(n12540) );
  OAI211_X1 U14804 ( .C1(n12542), .C2(n15030), .A(n12541), .B(n12540), .ZN(
        n12603) );
  MUX2_X1 U14805 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n12603), .S(n15096), .Z(
        P3_U3482) );
  INV_X1 U14806 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12545) );
  AOI21_X1 U14807 ( .B1(n14362), .B2(n12544), .A(n12543), .ZN(n12604) );
  MUX2_X1 U14808 ( .A(n12545), .B(n12604), .S(n15096), .Z(n12546) );
  OAI21_X1 U14809 ( .B1(n12606), .B2(n12585), .A(n12546), .ZN(P3_U3481) );
  INV_X1 U14810 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12549) );
  AOI21_X1 U14811 ( .B1(n14362), .B2(n12548), .A(n12547), .ZN(n12607) );
  MUX2_X1 U14812 ( .A(n12549), .B(n12607), .S(n15096), .Z(n12550) );
  OAI21_X1 U14813 ( .B1(n12610), .B2(n12585), .A(n12550), .ZN(P3_U3480) );
  INV_X1 U14814 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12553) );
  AOI21_X1 U14815 ( .B1(n12552), .B2(n14362), .A(n12551), .ZN(n12611) );
  MUX2_X1 U14816 ( .A(n12553), .B(n12611), .S(n15096), .Z(n12554) );
  OAI21_X1 U14817 ( .B1(n12614), .B2(n12585), .A(n12554), .ZN(P3_U3479) );
  INV_X1 U14818 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12557) );
  AOI21_X1 U14819 ( .B1(n14362), .B2(n12556), .A(n12555), .ZN(n12615) );
  MUX2_X1 U14820 ( .A(n12557), .B(n12615), .S(n15096), .Z(n12558) );
  OAI21_X1 U14821 ( .B1(n12585), .B2(n12618), .A(n12558), .ZN(P3_U3478) );
  AOI22_X1 U14822 ( .A1(n12560), .A2(n14362), .B1(n15023), .B2(n12559), .ZN(
        n12561) );
  NAND2_X1 U14823 ( .A1(n12562), .A2(n12561), .ZN(n12619) );
  MUX2_X1 U14824 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12619), .S(n15096), .Z(
        P3_U3477) );
  AOI21_X1 U14825 ( .B1(n14362), .B2(n12564), .A(n12563), .ZN(n12620) );
  MUX2_X1 U14826 ( .A(n12565), .B(n12620), .S(n15096), .Z(n12566) );
  OAI21_X1 U14827 ( .B1(n12623), .B2(n12585), .A(n12566), .ZN(P3_U3476) );
  AOI22_X1 U14828 ( .A1(n12568), .A2(n14362), .B1(n15023), .B2(n12567), .ZN(
        n12569) );
  AND2_X1 U14829 ( .A1(n12570), .A2(n12569), .ZN(n12624) );
  MUX2_X1 U14830 ( .A(n12571), .B(n12624), .S(n15096), .Z(n12572) );
  INV_X1 U14831 ( .A(n12572), .ZN(P3_U3475) );
  AOI21_X1 U14832 ( .B1(n14362), .B2(n12574), .A(n12573), .ZN(n12626) );
  MUX2_X1 U14833 ( .A(n12575), .B(n12626), .S(n15096), .Z(n12576) );
  OAI21_X1 U14834 ( .B1(n12629), .B2(n12585), .A(n12576), .ZN(P3_U3474) );
  INV_X1 U14835 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12579) );
  AOI21_X1 U14836 ( .B1(n14362), .B2(n12578), .A(n12577), .ZN(n12630) );
  MUX2_X1 U14837 ( .A(n12579), .B(n12630), .S(n15096), .Z(n12580) );
  OAI21_X1 U14838 ( .B1(n12633), .B2(n12585), .A(n12580), .ZN(P3_U3473) );
  AOI21_X1 U14839 ( .B1(n12582), .B2(n14362), .A(n12581), .ZN(n12634) );
  MUX2_X1 U14840 ( .A(n12583), .B(n12634), .S(n15096), .Z(n12584) );
  OAI21_X1 U14841 ( .B1(n12585), .B2(n12637), .A(n12584), .ZN(P3_U3472) );
  MUX2_X1 U14842 ( .A(n12587), .B(n12586), .S(n15081), .Z(n12588) );
  OAI21_X1 U14843 ( .B1(n12589), .B2(n12638), .A(n12588), .ZN(P3_U3455) );
  MUX2_X1 U14844 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12590), .S(n15081), .Z(
        P3_U3454) );
  MUX2_X1 U14845 ( .A(n12592), .B(n12591), .S(n15081), .Z(n12593) );
  OAI21_X1 U14846 ( .B1(n12594), .B2(n12638), .A(n12593), .ZN(P3_U3453) );
  MUX2_X1 U14847 ( .A(n12596), .B(n12595), .S(n15081), .Z(n12597) );
  OAI21_X1 U14848 ( .B1(n12598), .B2(n12638), .A(n12597), .ZN(P3_U3452) );
  MUX2_X1 U14849 ( .A(n12600), .B(n12599), .S(n15081), .Z(n12601) );
  OAI21_X1 U14850 ( .B1(n12602), .B2(n12638), .A(n12601), .ZN(P3_U3451) );
  MUX2_X1 U14851 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n12603), .S(n15081), .Z(
        P3_U3450) );
  MUX2_X1 U14852 ( .A(n15236), .B(n12604), .S(n15081), .Z(n12605) );
  OAI21_X1 U14853 ( .B1(n12606), .B2(n12638), .A(n12605), .ZN(P3_U3449) );
  MUX2_X1 U14854 ( .A(n12608), .B(n12607), .S(n15081), .Z(n12609) );
  OAI21_X1 U14855 ( .B1(n12610), .B2(n12638), .A(n12609), .ZN(P3_U3448) );
  MUX2_X1 U14856 ( .A(n12612), .B(n12611), .S(n15081), .Z(n12613) );
  OAI21_X1 U14857 ( .B1(n12614), .B2(n12638), .A(n12613), .ZN(P3_U3447) );
  MUX2_X1 U14858 ( .A(n12616), .B(n12615), .S(n15081), .Z(n12617) );
  OAI21_X1 U14859 ( .B1(n12638), .B2(n12618), .A(n12617), .ZN(P3_U3446) );
  MUX2_X1 U14860 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n12619), .S(n15081), .Z(
        P3_U3444) );
  MUX2_X1 U14861 ( .A(n12621), .B(n12620), .S(n15081), .Z(n12622) );
  OAI21_X1 U14862 ( .B1(n12623), .B2(n12638), .A(n12622), .ZN(P3_U3441) );
  MUX2_X1 U14863 ( .A(n15131), .B(n12624), .S(n15081), .Z(n12625) );
  INV_X1 U14864 ( .A(n12625), .ZN(P3_U3438) );
  MUX2_X1 U14865 ( .A(n12627), .B(n12626), .S(n15081), .Z(n12628) );
  OAI21_X1 U14866 ( .B1(n12629), .B2(n12638), .A(n12628), .ZN(P3_U3435) );
  MUX2_X1 U14867 ( .A(n12631), .B(n12630), .S(n15081), .Z(n12632) );
  OAI21_X1 U14868 ( .B1(n12633), .B2(n12638), .A(n12632), .ZN(P3_U3432) );
  MUX2_X1 U14869 ( .A(n12635), .B(n12634), .S(n15081), .Z(n12636) );
  OAI21_X1 U14870 ( .B1(n12638), .B2(n12637), .A(n12636), .ZN(P3_U3429) );
  MUX2_X1 U14871 ( .A(P3_D_REG_1__SCAN_IN), .B(n12639), .S(n12640), .Z(
        P3_U3377) );
  MUX2_X1 U14872 ( .A(P3_D_REG_0__SCAN_IN), .B(n7335), .S(n12640), .Z(P3_U3376) );
  INV_X1 U14873 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12641) );
  NAND3_X1 U14874 ( .A1(n12641), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n12643) );
  OAI22_X1 U14875 ( .A1(n12644), .A2(n12643), .B1(n12642), .B2(n11881), .ZN(
        n12645) );
  AOI21_X1 U14876 ( .B1(n12647), .B2(n12646), .A(n12645), .ZN(n12648) );
  INV_X1 U14877 ( .A(n12648), .ZN(P3_U3264) );
  OAI22_X1 U14878 ( .A1(n12957), .A2(n12773), .B1(n12654), .B2(n12771), .ZN(
        n13118) );
  OAI22_X1 U14879 ( .A1(n13126), .A2(n14384), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12655), .ZN(n12656) );
  AOI21_X1 U14880 ( .B1(n13118), .B2(n14378), .A(n12656), .ZN(n12657) );
  OAI211_X1 U14881 ( .C1(n13402), .C2(n12776), .A(n12658), .B(n12657), .ZN(
        P2_U3186) );
  INV_X1 U14882 ( .A(n12659), .ZN(n12758) );
  NOR3_X1 U14883 ( .A1(n12660), .A2(n12714), .A3(n12765), .ZN(n12661) );
  AOI21_X1 U14884 ( .B1(n12758), .B2(n14376), .A(n12661), .ZN(n12670) );
  NOR2_X1 U14885 ( .A1(n14384), .A2(n13252), .ZN(n12665) );
  AND2_X1 U14886 ( .A1(n13053), .A2(n13036), .ZN(n12662) );
  AOI21_X1 U14887 ( .B1(n12928), .B2(n12749), .A(n12662), .ZN(n13246) );
  OAI21_X1 U14888 ( .B1(n13246), .B2(n12751), .A(n12663), .ZN(n12664) );
  AOI211_X1 U14889 ( .C1(n13251), .C2(n14381), .A(n12665), .B(n12664), .ZN(
        n12668) );
  INV_X1 U14890 ( .A(n12666), .ZN(n12740) );
  NAND2_X1 U14891 ( .A1(n12740), .A2(n14376), .ZN(n12667) );
  OAI211_X1 U14892 ( .C1(n12670), .C2(n12669), .A(n12668), .B(n12667), .ZN(
        P2_U3191) );
  AOI21_X1 U14893 ( .B1(n12672), .B2(n12671), .A(n12759), .ZN(n12674) );
  NAND2_X1 U14894 ( .A1(n12674), .A2(n12673), .ZN(n12678) );
  AOI22_X1 U14895 ( .A1(n13050), .A2(n12749), .B1(n13036), .B2(n12928), .ZN(
        n13207) );
  OAI22_X1 U14896 ( .A1(n13207), .A2(n12751), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12675), .ZN(n12676) );
  AOI21_X1 U14897 ( .B1(n13213), .B2(n12770), .A(n12676), .ZN(n12677) );
  OAI211_X1 U14898 ( .C1(n13420), .C2(n12776), .A(n12678), .B(n12677), .ZN(
        P2_U3195) );
  AOI22_X1 U14899 ( .A1(n13046), .A2(n12749), .B1(n13036), .B2(n13048), .ZN(
        n13144) );
  AOI22_X1 U14900 ( .A1(n12770), .A2(n13149), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12679) );
  OAI21_X1 U14901 ( .B1(n13144), .B2(n12751), .A(n12679), .ZN(n12686) );
  NAND3_X1 U14902 ( .A1(n12680), .A2(n12744), .A3(n13048), .ZN(n12684) );
  OAI21_X1 U14903 ( .B1(n12726), .B2(n12681), .A(n14376), .ZN(n12683) );
  INV_X1 U14904 ( .A(n12682), .ZN(n12768) );
  AOI21_X1 U14905 ( .B1(n12684), .B2(n12683), .A(n12768), .ZN(n12685) );
  INV_X1 U14906 ( .A(n12687), .ZN(P2_U3197) );
  INV_X1 U14907 ( .A(n12690), .ZN(n12691) );
  AOI21_X1 U14908 ( .B1(n12692), .B2(n12688), .A(n12691), .ZN(n12699) );
  NAND2_X1 U14909 ( .A1(n14378), .A2(n12693), .ZN(n12695) );
  OAI211_X1 U14910 ( .C1(n14384), .C2(n12696), .A(n12695), .B(n12694), .ZN(
        n12697) );
  AOI21_X1 U14911 ( .B1(n13372), .B2(n14381), .A(n12697), .ZN(n12698) );
  OAI21_X1 U14912 ( .B1(n12699), .B2(n12759), .A(n12698), .ZN(P2_U3198) );
  OR2_X1 U14913 ( .A1(n12700), .A2(n12759), .ZN(n12712) );
  OAI22_X1 U14914 ( .A1(n12751), .A2(n12702), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12701), .ZN(n12703) );
  AOI21_X1 U14915 ( .B1(n12704), .B2(n12770), .A(n12703), .ZN(n12711) );
  INV_X1 U14916 ( .A(n12705), .ZN(n12706) );
  OAI22_X1 U14917 ( .A1(n12765), .A2(n6635), .B1(n12706), .B2(n12759), .ZN(
        n12707) );
  NAND3_X1 U14918 ( .A1(n12708), .A2(n6616), .A3(n12707), .ZN(n12710) );
  NAND2_X1 U14919 ( .A1(n14381), .A2(n12841), .ZN(n12709) );
  NAND4_X1 U14920 ( .A1(n12712), .A2(n12711), .A3(n12710), .A4(n12709), .ZN(
        P2_U3199) );
  INV_X1 U14921 ( .A(n13290), .ZN(n12716) );
  OAI22_X1 U14922 ( .A1(n12714), .A2(n12773), .B1(n12719), .B2(n12771), .ZN(
        n13279) );
  AOI22_X1 U14923 ( .A1(n14378), .A2(n13279), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12715) );
  OAI21_X1 U14924 ( .B1(n12716), .B2(n14384), .A(n12715), .ZN(n12717) );
  AOI21_X1 U14925 ( .B1(n13287), .B2(n14381), .A(n12717), .ZN(n12724) );
  INV_X1 U14926 ( .A(n12718), .ZN(n12722) );
  OAI22_X1 U14927 ( .A1(n12720), .A2(n12759), .B1(n12719), .B2(n12765), .ZN(
        n12721) );
  NAND3_X1 U14928 ( .A1(n12690), .A2(n12722), .A3(n12721), .ZN(n12723) );
  OAI211_X1 U14929 ( .C1(n12725), .C2(n12759), .A(n12724), .B(n12723), .ZN(
        P2_U3200) );
  AOI211_X1 U14930 ( .C1(n12728), .C2(n12727), .A(n12759), .B(n12726), .ZN(
        n12729) );
  INV_X1 U14931 ( .A(n12729), .ZN(n12733) );
  OAI22_X1 U14932 ( .A1(n12772), .A2(n12773), .B1(n12730), .B2(n12771), .ZN(
        n13160) );
  OAI22_X1 U14933 ( .A1(n14384), .A2(n13165), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15225), .ZN(n12731) );
  AOI21_X1 U14934 ( .B1(n13160), .B2(n14378), .A(n12731), .ZN(n12732) );
  OAI211_X1 U14935 ( .C1(n13408), .C2(n12776), .A(n12733), .B(n12732), .ZN(
        P2_U3201) );
  OAI22_X1 U14936 ( .A1(n12735), .A2(n12773), .B1(n12756), .B2(n12771), .ZN(
        n13224) );
  AOI22_X1 U14937 ( .A1(n13224), .A2(n14378), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12736) );
  OAI21_X1 U14938 ( .B1(n13227), .B2(n14384), .A(n12736), .ZN(n12742) );
  AOI22_X1 U14939 ( .A1(n12737), .A2(n14376), .B1(n12744), .B2(n13052), .ZN(
        n12739) );
  NOR3_X1 U14940 ( .A1(n12740), .A2(n12739), .A3(n12738), .ZN(n12741) );
  AOI211_X1 U14941 ( .C1(n13353), .C2(n14381), .A(n12742), .B(n12741), .ZN(
        n12743) );
  OAI21_X1 U14942 ( .B1(n12759), .B2(n12734), .A(n12743), .ZN(P2_U3205) );
  NAND2_X1 U14943 ( .A1(n12744), .A2(n13050), .ZN(n12748) );
  NAND2_X1 U14944 ( .A1(n12745), .A2(n14376), .ZN(n12747) );
  MUX2_X1 U14945 ( .A(n12748), .B(n12747), .S(n12746), .Z(n12754) );
  AOI22_X1 U14946 ( .A1(n13049), .A2(n12749), .B1(n13036), .B2(n13051), .ZN(
        n13202) );
  OAI22_X1 U14947 ( .A1(n13202), .A2(n12751), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12750), .ZN(n12752) );
  AOI21_X1 U14948 ( .B1(n13195), .B2(n12770), .A(n12752), .ZN(n12753) );
  OAI211_X1 U14949 ( .C1(n13416), .C2(n12776), .A(n12754), .B(n12753), .ZN(
        P2_U3207) );
  OAI22_X1 U14950 ( .A1(n12756), .A2(n12773), .B1(n12755), .B2(n12771), .ZN(
        n13261) );
  NAND2_X1 U14951 ( .A1(n14378), .A2(n13261), .ZN(n12757) );
  NAND2_X1 U14952 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14812)
         );
  OAI211_X1 U14953 ( .C1(n14384), .C2(n13270), .A(n12757), .B(n14812), .ZN(
        n12763) );
  AOI211_X1 U14954 ( .C1(n12761), .C2(n12760), .A(n12759), .B(n12758), .ZN(
        n12762) );
  AOI211_X1 U14955 ( .C1(n13269), .C2(n14381), .A(n12763), .B(n12762), .ZN(
        n12764) );
  INV_X1 U14956 ( .A(n12764), .ZN(P2_U3210) );
  NOR3_X1 U14957 ( .A1(n12766), .A2(n12772), .A3(n12765), .ZN(n12767) );
  AOI21_X1 U14958 ( .B1(n12768), .B2(n14376), .A(n12767), .ZN(n12781) );
  INV_X1 U14959 ( .A(n12769), .ZN(n12778) );
  AOI22_X1 U14960 ( .A1(n13135), .A2(n12770), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12775) );
  OAI22_X1 U14961 ( .A1(n12956), .A2(n12773), .B1(n12772), .B2(n12771), .ZN(
        n13132) );
  NAND2_X1 U14962 ( .A1(n13132), .A2(n14378), .ZN(n12774) );
  OAI211_X1 U14963 ( .C1(n13137), .C2(n12776), .A(n12775), .B(n12774), .ZN(
        n12777) );
  AOI21_X1 U14964 ( .B1(n12778), .B2(n14376), .A(n12777), .ZN(n12779) );
  OAI21_X1 U14965 ( .B1(n12781), .B2(n12780), .A(n12779), .ZN(P2_U3212) );
  INV_X1 U14966 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n12789) );
  NAND2_X1 U14967 ( .A1(n12785), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n12788) );
  NAND2_X1 U14968 ( .A1(n12786), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n12787) );
  OAI211_X1 U14969 ( .C1(n12790), .C2(n12789), .A(n12788), .B(n12787), .ZN(
        n13091) );
  NAND2_X1 U14970 ( .A1(n13029), .A2(n12982), .ZN(n12792) );
  AOI211_X1 U14971 ( .C1(n6461), .C2(n13091), .A(n12792), .B(n12978), .ZN(
        n12793) );
  OAI22_X1 U14972 ( .A1(n13022), .A2(n6461), .B1(n12794), .B2(n12793), .ZN(
        n12970) );
  MUX2_X1 U14973 ( .A(n12794), .B(n13022), .S(n6461), .Z(n12971) );
  INV_X1 U14974 ( .A(n12795), .ZN(n13043) );
  MUX2_X1 U14975 ( .A(n13043), .B(n13308), .S(n6461), .Z(n12805) );
  INV_X1 U14976 ( .A(n12805), .ZN(n12798) );
  INV_X1 U14977 ( .A(n12806), .ZN(n12797) );
  NAND2_X1 U14978 ( .A1(n12799), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n12800) );
  AND2_X1 U14979 ( .A1(n13088), .A2(n12804), .ZN(n12801) );
  OAI21_X1 U14980 ( .B1(n13038), .B2(n13026), .A(n7737), .ZN(n12809) );
  NAND2_X1 U14981 ( .A1(n12810), .A2(n12809), .ZN(n12813) );
  NAND2_X1 U14982 ( .A1(n12811), .A2(n6461), .ZN(n12812) );
  NAND2_X1 U14983 ( .A1(n12813), .A2(n12812), .ZN(n12818) );
  MUX2_X1 U14984 ( .A(n12815), .B(n13070), .S(n12814), .Z(n12819) );
  NAND2_X1 U14985 ( .A1(n12818), .A2(n12819), .ZN(n12817) );
  MUX2_X1 U14986 ( .A(n13070), .B(n12815), .S(n12814), .Z(n12816) );
  NAND2_X1 U14987 ( .A1(n12817), .A2(n12816), .ZN(n12823) );
  INV_X1 U14988 ( .A(n12818), .ZN(n12821) );
  INV_X1 U14989 ( .A(n12819), .ZN(n12820) );
  NAND2_X1 U14990 ( .A1(n12821), .A2(n12820), .ZN(n12822) );
  NAND2_X1 U14991 ( .A1(n12823), .A2(n12822), .ZN(n12827) );
  MUX2_X1 U14992 ( .A(n13069), .B(n12824), .S(n6461), .Z(n12828) );
  NAND2_X1 U14993 ( .A1(n12827), .A2(n12828), .ZN(n12826) );
  MUX2_X1 U14994 ( .A(n12824), .B(n13069), .S(n6461), .Z(n12825) );
  NAND2_X1 U14995 ( .A1(n12826), .A2(n12825), .ZN(n12832) );
  INV_X1 U14996 ( .A(n12827), .ZN(n12830) );
  INV_X1 U14997 ( .A(n12828), .ZN(n12829) );
  NAND2_X1 U14998 ( .A1(n12830), .A2(n12829), .ZN(n12831) );
  MUX2_X1 U14999 ( .A(n13068), .B(n12833), .S(n6461), .Z(n12834) );
  MUX2_X1 U15000 ( .A(n13067), .B(n12836), .S(n6461), .Z(n12839) );
  MUX2_X1 U15001 ( .A(n13067), .B(n12836), .S(n12872), .Z(n12837) );
  INV_X1 U15002 ( .A(n12839), .ZN(n12840) );
  MUX2_X1 U15003 ( .A(n13066), .B(n12841), .S(n12852), .Z(n12845) );
  MUX2_X1 U15004 ( .A(n13066), .B(n12841), .S(n6461), .Z(n12842) );
  INV_X1 U15005 ( .A(n12844), .ZN(n12847) );
  INV_X1 U15006 ( .A(n12845), .ZN(n12846) );
  MUX2_X1 U15007 ( .A(n13065), .B(n12849), .S(n6461), .Z(n12851) );
  MUX2_X1 U15008 ( .A(n13065), .B(n12849), .S(n12852), .Z(n12850) );
  MUX2_X1 U15009 ( .A(n13064), .B(n12853), .S(n12852), .Z(n12857) );
  NAND2_X1 U15010 ( .A1(n12856), .A2(n12857), .ZN(n12855) );
  MUX2_X1 U15011 ( .A(n13064), .B(n12853), .S(n6461), .Z(n12854) );
  NAND2_X1 U15012 ( .A1(n12855), .A2(n12854), .ZN(n12861) );
  INV_X1 U15013 ( .A(n12856), .ZN(n12859) );
  INV_X1 U15014 ( .A(n12857), .ZN(n12858) );
  NAND2_X1 U15015 ( .A1(n12859), .A2(n12858), .ZN(n12860) );
  MUX2_X1 U15016 ( .A(n13063), .B(n14885), .S(n6461), .Z(n12863) );
  MUX2_X1 U15017 ( .A(n13063), .B(n14885), .S(n12872), .Z(n12862) );
  INV_X1 U15018 ( .A(n12863), .ZN(n12864) );
  MUX2_X1 U15019 ( .A(n13062), .B(n12865), .S(n12872), .Z(n12868) );
  MUX2_X1 U15020 ( .A(n13062), .B(n12865), .S(n6461), .Z(n12866) );
  INV_X1 U15021 ( .A(n12867), .ZN(n12870) );
  INV_X1 U15022 ( .A(n12868), .ZN(n12869) );
  MUX2_X1 U15023 ( .A(n13061), .B(n14892), .S(n6461), .Z(n12874) );
  MUX2_X1 U15024 ( .A(n13061), .B(n14892), .S(n12872), .Z(n12873) );
  MUX2_X1 U15025 ( .A(n13060), .B(n12875), .S(n12872), .Z(n12879) );
  NAND2_X1 U15026 ( .A1(n12878), .A2(n12879), .ZN(n12877) );
  MUX2_X1 U15027 ( .A(n13060), .B(n12875), .S(n6461), .Z(n12876) );
  INV_X1 U15028 ( .A(n12878), .ZN(n12881) );
  INV_X1 U15029 ( .A(n12879), .ZN(n12880) );
  NAND2_X1 U15030 ( .A1(n12881), .A2(n12880), .ZN(n12882) );
  MUX2_X1 U15031 ( .A(n13059), .B(n12883), .S(n6461), .Z(n12885) );
  MUX2_X1 U15032 ( .A(n13059), .B(n12883), .S(n12872), .Z(n12884) );
  MUX2_X1 U15033 ( .A(n13058), .B(n13386), .S(n12872), .Z(n12898) );
  MUX2_X1 U15034 ( .A(n12887), .B(n12886), .S(n12872), .Z(n12902) );
  MUX2_X1 U15035 ( .A(n13056), .B(n13435), .S(n6461), .Z(n12903) );
  NAND2_X1 U15036 ( .A1(n12902), .A2(n12903), .ZN(n12891) );
  AND2_X1 U15037 ( .A1(n13055), .A2(n12872), .ZN(n12889) );
  OAI21_X1 U15038 ( .B1(n12872), .B2(n13055), .A(n13372), .ZN(n12888) );
  OAI21_X1 U15039 ( .B1(n12889), .B2(n13372), .A(n12888), .ZN(n12890) );
  AND2_X1 U15040 ( .A1(n13283), .A2(n12890), .ZN(n12907) );
  MUX2_X1 U15041 ( .A(n12893), .B(n12892), .S(n12872), .Z(n12910) );
  MUX2_X1 U15042 ( .A(n13057), .B(n14380), .S(n6461), .Z(n12909) );
  NAND2_X1 U15043 ( .A1(n12910), .A2(n12909), .ZN(n12894) );
  OAI211_X1 U15044 ( .C1(n12899), .C2(n12898), .A(n12908), .B(n12894), .ZN(
        n12901) );
  MUX2_X1 U15045 ( .A(n12896), .B(n12895), .S(n6461), .Z(n12897) );
  AOI21_X1 U15046 ( .B1(n12899), .B2(n12898), .A(n12897), .ZN(n12900) );
  INV_X1 U15047 ( .A(n12902), .ZN(n12906) );
  INV_X1 U15048 ( .A(n12903), .ZN(n12905) );
  AOI21_X1 U15049 ( .B1(n12906), .B2(n12905), .A(n12904), .ZN(n12917) );
  INV_X1 U15050 ( .A(n12907), .ZN(n12916) );
  INV_X1 U15051 ( .A(n12908), .ZN(n12911) );
  OR3_X1 U15052 ( .A1(n12911), .A2(n12910), .A3(n12909), .ZN(n12915) );
  MUX2_X1 U15053 ( .A(n12913), .B(n12912), .S(n6461), .Z(n12914) );
  OAI211_X1 U15054 ( .C1(n12917), .C2(n12916), .A(n12915), .B(n12914), .ZN(
        n12918) );
  INV_X1 U15055 ( .A(n12918), .ZN(n12919) );
  MUX2_X1 U15056 ( .A(n13053), .B(n13269), .S(n6461), .Z(n12920) );
  INV_X1 U15057 ( .A(n12920), .ZN(n12922) );
  MUX2_X1 U15058 ( .A(n13269), .B(n13053), .S(n6461), .Z(n12921) );
  MUX2_X1 U15059 ( .A(n13052), .B(n13251), .S(n12872), .Z(n12926) );
  NAND2_X1 U15060 ( .A1(n12925), .A2(n12926), .ZN(n12924) );
  MUX2_X1 U15061 ( .A(n13052), .B(n13251), .S(n6461), .Z(n12923) );
  MUX2_X1 U15062 ( .A(n13353), .B(n12928), .S(n12872), .Z(n12930) );
  MUX2_X1 U15063 ( .A(n13353), .B(n12928), .S(n6461), .Z(n12929) );
  MUX2_X1 U15064 ( .A(n13212), .B(n13051), .S(n6461), .Z(n12934) );
  NAND2_X1 U15065 ( .A1(n12933), .A2(n12934), .ZN(n12932) );
  MUX2_X1 U15066 ( .A(n13051), .B(n13212), .S(n6461), .Z(n12931) );
  NAND2_X1 U15067 ( .A1(n12932), .A2(n12931), .ZN(n12938) );
  INV_X1 U15068 ( .A(n12933), .ZN(n12936) );
  INV_X1 U15069 ( .A(n12934), .ZN(n12935) );
  NAND2_X1 U15070 ( .A1(n12936), .A2(n12935), .ZN(n12937) );
  MUX2_X1 U15071 ( .A(n13050), .B(n13194), .S(n6461), .Z(n12940) );
  MUX2_X1 U15072 ( .A(n13194), .B(n13050), .S(n6461), .Z(n12939) );
  INV_X1 U15073 ( .A(n12940), .ZN(n12941) );
  MUX2_X1 U15074 ( .A(n13182), .B(n13049), .S(n6461), .Z(n12944) );
  MUX2_X1 U15075 ( .A(n13049), .B(n13182), .S(n6461), .Z(n12942) );
  INV_X1 U15076 ( .A(n12944), .ZN(n12945) );
  MUX2_X1 U15077 ( .A(n12946), .B(n13048), .S(n12872), .Z(n12949) );
  MUX2_X1 U15078 ( .A(n12946), .B(n13048), .S(n6461), .Z(n12947) );
  NAND2_X1 U15079 ( .A1(n12948), .A2(n12947), .ZN(n12951) );
  MUX2_X1 U15080 ( .A(n13047), .B(n13327), .S(n12872), .Z(n12953) );
  MUX2_X1 U15081 ( .A(n13047), .B(n13327), .S(n6461), .Z(n12952) );
  MUX2_X1 U15082 ( .A(n13046), .B(n13322), .S(n6461), .Z(n12954) );
  MUX2_X1 U15083 ( .A(n13322), .B(n13046), .S(n6461), .Z(n12955) );
  MUX2_X1 U15084 ( .A(n13402), .B(n12956), .S(n6461), .Z(n12959) );
  MUX2_X1 U15085 ( .A(n13111), .B(n12957), .S(n6461), .Z(n12964) );
  MUX2_X1 U15086 ( .A(n13044), .B(n13314), .S(n6461), .Z(n12963) );
  AOI22_X1 U15087 ( .A1(n12960), .A2(n12959), .B1(n12964), .B2(n12963), .ZN(
        n12962) );
  MUX2_X1 U15088 ( .A(n13045), .B(n13124), .S(n6461), .Z(n12958) );
  OAI21_X1 U15089 ( .B1(n12960), .B2(n12959), .A(n12958), .ZN(n12961) );
  NAND3_X1 U15090 ( .A1(n6542), .A2(n12962), .A3(n12961), .ZN(n12968) );
  INV_X1 U15091 ( .A(n12963), .ZN(n12966) );
  INV_X1 U15092 ( .A(n12964), .ZN(n12965) );
  NAND3_X1 U15093 ( .A1(n6542), .A2(n12966), .A3(n12965), .ZN(n12967) );
  INV_X1 U15094 ( .A(n12970), .ZN(n12973) );
  INV_X1 U15095 ( .A(n12971), .ZN(n12972) );
  NAND2_X1 U15096 ( .A1(n12973), .A2(n12972), .ZN(n12977) );
  NOR3_X1 U15097 ( .A1(n13393), .A2(n12872), .A3(n13091), .ZN(n12975) );
  NOR3_X1 U15098 ( .A1(n13088), .A2(n12804), .A3(n6461), .ZN(n12974) );
  INV_X1 U15099 ( .A(n12978), .ZN(n12981) );
  NAND3_X1 U15100 ( .A1(n13029), .A2(n12979), .A3(n7734), .ZN(n12980) );
  NAND2_X1 U15101 ( .A1(n13029), .A2(n13026), .ZN(n12983) );
  OAI211_X1 U15102 ( .C1(n13038), .C2(n12984), .A(n12983), .B(n12982), .ZN(
        n12985) );
  NAND2_X1 U15103 ( .A1(n13031), .A2(n12985), .ZN(n12986) );
  OAI21_X1 U15104 ( .B1(n13031), .B2(n7508), .A(n12986), .ZN(n13033) );
  NAND2_X1 U15105 ( .A1(n12988), .A2(n12987), .ZN(n13138) );
  NAND4_X1 U15106 ( .A1(n12992), .A2(n7734), .A3(n6735), .A4(n14838), .ZN(
        n12993) );
  NOR2_X1 U15107 ( .A1(n12994), .A2(n12993), .ZN(n12995) );
  NAND2_X1 U15108 ( .A1(n12996), .A2(n12995), .ZN(n12997) );
  NOR2_X1 U15109 ( .A1(n12998), .A2(n12997), .ZN(n13001) );
  NAND4_X1 U15110 ( .A1(n13002), .A2(n13001), .A3(n13000), .A4(n12999), .ZN(
        n13003) );
  NOR2_X1 U15111 ( .A1(n13004), .A2(n13003), .ZN(n13006) );
  NAND4_X1 U15112 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13009) );
  NOR2_X1 U15113 ( .A1(n13010), .A2(n13009), .ZN(n13012) );
  NAND4_X1 U15114 ( .A1(n13283), .A2(n13013), .A3(n13012), .A4(n13011), .ZN(
        n13014) );
  NOR4_X1 U15115 ( .A1(n13242), .A2(n13266), .A3(n13015), .A4(n13014), .ZN(
        n13017) );
  NAND4_X1 U15116 ( .A1(n13201), .A2(n13017), .A3(n13220), .A4(n13016), .ZN(
        n13018) );
  NOR4_X1 U15117 ( .A1(n13138), .A2(n13179), .A3(n13163), .A4(n13018), .ZN(
        n13019) );
  NAND4_X1 U15118 ( .A1(n13112), .A2(n13019), .A3(n13152), .A4(n13120), .ZN(
        n13021) );
  INV_X1 U15119 ( .A(n13022), .ZN(n13023) );
  NAND3_X1 U15120 ( .A1(n13025), .A2(n13024), .A3(n7507), .ZN(n13027) );
  NOR2_X1 U15121 ( .A1(n13033), .A2(n13032), .ZN(n13041) );
  NAND4_X1 U15122 ( .A1(n14835), .A2(n13036), .A3(n13035), .A4(n13034), .ZN(
        n13037) );
  OAI211_X1 U15123 ( .C1(n13038), .C2(n13040), .A(n13037), .B(P2_B_REG_SCAN_IN), .ZN(n13039) );
  OAI21_X1 U15124 ( .B1(n13041), .B2(n13040), .A(n13039), .ZN(P2_U3328) );
  MUX2_X1 U15125 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13091), .S(n13071), .Z(
        P2_U3562) );
  MUX2_X1 U15126 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13042), .S(n13071), .Z(
        P2_U3561) );
  MUX2_X1 U15127 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13043), .S(n13071), .Z(
        P2_U3560) );
  MUX2_X1 U15128 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13044), .S(n13071), .Z(
        P2_U3559) );
  MUX2_X1 U15129 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13045), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15130 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13046), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15131 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13047), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15132 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13048), .S(n13071), .Z(
        P2_U3555) );
  MUX2_X1 U15133 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13049), .S(n13071), .Z(
        P2_U3554) );
  MUX2_X1 U15134 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13050), .S(n13071), .Z(
        P2_U3553) );
  MUX2_X1 U15135 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13051), .S(n13071), .Z(
        P2_U3552) );
  MUX2_X1 U15136 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13052), .S(n13071), .Z(
        P2_U3550) );
  MUX2_X1 U15137 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13053), .S(n13071), .Z(
        P2_U3549) );
  MUX2_X1 U15138 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13054), .S(n13071), .Z(
        P2_U3548) );
  MUX2_X1 U15139 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13055), .S(n13071), .Z(
        P2_U3547) );
  MUX2_X1 U15140 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13056), .S(n13071), .Z(
        P2_U3546) );
  MUX2_X1 U15141 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13057), .S(n13071), .Z(
        P2_U3545) );
  MUX2_X1 U15142 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13058), .S(n13071), .Z(
        P2_U3544) );
  MUX2_X1 U15143 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13059), .S(n13071), .Z(
        P2_U3543) );
  MUX2_X1 U15144 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13060), .S(n13071), .Z(
        P2_U3542) );
  MUX2_X1 U15145 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13061), .S(n13071), .Z(
        P2_U3541) );
  MUX2_X1 U15146 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13062), .S(n13071), .Z(
        P2_U3540) );
  MUX2_X1 U15147 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13063), .S(n13071), .Z(
        P2_U3539) );
  MUX2_X1 U15148 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13064), .S(n13071), .Z(
        P2_U3538) );
  MUX2_X1 U15149 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13065), .S(n13071), .Z(
        P2_U3537) );
  MUX2_X1 U15150 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13066), .S(n13071), .Z(
        P2_U3536) );
  MUX2_X1 U15151 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13067), .S(n13071), .Z(
        P2_U3535) );
  MUX2_X1 U15152 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13068), .S(n13071), .Z(
        P2_U3534) );
  MUX2_X1 U15153 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13069), .S(n13071), .Z(
        P2_U3533) );
  MUX2_X1 U15154 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13070), .S(n13071), .Z(
        P2_U3532) );
  MUX2_X1 U15155 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13072), .S(n13071), .Z(
        P2_U3531) );
  NOR2_X1 U15156 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13073), .ZN(n13075) );
  NOR2_X1 U15157 ( .A1(n14827), .A2(n13079), .ZN(n13074) );
  AOI211_X1 U15158 ( .C1(n14819), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n13075), .B(
        n13074), .ZN(n13087) );
  OAI211_X1 U15159 ( .C1(n13078), .C2(n13077), .A(n14784), .B(n13076), .ZN(
        n13086) );
  MUX2_X1 U15160 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10217), .S(n13079), .Z(
        n13080) );
  NAND3_X1 U15161 ( .A1(n13082), .A2(n13081), .A3(n13080), .ZN(n13083) );
  NAND3_X1 U15162 ( .A1(n14805), .A2(n13084), .A3(n13083), .ZN(n13085) );
  NAND3_X1 U15163 ( .A1(n13087), .A2(n13086), .A3(n13085), .ZN(P2_U3222) );
  NAND2_X1 U15164 ( .A1(n13300), .A2(n13288), .ZN(n13094) );
  AND2_X1 U15165 ( .A1(n13092), .A2(n13091), .ZN(n13299) );
  INV_X1 U15166 ( .A(n13299), .ZN(n13303) );
  NOR2_X1 U15167 ( .A1(n13298), .A2(n13303), .ZN(n13098) );
  AOI21_X1 U15168 ( .B1(n13298), .B2(P2_REG2_REG_31__SCAN_IN), .A(n13098), 
        .ZN(n13093) );
  OAI211_X1 U15169 ( .C1(n13393), .C2(n13293), .A(n13094), .B(n13093), .ZN(
        P2_U3234) );
  OAI211_X1 U15170 ( .C1(n13022), .C2(n13096), .A(n13106), .B(n13095), .ZN(
        n13304) );
  NOR2_X1 U15171 ( .A1(n13022), .A2(n13293), .ZN(n13097) );
  AOI211_X1 U15172 ( .C1(n13298), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13098), 
        .B(n13097), .ZN(n13099) );
  OAI21_X1 U15173 ( .B1(n13184), .B2(n13304), .A(n13099), .ZN(P2_U3235) );
  NAND2_X1 U15174 ( .A1(n13100), .A2(n13198), .ZN(n13104) );
  OAI21_X1 U15175 ( .B1(n13104), .B2(n13103), .A(n13102), .ZN(n13312) );
  AOI21_X1 U15176 ( .B1(n13105), .B2(n13289), .A(n13312), .ZN(n13115) );
  OAI21_X1 U15177 ( .B1(n13111), .B2(n13122), .A(n13106), .ZN(n13107) );
  OR2_X1 U15178 ( .A1(n13108), .A2(n13107), .ZN(n13109) );
  INV_X1 U15179 ( .A(n13109), .ZN(n13313) );
  OAI22_X1 U15180 ( .A1(n13111), .A2(n13293), .B1(n13248), .B2(n13110), .ZN(
        n13114) );
  OAI21_X1 U15181 ( .B1(n13117), .B2(n13120), .A(n13116), .ZN(n13119) );
  XNOR2_X1 U15182 ( .A(n13121), .B(n13120), .ZN(n13318) );
  NAND2_X1 U15183 ( .A1(n13318), .A2(n13295), .ZN(n13130) );
  INV_X1 U15184 ( .A(n13134), .ZN(n13123) );
  AOI211_X1 U15185 ( .C1(n13124), .C2(n13123), .A(n13089), .B(n13122), .ZN(
        n13317) );
  NOR2_X1 U15186 ( .A1(n13402), .A2(n13293), .ZN(n13128) );
  OAI22_X1 U15187 ( .A1(n13126), .A2(n13226), .B1(n13125), .B2(n13248), .ZN(
        n13127) );
  AOI211_X1 U15188 ( .C1(n13317), .C2(n13288), .A(n13128), .B(n13127), .ZN(
        n13129) );
  OAI211_X1 U15189 ( .C1(n13298), .C2(n13316), .A(n13130), .B(n13129), .ZN(
        P2_U3238) );
  XNOR2_X1 U15190 ( .A(n13131), .B(n13138), .ZN(n13133) );
  AOI21_X1 U15191 ( .B1(n13133), .B2(n13198), .A(n13132), .ZN(n13324) );
  AOI211_X1 U15192 ( .C1(n13322), .C2(n13147), .A(n13089), .B(n13134), .ZN(
        n13321) );
  AOI22_X1 U15193 ( .A1(n13135), .A2(n13289), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13298), .ZN(n13136) );
  OAI21_X1 U15194 ( .B1(n13137), .B2(n13293), .A(n13136), .ZN(n13141) );
  XNOR2_X1 U15195 ( .A(n13139), .B(n13138), .ZN(n13325) );
  NOR2_X1 U15196 ( .A1(n13325), .A2(n13238), .ZN(n13140) );
  AOI211_X1 U15197 ( .C1(n13321), .C2(n13288), .A(n13141), .B(n13140), .ZN(
        n13142) );
  OAI21_X1 U15198 ( .B1(n13298), .B2(n13324), .A(n13142), .ZN(P2_U3239) );
  XNOR2_X1 U15199 ( .A(n13143), .B(n13152), .ZN(n13146) );
  INV_X1 U15200 ( .A(n13144), .ZN(n13145) );
  AOI21_X1 U15201 ( .B1(n13146), .B2(n13198), .A(n13145), .ZN(n13328) );
  INV_X1 U15202 ( .A(n13147), .ZN(n13148) );
  AOI211_X1 U15203 ( .C1(n13327), .C2(n13168), .A(n13089), .B(n13148), .ZN(
        n13326) );
  AOI22_X1 U15204 ( .A1(n13149), .A2(n13289), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13298), .ZN(n13150) );
  OAI21_X1 U15205 ( .B1(n7044), .B2(n13293), .A(n13150), .ZN(n13154) );
  XOR2_X1 U15206 ( .A(n13151), .B(n13152), .Z(n13330) );
  NOR2_X1 U15207 ( .A1(n13330), .A2(n13238), .ZN(n13153) );
  AOI211_X1 U15208 ( .C1(n13326), .C2(n13288), .A(n13154), .B(n13153), .ZN(
        n13155) );
  OAI21_X1 U15209 ( .B1(n13298), .B2(n13328), .A(n13155), .ZN(P2_U3240) );
  AND2_X1 U15210 ( .A1(n7518), .A2(n13156), .ZN(n13158) );
  OAI21_X1 U15211 ( .B1(n13159), .B2(n13158), .A(n13157), .ZN(n13161) );
  AOI21_X1 U15212 ( .B1(n13161), .B2(n13198), .A(n13160), .ZN(n13332) );
  OAI21_X1 U15213 ( .B1(n13164), .B2(n13163), .A(n13162), .ZN(n13333) );
  INV_X1 U15214 ( .A(n13333), .ZN(n13171) );
  INV_X1 U15215 ( .A(n13165), .ZN(n13166) );
  AOI22_X1 U15216 ( .A1(n13166), .A2(n13289), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13298), .ZN(n13167) );
  OAI21_X1 U15217 ( .B1(n13408), .B2(n13293), .A(n13167), .ZN(n13170) );
  OAI211_X1 U15218 ( .C1(n13408), .C2(n6481), .A(n13106), .B(n13168), .ZN(
        n13331) );
  NOR2_X1 U15219 ( .A1(n13331), .A2(n13184), .ZN(n13169) );
  AOI211_X1 U15220 ( .C1(n13171), .C2(n13295), .A(n13170), .B(n13169), .ZN(
        n13172) );
  OAI21_X1 U15221 ( .B1(n13298), .B2(n13332), .A(n13172), .ZN(P2_U3241) );
  AOI21_X1 U15222 ( .B1(n13179), .B2(n6582), .A(n13281), .ZN(n13175) );
  INV_X1 U15223 ( .A(n13173), .ZN(n13174) );
  AOI21_X1 U15224 ( .B1(n13175), .B2(n7518), .A(n13174), .ZN(n13339) );
  INV_X1 U15225 ( .A(n13339), .ZN(n13176) );
  AOI21_X1 U15226 ( .B1(n13177), .B2(n13289), .A(n13176), .ZN(n13187) );
  XNOR2_X1 U15227 ( .A(n13179), .B(n13178), .ZN(n13336) );
  NAND2_X1 U15228 ( .A1(n13182), .A2(n13191), .ZN(n13180) );
  NAND2_X1 U15229 ( .A1(n13180), .A2(n13106), .ZN(n13181) );
  OR2_X1 U15230 ( .A1(n6481), .A2(n13181), .ZN(n13337) );
  AOI22_X1 U15231 ( .A1(n13182), .A2(n13230), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n13298), .ZN(n13183) );
  OAI21_X1 U15232 ( .B1(n13337), .B2(n13184), .A(n13183), .ZN(n13185) );
  AOI21_X1 U15233 ( .B1(n13295), .B2(n13336), .A(n13185), .ZN(n13186) );
  OAI21_X1 U15234 ( .B1(n13187), .B2(n13298), .A(n13186), .ZN(P2_U3242) );
  OAI21_X1 U15235 ( .B1(n13190), .B2(n13189), .A(n13188), .ZN(n13342) );
  INV_X1 U15236 ( .A(n13211), .ZN(n13193) );
  INV_X1 U15237 ( .A(n13191), .ZN(n13192) );
  AOI211_X1 U15238 ( .C1(n13194), .C2(n13193), .A(n13089), .B(n13192), .ZN(
        n13343) );
  AOI22_X1 U15239 ( .A1(n13298), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13195), 
        .B2(n13289), .ZN(n13196) );
  OAI21_X1 U15240 ( .B1(n13416), .B2(n13293), .A(n13196), .ZN(n13197) );
  AOI21_X1 U15241 ( .B1(n13343), .B2(n13288), .A(n13197), .ZN(n13205) );
  OAI211_X1 U15242 ( .C1(n13201), .C2(n13200), .A(n13199), .B(n13198), .ZN(
        n13203) );
  NAND2_X1 U15243 ( .A1(n13203), .A2(n13202), .ZN(n13344) );
  NAND2_X1 U15244 ( .A1(n13344), .A2(n13248), .ZN(n13204) );
  OAI211_X1 U15245 ( .C1(n13342), .C2(n13238), .A(n13205), .B(n13204), .ZN(
        P2_U3243) );
  XNOR2_X1 U15246 ( .A(n13210), .B(n13206), .ZN(n13208) );
  OAI21_X1 U15247 ( .B1(n13208), .B2(n13281), .A(n13207), .ZN(n13348) );
  INV_X1 U15248 ( .A(n13348), .ZN(n13218) );
  XNOR2_X1 U15249 ( .A(n13210), .B(n13209), .ZN(n13350) );
  AOI211_X1 U15250 ( .C1(n13212), .C2(n13232), .A(n13089), .B(n13211), .ZN(
        n13349) );
  NAND2_X1 U15251 ( .A1(n13349), .A2(n13288), .ZN(n13215) );
  AOI22_X1 U15252 ( .A1(n13298), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n13213), 
        .B2(n13289), .ZN(n13214) );
  OAI211_X1 U15253 ( .C1(n13420), .C2(n13293), .A(n13215), .B(n13214), .ZN(
        n13216) );
  AOI21_X1 U15254 ( .B1(n13295), .B2(n13350), .A(n13216), .ZN(n13217) );
  OAI21_X1 U15255 ( .B1(n13298), .B2(n13218), .A(n13217), .ZN(P2_U3244) );
  XNOR2_X1 U15256 ( .A(n13219), .B(n13220), .ZN(n13356) );
  INV_X1 U15257 ( .A(n13220), .ZN(n13221) );
  NAND3_X1 U15258 ( .A1(n13221), .A2(n13243), .A3(n13240), .ZN(n13223) );
  AOI21_X1 U15259 ( .B1(n13223), .B2(n13222), .A(n13281), .ZN(n13225) );
  NOR2_X1 U15260 ( .A1(n13225), .A2(n13224), .ZN(n13355) );
  OAI22_X1 U15261 ( .A1(n13248), .A2(n13228), .B1(n13227), .B2(n13226), .ZN(
        n13229) );
  AOI21_X1 U15262 ( .B1(n13353), .B2(n13230), .A(n13229), .ZN(n13235) );
  AOI21_X1 U15263 ( .B1(n13353), .B2(n13249), .A(n13231), .ZN(n13233) );
  AND2_X1 U15264 ( .A1(n13233), .A2(n13232), .ZN(n13352) );
  NAND2_X1 U15265 ( .A1(n13352), .A2(n13288), .ZN(n13234) );
  OAI211_X1 U15266 ( .C1(n13355), .C2(n13298), .A(n13235), .B(n13234), .ZN(
        n13236) );
  INV_X1 U15267 ( .A(n13236), .ZN(n13237) );
  OAI21_X1 U15268 ( .B1(n13238), .B2(n13356), .A(n13237), .ZN(P2_U3245) );
  XNOR2_X1 U15269 ( .A(n13239), .B(n13242), .ZN(n13359) );
  INV_X1 U15270 ( .A(n13359), .ZN(n13259) );
  INV_X1 U15271 ( .A(n13240), .ZN(n13244) );
  AOI22_X1 U15272 ( .A1(n13244), .A2(n13243), .B1(n13242), .B2(n13241), .ZN(
        n13247) );
  NAND2_X1 U15273 ( .A1(n13359), .A2(n14890), .ZN(n13245) );
  OAI211_X1 U15274 ( .C1(n13247), .C2(n13281), .A(n13246), .B(n13245), .ZN(
        n13357) );
  NAND2_X1 U15275 ( .A1(n13357), .A2(n13248), .ZN(n13257) );
  INV_X1 U15276 ( .A(n13249), .ZN(n13250) );
  AOI211_X1 U15277 ( .C1(n13251), .C2(n13267), .A(n13089), .B(n13250), .ZN(
        n13358) );
  INV_X1 U15278 ( .A(n13251), .ZN(n13425) );
  INV_X1 U15279 ( .A(n13252), .ZN(n13253) );
  AOI22_X1 U15280 ( .A1(n13298), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13253), 
        .B2(n13289), .ZN(n13254) );
  OAI21_X1 U15281 ( .B1(n13425), .B2(n13293), .A(n13254), .ZN(n13255) );
  AOI21_X1 U15282 ( .B1(n13358), .B2(n13288), .A(n13255), .ZN(n13256) );
  OAI211_X1 U15283 ( .C1(n13259), .C2(n13258), .A(n13257), .B(n13256), .ZN(
        P2_U3246) );
  XNOR2_X1 U15284 ( .A(n13260), .B(n13266), .ZN(n13263) );
  INV_X1 U15285 ( .A(n13261), .ZN(n13262) );
  OAI21_X1 U15286 ( .B1(n13263), .B2(n13281), .A(n13262), .ZN(n13361) );
  INV_X1 U15287 ( .A(n13361), .ZN(n13276) );
  OAI21_X1 U15288 ( .B1(n7095), .B2(n13266), .A(n13265), .ZN(n13363) );
  INV_X1 U15289 ( .A(n13267), .ZN(n13268) );
  AOI211_X1 U15290 ( .C1(n13269), .C2(n7043), .A(n13089), .B(n13268), .ZN(
        n13362) );
  NAND2_X1 U15291 ( .A1(n13362), .A2(n13288), .ZN(n13273) );
  INV_X1 U15292 ( .A(n13270), .ZN(n13271) );
  AOI22_X1 U15293 ( .A1(n13298), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13271), 
        .B2(n13289), .ZN(n13272) );
  OAI211_X1 U15294 ( .C1(n13429), .C2(n13293), .A(n13273), .B(n13272), .ZN(
        n13274) );
  AOI21_X1 U15295 ( .B1(n13295), .B2(n13363), .A(n13274), .ZN(n13275) );
  OAI21_X1 U15296 ( .B1(n13298), .B2(n13276), .A(n13275), .ZN(P2_U3247) );
  XNOR2_X1 U15297 ( .A(n13278), .B(n13277), .ZN(n13282) );
  INV_X1 U15298 ( .A(n13279), .ZN(n13280) );
  OAI21_X1 U15299 ( .B1(n13282), .B2(n13281), .A(n13280), .ZN(n13365) );
  INV_X1 U15300 ( .A(n13365), .ZN(n13297) );
  XNOR2_X1 U15301 ( .A(n13284), .B(n13283), .ZN(n13367) );
  AOI211_X1 U15302 ( .C1(n13287), .C2(n13286), .A(n13089), .B(n13285), .ZN(
        n13366) );
  NAND2_X1 U15303 ( .A1(n13366), .A2(n13288), .ZN(n13292) );
  AOI22_X1 U15304 ( .A1(n13298), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13290), 
        .B2(n13289), .ZN(n13291) );
  OAI211_X1 U15305 ( .C1(n7041), .C2(n13293), .A(n13292), .B(n13291), .ZN(
        n13294) );
  AOI21_X1 U15306 ( .B1(n13295), .B2(n13367), .A(n13294), .ZN(n13296) );
  OAI21_X1 U15307 ( .B1(n13298), .B2(n13297), .A(n13296), .ZN(P2_U3248) );
  INV_X1 U15308 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n13301) );
  NOR2_X1 U15309 ( .A1(n13300), .A2(n13299), .ZN(n13390) );
  MUX2_X1 U15310 ( .A(n13301), .B(n13390), .S(n14912), .Z(n13302) );
  OAI21_X1 U15311 ( .B1(n13393), .B2(n13370), .A(n13302), .ZN(P2_U3530) );
  NAND2_X1 U15312 ( .A1(n13304), .A2(n13303), .ZN(n13394) );
  MUX2_X1 U15313 ( .A(n13394), .B(P2_REG1_REG_30__SCAN_IN), .S(n14910), .Z(
        n13305) );
  INV_X1 U15314 ( .A(n13305), .ZN(n13306) );
  OAI21_X1 U15315 ( .B1(n13022), .B2(n13370), .A(n13306), .ZN(P2_U3529) );
  AOI21_X1 U15316 ( .B1(n13308), .B2(n14891), .A(n13307), .ZN(n13309) );
  OAI211_X1 U15317 ( .C1(n14851), .C2(n13311), .A(n13310), .B(n13309), .ZN(
        n13397) );
  MUX2_X1 U15318 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13397), .S(n14912), .Z(
        P2_U3528) );
  MUX2_X1 U15319 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13398), .S(n14912), .Z(
        P2_U3527) );
  INV_X1 U15320 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n13319) );
  MUX2_X1 U15321 ( .A(n13319), .B(n13399), .S(n14912), .Z(n13320) );
  OAI21_X1 U15322 ( .B1(n13402), .B2(n13370), .A(n13320), .ZN(P2_U3526) );
  AOI21_X1 U15323 ( .B1(n13322), .B2(n14891), .A(n13321), .ZN(n13323) );
  OAI211_X1 U15324 ( .C1(n13325), .C2(n14851), .A(n13324), .B(n13323), .ZN(
        n13403) );
  MUX2_X1 U15325 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13403), .S(n14912), .Z(
        P2_U3525) );
  AOI21_X1 U15326 ( .B1(n13327), .B2(n14891), .A(n13326), .ZN(n13329) );
  OAI211_X1 U15327 ( .C1(n14851), .C2(n13330), .A(n13329), .B(n13328), .ZN(
        n13404) );
  MUX2_X1 U15328 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13404), .S(n14912), .Z(
        P2_U3524) );
  OAI211_X1 U15329 ( .C1(n14851), .C2(n13333), .A(n13332), .B(n13331), .ZN(
        n13334) );
  INV_X1 U15330 ( .A(n13334), .ZN(n13405) );
  MUX2_X1 U15331 ( .A(n15208), .B(n13405), .S(n14912), .Z(n13335) );
  OAI21_X1 U15332 ( .B1(n13408), .B2(n13370), .A(n13335), .ZN(P2_U3523) );
  NAND2_X1 U15333 ( .A1(n13336), .A2(n14880), .ZN(n13338) );
  NAND3_X1 U15334 ( .A1(n13339), .A2(n13338), .A3(n13337), .ZN(n13409) );
  MUX2_X1 U15335 ( .A(n13409), .B(P2_REG1_REG_23__SCAN_IN), .S(n14910), .Z(
        n13340) );
  INV_X1 U15336 ( .A(n13340), .ZN(n13341) );
  OAI21_X1 U15337 ( .B1(n13412), .B2(n13370), .A(n13341), .ZN(P2_U3522) );
  INV_X1 U15338 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n13346) );
  INV_X1 U15339 ( .A(n13342), .ZN(n13345) );
  AOI211_X1 U15340 ( .C1(n13345), .C2(n14880), .A(n13344), .B(n13343), .ZN(
        n13413) );
  MUX2_X1 U15341 ( .A(n13346), .B(n13413), .S(n14912), .Z(n13347) );
  OAI21_X1 U15342 ( .B1(n13416), .B2(n13370), .A(n13347), .ZN(P2_U3521) );
  AOI211_X1 U15343 ( .C1(n14880), .C2(n13350), .A(n13349), .B(n13348), .ZN(
        n13417) );
  MUX2_X1 U15344 ( .A(n15128), .B(n13417), .S(n14912), .Z(n13351) );
  OAI21_X1 U15345 ( .B1(n13420), .B2(n13370), .A(n13351), .ZN(P2_U3520) );
  AOI21_X1 U15346 ( .B1(n13353), .B2(n14891), .A(n13352), .ZN(n13354) );
  OAI211_X1 U15347 ( .C1(n14851), .C2(n13356), .A(n13355), .B(n13354), .ZN(
        n13421) );
  MUX2_X1 U15348 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13421), .S(n14912), .Z(
        P2_U3519) );
  AOI211_X1 U15349 ( .C1(n13359), .C2(n14873), .A(n13358), .B(n13357), .ZN(
        n13422) );
  MUX2_X1 U15350 ( .A(n15252), .B(n13422), .S(n14912), .Z(n13360) );
  OAI21_X1 U15351 ( .B1(n13425), .B2(n13370), .A(n13360), .ZN(P2_U3518) );
  AOI211_X1 U15352 ( .C1(n14880), .C2(n13363), .A(n13362), .B(n13361), .ZN(
        n13426) );
  MUX2_X1 U15353 ( .A(n14815), .B(n13426), .S(n14912), .Z(n13364) );
  OAI21_X1 U15354 ( .B1(n13429), .B2(n13370), .A(n13364), .ZN(P2_U3517) );
  INV_X1 U15355 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13368) );
  AOI211_X1 U15356 ( .C1(n13367), .C2(n14880), .A(n13366), .B(n13365), .ZN(
        n13430) );
  MUX2_X1 U15357 ( .A(n13368), .B(n13430), .S(n14912), .Z(n13369) );
  OAI21_X1 U15358 ( .B1(n7041), .B2(n13370), .A(n13369), .ZN(P2_U3516) );
  AOI21_X1 U15359 ( .B1(n13372), .B2(n14891), .A(n13371), .ZN(n13374) );
  OAI211_X1 U15360 ( .C1(n14851), .C2(n13375), .A(n13374), .B(n13373), .ZN(
        n13433) );
  MUX2_X1 U15361 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13433), .S(n14912), .Z(
        P2_U3515) );
  AOI211_X1 U15362 ( .C1(n14880), .C2(n13378), .A(n13377), .B(n13376), .ZN(
        n13437) );
  AOI22_X1 U15363 ( .A1(n13435), .A2(n13379), .B1(P2_REG1_REG_15__SCAN_IN), 
        .B2(n14910), .ZN(n13380) );
  OAI21_X1 U15364 ( .B1(n13437), .B2(n14910), .A(n13380), .ZN(P2_U3514) );
  AOI21_X1 U15365 ( .B1(n14380), .B2(n14891), .A(n13381), .ZN(n13383) );
  OAI211_X1 U15366 ( .C1(n14851), .C2(n13384), .A(n13383), .B(n13382), .ZN(
        n13438) );
  MUX2_X1 U15367 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13438), .S(n14912), .Z(
        P2_U3513) );
  AOI21_X1 U15368 ( .B1(n13386), .B2(n14891), .A(n13385), .ZN(n13387) );
  OAI211_X1 U15369 ( .C1(n13389), .C2(n14851), .A(n13388), .B(n13387), .ZN(
        n13439) );
  MUX2_X1 U15370 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13439), .S(n14912), .Z(
        P2_U3512) );
  INV_X1 U15371 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n13391) );
  MUX2_X1 U15372 ( .A(n13391), .B(n13390), .S(n15282), .Z(n13392) );
  OAI21_X1 U15373 ( .B1(n13393), .B2(n13432), .A(n13392), .ZN(P2_U3498) );
  MUX2_X1 U15374 ( .A(n13394), .B(P2_REG0_REG_30__SCAN_IN), .S(n14899), .Z(
        n13395) );
  INV_X1 U15375 ( .A(n13395), .ZN(n13396) );
  OAI21_X1 U15376 ( .B1(n13022), .B2(n13432), .A(n13396), .ZN(P2_U3497) );
  MUX2_X1 U15377 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13397), .S(n15282), .Z(
        P2_U3496) );
  MUX2_X1 U15378 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13398), .S(n15282), .Z(
        P2_U3495) );
  INV_X1 U15379 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n13400) );
  MUX2_X1 U15380 ( .A(n13400), .B(n13399), .S(n15282), .Z(n13401) );
  OAI21_X1 U15381 ( .B1(n13402), .B2(n13432), .A(n13401), .ZN(P2_U3494) );
  MUX2_X1 U15382 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13403), .S(n15282), .Z(
        P2_U3493) );
  MUX2_X1 U15383 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13404), .S(n15282), .Z(
        P2_U3492) );
  INV_X1 U15384 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n13406) );
  MUX2_X1 U15385 ( .A(n13406), .B(n13405), .S(n15282), .Z(n13407) );
  OAI21_X1 U15386 ( .B1(n13408), .B2(n13432), .A(n13407), .ZN(P2_U3491) );
  MUX2_X1 U15387 ( .A(n13409), .B(P2_REG0_REG_23__SCAN_IN), .S(n14899), .Z(
        n13410) );
  INV_X1 U15388 ( .A(n13410), .ZN(n13411) );
  OAI21_X1 U15389 ( .B1(n13412), .B2(n13432), .A(n13411), .ZN(P2_U3490) );
  INV_X1 U15390 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n13414) );
  MUX2_X1 U15391 ( .A(n13414), .B(n13413), .S(n15282), .Z(n13415) );
  OAI21_X1 U15392 ( .B1(n13416), .B2(n13432), .A(n13415), .ZN(P2_U3489) );
  INV_X1 U15393 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n13418) );
  MUX2_X1 U15394 ( .A(n13418), .B(n13417), .S(n15282), .Z(n13419) );
  OAI21_X1 U15395 ( .B1(n13420), .B2(n13432), .A(n13419), .ZN(P2_U3488) );
  MUX2_X1 U15396 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13421), .S(n15282), .Z(
        P2_U3487) );
  INV_X1 U15397 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n13423) );
  MUX2_X1 U15398 ( .A(n13423), .B(n13422), .S(n15282), .Z(n13424) );
  OAI21_X1 U15399 ( .B1(n13425), .B2(n13432), .A(n13424), .ZN(P2_U3486) );
  INV_X1 U15400 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n13427) );
  MUX2_X1 U15401 ( .A(n13427), .B(n13426), .S(n15282), .Z(n13428) );
  OAI21_X1 U15402 ( .B1(n13429), .B2(n13432), .A(n13428), .ZN(P2_U3484) );
  MUX2_X1 U15403 ( .A(n15133), .B(n13430), .S(n15282), .Z(n13431) );
  OAI21_X1 U15404 ( .B1(n7041), .B2(n13432), .A(n13431), .ZN(P2_U3481) );
  MUX2_X1 U15405 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13433), .S(n15282), .Z(
        P2_U3478) );
  AOI22_X1 U15406 ( .A1(n13435), .A2(n13434), .B1(P2_REG0_REG_15__SCAN_IN), 
        .B2(n14899), .ZN(n13436) );
  OAI21_X1 U15407 ( .B1(n13437), .B2(n14899), .A(n13436), .ZN(P2_U3475) );
  MUX2_X1 U15408 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13438), .S(n15282), .Z(
        P2_U3472) );
  MUX2_X1 U15409 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13439), .S(n15282), .Z(
        P2_U3469) );
  INV_X1 U15410 ( .A(n13440), .ZN(n14153) );
  NAND3_X1 U15411 ( .A1(n13442), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n13444) );
  OAI22_X1 U15412 ( .A1(n13441), .A2(n13444), .B1(n13443), .B2(n13464), .ZN(
        n13445) );
  INV_X1 U15413 ( .A(n13445), .ZN(n13446) );
  OAI21_X1 U15414 ( .B1(n14153), .B2(n13459), .A(n13446), .ZN(P2_U3296) );
  INV_X1 U15415 ( .A(n13447), .ZN(n14154) );
  OAI222_X1 U15416 ( .A1(n13459), .A2(n14154), .B1(n13449), .B2(P2_U3088), 
        .C1(n13448), .C2(n13464), .ZN(P2_U3298) );
  NAND2_X1 U15417 ( .A1(n14156), .A2(n13450), .ZN(n13452) );
  OAI211_X1 U15418 ( .C1(n13464), .C2(n13453), .A(n13452), .B(n13451), .ZN(
        P2_U3299) );
  INV_X1 U15419 ( .A(n8225), .ZN(n14161) );
  OAI222_X1 U15420 ( .A1(n13464), .A2(n13455), .B1(n13459), .B2(n14161), .C1(
        P2_U3088), .C2(n13454), .ZN(P2_U3300) );
  INV_X1 U15421 ( .A(n13456), .ZN(n14165) );
  OAI222_X1 U15422 ( .A1(n13459), .A2(n14165), .B1(P2_U3088), .B2(n13458), 
        .C1(n13457), .C2(n13464), .ZN(P2_U3301) );
  INV_X1 U15423 ( .A(n13460), .ZN(n14170) );
  INV_X1 U15424 ( .A(n13461), .ZN(n13462) );
  OAI222_X1 U15425 ( .A1(n13464), .A2(n13463), .B1(n13459), .B2(n14170), .C1(
        n13462), .C2(P2_U3088), .ZN(P2_U3302) );
  MUX2_X1 U15426 ( .A(n13465), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15427 ( .A1(n14066), .A2(n13587), .ZN(n13467) );
  NAND2_X1 U15428 ( .A1(n13756), .A2(n13555), .ZN(n13466) );
  NAND2_X1 U15429 ( .A1(n13467), .A2(n13466), .ZN(n13468) );
  XNOR2_X1 U15430 ( .A(n13468), .B(n13625), .ZN(n13472) );
  NAND2_X1 U15431 ( .A1(n14066), .A2(n10153), .ZN(n13470) );
  NAND2_X1 U15432 ( .A1(n13756), .A2(n10463), .ZN(n13469) );
  NAND2_X1 U15433 ( .A1(n13470), .A2(n13469), .ZN(n13471) );
  NOR2_X1 U15434 ( .A1(n13472), .A2(n13471), .ZN(n13624) );
  AOI21_X1 U15435 ( .B1(n13472), .B2(n13471), .A(n13624), .ZN(n13597) );
  NAND2_X1 U15436 ( .A1(n14087), .A2(n13587), .ZN(n13474) );
  NAND2_X1 U15437 ( .A1(n13759), .A2(n10153), .ZN(n13473) );
  NAND2_X1 U15438 ( .A1(n13474), .A2(n13473), .ZN(n13475) );
  XNOR2_X1 U15439 ( .A(n13475), .B(n13561), .ZN(n13571) );
  AND2_X1 U15440 ( .A1(n13759), .A2(n10463), .ZN(n13476) );
  AOI21_X1 U15441 ( .B1(n14087), .B2(n6460), .A(n13476), .ZN(n13572) );
  NAND2_X1 U15442 ( .A1(n13571), .A2(n13572), .ZN(n13576) );
  INV_X1 U15443 ( .A(n13576), .ZN(n13649) );
  NAND2_X1 U15444 ( .A1(n14093), .A2(n13587), .ZN(n13478) );
  NAND2_X1 U15445 ( .A1(n13760), .A2(n10153), .ZN(n13477) );
  NAND2_X1 U15446 ( .A1(n13478), .A2(n13477), .ZN(n13479) );
  XNOR2_X1 U15447 ( .A(n13479), .B(n13561), .ZN(n13481) );
  AND2_X1 U15448 ( .A1(n13760), .A2(n10463), .ZN(n13480) );
  AOI21_X1 U15449 ( .B1(n14093), .B2(n6460), .A(n13480), .ZN(n13482) );
  NAND2_X1 U15450 ( .A1(n13481), .A2(n13482), .ZN(n13680) );
  INV_X1 U15451 ( .A(n13481), .ZN(n13484) );
  INV_X1 U15452 ( .A(n13482), .ZN(n13483) );
  NAND2_X1 U15453 ( .A1(n13484), .A2(n13483), .ZN(n13485) );
  AND2_X1 U15454 ( .A1(n13680), .A2(n13485), .ZN(n13607) );
  INV_X1 U15455 ( .A(n13488), .ZN(n13489) );
  NAND2_X1 U15456 ( .A1(n13490), .A2(n13489), .ZN(n13491) );
  NAND2_X1 U15457 ( .A1(n14414), .A2(n13587), .ZN(n13493) );
  NAND2_X1 U15458 ( .A1(n13769), .A2(n13555), .ZN(n13492) );
  NAND2_X1 U15459 ( .A1(n13493), .A2(n13492), .ZN(n13494) );
  XNOR2_X1 U15460 ( .A(n13494), .B(n13561), .ZN(n13497) );
  NOR2_X1 U15461 ( .A1(n13495), .A2(n11011), .ZN(n13496) );
  AOI21_X1 U15462 ( .B1(n14414), .B2(n6460), .A(n13496), .ZN(n13498) );
  NAND2_X1 U15463 ( .A1(n13497), .A2(n13498), .ZN(n13502) );
  INV_X1 U15464 ( .A(n13497), .ZN(n13500) );
  INV_X1 U15465 ( .A(n13498), .ZN(n13499) );
  NAND2_X1 U15466 ( .A1(n13500), .A2(n13499), .ZN(n13501) );
  NAND2_X1 U15467 ( .A1(n13502), .A2(n13501), .ZN(n14391) );
  NAND2_X1 U15468 ( .A1(n14439), .A2(n13587), .ZN(n13504) );
  OR2_X1 U15469 ( .A1(n14386), .A2(n13627), .ZN(n13503) );
  NAND2_X1 U15470 ( .A1(n13504), .A2(n13503), .ZN(n13505) );
  XNOR2_X1 U15471 ( .A(n13505), .B(n13561), .ZN(n13507) );
  NOR2_X1 U15472 ( .A1(n14386), .A2(n11011), .ZN(n13506) );
  AOI21_X1 U15473 ( .B1(n14439), .B2(n13555), .A(n13506), .ZN(n13743) );
  OR2_X1 U15474 ( .A1(n13508), .A2(n13507), .ZN(n13509) );
  NAND2_X1 U15475 ( .A1(n14430), .A2(n13587), .ZN(n13511) );
  NAND2_X1 U15476 ( .A1(n13767), .A2(n6460), .ZN(n13510) );
  NAND2_X1 U15477 ( .A1(n13511), .A2(n13510), .ZN(n13512) );
  XNOR2_X1 U15478 ( .A(n13512), .B(n13561), .ZN(n13514) );
  AND2_X1 U15479 ( .A1(n13767), .A2(n10463), .ZN(n13513) );
  AOI21_X1 U15480 ( .B1(n14430), .B2(n13555), .A(n13513), .ZN(n13515) );
  NAND2_X1 U15481 ( .A1(n13514), .A2(n13515), .ZN(n13673) );
  INV_X1 U15482 ( .A(n13514), .ZN(n13517) );
  INV_X1 U15483 ( .A(n13515), .ZN(n13516) );
  NAND2_X1 U15484 ( .A1(n13517), .A2(n13516), .ZN(n13518) );
  NAND2_X1 U15485 ( .A1(n13673), .A2(n13518), .ZN(n13663) );
  NAND2_X1 U15486 ( .A1(n14423), .A2(n13587), .ZN(n13520) );
  NAND2_X1 U15487 ( .A1(n13766), .A2(n6460), .ZN(n13519) );
  NAND2_X1 U15488 ( .A1(n13520), .A2(n13519), .ZN(n13521) );
  XNOR2_X1 U15489 ( .A(n13521), .B(n13561), .ZN(n13523) );
  AND2_X1 U15490 ( .A1(n13766), .A2(n10463), .ZN(n13522) );
  AOI21_X1 U15491 ( .B1(n14423), .B2(n13555), .A(n13522), .ZN(n13524) );
  NAND2_X1 U15492 ( .A1(n13523), .A2(n13524), .ZN(n13528) );
  INV_X1 U15493 ( .A(n13523), .ZN(n13526) );
  INV_X1 U15494 ( .A(n13524), .ZN(n13525) );
  NAND2_X1 U15495 ( .A1(n13526), .A2(n13525), .ZN(n13527) );
  AND2_X1 U15496 ( .A1(n13528), .A2(n13527), .ZN(n13671) );
  OAI22_X1 U15497 ( .A1(n14044), .A2(n13629), .B1(n13530), .B2(n13627), .ZN(
        n13529) );
  XNOR2_X1 U15498 ( .A(n13529), .B(n13561), .ZN(n13537) );
  OAI22_X1 U15499 ( .A1(n14044), .A2(n13627), .B1(n13530), .B2(n11011), .ZN(
        n13535) );
  XNOR2_X1 U15500 ( .A(n13537), .B(n13535), .ZN(n13709) );
  NAND2_X1 U15501 ( .A1(n14027), .A2(n13587), .ZN(n13532) );
  NAND2_X1 U15502 ( .A1(n13764), .A2(n6460), .ZN(n13531) );
  NAND2_X1 U15503 ( .A1(n13532), .A2(n13531), .ZN(n13533) );
  XNOR2_X1 U15504 ( .A(n13533), .B(n13625), .ZN(n13541) );
  NOR2_X1 U15505 ( .A1(n13711), .A2(n11011), .ZN(n13534) );
  AOI21_X1 U15506 ( .B1(n14027), .B2(n13555), .A(n13534), .ZN(n13539) );
  XNOR2_X1 U15507 ( .A(n13541), .B(n13539), .ZN(n13618) );
  INV_X1 U15508 ( .A(n13535), .ZN(n13536) );
  NAND2_X1 U15509 ( .A1(n13537), .A2(n13536), .ZN(n13616) );
  AND2_X1 U15510 ( .A1(n13618), .A2(n13616), .ZN(n13538) );
  NAND2_X1 U15511 ( .A1(n13707), .A2(n13538), .ZN(n13617) );
  INV_X1 U15512 ( .A(n13539), .ZN(n13540) );
  NAND2_X1 U15513 ( .A1(n13541), .A2(n13540), .ZN(n13542) );
  NAND2_X1 U15514 ( .A1(n14113), .A2(n13587), .ZN(n13544) );
  NAND2_X1 U15515 ( .A1(n13763), .A2(n13555), .ZN(n13543) );
  NAND2_X1 U15516 ( .A1(n13544), .A2(n13543), .ZN(n13545) );
  XNOR2_X1 U15517 ( .A(n13545), .B(n13625), .ZN(n13549) );
  AND2_X1 U15518 ( .A1(n13763), .A2(n10463), .ZN(n13546) );
  AOI21_X1 U15519 ( .B1(n14113), .B2(n13555), .A(n13546), .ZN(n13547) );
  XNOR2_X1 U15520 ( .A(n13549), .B(n13547), .ZN(n13692) );
  INV_X1 U15521 ( .A(n13547), .ZN(n13548) );
  NAND2_X1 U15522 ( .A1(n13549), .A2(n13548), .ZN(n13550) );
  NAND2_X1 U15523 ( .A1(n14108), .A2(n13587), .ZN(n13552) );
  NAND2_X1 U15524 ( .A1(n13762), .A2(n13555), .ZN(n13551) );
  NAND2_X1 U15525 ( .A1(n13552), .A2(n13551), .ZN(n13553) );
  XNOR2_X1 U15526 ( .A(n13553), .B(n13561), .ZN(n13556) );
  AND2_X1 U15527 ( .A1(n13762), .A2(n10463), .ZN(n13554) );
  AOI21_X1 U15528 ( .B1(n14108), .B2(n13555), .A(n13554), .ZN(n13557) );
  NAND2_X1 U15529 ( .A1(n13556), .A2(n13557), .ZN(n13699) );
  INV_X1 U15530 ( .A(n13556), .ZN(n13559) );
  INV_X1 U15531 ( .A(n13557), .ZN(n13558) );
  NAND2_X1 U15532 ( .A1(n13559), .A2(n13558), .ZN(n13560) );
  NAND2_X1 U15533 ( .A1(n13699), .A2(n13560), .ZN(n13640) );
  OAI22_X1 U15534 ( .A1(n14101), .A2(n13629), .B1(n13642), .B2(n13627), .ZN(
        n13562) );
  XNOR2_X1 U15535 ( .A(n13562), .B(n13561), .ZN(n13566) );
  OR2_X1 U15536 ( .A1(n14101), .A2(n13627), .ZN(n13564) );
  NAND2_X1 U15537 ( .A1(n13761), .A2(n10463), .ZN(n13563) );
  NAND2_X1 U15538 ( .A1(n13564), .A2(n13563), .ZN(n13567) );
  INV_X1 U15539 ( .A(n13567), .ZN(n13565) );
  NAND2_X1 U15540 ( .A1(n13566), .A2(n13565), .ZN(n13605) );
  INV_X1 U15541 ( .A(n13566), .ZN(n13568) );
  NAND2_X1 U15542 ( .A1(n13568), .A2(n13567), .ZN(n13569) );
  AND2_X1 U15543 ( .A1(n13605), .A2(n13569), .ZN(n13700) );
  NAND2_X1 U15544 ( .A1(n13607), .A2(n13570), .ZN(n13608) );
  INV_X1 U15545 ( .A(n13571), .ZN(n13574) );
  INV_X1 U15546 ( .A(n13572), .ZN(n13573) );
  NAND2_X1 U15547 ( .A1(n13574), .A2(n13573), .ZN(n13575) );
  AND2_X1 U15548 ( .A1(n13576), .A2(n13575), .ZN(n13683) );
  NAND2_X1 U15549 ( .A1(n14082), .A2(n13587), .ZN(n13579) );
  NAND2_X1 U15550 ( .A1(n13758), .A2(n10153), .ZN(n13578) );
  NAND2_X1 U15551 ( .A1(n13579), .A2(n13578), .ZN(n13580) );
  XNOR2_X1 U15552 ( .A(n13580), .B(n13625), .ZN(n13584) );
  NAND2_X1 U15553 ( .A1(n14082), .A2(n10153), .ZN(n13582) );
  NAND2_X1 U15554 ( .A1(n13758), .A2(n10463), .ZN(n13581) );
  NAND2_X1 U15555 ( .A1(n13582), .A2(n13581), .ZN(n13583) );
  NOR2_X1 U15556 ( .A1(n13584), .A2(n13583), .ZN(n13585) );
  AOI21_X1 U15557 ( .B1(n13584), .B2(n13583), .A(n13585), .ZN(n13650) );
  OAI21_X1 U15558 ( .B1(n13649), .B2(n13684), .A(n13650), .ZN(n13651) );
  INV_X1 U15559 ( .A(n13585), .ZN(n13586) );
  NAND2_X1 U15560 ( .A1(n13651), .A2(n13586), .ZN(n13729) );
  NAND2_X1 U15561 ( .A1(n13915), .A2(n13587), .ZN(n13589) );
  NAND2_X1 U15562 ( .A1(n13757), .A2(n10153), .ZN(n13588) );
  NAND2_X1 U15563 ( .A1(n13589), .A2(n13588), .ZN(n13590) );
  XNOR2_X1 U15564 ( .A(n13590), .B(n13625), .ZN(n13594) );
  NAND2_X1 U15565 ( .A1(n13915), .A2(n13555), .ZN(n13592) );
  NAND2_X1 U15566 ( .A1(n13757), .A2(n10463), .ZN(n13591) );
  NAND2_X1 U15567 ( .A1(n13592), .A2(n13591), .ZN(n13593) );
  NOR2_X1 U15568 ( .A1(n13594), .A2(n13593), .ZN(n13595) );
  AOI21_X1 U15569 ( .B1(n13594), .B2(n13593), .A(n13595), .ZN(n13730) );
  INV_X1 U15570 ( .A(n13595), .ZN(n13596) );
  NAND2_X1 U15571 ( .A1(n13598), .A2(n14395), .ZN(n13603) );
  OAI22_X1 U15572 ( .A1(n13628), .A2(n14385), .B1(n13599), .B2(n14633), .ZN(
        n13897) );
  AOI22_X1 U15573 ( .A1(n13897), .A2(n14397), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13602) );
  NAND2_X1 U15574 ( .A1(n14066), .A2(n14398), .ZN(n13601) );
  NAND2_X1 U15575 ( .A1(n13739), .A2(n13902), .ZN(n13600) );
  NAND4_X1 U15576 ( .A1(n13603), .A2(n13602), .A3(n13601), .A4(n13600), .ZN(
        P1_U3214) );
  INV_X1 U15577 ( .A(n14093), .ZN(n13964) );
  INV_X1 U15578 ( .A(n13604), .ZN(n13701) );
  INV_X1 U15579 ( .A(n13605), .ZN(n13606) );
  NOR3_X1 U15580 ( .A1(n13701), .A2(n13607), .A3(n13606), .ZN(n13609) );
  INV_X1 U15581 ( .A(n13608), .ZN(n13682) );
  OAI21_X1 U15582 ( .B1(n13609), .B2(n13682), .A(n14395), .ZN(n13615) );
  NAND2_X1 U15583 ( .A1(n13761), .A2(n14387), .ZN(n13611) );
  NAND2_X1 U15584 ( .A1(n13759), .A2(n13732), .ZN(n13610) );
  AND2_X1 U15585 ( .A1(n13611), .A2(n13610), .ZN(n13960) );
  OAI22_X1 U15586 ( .A1(n13737), .A2(n13960), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13612), .ZN(n13613) );
  AOI21_X1 U15587 ( .B1(n13961), .B2(n13739), .A(n13613), .ZN(n13614) );
  OAI211_X1 U15588 ( .C1(n13964), .C2(n13742), .A(n13615), .B(n13614), .ZN(
        P1_U3216) );
  INV_X1 U15589 ( .A(n14027), .ZN(n14123) );
  AND2_X1 U15590 ( .A1(n13707), .A2(n13616), .ZN(n13619) );
  OAI211_X1 U15591 ( .C1(n13619), .C2(n13618), .A(n14395), .B(n13617), .ZN(
        n13623) );
  INV_X1 U15592 ( .A(n13620), .ZN(n14026) );
  AOI22_X1 U15593 ( .A1(n13763), .A2(n13732), .B1(n14387), .B2(n13765), .ZN(
        n14121) );
  NAND2_X1 U15594 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13861)
         );
  OAI21_X1 U15595 ( .B1(n14121), .B2(n13737), .A(n13861), .ZN(n13621) );
  AOI21_X1 U15596 ( .B1(n14026), .B2(n13739), .A(n13621), .ZN(n13622) );
  OAI211_X1 U15597 ( .C1(n14123), .C2(n13742), .A(n13623), .B(n13622), .ZN(
        P1_U3219) );
  OAI22_X1 U15598 ( .A1(n6960), .A2(n13627), .B1(n13628), .B2(n11011), .ZN(
        n13626) );
  XNOR2_X1 U15599 ( .A(n13626), .B(n13625), .ZN(n13631) );
  OAI22_X1 U15600 ( .A1(n6960), .A2(n13629), .B1(n13628), .B2(n13627), .ZN(
        n13630) );
  XNOR2_X1 U15601 ( .A(n13631), .B(n13630), .ZN(n13632) );
  INV_X1 U15602 ( .A(n13633), .ZN(n13886) );
  OAI22_X1 U15603 ( .A1(n13635), .A2(n14385), .B1(n13634), .B2(n14633), .ZN(
        n13880) );
  AOI22_X1 U15604 ( .A1(n13880), .A2(n14397), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13636) );
  OAI21_X1 U15605 ( .B1(n13886), .B2(n14401), .A(n13636), .ZN(n13637) );
  AOI21_X1 U15606 ( .B1(n14061), .B2(n14398), .A(n13637), .ZN(n13638) );
  OAI21_X1 U15607 ( .B1(n13639), .B2(n13751), .A(n13638), .ZN(P1_U3220) );
  AOI21_X1 U15608 ( .B1(n13641), .B2(n13640), .A(n6502), .ZN(n13648) );
  INV_X1 U15609 ( .A(n13989), .ZN(n13645) );
  OAI22_X1 U15610 ( .A1(n13643), .A2(n14633), .B1(n13642), .B2(n14385), .ZN(
        n14107) );
  AOI22_X1 U15611 ( .A1(n14107), .A2(n14397), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13644) );
  OAI21_X1 U15612 ( .B1(n13645), .B2(n14401), .A(n13644), .ZN(n13646) );
  AOI21_X1 U15613 ( .B1(n14108), .B2(n14398), .A(n13646), .ZN(n13647) );
  OAI21_X1 U15614 ( .B1(n13648), .B2(n13751), .A(n13647), .ZN(P1_U3223) );
  NOR3_X1 U15615 ( .A1(n13650), .A2(n13649), .A3(n13684), .ZN(n13653) );
  INV_X1 U15616 ( .A(n13651), .ZN(n13652) );
  OAI21_X1 U15617 ( .B1(n13653), .B2(n13652), .A(n14395), .ZN(n13659) );
  NAND2_X1 U15618 ( .A1(n13759), .A2(n14387), .ZN(n13655) );
  NAND2_X1 U15619 ( .A1(n13757), .A2(n13732), .ZN(n13654) );
  NAND2_X1 U15620 ( .A1(n13655), .A2(n13654), .ZN(n14081) );
  INV_X1 U15621 ( .A(n14081), .ZN(n13933) );
  OAI22_X1 U15622 ( .A1(n13737), .A2(n13933), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13656), .ZN(n13657) );
  AOI21_X1 U15623 ( .B1(n13931), .B2(n13739), .A(n13657), .ZN(n13658) );
  OAI211_X1 U15624 ( .C1(n13660), .C2(n13742), .A(n13659), .B(n13658), .ZN(
        P1_U3225) );
  INV_X1 U15625 ( .A(n13674), .ZN(n13661) );
  AOI21_X1 U15626 ( .B1(n13663), .B2(n13662), .A(n13661), .ZN(n13668) );
  NAND2_X1 U15627 ( .A1(n14429), .A2(n14397), .ZN(n13664) );
  NAND2_X1 U15628 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14551)
         );
  OAI211_X1 U15629 ( .C1(n14401), .C2(n13665), .A(n13664), .B(n14551), .ZN(
        n13666) );
  AOI21_X1 U15630 ( .B1(n14430), .B2(n14398), .A(n13666), .ZN(n13667) );
  OAI21_X1 U15631 ( .B1(n13668), .B2(n13751), .A(n13667), .ZN(P1_U3226) );
  NAND2_X1 U15632 ( .A1(n14422), .A2(n14397), .ZN(n13669) );
  NAND2_X1 U15633 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14568)
         );
  OAI211_X1 U15634 ( .C1(n14401), .C2(n13670), .A(n13669), .B(n14568), .ZN(
        n13678) );
  INV_X1 U15635 ( .A(n13671), .ZN(n13672) );
  NAND3_X1 U15636 ( .A1(n13674), .A2(n13673), .A3(n13672), .ZN(n13675) );
  AOI21_X1 U15637 ( .B1(n13676), .B2(n13675), .A(n13751), .ZN(n13677) );
  AOI211_X1 U15638 ( .C1(n14423), .C2(n14398), .A(n13678), .B(n13677), .ZN(
        n13679) );
  INV_X1 U15639 ( .A(n13679), .ZN(P1_U3228) );
  INV_X1 U15640 ( .A(n13680), .ZN(n13681) );
  NOR3_X1 U15641 ( .A1(n13683), .A2(n13682), .A3(n13681), .ZN(n13685) );
  OAI21_X1 U15642 ( .B1(n13685), .B2(n13684), .A(n14395), .ZN(n13691) );
  NAND2_X1 U15643 ( .A1(n13760), .A2(n14387), .ZN(n13687) );
  NAND2_X1 U15644 ( .A1(n13758), .A2(n13732), .ZN(n13686) );
  NAND2_X1 U15645 ( .A1(n13687), .A2(n13686), .ZN(n13943) );
  INV_X1 U15646 ( .A(n13943), .ZN(n13688) );
  OAI22_X1 U15647 ( .A1(n13737), .A2(n13688), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15248), .ZN(n13689) );
  AOI21_X1 U15648 ( .B1(n13948), .B2(n13739), .A(n13689), .ZN(n13690) );
  OAI211_X1 U15649 ( .C1(n13950), .C2(n13742), .A(n13691), .B(n13690), .ZN(
        P1_U3229) );
  XNOR2_X1 U15650 ( .A(n13693), .B(n13692), .ZN(n13698) );
  NOR2_X1 U15651 ( .A1(n14401), .A2(n14006), .ZN(n13696) );
  AOI22_X1 U15652 ( .A1(n13762), .A2(n13732), .B1(n14387), .B2(n13764), .ZN(
        n14004) );
  OAI22_X1 U15653 ( .A1(n14004), .A2(n13737), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13694), .ZN(n13695) );
  AOI211_X1 U15654 ( .C1(n14113), .C2(n14398), .A(n13696), .B(n13695), .ZN(
        n13697) );
  OAI21_X1 U15655 ( .B1(n13698), .B2(n13751), .A(n13697), .ZN(P1_U3233) );
  NOR3_X1 U15656 ( .A1(n6502), .A2(n7396), .A3(n13700), .ZN(n13702) );
  OAI21_X1 U15657 ( .B1(n13702), .B2(n13701), .A(n14395), .ZN(n13706) );
  AOI22_X1 U15658 ( .A1(n13762), .A2(n14387), .B1(n13732), .B2(n13760), .ZN(
        n14099) );
  OAI22_X1 U15659 ( .A1(n14099), .A2(n13737), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13703), .ZN(n13704) );
  AOI21_X1 U15660 ( .B1(n13975), .B2(n13739), .A(n13704), .ZN(n13705) );
  OAI211_X1 U15661 ( .C1(n13742), .C2(n14101), .A(n13706), .B(n13705), .ZN(
        P1_U3235) );
  OAI21_X1 U15662 ( .B1(n13709), .B2(n13708), .A(n13707), .ZN(n13710) );
  NAND2_X1 U15663 ( .A1(n13710), .A2(n14395), .ZN(n13715) );
  OAI22_X1 U15664 ( .A1(n13711), .A2(n14385), .B1(n7279), .B2(n14633), .ZN(
        n13712) );
  INV_X1 U15665 ( .A(n13712), .ZN(n14036) );
  NAND2_X1 U15666 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14583)
         );
  OAI21_X1 U15667 ( .B1(n14036), .B2(n13737), .A(n14583), .ZN(n13713) );
  AOI21_X1 U15668 ( .B1(n14041), .B2(n13739), .A(n13713), .ZN(n13714) );
  OAI211_X1 U15669 ( .C1(n14044), .C2(n13742), .A(n13715), .B(n13714), .ZN(
        P1_U3238) );
  AND2_X1 U15670 ( .A1(n13717), .A2(n13716), .ZN(n13720) );
  OAI211_X1 U15671 ( .C1(n13720), .C2(n13719), .A(n14395), .B(n13718), .ZN(
        n13727) );
  NAND2_X1 U15672 ( .A1(n13777), .A2(n14387), .ZN(n13722) );
  NAND2_X1 U15673 ( .A1(n13775), .A2(n13732), .ZN(n13721) );
  NAND2_X1 U15674 ( .A1(n13722), .A2(n13721), .ZN(n14593) );
  AOI22_X1 U15675 ( .A1(n14397), .A2(n14593), .B1(P1_REG3_REG_6__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13726) );
  NAND2_X1 U15676 ( .A1(n14398), .A2(n13723), .ZN(n13725) );
  OR2_X1 U15677 ( .A1(n14401), .A2(n14594), .ZN(n13724) );
  NAND4_X1 U15678 ( .A1(n13727), .A2(n13726), .A3(n13725), .A4(n13724), .ZN(
        P1_U3239) );
  OAI21_X1 U15679 ( .B1(n13730), .B2(n13729), .A(n13728), .ZN(n13731) );
  NAND2_X1 U15680 ( .A1(n13731), .A2(n14395), .ZN(n13741) );
  NAND2_X1 U15681 ( .A1(n13756), .A2(n13732), .ZN(n13734) );
  NAND2_X1 U15682 ( .A1(n13758), .A2(n14387), .ZN(n13733) );
  NAND2_X1 U15683 ( .A1(n13734), .A2(n13733), .ZN(n14071) );
  INV_X1 U15684 ( .A(n14071), .ZN(n13736) );
  OAI22_X1 U15685 ( .A1(n13737), .A2(n13736), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13735), .ZN(n13738) );
  AOI21_X1 U15686 ( .B1(n13916), .B2(n13739), .A(n13738), .ZN(n13740) );
  OAI211_X1 U15687 ( .C1(n14070), .C2(n13742), .A(n13741), .B(n13740), .ZN(
        P1_U3240) );
  XNOR2_X1 U15688 ( .A(n13744), .B(n13743), .ZN(n13752) );
  INV_X1 U15689 ( .A(n13745), .ZN(n13748) );
  AOI21_X1 U15690 ( .B1(n14397), .B2(n14438), .A(n13746), .ZN(n13747) );
  OAI21_X1 U15691 ( .B1(n13748), .B2(n14401), .A(n13747), .ZN(n13749) );
  AOI21_X1 U15692 ( .B1(n14439), .B2(n14398), .A(n13749), .ZN(n13750) );
  OAI21_X1 U15693 ( .B1(n13752), .B2(n13751), .A(n13750), .ZN(P1_U3241) );
  MUX2_X1 U15694 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n13864), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15695 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13753), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15696 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13754), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15697 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13755), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15698 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13756), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15699 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13757), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15700 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n13758), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15701 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13759), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15702 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13760), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15703 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n13761), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15704 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13762), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15705 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13763), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15706 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13764), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15707 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13765), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15708 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13766), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15709 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13767), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15710 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13768), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15711 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13769), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15712 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14388), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15713 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13770), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15714 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13771), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15715 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13772), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15716 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13773), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15717 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13774), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15718 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13775), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15719 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13776), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15720 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13777), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15721 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13778), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15722 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13779), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15723 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13780), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15724 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14629), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15725 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n10017), .S(P1_U4016), .Z(
        P1_U3560) );
  MUX2_X1 U15726 ( .A(n13782), .B(n13781), .S(n6459), .Z(n13786) );
  OAI21_X1 U15727 ( .B1(n6459), .B2(P1_REG2_REG_0__SCAN_IN), .A(n13783), .ZN(
        n14487) );
  NAND2_X1 U15728 ( .A1(n14487), .A2(n13784), .ZN(n13785) );
  OAI211_X1 U15729 ( .C1(n13786), .C2(n14159), .A(P1_U4016), .B(n13785), .ZN(
        n13824) );
  INV_X1 U15730 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n14611) );
  OAI22_X1 U15731 ( .A1(n14585), .A2(n7031), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14611), .ZN(n13787) );
  AOI21_X1 U15732 ( .B1(n13788), .B2(n14582), .A(n13787), .ZN(n13798) );
  AOI211_X1 U15733 ( .C1(n13791), .C2(n13790), .A(n13789), .B(n14572), .ZN(
        n13792) );
  INV_X1 U15734 ( .A(n13792), .ZN(n13797) );
  OAI211_X1 U15735 ( .C1(n13795), .C2(n13794), .A(n14558), .B(n13793), .ZN(
        n13796) );
  NAND4_X1 U15736 ( .A1(n13824), .A2(n13798), .A3(n13797), .A4(n13796), .ZN(
        P1_U3245) );
  AOI211_X1 U15737 ( .C1(n13801), .C2(n13800), .A(n13799), .B(n14572), .ZN(
        n13802) );
  INV_X1 U15738 ( .A(n13802), .ZN(n13811) );
  NAND2_X1 U15739 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n13803) );
  OAI21_X1 U15740 ( .B1(n14585), .B2(n14182), .A(n13803), .ZN(n13804) );
  AOI21_X1 U15741 ( .B1(n13805), .B2(n14582), .A(n13804), .ZN(n13810) );
  OAI211_X1 U15742 ( .C1(n13808), .C2(n13807), .A(n14558), .B(n13806), .ZN(
        n13809) );
  NAND3_X1 U15743 ( .A1(n13811), .A2(n13810), .A3(n13809), .ZN(P1_U3246) );
  INV_X1 U15744 ( .A(n13812), .ZN(n13817) );
  AOI211_X1 U15745 ( .C1(n13815), .C2(n13814), .A(n14572), .B(n13813), .ZN(
        n13816) );
  AOI211_X1 U15746 ( .C1(n14491), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n13817), .B(
        n13816), .ZN(n13826) );
  NOR2_X1 U15747 ( .A1(n13819), .A2(n13818), .ZN(n13820) );
  NOR2_X1 U15748 ( .A1(n13821), .A2(n13820), .ZN(n13822) );
  AOI22_X1 U15749 ( .A1(n13823), .A2(n14582), .B1(n14558), .B2(n13822), .ZN(
        n13825) );
  NAND3_X1 U15750 ( .A1(n13826), .A2(n13825), .A3(n13824), .ZN(P1_U3247) );
  NAND2_X1 U15751 ( .A1(n13827), .A2(n13840), .ZN(n13829) );
  NAND2_X1 U15752 ( .A1(n14549), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13830) );
  OAI21_X1 U15753 ( .B1(n14549), .B2(P1_REG2_REG_16__SCAN_IN), .A(n13830), 
        .ZN(n14543) );
  NAND2_X1 U15754 ( .A1(n13844), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13831) );
  NAND2_X1 U15755 ( .A1(n14542), .A2(n13831), .ZN(n14557) );
  OR2_X1 U15756 ( .A1(n13849), .A2(n13832), .ZN(n13834) );
  NAND2_X1 U15757 ( .A1(n13849), .A2(n13832), .ZN(n13833) );
  NAND2_X1 U15758 ( .A1(n13834), .A2(n13833), .ZN(n14556) );
  NAND2_X1 U15759 ( .A1(n14557), .A2(n14556), .ZN(n14555) );
  NAND2_X1 U15760 ( .A1(n13849), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13835) );
  XNOR2_X1 U15761 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13838), .ZN(n13857) );
  INV_X1 U15762 ( .A(n13857), .ZN(n13855) );
  NAND2_X1 U15763 ( .A1(n13840), .A2(n13839), .ZN(n13842) );
  NAND2_X1 U15764 ( .A1(n14549), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n13843) );
  OAI21_X1 U15765 ( .B1(n14549), .B2(P1_REG1_REG_16__SCAN_IN), .A(n13843), 
        .ZN(n14545) );
  NAND2_X1 U15766 ( .A1(n13844), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n13845) );
  NAND2_X1 U15767 ( .A1(n14544), .A2(n13845), .ZN(n14560) );
  INV_X1 U15768 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13846) );
  OR2_X1 U15769 ( .A1(n13849), .A2(n13846), .ZN(n13848) );
  NAND2_X1 U15770 ( .A1(n13849), .A2(n13846), .ZN(n13847) );
  NAND2_X1 U15771 ( .A1(n13848), .A2(n13847), .ZN(n14559) );
  NOR2_X1 U15772 ( .A1(n13851), .A2(n13850), .ZN(n13852) );
  AOI21_X1 U15773 ( .B1(n13851), .B2(n13850), .A(n13852), .ZN(n14574) );
  AND2_X1 U15774 ( .A1(n14574), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14575) );
  NOR2_X1 U15775 ( .A1(n14575), .A2(n13852), .ZN(n13853) );
  XNOR2_X1 U15776 ( .A(n13853), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n13856) );
  OAI21_X1 U15777 ( .B1(n13856), .B2(n14576), .A(n14566), .ZN(n13854) );
  AOI21_X1 U15778 ( .B1(n13855), .B2(n14554), .A(n13854), .ZN(n13860) );
  AOI22_X1 U15779 ( .A1(n13857), .A2(n14554), .B1(n14558), .B2(n13856), .ZN(
        n13859) );
  OAI211_X1 U15780 ( .C1(n7520), .C2(n14585), .A(n13862), .B(n13861), .ZN(
        P1_U3262) );
  XNOR2_X1 U15781 ( .A(n13869), .B(n13866), .ZN(n13863) );
  NAND2_X1 U15782 ( .A1(n13863), .A2(n14617), .ZN(n14047) );
  NAND2_X1 U15783 ( .A1(n13865), .A2(n13864), .ZN(n14049) );
  NOR2_X1 U15784 ( .A1(n14638), .A2(n14049), .ZN(n13875) );
  INV_X1 U15785 ( .A(n13866), .ZN(n14048) );
  NOR2_X1 U15786 ( .A1(n14048), .A2(n14640), .ZN(n13867) );
  AOI211_X1 U15787 ( .C1(n14648), .C2(P1_REG2_REG_31__SCAN_IN), .A(n13875), 
        .B(n13867), .ZN(n13868) );
  OAI21_X1 U15788 ( .B1(n14047), .B2(n14011), .A(n13868), .ZN(P1_U3263) );
  INV_X1 U15789 ( .A(n13869), .ZN(n13873) );
  NOR2_X1 U15790 ( .A1(n6956), .A2(n14640), .ZN(n13874) );
  AOI211_X1 U15791 ( .C1(n14648), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13875), 
        .B(n13874), .ZN(n13876) );
  OAI21_X1 U15792 ( .B1(n14011), .B2(n14052), .A(n13876), .ZN(P1_U3264) );
  OAI21_X1 U15793 ( .B1(n13879), .B2(n13878), .A(n13877), .ZN(n13881) );
  AOI21_X1 U15794 ( .B1(n13881), .B2(n14630), .A(n13880), .ZN(n14063) );
  OAI21_X1 U15795 ( .B1(n13884), .B2(n13883), .A(n13882), .ZN(n14064) );
  NAND2_X1 U15796 ( .A1(n14638), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n13885) );
  OAI21_X1 U15797 ( .B1(n14612), .B2(n13886), .A(n13885), .ZN(n13887) );
  AOI21_X1 U15798 ( .B1(n14061), .B2(n14409), .A(n13887), .ZN(n13890) );
  AOI21_X1 U15799 ( .B1(n14061), .B2(n13899), .A(n14675), .ZN(n13888) );
  NAND2_X1 U15800 ( .A1(n14060), .A2(n14644), .ZN(n13889) );
  OAI211_X1 U15801 ( .C1(n14064), .C2(n14016), .A(n13890), .B(n13889), .ZN(
        n13891) );
  INV_X1 U15802 ( .A(n13891), .ZN(n13892) );
  OAI21_X1 U15803 ( .B1(n14648), .B2(n14063), .A(n13892), .ZN(P1_U3265) );
  INV_X1 U15804 ( .A(n13907), .ZN(n13894) );
  NAND2_X1 U15805 ( .A1(n13894), .A2(n13893), .ZN(n13896) );
  OAI21_X1 U15806 ( .B1(n13896), .B2(n13921), .A(n13895), .ZN(n13898) );
  AOI21_X1 U15807 ( .B1(n13898), .B2(n14630), .A(n13897), .ZN(n14068) );
  INV_X1 U15808 ( .A(n13914), .ZN(n13901) );
  INV_X1 U15809 ( .A(n13899), .ZN(n13900) );
  AOI211_X1 U15810 ( .C1(n14066), .C2(n13901), .A(n14675), .B(n13900), .ZN(
        n14065) );
  AOI22_X1 U15811 ( .A1(n14638), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14637), 
        .B2(n13902), .ZN(n13903) );
  OAI21_X1 U15812 ( .B1(n13904), .B2(n14640), .A(n13903), .ZN(n13909) );
  AOI21_X1 U15813 ( .B1(n13907), .B2(n13906), .A(n13905), .ZN(n14069) );
  NOR2_X1 U15814 ( .A1(n14069), .A2(n14016), .ZN(n13908) );
  OAI21_X1 U15815 ( .B1(n14648), .B2(n14068), .A(n13910), .ZN(P1_U3266) );
  OAI21_X1 U15816 ( .B1(n13913), .B2(n13912), .A(n13911), .ZN(n14077) );
  AOI21_X1 U15817 ( .B1(n13915), .B2(n13929), .A(n13914), .ZN(n14073) );
  AOI22_X1 U15818 ( .A1(n14008), .A2(n14071), .B1(n13916), .B2(n14637), .ZN(
        n13918) );
  NAND2_X1 U15819 ( .A1(n14638), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n13917) );
  OAI211_X1 U15820 ( .C1(n14070), .C2(n14640), .A(n13918), .B(n13917), .ZN(
        n13919) );
  AOI21_X1 U15821 ( .B1(n14073), .B2(n13920), .A(n13919), .ZN(n13925) );
  OAI21_X1 U15822 ( .B1(n13923), .B2(n13922), .A(n6840), .ZN(n14074) );
  NAND2_X1 U15823 ( .A1(n14074), .A2(n13987), .ZN(n13924) );
  OAI211_X1 U15824 ( .C1(n14077), .C2(n14016), .A(n13925), .B(n13924), .ZN(
        P1_U3267) );
  XOR2_X1 U15825 ( .A(n13926), .B(n13927), .Z(n14085) );
  OR2_X1 U15826 ( .A1(n13928), .A2(n13927), .ZN(n14079) );
  NAND3_X1 U15827 ( .A1(n14079), .A2(n14078), .A3(n14419), .ZN(n13940) );
  AOI21_X1 U15828 ( .B1(n13946), .B2(n14082), .A(n14675), .ZN(n13930) );
  AND2_X1 U15829 ( .A1(n13930), .A2(n13929), .ZN(n14080) );
  NAND2_X1 U15830 ( .A1(n14082), .A2(n14409), .ZN(n13937) );
  INV_X1 U15831 ( .A(n13931), .ZN(n13932) );
  OAI22_X1 U15832 ( .A1(n14648), .A2(n13933), .B1(n13932), .B2(n14612), .ZN(
        n13934) );
  INV_X1 U15833 ( .A(n13934), .ZN(n13936) );
  NAND2_X1 U15834 ( .A1(n14638), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n13935) );
  NAND3_X1 U15835 ( .A1(n13937), .A2(n13936), .A3(n13935), .ZN(n13938) );
  AOI21_X1 U15836 ( .B1(n14080), .B2(n14644), .A(n13938), .ZN(n13939) );
  OAI211_X1 U15837 ( .C1(n14032), .C2(n14085), .A(n13940), .B(n13939), .ZN(
        P1_U3268) );
  AOI21_X1 U15838 ( .B1(n13942), .B2(n13941), .A(n14608), .ZN(n13945) );
  AOI21_X1 U15839 ( .B1(n13945), .B2(n13944), .A(n13943), .ZN(n14088) );
  INV_X1 U15840 ( .A(n13946), .ZN(n13947) );
  AOI211_X1 U15841 ( .C1(n14087), .C2(n6954), .A(n14675), .B(n13947), .ZN(
        n14086) );
  AOI22_X1 U15842 ( .A1(n14638), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13948), 
        .B2(n14637), .ZN(n13949) );
  OAI21_X1 U15843 ( .B1(n13950), .B2(n14640), .A(n13949), .ZN(n13954) );
  AOI21_X1 U15844 ( .B1(n8683), .B2(n13952), .A(n13951), .ZN(n14090) );
  NOR2_X1 U15845 ( .A1(n14090), .A2(n14016), .ZN(n13953) );
  AOI211_X1 U15846 ( .C1(n14086), .C2(n14644), .A(n13954), .B(n13953), .ZN(
        n13955) );
  OAI21_X1 U15847 ( .B1(n14648), .B2(n14088), .A(n13955), .ZN(P1_U3269) );
  OAI21_X1 U15848 ( .B1(n13967), .B2(n13957), .A(n13956), .ZN(n13958) );
  INV_X1 U15849 ( .A(n13958), .ZN(n14098) );
  AOI211_X1 U15850 ( .C1(n14093), .C2(n13974), .A(n14675), .B(n13959), .ZN(
        n14091) );
  INV_X1 U15851 ( .A(n13960), .ZN(n14092) );
  AOI22_X1 U15852 ( .A1(n14008), .A2(n14092), .B1(n13961), .B2(n14637), .ZN(
        n13963) );
  NAND2_X1 U15853 ( .A1(n14638), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n13962) );
  OAI211_X1 U15854 ( .C1(n13964), .C2(n14640), .A(n13963), .B(n13962), .ZN(
        n13965) );
  AOI21_X1 U15855 ( .B1(n14091), .B2(n14644), .A(n13965), .ZN(n13969) );
  NAND2_X1 U15856 ( .A1(n13967), .A2(n13966), .ZN(n14094) );
  NAND3_X1 U15857 ( .A1(n14095), .A2(n14419), .A3(n14094), .ZN(n13968) );
  OAI211_X1 U15858 ( .C1(n14098), .C2(n14032), .A(n13969), .B(n13968), .ZN(
        P1_U3270) );
  XNOR2_X1 U15859 ( .A(n13971), .B(n13970), .ZN(n14105) );
  XNOR2_X1 U15860 ( .A(n13973), .B(n13972), .ZN(n14103) );
  OAI211_X1 U15861 ( .C1(n14101), .C2(n13988), .A(n14617), .B(n13974), .ZN(
        n14100) );
  INV_X1 U15862 ( .A(n13975), .ZN(n13976) );
  OAI22_X1 U15863 ( .A1(n14099), .A2(n14648), .B1(n13976), .B2(n14612), .ZN(
        n13978) );
  NOR2_X1 U15864 ( .A1(n14101), .A2(n14640), .ZN(n13977) );
  AOI211_X1 U15865 ( .C1(n14648), .C2(P1_REG2_REG_22__SCAN_IN), .A(n13978), 
        .B(n13977), .ZN(n13979) );
  OAI21_X1 U15866 ( .B1(n14011), .B2(n14100), .A(n13979), .ZN(n13980) );
  AOI21_X1 U15867 ( .B1(n14419), .B2(n14103), .A(n13980), .ZN(n13981) );
  OAI21_X1 U15868 ( .B1(n14105), .B2(n14032), .A(n13981), .ZN(P1_U3271) );
  INV_X1 U15869 ( .A(n13982), .ZN(n13983) );
  AOI21_X1 U15870 ( .B1(n13985), .B2(n13984), .A(n13983), .ZN(n14112) );
  XOR2_X1 U15871 ( .A(n13986), .B(n13985), .Z(n14109) );
  NAND2_X1 U15872 ( .A1(n14109), .A2(n13987), .ZN(n13995) );
  AOI211_X1 U15873 ( .C1(n14108), .C2(n14009), .A(n14675), .B(n13988), .ZN(
        n14106) );
  AOI22_X1 U15874 ( .A1(n14107), .A2(n14008), .B1(n13989), .B2(n14637), .ZN(
        n13991) );
  NAND2_X1 U15875 ( .A1(n14638), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n13990) );
  OAI211_X1 U15876 ( .C1(n13992), .C2(n14640), .A(n13991), .B(n13990), .ZN(
        n13993) );
  AOI21_X1 U15877 ( .B1(n14106), .B2(n14644), .A(n13993), .ZN(n13994) );
  OAI211_X1 U15878 ( .C1(n14112), .C2(n14016), .A(n13995), .B(n13994), .ZN(
        P1_U3272) );
  NAND2_X1 U15879 ( .A1(n13997), .A2(n13996), .ZN(n13998) );
  NAND2_X1 U15880 ( .A1(n13999), .A2(n13998), .ZN(n14116) );
  NAND2_X1 U15881 ( .A1(n14001), .A2(n14000), .ZN(n14002) );
  NAND3_X1 U15882 ( .A1(n14003), .A2(n14630), .A3(n14002), .ZN(n14005) );
  NAND2_X1 U15883 ( .A1(n14005), .A2(n14004), .ZN(n14118) );
  NAND2_X1 U15884 ( .A1(n14118), .A2(n14008), .ZN(n14015) );
  INV_X1 U15885 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n14007) );
  OAI22_X1 U15886 ( .A1(n14008), .A2(n14007), .B1(n14006), .B2(n14612), .ZN(
        n14013) );
  AOI21_X1 U15887 ( .B1(n14113), .B2(n14022), .A(n14675), .ZN(n14010) );
  NAND2_X1 U15888 ( .A1(n14010), .A2(n14009), .ZN(n14115) );
  NOR2_X1 U15889 ( .A1(n14115), .A2(n14011), .ZN(n14012) );
  AOI211_X1 U15890 ( .C1(n14409), .C2(n14113), .A(n14013), .B(n14012), .ZN(
        n14014) );
  OAI211_X1 U15891 ( .C1(n14116), .C2(n14016), .A(n14015), .B(n14014), .ZN(
        P1_U3273) );
  XNOR2_X1 U15892 ( .A(n14018), .B(n14017), .ZN(n14127) );
  XNOR2_X1 U15893 ( .A(n14020), .B(n14019), .ZN(n14125) );
  INV_X1 U15894 ( .A(n14121), .ZN(n14025) );
  INV_X1 U15895 ( .A(n14021), .ZN(n14039) );
  OAI211_X1 U15896 ( .C1(n14039), .C2(n14123), .A(n14617), .B(n14022), .ZN(
        n14122) );
  NOR2_X1 U15897 ( .A1(n14122), .A2(n14023), .ZN(n14024) );
  AOI211_X1 U15898 ( .C1(n14637), .C2(n14026), .A(n14025), .B(n14024), .ZN(
        n14029) );
  AOI22_X1 U15899 ( .A1(n14027), .A2(n14409), .B1(n14648), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n14028) );
  OAI21_X1 U15900 ( .B1(n14029), .B2(n14638), .A(n14028), .ZN(n14030) );
  AOI21_X1 U15901 ( .B1(n14419), .B2(n14125), .A(n14030), .ZN(n14031) );
  OAI21_X1 U15902 ( .B1(n14127), .B2(n14032), .A(n14031), .ZN(P1_U3274) );
  XNOR2_X1 U15903 ( .A(n14033), .B(n14034), .ZN(n14128) );
  XNOR2_X1 U15904 ( .A(n14035), .B(n14034), .ZN(n14037) );
  OAI21_X1 U15905 ( .B1(n14037), .B2(n14608), .A(n14036), .ZN(n14038) );
  AOI21_X1 U15906 ( .B1(n14712), .B2(n14128), .A(n14038), .ZN(n14132) );
  AOI211_X1 U15907 ( .C1(n14130), .C2(n14040), .A(n14675), .B(n14039), .ZN(
        n14129) );
  NAND2_X1 U15908 ( .A1(n14129), .A2(n14644), .ZN(n14043) );
  AOI22_X1 U15909 ( .A1(n14638), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14041), 
        .B2(n14637), .ZN(n14042) );
  OAI211_X1 U15910 ( .C1(n14044), .C2(n14640), .A(n14043), .B(n14042), .ZN(
        n14045) );
  AOI21_X1 U15911 ( .B1(n14645), .B2(n14128), .A(n14045), .ZN(n14046) );
  OAI21_X1 U15912 ( .B1(n14132), .B2(n14638), .A(n14046), .ZN(P1_U3275) );
  OAI211_X1 U15913 ( .C1(n14048), .C2(n14717), .A(n14047), .B(n14049), .ZN(
        n14135) );
  MUX2_X1 U15914 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14135), .S(n14740), .Z(
        P1_U3559) );
  INV_X1 U15915 ( .A(n14050), .ZN(n14051) );
  MUX2_X1 U15916 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14136), .S(n14740), .Z(
        P1_U3558) );
  OAI21_X1 U15917 ( .B1(n14054), .B2(n14717), .A(n14053), .ZN(n14055) );
  AOI21_X1 U15918 ( .B1(n14056), .B2(n14617), .A(n14055), .ZN(n14057) );
  AOI21_X1 U15919 ( .B1(n14706), .B2(n14061), .A(n14060), .ZN(n14062) );
  OAI211_X1 U15920 ( .C1(n14064), .C2(n14442), .A(n14063), .B(n14062), .ZN(
        n14137) );
  MUX2_X1 U15921 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14137), .S(n14740), .Z(
        P1_U3556) );
  AOI21_X1 U15922 ( .B1(n14706), .B2(n14066), .A(n14065), .ZN(n14067) );
  OAI211_X1 U15923 ( .C1(n14069), .C2(n14442), .A(n14068), .B(n14067), .ZN(
        n14138) );
  MUX2_X1 U15924 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14138), .S(n14740), .Z(
        P1_U3555) );
  NOR2_X1 U15925 ( .A1(n14070), .A2(n14717), .ZN(n14072) );
  AOI211_X1 U15926 ( .C1(n14073), .C2(n14617), .A(n14072), .B(n14071), .ZN(
        n14076) );
  NAND2_X1 U15927 ( .A1(n14074), .A2(n14630), .ZN(n14075) );
  OAI211_X1 U15928 ( .C1(n14077), .C2(n14442), .A(n14076), .B(n14075), .ZN(
        n14139) );
  MUX2_X1 U15929 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14139), .S(n14740), .Z(
        P1_U3554) );
  NAND3_X1 U15930 ( .A1(n14079), .A2(n14078), .A3(n14714), .ZN(n14084) );
  AOI211_X1 U15931 ( .C1(n14706), .C2(n14082), .A(n14081), .B(n14080), .ZN(
        n14083) );
  OAI211_X1 U15932 ( .C1(n14608), .C2(n14085), .A(n14084), .B(n14083), .ZN(
        n14140) );
  MUX2_X1 U15933 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14140), .S(n14740), .Z(
        P1_U3553) );
  AOI21_X1 U15934 ( .B1(n14706), .B2(n14087), .A(n14086), .ZN(n14089) );
  OAI211_X1 U15935 ( .C1(n14442), .C2(n14090), .A(n14089), .B(n14088), .ZN(
        n14141) );
  MUX2_X1 U15936 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14141), .S(n14740), .Z(
        P1_U3552) );
  AOI211_X1 U15937 ( .C1(n14706), .C2(n14093), .A(n14092), .B(n14091), .ZN(
        n14097) );
  NAND3_X1 U15938 ( .A1(n14095), .A2(n14714), .A3(n14094), .ZN(n14096) );
  OAI211_X1 U15939 ( .C1(n14608), .C2(n14098), .A(n14097), .B(n14096), .ZN(
        n14142) );
  MUX2_X1 U15940 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14142), .S(n14740), .Z(
        P1_U3551) );
  OAI211_X1 U15941 ( .C1(n14717), .C2(n14101), .A(n14100), .B(n14099), .ZN(
        n14102) );
  AOI21_X1 U15942 ( .B1(n14103), .B2(n14714), .A(n14102), .ZN(n14104) );
  OAI21_X1 U15943 ( .B1(n14105), .B2(n14608), .A(n14104), .ZN(n14143) );
  MUX2_X1 U15944 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14143), .S(n14740), .Z(
        P1_U3550) );
  AOI211_X1 U15945 ( .C1(n14706), .C2(n14108), .A(n14107), .B(n14106), .ZN(
        n14111) );
  NAND2_X1 U15946 ( .A1(n14109), .A2(n14630), .ZN(n14110) );
  OAI211_X1 U15947 ( .C1(n14112), .C2(n14442), .A(n14111), .B(n14110), .ZN(
        n14144) );
  MUX2_X1 U15948 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14144), .S(n14740), .Z(
        P1_U3549) );
  NAND2_X1 U15949 ( .A1(n14113), .A2(n14706), .ZN(n14114) );
  OAI211_X1 U15950 ( .C1(n14116), .C2(n14442), .A(n14115), .B(n14114), .ZN(
        n14117) );
  NOR2_X1 U15951 ( .A1(n14118), .A2(n14117), .ZN(n14145) );
  MUX2_X1 U15952 ( .A(n14119), .B(n14145), .S(n14740), .Z(n14120) );
  INV_X1 U15953 ( .A(n14120), .ZN(P1_U3548) );
  OAI211_X1 U15954 ( .C1(n14123), .C2(n14717), .A(n14122), .B(n14121), .ZN(
        n14124) );
  AOI21_X1 U15955 ( .B1(n14125), .B2(n14714), .A(n14124), .ZN(n14126) );
  OAI21_X1 U15956 ( .B1(n14127), .B2(n14608), .A(n14126), .ZN(n14148) );
  MUX2_X1 U15957 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14148), .S(n14740), .Z(
        P1_U3547) );
  INV_X1 U15958 ( .A(n14128), .ZN(n14133) );
  AOI21_X1 U15959 ( .B1(n14706), .B2(n14130), .A(n14129), .ZN(n14131) );
  OAI211_X1 U15960 ( .C1(n14133), .C2(n14709), .A(n14132), .B(n14131), .ZN(
        n14149) );
  MUX2_X1 U15961 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14149), .S(n14740), .Z(
        P1_U3546) );
  MUX2_X1 U15962 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n14134), .S(n14740), .Z(
        P1_U3528) );
  MUX2_X1 U15963 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14135), .S(n14724), .Z(
        P1_U3527) );
  MUX2_X1 U15964 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14136), .S(n14724), .Z(
        P1_U3526) );
  MUX2_X1 U15965 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14137), .S(n14724), .Z(
        P1_U3524) );
  MUX2_X1 U15966 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14138), .S(n14724), .Z(
        P1_U3523) );
  MUX2_X1 U15967 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14139), .S(n14724), .Z(
        P1_U3522) );
  MUX2_X1 U15968 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14140), .S(n14724), .Z(
        P1_U3521) );
  MUX2_X1 U15969 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14141), .S(n14724), .Z(
        P1_U3520) );
  MUX2_X1 U15970 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14142), .S(n14724), .Z(
        P1_U3519) );
  MUX2_X1 U15971 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14143), .S(n14724), .Z(
        P1_U3518) );
  MUX2_X1 U15972 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14144), .S(n14724), .Z(
        P1_U3517) );
  INV_X1 U15973 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n14146) );
  MUX2_X1 U15974 ( .A(n14146), .B(n14145), .S(n14724), .Z(n14147) );
  INV_X1 U15975 ( .A(n14147), .ZN(P1_U3516) );
  MUX2_X1 U15976 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14148), .S(n14724), .Z(
        P1_U3515) );
  MUX2_X1 U15977 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14149), .S(n14724), .Z(
        P1_U3513) );
  NOR4_X1 U15978 ( .A1(n6823), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8241), .A4(
        P1_U3086), .ZN(n14150) );
  AOI21_X1 U15979 ( .B1(n14151), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14150), 
        .ZN(n14152) );
  OAI21_X1 U15980 ( .B1(n14153), .B2(n14171), .A(n14152), .ZN(P1_U3324) );
  OAI222_X1 U15981 ( .A1(P1_U3086), .A2(n14155), .B1(n14166), .B2(n14154), 
        .C1(n15205), .C2(n14163), .ZN(P1_U3326) );
  INV_X1 U15982 ( .A(n14156), .ZN(n14158) );
  OAI222_X1 U15983 ( .A1(P1_U3086), .A2(n14159), .B1(n14166), .B2(n14158), 
        .C1(n14157), .C2(n14163), .ZN(P1_U3327) );
  OAI222_X1 U15984 ( .A1(n6459), .A2(P1_U3086), .B1(n14166), .B2(n14161), .C1(
        n14160), .C2(n14163), .ZN(P1_U3328) );
  INV_X1 U15985 ( .A(n14162), .ZN(n14167) );
  OAI222_X1 U15986 ( .A1(P1_U3086), .A2(n14167), .B1(n14166), .B2(n14165), 
        .C1(n14164), .C2(n14163), .ZN(P1_U3329) );
  INV_X1 U15987 ( .A(n14168), .ZN(n14173) );
  OAI222_X1 U15988 ( .A1(n14173), .A2(P1_U3086), .B1(n14171), .B2(n14170), 
        .C1(n14169), .C2(n14163), .ZN(P1_U3330) );
  MUX2_X1 U15989 ( .A(n14174), .B(n9504), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U15990 ( .A(n14175), .ZN(n14176) );
  MUX2_X1 U15991 ( .A(n14176), .B(n6720), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3355) );
  INV_X1 U15992 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14541) );
  XOR2_X1 U15993 ( .A(n14210), .B(n14541), .Z(n14220) );
  INV_X1 U15994 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14208) );
  INV_X1 U15995 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14206) );
  INV_X1 U15996 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14507) );
  INV_X1 U15997 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14199) );
  INV_X1 U15998 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14952) );
  XNOR2_X1 U15999 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n14226) );
  XOR2_X1 U16000 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n14180), .Z(n14236) );
  AND2_X1 U16001 ( .A1(n14179), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n14178) );
  INV_X1 U16002 ( .A(n14231), .ZN(n14177) );
  NAND2_X1 U16003 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14181), .ZN(n14184) );
  NAND2_X1 U16004 ( .A1(n14240), .A2(n14182), .ZN(n14183) );
  NAND2_X1 U16005 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14185), .ZN(n14187) );
  NAND2_X1 U16006 ( .A1(n14228), .A2(n14229), .ZN(n14186) );
  NAND2_X1 U16007 ( .A1(n14187), .A2(n14186), .ZN(n14188) );
  NAND2_X1 U16008 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14188), .ZN(n14190) );
  XOR2_X1 U16009 ( .A(n14188), .B(P3_ADDR_REG_5__SCAN_IN), .Z(n14248) );
  INV_X1 U16010 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14249) );
  NAND2_X1 U16011 ( .A1(n14248), .A2(n14249), .ZN(n14189) );
  NAND2_X1 U16012 ( .A1(n14190), .A2(n14189), .ZN(n14255) );
  NAND2_X1 U16013 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n14191), .ZN(n14192) );
  NAND2_X1 U16014 ( .A1(n14194), .A2(n10674), .ZN(n14196) );
  XNOR2_X1 U16015 ( .A(n14194), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14260) );
  NAND2_X1 U16016 ( .A1(n14260), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14195) );
  NAND2_X1 U16017 ( .A1(n14196), .A2(n14195), .ZN(n14227) );
  XNOR2_X1 U16018 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n14266) );
  NAND2_X1 U16019 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n14200), .ZN(n14203) );
  XOR2_X1 U16020 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(n14200), .Z(n14225) );
  INV_X1 U16021 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14201) );
  NAND2_X1 U16022 ( .A1(n14225), .A2(n14201), .ZN(n14202) );
  NAND2_X1 U16023 ( .A1(n14203), .A2(n14202), .ZN(n14270) );
  XNOR2_X1 U16024 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(n14507), .ZN(n14269) );
  NOR2_X1 U16025 ( .A1(n14270), .A2(n14269), .ZN(n14204) );
  XOR2_X1 U16026 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n14223) );
  NOR2_X1 U16027 ( .A1(n14224), .A2(n14223), .ZN(n14205) );
  INV_X1 U16028 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14524) );
  NOR2_X1 U16029 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14524), .ZN(n14207) );
  NOR2_X1 U16030 ( .A1(n14220), .A2(n14219), .ZN(n14209) );
  AOI21_X1 U16031 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n14210), .A(n14209), 
        .ZN(n14278) );
  NAND2_X1 U16032 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14211), .ZN(n14213) );
  INV_X1 U16033 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14212) );
  AOI22_X1 U16034 ( .A1(n14278), .A2(n14213), .B1(P3_ADDR_REG_15__SCAN_IN), 
        .B2(n14212), .ZN(n14282) );
  INV_X1 U16035 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14553) );
  NAND2_X1 U16036 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14553), .ZN(n14214) );
  AOI22_X1 U16037 ( .A1(n14282), .A2(n14214), .B1(P1_ADDR_REG_16__SCAN_IN), 
        .B2(n14281), .ZN(n14215) );
  INV_X1 U16038 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14570) );
  NAND2_X1 U16039 ( .A1(n14215), .A2(n14570), .ZN(n14217) );
  XNOR2_X1 U16040 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14215), .ZN(n14287) );
  NAND2_X1 U16041 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14287), .ZN(n14216) );
  NAND2_X1 U16042 ( .A1(n14217), .A2(n14216), .ZN(n14322) );
  NOR2_X1 U16043 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n14325), .ZN(n14218) );
  AOI21_X1 U16044 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n14325), .A(n14218), 
        .ZN(n14323) );
  XNOR2_X1 U16045 ( .A(n14322), .B(n14323), .ZN(n14319) );
  INV_X1 U16046 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14810) );
  XOR2_X1 U16047 ( .A(n14220), .B(n14219), .Z(n14478) );
  XNOR2_X1 U16048 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n14222) );
  XOR2_X1 U16049 ( .A(n14222), .B(n14221), .Z(n14273) );
  XNOR2_X1 U16050 ( .A(n14224), .B(n14223), .ZN(n14474) );
  INV_X1 U16051 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14303) );
  XNOR2_X1 U16052 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14225), .ZN(n14301) );
  INV_X1 U16053 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14796) );
  XOR2_X1 U16054 ( .A(n14227), .B(n14226), .Z(n14265) );
  NOR2_X1 U16055 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14245), .ZN(n14247) );
  XNOR2_X1 U16056 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14230) );
  XNOR2_X1 U16057 ( .A(n14230), .B(n14231), .ZN(n14233) );
  NAND2_X1 U16058 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14233), .ZN(n14235) );
  AOI21_X1 U16059 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14232), .A(n14231), .ZN(
        n15288) );
  NOR2_X1 U16060 ( .A1(n15288), .A2(n10179), .ZN(n15293) );
  NAND2_X1 U16061 ( .A1(n15293), .A2(n15292), .ZN(n14234) );
  NAND2_X1 U16062 ( .A1(n14235), .A2(n14234), .ZN(n14292) );
  XNOR2_X1 U16063 ( .A(n14237), .B(n14236), .ZN(n14291) );
  NOR2_X1 U16064 ( .A1(n14292), .A2(n14291), .ZN(n14239) );
  INV_X1 U16065 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14238) );
  NAND2_X1 U16066 ( .A1(n14292), .A2(n14291), .ZN(n14290) );
  OAI21_X1 U16067 ( .B1(n14239), .B2(n14238), .A(n14290), .ZN(n14242) );
  XOR2_X1 U16068 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14240), .Z(n14241) );
  NOR2_X1 U16069 ( .A1(n14242), .A2(n14241), .ZN(n14244) );
  XNOR2_X1 U16070 ( .A(n14242), .B(n14241), .ZN(n15291) );
  NOR2_X1 U16071 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15291), .ZN(n14243) );
  NOR2_X1 U16072 ( .A1(n14244), .A2(n14243), .ZN(n15286) );
  NOR2_X1 U16073 ( .A1(n15286), .A2(n15285), .ZN(n14246) );
  NOR2_X1 U16074 ( .A1(n14247), .A2(n14246), .ZN(n14251) );
  XNOR2_X1 U16075 ( .A(n14249), .B(n14248), .ZN(n14250) );
  NOR2_X1 U16076 ( .A1(n14251), .A2(n14250), .ZN(n14253) );
  XNOR2_X1 U16077 ( .A(n14251), .B(n14250), .ZN(n15287) );
  NOR2_X1 U16078 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15287), .ZN(n14252) );
  XOR2_X1 U16079 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), .Z(
        n14254) );
  XOR2_X1 U16080 ( .A(n14255), .B(n14254), .Z(n14294) );
  NAND2_X1 U16081 ( .A1(n14256), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14257) );
  NAND2_X1 U16082 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14259), .ZN(n14263) );
  INV_X1 U16083 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n14258) );
  XNOR2_X1 U16084 ( .A(n14261), .B(n14260), .ZN(n15289) );
  NAND2_X1 U16085 ( .A1(n15290), .A2(n15289), .ZN(n14262) );
  XNOR2_X1 U16086 ( .A(n14267), .B(n14266), .ZN(n14298) );
  NAND2_X1 U16087 ( .A1(n14299), .A2(n14298), .ZN(n14268) );
  NOR2_X1 U16088 ( .A1(n14299), .A2(n14298), .ZN(n14297) );
  XNOR2_X1 U16089 ( .A(n14270), .B(n14269), .ZN(n14470) );
  INV_X1 U16090 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14271) );
  NAND2_X1 U16091 ( .A1(n14469), .A2(n14470), .ZN(n14468) );
  NOR2_X1 U16092 ( .A1(n14273), .A2(n14274), .ZN(n14276) );
  NAND2_X1 U16093 ( .A1(n14478), .A2(n14479), .ZN(n14277) );
  XNOR2_X1 U16094 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14279) );
  XNOR2_X1 U16095 ( .A(n14279), .B(n14278), .ZN(n14481) );
  NAND2_X1 U16096 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14281), .ZN(n14280) );
  OAI21_X1 U16097 ( .B1(n14281), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14280), 
        .ZN(n14283) );
  XOR2_X1 U16098 ( .A(n14283), .B(n14282), .Z(n14284) );
  AND2_X1 U16099 ( .A1(n14285), .A2(n14284), .ZN(n14485) );
  NOR2_X1 U16100 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n14484), .ZN(n14286) );
  XNOR2_X1 U16101 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14287), .ZN(n14315) );
  XNOR2_X1 U16102 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14317), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16103 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14288) );
  OAI21_X1 U16104 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14288), 
        .ZN(U28) );
  AOI21_X1 U16105 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14289) );
  OAI21_X1 U16106 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14289), 
        .ZN(U29) );
  OAI21_X1 U16107 ( .B1(n14292), .B2(n14291), .A(n14290), .ZN(n14293) );
  XNOR2_X1 U16108 ( .A(n14293), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  XOR2_X1 U16109 ( .A(n14295), .B(n14294), .Z(SUB_1596_U57) );
  XNOR2_X1 U16110 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14296), .ZN(SUB_1596_U55)
         );
  AOI21_X1 U16111 ( .B1(n14299), .B2(n14298), .A(n14297), .ZN(n14300) );
  XNOR2_X1 U16112 ( .A(n14300), .B(n14796), .ZN(SUB_1596_U54) );
  AOI21_X1 U16113 ( .B1(n14302), .B2(n14301), .A(n6597), .ZN(n14304) );
  XNOR2_X1 U16114 ( .A(n14304), .B(n14303), .ZN(SUB_1596_U70) );
  AND2_X1 U16115 ( .A1(n14305), .A2(n14714), .ZN(n14308) );
  OAI22_X1 U16116 ( .A1(n14306), .A2(n14675), .B1(n6961), .B2(n14717), .ZN(
        n14307) );
  NOR3_X1 U16117 ( .A1(n14309), .A2(n14308), .A3(n14307), .ZN(n14312) );
  INV_X1 U16118 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14310) );
  AOI22_X1 U16119 ( .A1(n14724), .A2(n14312), .B1(n14310), .B2(n14722), .ZN(
        P1_U3495) );
  AOI22_X1 U16120 ( .A1(n14740), .A2(n14312), .B1(n14311), .B2(n14738), .ZN(
        P1_U3540) );
  OAI21_X1 U16121 ( .B1(n14315), .B2(n14314), .A(n14313), .ZN(n14316) );
  XNOR2_X1 U16122 ( .A(n14316), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  NOR2_X1 U16123 ( .A1(n14319), .A2(n14318), .ZN(n14320) );
  NOR2_X1 U16124 ( .A1(n14321), .A2(n14320), .ZN(n14330) );
  NAND2_X1 U16125 ( .A1(n14323), .A2(n14322), .ZN(n14324) );
  OAI21_X1 U16126 ( .B1(n14325), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n14324), 
        .ZN(n14328) );
  XNOR2_X1 U16127 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(n6894), .ZN(n14326) );
  XNOR2_X1 U16128 ( .A(n11994), .B(n14326), .ZN(n14327) );
  XNOR2_X1 U16129 ( .A(n14328), .B(n14327), .ZN(n14329) );
  XNOR2_X1 U16130 ( .A(n14330), .B(n14329), .ZN(SUB_1596_U4) );
  NOR2_X1 U16131 ( .A1(n14332), .A2(n14331), .ZN(n14354) );
  AOI22_X1 U16132 ( .A1(n14333), .A2(n15046), .B1(n14354), .B2(n15050), .ZN(
        n14338) );
  INV_X1 U16133 ( .A(n14958), .ZN(n14336) );
  AOI22_X1 U16134 ( .A1(n9315), .A2(n14336), .B1(n14334), .B2(
        P3_REG2_REG_31__SCAN_IN), .ZN(n14335) );
  NAND2_X1 U16135 ( .A1(n14338), .A2(n14335), .ZN(P3_U3202) );
  AOI22_X1 U16136 ( .A1(n14355), .A2(n14336), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n14334), .ZN(n14337) );
  NAND2_X1 U16137 ( .A1(n14338), .A2(n14337), .ZN(P3_U3203) );
  XNOR2_X1 U16138 ( .A(n14340), .B(n14339), .ZN(n14359) );
  OAI211_X1 U16139 ( .C1(n14343), .C2(n14342), .A(n14341), .B(n15039), .ZN(
        n14346) );
  NAND2_X1 U16140 ( .A1(n14344), .A2(n15035), .ZN(n14345) );
  OAI211_X1 U16141 ( .C1(n14347), .C2(n15019), .A(n14346), .B(n14345), .ZN(
        n14357) );
  AOI21_X1 U16142 ( .B1(n14359), .B2(n14953), .A(n14357), .ZN(n14352) );
  INV_X1 U16143 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n14351) );
  NOR2_X1 U16144 ( .A1(n14348), .A2(n15030), .ZN(n14358) );
  AOI22_X1 U16145 ( .A1(n14358), .A2(n15000), .B1(n15046), .B2(n14349), .ZN(
        n14350) );
  OAI221_X1 U16146 ( .B1(n14334), .B2(n14352), .C1(n15050), .C2(n14351), .A(
        n14350), .ZN(P3_U3221) );
  AOI21_X1 U16147 ( .B1(n9315), .B2(n15023), .A(n14354), .ZN(n14367) );
  INV_X1 U16148 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14353) );
  AOI22_X1 U16149 ( .A1(n15096), .A2(n14367), .B1(n14353), .B2(n15094), .ZN(
        P3_U3490) );
  AOI21_X1 U16150 ( .B1(n14355), .B2(n15023), .A(n14354), .ZN(n14369) );
  INV_X1 U16151 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14356) );
  AOI22_X1 U16152 ( .A1(n15096), .A2(n14369), .B1(n14356), .B2(n15094), .ZN(
        P3_U3489) );
  AOI211_X1 U16153 ( .C1(n14359), .C2(n14362), .A(n14358), .B(n14357), .ZN(
        n14370) );
  INV_X1 U16154 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14360) );
  AOI22_X1 U16155 ( .A1(n15096), .A2(n14370), .B1(n14360), .B2(n15094), .ZN(
        P3_U3471) );
  AOI21_X1 U16156 ( .B1(n14363), .B2(n14362), .A(n14361), .ZN(n14364) );
  AOI22_X1 U16157 ( .A1(n15096), .A2(n14371), .B1(n11520), .B2(n15094), .ZN(
        P3_U3470) );
  AOI22_X1 U16158 ( .A1(n15081), .A2(n14367), .B1(n14366), .B2(n15080), .ZN(
        P3_U3458) );
  AOI22_X1 U16159 ( .A1(n15081), .A2(n14369), .B1(n14368), .B2(n15080), .ZN(
        P3_U3457) );
  AOI22_X1 U16160 ( .A1(n15081), .A2(n14370), .B1(n8978), .B2(n15080), .ZN(
        P3_U3426) );
  AOI22_X1 U16161 ( .A1(n15081), .A2(n14371), .B1(n8955), .B2(n15080), .ZN(
        P3_U3423) );
  NAND2_X1 U16162 ( .A1(n14373), .A2(n14374), .ZN(n14375) );
  NAND2_X1 U16163 ( .A1(n14372), .A2(n14375), .ZN(n14377) );
  AOI222_X1 U16164 ( .A1(n14381), .A2(n14380), .B1(n14379), .B2(n14378), .C1(
        n14377), .C2(n14376), .ZN(n14382) );
  NAND2_X1 U16165 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14797)
         );
  OAI211_X1 U16166 ( .C1(n14384), .C2(n14383), .A(n14382), .B(n14797), .ZN(
        P2_U3187) );
  OR2_X1 U16167 ( .A1(n14386), .A2(n14385), .ZN(n14390) );
  NAND2_X1 U16168 ( .A1(n14388), .A2(n14387), .ZN(n14389) );
  NAND2_X1 U16169 ( .A1(n14390), .A2(n14389), .ZN(n14405) );
  NAND2_X1 U16170 ( .A1(n14392), .A2(n14391), .ZN(n14393) );
  NAND2_X1 U16171 ( .A1(n14394), .A2(n14393), .ZN(n14396) );
  AOI222_X1 U16172 ( .A1(n14398), .A2(n14414), .B1(n14405), .B2(n14397), .C1(
        n14396), .C2(n14395), .ZN(n14399) );
  NAND2_X1 U16173 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14539)
         );
  OAI211_X1 U16174 ( .C1(n14401), .C2(n14400), .A(n14399), .B(n14539), .ZN(
        P1_U3215) );
  INV_X1 U16175 ( .A(n14402), .ZN(n14404) );
  INV_X1 U16176 ( .A(n14413), .ZN(n14403) );
  AOI21_X1 U16177 ( .B1(n14404), .B2(n14403), .A(n14608), .ZN(n14407) );
  AOI21_X1 U16178 ( .B1(n14407), .B2(n14406), .A(n14405), .ZN(n14448) );
  AOI222_X1 U16179 ( .A1(n14414), .A2(n14409), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n14638), .C1(n14408), .C2(n14637), .ZN(n14421) );
  INV_X1 U16180 ( .A(n14410), .ZN(n14411) );
  AOI21_X1 U16181 ( .B1(n14413), .B2(n14412), .A(n14411), .ZN(n14451) );
  INV_X1 U16182 ( .A(n14414), .ZN(n14447) );
  INV_X1 U16183 ( .A(n14415), .ZN(n14417) );
  OAI211_X1 U16184 ( .C1(n14447), .C2(n14417), .A(n14617), .B(n14416), .ZN(
        n14446) );
  INV_X1 U16185 ( .A(n14446), .ZN(n14418) );
  AOI22_X1 U16186 ( .A1(n14451), .A2(n14419), .B1(n14644), .B2(n14418), .ZN(
        n14420) );
  OAI211_X1 U16187 ( .C1(n14648), .C2(n14448), .A(n14421), .B(n14420), .ZN(
        P1_U3279) );
  AOI21_X1 U16188 ( .B1(n14423), .B2(n14706), .A(n14422), .ZN(n14425) );
  OAI211_X1 U16189 ( .C1(n14426), .C2(n14442), .A(n14425), .B(n14424), .ZN(
        n14427) );
  AOI21_X1 U16190 ( .B1(n14630), .B2(n14428), .A(n14427), .ZN(n14460) );
  AOI22_X1 U16191 ( .A1(n14740), .A2(n14460), .B1(n13846), .B2(n14738), .ZN(
        P1_U3545) );
  AOI21_X1 U16192 ( .B1(n14430), .B2(n14706), .A(n14429), .ZN(n14432) );
  OAI211_X1 U16193 ( .C1(n14433), .C2(n14608), .A(n14432), .B(n14431), .ZN(
        n14434) );
  AOI21_X1 U16194 ( .B1(n14435), .B2(n14714), .A(n14434), .ZN(n14462) );
  INV_X1 U16195 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14436) );
  AOI22_X1 U16196 ( .A1(n14740), .A2(n14462), .B1(n14436), .B2(n14738), .ZN(
        P1_U3544) );
  AOI211_X1 U16197 ( .C1(n14706), .C2(n14439), .A(n14438), .B(n14437), .ZN(
        n14441) );
  OAI211_X1 U16198 ( .C1(n14443), .C2(n14442), .A(n14441), .B(n14440), .ZN(
        n14444) );
  INV_X1 U16199 ( .A(n14444), .ZN(n14464) );
  AOI22_X1 U16200 ( .A1(n14740), .A2(n14464), .B1(n14445), .B2(n14738), .ZN(
        P1_U3543) );
  OAI21_X1 U16201 ( .B1(n14447), .B2(n14717), .A(n14446), .ZN(n14450) );
  INV_X1 U16202 ( .A(n14448), .ZN(n14449) );
  AOI211_X1 U16203 ( .C1(n14451), .C2(n14714), .A(n14450), .B(n14449), .ZN(
        n14465) );
  AOI22_X1 U16204 ( .A1(n14740), .A2(n14465), .B1(n11861), .B2(n14738), .ZN(
        P1_U3542) );
  AND2_X1 U16205 ( .A1(n14452), .A2(n14714), .ZN(n14458) );
  NAND2_X1 U16206 ( .A1(n14453), .A2(n14706), .ZN(n14454) );
  NAND2_X1 U16207 ( .A1(n14455), .A2(n14454), .ZN(n14456) );
  NOR3_X1 U16208 ( .A1(n14458), .A2(n14457), .A3(n14456), .ZN(n14467) );
  AOI22_X1 U16209 ( .A1(n14740), .A2(n14467), .B1(n11429), .B2(n14738), .ZN(
        P1_U3539) );
  INV_X1 U16210 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14459) );
  AOI22_X1 U16211 ( .A1(n14724), .A2(n14460), .B1(n14459), .B2(n14722), .ZN(
        P1_U3510) );
  INV_X1 U16212 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14461) );
  AOI22_X1 U16213 ( .A1(n14724), .A2(n14462), .B1(n14461), .B2(n14722), .ZN(
        P1_U3507) );
  INV_X1 U16214 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14463) );
  AOI22_X1 U16215 ( .A1(n14724), .A2(n14464), .B1(n14463), .B2(n14722), .ZN(
        P1_U3504) );
  AOI22_X1 U16216 ( .A1(n14724), .A2(n14465), .B1(n8449), .B2(n14722), .ZN(
        P1_U3501) );
  INV_X1 U16217 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14466) );
  AOI22_X1 U16218 ( .A1(n14724), .A2(n14467), .B1(n14466), .B2(n14722), .ZN(
        P1_U3492) );
  OAI21_X1 U16219 ( .B1(n14470), .B2(n14469), .A(n14468), .ZN(n14471) );
  XNOR2_X1 U16220 ( .A(n14471), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16221 ( .B1(n14474), .B2(n14473), .A(n14472), .ZN(n14475) );
  XNOR2_X1 U16222 ( .A(n14475), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  XNOR2_X1 U16223 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14476), .ZN(SUB_1596_U67)
         );
  AOI21_X1 U16224 ( .B1(n14479), .B2(n14478), .A(n14477), .ZN(n14480) );
  XNOR2_X1 U16225 ( .A(n14480), .B(n14810), .ZN(SUB_1596_U66) );
  AOI21_X1 U16226 ( .B1(n14482), .B2(n14481), .A(n6557), .ZN(n14483) );
  XOR2_X1 U16227 ( .A(n14483), .B(P2_ADDR_REG_15__SCAN_IN), .Z(SUB_1596_U65)
         );
  NOR2_X1 U16228 ( .A1(n14485), .A2(n14484), .ZN(n14486) );
  XOR2_X1 U16229 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14486), .Z(SUB_1596_U64)
         );
  AOI21_X1 U16230 ( .B1(n6459), .B2(n14488), .A(n14487), .ZN(n14490) );
  XNOR2_X1 U16231 ( .A(n14490), .B(n6720), .ZN(n14494) );
  AOI22_X1 U16232 ( .A1(n14491), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14492) );
  OAI21_X1 U16233 ( .B1(n14494), .B2(n14493), .A(n14492), .ZN(P1_U3243) );
  OAI21_X1 U16234 ( .B1(n14497), .B2(n14496), .A(n14495), .ZN(n14504) );
  NOR2_X1 U16235 ( .A1(n14566), .A2(n14498), .ZN(n14503) );
  AOI211_X1 U16236 ( .C1(n14501), .C2(n14500), .A(n14572), .B(n14499), .ZN(
        n14502) );
  AOI211_X1 U16237 ( .C1(n14558), .C2(n14504), .A(n14503), .B(n14502), .ZN(
        n14506) );
  OAI211_X1 U16238 ( .C1(n14507), .C2(n14585), .A(n14506), .B(n14505), .ZN(
        P1_U3254) );
  NAND2_X1 U16239 ( .A1(n14509), .A2(n14508), .ZN(n14512) );
  NOR2_X1 U16240 ( .A1(n14576), .A2(n14510), .ZN(n14511) );
  NAND2_X1 U16241 ( .A1(n14512), .A2(n14511), .ZN(n14519) );
  NAND2_X1 U16242 ( .A1(n14514), .A2(n14513), .ZN(n14517) );
  NOR2_X1 U16243 ( .A1(n14572), .A2(n14515), .ZN(n14516) );
  NAND2_X1 U16244 ( .A1(n14517), .A2(n14516), .ZN(n14518) );
  OAI211_X1 U16245 ( .C1(n14566), .C2(n14520), .A(n14519), .B(n14518), .ZN(
        n14521) );
  INV_X1 U16246 ( .A(n14521), .ZN(n14523) );
  OAI211_X1 U16247 ( .C1(n14524), .C2(n14585), .A(n14523), .B(n14522), .ZN(
        P1_U3256) );
  INV_X1 U16248 ( .A(n14525), .ZN(n14537) );
  NAND2_X1 U16249 ( .A1(n14527), .A2(n14526), .ZN(n14530) );
  INV_X1 U16250 ( .A(n14528), .ZN(n14529) );
  NAND3_X1 U16251 ( .A1(n14554), .A2(n14530), .A3(n14529), .ZN(n14536) );
  OAI21_X1 U16252 ( .B1(n14533), .B2(n14532), .A(n14531), .ZN(n14534) );
  NAND2_X1 U16253 ( .A1(n14558), .A2(n14534), .ZN(n14535) );
  OAI211_X1 U16254 ( .C1(n14566), .C2(n14537), .A(n14536), .B(n14535), .ZN(
        n14538) );
  INV_X1 U16255 ( .A(n14538), .ZN(n14540) );
  OAI211_X1 U16256 ( .C1(n14541), .C2(n14585), .A(n14540), .B(n14539), .ZN(
        P1_U3257) );
  OAI211_X1 U16257 ( .C1(n7503), .C2(n14543), .A(n14542), .B(n14554), .ZN(
        n14548) );
  OAI211_X1 U16258 ( .C1(n14546), .C2(n14545), .A(n14544), .B(n14558), .ZN(
        n14547) );
  OAI211_X1 U16259 ( .C1(n14566), .C2(n14549), .A(n14548), .B(n14547), .ZN(
        n14550) );
  INV_X1 U16260 ( .A(n14550), .ZN(n14552) );
  OAI211_X1 U16261 ( .C1(n14553), .C2(n14585), .A(n14552), .B(n14551), .ZN(
        P1_U3259) );
  OAI211_X1 U16262 ( .C1(n14557), .C2(n14556), .A(n14555), .B(n14554), .ZN(
        n14564) );
  OAI21_X1 U16263 ( .B1(n14560), .B2(n14559), .A(n14558), .ZN(n14561) );
  OR2_X1 U16264 ( .A1(n14562), .A2(n14561), .ZN(n14563) );
  OAI211_X1 U16265 ( .C1(n14566), .C2(n14565), .A(n14564), .B(n14563), .ZN(
        n14567) );
  INV_X1 U16266 ( .A(n14567), .ZN(n14569) );
  OAI211_X1 U16267 ( .C1(n14570), .C2(n14585), .A(n14569), .B(n14568), .ZN(
        P1_U3260) );
  INV_X1 U16268 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14586) );
  AOI211_X1 U16269 ( .C1(n8501), .C2(n14573), .A(n14572), .B(n14571), .ZN(
        n14580) );
  INV_X1 U16270 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14578) );
  INV_X1 U16271 ( .A(n14574), .ZN(n14577) );
  AOI211_X1 U16272 ( .C1(n14578), .C2(n14577), .A(n14576), .B(n14575), .ZN(
        n14579) );
  AOI211_X1 U16273 ( .C1(n14582), .C2(n14581), .A(n14580), .B(n14579), .ZN(
        n14584) );
  OAI211_X1 U16274 ( .C1(n14586), .C2(n14585), .A(n14584), .B(n14583), .ZN(
        P1_U3261) );
  XNOR2_X1 U16275 ( .A(n14588), .B(n14589), .ZN(n14686) );
  XNOR2_X1 U16276 ( .A(n14590), .B(n14589), .ZN(n14591) );
  NOR2_X1 U16277 ( .A1(n14591), .A2(n14608), .ZN(n14592) );
  AOI211_X1 U16278 ( .C1(n14712), .C2(n14686), .A(n14593), .B(n14592), .ZN(
        n14683) );
  NOR2_X1 U16279 ( .A1(n14612), .A2(n14594), .ZN(n14595) );
  AOI21_X1 U16280 ( .B1(n14648), .B2(P1_REG2_REG_6__SCAN_IN), .A(n14595), .ZN(
        n14596) );
  OAI21_X1 U16281 ( .B1(n14640), .B2(n14682), .A(n14596), .ZN(n14597) );
  INV_X1 U16282 ( .A(n14597), .ZN(n14603) );
  INV_X1 U16283 ( .A(n14598), .ZN(n14599) );
  OAI211_X1 U16284 ( .C1(n14682), .C2(n14600), .A(n14599), .B(n14617), .ZN(
        n14681) );
  INV_X1 U16285 ( .A(n14681), .ZN(n14601) );
  AOI22_X1 U16286 ( .A1(n14686), .A2(n14645), .B1(n14644), .B2(n14601), .ZN(
        n14602) );
  OAI211_X1 U16287 ( .C1(n14648), .C2(n14683), .A(n14603), .B(n14602), .ZN(
        P1_U3287) );
  XNOR2_X1 U16288 ( .A(n14604), .B(n14605), .ZN(n14663) );
  XNOR2_X1 U16289 ( .A(n14606), .B(n14605), .ZN(n14609) );
  OAI21_X1 U16290 ( .B1(n14609), .B2(n14608), .A(n14607), .ZN(n14610) );
  AOI21_X1 U16291 ( .B1(n14712), .B2(n14663), .A(n14610), .ZN(n14660) );
  NOR2_X1 U16292 ( .A1(n14612), .A2(n14611), .ZN(n14613) );
  AOI21_X1 U16293 ( .B1(n14648), .B2(P1_REG2_REG_2__SCAN_IN), .A(n14613), .ZN(
        n14614) );
  OAI21_X1 U16294 ( .B1(n14640), .B2(n14659), .A(n14614), .ZN(n14615) );
  INV_X1 U16295 ( .A(n14615), .ZN(n14622) );
  INV_X1 U16296 ( .A(n14627), .ZN(n14619) );
  INV_X1 U16297 ( .A(n14616), .ZN(n14618) );
  OAI211_X1 U16298 ( .C1(n14659), .C2(n14619), .A(n14618), .B(n14617), .ZN(
        n14658) );
  INV_X1 U16299 ( .A(n14658), .ZN(n14620) );
  AOI22_X1 U16300 ( .A1(n14663), .A2(n14645), .B1(n14644), .B2(n14620), .ZN(
        n14621) );
  OAI211_X1 U16301 ( .C1(n14648), .C2(n14660), .A(n14622), .B(n14621), .ZN(
        P1_U3291) );
  XNOR2_X1 U16302 ( .A(n14624), .B(n14623), .ZN(n14656) );
  INV_X1 U16303 ( .A(n14624), .ZN(n14626) );
  OAI21_X1 U16304 ( .B1(n14626), .B2(n14625), .A(n14630), .ZN(n14634) );
  OAI21_X1 U16305 ( .B1(n14652), .B2(n14628), .A(n14627), .ZN(n14642) );
  XNOR2_X1 U16306 ( .A(n14642), .B(n14629), .ZN(n14631) );
  AOI21_X1 U16307 ( .B1(n14631), .B2(n14630), .A(n10017), .ZN(n14632) );
  AOI21_X1 U16308 ( .B1(n14634), .B2(n14633), .A(n14632), .ZN(n14635) );
  AOI211_X1 U16309 ( .C1(n14712), .C2(n14656), .A(n14636), .B(n14635), .ZN(
        n14653) );
  AOI22_X1 U16310 ( .A1(n14638), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n14637), .ZN(n14639) );
  OAI21_X1 U16311 ( .B1(n14640), .B2(n14652), .A(n14639), .ZN(n14641) );
  INV_X1 U16312 ( .A(n14641), .ZN(n14647) );
  OR2_X1 U16313 ( .A1(n14642), .A2(n14675), .ZN(n14651) );
  INV_X1 U16314 ( .A(n14651), .ZN(n14643) );
  AOI22_X1 U16315 ( .A1(n14645), .A2(n14656), .B1(n14644), .B2(n14643), .ZN(
        n14646) );
  OAI211_X1 U16316 ( .C1(n14648), .C2(n14653), .A(n14647), .B(n14646), .ZN(
        P1_U3292) );
  AND2_X1 U16317 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14650), .ZN(P1_U3294) );
  AND2_X1 U16318 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14650), .ZN(P1_U3295) );
  AND2_X1 U16319 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14650), .ZN(P1_U3296) );
  AND2_X1 U16320 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14650), .ZN(P1_U3297) );
  AND2_X1 U16321 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14650), .ZN(P1_U3298) );
  AND2_X1 U16322 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14650), .ZN(P1_U3299) );
  AND2_X1 U16323 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14650), .ZN(P1_U3300) );
  AND2_X1 U16324 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14650), .ZN(P1_U3301) );
  INV_X1 U16325 ( .A(n14650), .ZN(n14649) );
  INV_X1 U16326 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15234) );
  NOR2_X1 U16327 ( .A1(n14649), .A2(n15234), .ZN(P1_U3302) );
  AND2_X1 U16328 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14650), .ZN(P1_U3303) );
  AND2_X1 U16329 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14650), .ZN(P1_U3304) );
  AND2_X1 U16330 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14650), .ZN(P1_U3305) );
  AND2_X1 U16331 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14650), .ZN(P1_U3306) );
  AND2_X1 U16332 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14650), .ZN(P1_U3307) );
  AND2_X1 U16333 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14650), .ZN(P1_U3308) );
  AND2_X1 U16334 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14650), .ZN(P1_U3309) );
  AND2_X1 U16335 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14650), .ZN(P1_U3310) );
  AND2_X1 U16336 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14650), .ZN(P1_U3311) );
  AND2_X1 U16337 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14650), .ZN(P1_U3312) );
  AND2_X1 U16338 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14650), .ZN(P1_U3313) );
  AND2_X1 U16339 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14650), .ZN(P1_U3314) );
  AND2_X1 U16340 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14650), .ZN(P1_U3315) );
  AND2_X1 U16341 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14650), .ZN(P1_U3316) );
  AND2_X1 U16342 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14650), .ZN(P1_U3317) );
  AND2_X1 U16343 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14650), .ZN(P1_U3318) );
  AND2_X1 U16344 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14650), .ZN(P1_U3319) );
  AND2_X1 U16345 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14650), .ZN(P1_U3320) );
  AND2_X1 U16346 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14650), .ZN(P1_U3321) );
  AND2_X1 U16347 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14650), .ZN(P1_U3322) );
  AND2_X1 U16348 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14650), .ZN(P1_U3323) );
  INV_X1 U16349 ( .A(n14709), .ZN(n14687) );
  OAI21_X1 U16350 ( .B1(n14652), .B2(n14717), .A(n14651), .ZN(n14655) );
  INV_X1 U16351 ( .A(n14653), .ZN(n14654) );
  AOI211_X1 U16352 ( .C1(n14687), .C2(n14656), .A(n14655), .B(n14654), .ZN(
        n14726) );
  INV_X1 U16353 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14657) );
  AOI22_X1 U16354 ( .A1(n14724), .A2(n14726), .B1(n14657), .B2(n14722), .ZN(
        P1_U3462) );
  OAI21_X1 U16355 ( .B1(n14659), .B2(n14717), .A(n14658), .ZN(n14662) );
  INV_X1 U16356 ( .A(n14660), .ZN(n14661) );
  AOI211_X1 U16357 ( .C1(n14687), .C2(n14663), .A(n14662), .B(n14661), .ZN(
        n14728) );
  INV_X1 U16358 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14664) );
  AOI22_X1 U16359 ( .A1(n14724), .A2(n14728), .B1(n14664), .B2(n14722), .ZN(
        P1_U3465) );
  OAI22_X1 U16360 ( .A1(n14665), .A2(n14675), .B1(n8301), .B2(n14717), .ZN(
        n14667) );
  AOI211_X1 U16361 ( .C1(n14714), .C2(n14668), .A(n14667), .B(n14666), .ZN(
        n14730) );
  AOI22_X1 U16362 ( .A1(n14724), .A2(n14730), .B1(n8296), .B2(n14722), .ZN(
        P1_U3468) );
  OAI21_X1 U16363 ( .B1(n14670), .B2(n14717), .A(n14669), .ZN(n14672) );
  AOI211_X1 U16364 ( .C1(n14673), .C2(n14714), .A(n14672), .B(n14671), .ZN(
        n14731) );
  AOI22_X1 U16365 ( .A1(n14724), .A2(n14731), .B1(n8306), .B2(n14722), .ZN(
        P1_U3471) );
  OAI22_X1 U16366 ( .A1(n14676), .A2(n14675), .B1(n14674), .B2(n14717), .ZN(
        n14678) );
  AOI211_X1 U16367 ( .C1(n14687), .C2(n14679), .A(n14678), .B(n14677), .ZN(
        n14733) );
  INV_X1 U16368 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14680) );
  AOI22_X1 U16369 ( .A1(n14724), .A2(n14733), .B1(n14680), .B2(n14722), .ZN(
        P1_U3474) );
  OAI21_X1 U16370 ( .B1(n14682), .B2(n14717), .A(n14681), .ZN(n14685) );
  INV_X1 U16371 ( .A(n14683), .ZN(n14684) );
  AOI211_X1 U16372 ( .C1(n14687), .C2(n14686), .A(n14685), .B(n14684), .ZN(
        n14734) );
  INV_X1 U16373 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14688) );
  AOI22_X1 U16374 ( .A1(n14724), .A2(n14734), .B1(n14688), .B2(n14722), .ZN(
        P1_U3477) );
  AOI21_X1 U16375 ( .B1(n14709), .B2(n14690), .A(n14689), .ZN(n14695) );
  OAI21_X1 U16376 ( .B1(n14692), .B2(n14717), .A(n14691), .ZN(n14693) );
  NOR3_X1 U16377 ( .A1(n14695), .A2(n14694), .A3(n14693), .ZN(n14735) );
  INV_X1 U16378 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14696) );
  AOI22_X1 U16379 ( .A1(n14724), .A2(n14735), .B1(n14696), .B2(n14722), .ZN(
        P1_U3480) );
  OAI211_X1 U16380 ( .C1(n14699), .C2(n14717), .A(n14698), .B(n14697), .ZN(
        n14700) );
  AOI21_X1 U16381 ( .B1(n14701), .B2(n14714), .A(n14700), .ZN(n14736) );
  INV_X1 U16382 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14702) );
  AOI22_X1 U16383 ( .A1(n14724), .A2(n14736), .B1(n14702), .B2(n14722), .ZN(
        P1_U3483) );
  INV_X1 U16384 ( .A(n14708), .ZN(n14711) );
  AOI211_X1 U16385 ( .C1(n14706), .C2(n14705), .A(n14704), .B(n14703), .ZN(
        n14707) );
  OAI21_X1 U16386 ( .B1(n14709), .B2(n14708), .A(n14707), .ZN(n14710) );
  AOI21_X1 U16387 ( .B1(n14712), .B2(n14711), .A(n14710), .ZN(n14737) );
  INV_X1 U16388 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14713) );
  AOI22_X1 U16389 ( .A1(n14724), .A2(n14737), .B1(n14713), .B2(n14722), .ZN(
        P1_U3486) );
  AND2_X1 U16390 ( .A1(n14715), .A2(n14714), .ZN(n14721) );
  OAI21_X1 U16391 ( .B1(n14718), .B2(n14717), .A(n14716), .ZN(n14719) );
  NOR3_X1 U16392 ( .A1(n14721), .A2(n14720), .A3(n14719), .ZN(n14739) );
  INV_X1 U16393 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14723) );
  AOI22_X1 U16394 ( .A1(n14724), .A2(n14739), .B1(n14723), .B2(n14722), .ZN(
        P1_U3489) );
  AOI22_X1 U16395 ( .A1(n14740), .A2(n14726), .B1(n14725), .B2(n14738), .ZN(
        P1_U3529) );
  AOI22_X1 U16396 ( .A1(n14740), .A2(n14728), .B1(n14727), .B2(n14738), .ZN(
        P1_U3530) );
  INV_X1 U16397 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n14729) );
  AOI22_X1 U16398 ( .A1(n14740), .A2(n14730), .B1(n14729), .B2(n14738), .ZN(
        P1_U3531) );
  AOI22_X1 U16399 ( .A1(n14740), .A2(n14731), .B1(n15265), .B2(n14738), .ZN(
        P1_U3532) );
  INV_X1 U16400 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14732) );
  AOI22_X1 U16401 ( .A1(n14740), .A2(n14733), .B1(n14732), .B2(n14738), .ZN(
        P1_U3533) );
  AOI22_X1 U16402 ( .A1(n14740), .A2(n14734), .B1(n10042), .B2(n14738), .ZN(
        P1_U3534) );
  AOI22_X1 U16403 ( .A1(n14740), .A2(n14735), .B1(n10253), .B2(n14738), .ZN(
        P1_U3535) );
  AOI22_X1 U16404 ( .A1(n14740), .A2(n14736), .B1(n10426), .B2(n14738), .ZN(
        P1_U3536) );
  AOI22_X1 U16405 ( .A1(n14740), .A2(n14737), .B1(n10727), .B2(n14738), .ZN(
        P1_U3537) );
  AOI22_X1 U16406 ( .A1(n14740), .A2(n14739), .B1(n10985), .B2(n14738), .ZN(
        P1_U3538) );
  NOR2_X1 U16407 ( .A1(n14819), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16408 ( .A1(n14819), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14753) );
  OAI211_X1 U16409 ( .C1(n14743), .C2(n14742), .A(n14784), .B(n14741), .ZN(
        n14744) );
  OAI21_X1 U16410 ( .B1(n14827), .B2(n14745), .A(n14744), .ZN(n14746) );
  INV_X1 U16411 ( .A(n14746), .ZN(n14752) );
  OAI21_X1 U16412 ( .B1(n14748), .B2(n6915), .A(n14747), .ZN(n14749) );
  NAND3_X1 U16413 ( .A1(n14805), .A2(n14750), .A3(n14749), .ZN(n14751) );
  NAND3_X1 U16414 ( .A1(n14753), .A2(n14752), .A3(n14751), .ZN(P2_U3215) );
  AOI22_X1 U16415 ( .A1(n14819), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14765) );
  OAI211_X1 U16416 ( .C1(n14756), .C2(n14755), .A(n14784), .B(n14754), .ZN(
        n14757) );
  OAI21_X1 U16417 ( .B1(n14827), .B2(n14758), .A(n14757), .ZN(n14759) );
  INV_X1 U16418 ( .A(n14759), .ZN(n14764) );
  XOR2_X1 U16419 ( .A(n14761), .B(n14760), .Z(n14762) );
  NAND2_X1 U16420 ( .A1(n14805), .A2(n14762), .ZN(n14763) );
  NAND3_X1 U16421 ( .A1(n14765), .A2(n14764), .A3(n14763), .ZN(P2_U3216) );
  INV_X1 U16422 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14779) );
  OAI211_X1 U16423 ( .C1(n14768), .C2(n14767), .A(n14784), .B(n14766), .ZN(
        n14770) );
  OAI211_X1 U16424 ( .C1(n14772), .C2(n14771), .A(n14770), .B(n14769), .ZN(
        n14773) );
  INV_X1 U16425 ( .A(n14773), .ZN(n14778) );
  OAI211_X1 U16426 ( .C1(n14776), .C2(n14775), .A(n14805), .B(n14774), .ZN(
        n14777) );
  OAI211_X1 U16427 ( .C1(n14811), .C2(n14779), .A(n14778), .B(n14777), .ZN(
        P2_U3218) );
  NAND2_X1 U16428 ( .A1(n14781), .A2(n14780), .ZN(n14782) );
  NAND2_X1 U16429 ( .A1(n14783), .A2(n14782), .ZN(n14785) );
  NAND2_X1 U16430 ( .A1(n14785), .A2(n14784), .ZN(n14791) );
  OAI21_X1 U16431 ( .B1(n14788), .B2(n14787), .A(n14786), .ZN(n14789) );
  NAND2_X1 U16432 ( .A1(n14789), .A2(n14805), .ZN(n14790) );
  OAI211_X1 U16433 ( .C1(n14827), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        n14793) );
  INV_X1 U16434 ( .A(n14793), .ZN(n14795) );
  OAI211_X1 U16435 ( .C1(n14796), .C2(n14811), .A(n14795), .B(n14794), .ZN(
        P2_U3223) );
  INV_X1 U16436 ( .A(n14797), .ZN(n14802) );
  AOI211_X1 U16437 ( .C1(n14800), .C2(n14799), .A(n14798), .B(n14813), .ZN(
        n14801) );
  AOI211_X1 U16438 ( .C1(n14804), .C2(n14803), .A(n14802), .B(n14801), .ZN(
        n14809) );
  OAI211_X1 U16439 ( .C1(n14807), .C2(P2_REG2_REG_14__SCAN_IN), .A(n14806), 
        .B(n14805), .ZN(n14808) );
  OAI211_X1 U16440 ( .C1(n14811), .C2(n14810), .A(n14809), .B(n14808), .ZN(
        P2_U3228) );
  INV_X1 U16441 ( .A(n14812), .ZN(n14818) );
  AOI211_X1 U16442 ( .C1(n14816), .C2(n14815), .A(n14814), .B(n14813), .ZN(
        n14817) );
  AOI211_X1 U16443 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n14819), .A(n14818), 
        .B(n14817), .ZN(n14825) );
  AOI21_X1 U16444 ( .B1(n14821), .B2(P2_REG2_REG_18__SCAN_IN), .A(n14820), 
        .ZN(n14822) );
  OR2_X1 U16445 ( .A1(n14823), .A2(n14822), .ZN(n14824) );
  OAI211_X1 U16446 ( .C1(n14827), .C2(n14826), .A(n14825), .B(n14824), .ZN(
        P2_U3232) );
  AND2_X1 U16447 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14829), .ZN(P2_U3266) );
  AND2_X1 U16448 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14829), .ZN(P2_U3267) );
  AND2_X1 U16449 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14829), .ZN(P2_U3268) );
  AND2_X1 U16450 ( .A1(n14829), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3269) );
  AND2_X1 U16451 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14829), .ZN(P2_U3270) );
  AND2_X1 U16452 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14829), .ZN(P2_U3271) );
  AND2_X1 U16453 ( .A1(n14829), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3272) );
  AND2_X1 U16454 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14829), .ZN(P2_U3273) );
  AND2_X1 U16455 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14829), .ZN(P2_U3274) );
  AND2_X1 U16456 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14829), .ZN(P2_U3275) );
  AND2_X1 U16457 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14829), .ZN(P2_U3276) );
  AND2_X1 U16458 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14829), .ZN(P2_U3277) );
  AND2_X1 U16459 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14829), .ZN(P2_U3278) );
  AND2_X1 U16460 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14829), .ZN(P2_U3279) );
  AND2_X1 U16461 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14829), .ZN(P2_U3280) );
  AND2_X1 U16462 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14829), .ZN(P2_U3281) );
  AND2_X1 U16463 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14829), .ZN(P2_U3282) );
  AND2_X1 U16464 ( .A1(n14829), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3283) );
  AND2_X1 U16465 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14829), .ZN(P2_U3284) );
  AND2_X1 U16466 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14829), .ZN(P2_U3285) );
  AND2_X1 U16467 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14829), .ZN(P2_U3286) );
  AND2_X1 U16468 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14829), .ZN(P2_U3287) );
  AND2_X1 U16469 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14829), .ZN(P2_U3288) );
  AND2_X1 U16470 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14829), .ZN(P2_U3289) );
  AND2_X1 U16471 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14829), .ZN(P2_U3290) );
  AND2_X1 U16472 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14829), .ZN(P2_U3291) );
  AND2_X1 U16473 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14829), .ZN(P2_U3292) );
  AND2_X1 U16474 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14829), .ZN(P2_U3293) );
  AND2_X1 U16475 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14829), .ZN(P2_U3294) );
  AND2_X1 U16476 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14829), .ZN(P2_U3295) );
  INV_X1 U16477 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14830) );
  AOI22_X1 U16478 ( .A1(n14835), .A2(n14831), .B1(n14830), .B2(n14832), .ZN(
        P2_U3416) );
  INV_X1 U16479 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14833) );
  AOI22_X1 U16480 ( .A1(n14835), .A2(n14834), .B1(n14833), .B2(n14832), .ZN(
        P2_U3417) );
  OAI211_X1 U16481 ( .C1(n14895), .C2(n14838), .A(n14837), .B(n14836), .ZN(
        n14839) );
  INV_X1 U16482 ( .A(n14839), .ZN(n14901) );
  INV_X1 U16483 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14840) );
  AOI22_X1 U16484 ( .A1(n15282), .A2(n14901), .B1(n14840), .B2(n14899), .ZN(
        P2_U3430) );
  INV_X1 U16485 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14841) );
  AOI22_X1 U16486 ( .A1(n15282), .A2(n14842), .B1(n14841), .B2(n14899), .ZN(
        P2_U3433) );
  OAI21_X1 U16487 ( .B1(n14876), .B2(n14844), .A(n14843), .ZN(n14848) );
  INV_X1 U16488 ( .A(n14849), .ZN(n14846) );
  OAI21_X1 U16489 ( .B1(n14846), .B2(n10336), .A(n14845), .ZN(n14847) );
  AOI211_X1 U16490 ( .C1(n14873), .C2(n14849), .A(n14848), .B(n14847), .ZN(
        n14902) );
  INV_X1 U16491 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14850) );
  AOI22_X1 U16492 ( .A1(n15282), .A2(n14902), .B1(n14850), .B2(n14899), .ZN(
        P2_U3436) );
  NOR2_X1 U16493 ( .A1(n14852), .A2(n14851), .ZN(n14856) );
  OAI21_X1 U16494 ( .B1(n10566), .B2(n14876), .A(n14853), .ZN(n14854) );
  NOR4_X1 U16495 ( .A1(n14857), .A2(n14856), .A3(n14855), .A4(n14854), .ZN(
        n14903) );
  INV_X1 U16496 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n15264) );
  AOI22_X1 U16497 ( .A1(n15282), .A2(n14903), .B1(n15264), .B2(n14899), .ZN(
        P2_U3439) );
  NAND2_X1 U16498 ( .A1(n14863), .A2(n14873), .ZN(n14859) );
  OAI211_X1 U16499 ( .C1(n14860), .C2(n14876), .A(n14859), .B(n14858), .ZN(
        n14861) );
  AOI211_X1 U16500 ( .C1(n14890), .C2(n14863), .A(n14862), .B(n14861), .ZN(
        n14904) );
  INV_X1 U16501 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14864) );
  AOI22_X1 U16502 ( .A1(n15282), .A2(n14904), .B1(n14864), .B2(n14899), .ZN(
        P2_U3442) );
  INV_X1 U16503 ( .A(n14866), .ZN(n14872) );
  OAI21_X1 U16504 ( .B1(n10336), .B2(n14866), .A(n14865), .ZN(n14871) );
  INV_X1 U16505 ( .A(n14867), .ZN(n14868) );
  OAI21_X1 U16506 ( .B1(n14869), .B2(n14876), .A(n14868), .ZN(n14870) );
  AOI211_X1 U16507 ( .C1(n14873), .C2(n14872), .A(n14871), .B(n14870), .ZN(
        n14905) );
  INV_X1 U16508 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14874) );
  AOI22_X1 U16509 ( .A1(n15282), .A2(n14905), .B1(n14874), .B2(n14899), .ZN(
        P2_U3445) );
  OAI21_X1 U16510 ( .B1(n14877), .B2(n14876), .A(n14875), .ZN(n14879) );
  AOI211_X1 U16511 ( .C1(n14881), .C2(n14880), .A(n14879), .B(n14878), .ZN(
        n14907) );
  INV_X1 U16512 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14882) );
  AOI22_X1 U16513 ( .A1(n15282), .A2(n14907), .B1(n14882), .B2(n14899), .ZN(
        P2_U3451) );
  INV_X1 U16514 ( .A(n14887), .ZN(n14889) );
  AOI211_X1 U16515 ( .C1(n14885), .C2(n14891), .A(n14884), .B(n14883), .ZN(
        n14886) );
  OAI21_X1 U16516 ( .B1(n14887), .B2(n14895), .A(n14886), .ZN(n14888) );
  AOI21_X1 U16517 ( .B1(n14890), .B2(n14889), .A(n14888), .ZN(n14909) );
  INV_X1 U16518 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15222) );
  AOI22_X1 U16519 ( .A1(n15282), .A2(n14909), .B1(n15222), .B2(n14899), .ZN(
        P2_U3454) );
  NAND2_X1 U16520 ( .A1(n14892), .A2(n14891), .ZN(n14893) );
  OAI211_X1 U16521 ( .C1(n14896), .C2(n14895), .A(n14894), .B(n14893), .ZN(
        n14897) );
  NOR2_X1 U16522 ( .A1(n14898), .A2(n14897), .ZN(n14911) );
  INV_X1 U16523 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14900) );
  AOI22_X1 U16524 ( .A1(n15282), .A2(n14911), .B1(n14900), .B2(n14899), .ZN(
        P2_U3460) );
  AOI22_X1 U16525 ( .A1(n14912), .A2(n14901), .B1(n10174), .B2(n14910), .ZN(
        P2_U3499) );
  AOI22_X1 U16526 ( .A1(n14912), .A2(n14902), .B1(n10076), .B2(n14910), .ZN(
        P2_U3501) );
  AOI22_X1 U16527 ( .A1(n14912), .A2(n14903), .B1(n10082), .B2(n14910), .ZN(
        P2_U3502) );
  AOI22_X1 U16528 ( .A1(n14912), .A2(n14904), .B1(n10085), .B2(n14910), .ZN(
        P2_U3503) );
  AOI22_X1 U16529 ( .A1(n14912), .A2(n14905), .B1(n10075), .B2(n14910), .ZN(
        P2_U3504) );
  AOI22_X1 U16530 ( .A1(n14912), .A2(n14907), .B1(n14906), .B2(n14910), .ZN(
        P2_U3506) );
  AOI22_X1 U16531 ( .A1(n14912), .A2(n14909), .B1(n14908), .B2(n14910), .ZN(
        P2_U3507) );
  AOI22_X1 U16532 ( .A1(n14912), .A2(n14911), .B1(n10208), .B2(n14910), .ZN(
        P2_U3509) );
  NOR2_X1 U16533 ( .A1(P3_U3897), .A2(n14921), .ZN(P3_U3150) );
  INV_X1 U16534 ( .A(n14913), .ZN(n14915) );
  AOI222_X1 U16535 ( .A1(n14918), .A2(n14917), .B1(n7333), .B2(n14916), .C1(
        n14915), .C2(n14914), .ZN(n14919) );
  OAI21_X1 U16536 ( .B1(n14920), .B2(n10288), .A(n14919), .ZN(P3_U3172) );
  AOI22_X1 U16537 ( .A1(n14948), .A2(P3_IR_REG_0__SCAN_IN), .B1(n14921), .B2(
        P3_ADDR_REG_0__SCAN_IN), .ZN(n14930) );
  NOR3_X1 U16538 ( .A1(n14924), .A2(n14923), .A3(n14922), .ZN(n14928) );
  AOI21_X1 U16539 ( .B1(n15207), .B2(n14926), .A(n14925), .ZN(n14927) );
  OR2_X1 U16540 ( .A1(n14928), .A2(n14927), .ZN(n14929) );
  OAI211_X1 U16541 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n10288), .A(n14930), .B(
        n14929), .ZN(P3_U3182) );
  AOI21_X1 U16542 ( .B1(n14933), .B2(n14932), .A(n14931), .ZN(n14939) );
  AOI21_X1 U16543 ( .B1(n14936), .B2(n14935), .A(n14934), .ZN(n14938) );
  OAI22_X1 U16544 ( .A1(n14940), .A2(n14939), .B1(n14938), .B2(n14937), .ZN(
        n14946) );
  XOR2_X1 U16545 ( .A(n14942), .B(n14941), .Z(n14944) );
  NOR2_X1 U16546 ( .A1(n14944), .A2(n14943), .ZN(n14945) );
  AOI211_X1 U16547 ( .C1(n14948), .C2(n14947), .A(n14946), .B(n14945), .ZN(
        n14950) );
  OAI211_X1 U16548 ( .C1(n14952), .C2(n14951), .A(n14950), .B(n14949), .ZN(
        P3_U3190) );
  INV_X1 U16549 ( .A(n14953), .ZN(n14956) );
  OAI21_X1 U16550 ( .B1(n14956), .B2(n14955), .A(n14954), .ZN(n14960) );
  OAI22_X1 U16551 ( .A1(n14958), .A2(n14957), .B1(n11058), .B2(n15050), .ZN(
        n14959) );
  AOI21_X1 U16552 ( .B1(n14960), .B2(n15050), .A(n14959), .ZN(n14961) );
  OAI21_X1 U16553 ( .B1(n14962), .B2(n15012), .A(n14961), .ZN(P3_U3224) );
  XNOR2_X1 U16554 ( .A(n14964), .B(n14963), .ZN(n14972) );
  INV_X1 U16555 ( .A(n14972), .ZN(n15075) );
  XNOR2_X1 U16556 ( .A(n14966), .B(n14965), .ZN(n14967) );
  NAND2_X1 U16557 ( .A1(n14967), .A2(n15039), .ZN(n14971) );
  AOI22_X1 U16558 ( .A1(n14969), .A2(n15034), .B1(n15035), .B2(n14968), .ZN(
        n14970) );
  OAI211_X1 U16559 ( .C1(n15043), .C2(n14972), .A(n14971), .B(n14970), .ZN(
        n15073) );
  AOI21_X1 U16560 ( .B1(n14993), .B2(n15075), .A(n15073), .ZN(n14977) );
  NOR2_X1 U16561 ( .A1(n14973), .A2(n15030), .ZN(n15074) );
  AOI22_X1 U16562 ( .A1(n15074), .A2(n15000), .B1(n15046), .B2(n14974), .ZN(
        n14975) );
  OAI221_X1 U16563 ( .B1(n14334), .B2(n14977), .C1(n15050), .C2(n14976), .A(
        n14975), .ZN(P3_U3226) );
  XOR2_X1 U16564 ( .A(n14978), .B(n14981), .Z(n14992) );
  INV_X1 U16565 ( .A(n14992), .ZN(n15069) );
  NAND2_X1 U16566 ( .A1(n15003), .A2(n15001), .ZN(n14983) );
  AND2_X1 U16567 ( .A1(n14983), .A2(n14980), .ZN(n14986) );
  INV_X1 U16568 ( .A(n14981), .ZN(n14985) );
  NAND2_X1 U16569 ( .A1(n14983), .A2(n14982), .ZN(n14984) );
  OAI21_X1 U16570 ( .B1(n14986), .B2(n14985), .A(n14984), .ZN(n14990) );
  OAI22_X1 U16571 ( .A1(n14988), .A2(n15019), .B1(n14987), .B2(n15017), .ZN(
        n14989) );
  AOI21_X1 U16572 ( .B1(n14990), .B2(n15039), .A(n14989), .ZN(n14991) );
  OAI21_X1 U16573 ( .B1(n15043), .B2(n14992), .A(n14991), .ZN(n15067) );
  AOI21_X1 U16574 ( .B1(n14993), .B2(n15069), .A(n15067), .ZN(n14998) );
  AND2_X1 U16575 ( .A1(n14994), .A2(n15023), .ZN(n15068) );
  AOI22_X1 U16576 ( .A1(n15000), .A2(n15068), .B1(n15046), .B2(n14995), .ZN(
        n14996) );
  OAI221_X1 U16577 ( .B1(n14334), .B2(n14998), .C1(n15050), .C2(n14997), .A(
        n14996), .ZN(P3_U3228) );
  AND2_X1 U16578 ( .A1(n14999), .A2(n15023), .ZN(n15065) );
  AOI22_X1 U16579 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n14334), .B1(n15000), 
        .B2(n15065), .ZN(n15011) );
  XNOR2_X1 U16580 ( .A(n15002), .B(n15001), .ZN(n15063) );
  XNOR2_X1 U16581 ( .A(n15004), .B(n15003), .ZN(n15007) );
  OAI22_X1 U16582 ( .A1(n15005), .A2(n15017), .B1(n15018), .B2(n15019), .ZN(
        n15006) );
  AOI21_X1 U16583 ( .B1(n15007), .B2(n15039), .A(n15006), .ZN(n15008) );
  OAI21_X1 U16584 ( .B1(n15043), .B2(n15063), .A(n15008), .ZN(n15064) );
  NOR2_X1 U16585 ( .A1(n15063), .A2(n15026), .ZN(n15009) );
  OAI21_X1 U16586 ( .B1(n15064), .B2(n15009), .A(n15050), .ZN(n15010) );
  OAI211_X1 U16587 ( .C1(n15013), .C2(n15012), .A(n15011), .B(n15010), .ZN(
        P3_U3229) );
  OAI21_X1 U16588 ( .B1(n15016), .B2(n15015), .A(n15014), .ZN(n15021) );
  OAI22_X1 U16589 ( .A1(n8829), .A2(n15019), .B1(n15018), .B2(n15017), .ZN(
        n15020) );
  AOI21_X1 U16590 ( .B1(n15021), .B2(n15039), .A(n15020), .ZN(n15022) );
  OAI21_X1 U16591 ( .B1(n15043), .B2(n15056), .A(n15022), .ZN(n15057) );
  AND2_X1 U16592 ( .A1(n15024), .A2(n15023), .ZN(n15058) );
  AOI22_X1 U16593 ( .A1(n15058), .A2(n15044), .B1(P3_REG3_REG_2__SCAN_IN), 
        .B2(n15046), .ZN(n15025) );
  OAI21_X1 U16594 ( .B1(n15056), .B2(n15026), .A(n15025), .ZN(n15027) );
  NOR2_X1 U16595 ( .A1(n15057), .A2(n15027), .ZN(n15028) );
  AOI22_X1 U16596 ( .A1(n14334), .A2(n15029), .B1(n15028), .B2(n15050), .ZN(
        P3_U3231) );
  NOR2_X1 U16597 ( .A1(n15031), .A2(n15030), .ZN(n15054) );
  XNOR2_X1 U16598 ( .A(n15038), .B(n15032), .ZN(n15045) );
  AOI22_X1 U16599 ( .A1(n15036), .A2(n15035), .B1(n15034), .B2(n15033), .ZN(
        n15042) );
  XNOR2_X1 U16600 ( .A(n15038), .B(n15037), .ZN(n15040) );
  NAND2_X1 U16601 ( .A1(n15040), .A2(n15039), .ZN(n15041) );
  OAI211_X1 U16602 ( .C1(n15045), .C2(n15043), .A(n15042), .B(n15041), .ZN(
        n15053) );
  AOI21_X1 U16603 ( .B1(n15054), .B2(n15044), .A(n15053), .ZN(n15051) );
  INV_X1 U16604 ( .A(n15045), .ZN(n15055) );
  AOI22_X1 U16605 ( .A1(n15055), .A2(n15047), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15046), .ZN(n15048) );
  OAI221_X1 U16606 ( .B1(n14334), .B2(n15051), .C1(n15050), .C2(n15049), .A(
        n15048), .ZN(P3_U3232) );
  AOI211_X1 U16607 ( .C1(n15079), .C2(n15055), .A(n15054), .B(n15053), .ZN(
        n15083) );
  AOI22_X1 U16608 ( .A1(n15081), .A2(n15083), .B1(n8803), .B2(n15080), .ZN(
        P3_U3393) );
  INV_X1 U16609 ( .A(n15056), .ZN(n15059) );
  AOI211_X1 U16610 ( .C1(n15059), .C2(n15079), .A(n15058), .B(n15057), .ZN(
        n15084) );
  AOI22_X1 U16611 ( .A1(n15081), .A2(n15084), .B1(n8798), .B2(n15080), .ZN(
        P3_U3396) );
  AOI211_X1 U16612 ( .C1(n15079), .C2(n15062), .A(n15061), .B(n15060), .ZN(
        n15086) );
  AOI22_X1 U16613 ( .A1(n15081), .A2(n15086), .B1(n8832), .B2(n15080), .ZN(
        P3_U3399) );
  INV_X1 U16614 ( .A(n15063), .ZN(n15066) );
  AOI211_X1 U16615 ( .C1(n15066), .C2(n15079), .A(n15065), .B(n15064), .ZN(
        n15088) );
  AOI22_X1 U16616 ( .A1(n15081), .A2(n15088), .B1(n8848), .B2(n15080), .ZN(
        P3_U3402) );
  AOI211_X1 U16617 ( .C1(n15069), .C2(n15079), .A(n15068), .B(n15067), .ZN(
        n15090) );
  AOI22_X1 U16618 ( .A1(n15081), .A2(n15090), .B1(n8870), .B2(n15080), .ZN(
        P3_U3405) );
  AOI211_X1 U16619 ( .C1(n15079), .C2(n15072), .A(n15071), .B(n15070), .ZN(
        n15092) );
  AOI22_X1 U16620 ( .A1(n15081), .A2(n15092), .B1(n8880), .B2(n15080), .ZN(
        P3_U3408) );
  AOI211_X1 U16621 ( .C1(n15075), .C2(n15079), .A(n15074), .B(n15073), .ZN(
        n15093) );
  AOI22_X1 U16622 ( .A1(n15081), .A2(n15093), .B1(n8896), .B2(n15080), .ZN(
        P3_U3411) );
  AOI211_X1 U16623 ( .C1(n15079), .C2(n15078), .A(n15077), .B(n15076), .ZN(
        n15095) );
  AOI22_X1 U16624 ( .A1(n15081), .A2(n15095), .B1(n8909), .B2(n15080), .ZN(
        P3_U3414) );
  AOI22_X1 U16625 ( .A1(n15096), .A2(n15083), .B1(n15082), .B2(n15094), .ZN(
        P3_U3460) );
  AOI22_X1 U16626 ( .A1(n15096), .A2(n15084), .B1(n15261), .B2(n15094), .ZN(
        P3_U3461) );
  AOI22_X1 U16627 ( .A1(n15096), .A2(n15086), .B1(n15085), .B2(n15094), .ZN(
        P3_U3462) );
  INV_X1 U16628 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15087) );
  AOI22_X1 U16629 ( .A1(n15096), .A2(n15088), .B1(n15087), .B2(n15094), .ZN(
        P3_U3463) );
  AOI22_X1 U16630 ( .A1(n15096), .A2(n15090), .B1(n15089), .B2(n15094), .ZN(
        P3_U3464) );
  AOI22_X1 U16631 ( .A1(n15096), .A2(n15092), .B1(n15091), .B2(n15094), .ZN(
        P3_U3465) );
  AOI22_X1 U16632 ( .A1(n15096), .A2(n15093), .B1(n15098), .B2(n15094), .ZN(
        P3_U3466) );
  AOI22_X1 U16633 ( .A1(n15096), .A2(n15095), .B1(n11074), .B2(n15094), .ZN(
        P3_U3467) );
  AOI22_X1 U16634 ( .A1(n15098), .A2(keyinput87), .B1(keyinput120), .B2(n8832), 
        .ZN(n15097) );
  OAI221_X1 U16635 ( .B1(n15098), .B2(keyinput87), .C1(n8832), .C2(keyinput120), .A(n15097), .ZN(n15108) );
  INV_X1 U16636 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15100) );
  AOI22_X1 U16637 ( .A1(n9995), .A2(keyinput74), .B1(n15100), .B2(keyinput95), 
        .ZN(n15099) );
  OAI221_X1 U16638 ( .B1(n9995), .B2(keyinput74), .C1(n15100), .C2(keyinput95), 
        .A(n15099), .ZN(n15107) );
  AOI22_X1 U16639 ( .A1(n15264), .A2(keyinput65), .B1(n15225), .B2(keyinput100), .ZN(n15101) );
  OAI221_X1 U16640 ( .B1(n15264), .B2(keyinput65), .C1(n15225), .C2(
        keyinput100), .A(n15101), .ZN(n15106) );
  AOI22_X1 U16641 ( .A1(n15104), .A2(keyinput115), .B1(n15103), .B2(
        keyinput116), .ZN(n15102) );
  OAI221_X1 U16642 ( .B1(n15104), .B2(keyinput115), .C1(n15103), .C2(
        keyinput116), .A(n15102), .ZN(n15105) );
  NOR4_X1 U16643 ( .A1(n15108), .A2(n15107), .A3(n15106), .A4(n15105), .ZN(
        n15141) );
  AOI22_X1 U16644 ( .A1(P1_REG0_REG_21__SCAN_IN), .A2(keyinput112), .B1(
        P3_REG0_REG_22__SCAN_IN), .B2(keyinput82), .ZN(n15109) );
  OAI221_X1 U16645 ( .B1(P1_REG0_REG_21__SCAN_IN), .B2(keyinput112), .C1(
        P3_REG0_REG_22__SCAN_IN), .C2(keyinput82), .A(n15109), .ZN(n15116) );
  AOI22_X1 U16646 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(keyinput73), .B1(
        P3_REG2_REG_13__SCAN_IN), .B2(keyinput71), .ZN(n15110) );
  OAI221_X1 U16647 ( .B1(P2_IR_REG_16__SCAN_IN), .B2(keyinput73), .C1(
        P3_REG2_REG_13__SCAN_IN), .C2(keyinput71), .A(n15110), .ZN(n15115) );
  AOI22_X1 U16648 ( .A1(n15249), .A2(keyinput68), .B1(n15218), .B2(keyinput105), .ZN(n15111) );
  OAI221_X1 U16649 ( .B1(n15249), .B2(keyinput68), .C1(n15218), .C2(
        keyinput105), .A(n15111), .ZN(n15114) );
  AOI22_X1 U16650 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(keyinput103), .B1(n8426), 
        .B2(keyinput83), .ZN(n15112) );
  OAI221_X1 U16651 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(keyinput103), .C1(n8426), 
        .C2(keyinput83), .A(n15112), .ZN(n15113) );
  NOR4_X1 U16652 ( .A1(n15116), .A2(n15115), .A3(n15114), .A4(n15113), .ZN(
        n15140) );
  AOI22_X1 U16653 ( .A1(n7031), .A2(keyinput117), .B1(n10039), .B2(keyinput81), 
        .ZN(n15117) );
  OAI221_X1 U16654 ( .B1(n7031), .B2(keyinput117), .C1(n10039), .C2(keyinput81), .A(n15117), .ZN(n15125) );
  AOI22_X1 U16655 ( .A1(n10174), .A2(keyinput78), .B1(n15119), .B2(keyinput106), .ZN(n15118) );
  OAI221_X1 U16656 ( .B1(n10174), .B2(keyinput78), .C1(n15119), .C2(
        keyinput106), .A(n15118), .ZN(n15124) );
  AOI22_X1 U16657 ( .A1(n15252), .A2(keyinput90), .B1(n15221), .B2(keyinput67), 
        .ZN(n15120) );
  OAI221_X1 U16658 ( .B1(n15252), .B2(keyinput90), .C1(n15221), .C2(keyinput67), .A(n15120), .ZN(n15123) );
  AOI22_X1 U16659 ( .A1(n15265), .A2(keyinput101), .B1(n15251), .B2(
        keyinput113), .ZN(n15121) );
  OAI221_X1 U16660 ( .B1(n15265), .B2(keyinput101), .C1(n15251), .C2(
        keyinput113), .A(n15121), .ZN(n15122) );
  NOR4_X1 U16661 ( .A1(n15125), .A2(n15124), .A3(n15123), .A4(n15122), .ZN(
        n15139) );
  AOI22_X1 U16662 ( .A1(n15207), .A2(keyinput84), .B1(keyinput122), .B2(n15245), .ZN(n15126) );
  OAI221_X1 U16663 ( .B1(n15207), .B2(keyinput84), .C1(n15245), .C2(
        keyinput122), .A(n15126), .ZN(n15137) );
  AOI22_X1 U16664 ( .A1(n15260), .A2(keyinput104), .B1(n15128), .B2(
        keyinput119), .ZN(n15127) );
  OAI221_X1 U16665 ( .B1(n15260), .B2(keyinput104), .C1(n15128), .C2(
        keyinput119), .A(n15127), .ZN(n15136) );
  AOI22_X1 U16666 ( .A1(n15131), .A2(keyinput91), .B1(keyinput89), .B2(n15130), 
        .ZN(n15129) );
  OAI221_X1 U16667 ( .B1(n15131), .B2(keyinput91), .C1(n15130), .C2(keyinput89), .A(n15129), .ZN(n15135) );
  AOI22_X1 U16668 ( .A1(n15133), .A2(keyinput80), .B1(keyinput93), .B2(n15234), 
        .ZN(n15132) );
  OAI221_X1 U16669 ( .B1(n15133), .B2(keyinput80), .C1(n15234), .C2(keyinput93), .A(n15132), .ZN(n15134) );
  NOR4_X1 U16670 ( .A1(n15137), .A2(n15136), .A3(n15135), .A4(n15134), .ZN(
        n15138) );
  AND4_X1 U16671 ( .A1(n15141), .A2(n15140), .A3(n15139), .A4(n15138), .ZN(
        n15279) );
  OAI22_X1 U16672 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput69), .B1(
        keyinput77), .B2(P1_IR_REG_25__SCAN_IN), .ZN(n15142) );
  AOI221_X1 U16673 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput69), .C1(
        P1_IR_REG_25__SCAN_IN), .C2(keyinput77), .A(n15142), .ZN(n15149) );
  OAI22_X1 U16674 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput126), .B1(
        keyinput85), .B2(P2_REG0_REG_8__SCAN_IN), .ZN(n15143) );
  AOI221_X1 U16675 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput126), .C1(
        P2_REG0_REG_8__SCAN_IN), .C2(keyinput85), .A(n15143), .ZN(n15148) );
  OAI22_X1 U16676 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(keyinput92), .B1(
        keyinput124), .B2(P3_REG1_REG_2__SCAN_IN), .ZN(n15144) );
  AOI221_X1 U16677 ( .B1(P1_DATAO_REG_7__SCAN_IN), .B2(keyinput92), .C1(
        P3_REG1_REG_2__SCAN_IN), .C2(keyinput124), .A(n15144), .ZN(n15147) );
  OAI22_X1 U16678 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput108), .B1(
        keyinput121), .B2(P2_REG1_REG_9__SCAN_IN), .ZN(n15145) );
  AOI221_X1 U16679 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput108), .C1(
        P2_REG1_REG_9__SCAN_IN), .C2(keyinput121), .A(n15145), .ZN(n15146) );
  NAND4_X1 U16680 ( .A1(n15149), .A2(n15148), .A3(n15147), .A4(n15146), .ZN(
        n15177) );
  OAI22_X1 U16681 ( .A1(P3_ADDR_REG_19__SCAN_IN), .A2(keyinput79), .B1(
        keyinput125), .B2(SI_2_), .ZN(n15150) );
  AOI221_X1 U16682 ( .B1(P3_ADDR_REG_19__SCAN_IN), .B2(keyinput79), .C1(SI_2_), 
        .C2(keyinput125), .A(n15150), .ZN(n15157) );
  OAI22_X1 U16683 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(keyinput111), .B1(
        keyinput97), .B2(P2_REG1_REG_24__SCAN_IN), .ZN(n15151) );
  AOI221_X1 U16684 ( .B1(P3_IR_REG_2__SCAN_IN), .B2(keyinput111), .C1(
        P2_REG1_REG_24__SCAN_IN), .C2(keyinput97), .A(n15151), .ZN(n15156) );
  OAI22_X1 U16685 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(keyinput127), .B1(
        SI_31_), .B2(keyinput88), .ZN(n15152) );
  AOI221_X1 U16686 ( .B1(P2_DATAO_REG_11__SCAN_IN), .B2(keyinput127), .C1(
        keyinput88), .C2(SI_31_), .A(n15152), .ZN(n15155) );
  OAI22_X1 U16687 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(keyinput102), .B1(
        P2_IR_REG_23__SCAN_IN), .B2(keyinput114), .ZN(n15153) );
  AOI221_X1 U16688 ( .B1(P2_DATAO_REG_3__SCAN_IN), .B2(keyinput102), .C1(
        keyinput114), .C2(P2_IR_REG_23__SCAN_IN), .A(n15153), .ZN(n15154) );
  NAND4_X1 U16689 ( .A1(n15157), .A2(n15156), .A3(n15155), .A4(n15154), .ZN(
        n15176) );
  OAI22_X1 U16690 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(keyinput75), .B1(
        keyinput76), .B2(SI_16_), .ZN(n15158) );
  AOI221_X1 U16691 ( .B1(P1_DATAO_REG_17__SCAN_IN), .B2(keyinput75), .C1(
        SI_16_), .C2(keyinput76), .A(n15158), .ZN(n15165) );
  OAI22_X1 U16692 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(keyinput110), .B1(
        keyinput86), .B2(P2_D_REG_28__SCAN_IN), .ZN(n15159) );
  AOI221_X1 U16693 ( .B1(P2_IR_REG_19__SCAN_IN), .B2(keyinput110), .C1(
        P2_D_REG_28__SCAN_IN), .C2(keyinput86), .A(n15159), .ZN(n15164) );
  OAI22_X1 U16694 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput96), .B1(
        P1_REG3_REG_24__SCAN_IN), .B2(keyinput123), .ZN(n15160) );
  AOI221_X1 U16695 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput96), .C1(
        keyinput123), .C2(P1_REG3_REG_24__SCAN_IN), .A(n15160), .ZN(n15163) );
  OAI22_X1 U16696 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput66), .B1(
        P1_REG2_REG_18__SCAN_IN), .B2(keyinput94), .ZN(n15161) );
  AOI221_X1 U16697 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput66), .C1(
        keyinput94), .C2(P1_REG2_REG_18__SCAN_IN), .A(n15161), .ZN(n15162) );
  NAND4_X1 U16698 ( .A1(n15165), .A2(n15164), .A3(n15163), .A4(n15162), .ZN(
        n15175) );
  OAI22_X1 U16699 ( .A1(P2_REG1_REG_1__SCAN_IN), .A2(keyinput118), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput107), .ZN(n15166) );
  AOI221_X1 U16700 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(keyinput118), .C1(
        keyinput107), .C2(P1_IR_REG_19__SCAN_IN), .A(n15166), .ZN(n15173) );
  OAI22_X1 U16701 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(keyinput98), .B1(keyinput64), .B2(P3_REG1_REG_16__SCAN_IN), .ZN(n15167) );
  AOI221_X1 U16702 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(keyinput98), .C1(
        P3_REG1_REG_16__SCAN_IN), .C2(keyinput64), .A(n15167), .ZN(n15172) );
  OAI22_X1 U16703 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(keyinput109), .B1(
        SI_25_), .B2(keyinput99), .ZN(n15168) );
  AOI221_X1 U16704 ( .B1(P2_DATAO_REG_29__SCAN_IN), .B2(keyinput109), .C1(
        keyinput99), .C2(SI_25_), .A(n15168), .ZN(n15171) );
  OAI22_X1 U16705 ( .A1(P2_REG0_REG_23__SCAN_IN), .A2(keyinput72), .B1(
        P1_REG1_REG_30__SCAN_IN), .B2(keyinput70), .ZN(n15169) );
  AOI221_X1 U16706 ( .B1(P2_REG0_REG_23__SCAN_IN), .B2(keyinput72), .C1(
        keyinput70), .C2(P1_REG1_REG_30__SCAN_IN), .A(n15169), .ZN(n15170) );
  NAND4_X1 U16707 ( .A1(n15173), .A2(n15172), .A3(n15171), .A4(n15170), .ZN(
        n15174) );
  NOR4_X1 U16708 ( .A1(n15177), .A2(n15176), .A3(n15175), .A4(n15174), .ZN(
        n15278) );
  AOI22_X1 U16709 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput52), .B1(
        P3_ADDR_REG_19__SCAN_IN), .B2(keyinput15), .ZN(n15178) );
  OAI221_X1 U16710 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput52), .C1(
        P3_ADDR_REG_19__SCAN_IN), .C2(keyinput15), .A(n15178), .ZN(n15185) );
  AOI22_X1 U16711 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(keyinput10), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(keyinput14), .ZN(n15179) );
  OAI221_X1 U16712 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(keyinput10), .C1(
        P2_REG1_REG_0__SCAN_IN), .C2(keyinput14), .A(n15179), .ZN(n15184) );
  AOI22_X1 U16713 ( .A1(P1_REG0_REG_21__SCAN_IN), .A2(keyinput48), .B1(
        P1_REG3_REG_15__SCAN_IN), .B2(keyinput51), .ZN(n15180) );
  OAI221_X1 U16714 ( .B1(P1_REG0_REG_21__SCAN_IN), .B2(keyinput48), .C1(
        P1_REG3_REG_15__SCAN_IN), .C2(keyinput51), .A(n15180), .ZN(n15183) );
  AOI22_X1 U16715 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(keyinput5), .B1(
        P3_REG1_REG_7__SCAN_IN), .B2(keyinput23), .ZN(n15181) );
  OAI221_X1 U16716 ( .B1(P1_IR_REG_20__SCAN_IN), .B2(keyinput5), .C1(
        P3_REG1_REG_7__SCAN_IN), .C2(keyinput23), .A(n15181), .ZN(n15182) );
  NOR4_X1 U16717 ( .A1(n15185), .A2(n15184), .A3(n15183), .A4(n15182), .ZN(
        n15216) );
  AOI22_X1 U16718 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput32), .B1(
        P3_IR_REG_2__SCAN_IN), .B2(keyinput47), .ZN(n15186) );
  OAI221_X1 U16719 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput32), .C1(
        P3_IR_REG_2__SCAN_IN), .C2(keyinput47), .A(n15186), .ZN(n15193) );
  AOI22_X1 U16720 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(keyinput53), .B1(
        P1_REG1_REG_30__SCAN_IN), .B2(keyinput6), .ZN(n15187) );
  OAI221_X1 U16721 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(keyinput53), .C1(
        P1_REG1_REG_30__SCAN_IN), .C2(keyinput6), .A(n15187), .ZN(n15192) );
  AOI22_X1 U16722 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(keyinput9), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(keyinput42), .ZN(n15188) );
  OAI221_X1 U16723 ( .B1(P2_IR_REG_16__SCAN_IN), .B2(keyinput9), .C1(
        P2_DATAO_REG_24__SCAN_IN), .C2(keyinput42), .A(n15188), .ZN(n15191) );
  AOI22_X1 U16724 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(keyinput57), .B1(
        P3_REG2_REG_13__SCAN_IN), .B2(keyinput7), .ZN(n15189) );
  OAI221_X1 U16725 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(keyinput57), .C1(
        P3_REG2_REG_13__SCAN_IN), .C2(keyinput7), .A(n15189), .ZN(n15190) );
  NOR4_X1 U16726 ( .A1(n15193), .A2(n15192), .A3(n15191), .A4(n15190), .ZN(
        n15215) );
  AOI22_X1 U16727 ( .A1(P2_D_REG_25__SCAN_IN), .A2(keyinput2), .B1(SI_31_), 
        .B2(keyinput24), .ZN(n15194) );
  OAI221_X1 U16728 ( .B1(P2_D_REG_25__SCAN_IN), .B2(keyinput2), .C1(SI_31_), 
        .C2(keyinput24), .A(n15194), .ZN(n15201) );
  AOI22_X1 U16729 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(keyinput50), .B1(
        P3_REG0_REG_16__SCAN_IN), .B2(keyinput27), .ZN(n15195) );
  OAI221_X1 U16730 ( .B1(P2_IR_REG_23__SCAN_IN), .B2(keyinput50), .C1(
        P3_REG0_REG_16__SCAN_IN), .C2(keyinput27), .A(n15195), .ZN(n15200) );
  AOI22_X1 U16731 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(keyinput39), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(keyinput62), .ZN(n15196) );
  OAI221_X1 U16732 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(keyinput39), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput62), .A(n15196), .ZN(n15199) );
  AOI22_X1 U16733 ( .A1(P2_D_REG_14__SCAN_IN), .A2(keyinput31), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(keyinput28), .ZN(n15197) );
  OAI221_X1 U16734 ( .B1(P2_D_REG_14__SCAN_IN), .B2(keyinput31), .C1(
        P1_DATAO_REG_7__SCAN_IN), .C2(keyinput28), .A(n15197), .ZN(n15198) );
  NOR4_X1 U16735 ( .A1(n15201), .A2(n15200), .A3(n15199), .A4(n15198), .ZN(
        n15214) );
  AOI22_X1 U16736 ( .A1(P2_REG0_REG_17__SCAN_IN), .A2(keyinput16), .B1(
        P2_D_REG_28__SCAN_IN), .B2(keyinput22), .ZN(n15202) );
  OAI221_X1 U16737 ( .B1(P2_REG0_REG_17__SCAN_IN), .B2(keyinput16), .C1(
        P2_D_REG_28__SCAN_IN), .C2(keyinput22), .A(n15202), .ZN(n15212) );
  AOI22_X1 U16738 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(keyinput17), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput43), .ZN(n15203) );
  OAI221_X1 U16739 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(keyinput17), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput43), .A(n15203), .ZN(n15211) );
  AOI22_X1 U16740 ( .A1(P1_REG0_REG_30__SCAN_IN), .A2(keyinput25), .B1(n15205), 
        .B2(keyinput45), .ZN(n15204) );
  OAI221_X1 U16741 ( .B1(P1_REG0_REG_30__SCAN_IN), .B2(keyinput25), .C1(n15205), .C2(keyinput45), .A(n15204), .ZN(n15210) );
  AOI22_X1 U16742 ( .A1(n15208), .A2(keyinput33), .B1(n15207), .B2(keyinput20), 
        .ZN(n15206) );
  OAI221_X1 U16743 ( .B1(n15208), .B2(keyinput33), .C1(n15207), .C2(keyinput20), .A(n15206), .ZN(n15209) );
  NOR4_X1 U16744 ( .A1(n15212), .A2(n15211), .A3(n15210), .A4(n15209), .ZN(
        n15213) );
  NAND4_X1 U16745 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        n15277) );
  AOI22_X1 U16746 ( .A1(n15219), .A2(keyinput11), .B1(keyinput41), .B2(n15218), 
        .ZN(n15217) );
  OAI221_X1 U16747 ( .B1(n15219), .B2(keyinput11), .C1(n15218), .C2(keyinput41), .A(n15217), .ZN(n15231) );
  AOI22_X1 U16748 ( .A1(n15222), .A2(keyinput21), .B1(n15221), .B2(keyinput3), 
        .ZN(n15220) );
  OAI221_X1 U16749 ( .B1(n15222), .B2(keyinput21), .C1(n15221), .C2(keyinput3), 
        .A(n15220), .ZN(n15230) );
  AOI22_X1 U16750 ( .A1(n15225), .A2(keyinput36), .B1(n15224), .B2(keyinput63), 
        .ZN(n15223) );
  OAI221_X1 U16751 ( .B1(n15225), .B2(keyinput36), .C1(n15224), .C2(keyinput63), .A(n15223), .ZN(n15229) );
  XNOR2_X1 U16752 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput38), .ZN(n15227)
         );
  XNOR2_X1 U16753 ( .A(P3_REG3_REG_23__SCAN_IN), .B(keyinput44), .ZN(n15226)
         );
  NAND2_X1 U16754 ( .A1(n15227), .A2(n15226), .ZN(n15228) );
  NOR4_X1 U16755 ( .A1(n15231), .A2(n15230), .A3(n15229), .A4(n15228), .ZN(
        n15275) );
  AOI22_X1 U16756 ( .A1(n15234), .A2(keyinput29), .B1(n15233), .B2(keyinput35), 
        .ZN(n15232) );
  OAI221_X1 U16757 ( .B1(n15234), .B2(keyinput29), .C1(n15233), .C2(keyinput35), .A(n15232), .ZN(n15243) );
  AOI22_X1 U16758 ( .A1(n8501), .A2(keyinput30), .B1(n15236), .B2(keyinput18), 
        .ZN(n15235) );
  OAI221_X1 U16759 ( .B1(n8501), .B2(keyinput30), .C1(n15236), .C2(keyinput18), 
        .A(n15235), .ZN(n15242) );
  XNOR2_X1 U16760 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput13), .ZN(n15240) );
  XNOR2_X1 U16761 ( .A(P3_REG1_REG_16__SCAN_IN), .B(keyinput0), .ZN(n15239) );
  XNOR2_X1 U16762 ( .A(SI_2_), .B(keyinput61), .ZN(n15238) );
  XNOR2_X1 U16763 ( .A(SI_16_), .B(keyinput12), .ZN(n15237) );
  NAND4_X1 U16764 ( .A1(n15240), .A2(n15239), .A3(n15238), .A4(n15237), .ZN(
        n15241) );
  NOR3_X1 U16765 ( .A1(n15243), .A2(n15242), .A3(n15241), .ZN(n15274) );
  AOI22_X1 U16766 ( .A1(n15246), .A2(keyinput8), .B1(n15245), .B2(keyinput58), 
        .ZN(n15244) );
  OAI221_X1 U16767 ( .B1(n15246), .B2(keyinput8), .C1(n15245), .C2(keyinput58), 
        .A(n15244), .ZN(n15258) );
  AOI22_X1 U16768 ( .A1(n15249), .A2(keyinput4), .B1(keyinput59), .B2(n15248), 
        .ZN(n15247) );
  OAI221_X1 U16769 ( .B1(n15249), .B2(keyinput4), .C1(n15248), .C2(keyinput59), 
        .A(n15247), .ZN(n15257) );
  AOI22_X1 U16770 ( .A1(n15252), .A2(keyinput26), .B1(n15251), .B2(keyinput49), 
        .ZN(n15250) );
  OAI221_X1 U16771 ( .B1(n15252), .B2(keyinput26), .C1(n15251), .C2(keyinput49), .A(n15250), .ZN(n15256) );
  XNOR2_X1 U16772 ( .A(P2_REG1_REG_21__SCAN_IN), .B(keyinput55), .ZN(n15254)
         );
  XNOR2_X1 U16773 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput46), .ZN(n15253) );
  NAND2_X1 U16774 ( .A1(n15254), .A2(n15253), .ZN(n15255) );
  NOR4_X1 U16775 ( .A1(n15258), .A2(n15257), .A3(n15256), .A4(n15255), .ZN(
        n15273) );
  AOI22_X1 U16776 ( .A1(n15261), .A2(keyinput60), .B1(keyinput40), .B2(n15260), 
        .ZN(n15259) );
  OAI221_X1 U16777 ( .B1(n15261), .B2(keyinput60), .C1(n15260), .C2(keyinput40), .A(n15259), .ZN(n15271) );
  AOI22_X1 U16778 ( .A1(n8832), .A2(keyinput56), .B1(keyinput19), .B2(n8426), 
        .ZN(n15262) );
  OAI221_X1 U16779 ( .B1(n8832), .B2(keyinput56), .C1(n8426), .C2(keyinput19), 
        .A(n15262), .ZN(n15270) );
  AOI22_X1 U16780 ( .A1(n15264), .A2(keyinput1), .B1(n8811), .B2(keyinput34), 
        .ZN(n15263) );
  OAI221_X1 U16781 ( .B1(n15264), .B2(keyinput1), .C1(n8811), .C2(keyinput34), 
        .A(n15263), .ZN(n15269) );
  XOR2_X1 U16782 ( .A(n15265), .B(keyinput37), .Z(n15267) );
  XNOR2_X1 U16783 ( .A(P2_REG1_REG_1__SCAN_IN), .B(keyinput54), .ZN(n15266) );
  NAND2_X1 U16784 ( .A1(n15267), .A2(n15266), .ZN(n15268) );
  NOR4_X1 U16785 ( .A1(n15271), .A2(n15270), .A3(n15269), .A4(n15268), .ZN(
        n15272) );
  NAND4_X1 U16786 ( .A1(n15275), .A2(n15274), .A3(n15273), .A4(n15272), .ZN(
        n15276) );
  AOI211_X1 U16787 ( .C1(n15279), .C2(n15278), .A(n15277), .B(n15276), .ZN(
        n15284) );
  NAND2_X1 U16788 ( .A1(n15280), .A2(n15282), .ZN(n15281) );
  OAI21_X1 U16789 ( .B1(P2_REG0_REG_6__SCAN_IN), .B2(n15282), .A(n15281), .ZN(
        n15283) );
  XNOR2_X1 U16790 ( .A(n15284), .B(n15283), .ZN(P2_U3448) );
  XNOR2_X1 U16791 ( .A(n15286), .B(n15285), .ZN(SUB_1596_U59) );
  XNOR2_X1 U16792 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15287), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16793 ( .B1(n15288), .B2(n10179), .A(n15293), .ZN(SUB_1596_U53) );
  XOR2_X1 U16794 ( .A(n15290), .B(n15289), .Z(SUB_1596_U56) );
  XNOR2_X1 U16795 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15291), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U16796 ( .A(n15293), .B(n15292), .Z(SUB_1596_U5) );
  CLKBUF_X2 U7274 ( .A(n14489), .Z(n6459) );
  INV_X2 U7294 ( .A(n8312), .ZN(n9656) );
  CLKBUF_X1 U7601 ( .A(n8839), .Z(n9088) );
  CLKBUF_X1 U11285 ( .A(n9088), .Z(n9295) );
endmodule

