

module b21_C_SARLock_k_128_9 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4402, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235;

  NAND2_X1 U4896 ( .A1(n4938), .A2(n4939), .ZN(n8495) );
  INV_X1 U4897 ( .A(n5411), .ZN(n5456) );
  CLKBUF_X2 U4898 ( .A(n5399), .Z(n5540) );
  OR2_X1 U4899 ( .A1(n6041), .A2(n6398), .ZN(n5909) );
  AND2_X1 U4900 ( .A1(n6293), .A2(n8219), .ZN(n8224) );
  OR2_X1 U4901 ( .A1(n6649), .A2(n6760), .ZN(n7007) );
  CLKBUF_X2 U4902 ( .A(n8490), .Z(n4394) );
  NAND2_X1 U4903 ( .A1(n8224), .A2(n4394), .ZN(n8214) );
  OR2_X1 U4904 ( .A1(n8485), .A2(n8484), .ZN(n4801) );
  INV_X1 U4905 ( .A(n5846), .ZN(n5906) );
  NAND2_X1 U4906 ( .A1(n7774), .A2(n7773), .ZN(n8242) );
  INV_X1 U4908 ( .A(n5910), .ZN(n8025) );
  NAND2_X1 U4909 ( .A1(n8226), .A2(n4504), .ZN(n6305) );
  INV_X1 U4910 ( .A(n7994), .ZN(n7963) );
  INV_X1 U4911 ( .A(n7955), .ZN(n7992) );
  AOI21_X1 U4912 ( .B1(n8455), .B2(n6238), .A(n6237), .ZN(n8471) );
  INV_X1 U4913 ( .A(n5390), .ZN(n5562) );
  AND4_X1 U4914 ( .A1(n5446), .A2(n5445), .A3(n5444), .A4(n5443), .ZN(n7378)
         );
  OAI22_X2 U4915 ( .A1(n8495), .A2(n8498), .B1(n8505), .B2(n8356), .ZN(n8482)
         );
  NAND2_X2 U4916 ( .A1(n7139), .A2(n7138), .ZN(n7194) );
  NAND2_X2 U4917 ( .A1(n8011), .A2(n8148), .ZN(n8598) );
  INV_X1 U4918 ( .A(n5846), .ZN(n4390) );
  NAND4_X2 U4919 ( .A1(n5834), .A2(n5833), .A3(n5832), .A4(n5831), .ZN(n6649)
         );
  XNOR2_X2 U4920 ( .A(n6263), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8235) );
  INV_X2 U4921 ( .A(n7115), .ZN(n8631) );
  OAI21_X2 U4922 ( .B1(n8892), .B2(n8890), .A(n8888), .ZN(n8821) );
  XNOR2_X1 U4924 ( .A(n5111), .B(n5114), .ZN(n5765) );
  AOI21_X2 U4925 ( .B1(n4736), .B2(n4733), .A(n4732), .ZN(n4731) );
  AOI21_X2 U4926 ( .B1(n8814), .B2(n8815), .A(n4968), .ZN(n8892) );
  NAND2_X1 U4927 ( .A1(n4888), .A2(n4438), .ZN(n8285) );
  NOR2_X1 U4928 ( .A1(n5593), .A2(n5625), .ZN(n9131) );
  NAND2_X1 U4929 ( .A1(n4516), .A2(n4892), .ZN(n4888) );
  NAND2_X1 U4930 ( .A1(n5225), .A2(n5224), .ZN(n9419) );
  NAND2_X1 U4931 ( .A1(n7119), .A2(n7118), .ZN(n9729) );
  NAND2_X1 U4932 ( .A1(n7018), .A2(n7017), .ZN(n7040) );
  INV_X2 U4933 ( .A(n9785), .ZN(n4392) );
  INV_X2 U4934 ( .A(n9614), .ZN(n4393) );
  OAI211_X1 U4935 ( .C1(n6482), .C2(n6397), .A(n5909), .B(n5908), .ZN(n7115)
         );
  NAND2_X1 U4936 ( .A1(n6893), .A2(n6890), .ZN(n8073) );
  INV_X1 U4937 ( .A(n6891), .ZN(n6893) );
  XNOR2_X1 U4938 ( .A(n9772), .B(n9806), .ZN(n8086) );
  INV_X1 U4939 ( .A(n6892), .ZN(n6890) );
  CLKBUF_X2 U4940 ( .A(n5412), .Z(n5560) );
  INV_X2 U4941 ( .A(n8039), .ZN(n6759) );
  INV_X1 U4942 ( .A(n7208), .ZN(n7158) );
  BUF_X1 U4943 ( .A(n6424), .Z(n4402) );
  NAND2_X2 U4944 ( .A1(n5766), .A2(n5765), .ZN(n5408) );
  INV_X2 U4945 ( .A(n6384), .ZN(n4556) );
  NAND2_X1 U4946 ( .A1(n5420), .A2(n4584), .ZN(n5481) );
  INV_X4 U4947 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  INV_X1 U4948 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4974) );
  OAI21_X1 U4949 ( .B1(n8778), .B2(n8777), .A(n8944), .ZN(n8782) );
  NAND2_X1 U4950 ( .A1(n8840), .A2(n7976), .ZN(n8943) );
  AND2_X1 U4951 ( .A1(n8265), .A2(n8264), .ZN(n8646) );
  AND2_X1 U4952 ( .A1(n4908), .A2(n4905), .ZN(n8339) );
  NAND2_X1 U4953 ( .A1(n8451), .A2(n8458), .ZN(n8450) );
  AOI21_X1 U4954 ( .B1(n4512), .B2(n9774), .A(n4509), .ZN(n8655) );
  NAND2_X1 U4955 ( .A1(n4414), .A2(n9147), .ZN(n9146) );
  NAND2_X1 U4956 ( .A1(n8466), .A2(n8469), .ZN(n8465) );
  NAND2_X1 U4957 ( .A1(n4606), .A2(n4605), .ZN(n8868) );
  AND2_X1 U4958 ( .A1(n6202), .A2(n6203), .ZN(n4515) );
  INV_X1 U4959 ( .A(n9074), .ZN(n9354) );
  OR2_X1 U4960 ( .A1(n5593), .A2(n5698), .ZN(n5722) );
  NAND2_X1 U4961 ( .A1(n5133), .A2(n5132), .ZN(n9367) );
  NAND2_X1 U4962 ( .A1(n7788), .A2(n6092), .ZN(n7813) );
  NAND2_X1 U4963 ( .A1(n5536), .A2(n5535), .ZN(n9373) );
  XNOR2_X1 U4964 ( .A(n5131), .B(n5130), .ZN(n9475) );
  XNOR2_X1 U4965 ( .A(n5534), .B(n5533), .ZN(n8766) );
  NAND2_X1 U4966 ( .A1(n5534), .A2(n5533), .ZN(n5098) );
  OAI21_X1 U4967 ( .B1(n5163), .B2(n5162), .A(n5086), .ZN(n5522) );
  NAND2_X1 U4968 ( .A1(n5185), .A2(n5184), .ZN(n9405) );
  OAI21_X1 U4969 ( .B1(n7345), .B2(n4791), .A(n4789), .ZN(n4794) );
  XNOR2_X1 U4970 ( .A(n5193), .B(n5192), .ZN(n7359) );
  AOI21_X1 U4971 ( .B1(n9481), .B2(n9486), .A(n7635), .ZN(n7749) );
  NAND2_X1 U4972 ( .A1(n6121), .A2(n6120), .ZN(n8696) );
  OAI21_X1 U4973 ( .B1(n7281), .B2(n4929), .A(n4926), .ZN(n7634) );
  NAND2_X1 U4974 ( .A1(n5251), .A2(n5250), .ZN(n5047) );
  OR2_X1 U4975 ( .A1(n7451), .A2(n7446), .ZN(n8119) );
  INV_X1 U4976 ( .A(n8122), .ZN(n4395) );
  NAND2_X1 U4977 ( .A1(n5296), .A2(n5295), .ZN(n8837) );
  AND2_X1 U4978 ( .A1(n5996), .A2(n5995), .ZN(n7450) );
  NAND2_X2 U4979 ( .A1(n6805), .A2(n9750), .ZN(n9785) );
  AND2_X1 U4980 ( .A1(n4435), .A2(n6831), .ZN(n6876) );
  AND2_X1 U4981 ( .A1(n7197), .A2(n7196), .ZN(n7368) );
  NAND2_X2 U4982 ( .A1(n7287), .A2(n9605), .ZN(n9614) );
  NAND2_X1 U4983 ( .A1(n5362), .A2(n5361), .ZN(n7537) );
  INV_X1 U4984 ( .A(n7415), .ZN(n7387) );
  INV_X1 U4985 ( .A(n9660), .ZN(n7326) );
  AND3_X1 U4986 ( .A1(n5454), .A2(n5453), .A3(n5452), .ZN(n9660) );
  INV_X4 U4987 ( .A(n7848), .ZN(n7990) );
  AND2_X1 U4988 ( .A1(n5504), .A2(n5503), .ZN(n7415) );
  OR2_X1 U4989 ( .A1(n7068), .A2(n7265), .ZN(n5629) );
  CLKBUF_X3 U4990 ( .A(n6828), .Z(n7994) );
  NAND2_X1 U4991 ( .A1(n8073), .A2(n8080), .ZN(n7008) );
  AND4_X2 U4992 ( .A1(n5460), .A2(n5459), .A3(n5458), .A4(n5457), .ZN(n7297)
         );
  AND4_X1 U4993 ( .A1(n5496), .A2(n5495), .A3(n5494), .A4(n5493), .ZN(n7423)
         );
  CLKBUF_X1 U4994 ( .A(n6814), .Z(n7151) );
  AND2_X2 U4995 ( .A1(n6350), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  INV_X1 U4996 ( .A(n9649), .ZN(n7305) );
  INV_X1 U4997 ( .A(n7838), .ZN(n6973) );
  AND4_X1 U4998 ( .A1(n5917), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(n7117)
         );
  NAND4_X1 U4999 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n9772)
         );
  INV_X1 U5000 ( .A(n9214), .ZN(n6978) );
  INV_X1 U5001 ( .A(n5419), .ZN(n5502) );
  INV_X2 U5002 ( .A(n5480), .ZN(n5581) );
  OR3_X2 U5003 ( .A1(n7826), .A2(n7739), .A3(n7689), .ZN(n6785) );
  XNOR2_X1 U5004 ( .A(n5768), .B(n9938), .ZN(n7826) );
  INV_X1 U5005 ( .A(n8490), .ZN(n4504) );
  NAND2_X1 U5006 ( .A1(n5772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5768) );
  INV_X2 U5007 ( .A(n6213), .ZN(n4396) );
  INV_X1 U5008 ( .A(n8762), .ZN(n5824) );
  XNOR2_X1 U5009 ( .A(n5810), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U5010 ( .A1(n8756), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4802) );
  NAND2_X1 U5011 ( .A1(n4569), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U5012 ( .A1(n5110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5111) );
  OAI21_X1 U5013 ( .B1(n5767), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5770) );
  OR2_X1 U5014 ( .A1(n5819), .A2(n5795), .ZN(n5820) );
  XNOR2_X1 U5015 ( .A(n5794), .B(n5793), .ZN(n8765) );
  OR2_X1 U5016 ( .A1(n5811), .A2(n5795), .ZN(n5813) );
  AND2_X1 U5017 ( .A1(n5277), .A2(n5204), .ZN(n5267) );
  AND2_X1 U5018 ( .A1(n5806), .A2(n4646), .ZN(n5811) );
  AND2_X1 U5019 ( .A1(n5108), .A2(n4695), .ZN(n4694) );
  OR2_X2 U5020 ( .A1(n6384), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8769) );
  AND2_X1 U5021 ( .A1(n4972), .A2(n4969), .ZN(n5108) );
  AND2_X1 U5022 ( .A1(n5398), .A2(n4582), .ZN(n5420) );
  NAND4_X1 U5023 ( .A1(n4518), .A2(n5103), .A3(n4517), .A4(n5359), .ZN(n4583)
         );
  NAND2_X1 U5024 ( .A1(n7504), .A2(n4974), .ZN(n4977) );
  NAND2_X1 U5025 ( .A1(n7505), .A2(n4975), .ZN(n4976) );
  INV_X1 U5026 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5812) );
  INV_X1 U5027 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5755) );
  NOR2_X1 U5028 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4584) );
  INV_X1 U5029 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6266) );
  INV_X1 U5030 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5753) );
  INV_X1 U5031 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5104) );
  NOR2_X1 U5032 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4518) );
  INV_X1 U5033 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5103) );
  INV_X1 U5034 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4517) );
  INV_X4 U5035 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5036 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5359) );
  INV_X1 U5037 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4962) );
  INV_X1 U5038 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5958) );
  AND2_X1 U5039 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7505) );
  NOR2_X2 U5040 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7504) );
  AOI21_X2 U5041 ( .B1(n4601), .B2(n4870), .A(n4599), .ZN(n4598) );
  INV_X2 U5042 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4618) );
  XNOR2_X1 U5043 ( .A(n5813), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8490) );
  INV_X1 U5044 ( .A(n7521), .ZN(n4397) );
  AND2_X1 U5045 ( .A1(n6785), .A2(n6814), .ZN(n7521) );
  NAND2_X1 U5046 ( .A1(n5797), .A2(n5817), .ZN(n8767) );
  NOR2_X2 U5047 ( .A1(n8016), .A2(n8015), .ZN(n8485) );
  NOR3_X2 U5048 ( .A1(n8496), .A2(n8497), .A3(n8041), .ZN(n8016) );
  AND2_X1 U5049 ( .A1(n5887), .A2(n5786), .ZN(n5806) );
  AND3_X2 U5050 ( .A1(n5805), .A2(n5804), .A3(n5803), .ZN(n6892) );
  AND2_X1 U5051 ( .A1(n8224), .A2(n8038), .ZN(n4398) );
  NAND4_X2 U5052 ( .A1(n5786), .A2(n5792), .A3(n4813), .A4(n5887), .ZN(n5817)
         );
  OAI21_X2 U5053 ( .B1(n7040), .B2(n4964), .A(n4963), .ZN(n7114) );
  BUF_X4 U5054 ( .A(n4396), .Z(n4399) );
  AOI21_X2 U5055 ( .B1(n8469), .B2(n8468), .A(n8467), .ZN(n8470) );
  OR2_X2 U5056 ( .A1(n8614), .A2(n8618), .ZN(n8616) );
  NAND2_X1 U5057 ( .A1(n5823), .A2(n8762), .ZN(n6213) );
  AND2_X1 U5058 ( .A1(n6482), .A2(n6384), .ZN(n4400) );
  BUF_X4 U5059 ( .A(n6119), .Z(n6205) );
  NOR3_X2 U5060 ( .A1(n8514), .A2(n8179), .A3(n8512), .ZN(n8496) );
  NOR3_X4 U5061 ( .A1(n8550), .A2(n8530), .A3(n8529), .ZN(n8514) );
  AND2_X1 U5064 ( .A1(n4737), .A2(n5334), .ZN(n4736) );
  OR2_X1 U5065 ( .A1(n9258), .A2(n9257), .ZN(n4664) );
  NAND2_X1 U5066 ( .A1(n5408), .A2(n6384), .ZN(n5480) );
  AND2_X1 U5067 ( .A1(n9354), .A2(n9076), .ZN(n5718) );
  NOR2_X1 U5068 ( .A1(n4548), .A2(n4547), .ZN(n4546) );
  INV_X1 U5069 ( .A(n5661), .ZN(n4548) );
  INV_X1 U5070 ( .A(n9344), .ZN(n4547) );
  NOR2_X1 U5071 ( .A1(n8245), .A2(n8012), .ZN(n8014) );
  NAND2_X1 U5072 ( .A1(n4710), .A2(n9165), .ZN(n4709) );
  NAND2_X1 U5073 ( .A1(n4765), .A2(n4763), .ZN(n5577) );
  AOI21_X1 U5074 ( .B1(n4420), .B2(n4764), .A(n4494), .ZN(n4763) );
  NAND2_X1 U5075 ( .A1(n5098), .A2(n4766), .ZN(n4765) );
  NAND2_X1 U5076 ( .A1(n5009), .A2(n5008), .ZN(n5012) );
  OAI21_X1 U5077 ( .B1(n6380), .B2(P1_DATAO_REG_8__SCAN_IN), .A(n4498), .ZN(
        n5004) );
  NAND2_X1 U5078 ( .A1(n6380), .A2(n10091), .ZN(n4498) );
  NAND2_X1 U5079 ( .A1(n7812), .A2(n4894), .ZN(n4893) );
  OR2_X1 U5080 ( .A1(n8421), .A2(n8423), .ZN(n8215) );
  NAND2_X1 U5081 ( .A1(n6194), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U5082 ( .A1(n8739), .A2(n8551), .ZN(n4948) );
  NAND2_X1 U5083 ( .A1(n7607), .A2(n8131), .ZN(n7608) );
  INV_X1 U5084 ( .A(n4722), .ZN(n4721) );
  NAND2_X1 U5085 ( .A1(n7453), .A2(n7452), .ZN(n7455) );
  OAI21_X1 U5086 ( .B1(n7371), .B2(n4873), .A(n7526), .ZN(n4872) );
  AOI21_X1 U5087 ( .B1(n4870), .B2(n4871), .A(n4465), .ZN(n4596) );
  INV_X1 U5088 ( .A(n7846), .ZN(n4599) );
  NAND2_X1 U5089 ( .A1(n9419), .A2(n9288), .ZN(n4691) );
  NAND2_X1 U5090 ( .A1(n4457), .A2(n7701), .ZN(n7700) );
  NAND2_X1 U5091 ( .A1(n8837), .A2(n8906), .ZN(n5637) );
  OR2_X1 U5092 ( .A1(n7527), .A2(n7537), .ZN(n7512) );
  NAND2_X1 U5093 ( .A1(n4549), .A2(n5766), .ZN(n4557) );
  INV_X1 U5094 ( .A(n4553), .ZN(n4549) );
  XNOR2_X1 U5095 ( .A(n5577), .B(n5576), .ZN(n5575) );
  NAND2_X1 U5096 ( .A1(n5752), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5717) );
  AND2_X1 U5097 ( .A1(n5032), .A2(n5031), .ZN(n5275) );
  AND2_X1 U5098 ( .A1(n4434), .A2(n5105), .ZN(n4931) );
  INV_X1 U5099 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5105) );
  INV_X1 U5100 ( .A(n5305), .ZN(n5021) );
  NAND2_X1 U5101 ( .A1(n4729), .A2(n4680), .ZN(n4674) );
  NAND2_X1 U5102 ( .A1(n5004), .A2(n9950), .ZN(n5007) );
  INV_X1 U5103 ( .A(n6238), .ZN(n6295) );
  NOR2_X1 U5104 ( .A1(n8442), .A2(n8453), .ZN(n8441) );
  OR2_X1 U5105 ( .A1(n8664), .A2(n8501), .ZN(n8192) );
  AOI21_X1 U5106 ( .B1(n4941), .B2(n4943), .A(n4459), .ZN(n4939) );
  OR2_X1 U5107 ( .A1(n8537), .A2(n8551), .ZN(n8515) );
  AOI21_X1 U5108 ( .B1(n4944), .B2(n4946), .A(n4942), .ZN(n4941) );
  INV_X1 U5109 ( .A(n4944), .ZN(n4943) );
  NOR2_X1 U5110 ( .A1(n4956), .A2(n8244), .ZN(n4955) );
  INV_X1 U5111 ( .A(n8243), .ZN(n4956) );
  INV_X1 U5112 ( .A(n9770), .ZN(n9745) );
  OR2_X1 U5113 ( .A1(n6650), .A2(n6304), .ZN(n9743) );
  INV_X1 U5114 ( .A(n9774), .ZN(n9740) );
  AND2_X1 U5115 ( .A1(n4871), .A2(n4465), .ZN(n4601) );
  NAND2_X1 U5116 ( .A1(n8926), .A2(n8925), .ZN(n4585) );
  NAND2_X1 U5117 ( .A1(n5390), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U5119 ( .A1(n8005), .A2(n5124), .ZN(n5412) );
  AND2_X1 U5120 ( .A1(n8005), .A2(n9470), .ZN(n5411) );
  NAND2_X1 U5121 ( .A1(n5583), .A2(n5582), .ZN(n9074) );
  NAND2_X1 U5122 ( .A1(n9091), .A2(n4919), .ZN(n9258) );
  OR2_X1 U5123 ( .A1(n9411), .A2(n9289), .ZN(n4919) );
  NAND2_X1 U5124 ( .A1(n4685), .A2(n4691), .ZN(n4684) );
  INV_X1 U5125 ( .A(n4687), .ZN(n4685) );
  AOI21_X1 U5126 ( .B1(n4689), .B2(n9088), .A(n4688), .ZN(n4687) );
  INV_X1 U5127 ( .A(n9302), .ZN(n4688) );
  OR2_X1 U5128 ( .A1(n9084), .A2(n9348), .ZN(n9107) );
  AOI21_X1 U5129 ( .B1(n7754), .B2(n7753), .A(n7752), .ZN(n9109) );
  NOR2_X1 U5130 ( .A1(n9344), .A2(n4922), .ZN(n4921) );
  INV_X1 U5131 ( .A(n4924), .ZN(n4922) );
  OR2_X1 U5132 ( .A1(n9084), .A2(n10214), .ZN(n4924) );
  INV_X1 U5133 ( .A(n5408), .ZN(n5501) );
  INV_X1 U5134 ( .A(n9488), .ZN(n9308) );
  AOI21_X1 U5135 ( .B1(n4460), .B2(n4529), .A(n5777), .ZN(n4528) );
  INV_X1 U5136 ( .A(n4531), .ZN(n4529) );
  NAND2_X1 U5137 ( .A1(n4530), .A2(n4527), .ZN(n4526) );
  AOI21_X1 U5138 ( .B1(n5715), .B2(n6981), .A(n9607), .ZN(n4527) );
  NAND2_X1 U5139 ( .A1(n4561), .A2(n4559), .ZN(n5641) );
  NAND2_X1 U5140 ( .A1(n5635), .A2(n4562), .ZN(n4561) );
  OAI21_X1 U5141 ( .B1(n7314), .B2(n7311), .A(n4441), .ZN(n4560) );
  NAND2_X1 U5142 ( .A1(n4626), .A2(n4628), .ZN(n4621) );
  NAND2_X1 U5143 ( .A1(n4625), .A2(n8127), .ZN(n4622) );
  INV_X1 U5144 ( .A(n8135), .ZN(n4629) );
  INV_X1 U5145 ( .A(n4626), .ZN(n4623) );
  INV_X1 U5146 ( .A(n4625), .ZN(n4624) );
  NAND2_X1 U5147 ( .A1(n4541), .A2(n4539), .ZN(n5676) );
  AND2_X1 U5148 ( .A1(n5666), .A2(n4540), .ZN(n4539) );
  OAI21_X1 U5149 ( .B1(n4650), .B2(n4649), .A(n4648), .ZN(n8157) );
  AOI21_X1 U5150 ( .B1(n8146), .B2(n4442), .A(n4651), .ZN(n4650) );
  INV_X1 U5151 ( .A(n8618), .ZN(n4649) );
  NOR2_X1 U5152 ( .A1(n8155), .A2(n4811), .ZN(n4648) );
  AOI211_X1 U5153 ( .C1(n8177), .C2(n8214), .A(n4430), .B(n8512), .ZN(n4656)
         );
  INV_X1 U5154 ( .A(n8188), .ZN(n4655) );
  AOI21_X1 U5155 ( .B1(n4566), .B2(n4565), .A(n4563), .ZN(n5694) );
  OR2_X1 U5156 ( .A1(n5690), .A2(n4564), .ZN(n4563) );
  INV_X1 U5157 ( .A(n5688), .ZN(n4565) );
  OAI211_X1 U5158 ( .C1(n4568), .C2(n6701), .A(n4567), .B(n9123), .ZN(n4566)
         );
  NOR2_X1 U5159 ( .A1(n8505), .A2(n8664), .ZN(n4726) );
  AOI21_X1 U5160 ( .B1(n4778), .B2(n4776), .A(n4775), .ZN(n4774) );
  INV_X1 U5161 ( .A(n5275), .ZN(n4775) );
  INV_X1 U5162 ( .A(n4780), .ZN(n4776) );
  INV_X1 U5163 ( .A(n4778), .ZN(n4777) );
  INV_X1 U5164 ( .A(n4736), .ZN(n4734) );
  NOR2_X1 U5165 ( .A1(n6154), .A2(n8295), .ZN(n6159) );
  AND2_X1 U5166 ( .A1(n4643), .A2(n4633), .ZN(n4632) );
  NOR2_X1 U5167 ( .A1(n8205), .A2(n8197), .ZN(n4633) );
  OAI21_X1 U5168 ( .B1(n8218), .B2(n4638), .A(n8217), .ZN(n4637) );
  NOR2_X1 U5169 ( .A1(n4644), .A2(n4639), .ZN(n4638) );
  NOR3_X1 U5170 ( .A1(n8257), .A2(n8208), .A3(n8256), .ZN(n4639) );
  INV_X1 U5171 ( .A(n8218), .ZN(n4643) );
  NOR2_X1 U5172 ( .A1(n8218), .A2(n4640), .ZN(n4635) );
  NAND2_X1 U5173 ( .A1(n4642), .A2(n4641), .ZN(n4640) );
  INV_X1 U5174 ( .A(n8208), .ZN(n4642) );
  NOR2_X1 U5175 ( .A1(n8206), .A2(n8197), .ZN(n4636) );
  NOR2_X1 U5176 ( .A1(n8477), .A2(n4725), .ZN(n4724) );
  INV_X1 U5177 ( .A(n4726), .ZN(n4725) );
  OR2_X1 U5178 ( .A1(n8505), .A2(n8518), .ZN(n8184) );
  NAND2_X1 U5179 ( .A1(n6180), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U5180 ( .A1(n4808), .A2(n8013), .ZN(n4807) );
  NAND2_X1 U5181 ( .A1(n8014), .A2(n4809), .ZN(n4808) );
  INV_X1 U5182 ( .A(n6137), .ZN(n6136) );
  OR2_X1 U5183 ( .A1(n7798), .A2(n8359), .ZN(n8147) );
  NAND2_X1 U5184 ( .A1(n4395), .A2(n8119), .ZN(n4791) );
  NAND2_X1 U5185 ( .A1(n7228), .A2(n4449), .ZN(n7349) );
  INV_X1 U5186 ( .A(n8052), .ZN(n7229) );
  OR2_X1 U5187 ( .A1(n7346), .A2(n7226), .ZN(n4722) );
  NOR2_X1 U5188 ( .A1(n8544), .A2(n8537), .ZN(n8536) );
  NAND2_X1 U5189 ( .A1(n4405), .A2(n4957), .ZN(n4954) );
  AOI21_X1 U5190 ( .B1(n4405), .B2(n4953), .A(n4454), .ZN(n4952) );
  INV_X1 U5191 ( .A(n7524), .ZN(n4873) );
  NOR2_X1 U5192 ( .A1(n4431), .A2(n4613), .ZN(n4611) );
  INV_X1 U5193 ( .A(n7950), .ZN(n4879) );
  AOI21_X1 U5194 ( .B1(n4611), .B2(n4609), .A(n4608), .ZN(n4607) );
  INV_X1 U5195 ( .A(n4876), .ZN(n4608) );
  INV_X1 U5196 ( .A(n8822), .ZN(n4609) );
  INV_X1 U5197 ( .A(n4601), .ZN(n4600) );
  AND2_X1 U5198 ( .A1(n6783), .A2(n7521), .ZN(n6828) );
  AND2_X1 U5199 ( .A1(n4863), .A2(n4423), .ZN(n4862) );
  NOR2_X1 U5200 ( .A1(n4535), .A2(n4534), .ZN(n4533) );
  INV_X1 U5201 ( .A(n9129), .ZN(n4534) );
  NOR2_X1 U5202 ( .A1(n5703), .A2(n4536), .ZN(n4535) );
  NAND2_X1 U5203 ( .A1(n5705), .A2(n5704), .ZN(n4536) );
  INV_X1 U5204 ( .A(n5718), .ZN(n5750) );
  NOR2_X1 U5205 ( .A1(n5749), .A2(n9354), .ZN(n5707) );
  NOR2_X1 U5206 ( .A1(n4709), .A2(n5551), .ZN(n4708) );
  AND2_X1 U5207 ( .A1(n5704), .A2(n5720), .ZN(n4830) );
  NOR2_X1 U5208 ( .A1(n9389), .A2(n9095), .ZN(n9124) );
  INV_X1 U5209 ( .A(n9227), .ZN(n4839) );
  OR2_X1 U5210 ( .A1(n9411), .A2(n9254), .ZN(n9117) );
  NAND2_X1 U5211 ( .A1(n4819), .A2(n4818), .ZN(n4817) );
  INV_X1 U5212 ( .A(n4825), .ZN(n4818) );
  NOR2_X1 U5213 ( .A1(n9112), .A2(n4826), .ZN(n4825) );
  INV_X1 U5214 ( .A(n9107), .ZN(n4826) );
  OR2_X1 U5215 ( .A1(n7315), .A2(n7137), .ZN(n5631) );
  AND2_X1 U5216 ( .A1(n5205), .A2(n10005), .ZN(n4883) );
  NAND2_X1 U5217 ( .A1(n4827), .A2(n7208), .ZN(n4828) );
  INV_X1 U5218 ( .A(n4709), .ZN(n4707) );
  OR2_X1 U5219 ( .A1(n5097), .A2(n4769), .ZN(n4768) );
  AOI21_X1 U5220 ( .B1(n4759), .B2(n4760), .A(n4486), .ZN(n4758) );
  NAND2_X1 U5221 ( .A1(n5589), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5590) );
  AOI21_X1 U5222 ( .B1(n4750), .B2(n4752), .A(n4485), .ZN(n4748) );
  NOR2_X1 U5223 ( .A1(n5052), .A2(n4754), .ZN(n4753) );
  INV_X1 U5224 ( .A(n5046), .ZN(n4754) );
  NOR2_X1 U5225 ( .A1(n5291), .A2(n4781), .ZN(n4780) );
  INV_X1 U5226 ( .A(n5020), .ZN(n4781) );
  AOI21_X1 U5227 ( .B1(n4780), .B2(n5021), .A(n4779), .ZN(n4778) );
  INV_X1 U5228 ( .A(n5026), .ZN(n4779) );
  INV_X1 U5229 ( .A(n5007), .ZN(n4733) );
  INV_X1 U5230 ( .A(n5012), .ZN(n4732) );
  AND2_X1 U5231 ( .A1(n5017), .A2(n5016), .ZN(n5318) );
  NAND2_X1 U5232 ( .A1(n5007), .A2(n5006), .ZN(n5357) );
  XNOR2_X1 U5233 ( .A(n5001), .B(SI_7_), .ZN(n5497) );
  INV_X1 U5234 ( .A(n4996), .ZN(n4662) );
  OR2_X1 U5235 ( .A1(n6232), .A2(n6231), .ZN(n6244) );
  NOR2_X1 U5236 ( .A1(n7434), .A2(n4917), .ZN(n4916) );
  INV_X1 U5237 ( .A(n6028), .ZN(n4917) );
  NOR2_X1 U5238 ( .A1(n7095), .A2(n4912), .ZN(n4911) );
  INV_X1 U5239 ( .A(n5957), .ZN(n4912) );
  INV_X1 U5240 ( .A(n8287), .ZN(n4887) );
  NAND2_X1 U5241 ( .A1(n6032), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6048) );
  INV_X1 U5242 ( .A(n6033), .ZN(n6032) );
  NAND2_X1 U5243 ( .A1(n4915), .A2(n4914), .ZN(n7591) );
  AND2_X1 U5244 ( .A1(n7593), .A2(n4433), .ZN(n4914) );
  INV_X1 U5245 ( .A(n5857), .ZN(n5910) );
  OR3_X1 U5246 ( .A1(n7687), .A2(n7821), .A3(n7741), .ZN(n6460) );
  AND4_X1 U5247 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n7670)
         );
  AND4_X1 U5248 ( .A1(n5953), .A2(n5952), .A3(n5951), .A4(n5950), .ZN(n7225)
         );
  AND2_X1 U5249 ( .A1(n8255), .A2(n8441), .ZN(n8428) );
  NAND2_X1 U5250 ( .A1(n8450), .A2(n4950), .ZN(n8434) );
  OR2_X1 U5251 ( .A1(n8652), .A2(n8353), .ZN(n4950) );
  NAND2_X1 U5252 ( .A1(n8434), .A2(n8436), .ZN(n8433) );
  NAND2_X1 U5253 ( .A1(n4461), .A2(n8018), .ZN(n4796) );
  NAND2_X1 U5254 ( .A1(n8460), .A2(n9771), .ZN(n4511) );
  NAND2_X1 U5255 ( .A1(n8018), .A2(n8198), .ZN(n8458) );
  OR2_X1 U5256 ( .A1(n8664), .A2(n8355), .ZN(n8248) );
  AND2_X1 U5257 ( .A1(n6225), .A2(n6224), .ZN(n8487) );
  NAND2_X1 U5258 ( .A1(n4463), .A2(n4948), .ZN(n4944) );
  OR2_X1 U5259 ( .A1(n8569), .A2(n8559), .ZN(n8544) );
  NAND2_X1 U5260 ( .A1(n6122), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6137) );
  INV_X1 U5261 ( .A(n6123), .ZN(n6122) );
  XNOR2_X1 U5262 ( .A(n8706), .B(n8358), .ZN(n8618) );
  AND2_X1 U5263 ( .A1(n8135), .A2(n7560), .ZN(n4959) );
  OR2_X1 U5264 ( .A1(n7467), .A2(n7559), .ZN(n7565) );
  AND4_X1 U5265 ( .A1(n6022), .A2(n6021), .A3(n6020), .A4(n6019), .ZN(n7461)
         );
  NOR2_X1 U5266 ( .A1(n8048), .A2(n4793), .ZN(n4792) );
  AND4_X1 U5267 ( .A1(n5988), .A2(n5987), .A3(n5986), .A4(n5985), .ZN(n7446)
         );
  AND2_X1 U5268 ( .A1(n8116), .A2(n8112), .ZN(n8052) );
  AND2_X1 U5269 ( .A1(n8100), .A2(n8101), .ZN(n4806) );
  NOR2_X1 U5270 ( .A1(n8370), .A2(n7041), .ZN(n4964) );
  OR2_X1 U5271 ( .A1(n8045), .A2(n9821), .ZN(n4963) );
  NAND2_X1 U5272 ( .A1(n7023), .A2(n8046), .ZN(n7110) );
  NAND2_X1 U5273 ( .A1(n6891), .A2(n6892), .ZN(n8080) );
  INV_X1 U5274 ( .A(n6904), .ZN(n9769) );
  NAND2_X1 U5275 ( .A1(n8081), .A2(n8079), .ZN(n6904) );
  NAND2_X1 U5276 ( .A1(n8024), .A2(n8023), .ZN(n8429) );
  NAND2_X1 U5277 ( .A1(n8020), .A2(n8019), .ZN(n8643) );
  NAND2_X1 U5278 ( .A1(n6031), .A2(n6030), .ZN(n7602) );
  AND2_X1 U5279 ( .A1(n4965), .A2(n4814), .ZN(n4813) );
  NOR2_X1 U5280 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4814) );
  INV_X4 U5281 ( .A(n4556), .ZN(n6380) );
  NAND2_X1 U5282 ( .A1(n8943), .A2(n7987), .ZN(n8774) );
  OR2_X1 U5283 ( .A1(n5312), .A2(n5298), .ZN(n5300) );
  NAND2_X1 U5284 ( .A1(n8865), .A2(n7965), .ZN(n8841) );
  AND2_X1 U5285 ( .A1(n7915), .A2(n7916), .ZN(n8850) );
  NOR2_X1 U5286 ( .A1(n4596), .A2(n4598), .ZN(n4589) );
  NOR2_X1 U5287 ( .A1(n4590), .A2(n4588), .ZN(n4587) );
  AND2_X1 U5288 ( .A1(n4596), .A2(n4597), .ZN(n4588) );
  NOR2_X1 U5289 ( .A1(n4604), .A2(n4600), .ZN(n4593) );
  NAND2_X1 U5290 ( .A1(n7373), .A2(n4871), .ZN(n4586) );
  INV_X1 U5291 ( .A(n4598), .ZN(n4595) );
  NAND2_X1 U5292 ( .A1(n4585), .A2(n4448), .ZN(n8829) );
  AOI22_X1 U5293 ( .A1(n4866), .A2(n8850), .B1(n4865), .B2(n4427), .ZN(n4863)
         );
  INV_X1 U5294 ( .A(n8858), .ZN(n4865) );
  AND4_X1 U5295 ( .A1(n5356), .A2(n5355), .A3(n5354), .A4(n5353), .ZN(n7527)
         );
  NAND2_X1 U5296 ( .A1(n6865), .A2(n4497), .ZN(n6569) );
  OR2_X1 U5297 ( .A1(n6861), .A2(n6335), .ZN(n4497) );
  NAND2_X1 U5298 ( .A1(n9571), .A2(n4570), .ZN(n6630) );
  NAND2_X1 U5299 ( .A1(n9568), .A2(n5428), .ZN(n4570) );
  NAND2_X1 U5300 ( .A1(n8997), .A2(n8998), .ZN(n8996) );
  OR2_X1 U5301 ( .A1(n6921), .A2(n6920), .ZN(n4578) );
  AND2_X1 U5302 ( .A1(n4578), .A2(n4577), .ZN(n7087) );
  NAND2_X1 U5303 ( .A1(n6642), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4577) );
  OR2_X1 U5304 ( .A1(n7087), .A2(n7086), .ZN(n4576) );
  OR2_X1 U5305 ( .A1(n9015), .A2(n9014), .ZN(n4573) );
  AND2_X1 U5306 ( .A1(n4573), .A2(n4572), .ZN(n9032) );
  NAND2_X1 U5307 ( .A1(n9034), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4572) );
  AOI21_X1 U5308 ( .B1(n9034), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9033), .ZN(
        n9036) );
  NAND2_X1 U5309 ( .A1(n9199), .A2(n5720), .ZN(n4832) );
  NAND2_X1 U5310 ( .A1(n4933), .A2(n4447), .ZN(n4672) );
  INV_X1 U5311 ( .A(n9100), .ZN(n4673) );
  OR2_X1 U5312 ( .A1(n9382), .A2(n9210), .ZN(n9180) );
  NAND2_X1 U5313 ( .A1(n9191), .A2(n9200), .ZN(n4933) );
  NOR2_X1 U5314 ( .A1(n9220), .A2(n9389), .ZN(n9211) );
  NAND2_X1 U5315 ( .A1(n9180), .A2(n5626), .ZN(n9200) );
  AOI21_X1 U5316 ( .B1(n9219), .B2(n9094), .A(n9093), .ZN(n9206) );
  NAND2_X1 U5317 ( .A1(n9257), .A2(n5248), .ZN(n4843) );
  INV_X1 U5318 ( .A(n4842), .ZN(n4841) );
  OAI21_X1 U5319 ( .B1(n9121), .B2(n5672), .A(n9120), .ZN(n4842) );
  NAND2_X1 U5320 ( .A1(n4664), .A2(n4451), .ZN(n4918) );
  OR2_X1 U5321 ( .A1(n9251), .A2(n9252), .ZN(n4844) );
  OR2_X1 U5322 ( .A1(n5210), .A2(n9992), .ZN(n5197) );
  AND2_X1 U5323 ( .A1(n9090), .A2(n9089), .ZN(n9263) );
  AND2_X1 U5324 ( .A1(n4684), .A2(n4464), .ZN(n4682) );
  AND2_X1 U5325 ( .A1(n5677), .A2(n9116), .ZN(n9287) );
  NOR2_X1 U5326 ( .A1(n4690), .A2(n4453), .ZN(n4689) );
  NOR2_X1 U5327 ( .A1(n9088), .A2(n4426), .ZN(n4690) );
  INV_X1 U5328 ( .A(n4823), .ZN(n4822) );
  OAI21_X1 U5329 ( .B1(n9112), .B2(n4824), .A(n9111), .ZN(n4823) );
  NAND2_X1 U5330 ( .A1(n9108), .A2(n9107), .ZN(n4824) );
  NAND2_X1 U5331 ( .A1(n9109), .A2(n4825), .ZN(n4821) );
  NAND2_X1 U5332 ( .A1(n7751), .A2(n4440), .ZN(n4923) );
  INV_X1 U5333 ( .A(n7750), .ZN(n4925) );
  INV_X1 U5334 ( .A(n10214), .ZN(n9348) );
  OAI21_X1 U5335 ( .B1(n7692), .B2(n4458), .A(n4845), .ZN(n7754) );
  OR2_X1 U5336 ( .A1(n4406), .A2(n4846), .ZN(n4845) );
  INV_X1 U5337 ( .A(n7694), .ZN(n4846) );
  OR2_X1 U5338 ( .A1(n7704), .A2(n7703), .ZN(n7746) );
  AND2_X1 U5339 ( .A1(n7714), .A2(n4436), .ZN(n7703) );
  AND2_X1 U5340 ( .A1(n5599), .A2(n7694), .ZN(n7719) );
  NOR2_X1 U5341 ( .A1(n7647), .A2(n9501), .ZN(n9502) );
  OAI21_X1 U5342 ( .B1(n7634), .B2(n7633), .A(n7632), .ZN(n9481) );
  AND2_X1 U5343 ( .A1(n7278), .A2(n7277), .ZN(n7312) );
  AND4_X1 U5344 ( .A1(n5477), .A2(n5476), .A3(n5475), .A4(n5474), .ZN(n7068)
         );
  AND2_X1 U5345 ( .A1(n5631), .A2(n5630), .ZN(n7066) );
  NAND2_X1 U5346 ( .A1(n7257), .A2(n7267), .ZN(n7259) );
  NAND2_X1 U5347 ( .A1(n5763), .A2(n4867), .ZN(n6980) );
  INV_X1 U5348 ( .A(n9607), .ZN(n4867) );
  OR2_X1 U5349 ( .A1(n5412), .A2(n6335), .ZN(n5413) );
  OR2_X1 U5350 ( .A1(n6981), .A2(n4391), .ZN(n9491) );
  INV_X1 U5351 ( .A(n9492), .ZN(n9305) );
  NAND2_X1 U5352 ( .A1(n5524), .A2(n5523), .ZN(n9377) );
  NAND2_X1 U5353 ( .A1(n7819), .A2(n5581), .ZN(n5524) );
  AND3_X1 U5354 ( .A1(n5487), .A2(n5486), .A3(n5485), .ZN(n9654) );
  AND3_X1 U5355 ( .A1(n5468), .A2(n5467), .A3(n5466), .ZN(n7838) );
  NAND2_X1 U5356 ( .A1(n4551), .A2(n4550), .ZN(n9645) );
  NAND2_X1 U5357 ( .A1(n4557), .A2(n4552), .ZN(n4551) );
  NOR2_X1 U5358 ( .A1(n4555), .A2(n4415), .ZN(n4552) );
  NAND2_X1 U5359 ( .A1(n5619), .A2(n5714), .ZN(n7206) );
  INV_X1 U5360 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4936) );
  INV_X1 U5361 ( .A(n4937), .ZN(n4934) );
  NAND2_X1 U5362 ( .A1(n5092), .A2(n5091), .ZN(n5534) );
  OAI21_X1 U5363 ( .B1(n5172), .B2(n5171), .A(n5073), .ZN(n5152) );
  NAND2_X1 U5364 ( .A1(n4762), .A2(n5066), .ZN(n5182) );
  NAND2_X1 U5365 ( .A1(n5193), .A2(n5192), .ZN(n4762) );
  INV_X1 U5366 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4930) );
  XNOR2_X1 U5367 ( .A(n5292), .B(n5291), .ZN(n6641) );
  NAND2_X1 U5368 ( .A1(n4681), .A2(n5020), .ZN(n5292) );
  NOR2_X1 U5369 ( .A1(n5021), .A2(n4679), .ZN(n4675) );
  NAND2_X1 U5370 ( .A1(n4514), .A2(n4513), .ZN(n8279) );
  NAND2_X1 U5371 ( .A1(n6178), .A2(n6179), .ZN(n4513) );
  OR2_X1 U5372 ( .A1(n6178), .A2(n4462), .ZN(n4514) );
  NAND2_X1 U5373 ( .A1(n6242), .A2(n6241), .ZN(n8442) );
  NAND2_X1 U5374 ( .A1(n9475), .A2(n6204), .ZN(n6242) );
  NOR2_X1 U5375 ( .A1(n8327), .A2(n8326), .ZN(n8325) );
  XNOR2_X1 U5376 ( .A(n6178), .B(n6171), .ZN(n8327) );
  NAND2_X1 U5377 ( .A1(n6109), .A2(n6108), .ZN(n8604) );
  INV_X1 U5378 ( .A(n8332), .ZN(n8344) );
  AND2_X1 U5379 ( .A1(n6462), .A2(n6304), .ZN(n9770) );
  INV_X1 U5380 ( .A(n8249), .ZN(n8460) );
  NAND2_X1 U5381 ( .A1(n4507), .A2(n4506), .ZN(n7574) );
  NAND2_X1 U5382 ( .A1(n7573), .A2(n7588), .ZN(n4506) );
  INV_X1 U5383 ( .A(n8404), .ZN(n4507) );
  NAND2_X1 U5384 ( .A1(n4502), .A2(n4501), .ZN(n4500) );
  NOR2_X1 U5385 ( .A1(n9709), .A2(n4504), .ZN(n4501) );
  NAND2_X1 U5386 ( .A1(n8414), .A2(n9711), .ZN(n4502) );
  NAND2_X1 U5387 ( .A1(n8415), .A2(n4504), .ZN(n4503) );
  NAND2_X1 U5388 ( .A1(n4801), .A2(n8192), .ZN(n8468) );
  NAND2_X1 U5389 ( .A1(n9475), .A2(n5581), .ZN(n5133) );
  NAND2_X1 U5390 ( .A1(n5255), .A2(n5254), .ZN(n9431) );
  NAND2_X1 U5391 ( .A1(n5236), .A2(n5235), .ZN(n9426) );
  INV_X1 U5392 ( .A(n9389), .ZN(n9096) );
  INV_X1 U5393 ( .A(n8971), .ZN(n9238) );
  OR2_X1 U5394 ( .A1(n5412), .A2(n6591), .ZN(n5391) );
  NAND2_X1 U5395 ( .A1(n5377), .A2(n5376), .ZN(n9084) );
  NAND2_X1 U5396 ( .A1(n4744), .A2(n4743), .ZN(n5719) );
  OR2_X1 U5397 ( .A1(n5711), .A2(n5712), .ZN(n4743) );
  AND2_X1 U5398 ( .A1(n4524), .A2(n5776), .ZN(n4523) );
  NAND2_X1 U5399 ( .A1(n4528), .A2(n4531), .ZN(n4525) );
  OR2_X1 U5400 ( .A1(n5399), .A2(n7209), .ZN(n5402) );
  OR2_X1 U5401 ( .A1(n5412), .A2(n8988), .ZN(n5401) );
  INV_X1 U5402 ( .A(n8129), .ZN(n4628) );
  AOI21_X1 U5403 ( .B1(n4417), .B2(n8130), .A(n8197), .ZN(n4625) );
  AND2_X1 U5404 ( .A1(n4630), .A2(n4627), .ZN(n4626) );
  NAND2_X1 U5405 ( .A1(n8122), .A2(n8129), .ZN(n4627) );
  NOR2_X1 U5406 ( .A1(n8127), .A2(n8214), .ZN(n4630) );
  AOI21_X1 U5407 ( .B1(n5641), .B2(n7512), .A(n4558), .ZN(n5639) );
  OR2_X1 U5408 ( .A1(n5636), .A2(n5643), .ZN(n4558) );
  AOI21_X1 U5409 ( .B1(n4546), .B2(n4544), .A(n4543), .ZN(n4542) );
  NAND2_X1 U5410 ( .A1(n5658), .A2(n7755), .ZN(n4544) );
  NAND2_X1 U5411 ( .A1(n9315), .A2(n5662), .ZN(n4543) );
  NAND2_X1 U5412 ( .A1(n4542), .A2(n4545), .ZN(n4540) );
  INV_X1 U5413 ( .A(n4546), .ZN(n4545) );
  NAND2_X1 U5414 ( .A1(n4409), .A2(n4452), .ZN(n4619) );
  NOR2_X1 U5415 ( .A1(n8147), .A2(n8197), .ZN(n4651) );
  INV_X1 U5416 ( .A(n8157), .ZN(n8167) );
  OR2_X1 U5417 ( .A1(n5685), .A2(n4562), .ZN(n4567) );
  AOI21_X1 U5418 ( .B1(n5675), .B2(n9120), .A(n5674), .ZN(n4568) );
  AND2_X1 U5419 ( .A1(n9125), .A2(n6701), .ZN(n4564) );
  INV_X1 U5420 ( .A(n7154), .ZN(n5602) );
  AND2_X1 U5421 ( .A1(n4420), .A2(n4767), .ZN(n4766) );
  INV_X1 U5422 ( .A(n5569), .ZN(n4767) );
  NOR2_X1 U5423 ( .A1(n5569), .A2(n5130), .ZN(n4764) );
  NAND2_X1 U5424 ( .A1(n8207), .A2(n8197), .ZN(n4645) );
  OR2_X1 U5425 ( .A1(n4656), .A2(n8188), .ZN(n4653) );
  OR2_X1 U5426 ( .A1(n8643), .A2(n8438), .ZN(n8204) );
  INV_X1 U5427 ( .A(n4810), .ZN(n4809) );
  NOR2_X1 U5428 ( .A1(n4955), .A2(n4958), .ZN(n4953) );
  OAI21_X1 U5429 ( .B1(n4538), .B2(n6701), .A(n4537), .ZN(n5703) );
  NAND2_X1 U5430 ( .A1(n5695), .A2(n6701), .ZN(n4537) );
  INV_X1 U5431 ( .A(n5696), .ZN(n4538) );
  OR2_X1 U5432 ( .A1(n9367), .A2(n9168), .ZN(n5705) );
  NOR2_X1 U5433 ( .A1(n4761), .A2(n4757), .ZN(n4756) );
  INV_X1 U5434 ( .A(n5061), .ZN(n4757) );
  INV_X1 U5435 ( .A(n5192), .ZN(n4759) );
  INV_X1 U5436 ( .A(n4751), .ZN(n4750) );
  OAI21_X1 U5437 ( .B1(n4753), .B2(n4752), .A(n5053), .ZN(n4751) );
  INV_X1 U5438 ( .A(n5051), .ZN(n4752) );
  INV_X1 U5439 ( .A(n5497), .ZN(n5000) );
  INV_X1 U5440 ( .A(n6228), .ZN(n4902) );
  OR2_X1 U5441 ( .A1(n8303), .A2(n8302), .ZN(n4909) );
  NOR2_X1 U5442 ( .A1(n8469), .A2(n4798), .ZN(n4797) );
  NAND2_X1 U5443 ( .A1(n8484), .A2(n8192), .ZN(n4798) );
  OR2_X1 U5444 ( .A1(n8442), .A2(n8249), .ZN(n8256) );
  NOR2_X1 U5445 ( .A1(n8469), .A2(n4800), .ZN(n4799) );
  INV_X1 U5446 ( .A(n8192), .ZN(n4800) );
  OR2_X1 U5447 ( .A1(n8477), .A2(n8487), .ZN(n8194) );
  NOR2_X1 U5448 ( .A1(n8589), .A2(n4811), .ZN(n4810) );
  NOR2_X1 U5449 ( .A1(n7671), .A2(n8141), .ZN(n4717) );
  NAND2_X1 U5450 ( .A1(n8598), .A2(n8599), .ZN(n4812) );
  NAND2_X1 U5451 ( .A1(n9779), .A2(n9778), .ZN(n6899) );
  INV_X1 U5452 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4965) );
  AND2_X1 U5453 ( .A1(n4425), .A2(n5787), .ZN(n4646) );
  NAND2_X1 U5454 ( .A1(n4877), .A2(n7950), .ZN(n4876) );
  INV_X1 U5455 ( .A(n8913), .ZN(n4877) );
  NAND2_X1 U5456 ( .A1(n4598), .A2(n4600), .ZN(n4591) );
  AND2_X1 U5457 ( .A1(n4576), .A2(n4575), .ZN(n6362) );
  NAND2_X1 U5458 ( .A1(n7083), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4575) );
  AND2_X1 U5459 ( .A1(n5551), .A2(n5550), .ZN(n5625) );
  OR2_X1 U5460 ( .A1(n9244), .A2(n9228), .ZN(n9120) );
  NOR2_X1 U5461 ( .A1(n9405), .A2(n9411), .ZN(n4701) );
  NOR2_X1 U5462 ( .A1(n8837), .A2(n8930), .ZN(n4699) );
  NOR2_X1 U5463 ( .A1(n7387), .A2(n7326), .ZN(n4705) );
  OR2_X1 U5464 ( .A1(n7423), .A2(n7387), .ZN(n5735) );
  NAND2_X1 U5465 ( .A1(n5762), .A2(n7362), .ZN(n6814) );
  NAND2_X1 U5466 ( .A1(n4391), .A2(n4554), .ZN(n4553) );
  INV_X1 U5467 ( .A(n6590), .ZN(n4554) );
  NOR2_X1 U5468 ( .A1(n6385), .A2(n4556), .ZN(n4555) );
  INV_X1 U5469 ( .A(SI_30_), .ZN(n4746) );
  AND2_X1 U5470 ( .A1(n9923), .A2(n5114), .ZN(n4937) );
  AND2_X1 U5471 ( .A1(n4883), .A2(n5587), .ZN(n4882) );
  NAND2_X1 U5472 ( .A1(n5062), .A2(n5061), .ZN(n5193) );
  AOI21_X1 U5473 ( .B1(n4774), .B2(n4777), .A(n4772), .ZN(n4771) );
  INV_X1 U5474 ( .A(n5032), .ZN(n4772) );
  INV_X1 U5475 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n4932) );
  XNOR2_X1 U5476 ( .A(n5018), .B(SI_11_), .ZN(n5305) );
  OR2_X1 U5477 ( .A1(n5358), .A2(n4734), .ZN(n4728) );
  INV_X1 U5478 ( .A(n5318), .ZN(n4730) );
  OR2_X1 U5479 ( .A1(n4671), .A2(n4421), .ZN(n4669) );
  INV_X1 U5480 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4582) );
  INV_X1 U5481 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4975) );
  AOI21_X1 U5482 ( .B1(n4892), .B2(n4890), .A(n4456), .ZN(n4889) );
  INV_X1 U5483 ( .A(n4894), .ZN(n4890) );
  INV_X1 U5484 ( .A(n7813), .ZN(n4516) );
  INV_X1 U5485 ( .A(n4910), .ZN(n8271) );
  OAI21_X1 U5486 ( .B1(n8305), .B2(n4906), .A(n4901), .ZN(n4910) );
  AOI21_X1 U5487 ( .B1(n4903), .B2(n4905), .A(n4902), .ZN(n4901) );
  INV_X1 U5488 ( .A(n4909), .ZN(n4903) );
  OR2_X1 U5489 ( .A1(n6073), .A2(n4900), .ZN(n4897) );
  INV_X1 U5490 ( .A(n7620), .ZN(n4900) );
  NAND2_X1 U5491 ( .A1(n4899), .A2(n4443), .ZN(n4898) );
  INV_X1 U5492 ( .A(n7623), .ZN(n4899) );
  OAI21_X1 U5493 ( .B1(n6730), .B2(n6731), .A(n4886), .ZN(n4885) );
  NAND2_X1 U5494 ( .A1(n4898), .A2(n4895), .ZN(n7788) );
  NOR2_X1 U5495 ( .A1(n7791), .A2(n4896), .ZN(n4895) );
  INV_X1 U5496 ( .A(n4897), .ZN(n4896) );
  INV_X1 U5497 ( .A(n6017), .ZN(n6014) );
  OR2_X1 U5498 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  OR2_X1 U5499 ( .A1(n8318), .A2(n6159), .ZN(n6161) );
  OR2_X1 U5500 ( .A1(n6105), .A2(n6104), .ZN(n4894) );
  AND2_X1 U5501 ( .A1(n8303), .A2(n8302), .ZN(n4907) );
  OR2_X1 U5502 ( .A1(n6048), .A2(n6047), .ZN(n6067) );
  NAND2_X1 U5503 ( .A1(n6066), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6081) );
  INV_X1 U5504 ( .A(n6067), .ZN(n6066) );
  OAI21_X1 U5505 ( .B1(n8209), .B2(n4634), .A(n4631), .ZN(n8227) );
  AOI21_X1 U5506 ( .B1(n4643), .B2(n4636), .A(n4635), .ZN(n4634) );
  NOR2_X1 U5507 ( .A1(n4632), .A2(n4637), .ZN(n4631) );
  AND4_X1 U5508 ( .A1(n6038), .A2(n6037), .A3(n6036), .A4(n6035), .ZN(n7596)
         );
  AOI21_X1 U5509 ( .B1(n8375), .B2(n8374), .A(n8373), .ZN(n6533) );
  OR2_X1 U5510 ( .A1(n5923), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5942) );
  OR3_X1 U5511 ( .A1(n6009), .A2(P2_IR_REG_10__SCAN_IN), .A3(n6008), .ZN(n6029) );
  NOR2_X1 U5512 ( .A1(n7048), .A2(n7047), .ZN(n7173) );
  NAND2_X1 U5513 ( .A1(n8519), .A2(n4724), .ZN(n8472) );
  NAND2_X1 U5514 ( .A1(n8519), .A2(n4413), .ZN(n8453) );
  NAND2_X1 U5515 ( .A1(n8465), .A2(n4508), .ZN(n8451) );
  OR2_X1 U5516 ( .A1(n8477), .A2(n8461), .ZN(n4508) );
  NAND2_X1 U5517 ( .A1(n8194), .A2(n8017), .ZN(n8469) );
  NAND2_X1 U5518 ( .A1(n8192), .A2(n8189), .ZN(n8484) );
  AND2_X1 U5519 ( .A1(n8536), .A2(n8525), .ZN(n8519) );
  NAND2_X1 U5520 ( .A1(n8519), .A2(n8734), .ZN(n8502) );
  INV_X1 U5521 ( .A(n8041), .ZN(n8498) );
  AND2_X1 U5522 ( .A1(n8603), .A2(n8250), .ZN(n8584) );
  NAND2_X1 U5523 ( .A1(n8584), .A2(n8570), .ZN(n8569) );
  NAND2_X1 U5524 ( .A1(n4812), .A2(n4810), .ZN(n8587) );
  OR2_X1 U5525 ( .A1(n6110), .A2(n7830), .ZN(n6123) );
  OR2_X1 U5526 ( .A1(n6081), .A2(n6080), .ZN(n6098) );
  NAND2_X1 U5527 ( .A1(n6096), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6110) );
  INV_X1 U5528 ( .A(n6098), .ZN(n6096) );
  AND2_X1 U5529 ( .A1(n8147), .A2(n8149), .ZN(n8241) );
  NAND2_X1 U5530 ( .A1(n7612), .A2(n4410), .ZN(n8613) );
  AND2_X1 U5531 ( .A1(n7612), .A2(n4717), .ZN(n7781) );
  INV_X1 U5532 ( .A(n4786), .ZN(n4785) );
  OAI21_X1 U5533 ( .B1(n8134), .B2(n4787), .A(n8139), .ZN(n4786) );
  AND2_X1 U5534 ( .A1(n7612), .A2(n9518), .ZN(n7678) );
  INV_X1 U5535 ( .A(n7608), .ZN(n7609) );
  NAND2_X1 U5536 ( .A1(n7609), .A2(n8134), .ZN(n7674) );
  NOR2_X1 U5537 ( .A1(n7565), .A2(n7602), .ZN(n7612) );
  INV_X1 U5538 ( .A(n4794), .ZN(n7554) );
  INV_X1 U5539 ( .A(n4790), .ZN(n4789) );
  NOR2_X1 U5540 ( .A1(n8053), .A2(n4961), .ZN(n4960) );
  INV_X1 U5541 ( .A(n7464), .ZN(n4961) );
  NOR2_X1 U5542 ( .A1(n7451), .A2(n9843), .ZN(n4719) );
  NAND2_X1 U5543 ( .A1(n4720), .A2(n4721), .ZN(n7448) );
  NOR2_X1 U5544 ( .A1(n7451), .A2(n9731), .ZN(n4720) );
  NAND2_X1 U5545 ( .A1(n7345), .A2(n8112), .ZN(n7443) );
  NAND2_X1 U5546 ( .A1(n7349), .A2(n7348), .ZN(n7453) );
  NAND2_X1 U5547 ( .A1(n7228), .A2(n7227), .ZN(n7231) );
  NOR2_X1 U5548 ( .A1(n4722), .A2(n9731), .ZN(n7344) );
  INV_X1 U5549 ( .A(n4806), .ZN(n4805) );
  NOR2_X1 U5550 ( .A1(n9731), .A2(n7226), .ZN(n7241) );
  OR2_X1 U5551 ( .A1(n9730), .A2(n9727), .ZN(n9731) );
  AND2_X1 U5552 ( .A1(n9760), .A2(n9821), .ZN(n7030) );
  NAND2_X1 U5553 ( .A1(n8093), .A2(n4715), .ZN(n9758) );
  INV_X1 U5554 ( .A(n6899), .ZN(n4715) );
  NAND2_X1 U5555 ( .A1(n6895), .A2(n6894), .ZN(n9781) );
  OR2_X1 U5556 ( .A1(n6293), .A2(n6292), .ZN(n9838) );
  AND2_X1 U5557 ( .A1(n6653), .A2(n6305), .ZN(n9844) );
  NOR2_X1 U5558 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5800) );
  NAND2_X1 U5559 ( .A1(n4878), .A2(n4875), .ZN(n8796) );
  AND2_X1 U5560 ( .A1(n4876), .A2(n4479), .ZN(n4875) );
  NAND2_X1 U5561 ( .A1(n4612), .A2(n4611), .ZN(n4878) );
  AOI21_X1 U5562 ( .B1(n4607), .B2(n4610), .A(n4479), .ZN(n4605) );
  INV_X1 U5563 ( .A(n4611), .ZN(n4610) );
  AND2_X1 U5564 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5470) );
  NOR2_X1 U5565 ( .A1(n5351), .A2(n5339), .ZN(n5340) );
  NAND2_X1 U5566 ( .A1(n6825), .A2(n7208), .ZN(n6786) );
  AND2_X1 U5567 ( .A1(n6839), .A2(n6795), .ZN(n7150) );
  NAND2_X1 U5568 ( .A1(n4862), .A2(n4864), .ZN(n4861) );
  AND2_X1 U5569 ( .A1(n5257), .A2(n5122), .ZN(n5227) );
  NOR2_X1 U5570 ( .A1(n5440), .A2(n5439), .ZN(n5490) );
  INV_X1 U5571 ( .A(n9186), .ZN(n9103) );
  INV_X1 U5572 ( .A(n5707), .ZN(n4742) );
  NOR2_X1 U5573 ( .A1(n4533), .A2(n4432), .ZN(n5708) );
  NAND2_X1 U5574 ( .A1(n5620), .A2(n4741), .ZN(n4740) );
  NOR2_X1 U5575 ( .A1(n9354), .A2(n4562), .ZN(n4741) );
  NAND2_X1 U5576 ( .A1(n4532), .A2(n6700), .ZN(n4531) );
  NAND2_X1 U5577 ( .A1(n5716), .A2(n9607), .ZN(n4532) );
  OR2_X1 U5578 ( .A1(n4526), .A2(n5715), .ZN(n4524) );
  NOR3_X1 U5579 ( .A1(n6334), .A2(n8988), .A3(n8986), .ZN(n6867) );
  NAND2_X1 U5580 ( .A1(n6569), .A2(n6568), .ZN(n6337) );
  OR2_X1 U5581 ( .A1(n9559), .A2(n4571), .ZN(n9573) );
  NOR2_X1 U5582 ( .A1(n6326), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4571) );
  NAND2_X1 U5583 ( .A1(n9573), .A2(n9572), .ZN(n9571) );
  NOR2_X1 U5584 ( .A1(n6342), .A2(n6631), .ZN(n6438) );
  AOI21_X1 U5585 ( .B1(n5489), .B2(n6440), .A(n6436), .ZN(n6498) );
  NOR2_X1 U5586 ( .A1(n6360), .A2(n4480), .ZN(n9594) );
  NOR2_X1 U5587 ( .A1(n9594), .A2(n9593), .ZN(n9592) );
  NAND2_X1 U5588 ( .A1(n9588), .A2(n4492), .ZN(n9004) );
  NOR2_X1 U5589 ( .A1(n9592), .A2(n4579), .ZN(n8997) );
  AND2_X1 U5590 ( .A1(n6370), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4579) );
  NAND2_X1 U5591 ( .A1(n9004), .A2(n9005), .ZN(n9003) );
  NAND2_X1 U5592 ( .A1(n6913), .A2(n4491), .ZN(n7081) );
  NAND2_X1 U5593 ( .A1(n7081), .A2(n7082), .ZN(n7080) );
  NOR2_X1 U5594 ( .A1(n9032), .A2(n9031), .ZN(n9049) );
  AND2_X1 U5595 ( .A1(n9176), .A2(n4470), .ZN(n9079) );
  NAND2_X1 U5596 ( .A1(n9367), .A2(n9168), .ZN(n9129) );
  INV_X1 U5597 ( .A(n9132), .ZN(n9168) );
  NOR2_X1 U5598 ( .A1(n4834), .A2(n9167), .ZN(n4831) );
  NAND2_X1 U5599 ( .A1(n4832), .A2(n4833), .ZN(n9166) );
  NOR2_X1 U5600 ( .A1(n9192), .A2(n9377), .ZN(n9176) );
  NAND2_X1 U5601 ( .A1(n9211), .A2(n9198), .ZN(n9192) );
  NAND2_X1 U5602 ( .A1(n4837), .A2(n4835), .ZN(n9208) );
  AOI21_X1 U5603 ( .B1(n4838), .B2(n4843), .A(n4836), .ZN(n4835) );
  AND2_X1 U5604 ( .A1(n4839), .A2(n4841), .ZN(n4838) );
  NAND2_X1 U5605 ( .A1(n9280), .A2(n4700), .ZN(n9220) );
  AND2_X1 U5606 ( .A1(n4411), .A2(n9225), .ZN(n4700) );
  NAND2_X1 U5607 ( .A1(n4663), .A2(n4483), .ZN(n9219) );
  NAND2_X1 U5608 ( .A1(n4918), .A2(n4439), .ZN(n4663) );
  NAND2_X1 U5609 ( .A1(n9280), .A2(n4701), .ZN(n9247) );
  NAND2_X1 U5610 ( .A1(n9280), .A2(n9267), .ZN(n9264) );
  NAND2_X1 U5611 ( .A1(n4816), .A2(n4815), .ZN(n9286) );
  AOI21_X1 U5612 ( .B1(n4408), .B2(n4820), .A(n5663), .ZN(n4815) );
  AND2_X1 U5613 ( .A1(n9296), .A2(n9284), .ZN(n9280) );
  OR2_X1 U5614 ( .A1(n9335), .A2(n9426), .ZN(n9317) );
  NOR2_X1 U5615 ( .A1(n5378), .A2(n5121), .ZN(n5380) );
  AND2_X1 U5616 ( .A1(n5380), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U5617 ( .A1(n9502), .A2(n4696), .ZN(n7762) );
  AND2_X1 U5618 ( .A1(n4407), .A2(n4697), .ZN(n4696) );
  NOR2_X1 U5619 ( .A1(n7762), .A2(n9084), .ZN(n9334) );
  INV_X1 U5620 ( .A(n8973), .ZN(n8788) );
  NAND2_X1 U5621 ( .A1(n7700), .A2(n4446), .ZN(n7714) );
  NAND2_X1 U5622 ( .A1(n9502), .A2(n4407), .ZN(n7726) );
  NAND2_X1 U5623 ( .A1(n4847), .A2(n4406), .ZN(n7717) );
  AND2_X1 U5624 ( .A1(n4847), .A2(n7693), .ZN(n7718) );
  NAND2_X1 U5625 ( .A1(n4848), .A2(n4849), .ZN(n4847) );
  NAND2_X1 U5626 ( .A1(n9502), .A2(n4699), .ZN(n7724) );
  AND2_X1 U5627 ( .A1(n9502), .A2(n9542), .ZN(n7664) );
  AND2_X1 U5628 ( .A1(n5340), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U5629 ( .A1(n7639), .A2(n7638), .ZN(n7692) );
  NAND2_X1 U5630 ( .A1(n7513), .A2(n4856), .ZN(n7639) );
  AND2_X1 U5631 ( .A1(n4858), .A2(n7512), .ZN(n4856) );
  INV_X1 U5632 ( .A(n7637), .ZN(n4858) );
  NAND2_X1 U5633 ( .A1(n4703), .A2(n4404), .ZN(n7516) );
  NAND2_X1 U5634 ( .A1(n7513), .A2(n7512), .ZN(n9485) );
  AOI21_X1 U5635 ( .B1(n4928), .B2(n4927), .A(n4450), .ZN(n4926) );
  OR2_X1 U5636 ( .A1(n5492), .A2(n5349), .ZN(n5351) );
  NAND2_X1 U5637 ( .A1(n7420), .A2(n4857), .ZN(n7513) );
  NOR2_X1 U5638 ( .A1(n7421), .A2(n5633), .ZN(n4857) );
  NAND2_X1 U5639 ( .A1(n7420), .A2(n7419), .ZN(n7422) );
  NOR2_X1 U5640 ( .A1(n7321), .A2(n7326), .ZN(n7322) );
  NOR2_X1 U5641 ( .A1(n7321), .A2(n4704), .ZN(n7429) );
  INV_X1 U5642 ( .A(n4705), .ZN(n4704) );
  NAND2_X1 U5643 ( .A1(n7281), .A2(n7280), .ZN(n7417) );
  AND3_X1 U5644 ( .A1(n5438), .A2(n5437), .A3(n5436), .ZN(n9603) );
  OAI21_X1 U5645 ( .B1(n7268), .B2(n5628), .A(n5629), .ZN(n7067) );
  INV_X1 U5646 ( .A(n7066), .ZN(n7062) );
  INV_X1 U5647 ( .A(n9654), .ZN(n7265) );
  NAND2_X1 U5648 ( .A1(n6975), .A2(n5627), .ZN(n7268) );
  NOR2_X1 U5649 ( .A1(n6973), .A2(n7303), .ZN(n7260) );
  NAND2_X1 U5650 ( .A1(n6977), .A2(n6976), .ZN(n6975) );
  NAND2_X1 U5651 ( .A1(n4693), .A2(n9649), .ZN(n7303) );
  INV_X1 U5652 ( .A(n7301), .ZN(n4693) );
  XNOR2_X1 U5653 ( .A(n6826), .B(n9649), .ZN(n7293) );
  OAI21_X1 U5654 ( .B1(n7154), .B2(n4828), .A(n5409), .ZN(n7292) );
  AND2_X1 U5655 ( .A1(n6791), .A2(n7208), .ZN(n7146) );
  OR2_X1 U5656 ( .A1(n6701), .A2(n6700), .ZN(n7065) );
  CLKBUF_X1 U5657 ( .A(n6965), .Z(n7154) );
  INV_X1 U5658 ( .A(n4828), .ZN(n7153) );
  NAND2_X1 U5659 ( .A1(n5165), .A2(n5164), .ZN(n9382) );
  INV_X1 U5660 ( .A(n4664), .ZN(n9408) );
  INV_X1 U5661 ( .A(n9668), .ZN(n9503) );
  AND2_X1 U5662 ( .A1(n6405), .A2(n6407), .ZN(n9616) );
  XNOR2_X1 U5663 ( .A(n4745), .B(n5580), .ZN(n8032) );
  OAI21_X1 U5664 ( .B1(n5575), .B2(n4746), .A(n5578), .ZN(n4745) );
  OR2_X1 U5665 ( .A1(n5118), .A2(n5449), .ZN(n5115) );
  XNOR2_X1 U5666 ( .A(n5575), .B(SI_30_), .ZN(n8022) );
  XNOR2_X1 U5667 ( .A(n5570), .B(n5102), .ZN(n8760) );
  OAI21_X1 U5668 ( .B1(n5098), .B2(n4769), .A(n4420), .ZN(n5570) );
  NAND2_X1 U5669 ( .A1(n4694), .A2(n5277), .ZN(n4569) );
  XNOR2_X1 U5670 ( .A(n5522), .B(n5521), .ZN(n7819) );
  NAND2_X1 U5671 ( .A1(n4749), .A2(n5051), .ZN(n5219) );
  NAND2_X1 U5672 ( .A1(n5047), .A2(n4753), .ZN(n4749) );
  AND2_X1 U5673 ( .A1(n5267), .A2(n5205), .ZN(n5252) );
  NAND2_X1 U5674 ( .A1(n4773), .A2(n4778), .ZN(n5276) );
  NAND2_X1 U5675 ( .A1(n5306), .A2(n4780), .ZN(n4773) );
  NAND2_X1 U5676 ( .A1(n4735), .A2(n5007), .ZN(n5333) );
  OR2_X1 U5677 ( .A1(n5358), .A2(n5357), .ZN(n4735) );
  OAI21_X1 U5678 ( .B1(n4997), .B2(n4658), .A(n4657), .ZN(n5498) );
  XNOR2_X1 U5679 ( .A(n4994), .B(SI_5_), .ZN(n5433) );
  INV_X1 U5680 ( .A(n4986), .ZN(n4671) );
  NAND2_X1 U5681 ( .A1(n4581), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5422) );
  INV_X1 U5682 ( .A(n5420), .ZN(n4581) );
  NAND2_X1 U5683 ( .A1(n6767), .A2(n5922), .ZN(n6942) );
  AND2_X1 U5684 ( .A1(n6244), .A2(n6233), .ZN(n8455) );
  NAND2_X1 U5685 ( .A1(n8766), .A2(n6204), .ZN(n6230) );
  AND2_X1 U5686 ( .A1(n4915), .A2(n4433), .ZN(n7592) );
  NAND2_X1 U5687 ( .A1(n6173), .A2(n6172), .ZN(n8674) );
  AND4_X1 U5688 ( .A1(n5968), .A2(n5967), .A3(n5966), .A4(n5965), .ZN(n7224)
         );
  AND4_X1 U5689 ( .A1(n6115), .A2(n6114), .A3(n6113), .A4(n6112), .ZN(n8591)
         );
  NAND2_X1 U5690 ( .A1(n4888), .A2(n4889), .ZN(n8288) );
  OR2_X1 U5691 ( .A1(n7002), .A2(n6759), .ZN(n5839) );
  AND3_X1 U5692 ( .A1(n6141), .A2(n6140), .A3(n6139), .ZN(n8592) );
  NAND2_X1 U5693 ( .A1(n6012), .A2(n6011), .ZN(n7559) );
  AND2_X1 U5694 ( .A1(n6201), .A2(n6200), .ZN(n8518) );
  AND2_X1 U5695 ( .A1(n6311), .A2(n6310), .ZN(n8332) );
  NAND2_X1 U5696 ( .A1(n4898), .A2(n4897), .ZN(n7790) );
  NAND2_X1 U5697 ( .A1(n6079), .A2(n6078), .ZN(n7798) );
  AND4_X1 U5698 ( .A1(n6086), .A2(n6085), .A3(n6084), .A4(n6083), .ZN(n8359)
         );
  AND3_X1 U5699 ( .A1(n6127), .A2(n6126), .A3(n6125), .ZN(n8602) );
  NAND2_X1 U5700 ( .A1(n7405), .A2(n6028), .ZN(n7435) );
  NAND2_X1 U5701 ( .A1(n6163), .A2(n6162), .ZN(n8537) );
  OR2_X1 U5702 ( .A1(n7627), .A2(n9745), .ZN(n8330) );
  NAND2_X1 U5703 ( .A1(n4891), .A2(n4894), .ZN(n7829) );
  OR2_X1 U5704 ( .A1(n7813), .A2(n7812), .ZN(n4891) );
  NAND2_X1 U5705 ( .A1(n5905), .A2(n5904), .ZN(n6769) );
  NAND2_X1 U5706 ( .A1(n4908), .A2(n4904), .ZN(n8341) );
  INV_X1 U5707 ( .A(n4907), .ZN(n4904) );
  OAI21_X1 U5708 ( .B1(n8036), .B2(n8213), .A(n8216), .ZN(n8037) );
  AND2_X1 U5709 ( .A1(n6188), .A2(n6187), .ZN(n8535) );
  AND2_X1 U5710 ( .A1(n6170), .A2(n6169), .ZN(n8551) );
  OR2_X1 U5711 ( .A1(n6318), .A2(n6460), .ZN(n8354) );
  AOI21_X1 U5712 ( .B1(n6539), .B2(n6522), .A(n6521), .ZN(n6615) );
  NOR2_X1 U5713 ( .A1(n6683), .A2(n6682), .ZN(n8392) );
  AOI21_X1 U5714 ( .B1(n6948), .B2(n6955), .A(n6947), .ZN(n6951) );
  AND2_X1 U5715 ( .A1(n6484), .A2(n6483), .ZN(n9711) );
  NAND2_X1 U5716 ( .A1(n7182), .A2(n4505), .ZN(n7336) );
  AND2_X1 U5717 ( .A1(n7180), .A2(n4496), .ZN(n4505) );
  NAND2_X1 U5718 ( .A1(n7336), .A2(n4496), .ZN(n7339) );
  XNOR2_X1 U5719 ( .A(n8420), .B(n4714), .ZN(n8636) );
  AOI21_X1 U5720 ( .B1(n8460), .B2(n9770), .A(n8263), .ZN(n8264) );
  NAND2_X1 U5721 ( .A1(n8433), .A2(n4973), .ZN(n4949) );
  NAND2_X1 U5722 ( .A1(n4511), .A2(n4510), .ZN(n4509) );
  XNOR2_X1 U5723 ( .A(n8459), .B(n8458), .ZN(n4512) );
  NAND2_X1 U5724 ( .A1(n8461), .A2(n9770), .ZN(n4510) );
  NAND2_X1 U5725 ( .A1(n6207), .A2(n6206), .ZN(n8664) );
  NAND2_X1 U5726 ( .A1(n4940), .A2(n4944), .ZN(n8513) );
  OAI21_X1 U5727 ( .B1(n8546), .B2(n4943), .A(n4941), .ZN(n8511) );
  NAND2_X1 U5728 ( .A1(n8546), .A2(n4945), .ZN(n4940) );
  AND2_X1 U5729 ( .A1(n4947), .A2(n4424), .ZN(n8528) );
  NAND2_X1 U5730 ( .A1(n8546), .A2(n8247), .ZN(n4947) );
  NAND2_X1 U5731 ( .A1(n6143), .A2(n6142), .ZN(n8559) );
  NAND2_X1 U5732 ( .A1(n4951), .A2(n4957), .ZN(n8581) );
  NAND2_X1 U5733 ( .A1(n8616), .A2(n4955), .ZN(n4951) );
  NAND2_X1 U5734 ( .A1(n8616), .A2(n8243), .ZN(n8597) );
  NAND2_X1 U5735 ( .A1(n4788), .A2(n8119), .ZN(n7460) );
  NAND2_X1 U5736 ( .A1(n7345), .A2(n4792), .ZN(n4788) );
  NAND2_X1 U5737 ( .A1(n7110), .A2(n4806), .ZN(n9723) );
  AND2_X1 U5738 ( .A1(n8077), .A2(n8080), .ZN(n9768) );
  INV_X1 U5739 ( .A(n9757), .ZN(n9726) );
  INV_X1 U5740 ( .A(n9879), .ZN(n9877) );
  AOI21_X1 U5741 ( .B1(n8636), .B2(n9845), .A(n8639), .ZN(n8714) );
  INV_X1 U5742 ( .A(n8429), .ZN(n8719) );
  INV_X1 U5743 ( .A(n8537), .ZN(n8739) );
  AND2_X1 U5744 ( .A1(n6423), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9794) );
  XNOR2_X1 U5745 ( .A(n6267), .B(n6266), .ZN(n7687) );
  NAND2_X1 U5746 ( .A1(n5806), .A2(n4425), .ZN(n6106) );
  INV_X1 U5747 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6387) );
  INV_X1 U5748 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6383) );
  INV_X1 U5749 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6381) );
  CLKBUF_X1 U5750 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n9691) );
  NAND2_X1 U5751 ( .A1(n4874), .A2(n7371), .ZN(n7525) );
  OR2_X1 U5752 ( .A1(n7373), .A2(n7372), .ZN(n4874) );
  NAND2_X1 U5753 ( .A1(n5209), .A2(n5208), .ZN(n9415) );
  NAND2_X1 U5754 ( .A1(n4604), .A2(n4603), .ZN(n4602) );
  NAND2_X1 U5755 ( .A1(n4585), .A2(n7871), .ZN(n8831) );
  NAND2_X1 U5756 ( .A1(n4487), .A2(n8849), .ZN(n8859) );
  NAND2_X1 U5757 ( .A1(n4594), .A2(n4592), .ZN(n8877) );
  NAND2_X1 U5758 ( .A1(n7845), .A2(n4595), .ZN(n4594) );
  NAND2_X1 U5759 ( .A1(n7845), .A2(n4593), .ZN(n4592) );
  INV_X1 U5760 ( .A(n8974), .ZN(n8906) );
  NOR2_X1 U5761 ( .A1(n8901), .A2(n4881), .ZN(n4880) );
  INV_X1 U5762 ( .A(n7882), .ZN(n4881) );
  NAND2_X1 U5763 ( .A1(n8829), .A2(n7882), .ZN(n8900) );
  NAND2_X1 U5764 ( .A1(n7951), .A2(n7950), .ZN(n8912) );
  AND2_X1 U5765 ( .A1(n4612), .A2(n4614), .ZN(n7951) );
  INV_X1 U5766 ( .A(n8921), .ZN(n8960) );
  NAND2_X1 U5767 ( .A1(n8848), .A2(n4866), .ZN(n4615) );
  AND2_X1 U5768 ( .A1(n8945), .A2(n8942), .ZN(n7976) );
  OR2_X1 U5769 ( .A1(n5201), .A2(n5200), .ZN(n9289) );
  AOI21_X1 U5770 ( .B1(n6332), .B2(n9562), .A(n9553), .ZN(n9578) );
  NOR2_X1 U5771 ( .A1(n6628), .A2(n4428), .ZN(n6434) );
  NAND2_X1 U5772 ( .A1(n6434), .A2(n6435), .ZN(n6433) );
  NAND2_X1 U5773 ( .A1(n6433), .A2(n4574), .ZN(n6493) );
  OR2_X1 U5774 ( .A1(n6343), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4574) );
  NAND2_X1 U5775 ( .A1(n6493), .A2(n6494), .ZN(n6492) );
  INV_X1 U5776 ( .A(n4578), .ZN(n6919) );
  INV_X1 U5777 ( .A(n4576), .ZN(n7085) );
  XNOR2_X1 U5778 ( .A(n9017), .B(n9016), .ZN(n6374) );
  NOR2_X1 U5779 ( .A1(n9011), .A2(n9012), .ZN(n9015) );
  INV_X1 U5780 ( .A(n4573), .ZN(n9029) );
  AOI21_X1 U5781 ( .B1(n9050), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9044), .ZN(
        n9045) );
  AOI21_X1 U5782 ( .B1(n9368), .B2(n9313), .A(n9157), .ZN(n4852) );
  AND2_X1 U5783 ( .A1(n4855), .A2(n4854), .ZN(n9370) );
  AOI21_X1 U5784 ( .B1(n9155), .B2(n9305), .A(n4481), .ZN(n4854) );
  NAND2_X1 U5785 ( .A1(n9156), .A2(n9308), .ZN(n4855) );
  INV_X1 U5786 ( .A(n9373), .ZN(n9165) );
  NAND2_X1 U5787 ( .A1(n4672), .A2(n9101), .ZN(n9158) );
  NAND2_X1 U5788 ( .A1(n4933), .A2(n9099), .ZN(n9175) );
  NAND2_X1 U5789 ( .A1(n5144), .A2(n5143), .ZN(n9389) );
  NAND2_X1 U5790 ( .A1(n4840), .A2(n4841), .ZN(n9226) );
  OR2_X1 U5791 ( .A1(n9251), .A2(n4843), .ZN(n4840) );
  AND2_X1 U5792 ( .A1(n4844), .A2(n5672), .ZN(n9235) );
  INV_X1 U5793 ( .A(n4918), .ZN(n9234) );
  NAND2_X1 U5794 ( .A1(n4683), .A2(n4684), .ZN(n9279) );
  NAND2_X1 U5795 ( .A1(n4686), .A2(n4689), .ZN(n9294) );
  OR2_X1 U5796 ( .A1(n4920), .A2(n9088), .ZN(n4686) );
  NAND2_X1 U5797 ( .A1(n4821), .A2(n4822), .ZN(n9325) );
  AND2_X1 U5798 ( .A1(n4920), .A2(n4426), .ZN(n9316) );
  OAI21_X1 U5799 ( .B1(n9109), .B2(n9108), .A(n9107), .ZN(n9345) );
  NAND2_X1 U5800 ( .A1(n4923), .A2(n4924), .ZN(n9332) );
  INV_X1 U5801 ( .A(n4920), .ZN(n9331) );
  NAND2_X1 U5802 ( .A1(n7751), .A2(n7750), .ZN(n9086) );
  NAND2_X1 U5803 ( .A1(n5324), .A2(n5323), .ZN(n9501) );
  NAND2_X1 U5804 ( .A1(n7259), .A2(n7061), .ZN(n7063) );
  INV_X1 U5805 ( .A(n9338), .ZN(n9500) );
  NAND2_X1 U5806 ( .A1(n5119), .A2(n9463), .ZN(n9470) );
  OR2_X1 U5807 ( .A1(n5767), .A2(n4469), .ZN(n5116) );
  NAND2_X1 U5808 ( .A1(n5767), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5774) );
  XNOR2_X1 U5809 ( .A(n5152), .B(n5151), .ZN(n7542) );
  NAND2_X1 U5810 ( .A1(n5623), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5624) );
  CLKBUF_X1 U5811 ( .A(n6978), .Z(n9607) );
  INV_X1 U5812 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9976) );
  INV_X1 U5813 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10091) );
  INV_X1 U5814 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6394) );
  INV_X1 U5815 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U5816 ( .A1(n4987), .A2(n4986), .ZN(n5462) );
  INV_X1 U5817 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U5818 ( .A1(n5463), .A2(n4580), .ZN(n6861) );
  OR2_X1 U5819 ( .A1(n5422), .A2(n5421), .ZN(n4580) );
  NAND2_X1 U5820 ( .A1(n4913), .A2(n5957), .ZN(n7096) );
  NAND2_X1 U5821 ( .A1(n4503), .A2(n4499), .ZN(n8417) );
  OR2_X1 U5822 ( .A1(n8413), .A2(n4500), .ZN(n4499) );
  OAI21_X1 U5823 ( .B1(n8714), .B2(n9860), .A(n4711), .ZN(P2_U3519) );
  AOI21_X1 U5824 ( .B1(n8421), .B2(n4713), .A(n4712), .ZN(n4711) );
  NOR2_X1 U5825 ( .A1(n9861), .A2(n8715), .ZN(n4712) );
  INV_X1 U5826 ( .A(n8754), .ZN(n4713) );
  NAND2_X1 U5827 ( .A1(n5719), .A2(n4528), .ZN(n4520) );
  NOR2_X1 U5828 ( .A1(n5719), .A2(n4526), .ZN(n4519) );
  NAND2_X1 U5829 ( .A1(n4853), .A2(n4850), .ZN(P1_U3263) );
  OR2_X1 U5830 ( .A1(n9370), .A2(n4393), .ZN(n4853) );
  INV_X1 U5831 ( .A(n4851), .ZN(n4850) );
  OAI21_X1 U5832 ( .B1(n9371), .B2(n9351), .A(n4852), .ZN(n4851) );
  OAI21_X1 U5833 ( .B1(n8007), .B2(n9473), .A(n4868), .ZN(P1_U3331) );
  INV_X1 U5834 ( .A(n4869), .ZN(n4868) );
  OAI22_X1 U5835 ( .A1(n5714), .A2(P1_U3084), .B1(n9479), .B2(n8008), .ZN(
        n4869) );
  NOR2_X1 U5836 ( .A1(n5767), .A2(n4935), .ZN(n5118) );
  AND2_X1 U5837 ( .A1(n9667), .A2(n4705), .ZN(n4404) );
  AND2_X1 U5838 ( .A1(n4427), .A2(n8849), .ZN(n4866) );
  NAND2_X1 U5839 ( .A1(n8696), .A2(n8566), .ZN(n4405) );
  AND2_X1 U5840 ( .A1(n7693), .A2(n7719), .ZN(n4406) );
  AND2_X1 U5841 ( .A1(n4699), .A2(n4698), .ZN(n4407) );
  AND2_X1 U5842 ( .A1(n5664), .A2(n4817), .ZN(n4408) );
  AND3_X1 U5843 ( .A1(n4622), .A2(n4629), .A3(n4621), .ZN(n4409) );
  AND2_X1 U5844 ( .A1(n4717), .A2(n8755), .ZN(n4410) );
  INV_X1 U5845 ( .A(n8512), .ZN(n4942) );
  INV_X1 U5846 ( .A(n7280), .ZN(n4927) );
  OR2_X1 U5847 ( .A1(n8652), .A2(n8471), .ZN(n8018) );
  NAND2_X1 U5848 ( .A1(n6065), .A2(n6064), .ZN(n8141) );
  AND2_X1 U5849 ( .A1(n4701), .A2(n9244), .ZN(n4411) );
  AND2_X1 U5850 ( .A1(n9828), .A2(n8368), .ZN(n4412) );
  AND2_X1 U5851 ( .A1(n4724), .A2(n4723), .ZN(n4413) );
  AND2_X1 U5852 ( .A1(n9105), .A2(n9104), .ZN(n4414) );
  AND2_X1 U5853 ( .A1(n4556), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4415) );
  NAND2_X1 U5854 ( .A1(n8369), .A2(n7115), .ZN(n4416) );
  INV_X1 U5855 ( .A(n4870), .ZN(n4603) );
  OR2_X1 U5856 ( .A1(n7372), .A2(n4873), .ZN(n4870) );
  NAND2_X1 U5857 ( .A1(n8129), .A2(n8128), .ZN(n4417) );
  AND2_X1 U5858 ( .A1(n7062), .A2(n7061), .ZN(n4418) );
  AND2_X1 U5859 ( .A1(n4706), .A2(n4404), .ZN(n4419) );
  AND2_X1 U5860 ( .A1(n8719), .A2(n8352), .ZN(n8211) );
  NAND2_X1 U5861 ( .A1(n8034), .A2(n8033), .ZN(n8421) );
  INV_X1 U5862 ( .A(n8421), .ZN(n4714) );
  NAND2_X1 U5863 ( .A1(n7417), .A2(n4928), .ZN(n7511) );
  AND2_X1 U5864 ( .A1(n4768), .A2(n5101), .ZN(n4420) );
  INV_X1 U5865 ( .A(n4872), .ZN(n4871) );
  NAND2_X2 U5866 ( .A1(n5408), .A2(n4556), .ZN(n5419) );
  NAND2_X1 U5867 ( .A1(n6135), .A2(n6134), .ZN(n8689) );
  OAI211_X1 U5868 ( .C1(n6041), .C2(n6389), .A(n5856), .B(n5855), .ZN(n9806)
         );
  AND2_X1 U5869 ( .A1(n4989), .A2(SI_3_), .ZN(n4421) );
  AOI21_X1 U5870 ( .B1(n8760), .B2(n5581), .A(n5113), .ZN(n9361) );
  AND2_X1 U5871 ( .A1(n4999), .A2(SI_6_), .ZN(n4422) );
  NAND2_X1 U5872 ( .A1(n8841), .A2(n8842), .ZN(n8840) );
  INV_X1 U5873 ( .A(n4929), .ZN(n4928) );
  NAND2_X1 U5874 ( .A1(n7421), .A2(n7416), .ZN(n4929) );
  XNOR2_X1 U5875 ( .A(n5115), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5123) );
  INV_X1 U5876 ( .A(n8112), .ZN(n4793) );
  XOR2_X1 U5877 ( .A(n7928), .B(n7992), .Z(n4423) );
  NAND2_X1 U5878 ( .A1(n8559), .A2(n8567), .ZN(n4424) );
  AND2_X1 U5879 ( .A1(n5807), .A2(n4647), .ZN(n4425) );
  NAND2_X1 U5880 ( .A1(n9431), .A2(n9087), .ZN(n4426) );
  NAND2_X1 U5881 ( .A1(n7925), .A2(n7924), .ZN(n4427) );
  OR2_X1 U5882 ( .A1(n9373), .A2(n9103), .ZN(n5704) );
  AND2_X1 U5883 ( .A1(n6341), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4428) );
  NAND2_X1 U5884 ( .A1(n6095), .A2(n6094), .ZN(n8706) );
  OR2_X1 U5885 ( .A1(n7951), .A2(n7950), .ZN(n4429) );
  AND2_X1 U5886 ( .A1(n8179), .A2(n8214), .ZN(n4430) );
  INV_X1 U5887 ( .A(n5109), .ZN(n4695) );
  INV_X1 U5888 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5818) );
  AND2_X1 U5889 ( .A1(n8913), .A2(n4879), .ZN(n4431) );
  OR2_X1 U5890 ( .A1(n5706), .A2(n6701), .ZN(n4432) );
  NAND2_X1 U5891 ( .A1(n6192), .A2(n6191), .ZN(n8505) );
  NAND2_X1 U5892 ( .A1(n4812), .A2(n8156), .ZN(n8586) );
  NAND2_X1 U5893 ( .A1(n8204), .A2(n8205), .ZN(n8257) );
  INV_X1 U5894 ( .A(n8257), .ZN(n4641) );
  NAND2_X1 U5895 ( .A1(n5800), .A2(n4962), .ZN(n5853) );
  NAND2_X1 U5896 ( .A1(n6040), .A2(n6039), .ZN(n4433) );
  AND2_X1 U5897 ( .A1(n5104), .A2(n4932), .ZN(n4434) );
  OR2_X1 U5898 ( .A1(n6830), .A2(n6829), .ZN(n4435) );
  INV_X1 U5899 ( .A(n8045), .ZN(n7021) );
  NAND2_X1 U5900 ( .A1(n8898), .A2(n8973), .ZN(n4436) );
  AND2_X1 U5901 ( .A1(n8079), .A2(n8080), .ZN(n4437) );
  AND2_X1 U5902 ( .A1(n4889), .A2(n4887), .ZN(n4438) );
  NAND2_X1 U5903 ( .A1(n5572), .A2(n5571), .ZN(n9080) );
  INV_X1 U5904 ( .A(n9080), .ZN(n9359) );
  OR2_X1 U5905 ( .A1(n9399), .A2(n9228), .ZN(n4439) );
  INV_X1 U5906 ( .A(n7311), .ZN(n7313) );
  NAND2_X1 U5907 ( .A1(n6046), .A2(n6045), .ZN(n7671) );
  NAND2_X1 U5908 ( .A1(n5195), .A2(n5194), .ZN(n9411) );
  OR2_X1 U5909 ( .A1(n8604), .A2(n8591), .ZN(n8156) );
  INV_X1 U5910 ( .A(n8156), .ZN(n4811) );
  AND2_X1 U5911 ( .A1(n9855), .A2(n8363), .ZN(n8127) );
  NOR2_X1 U5912 ( .A1(n9085), .A2(n4925), .ZN(n4440) );
  AND2_X1 U5913 ( .A1(n7419), .A2(n5727), .ZN(n4441) );
  INV_X1 U5914 ( .A(n9244), .ZN(n9399) );
  AND2_X1 U5915 ( .A1(n5174), .A2(n5173), .ZN(n9244) );
  AND2_X1 U5916 ( .A1(n8145), .A2(n8241), .ZN(n4442) );
  NAND2_X1 U5917 ( .A1(n8519), .A2(n4726), .ZN(n4727) );
  OR2_X1 U5918 ( .A1(n7621), .A2(n7620), .ZN(n4443) );
  AND2_X1 U5919 ( .A1(n4832), .A2(n4831), .ZN(n4444) );
  NAND2_X1 U5920 ( .A1(n6216), .A2(n6215), .ZN(n8477) );
  INV_X1 U5921 ( .A(n4820), .ZN(n4819) );
  NAND2_X1 U5922 ( .A1(n4822), .A2(n5598), .ZN(n4820) );
  AND2_X1 U5923 ( .A1(n5705), .A2(n9129), .ZN(n9154) );
  OR2_X1 U5924 ( .A1(n8458), .A2(n8457), .ZN(n4445) );
  NAND2_X1 U5925 ( .A1(n7702), .A2(n7701), .ZN(n4446) );
  INV_X1 U5926 ( .A(n7691), .ZN(n4849) );
  INV_X1 U5927 ( .A(n4946), .ZN(n4945) );
  NAND2_X1 U5928 ( .A1(n4948), .A2(n8247), .ZN(n4946) );
  AND2_X1 U5929 ( .A1(n4673), .A2(n9099), .ZN(n4447) );
  AND2_X1 U5930 ( .A1(n7881), .A2(n7871), .ZN(n4448) );
  AND2_X1 U5931 ( .A1(n7229), .A2(n7227), .ZN(n4449) );
  INV_X1 U5932 ( .A(n4834), .ZN(n4833) );
  OAI21_X1 U5933 ( .B1(n9127), .B2(n5626), .A(n9126), .ZN(n4834) );
  AND2_X1 U5934 ( .A1(n8978), .A2(n7537), .ZN(n4450) );
  OR2_X1 U5935 ( .A1(n8689), .A2(n8592), .ZN(n8013) );
  NAND2_X1 U5936 ( .A1(n9405), .A2(n9092), .ZN(n4451) );
  AND2_X1 U5937 ( .A1(n8130), .A2(n8129), .ZN(n8053) );
  AND2_X1 U5938 ( .A1(n4624), .A2(n4623), .ZN(n4452) );
  NOR2_X1 U5939 ( .A1(n9319), .A2(n9347), .ZN(n4453) );
  NOR2_X1 U5940 ( .A1(n8696), .A2(n8566), .ZN(n4454) );
  AND2_X1 U5941 ( .A1(n4893), .A2(n7828), .ZN(n4892) );
  AND2_X1 U5942 ( .A1(n8126), .A2(n8125), .ZN(n4455) );
  INV_X1 U5943 ( .A(n4866), .ZN(n4864) );
  AND2_X1 U5944 ( .A1(n6118), .A2(n6117), .ZN(n4456) );
  INV_X1 U5945 ( .A(n4958), .ZN(n4957) );
  NOR2_X1 U5946 ( .A1(n8749), .A2(n8591), .ZN(n4958) );
  INV_X1 U5947 ( .A(n7450), .ZN(n9843) );
  AND2_X1 U5948 ( .A1(n5647), .A2(n5637), .ZN(n4457) );
  INV_X1 U5949 ( .A(n9367), .ZN(n4710) );
  AND2_X1 U5950 ( .A1(n5709), .A2(n5585), .ZN(n5749) );
  INV_X1 U5951 ( .A(n4906), .ZN(n4905) );
  OR2_X1 U5952 ( .A1(n8342), .A2(n4907), .ZN(n4906) );
  OR2_X1 U5953 ( .A1(n7691), .A2(n4846), .ZN(n4458) );
  NOR2_X1 U5954 ( .A1(n8525), .A2(n8535), .ZN(n4459) );
  AND2_X1 U5955 ( .A1(n5596), .A2(n5672), .ZN(n9257) );
  OR3_X1 U5956 ( .A1(n5718), .A2(n5763), .A3(n5619), .ZN(n4460) );
  OR2_X1 U5957 ( .A1(n4445), .A2(n4797), .ZN(n4461) );
  XOR2_X1 U5958 ( .A(n6176), .B(n8525), .Z(n4462) );
  NAND2_X1 U5959 ( .A1(n8529), .A2(n4424), .ZN(n4463) );
  OR2_X1 U5960 ( .A1(n9392), .A2(n9238), .ZN(n9122) );
  INV_X1 U5961 ( .A(n9122), .ZN(n4836) );
  OR2_X1 U5962 ( .A1(n9415), .A2(n9306), .ZN(n4464) );
  AND2_X1 U5963 ( .A1(n7529), .A2(n7528), .ZN(n4465) );
  AND2_X1 U5964 ( .A1(n4689), .A2(n4691), .ZN(n4466) );
  AND2_X1 U5965 ( .A1(n9167), .A2(n9101), .ZN(n4467) );
  AND3_X1 U5966 ( .A1(n5893), .A2(n5892), .A3(n5891), .ZN(n9821) );
  AND2_X1 U5967 ( .A1(n8014), .A2(n8599), .ZN(n4468) );
  OR2_X1 U5968 ( .A1(n4934), .A2(n5109), .ZN(n4469) );
  AND2_X1 U5969 ( .A1(n4708), .A2(n9359), .ZN(n4470) );
  OR2_X1 U5970 ( .A1(n4831), .A2(n9128), .ZN(n4471) );
  AND2_X1 U5971 ( .A1(n8133), .A2(n8134), .ZN(n4472) );
  AND2_X1 U5972 ( .A1(n5935), .A2(n5922), .ZN(n4473) );
  AND2_X1 U5973 ( .A1(n4862), .A2(n7908), .ZN(n4474) );
  INV_X1 U5974 ( .A(n9392), .ZN(n9225) );
  NAND2_X1 U5975 ( .A1(n5154), .A2(n5153), .ZN(n9392) );
  AND2_X1 U5976 ( .A1(n4410), .A2(n8152), .ZN(n4475) );
  INV_X1 U5977 ( .A(n8136), .ZN(n4787) );
  OR2_X1 U5978 ( .A1(n7671), .A2(n7670), .ZN(n8136) );
  AND2_X1 U5979 ( .A1(n8187), .A2(n8186), .ZN(n4476) );
  INV_X1 U5980 ( .A(n4871), .ZN(n4597) );
  INV_X1 U5981 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5795) );
  AND2_X1 U5982 ( .A1(n8018), .A2(n4799), .ZN(n4477) );
  OR2_X1 U5983 ( .A1(n4422), .A2(n4662), .ZN(n4478) );
  AND2_X2 U5984 ( .A1(n6482), .A2(n4556), .ZN(n5862) );
  INV_X2 U5985 ( .A(n6041), .ZN(n6204) );
  AND2_X2 U5986 ( .A1(n6482), .A2(n6384), .ZN(n6119) );
  NAND2_X1 U5987 ( .A1(n5806), .A2(n5807), .ZN(n6075) );
  XNOR2_X1 U5988 ( .A(n7992), .B(n7952), .ZN(n4479) );
  AND2_X1 U5989 ( .A1(n6369), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4480) );
  NAND2_X1 U5990 ( .A1(n7909), .A2(n7908), .ZN(n8848) );
  AND2_X1 U5991 ( .A1(n9186), .A2(n9303), .ZN(n4481) );
  NAND2_X1 U5992 ( .A1(n6230), .A2(n6229), .ZN(n8652) );
  INV_X1 U5993 ( .A(n8652), .ZN(n4723) );
  AND2_X1 U5994 ( .A1(n4821), .A2(n4819), .ZN(n4482) );
  NAND2_X1 U5995 ( .A1(n5335), .A2(n4931), .ZN(n5293) );
  NAND2_X1 U5996 ( .A1(n5335), .A2(n5104), .ZN(n5321) );
  OR2_X1 U5997 ( .A1(n9244), .A2(n9255), .ZN(n4483) );
  NAND2_X1 U5998 ( .A1(n9280), .A2(n4411), .ZN(n4702) );
  INV_X1 U5999 ( .A(n4761), .ZN(n4760) );
  NAND2_X1 U6000 ( .A1(n5066), .A2(n5181), .ZN(n4761) );
  AND2_X1 U6001 ( .A1(n5267), .A2(n4883), .ZN(n5588) );
  NAND2_X1 U6002 ( .A1(n5335), .A2(n4434), .ZN(n4484) );
  AND2_X1 U6003 ( .A1(n5054), .A2(SI_18_), .ZN(n4485) );
  AND2_X1 U6004 ( .A1(n5068), .A2(SI_21_), .ZN(n4486) );
  OR2_X1 U6005 ( .A1(n8848), .A2(n8850), .ZN(n4487) );
  AND2_X1 U6006 ( .A1(n5141), .A2(n5078), .ZN(n4488) );
  AND2_X1 U6007 ( .A1(n7417), .A2(n7416), .ZN(n4489) );
  INV_X1 U6008 ( .A(n4614), .ZN(n4613) );
  AND2_X1 U6009 ( .A1(n7561), .A2(n7560), .ZN(n4490) );
  INV_X1 U6010 ( .A(n7373), .ZN(n4604) );
  NAND2_X1 U6011 ( .A1(n5714), .A2(n9214), .ZN(n6701) );
  INV_X1 U6012 ( .A(n6701), .ZN(n4562) );
  NAND2_X1 U6013 ( .A1(n5280), .A2(n5279), .ZN(n8898) );
  INV_X1 U6014 ( .A(n8898), .ZN(n4698) );
  NAND2_X1 U6015 ( .A1(n5269), .A2(n5268), .ZN(n8793) );
  INV_X1 U6016 ( .A(n8793), .ZN(n4697) );
  OR2_X1 U6017 ( .A1(n6642), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n4491) );
  OR2_X1 U6018 ( .A1(n6370), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4492) );
  AND2_X1 U6019 ( .A1(n8101), .A2(n8098), .ZN(n8046) );
  INV_X1 U6020 ( .A(n8046), .ZN(n4804) );
  INV_X1 U6021 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4647) );
  INV_X1 U6022 ( .A(n6814), .ZN(n6784) );
  INV_X1 U6023 ( .A(n5130), .ZN(n4769) );
  NAND2_X1 U6024 ( .A1(n4586), .A2(n4596), .ZN(n7845) );
  NAND2_X1 U6025 ( .A1(n7110), .A2(n8101), .ZN(n4493) );
  AND2_X1 U6026 ( .A1(n5568), .A2(SI_29_), .ZN(n4494) );
  AND2_X1 U6027 ( .A1(n7465), .A2(n7464), .ZN(n4495) );
  INV_X1 U6028 ( .A(n6791), .ZN(n4827) );
  OR2_X1 U6029 ( .A1(n7337), .A2(n7179), .ZN(n4496) );
  NAND2_X1 U6030 ( .A1(n6875), .A2(n6831), .ZN(n6993) );
  NAND2_X1 U6031 ( .A1(n5338), .A2(n5337), .ZN(n8885) );
  INV_X1 U6032 ( .A(n8885), .ZN(n4706) );
  OAI21_X1 U6033 ( .B1(n6992), .B2(n6993), .A(n6994), .ZN(n6996) );
  OR2_X1 U6034 ( .A1(n7262), .A2(n7137), .ZN(n7321) );
  INV_X1 U6035 ( .A(n7321), .ZN(n4703) );
  INV_X1 U6036 ( .A(n4716), .ZN(n9778) );
  NAND2_X1 U6037 ( .A1(n6892), .A2(n6760), .ZN(n4716) );
  XNOR2_X1 U6038 ( .A(n5207), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9214) );
  XNOR2_X1 U6039 ( .A(n5717), .B(P1_IR_REG_20__SCAN_IN), .ZN(n6700) );
  AOI211_X1 U6040 ( .C1(n8342), .C2(n8341), .A(n8340), .B(n8339), .ZN(n8351)
         );
  NAND4_X2 U6041 ( .A1(n4962), .A2(n4618), .A3(n4617), .A4(n4616), .ZN(n5864)
         );
  NOR2_X4 U6042 ( .A1(n5864), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5887) );
  NAND2_X4 U6043 ( .A1(n8765), .A2(n8767), .ZN(n6482) );
  XNOR2_X1 U6044 ( .A(n6202), .B(n6193), .ZN(n8311) );
  OR2_X1 U6045 ( .A1(n5881), .A2(n5880), .ZN(n5882) );
  NAND2_X1 U6046 ( .A1(n5941), .A2(n5940), .ZN(n6927) );
  NAND2_X2 U6047 ( .A1(n7121), .A2(n8102), .ZN(n7228) );
  AOI21_X2 U6048 ( .B1(n9729), .B2(n9728), .A(n7120), .ZN(n7121) );
  NOR2_X2 U6049 ( .A1(n5817), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5819) );
  NAND2_X1 U6050 ( .A1(n5357), .A2(n5007), .ZN(n4737) );
  AOI21_X1 U6051 ( .B1(n8598), .B2(n4468), .A(n4807), .ZN(n8545) );
  OAI21_X2 U6052 ( .B1(n5266), .B2(n5036), .A(n5035), .ZN(n5369) );
  NOR2_X2 U6053 ( .A1(n8437), .A2(n8436), .ZN(n8435) );
  NAND2_X1 U6054 ( .A1(n5418), .A2(n5417), .ZN(n4987) );
  NAND2_X1 U6055 ( .A1(n4997), .A2(n4996), .ZN(n5448) );
  OAI21_X1 U6056 ( .B1(n7023), .B2(n4805), .A(n4803), .ZN(n7113) );
  NAND2_X1 U6057 ( .A1(n8485), .A2(n4477), .ZN(n4795) );
  NAND2_X1 U6058 ( .A1(n5152), .A2(n5151), .ZN(n4782) );
  INV_X1 U6059 ( .A(n5777), .ZN(n4530) );
  NAND2_X1 U6060 ( .A1(n4677), .A2(n4729), .ZN(n4676) );
  NAND2_X1 U6061 ( .A1(n5522), .A2(n5521), .ZN(n5092) );
  NAND2_X1 U6062 ( .A1(n5082), .A2(n5081), .ZN(n5163) );
  INV_X1 U6063 ( .A(n4997), .ZN(n4661) );
  NAND2_X1 U6064 ( .A1(n5003), .A2(n5002), .ZN(n5358) );
  NAND2_X1 U6065 ( .A1(n4525), .A2(n4523), .ZN(n4522) );
  OAI21_X2 U6066 ( .B1(n8616), .B2(n4954), .A(n4952), .ZN(n8572) );
  NAND2_X2 U6067 ( .A1(n7455), .A2(n7454), .ZN(n7465) );
  AND2_X2 U6068 ( .A1(n4801), .A2(n4799), .ZN(n8467) );
  NAND2_X1 U6069 ( .A1(n4784), .A2(n4785), .ZN(n7776) );
  OAI21_X1 U6070 ( .B1(n4792), .B2(n4791), .A(n8128), .ZN(n4790) );
  NAND2_X1 U6071 ( .A1(n4728), .A2(n4731), .ZN(n5319) );
  INV_X1 U6072 ( .A(n4660), .ZN(n4659) );
  AOI21_X2 U6073 ( .B1(n8311), .B2(n8312), .A(n4515), .ZN(n8305) );
  NAND2_X2 U6074 ( .A1(n5921), .A2(n5920), .ZN(n6767) );
  NAND2_X1 U6075 ( .A1(n6927), .A2(n6926), .ZN(n4913) );
  OAI21_X1 U6076 ( .B1(n6270), .B2(P2_IR_REG_26__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U6077 ( .A1(n5874), .A2(n4885), .ZN(n5883) );
  NOR2_X1 U6078 ( .A1(n4522), .A2(n4519), .ZN(n4521) );
  NAND2_X1 U6079 ( .A1(n4521), .A2(n4520), .ZN(P1_U3240) );
  NAND2_X1 U6080 ( .A1(n5659), .A2(n4542), .ZN(n4541) );
  NAND3_X1 U6081 ( .A1(n5766), .A2(n4391), .A3(n4553), .ZN(n4550) );
  NAND3_X1 U6082 ( .A1(n4560), .A2(n6701), .A3(n5735), .ZN(n4559) );
  NOR2_X4 U6083 ( .A1(n5481), .A2(n4583), .ZN(n5335) );
  OAI21_X2 U6084 ( .B1(n7373), .B2(n4589), .A(n4587), .ZN(n8876) );
  NAND2_X1 U6085 ( .A1(n4591), .A2(n8878), .ZN(n4590) );
  NAND2_X1 U6086 ( .A1(n4602), .A2(n4601), .ZN(n7847) );
  NAND2_X1 U6087 ( .A1(n8821), .A2(n4607), .ZN(n4606) );
  NAND2_X1 U6088 ( .A1(n8821), .A2(n8822), .ZN(n4612) );
  NAND2_X1 U6089 ( .A1(n7948), .A2(n7947), .ZN(n4614) );
  AOI21_X2 U6090 ( .B1(n4615), .B2(n4863), .A(n4423), .ZN(n8936) );
  INV_X2 U6091 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4616) );
  INV_X2 U6092 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4617) );
  NAND2_X1 U6093 ( .A1(n4455), .A2(n4409), .ZN(n4620) );
  NAND3_X1 U6094 ( .A1(n4620), .A2(n4472), .A3(n4619), .ZN(n8140) );
  NAND3_X1 U6095 ( .A1(n8040), .A2(n4645), .A3(n8210), .ZN(n4644) );
  NAND2_X1 U6096 ( .A1(n4652), .A2(n8191), .ZN(n8195) );
  NAND3_X1 U6097 ( .A1(n4654), .A2(n4476), .A3(n4653), .ZN(n4652) );
  NAND3_X1 U6098 ( .A1(n8178), .A2(n8197), .A3(n4655), .ZN(n4654) );
  AOI21_X1 U6099 ( .B1(n5447), .B2(n4662), .A(n4422), .ZN(n4657) );
  INV_X1 U6100 ( .A(n5447), .ZN(n4658) );
  OAI21_X1 U6101 ( .B1(n4661), .B2(n4478), .A(n4659), .ZN(n5003) );
  OAI21_X1 U6102 ( .B1(n5447), .B2(n4422), .A(n5000), .ZN(n4660) );
  INV_X1 U6103 ( .A(n4987), .ZN(n4670) );
  OAI21_X1 U6104 ( .B1(n4987), .B2(n4666), .A(n4665), .ZN(n5479) );
  AOI21_X1 U6105 ( .B1(n4671), .B2(n5461), .A(n4421), .ZN(n4665) );
  INV_X1 U6106 ( .A(n5461), .ZN(n4666) );
  OAI21_X1 U6107 ( .B1(n4670), .B2(n4669), .A(n4667), .ZN(n4993) );
  INV_X1 U6108 ( .A(n4668), .ZN(n4667) );
  OAI21_X1 U6109 ( .B1(n5461), .B2(n4421), .A(n5478), .ZN(n4668) );
  NAND2_X1 U6110 ( .A1(n4672), .A2(n4467), .ZN(n9105) );
  INV_X1 U6111 ( .A(n5358), .ZN(n4677) );
  NAND3_X1 U6112 ( .A1(n4676), .A2(n4674), .A3(n5017), .ZN(n5306) );
  NAND3_X1 U6113 ( .A1(n4676), .A2(n4675), .A3(n4674), .ZN(n4681) );
  NAND2_X1 U6114 ( .A1(n4678), .A2(n4729), .ZN(n5317) );
  NAND2_X1 U6115 ( .A1(n5358), .A2(n4731), .ZN(n4678) );
  INV_X1 U6116 ( .A(n5017), .ZN(n4679) );
  INV_X1 U6117 ( .A(n4731), .ZN(n4680) );
  NAND2_X1 U6118 ( .A1(n4920), .A2(n4466), .ZN(n4683) );
  NAND2_X1 U6119 ( .A1(n4683), .A2(n4682), .ZN(n9090) );
  AND2_X2 U6120 ( .A1(n5423), .A2(n4692), .ZN(n9649) );
  AND2_X1 U6121 ( .A1(n5425), .A2(n5424), .ZN(n4692) );
  NAND2_X1 U6122 ( .A1(n5277), .A2(n5108), .ZN(n5767) );
  NAND3_X1 U6123 ( .A1(n5277), .A2(n4694), .A3(n9923), .ZN(n5110) );
  INV_X1 U6124 ( .A(n4702), .ZN(n9239) );
  NAND2_X1 U6125 ( .A1(n4419), .A2(n4703), .ZN(n7647) );
  AND2_X1 U6126 ( .A1(n9176), .A2(n4707), .ZN(n9148) );
  NAND2_X1 U6127 ( .A1(n9176), .A2(n4708), .ZN(n9137) );
  NAND2_X1 U6128 ( .A1(n9176), .A2(n9165), .ZN(n9159) );
  NAND4_X1 U6129 ( .A1(n5786), .A2(n5792), .A3(n4965), .A4(n5887), .ZN(n6270)
         );
  NOR2_X2 U6130 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  NOR2_X2 U6131 ( .A1(n5785), .A2(n5784), .ZN(n5786) );
  NAND2_X1 U6132 ( .A1(n7612), .A2(n4475), .ZN(n8611) );
  INV_X1 U6133 ( .A(n9731), .ZN(n4718) );
  NAND3_X1 U6134 ( .A1(n4721), .A2(n4719), .A3(n4718), .ZN(n7467) );
  INV_X1 U6135 ( .A(n4727), .ZN(n8488) );
  AOI21_X2 U6136 ( .B1(n4731), .B2(n4734), .A(n4730), .ZN(n4729) );
  INV_X1 U6137 ( .A(n5713), .ZN(n4738) );
  NAND2_X1 U6138 ( .A1(n5708), .A2(n4742), .ZN(n4739) );
  NAND3_X1 U6139 ( .A1(n4739), .A2(n4740), .A3(n4738), .ZN(n4744) );
  NAND2_X1 U6140 ( .A1(n5047), .A2(n4750), .ZN(n4747) );
  NAND2_X1 U6141 ( .A1(n4747), .A2(n4748), .ZN(n5203) );
  NAND2_X1 U6142 ( .A1(n5047), .A2(n5046), .ZN(n5233) );
  NAND2_X1 U6143 ( .A1(n5062), .A2(n4756), .ZN(n4755) );
  NAND2_X1 U6144 ( .A1(n4755), .A2(n4758), .ZN(n5172) );
  NAND2_X1 U6145 ( .A1(n5098), .A2(n5097), .ZN(n5131) );
  NAND2_X1 U6146 ( .A1(n5306), .A2(n4774), .ZN(n4770) );
  NAND2_X1 U6147 ( .A1(n4770), .A2(n4771), .ZN(n5266) );
  NAND2_X1 U6148 ( .A1(n4782), .A2(n5078), .ZN(n5142) );
  NAND2_X1 U6149 ( .A1(n4782), .A2(n4488), .ZN(n5082) );
  NAND2_X1 U6150 ( .A1(n9767), .A2(n8081), .ZN(n6905) );
  NAND2_X1 U6151 ( .A1(n4783), .A2(n4437), .ZN(n9767) );
  AND2_X1 U6152 ( .A1(n8077), .A2(n8081), .ZN(n4783) );
  NAND2_X1 U6153 ( .A1(n8073), .A2(n7007), .ZN(n8077) );
  NAND2_X1 U6154 ( .A1(n7608), .A2(n8136), .ZN(n4784) );
  NAND2_X1 U6155 ( .A1(n4795), .A2(n4796), .ZN(n8437) );
  XNOR2_X2 U6156 ( .A(n4802), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5823) );
  XNOR2_X2 U6157 ( .A(n5820), .B(n5818), .ZN(n8762) );
  AOI21_X1 U6158 ( .B1(n4806), .B2(n4804), .A(n4412), .ZN(n4803) );
  NAND2_X1 U6159 ( .A1(n9109), .A2(n4408), .ZN(n4816) );
  NAND2_X1 U6160 ( .A1(n7292), .A2(n7293), .ZN(n5427) );
  NAND2_X1 U6161 ( .A1(n9199), .A2(n4830), .ZN(n4829) );
  NOR2_X1 U6162 ( .A1(n9199), .A2(n9125), .ZN(n9182) );
  NAND2_X1 U6163 ( .A1(n4829), .A2(n4471), .ZN(n9153) );
  NAND2_X1 U6164 ( .A1(n9251), .A2(n4838), .ZN(n4837) );
  INV_X1 U6165 ( .A(n4844), .ZN(n9250) );
  AND2_X2 U6166 ( .A1(n9470), .A2(n5123), .ZN(n5390) );
  INV_X1 U6167 ( .A(n7692), .ZN(n4848) );
  AND3_X2 U6168 ( .A1(n5335), .A2(n4930), .A3(n4931), .ZN(n5277) );
  OAI21_X2 U6169 ( .B1(n8809), .B2(n7863), .A(n4859), .ZN(n8926) );
  OR2_X1 U6170 ( .A1(n8807), .A2(n8806), .ZN(n4859) );
  NAND2_X1 U6171 ( .A1(n8876), .A2(n7857), .ZN(n8809) );
  NAND2_X1 U6172 ( .A1(n7909), .A2(n4474), .ZN(n4860) );
  NAND2_X1 U6173 ( .A1(n4860), .A2(n4861), .ZN(n8934) );
  NAND2_X1 U6174 ( .A1(n6985), .A2(n5714), .ZN(n6783) );
  NAND3_X1 U6175 ( .A1(n6985), .A2(n5714), .A3(n5762), .ZN(n6986) );
  NAND2_X1 U6176 ( .A1(n8829), .A2(n4880), .ZN(n8904) );
  NAND2_X1 U6177 ( .A1(n6874), .A2(n6876), .ZN(n6875) );
  NAND2_X1 U6178 ( .A1(n5267), .A2(n4882), .ZN(n5752) );
  CLKBUF_X1 U6179 ( .A(n4885), .Z(n4884) );
  NAND2_X1 U6180 ( .A1(n4884), .A2(n6745), .ZN(n6672) );
  XNOR2_X1 U6181 ( .A(n4884), .B(n6745), .ZN(n6750) );
  OR2_X1 U6182 ( .A1(n5852), .A2(n5851), .ZN(n4886) );
  NAND2_X1 U6183 ( .A1(n8305), .A2(n4909), .ZN(n4908) );
  NAND2_X1 U6184 ( .A1(n4913), .A2(n4911), .ZN(n7093) );
  NAND2_X1 U6185 ( .A1(n7405), .A2(n4916), .ZN(n4915) );
  NAND2_X1 U6186 ( .A1(n6767), .A2(n4473), .ZN(n5941) );
  NAND2_X1 U6187 ( .A1(n4923), .A2(n4921), .ZN(n4920) );
  NAND2_X1 U6188 ( .A1(n7259), .A2(n4418), .ZN(n7278) );
  NAND3_X1 U6189 ( .A1(n4695), .A2(n4937), .A3(n4936), .ZN(n4935) );
  NAND2_X1 U6190 ( .A1(n8546), .A2(n4941), .ZN(n4938) );
  XNOR2_X2 U6191 ( .A(n4949), .B(n4641), .ZN(n8647) );
  NAND2_X2 U6192 ( .A1(n7561), .A2(n4959), .ZN(n7605) );
  NAND2_X2 U6193 ( .A1(n7465), .A2(n4960), .ZN(n7561) );
  INV_X1 U6194 ( .A(n7114), .ZN(n7116) );
  NAND3_X1 U6195 ( .A1(n5887), .A2(n5786), .A3(n5792), .ZN(n6268) );
  AND2_X1 U6196 ( .A1(n5830), .A2(n5840), .ZN(n6739) );
  OR2_X1 U6197 ( .A1(n5829), .A2(n5828), .ZN(n5830) );
  AND2_X4 U6198 ( .A1(n8224), .A2(n8038), .ZN(n5846) );
  NAND2_X1 U6199 ( .A1(n8261), .A2(n9774), .ZN(n8265) );
  OR2_X1 U6200 ( .A1(n6815), .A2(n7955), .ZN(n6816) );
  NAND2_X1 U6201 ( .A1(n6739), .A2(n6738), .ZN(n6737) );
  AOI211_X2 U6202 ( .C1(n8644), .C2(n9761), .A(n8267), .B(n8266), .ZN(n8268)
         );
  OAI21_X1 U6203 ( .B1(n4414), .B2(n9147), .A(n9146), .ZN(n9371) );
  OAI22_X1 U6204 ( .A1(n6818), .A2(n7848), .B1(n6832), .B2(n9645), .ZN(n6819)
         );
  NAND2_X1 U6205 ( .A1(n7605), .A2(n7604), .ZN(n7673) );
  NAND2_X2 U6206 ( .A1(n7194), .A2(n7193), .ZN(n7373) );
  OAI22_X1 U6207 ( .A1(n8242), .A2(n8241), .B1(n8359), .B2(n8755), .ZN(n8614)
         );
  INV_X2 U6208 ( .A(n5823), .ZN(n8240) );
  NOR2_X2 U6209 ( .A1(n8932), .A2(n8936), .ZN(n8814) );
  AND2_X4 U6210 ( .A1(n8240), .A2(n8762), .ZN(n5857) );
  NOR2_X1 U6211 ( .A1(n7747), .A2(n7746), .ZN(n4966) );
  OR2_X1 U6212 ( .A1(n6785), .A2(n8986), .ZN(n4967) );
  AND2_X1 U6213 ( .A1(n7936), .A2(n7935), .ZN(n4968) );
  AND4_X1 U6214 ( .A1(n5204), .A2(n5755), .A3(n5754), .A4(n5753), .ZN(n4969)
         );
  AND3_X1 U6215 ( .A1(n6287), .A2(n6289), .A3(n7594), .ZN(n4970) );
  AND2_X1 U6216 ( .A1(n8229), .A2(n8228), .ZN(n4971) );
  INV_X1 U6217 ( .A(n5862), .ZN(n6041) );
  AND4_X1 U6218 ( .A1(n5205), .A2(n5107), .A3(n5106), .A4(n5757), .ZN(n4972)
         );
  OR2_X1 U6219 ( .A1(n8442), .A2(n8460), .ZN(n4973) );
  INV_X1 U6220 ( .A(n8102), .ZN(n7111) );
  INV_X1 U6221 ( .A(n7521), .ZN(n6832) );
  INV_X1 U6222 ( .A(n6195), .ZN(n6194) );
  INV_X1 U6223 ( .A(n6181), .ZN(n6180) );
  INV_X1 U6224 ( .A(n8018), .ZN(n8201) );
  AND2_X1 U6225 ( .A1(n7862), .A2(n7861), .ZN(n8806) );
  INV_X1 U6226 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5439) );
  OR2_X1 U6227 ( .A1(n6175), .A2(n6174), .ZN(n6190) );
  INV_X1 U6228 ( .A(n6203), .ZN(n6193) );
  NAND2_X1 U6229 ( .A1(n6136), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6144) );
  OR2_X1 U6230 ( .A1(n6208), .A2(n9935), .ZN(n6219) );
  OR2_X1 U6231 ( .A1(n6164), .A2(n8328), .ZN(n6181) );
  AND2_X1 U6232 ( .A1(n8398), .A2(n8397), .ZN(n8395) );
  OR2_X1 U6233 ( .A1(n6144), .A2(n8297), .ZN(n6164) );
  AND2_X1 U6234 ( .A1(n8775), .A2(n8776), .ZN(n7987) );
  INV_X1 U6235 ( .A(n8832), .ZN(n7881) );
  NAND2_X1 U6236 ( .A1(n6786), .A2(n4967), .ZN(n6787) );
  NOR2_X1 U6237 ( .A1(n5197), .A2(n8823), .ZN(n5186) );
  OR2_X1 U6238 ( .A1(n5399), .A2(n7159), .ZN(n5393) );
  OR2_X1 U6239 ( .A1(n5300), .A2(n5281), .ZN(n5378) );
  OAI21_X1 U6240 ( .B1(n9208), .B2(n9124), .A(n9123), .ZN(n9199) );
  INV_X1 U6241 ( .A(n9603), .ZN(n7137) );
  NAND2_X1 U6242 ( .A1(n5629), .A2(n5600), .ZN(n7267) );
  INV_X1 U6243 ( .A(n5588), .ZN(n5220) );
  NAND2_X1 U6244 ( .A1(n6014), .A2(n6013), .ZN(n6033) );
  OR2_X1 U6245 ( .A1(n5963), .A2(n5962), .ZN(n5983) );
  OR2_X1 U6246 ( .A1(n7627), .A2(n9743), .ZN(n8333) );
  OR2_X1 U6247 ( .A1(n6309), .A2(n9788), .ZN(n6301) );
  OR2_X1 U6248 ( .A1(n8443), .A2(n6295), .ZN(n6250) );
  NAND2_X1 U6249 ( .A1(n8256), .A2(n8199), .ZN(n8436) );
  INV_X1 U6250 ( .A(n8674), .ZN(n8525) );
  INV_X1 U6251 ( .A(n8245), .ZN(n8571) );
  AND2_X1 U6252 ( .A1(n8156), .A2(n8164), .ZN(n8599) );
  OR2_X1 U6253 ( .A1(n5983), .A2(n5982), .ZN(n6017) );
  OR2_X1 U6254 ( .A1(n6646), .A2(n6645), .ZN(n6803) );
  INV_X1 U6255 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5977) );
  AND2_X1 U6256 ( .A1(n7367), .A2(n7368), .ZN(n7372) );
  AND2_X1 U6257 ( .A1(n7965), .A2(n7962), .ZN(n8866) );
  NOR2_X1 U6258 ( .A1(n8934), .A2(n8933), .ZN(n8932) );
  NOR2_X1 U6259 ( .A1(n5155), .A2(n8871), .ZN(n5166) );
  OR2_X1 U6260 ( .A1(n5540), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5459) );
  AND4_X2 U6261 ( .A1(n5394), .A2(n5393), .A3(n5392), .A4(n5391), .ZN(n6818)
         );
  NAND2_X1 U6262 ( .A1(n9415), .A2(n9306), .ZN(n9089) );
  AND2_X1 U6263 ( .A1(n9110), .A2(n9111), .ZN(n9344) );
  AND2_X1 U6264 ( .A1(n5660), .A2(n9107), .ZN(n7755) );
  INV_X1 U6265 ( .A(n8975), .ZN(n9493) );
  OR2_X1 U6266 ( .A1(n6981), .A2(n6854), .ZN(n9492) );
  AND2_X1 U6267 ( .A1(n7362), .A2(n6978), .ZN(n6985) );
  AND2_X1 U6268 ( .A1(n6980), .A2(n6979), .ZN(n9488) );
  AND2_X1 U6269 ( .A1(n5046), .A2(n5045), .ZN(n5250) );
  AND2_X1 U6270 ( .A1(n5012), .A2(n5011), .ZN(n5334) );
  NAND2_X1 U6271 ( .A1(n4991), .A2(SI_4_), .ZN(n4992) );
  INV_X1 U6272 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5449) );
  AND2_X1 U6273 ( .A1(n6250), .A2(n6249), .ZN(n8249) );
  INV_X1 U6274 ( .A(n9686), .ZN(n9715) );
  NOR2_X1 U6275 ( .A1(n8646), .A2(n4392), .ZN(n8266) );
  AND2_X1 U6276 ( .A1(n9734), .A2(n9845), .ZN(n9761) );
  OR2_X1 U6277 ( .A1(n9788), .A2(n6647), .ZN(n9750) );
  INV_X1 U6278 ( .A(n9838), .ZN(n9845) );
  INV_X1 U6279 ( .A(n9848), .ZN(n9859) );
  AND2_X1 U6280 ( .A1(n6276), .A2(n6275), .ZN(n9787) );
  AND2_X1 U6281 ( .A1(n6843), .A2(n6854), .ZN(n8962) );
  AND2_X1 U6282 ( .A1(n6843), .A2(n4391), .ZN(n8921) );
  INV_X1 U6283 ( .A(n8969), .ZN(n8944) );
  AND4_X1 U6284 ( .A1(n5180), .A2(n5179), .A3(n5178), .A4(n5177), .ZN(n9255)
         );
  INV_X1 U6285 ( .A(n9102), .ZN(n9167) );
  AND2_X1 U6286 ( .A1(n5597), .A2(n9117), .ZN(n9273) );
  AND2_X1 U6287 ( .A1(n5598), .A2(n9299), .ZN(n9315) );
  INV_X1 U6288 ( .A(n9491), .ZN(n9303) );
  INV_X1 U6289 ( .A(n9645), .ZN(n7162) );
  OR2_X1 U6290 ( .A1(n7065), .A2(n6796), .ZN(n9605) );
  OR2_X1 U6291 ( .A1(n7206), .A2(n6985), .ZN(n9666) );
  INV_X1 U6292 ( .A(n9528), .ZN(n9434) );
  INV_X1 U6293 ( .A(n5762), .ZN(n5619) );
  XNOR2_X1 U6294 ( .A(n4999), .B(n4998), .ZN(n5447) );
  XNOR2_X1 U6295 ( .A(n4988), .B(SI_3_), .ZN(n5461) );
  INV_X1 U6296 ( .A(n8336), .ZN(n8349) );
  INV_X1 U6297 ( .A(n7594), .ZN(n8340) );
  AND2_X1 U6298 ( .A1(n6300), .A2(n6299), .ZN(n8438) );
  AND2_X1 U6299 ( .A1(n6427), .A2(n6426), .ZN(n8419) );
  INV_X1 U6300 ( .A(n8477), .ZN(n8729) );
  INV_X1 U6301 ( .A(n7798), .ZN(n8755) );
  INV_X1 U6302 ( .A(n9861), .ZN(n9860) );
  INV_X1 U6303 ( .A(n9789), .ZN(n9792) );
  INV_X1 U6304 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6390) );
  INV_X1 U6305 ( .A(n9382), .ZN(n9198) );
  AND2_X1 U6306 ( .A1(n6842), .A2(n6841), .ZN(n8965) );
  INV_X1 U6307 ( .A(n8967), .ZN(n8954) );
  INV_X1 U6308 ( .A(n9255), .ZN(n9228) );
  OR2_X1 U6309 ( .A1(P1_U3083), .A2(n6350), .ZN(n9586) );
  AND2_X1 U6310 ( .A1(n7723), .A2(n7722), .ZN(n9534) );
  OR2_X1 U6311 ( .A1(n6780), .A2(n6727), .ZN(n9680) );
  AND2_X1 U6312 ( .A1(n9534), .A2(n9533), .ZN(n9549) );
  OR2_X1 U6313 ( .A1(n6780), .A2(n6716), .ZN(n9674) );
  CLKBUF_X1 U6314 ( .A(n9643), .Z(n9633) );
  AND2_X1 U6315 ( .A1(n6838), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6795) );
  INV_X1 U6316 ( .A(n5123), .ZN(n8005) );
  INV_X1 U6317 ( .A(n6700), .ZN(n7362) );
  INV_X1 U6318 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6392) );
  NAND2_X4 U6319 ( .A1(n4977), .A2(n4976), .ZN(n6384) );
  NAND2_X1 U6320 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4979) );
  AND2_X1 U6321 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4978) );
  NAND2_X1 U6322 ( .A1(n6384), .A2(n4978), .ZN(n5406) );
  OAI21_X1 U6323 ( .B1(n6384), .B2(n4979), .A(n5406), .ZN(n4981) );
  INV_X1 U6324 ( .A(SI_1_), .ZN(n4980) );
  XNOR2_X1 U6325 ( .A(n4981), .B(n4980), .ZN(n5396) );
  MUX2_X1 U6326 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6384), .Z(n5395) );
  NAND2_X1 U6327 ( .A1(n5396), .A2(n5395), .ZN(n4983) );
  NAND2_X1 U6328 ( .A1(n4981), .A2(SI_1_), .ZN(n4982) );
  NAND2_X1 U6329 ( .A1(n4983), .A2(n4982), .ZN(n5418) );
  MUX2_X1 U6330 ( .A(n6381), .B(n6396), .S(n6384), .Z(n4984) );
  XNOR2_X1 U6331 ( .A(n4984), .B(SI_2_), .ZN(n5417) );
  INV_X1 U6332 ( .A(n4984), .ZN(n4985) );
  NAND2_X1 U6333 ( .A1(n4985), .A2(SI_2_), .ZN(n4986) );
  MUX2_X1 U6334 ( .A(n6383), .B(n6388), .S(n6384), .Z(n4988) );
  INV_X1 U6335 ( .A(n4988), .ZN(n4989) );
  MUX2_X1 U6336 ( .A(n6387), .B(n6394), .S(n6384), .Z(n4990) );
  XNOR2_X1 U6337 ( .A(n4990), .B(SI_4_), .ZN(n5478) );
  INV_X1 U6338 ( .A(n4990), .ZN(n4991) );
  NAND2_X1 U6339 ( .A1(n4993), .A2(n4992), .ZN(n5434) );
  MUX2_X1 U6340 ( .A(n6390), .B(n6392), .S(n6384), .Z(n4994) );
  NAND2_X1 U6341 ( .A1(n5434), .A2(n5433), .ZN(n4997) );
  INV_X1 U6342 ( .A(n4994), .ZN(n4995) );
  NAND2_X1 U6343 ( .A1(n4995), .A2(SI_5_), .ZN(n4996) );
  MUX2_X1 U6344 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6380), .Z(n4999) );
  INV_X1 U6345 ( .A(SI_6_), .ZN(n4998) );
  MUX2_X1 U6346 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6380), .Z(n5001) );
  NAND2_X1 U6347 ( .A1(n5001), .A2(SI_7_), .ZN(n5002) );
  INV_X1 U6348 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6411) );
  INV_X1 U6349 ( .A(SI_8_), .ZN(n9950) );
  INV_X1 U6350 ( .A(n5004), .ZN(n5005) );
  NAND2_X1 U6351 ( .A1(n5005), .A2(SI_8_), .ZN(n5006) );
  INV_X1 U6352 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6415) );
  MUX2_X1 U6353 ( .A(n6415), .B(n9976), .S(n6380), .Z(n5009) );
  INV_X1 U6354 ( .A(SI_9_), .ZN(n5008) );
  INV_X1 U6355 ( .A(n5009), .ZN(n5010) );
  NAND2_X1 U6356 ( .A1(n5010), .A2(SI_9_), .ZN(n5011) );
  INV_X1 U6357 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6419) );
  INV_X1 U6358 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6421) );
  MUX2_X1 U6359 ( .A(n6419), .B(n6421), .S(n6380), .Z(n5014) );
  INV_X1 U6360 ( .A(SI_10_), .ZN(n5013) );
  NAND2_X1 U6361 ( .A1(n5014), .A2(n5013), .ZN(n5017) );
  INV_X1 U6362 ( .A(n5014), .ZN(n5015) );
  NAND2_X1 U6363 ( .A1(n5015), .A2(SI_10_), .ZN(n5016) );
  INV_X1 U6364 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6429) );
  INV_X1 U6365 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6431) );
  MUX2_X1 U6366 ( .A(n6429), .B(n6431), .S(n6380), .Z(n5018) );
  INV_X1 U6367 ( .A(n5018), .ZN(n5019) );
  NAND2_X1 U6368 ( .A1(n5019), .A2(SI_11_), .ZN(n5020) );
  INV_X1 U6369 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10181) );
  INV_X1 U6370 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9953) );
  MUX2_X1 U6371 ( .A(n10181), .B(n9953), .S(n6380), .Z(n5023) );
  INV_X1 U6372 ( .A(SI_12_), .ZN(n5022) );
  NAND2_X1 U6373 ( .A1(n5023), .A2(n5022), .ZN(n5026) );
  INV_X1 U6374 ( .A(n5023), .ZN(n5024) );
  NAND2_X1 U6375 ( .A1(n5024), .A2(SI_12_), .ZN(n5025) );
  NAND2_X1 U6376 ( .A1(n5026), .A2(n5025), .ZN(n5291) );
  INV_X1 U6377 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6661) );
  INV_X1 U6378 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5027) );
  MUX2_X1 U6379 ( .A(n6661), .B(n5027), .S(n6380), .Z(n5029) );
  INV_X1 U6380 ( .A(SI_13_), .ZN(n5028) );
  NAND2_X1 U6381 ( .A1(n5029), .A2(n5028), .ZN(n5032) );
  INV_X1 U6382 ( .A(n5029), .ZN(n5030) );
  NAND2_X1 U6383 ( .A1(n5030), .A2(SI_13_), .ZN(n5031) );
  MUX2_X1 U6384 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6380), .Z(n5034) );
  INV_X1 U6385 ( .A(SI_14_), .ZN(n5033) );
  XNOR2_X1 U6386 ( .A(n5034), .B(n5033), .ZN(n5265) );
  INV_X1 U6387 ( .A(n5265), .ZN(n5036) );
  NAND2_X1 U6388 ( .A1(n5034), .A2(SI_14_), .ZN(n5035) );
  INV_X1 U6389 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5037) );
  INV_X1 U6390 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6777) );
  MUX2_X1 U6391 ( .A(n5037), .B(n6777), .S(n6380), .Z(n5039) );
  INV_X1 U6392 ( .A(SI_15_), .ZN(n5038) );
  NAND2_X1 U6393 ( .A1(n5039), .A2(n5038), .ZN(n5042) );
  INV_X1 U6394 ( .A(n5039), .ZN(n5040) );
  NAND2_X1 U6395 ( .A1(n5040), .A2(SI_15_), .ZN(n5041) );
  NAND2_X1 U6396 ( .A1(n5042), .A2(n5041), .ZN(n5368) );
  OAI21_X2 U6397 ( .B1(n5369), .B2(n5368), .A(n5042), .ZN(n5251) );
  INV_X1 U6398 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6934) );
  INV_X1 U6399 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6933) );
  MUX2_X1 U6400 ( .A(n6934), .B(n6933), .S(n6380), .Z(n5043) );
  INV_X1 U6401 ( .A(SI_16_), .ZN(n10127) );
  NAND2_X1 U6402 ( .A1(n5043), .A2(n10127), .ZN(n5046) );
  INV_X1 U6403 ( .A(n5043), .ZN(n5044) );
  NAND2_X1 U6404 ( .A1(n5044), .A2(SI_16_), .ZN(n5045) );
  INV_X1 U6405 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6963) );
  INV_X1 U6406 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5048) );
  MUX2_X1 U6407 ( .A(n6963), .B(n5048), .S(n6380), .Z(n5049) );
  XNOR2_X1 U6408 ( .A(n5049), .B(SI_17_), .ZN(n5232) );
  INV_X1 U6409 ( .A(n5232), .ZN(n5052) );
  INV_X1 U6410 ( .A(n5049), .ZN(n5050) );
  NAND2_X1 U6411 ( .A1(n5050), .A2(SI_17_), .ZN(n5051) );
  MUX2_X1 U6412 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6380), .Z(n5054) );
  XNOR2_X1 U6413 ( .A(n5054), .B(SI_18_), .ZN(n5218) );
  INV_X1 U6414 ( .A(n5218), .ZN(n5053) );
  INV_X1 U6415 ( .A(n5203), .ZN(n5060) );
  INV_X1 U6416 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7187) );
  INV_X1 U6417 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7189) );
  MUX2_X1 U6418 ( .A(n7187), .B(n7189), .S(n6380), .Z(n5056) );
  INV_X1 U6419 ( .A(SI_19_), .ZN(n5055) );
  NAND2_X1 U6420 ( .A1(n5056), .A2(n5055), .ZN(n5061) );
  INV_X1 U6421 ( .A(n5056), .ZN(n5057) );
  NAND2_X1 U6422 ( .A1(n5057), .A2(SI_19_), .ZN(n5058) );
  NAND2_X1 U6423 ( .A1(n5061), .A2(n5058), .ZN(n5202) );
  INV_X1 U6424 ( .A(n5202), .ZN(n5059) );
  NAND2_X1 U6425 ( .A1(n5060), .A2(n5059), .ZN(n5062) );
  INV_X1 U6426 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7360) );
  INV_X1 U6427 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7363) );
  MUX2_X1 U6428 ( .A(n7360), .B(n7363), .S(n6380), .Z(n5063) );
  INV_X1 U6429 ( .A(SI_20_), .ZN(n9997) );
  NAND2_X1 U6430 ( .A1(n5063), .A2(n9997), .ZN(n5066) );
  INV_X1 U6431 ( .A(n5063), .ZN(n5064) );
  NAND2_X1 U6432 ( .A1(n5064), .A2(SI_20_), .ZN(n5065) );
  AND2_X1 U6433 ( .A1(n5066), .A2(n5065), .ZN(n5192) );
  INV_X1 U6434 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7385) );
  INV_X1 U6435 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n5183) );
  MUX2_X1 U6436 ( .A(n7385), .B(n5183), .S(n6384), .Z(n5067) );
  XNOR2_X1 U6437 ( .A(n5067), .B(SI_21_), .ZN(n5181) );
  INV_X1 U6438 ( .A(n5067), .ZN(n5068) );
  INV_X1 U6439 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7510) );
  INV_X1 U6440 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8008) );
  MUX2_X1 U6441 ( .A(n7510), .B(n8008), .S(n6380), .Z(n5070) );
  INV_X1 U6442 ( .A(SI_22_), .ZN(n5069) );
  NAND2_X1 U6443 ( .A1(n5070), .A2(n5069), .ZN(n5073) );
  INV_X1 U6444 ( .A(n5070), .ZN(n5071) );
  NAND2_X1 U6445 ( .A1(n5071), .A2(SI_22_), .ZN(n5072) );
  NAND2_X1 U6446 ( .A1(n5073), .A2(n5072), .ZN(n5171) );
  INV_X1 U6447 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5074) );
  INV_X1 U6448 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7545) );
  MUX2_X1 U6449 ( .A(n5074), .B(n7545), .S(n6384), .Z(n5075) );
  INV_X1 U6450 ( .A(SI_23_), .ZN(n9946) );
  NAND2_X1 U6451 ( .A1(n5075), .A2(n9946), .ZN(n5078) );
  INV_X1 U6452 ( .A(n5075), .ZN(n5076) );
  NAND2_X1 U6453 ( .A1(n5076), .A2(SI_23_), .ZN(n5077) );
  AND2_X1 U6454 ( .A1(n5078), .A2(n5077), .ZN(n5151) );
  INV_X1 U6455 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9911) );
  INV_X1 U6456 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7690) );
  MUX2_X1 U6457 ( .A(n9911), .B(n7690), .S(n6380), .Z(n5079) );
  XNOR2_X1 U6458 ( .A(n5079), .B(SI_24_), .ZN(n5141) );
  INV_X1 U6459 ( .A(n5079), .ZN(n5080) );
  NAND2_X1 U6460 ( .A1(n5080), .A2(SI_24_), .ZN(n5081) );
  INV_X1 U6461 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7743) );
  INV_X1 U6462 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7740) );
  MUX2_X1 U6463 ( .A(n7743), .B(n7740), .S(n6380), .Z(n5083) );
  INV_X1 U6464 ( .A(SI_25_), .ZN(n10196) );
  NAND2_X1 U6465 ( .A1(n5083), .A2(n10196), .ZN(n5086) );
  INV_X1 U6466 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6467 ( .A1(n5084), .A2(SI_25_), .ZN(n5085) );
  NAND2_X1 U6468 ( .A1(n5086), .A2(n5085), .ZN(n5162) );
  INV_X1 U6469 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7820) );
  INV_X1 U6470 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7827) );
  MUX2_X1 U6471 ( .A(n7820), .B(n7827), .S(n6384), .Z(n5088) );
  INV_X1 U6472 ( .A(SI_26_), .ZN(n5087) );
  NAND2_X1 U6473 ( .A1(n5088), .A2(n5087), .ZN(n5091) );
  INV_X1 U6474 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6475 ( .A1(n5089), .A2(SI_26_), .ZN(n5090) );
  AND2_X1 U6476 ( .A1(n5091), .A2(n5090), .ZN(n5521) );
  INV_X1 U6477 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8770) );
  INV_X1 U6478 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7824) );
  MUX2_X1 U6479 ( .A(n8770), .B(n7824), .S(n6380), .Z(n5094) );
  INV_X1 U6480 ( .A(SI_27_), .ZN(n5093) );
  NAND2_X1 U6481 ( .A1(n5094), .A2(n5093), .ZN(n5097) );
  INV_X1 U6482 ( .A(n5094), .ZN(n5095) );
  NAND2_X1 U6483 ( .A1(n5095), .A2(SI_27_), .ZN(n5096) );
  AND2_X1 U6484 ( .A1(n5097), .A2(n5096), .ZN(n5533) );
  INV_X1 U6485 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8763) );
  INV_X1 U6486 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9478) );
  MUX2_X1 U6487 ( .A(n8763), .B(n9478), .S(n6384), .Z(n5100) );
  XNOR2_X1 U6488 ( .A(n5100), .B(SI_28_), .ZN(n5130) );
  INV_X1 U6489 ( .A(SI_28_), .ZN(n5099) );
  NAND2_X1 U6490 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  INV_X1 U6491 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8761) );
  INV_X1 U6492 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9469) );
  MUX2_X1 U6493 ( .A(n8761), .B(n9469), .S(n6380), .Z(n5567) );
  XNOR2_X1 U6494 ( .A(n5567), .B(SI_29_), .ZN(n5102) );
  NOR2_X1 U6495 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5205) );
  NOR2_X1 U6496 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5107) );
  NOR2_X1 U6497 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5106) );
  INV_X1 U6498 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5757) );
  INV_X1 U6499 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5204) );
  INV_X1 U6500 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5754) );
  INV_X1 U6501 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5773) );
  INV_X1 U6502 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9938) );
  INV_X1 U6503 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5769) );
  NAND3_X1 U6504 ( .A1(n5773), .A2(n9938), .A3(n5769), .ZN(n5109) );
  INV_X1 U6505 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9923) );
  INV_X1 U6506 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5114) );
  XNOR2_X2 U6507 ( .A(n5112), .B(n9923), .ZN(n5766) );
  NOR2_X1 U6508 ( .A1(n5419), .A2(n9469), .ZN(n5113) );
  INV_X1 U6509 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U6510 ( .A1(n5116), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5117) );
  MUX2_X1 U6511 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5117), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5119) );
  INV_X1 U6512 ( .A(n5118), .ZN(n9463) );
  NAND2_X1 U6513 ( .A1(n5390), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5129) );
  INV_X1 U6514 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5120) );
  OR2_X1 U6515 ( .A1(n5456), .A2(n5120), .ZN(n5128) );
  NAND2_X1 U6516 ( .A1(n5124), .A2(n5123), .ZN(n5399) );
  NAND2_X1 U6517 ( .A1(n5470), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6518 ( .A1(n5490), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5492) );
  INV_X1 U6519 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5349) );
  INV_X1 U6520 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6521 ( .A1(n5327), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5312) );
  INV_X1 U6522 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5298) );
  INV_X1 U6523 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6524 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n5121) );
  AND2_X1 U6525 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n5122) );
  NAND2_X1 U6526 ( .A1(n5227), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5210) );
  INV_X1 U6527 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9992) );
  INV_X1 U6528 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8823) );
  NAND2_X1 U6529 ( .A1(n5186), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5176) );
  INV_X1 U6530 ( .A(n5176), .ZN(n5156) );
  NAND2_X1 U6531 ( .A1(n5156), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5155) );
  INV_X1 U6532 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U6533 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n5166), .ZN(n5525) );
  INV_X1 U6534 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8947) );
  NOR2_X1 U6535 ( .A1(n5525), .A2(n8947), .ZN(n5539) );
  NAND2_X1 U6536 ( .A1(n5539), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5538) );
  INV_X1 U6537 ( .A(n5538), .ZN(n5135) );
  NAND2_X1 U6538 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(n5135), .ZN(n9139) );
  OR2_X1 U6539 ( .A1(n5540), .A2(n9139), .ZN(n5127) );
  INV_X1 U6540 ( .A(n9470), .ZN(n5124) );
  INV_X1 U6541 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5125) );
  OR2_X1 U6542 ( .A1(n5560), .A2(n5125), .ZN(n5126) );
  NAND4_X1 U6543 ( .A1(n5129), .A2(n5128), .A3(n5127), .A4(n5126), .ZN(n9155)
         );
  AND2_X1 U6544 ( .A1(n9361), .A2(n9155), .ZN(n5593) );
  OR2_X1 U6545 ( .A1(n5419), .A2(n9478), .ZN(n5132) );
  INV_X1 U6546 ( .A(n5560), .ZN(n5526) );
  NAND2_X1 U6547 ( .A1(n5526), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5140) );
  INV_X1 U6548 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5134) );
  OR2_X1 U6549 ( .A1(n5562), .A2(n5134), .ZN(n5139) );
  OAI21_X1 U6550 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(n5135), .A(n9139), .ZN(
        n9149) );
  OR2_X1 U6551 ( .A1(n5540), .A2(n9149), .ZN(n5138) );
  INV_X1 U6552 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n5136) );
  OR2_X1 U6553 ( .A1(n5456), .A2(n5136), .ZN(n5137) );
  NAND4_X1 U6554 ( .A1(n5140), .A2(n5139), .A3(n5138), .A4(n5137), .ZN(n9132)
         );
  INV_X1 U6555 ( .A(n5705), .ZN(n5698) );
  INV_X1 U6556 ( .A(n5722), .ZN(n5574) );
  XNOR2_X1 U6557 ( .A(n5142), .B(n5141), .ZN(n7686) );
  NAND2_X1 U6558 ( .A1(n7686), .A2(n5581), .ZN(n5144) );
  OR2_X1 U6559 ( .A1(n5419), .A2(n7690), .ZN(n5143) );
  AOI21_X1 U6560 ( .B1(n5155), .B2(n8871), .A(n5166), .ZN(n9212) );
  INV_X1 U6561 ( .A(n5399), .ZN(n5410) );
  NAND2_X1 U6562 ( .A1(n9212), .A2(n5410), .ZN(n5150) );
  INV_X1 U6563 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6564 ( .A1(n5526), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5146) );
  NAND2_X1 U6565 ( .A1(n5558), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5145) );
  OAI211_X1 U6566 ( .C1(n5562), .C2(n5147), .A(n5146), .B(n5145), .ZN(n5148)
         );
  INV_X1 U6567 ( .A(n5148), .ZN(n5149) );
  NAND2_X1 U6568 ( .A1(n5150), .A2(n5149), .ZN(n9229) );
  INV_X1 U6569 ( .A(n9229), .ZN(n9095) );
  NAND2_X1 U6570 ( .A1(n7542), .A2(n5581), .ZN(n5154) );
  OR2_X1 U6571 ( .A1(n5419), .A2(n7545), .ZN(n5153) );
  NAND2_X1 U6572 ( .A1(n5390), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5161) );
  INV_X1 U6573 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10094) );
  OR2_X1 U6574 ( .A1(n5560), .A2(n10094), .ZN(n5160) );
  OAI21_X1 U6575 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n5156), .A(n5155), .ZN(
        n9222) );
  OR2_X1 U6576 ( .A1(n5540), .A2(n9222), .ZN(n5159) );
  INV_X1 U6577 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n5157) );
  OR2_X1 U6578 ( .A1(n5456), .A2(n5157), .ZN(n5158) );
  NAND4_X1 U6579 ( .A1(n5161), .A2(n5160), .A3(n5159), .A4(n5158), .ZN(n8971)
         );
  NAND2_X1 U6580 ( .A1(n9392), .A2(n9238), .ZN(n5681) );
  XNOR2_X1 U6581 ( .A(n5163), .B(n5162), .ZN(n7738) );
  NAND2_X1 U6582 ( .A1(n7738), .A2(n5581), .ZN(n5165) );
  OR2_X1 U6583 ( .A1(n5419), .A2(n7740), .ZN(n5164) );
  OAI21_X1 U6584 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n5166), .A(n5525), .ZN(
        n9195) );
  INV_X1 U6585 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10118) );
  NAND2_X1 U6586 ( .A1(n5390), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5168) );
  INV_X1 U6587 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n10148) );
  OR2_X1 U6588 ( .A1(n5560), .A2(n10148), .ZN(n5167) );
  OAI211_X1 U6589 ( .C1(n10118), .C2(n5456), .A(n5168), .B(n5167), .ZN(n5169)
         );
  INV_X1 U6590 ( .A(n5169), .ZN(n5170) );
  OAI21_X1 U6591 ( .B1(n9195), .B2(n5540), .A(n5170), .ZN(n9185) );
  INV_X1 U6592 ( .A(n9185), .ZN(n9210) );
  NAND2_X1 U6593 ( .A1(n9382), .A2(n9210), .ZN(n5626) );
  NAND2_X1 U6594 ( .A1(n9389), .A2(n9095), .ZN(n9123) );
  OAI211_X1 U6595 ( .C1(n9124), .C2(n5681), .A(n5626), .B(n9123), .ZN(n5741)
         );
  INV_X1 U6596 ( .A(n5741), .ZN(n5547) );
  OR2_X1 U6597 ( .A1(n9124), .A2(n4836), .ZN(n5674) );
  INV_X1 U6598 ( .A(n5674), .ZN(n5520) );
  XNOR2_X1 U6599 ( .A(n5172), .B(n5171), .ZN(n7508) );
  NAND2_X1 U6600 ( .A1(n7508), .A2(n5581), .ZN(n5174) );
  OR2_X1 U6601 ( .A1(n5419), .A2(n8008), .ZN(n5173) );
  NAND2_X1 U6602 ( .A1(n5390), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5180) );
  INV_X1 U6603 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9999) );
  OR2_X1 U6604 ( .A1(n5560), .A2(n9999), .ZN(n5179) );
  INV_X1 U6605 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n5175) );
  OR2_X1 U6606 ( .A1(n5456), .A2(n5175), .ZN(n5178) );
  OAI21_X1 U6607 ( .B1(n5186), .B2(P1_REG3_REG_22__SCAN_IN), .A(n5176), .ZN(
        n9240) );
  OR2_X1 U6608 ( .A1(n5540), .A2(n9240), .ZN(n5177) );
  AND2_X1 U6609 ( .A1(n9244), .A2(n9228), .ZN(n9121) );
  XNOR2_X1 U6610 ( .A(n5182), .B(n5181), .ZN(n7383) );
  NAND2_X1 U6611 ( .A1(n7383), .A2(n5581), .ZN(n5185) );
  OR2_X1 U6612 ( .A1(n5419), .A2(n5183), .ZN(n5184) );
  NAND2_X1 U6613 ( .A1(n5197), .A2(n8823), .ZN(n5188) );
  INV_X1 U6614 ( .A(n5186), .ZN(n5187) );
  NAND2_X1 U6615 ( .A1(n5188), .A2(n5187), .ZN(n9249) );
  AOI22_X1 U6616 ( .A1(n5390), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n5558), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6617 ( .A1(n5526), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5189) );
  OAI211_X1 U6618 ( .C1(n9249), .C2(n5540), .A(n5190), .B(n5189), .ZN(n9092)
         );
  INV_X1 U6619 ( .A(n9092), .ZN(n9275) );
  OR2_X1 U6620 ( .A1(n9405), .A2(n9275), .ZN(n5596) );
  INV_X1 U6621 ( .A(n5596), .ZN(n5191) );
  NOR2_X1 U6622 ( .A1(n9121), .A2(n5191), .ZN(n5678) );
  INV_X1 U6623 ( .A(n5678), .ZN(n5245) );
  NAND2_X1 U6624 ( .A1(n7359), .A2(n5581), .ZN(n5195) );
  OR2_X1 U6625 ( .A1(n5419), .A2(n7363), .ZN(n5194) );
  NAND2_X1 U6626 ( .A1(n5210), .A2(n9992), .ZN(n5196) );
  NAND2_X1 U6627 ( .A1(n5197), .A2(n5196), .ZN(n9268) );
  NAND2_X1 U6628 ( .A1(n5526), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5198) );
  OAI21_X1 U6629 ( .B1(n9268), .B2(n5540), .A(n5198), .ZN(n5201) );
  INV_X1 U6630 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9269) );
  NAND2_X1 U6631 ( .A1(n5558), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5199) );
  OAI21_X1 U6632 ( .B1(n9269), .B2(n5562), .A(n5199), .ZN(n5200) );
  INV_X1 U6633 ( .A(n9289), .ZN(n9254) );
  XNOR2_X1 U6634 ( .A(n5203), .B(n5202), .ZN(n7186) );
  NAND2_X1 U6635 ( .A1(n7186), .A2(n5581), .ZN(n5209) );
  INV_X1 U6636 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10005) );
  NOR2_X1 U6637 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5586) );
  NAND2_X1 U6638 ( .A1(n5588), .A2(n5586), .ZN(n5206) );
  NAND2_X1 U6639 ( .A1(n5206), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5207) );
  AOI22_X1 U6640 ( .A1(n5502), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9214), .B2(
        n5501), .ZN(n5208) );
  OR2_X1 U6641 ( .A1(n5227), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5211) );
  AND2_X1 U6642 ( .A1(n5211), .A2(n5210), .ZN(n9282) );
  NAND2_X1 U6643 ( .A1(n5410), .A2(n9282), .ZN(n5217) );
  INV_X1 U6644 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5212) );
  OR2_X1 U6645 ( .A1(n5562), .A2(n5212), .ZN(n5216) );
  INV_X1 U6646 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9968) );
  OR2_X1 U6647 ( .A1(n5560), .A2(n9968), .ZN(n5215) );
  INV_X1 U6648 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n5213) );
  OR2_X1 U6649 ( .A1(n5456), .A2(n5213), .ZN(n5214) );
  NAND4_X1 U6650 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n9306)
         );
  INV_X1 U6651 ( .A(n9306), .ZN(n9276) );
  OR2_X1 U6652 ( .A1(n9415), .A2(n9276), .ZN(n5677) );
  NAND2_X1 U6653 ( .A1(n9415), .A2(n9276), .ZN(n9116) );
  XNOR2_X1 U6654 ( .A(n5219), .B(n5218), .ZN(n7077) );
  NAND2_X1 U6655 ( .A1(n7077), .A2(n5581), .ZN(n5225) );
  NAND2_X1 U6656 ( .A1(n5220), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5234) );
  INV_X1 U6657 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6658 ( .A1(n5234), .A2(n5221), .ZN(n5222) );
  NAND2_X1 U6659 ( .A1(n5222), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5223) );
  XNOR2_X1 U6660 ( .A(n5223), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9062) );
  AOI22_X1 U6661 ( .A1(n5502), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9062), .B2(
        n5501), .ZN(n5224) );
  AOI21_X1 U6662 ( .B1(n5257), .B2(P1_REG3_REG_17__SCAN_IN), .A(
        P1_REG3_REG_18__SCAN_IN), .ZN(n5226) );
  NOR2_X1 U6663 ( .A1(n5227), .A2(n5226), .ZN(n9309) );
  NAND2_X1 U6664 ( .A1(n5410), .A2(n9309), .ZN(n5231) );
  INV_X1 U6665 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9297) );
  OR2_X1 U6666 ( .A1(n5562), .A2(n9297), .ZN(n5230) );
  INV_X1 U6667 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10163) );
  OR2_X1 U6668 ( .A1(n5456), .A2(n10163), .ZN(n5229) );
  INV_X1 U6669 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10164) );
  OR2_X1 U6670 ( .A1(n5560), .A2(n10164), .ZN(n5228) );
  NAND4_X1 U6671 ( .A1(n5231), .A2(n5230), .A3(n5229), .A4(n5228), .ZN(n9288)
         );
  INV_X1 U6672 ( .A(n9288), .ZN(n9328) );
  NAND2_X1 U6673 ( .A1(n9419), .A2(n9328), .ZN(n9114) );
  OR2_X1 U6674 ( .A1(n9419), .A2(n9328), .ZN(n5667) );
  XNOR2_X1 U6675 ( .A(n5233), .B(n5232), .ZN(n6911) );
  NAND2_X1 U6676 ( .A1(n6911), .A2(n5581), .ZN(n5236) );
  XNOR2_X1 U6677 ( .A(n5234), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9050) );
  AOI22_X1 U6678 ( .A1(n5502), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5501), .B2(
        n9050), .ZN(n5235) );
  NAND2_X1 U6679 ( .A1(n5390), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5242) );
  INV_X1 U6680 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n5237) );
  OR2_X1 U6681 ( .A1(n5456), .A2(n5237), .ZN(n5241) );
  XNOR2_X1 U6682 ( .A(n5257), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9320) );
  OR2_X1 U6683 ( .A1(n5540), .A2(n9320), .ZN(n5240) );
  INV_X1 U6684 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5238) );
  OR2_X1 U6685 ( .A1(n5560), .A2(n5238), .ZN(n5239) );
  NAND4_X1 U6686 ( .A1(n5242), .A2(n5241), .A3(n5240), .A4(n5239), .ZN(n9304)
         );
  INV_X1 U6687 ( .A(n9304), .ZN(n9347) );
  OR2_X1 U6688 ( .A1(n9426), .A2(n9347), .ZN(n9299) );
  NAND2_X1 U6689 ( .A1(n5667), .A2(n9299), .ZN(n9115) );
  NAND3_X1 U6690 ( .A1(n9116), .A2(n9114), .A3(n9115), .ZN(n5243) );
  NAND3_X1 U6691 ( .A1(n9117), .A2(n5677), .A3(n5243), .ZN(n5244) );
  OR2_X1 U6692 ( .A1(n5245), .A2(n5244), .ZN(n5249) );
  INV_X1 U6693 ( .A(n9121), .ZN(n5248) );
  AND2_X1 U6694 ( .A1(n9411), .A2(n9254), .ZN(n9118) );
  NAND2_X1 U6695 ( .A1(n5596), .A2(n9118), .ZN(n5246) );
  NAND2_X1 U6696 ( .A1(n9405), .A2(n9275), .ZN(n5672) );
  AND2_X1 U6697 ( .A1(n5246), .A2(n5672), .ZN(n5247) );
  NAND2_X1 U6698 ( .A1(n9120), .A2(n5247), .ZN(n5517) );
  NAND2_X1 U6699 ( .A1(n5248), .A2(n5517), .ZN(n5680) );
  NAND2_X1 U6700 ( .A1(n5249), .A2(n5680), .ZN(n5723) );
  AND2_X1 U6701 ( .A1(n9426), .A2(n9347), .ZN(n9113) );
  XNOR2_X1 U6702 ( .A(n5251), .B(n5250), .ZN(n6932) );
  NAND2_X1 U6703 ( .A1(n6932), .A2(n5581), .ZN(n5255) );
  OR2_X1 U6704 ( .A1(n5252), .A2(n5449), .ZN(n5253) );
  XNOR2_X1 U6705 ( .A(n5253), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9034) );
  AOI22_X1 U6706 ( .A1(n5502), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5501), .B2(
        n9034), .ZN(n5254) );
  NAND2_X1 U6707 ( .A1(n5390), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5262) );
  INV_X1 U6708 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10096) );
  OR2_X1 U6709 ( .A1(n5456), .A2(n10096), .ZN(n5261) );
  NOR2_X1 U6710 ( .A1(n5380), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5256) );
  OR2_X1 U6711 ( .A1(n5257), .A2(n5256), .ZN(n9340) );
  OR2_X1 U6712 ( .A1(n5540), .A2(n9340), .ZN(n5260) );
  INV_X1 U6713 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n5258) );
  OR2_X1 U6714 ( .A1(n5560), .A2(n5258), .ZN(n5259) );
  NAND4_X1 U6715 ( .A1(n5262), .A2(n5261), .A3(n5260), .A4(n5259), .ZN(n9087)
         );
  INV_X1 U6716 ( .A(n9087), .ZN(n9327) );
  NAND2_X1 U6717 ( .A1(n9431), .A2(n9327), .ZN(n9111) );
  INV_X1 U6718 ( .A(n9111), .ZN(n5263) );
  NOR2_X1 U6719 ( .A1(n9113), .A2(n5263), .ZN(n5264) );
  NAND2_X1 U6720 ( .A1(n5264), .A2(n9114), .ZN(n5514) );
  XNOR2_X1 U6721 ( .A(n5266), .B(n5265), .ZN(n6662) );
  NAND2_X1 U6722 ( .A1(n6662), .A2(n5581), .ZN(n5269) );
  OR2_X1 U6723 ( .A1(n5267), .A2(n5449), .ZN(n5371) );
  XNOR2_X1 U6724 ( .A(n5371), .B(P1_IR_REG_14__SCAN_IN), .ZN(n6373) );
  AOI22_X1 U6725 ( .A1(n5502), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5501), .B2(
        n6373), .ZN(n5268) );
  NAND2_X1 U6726 ( .A1(n5558), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5274) );
  INV_X1 U6727 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7707) );
  OR2_X1 U6728 ( .A1(n5562), .A2(n7707), .ZN(n5273) );
  INV_X1 U6729 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5270) );
  XNOR2_X1 U6730 ( .A(n5378), .B(n5270), .ZN(n8791) );
  OR2_X1 U6731 ( .A1(n5540), .A2(n8791), .ZN(n5272) );
  INV_X1 U6732 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6372) );
  OR2_X1 U6733 ( .A1(n5560), .A2(n6372), .ZN(n5271) );
  NAND4_X1 U6734 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n8972)
         );
  INV_X1 U6735 ( .A(n8972), .ZN(n7757) );
  NOR2_X1 U6736 ( .A1(n8793), .A2(n7757), .ZN(n7752) );
  XNOR2_X1 U6737 ( .A(n5276), .B(n5275), .ZN(n6656) );
  NAND2_X1 U6738 ( .A1(n6656), .A2(n5581), .ZN(n5280) );
  OR2_X1 U6739 ( .A1(n5277), .A2(n5449), .ZN(n5278) );
  XNOR2_X1 U6740 ( .A(n5278), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7083) );
  AOI22_X1 U6741 ( .A1(n5502), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5501), .B2(
        n7083), .ZN(n5279) );
  NAND2_X1 U6742 ( .A1(n5390), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5287) );
  INV_X1 U6743 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6366) );
  OR2_X1 U6744 ( .A1(n5560), .A2(n6366), .ZN(n5286) );
  NAND2_X1 U6745 ( .A1(n5300), .A2(n5281), .ZN(n5282) );
  NAND2_X1 U6746 ( .A1(n5378), .A2(n5282), .ZN(n8907) );
  OR2_X1 U6747 ( .A1(n5540), .A2(n8907), .ZN(n5285) );
  INV_X1 U6748 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5283) );
  OR2_X1 U6749 ( .A1(n5456), .A2(n5283), .ZN(n5284) );
  NAND4_X1 U6750 ( .A1(n5287), .A2(n5286), .A3(n5285), .A4(n5284), .ZN(n8973)
         );
  OR2_X1 U6751 ( .A1(n8898), .A2(n8788), .ZN(n5599) );
  INV_X1 U6752 ( .A(n5599), .ZN(n5288) );
  NOR2_X1 U6753 ( .A1(n7752), .A2(n5288), .ZN(n5648) );
  INV_X1 U6754 ( .A(n5648), .ZN(n5289) );
  NAND2_X1 U6755 ( .A1(n8793), .A2(n7757), .ZN(n5290) );
  NAND2_X1 U6756 ( .A1(n5289), .A2(n5290), .ZN(n5657) );
  NAND2_X1 U6757 ( .A1(n8898), .A2(n8788), .ZN(n7694) );
  NAND2_X1 U6758 ( .A1(n5290), .A2(n7694), .ZN(n5654) );
  INV_X1 U6759 ( .A(n5654), .ZN(n5366) );
  NAND2_X1 U6760 ( .A1(n6641), .A2(n5581), .ZN(n5296) );
  NAND2_X1 U6761 ( .A1(n5293), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5294) );
  XNOR2_X1 U6762 ( .A(n5294), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6642) );
  AOI22_X1 U6763 ( .A1(n5502), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5501), .B2(
        n6642), .ZN(n5295) );
  NAND2_X1 U6764 ( .A1(n5390), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5304) );
  INV_X1 U6765 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5297) );
  OR2_X1 U6766 ( .A1(n5456), .A2(n5297), .ZN(n5303) );
  NAND2_X1 U6767 ( .A1(n5312), .A2(n5298), .ZN(n5299) );
  NAND2_X1 U6768 ( .A1(n5300), .A2(n5299), .ZN(n8835) );
  OR2_X1 U6769 ( .A1(n5540), .A2(n8835), .ZN(n5302) );
  INV_X1 U6770 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6367) );
  OR2_X1 U6771 ( .A1(n5560), .A2(n6367), .ZN(n5301) );
  NAND4_X1 U6772 ( .A1(n5304), .A2(n5303), .A3(n5302), .A4(n5301), .ZN(n8974)
         );
  XNOR2_X1 U6773 ( .A(n5306), .B(n5305), .ZN(n6428) );
  NAND2_X1 U6774 ( .A1(n6428), .A2(n5581), .ZN(n5309) );
  NAND2_X1 U6775 ( .A1(n4484), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5307) );
  XNOR2_X1 U6776 ( .A(n5307), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6371) );
  AOI22_X1 U6777 ( .A1(n5502), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5501), .B2(
        n6371), .ZN(n5308) );
  NAND2_X1 U6778 ( .A1(n5309), .A2(n5308), .ZN(n8930) );
  NAND2_X1 U6779 ( .A1(n5558), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5316) );
  INV_X1 U6780 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7646) );
  OR2_X1 U6781 ( .A1(n5562), .A2(n7646), .ZN(n5315) );
  INV_X1 U6782 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5310) );
  OR2_X1 U6783 ( .A1(n5560), .A2(n5310), .ZN(n5314) );
  OR2_X1 U6784 ( .A1(n5327), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U6785 ( .A1(n5312), .A2(n5311), .ZN(n8924) );
  OR2_X1 U6786 ( .A1(n5540), .A2(n8924), .ZN(n5313) );
  NAND4_X1 U6787 ( .A1(n5316), .A2(n5315), .A3(n5314), .A4(n5313), .ZN(n8975)
         );
  NAND2_X1 U6788 ( .A1(n8930), .A2(n9493), .ZN(n7656) );
  NAND2_X1 U6789 ( .A1(n5637), .A2(n7656), .ZN(n7691) );
  OR2_X1 U6790 ( .A1(n5319), .A2(n5318), .ZN(n5320) );
  NAND2_X1 U6791 ( .A1(n5317), .A2(n5320), .ZN(n6418) );
  NAND2_X1 U6792 ( .A1(n6418), .A2(n5581), .ZN(n5324) );
  NAND2_X1 U6793 ( .A1(n5321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5322) );
  XNOR2_X1 U6794 ( .A(n5322), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6370) );
  AOI22_X1 U6795 ( .A1(n5502), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5501), .B2(
        n6370), .ZN(n5323) );
  NAND2_X1 U6796 ( .A1(n5390), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5332) );
  INV_X1 U6797 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5325) );
  OR2_X1 U6798 ( .A1(n5456), .A2(n5325), .ZN(n5331) );
  NOR2_X1 U6799 ( .A1(n5340), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5326) );
  OR2_X1 U6800 ( .A1(n5327), .A2(n5326), .ZN(n9497) );
  OR2_X1 U6801 ( .A1(n5540), .A2(n9497), .ZN(n5330) );
  INV_X1 U6802 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5328) );
  OR2_X1 U6803 ( .A1(n5560), .A2(n5328), .ZN(n5329) );
  NAND4_X1 U6804 ( .A1(n5332), .A2(n5331), .A3(n5330), .A4(n5329), .ZN(n8976)
         );
  INV_X1 U6805 ( .A(n8976), .ZN(n7641) );
  NAND2_X1 U6806 ( .A1(n9501), .A2(n7641), .ZN(n5638) );
  XNOR2_X1 U6807 ( .A(n5333), .B(n5334), .ZN(n6414) );
  NAND2_X1 U6808 ( .A1(n6414), .A2(n5581), .ZN(n5338) );
  OR2_X1 U6809 ( .A1(n5335), .A2(n5449), .ZN(n5336) );
  XNOR2_X1 U6810 ( .A(n5336), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6369) );
  AOI22_X1 U6811 ( .A1(n5502), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5501), .B2(
        n6369), .ZN(n5337) );
  NAND2_X1 U6812 ( .A1(n5390), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5346) );
  AND2_X1 U6813 ( .A1(n5351), .A2(n5339), .ZN(n5341) );
  OR2_X1 U6814 ( .A1(n5341), .A2(n5340), .ZN(n8883) );
  OR2_X1 U6815 ( .A1(n5540), .A2(n8883), .ZN(n5345) );
  INV_X1 U6816 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5342) );
  OR2_X1 U6817 ( .A1(n5456), .A2(n5342), .ZN(n5344) );
  INV_X1 U6818 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6345) );
  OR2_X1 U6819 ( .A1(n5560), .A2(n6345), .ZN(n5343) );
  NAND4_X1 U6820 ( .A1(n5346), .A2(n5345), .A3(n5344), .A4(n5343), .ZN(n8977)
         );
  INV_X1 U6821 ( .A(n8977), .ZN(n9490) );
  NAND2_X1 U6822 ( .A1(n8885), .A2(n9490), .ZN(n9484) );
  NAND2_X1 U6823 ( .A1(n5638), .A2(n9484), .ZN(n5347) );
  OR2_X1 U6824 ( .A1(n9501), .A2(n7641), .ZN(n5606) );
  NAND2_X1 U6825 ( .A1(n5347), .A2(n5606), .ZN(n7638) );
  INV_X1 U6826 ( .A(n7638), .ZN(n5348) );
  OR2_X1 U6827 ( .A1(n7691), .A2(n5348), .ZN(n5510) );
  OR2_X1 U6828 ( .A1(n8885), .A2(n9490), .ZN(n9482) );
  NAND2_X1 U6829 ( .A1(n5606), .A2(n9482), .ZN(n7637) );
  NAND2_X1 U6830 ( .A1(n5526), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5356) );
  INV_X1 U6831 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7428) );
  OR2_X1 U6832 ( .A1(n5562), .A2(n7428), .ZN(n5355) );
  NAND2_X1 U6833 ( .A1(n5492), .A2(n5349), .ZN(n5350) );
  NAND2_X1 U6834 ( .A1(n5351), .A2(n5350), .ZN(n7534) );
  OR2_X1 U6835 ( .A1(n5540), .A2(n7534), .ZN(n5354) );
  INV_X1 U6836 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5352) );
  OR2_X1 U6837 ( .A1(n5456), .A2(n5352), .ZN(n5353) );
  XNOR2_X1 U6838 ( .A(n5358), .B(n5357), .ZN(n6409) );
  NAND2_X1 U6839 ( .A1(n6409), .A2(n5581), .ZN(n5362) );
  OR2_X1 U6840 ( .A1(n5481), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5483) );
  NOR2_X1 U6841 ( .A1(n5483), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6842 ( .A1(n5450), .A2(n5359), .ZN(n5499) );
  OAI21_X1 U6843 ( .B1(n5499), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5360) );
  XNOR2_X1 U6844 ( .A(n5360), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6344) );
  AOI22_X1 U6845 ( .A1(n5502), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5501), .B2(
        n6344), .ZN(n5361) );
  INV_X1 U6846 ( .A(n7512), .ZN(n5363) );
  NOR2_X1 U6847 ( .A1(n7637), .A2(n5363), .ZN(n5642) );
  OR2_X1 U6848 ( .A1(n8837), .A2(n8906), .ZN(n5647) );
  OR2_X1 U6849 ( .A1(n8930), .A2(n9493), .ZN(n7657) );
  NAND2_X1 U6850 ( .A1(n5647), .A2(n7657), .ZN(n5364) );
  NAND2_X1 U6851 ( .A1(n5364), .A2(n5637), .ZN(n7693) );
  OAI21_X1 U6852 ( .B1(n5510), .B2(n5642), .A(n7693), .ZN(n5365) );
  NAND2_X1 U6853 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  NAND2_X1 U6854 ( .A1(n5657), .A2(n5367), .ZN(n5387) );
  XNOR2_X1 U6855 ( .A(n5369), .B(n5368), .ZN(n6743) );
  NAND2_X1 U6856 ( .A1(n6743), .A2(n5581), .ZN(n5377) );
  INV_X1 U6857 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5370) );
  NAND2_X1 U6858 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  NAND2_X1 U6859 ( .A1(n5372), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5374) );
  INV_X1 U6860 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5373) );
  XNOR2_X1 U6861 ( .A(n5374), .B(n5373), .ZN(n9017) );
  INV_X1 U6862 ( .A(n9017), .ZN(n5375) );
  AOI22_X1 U6863 ( .A1(n5502), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5501), .B2(
        n5375), .ZN(n5376) );
  NAND2_X1 U6864 ( .A1(n5526), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5386) );
  INV_X1 U6865 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7764) );
  OR2_X1 U6866 ( .A1(n5562), .A2(n7764), .ZN(n5385) );
  INV_X1 U6867 ( .A(n5378), .ZN(n5379) );
  AOI21_X1 U6868 ( .B1(n5379), .B2(P1_REG3_REG_14__SCAN_IN), .A(
        P1_REG3_REG_15__SCAN_IN), .ZN(n5381) );
  OR2_X1 U6869 ( .A1(n5381), .A2(n5380), .ZN(n8964) );
  OR2_X1 U6870 ( .A1(n5540), .A2(n8964), .ZN(n5384) );
  INV_X1 U6871 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5382) );
  OR2_X1 U6872 ( .A1(n5456), .A2(n5382), .ZN(n5383) );
  NAND4_X1 U6873 ( .A1(n5386), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(n10214)
         );
  AND2_X1 U6874 ( .A1(n9084), .A2(n9348), .ZN(n9108) );
  INV_X1 U6875 ( .A(n9108), .ZN(n5660) );
  NAND2_X1 U6876 ( .A1(n5387), .A2(n5660), .ZN(n5388) );
  OR2_X1 U6877 ( .A1(n9431), .A2(n9327), .ZN(n9110) );
  AND3_X1 U6878 ( .A1(n5388), .A2(n9110), .A3(n9107), .ZN(n5389) );
  OR2_X1 U6879 ( .A1(n5514), .A2(n5389), .ZN(n5512) );
  INV_X1 U6880 ( .A(n5512), .ZN(n5738) );
  INV_X1 U6881 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7159) );
  NAND2_X1 U6882 ( .A1(n5411), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5392) );
  INV_X1 U6883 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6591) );
  XNOR2_X1 U6884 ( .A(n5396), .B(n5395), .ZN(n6385) );
  INV_X1 U6885 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6386) );
  INV_X1 U6886 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6887 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5397) );
  XNOR2_X1 U6888 ( .A(n5397), .B(n5398), .ZN(n6590) );
  XNOR2_X1 U6889 ( .A(n6818), .B(n7162), .ZN(n6965) );
  NAND2_X1 U6890 ( .A1(n5390), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5403) );
  INV_X1 U6891 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7209) );
  NAND2_X1 U6892 ( .A1(n5411), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5400) );
  NAND4_X1 U6893 ( .A1(n5403), .A2(n5402), .A3(n5401), .A4(n5400), .ZN(n6791)
         );
  NAND2_X1 U6894 ( .A1(n6384), .A2(SI_0_), .ZN(n5405) );
  INV_X1 U6895 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6896 ( .A1(n5405), .A2(n5404), .ZN(n5407) );
  AND2_X1 U6897 ( .A1(n5407), .A2(n5406), .ZN(n9480) );
  MUX2_X1 U6898 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9480), .S(n5408), .Z(n7208) );
  NAND2_X1 U6899 ( .A1(n6818), .A2(n7162), .ZN(n5409) );
  NAND2_X1 U6900 ( .A1(n5390), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6901 ( .A1(n5410), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6902 ( .A1(n5411), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5414) );
  INV_X1 U6903 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6335) );
  AND4_X2 U6904 ( .A1(n5416), .A2(n5415), .A3(n5414), .A4(n5413), .ZN(n6826)
         );
  XNOR2_X1 U6905 ( .A(n5418), .B(n5417), .ZN(n6395) );
  OR2_X1 U6906 ( .A1(n5480), .A2(n6395), .ZN(n5425) );
  OR2_X1 U6907 ( .A1(n5419), .A2(n6396), .ZN(n5424) );
  INV_X1 U6908 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6909 ( .A1(n5422), .A2(n5421), .ZN(n5463) );
  OR2_X1 U6910 ( .A1(n5408), .A2(n6861), .ZN(n5423) );
  INV_X1 U6911 ( .A(n6826), .ZN(n8984) );
  NAND2_X1 U6912 ( .A1(n6826), .A2(n7305), .ZN(n5426) );
  NAND2_X1 U6913 ( .A1(n5427), .A2(n5426), .ZN(n6977) );
  NAND2_X1 U6914 ( .A1(n5558), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5432) );
  INV_X1 U6915 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5428) );
  OR2_X1 U6916 ( .A1(n5562), .A2(n5428), .ZN(n5431) );
  OAI21_X1 U6917 ( .B1(n5470), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5440), .ZN(
        n9604) );
  OR2_X1 U6918 ( .A1(n5540), .A2(n9604), .ZN(n5430) );
  INV_X1 U6919 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6339) );
  OR2_X1 U6920 ( .A1(n5560), .A2(n6339), .ZN(n5429) );
  AND4_X2 U6921 ( .A1(n5432), .A2(n5431), .A3(n5430), .A4(n5429), .ZN(n7315)
         );
  XNOR2_X1 U6922 ( .A(n5434), .B(n5433), .ZN(n6391) );
  OR2_X1 U6923 ( .A1(n5480), .A2(n6391), .ZN(n5438) );
  OR2_X1 U6924 ( .A1(n5419), .A2(n6392), .ZN(n5437) );
  NAND2_X1 U6925 ( .A1(n5483), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5435) );
  XNOR2_X1 U6926 ( .A(n5435), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6338) );
  INV_X1 U6927 ( .A(n6338), .ZN(n9568) );
  OR2_X1 U6928 ( .A1(n5408), .A2(n9568), .ZN(n5436) );
  NAND2_X1 U6929 ( .A1(n5558), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5446) );
  INV_X1 U6930 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7320) );
  OR2_X1 U6931 ( .A1(n5562), .A2(n7320), .ZN(n5445) );
  AND2_X1 U6932 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  OR2_X1 U6933 ( .A1(n5441), .A2(n5490), .ZN(n7319) );
  OR2_X1 U6934 ( .A1(n5540), .A2(n7319), .ZN(n5444) );
  INV_X1 U6935 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5442) );
  OR2_X1 U6936 ( .A1(n5560), .A2(n5442), .ZN(n5443) );
  XNOR2_X1 U6937 ( .A(n5448), .B(n5447), .ZN(n6398) );
  OR2_X1 U6938 ( .A1(n6398), .A2(n5480), .ZN(n5454) );
  INV_X1 U6939 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9989) );
  OR2_X1 U6940 ( .A1(n5419), .A2(n9989), .ZN(n5453) );
  OR2_X1 U6941 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  XNOR2_X1 U6942 ( .A(n5451), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6341) );
  INV_X1 U6943 ( .A(n6341), .ZN(n6635) );
  OR2_X1 U6944 ( .A1(n5408), .A2(n6635), .ZN(n5452) );
  OR2_X1 U6945 ( .A1(n7378), .A2(n7326), .ZN(n5603) );
  AND2_X1 U6946 ( .A1(n5631), .A2(n5603), .ZN(n5725) );
  NAND2_X1 U6947 ( .A1(n5390), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5460) );
  INV_X1 U6948 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5455) );
  OR2_X1 U6949 ( .A1(n5456), .A2(n5455), .ZN(n5458) );
  INV_X1 U6950 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6333) );
  OR2_X1 U6951 ( .A1(n5560), .A2(n6333), .ZN(n5457) );
  OR2_X1 U6952 ( .A1(n5419), .A2(n6388), .ZN(n5468) );
  XNOR2_X1 U6953 ( .A(n5462), .B(n5461), .ZN(n6389) );
  OR2_X1 U6954 ( .A1(n5480), .A2(n6389), .ZN(n5467) );
  NAND2_X1 U6955 ( .A1(n5463), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5465) );
  INV_X1 U6956 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5464) );
  XNOR2_X1 U6957 ( .A(n5465), .B(n5464), .ZN(n6567) );
  OR2_X1 U6958 ( .A1(n5408), .A2(n6567), .ZN(n5466) );
  NAND2_X1 U6959 ( .A1(n5558), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5477) );
  INV_X1 U6960 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6332) );
  OR2_X1 U6961 ( .A1(n5560), .A2(n6332), .ZN(n5476) );
  INV_X1 U6962 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5469) );
  OR2_X1 U6963 ( .A1(n5562), .A2(n5469), .ZN(n5475) );
  INV_X1 U6964 ( .A(n5470), .ZN(n5473) );
  INV_X1 U6965 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6844) );
  INV_X1 U6966 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U6967 ( .A1(n6844), .A2(n5471), .ZN(n5472) );
  NAND2_X1 U6968 ( .A1(n5473), .A2(n5472), .ZN(n7263) );
  OR2_X1 U6969 ( .A1(n5540), .A2(n7263), .ZN(n5474) );
  XNOR2_X1 U6970 ( .A(n5479), .B(n5478), .ZN(n6393) );
  OR2_X1 U6971 ( .A1(n5480), .A2(n6393), .ZN(n5487) );
  OR2_X1 U6972 ( .A1(n5419), .A2(n6394), .ZN(n5486) );
  NAND2_X1 U6973 ( .A1(n5481), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5482) );
  MUX2_X1 U6974 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5482), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5484) );
  NAND2_X1 U6975 ( .A1(n5484), .A2(n5483), .ZN(n9562) );
  OR2_X1 U6976 ( .A1(n5408), .A2(n9562), .ZN(n5485) );
  OAI21_X1 U6977 ( .B1(n7297), .B2(n6973), .A(n5629), .ZN(n5488) );
  INV_X1 U6978 ( .A(n5488), .ZN(n5505) );
  NAND2_X1 U6979 ( .A1(n5558), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5496) );
  INV_X1 U6980 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5489) );
  OR2_X1 U6981 ( .A1(n5560), .A2(n5489), .ZN(n5495) );
  INV_X1 U6982 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7284) );
  OR2_X1 U6983 ( .A1(n5562), .A2(n7284), .ZN(n5494) );
  OR2_X1 U6984 ( .A1(n5490), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5491) );
  NAND2_X1 U6985 ( .A1(n5492), .A2(n5491), .ZN(n7375) );
  OR2_X1 U6986 ( .A1(n5540), .A2(n7375), .ZN(n5493) );
  XNOR2_X1 U6987 ( .A(n5498), .B(n5497), .ZN(n6400) );
  NAND2_X1 U6988 ( .A1(n6400), .A2(n5581), .ZN(n5504) );
  NAND2_X1 U6989 ( .A1(n5499), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5500) );
  XNOR2_X1 U6990 ( .A(n5500), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6343) );
  AOI22_X1 U6991 ( .A1(n5502), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5501), .B2(
        n6343), .ZN(n5503) );
  AND3_X1 U6992 ( .A1(n5725), .A2(n5505), .A3(n5735), .ZN(n5733) );
  NAND2_X1 U6993 ( .A1(n5735), .A2(n5603), .ZN(n5632) );
  INV_X1 U6994 ( .A(n5632), .ZN(n5509) );
  NAND2_X1 U6995 ( .A1(n7068), .A2(n7265), .ZN(n5600) );
  INV_X1 U6996 ( .A(n5600), .ZN(n5628) );
  NAND2_X1 U6997 ( .A1(n7297), .A2(n6973), .ZN(n5627) );
  INV_X1 U6998 ( .A(n5627), .ZN(n5506) );
  OAI211_X1 U6999 ( .C1(n5628), .C2(n5506), .A(n5631), .B(n5629), .ZN(n5507)
         );
  NAND2_X1 U7000 ( .A1(n7378), .A2(n7326), .ZN(n5727) );
  NAND2_X1 U7001 ( .A1(n7315), .A2(n7137), .ZN(n5630) );
  NAND3_X1 U7002 ( .A1(n5507), .A2(n5727), .A3(n5630), .ZN(n5508) );
  AOI22_X1 U7003 ( .A1(n6977), .A2(n5733), .B1(n5509), .B2(n5508), .ZN(n5518)
         );
  NAND2_X1 U7004 ( .A1(n7527), .A2(n7537), .ZN(n5607) );
  INV_X1 U7005 ( .A(n5607), .ZN(n5643) );
  NAND2_X1 U7006 ( .A1(n7423), .A2(n7387), .ZN(n7419) );
  INV_X1 U7007 ( .A(n7419), .ZN(n5633) );
  OR3_X1 U7008 ( .A1(n5510), .A2(n5643), .A3(n5633), .ZN(n5511) );
  OR3_X1 U7009 ( .A1(n9108), .A2(n5511), .A3(n5654), .ZN(n5513) );
  OAI21_X1 U7010 ( .B1(n5514), .B2(n5513), .A(n5512), .ZN(n5515) );
  NAND2_X1 U7011 ( .A1(n5515), .A2(n9116), .ZN(n5516) );
  NOR2_X1 U7012 ( .A1(n5517), .A2(n5516), .ZN(n5736) );
  OAI21_X1 U7013 ( .B1(n5738), .B2(n5518), .A(n5736), .ZN(n5519) );
  NAND3_X1 U7014 ( .A1(n5520), .A2(n5723), .A3(n5519), .ZN(n5546) );
  OR2_X1 U7015 ( .A1(n5419), .A2(n7827), .ZN(n5523) );
  AOI21_X1 U7016 ( .B1(n5525), .B2(n8947), .A(n5539), .ZN(n9177) );
  NAND2_X1 U7017 ( .A1(n9177), .A2(n5410), .ZN(n5532) );
  INV_X1 U7018 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5529) );
  NAND2_X1 U7019 ( .A1(n5526), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5528) );
  NAND2_X1 U7020 ( .A1(n5558), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5527) );
  OAI211_X1 U7021 ( .C1(n5562), .C2(n5529), .A(n5528), .B(n5527), .ZN(n5530)
         );
  INV_X1 U7022 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U7023 ( .A1(n5532), .A2(n5531), .ZN(n9201) );
  INV_X1 U7024 ( .A(n9201), .ZN(n9169) );
  OR2_X1 U7025 ( .A1(n9377), .A2(n9169), .ZN(n5692) );
  NAND2_X1 U7026 ( .A1(n5692), .A2(n9180), .ZN(n9127) );
  NAND2_X1 U7027 ( .A1(n8766), .A2(n5581), .ZN(n5536) );
  OR2_X1 U7028 ( .A1(n5419), .A2(n7824), .ZN(n5535) );
  NAND2_X1 U7029 ( .A1(n5558), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5545) );
  INV_X1 U7030 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5537) );
  OR2_X1 U7031 ( .A1(n5562), .A2(n5537), .ZN(n5544) );
  OAI21_X1 U7032 ( .B1(P1_REG3_REG_27__SCAN_IN), .B2(n5539), .A(n5538), .ZN(
        n9162) );
  OR2_X1 U7033 ( .A1(n5540), .A2(n9162), .ZN(n5543) );
  INV_X1 U7034 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5541) );
  OR2_X1 U7035 ( .A1(n5560), .A2(n5541), .ZN(n5542) );
  NAND4_X1 U7036 ( .A1(n5545), .A2(n5544), .A3(n5543), .A4(n5542), .ZN(n9186)
         );
  INV_X1 U7037 ( .A(n5704), .ZN(n9128) );
  AOI211_X1 U7038 ( .C1(n5547), .C2(n5546), .A(n9127), .B(n9128), .ZN(n5573)
         );
  NAND2_X1 U7039 ( .A1(n9373), .A2(n9103), .ZN(n5689) );
  NAND2_X1 U7040 ( .A1(n9129), .A2(n5689), .ZN(n5697) );
  NAND2_X1 U7041 ( .A1(n9377), .A2(n9169), .ZN(n9126) );
  INV_X1 U7042 ( .A(n9126), .ZN(n5690) );
  AND2_X1 U7043 ( .A1(n5704), .A2(n5690), .ZN(n5548) );
  NOR2_X1 U7044 ( .A1(n5697), .A2(n5548), .ZN(n5549) );
  OR2_X1 U7045 ( .A1(n5722), .A2(n5549), .ZN(n5553) );
  INV_X1 U7046 ( .A(n9361), .ZN(n5551) );
  INV_X1 U7047 ( .A(n9155), .ZN(n5550) );
  INV_X1 U7048 ( .A(n5625), .ZN(n5552) );
  NAND2_X1 U7049 ( .A1(n5553), .A2(n5552), .ZN(n5743) );
  INV_X1 U7050 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U7051 ( .A1(n5558), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5556) );
  INV_X1 U7052 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5554) );
  OR2_X1 U7053 ( .A1(n5560), .A2(n5554), .ZN(n5555) );
  OAI211_X1 U7054 ( .C1(n5562), .C2(n5557), .A(n5556), .B(n5555), .ZN(n9133)
         );
  NAND2_X1 U7055 ( .A1(n5558), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5565) );
  INV_X1 U7056 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5559) );
  OR2_X1 U7057 ( .A1(n5560), .A2(n5559), .ZN(n5564) );
  INV_X1 U7058 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n5561) );
  OR2_X1 U7059 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  AND3_X1 U7060 ( .A1(n5565), .A2(n5564), .A3(n5563), .ZN(n5584) );
  INV_X1 U7061 ( .A(n5584), .ZN(n9076) );
  INV_X1 U7062 ( .A(SI_29_), .ZN(n5566) );
  AND2_X1 U7063 ( .A1(n5567), .A2(n5566), .ZN(n5569) );
  INV_X1 U7064 ( .A(n5567), .ZN(n5568) );
  MUX2_X1 U7065 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6384), .Z(n5576) );
  NAND2_X1 U7066 ( .A1(n8022), .A2(n5581), .ZN(n5572) );
  INV_X1 U7067 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8006) );
  OR2_X1 U7068 ( .A1(n5419), .A2(n8006), .ZN(n5571) );
  AOI21_X1 U7069 ( .B1(n9133), .B2(n9076), .A(n9359), .ZN(n5710) );
  AOI211_X1 U7070 ( .C1(n5574), .C2(n5573), .A(n5743), .B(n5710), .ZN(n5592)
         );
  NAND2_X1 U7071 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  MUX2_X1 U7072 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6380), .Z(n5579) );
  XNOR2_X1 U7073 ( .A(n5579), .B(SI_31_), .ZN(n5580) );
  NAND2_X1 U7074 ( .A1(n8032), .A2(n5581), .ZN(n5583) );
  INV_X1 U7075 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9461) );
  OR2_X1 U7076 ( .A1(n5419), .A2(n9461), .ZN(n5582) );
  NAND2_X1 U7077 ( .A1(n9074), .A2(n5584), .ZN(n5709) );
  INV_X1 U7078 ( .A(n9133), .ZN(n5617) );
  OR2_X1 U7079 ( .A1(n9080), .A2(n5617), .ZN(n5585) );
  AND2_X1 U7080 ( .A1(n5586), .A2(n10146), .ZN(n5587) );
  NAND2_X1 U7081 ( .A1(n5717), .A2(n5754), .ZN(n5589) );
  OR2_X1 U7082 ( .A1(n5590), .A2(n5755), .ZN(n5591) );
  NAND2_X1 U7083 ( .A1(n5590), .A2(n5755), .ZN(n5623) );
  AND2_X2 U7084 ( .A1(n5591), .A2(n5623), .ZN(n5762) );
  OAI211_X1 U7085 ( .C1(n5592), .C2(n5707), .A(n5762), .B(n5750), .ZN(n5622)
         );
  INV_X1 U7086 ( .A(n9154), .ZN(n9147) );
  AND2_X1 U7087 ( .A1(n5704), .A2(n5689), .ZN(n9102) );
  NOR2_X1 U7088 ( .A1(n9377), .A2(n9201), .ZN(n9100) );
  NAND2_X1 U7089 ( .A1(n9377), .A2(n9201), .ZN(n9101) );
  INV_X1 U7090 ( .A(n9101), .ZN(n5594) );
  OR2_X1 U7091 ( .A1(n9100), .A2(n5594), .ZN(n9183) );
  INV_X1 U7092 ( .A(n9200), .ZN(n5615) );
  NAND2_X1 U7093 ( .A1(n9122), .A2(n5681), .ZN(n9227) );
  INV_X1 U7094 ( .A(n9120), .ZN(n5595) );
  OR2_X1 U7095 ( .A1(n5595), .A2(n9121), .ZN(n9236) );
  INV_X1 U7096 ( .A(n9118), .ZN(n5597) );
  NAND2_X1 U7097 ( .A1(n5667), .A2(n9114), .ZN(n9302) );
  INV_X1 U7098 ( .A(n9113), .ZN(n5598) );
  INV_X1 U7099 ( .A(n9315), .ZN(n9324) );
  NAND2_X1 U7100 ( .A1(n7657), .A2(n7656), .ZN(n7636) );
  INV_X1 U7101 ( .A(n7636), .ZN(n7640) );
  INV_X1 U7102 ( .A(n7267), .ZN(n5601) );
  AND2_X1 U7103 ( .A1(n6791), .A2(n7158), .ZN(n5729) );
  NOR2_X1 U7104 ( .A1(n7153), .A2(n5729), .ZN(n6718) );
  AND4_X1 U7105 ( .A1(n7066), .A2(n5602), .A3(n5601), .A4(n6718), .ZN(n5605)
         );
  NAND2_X1 U7106 ( .A1(n5735), .A2(n7419), .ZN(n7280) );
  NAND2_X1 U7107 ( .A1(n5603), .A2(n5727), .ZN(n7311) );
  XNOR2_X1 U7108 ( .A(n7297), .B(n6973), .ZN(n6970) );
  INV_X1 U7109 ( .A(n6970), .ZN(n6976) );
  AND2_X1 U7110 ( .A1(n6976), .A2(n7293), .ZN(n5604) );
  NAND4_X1 U7111 ( .A1(n5605), .A2(n4927), .A3(n7313), .A4(n5604), .ZN(n5608)
         );
  NAND2_X1 U7112 ( .A1(n5606), .A2(n5638), .ZN(n9486) );
  NAND2_X1 U7113 ( .A1(n7512), .A2(n5607), .ZN(n7421) );
  NAND2_X1 U7114 ( .A1(n9482), .A2(n9484), .ZN(n7514) );
  NOR4_X1 U7115 ( .A1(n5608), .A2(n9486), .A3(n7421), .A4(n7514), .ZN(n5609)
         );
  AND4_X1 U7116 ( .A1(n7719), .A2(n4457), .A3(n7640), .A4(n5609), .ZN(n5610)
         );
  XNOR2_X1 U7117 ( .A(n8793), .B(n8972), .ZN(n7753) );
  NAND4_X1 U7118 ( .A1(n9344), .A2(n7755), .A3(n5610), .A4(n7753), .ZN(n5611)
         );
  NOR3_X1 U7119 ( .A1(n9302), .A2(n9324), .A3(n5611), .ZN(n5612) );
  NAND4_X1 U7120 ( .A1(n9257), .A2(n9287), .A3(n9273), .A4(n5612), .ZN(n5613)
         );
  NOR3_X1 U7121 ( .A1(n9227), .A2(n9236), .A3(n5613), .ZN(n5614) );
  XNOR2_X1 U7122 ( .A(n9389), .B(n9229), .ZN(n9207) );
  NAND4_X1 U7123 ( .A1(n9183), .A2(n5615), .A3(n5614), .A4(n9207), .ZN(n5616)
         );
  NOR3_X1 U7124 ( .A1(n9147), .A2(n9167), .A3(n5616), .ZN(n5618) );
  NAND2_X1 U7125 ( .A1(n9080), .A2(n5617), .ZN(n5744) );
  NAND4_X1 U7126 ( .A1(n5750), .A2(n9131), .A3(n5618), .A4(n5744), .ZN(n5621)
         );
  INV_X1 U7127 ( .A(n5749), .ZN(n5620) );
  OAI21_X1 U7128 ( .B1(n5621), .B2(n5620), .A(n5619), .ZN(n5715) );
  AND2_X1 U7129 ( .A1(n5622), .A2(n5715), .ZN(n5716) );
  XNOR2_X2 U7130 ( .A(n5624), .B(n5753), .ZN(n5714) );
  AOI21_X1 U7131 ( .B1(n5625), .B2(n4562), .A(n5710), .ZN(n5702) );
  INV_X1 U7132 ( .A(n5626), .ZN(n9125) );
  NAND2_X1 U7133 ( .A1(n7067), .A2(n5630), .ZN(n5726) );
  NAND2_X1 U7134 ( .A1(n5726), .A2(n5631), .ZN(n7314) );
  AOI21_X1 U7135 ( .B1(n7314), .B2(n7313), .A(n5632), .ZN(n5634) );
  NOR2_X1 U7136 ( .A1(n5634), .A2(n5633), .ZN(n5635) );
  INV_X1 U7137 ( .A(n9484), .ZN(n5636) );
  OAI211_X1 U7138 ( .C1(n5639), .C2(n7637), .A(n5638), .B(n5637), .ZN(n5640)
         );
  AOI21_X1 U7139 ( .B1(n5640), .B2(n6701), .A(n7636), .ZN(n5650) );
  INV_X1 U7140 ( .A(n5641), .ZN(n5644) );
  OAI21_X1 U7141 ( .B1(n5644), .B2(n5643), .A(n5642), .ZN(n5645) );
  NAND2_X1 U7142 ( .A1(n5645), .A2(n7638), .ZN(n5646) );
  AOI22_X1 U7143 ( .A1(n5650), .A2(n5646), .B1(n4562), .B2(n7691), .ZN(n5653)
         );
  INV_X1 U7144 ( .A(n5647), .ZN(n5652) );
  NAND2_X1 U7145 ( .A1(n5648), .A2(n7693), .ZN(n5649) );
  OAI22_X1 U7146 ( .A1(n5650), .A2(n5649), .B1(n6701), .B2(n5654), .ZN(n5651)
         );
  OAI21_X1 U7147 ( .B1(n5653), .B2(n5652), .A(n5651), .ZN(n5659) );
  INV_X1 U7148 ( .A(n7752), .ZN(n5655) );
  NAND2_X1 U7149 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  MUX2_X1 U7150 ( .A(n5657), .B(n5656), .S(n6701), .Z(n5658) );
  MUX2_X1 U7151 ( .A(n5660), .B(n9107), .S(n6701), .Z(n5661) );
  MUX2_X1 U7152 ( .A(n9110), .B(n9111), .S(n6701), .Z(n5662) );
  INV_X1 U7153 ( .A(n9114), .ZN(n5663) );
  NOR2_X1 U7154 ( .A1(n5663), .A2(n9113), .ZN(n5665) );
  INV_X1 U7155 ( .A(n9115), .ZN(n5664) );
  MUX2_X1 U7156 ( .A(n5665), .B(n5664), .S(n6701), .Z(n5666) );
  NAND3_X1 U7157 ( .A1(n5676), .A2(n5667), .A3(n5677), .ZN(n5671) );
  INV_X1 U7158 ( .A(n9116), .ZN(n5668) );
  NOR2_X1 U7159 ( .A1(n9118), .A2(n5668), .ZN(n5670) );
  INV_X1 U7160 ( .A(n9117), .ZN(n5669) );
  AOI21_X1 U7161 ( .B1(n5671), .B2(n5670), .A(n5669), .ZN(n5673) );
  INV_X1 U7162 ( .A(n5672), .ZN(n9119) );
  OAI21_X1 U7163 ( .B1(n5673), .B2(n9119), .A(n5678), .ZN(n5675) );
  NAND3_X1 U7164 ( .A1(n5676), .A2(n9114), .A3(n9116), .ZN(n5679) );
  NAND4_X1 U7165 ( .A1(n5679), .A2(n5678), .A3(n9117), .A4(n5677), .ZN(n5682)
         );
  NAND3_X1 U7166 ( .A1(n5682), .A2(n5681), .A3(n5680), .ZN(n5684) );
  INV_X1 U7167 ( .A(n9124), .ZN(n5683) );
  NAND2_X1 U7168 ( .A1(n5684), .A2(n5683), .ZN(n5685) );
  INV_X1 U7169 ( .A(n9123), .ZN(n5686) );
  OAI21_X1 U7170 ( .B1(n5686), .B2(n9122), .A(n9180), .ZN(n5687) );
  MUX2_X1 U7171 ( .A(n5741), .B(n5687), .S(n6701), .Z(n5688) );
  INV_X1 U7172 ( .A(n9127), .ZN(n5720) );
  INV_X1 U7173 ( .A(n5689), .ZN(n5691) );
  AOI211_X1 U7174 ( .C1(n5694), .C2(n5720), .A(n5691), .B(n5690), .ZN(n5696)
         );
  INV_X1 U7175 ( .A(n5692), .ZN(n5693) );
  NOR2_X1 U7176 ( .A1(n5694), .A2(n5693), .ZN(n5695) );
  AOI21_X1 U7177 ( .B1(n5703), .B2(n5704), .A(n5697), .ZN(n5699) );
  OAI211_X1 U7178 ( .C1(n5699), .C2(n5698), .A(n9131), .B(n6701), .ZN(n5701)
         );
  NAND3_X1 U7179 ( .A1(n9361), .A2(n6701), .A3(n9155), .ZN(n5700) );
  OAI211_X1 U7180 ( .C1(n5707), .C2(n5702), .A(n5701), .B(n5700), .ZN(n5713)
         );
  INV_X1 U7181 ( .A(n9131), .ZN(n5706) );
  INV_X1 U7182 ( .A(n5709), .ZN(n5712) );
  AOI21_X1 U7183 ( .B1(n5710), .B2(n6701), .A(n5718), .ZN(n5711) );
  INV_X1 U7184 ( .A(n5714), .ZN(n5763) );
  NAND2_X1 U7185 ( .A1(n5763), .A2(n5762), .ZN(n6981) );
  NAND2_X1 U7186 ( .A1(n9102), .A2(n5720), .ZN(n5721) );
  NOR2_X1 U7187 ( .A1(n5722), .A2(n5721), .ZN(n5742) );
  INV_X1 U7188 ( .A(n5723), .ZN(n5724) );
  NOR2_X1 U7189 ( .A1(n5724), .A2(n9124), .ZN(n5740) );
  NAND2_X1 U7190 ( .A1(n5726), .A2(n5725), .ZN(n5728) );
  NAND2_X1 U7191 ( .A1(n5728), .A2(n5727), .ZN(n7418) );
  OAI21_X1 U7192 ( .B1(n6818), .B2(n7162), .A(n5762), .ZN(n5732) );
  INV_X1 U7193 ( .A(n5729), .ZN(n5730) );
  OAI21_X1 U7194 ( .B1(n6826), .B2(n7305), .A(n5730), .ZN(n5731) );
  NOR2_X1 U7195 ( .A1(n5732), .A2(n5731), .ZN(n5734) );
  AOI22_X1 U7196 ( .A1(n7418), .A2(n5735), .B1(n5734), .B2(n5733), .ZN(n5737)
         );
  OAI21_X1 U7197 ( .B1(n5738), .B2(n5737), .A(n5736), .ZN(n5739) );
  NAND4_X1 U7198 ( .A1(n5742), .A2(n5740), .A3(n9122), .A4(n5739), .ZN(n5747)
         );
  NAND2_X1 U7199 ( .A1(n5742), .A2(n5741), .ZN(n5746) );
  INV_X1 U7200 ( .A(n5743), .ZN(n5745) );
  NAND4_X1 U7201 ( .A1(n5745), .A2(n5746), .A3(n5747), .A4(n5744), .ZN(n5748)
         );
  NAND2_X1 U7202 ( .A1(n5749), .A2(n5748), .ZN(n5751) );
  NAND2_X1 U7203 ( .A1(n5751), .A2(n5750), .ZN(n5761) );
  INV_X1 U7204 ( .A(n6985), .ZN(n7205) );
  NAND3_X1 U7205 ( .A1(n5761), .A2(n9214), .A3(n7362), .ZN(n5760) );
  NAND3_X1 U7206 ( .A1(n5755), .A2(n5754), .A3(n5753), .ZN(n5756) );
  OAI21_X1 U7207 ( .B1(n5752), .B2(n5756), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5758) );
  XNOR2_X1 U7208 ( .A(n5758), .B(n5757), .ZN(n6319) );
  OR2_X1 U7209 ( .A1(n6319), .A2(P1_U3084), .ZN(n7543) );
  INV_X1 U7210 ( .A(n7543), .ZN(n5759) );
  OAI211_X1 U7211 ( .C1(n5761), .C2(n7205), .A(n5760), .B(n5759), .ZN(n5777)
         );
  NAND2_X1 U7212 ( .A1(n5763), .A2(n6978), .ZN(n6984) );
  INV_X1 U7213 ( .A(n6984), .ZN(n5764) );
  AND2_X1 U7214 ( .A1(n6784), .A2(n5764), .ZN(n7283) );
  INV_X1 U7215 ( .A(n4391), .ZN(n6854) );
  INV_X1 U7216 ( .A(n5766), .ZN(n9075) );
  NAND2_X1 U7217 ( .A1(n5770), .A2(n5769), .ZN(n5772) );
  OR2_X1 U7218 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  NAND2_X1 U7219 ( .A1(n5772), .A2(n5771), .ZN(n7739) );
  XNOR2_X1 U7220 ( .A(n5774), .B(n5773), .ZN(n7689) );
  AND2_X1 U7221 ( .A1(n6319), .A2(n6785), .ZN(n6838) );
  NAND4_X1 U7222 ( .A1(n7283), .A2(n6854), .A3(n9075), .A4(n6795), .ZN(n5775)
         );
  OAI211_X1 U7223 ( .C1(n5763), .C2(n7543), .A(n5775), .B(P1_B_REG_SCAN_IN), 
        .ZN(n5776) );
  NOR2_X1 U7224 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5780) );
  NOR2_X1 U7225 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5779) );
  NOR2_X1 U7226 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5778) );
  NAND4_X1 U7227 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5977), .ZN(n5785)
         );
  INV_X1 U7228 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5783) );
  INV_X1 U7229 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5782) );
  INV_X1 U7230 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5781) );
  NAND4_X1 U7231 ( .A1(n5958), .A2(n5783), .A3(n5782), .A4(n5781), .ZN(n5784)
         );
  NOR2_X1 U7232 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5788) );
  INV_X1 U7233 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6284) );
  INV_X1 U7234 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5787) );
  NAND4_X1 U7235 ( .A1(n5788), .A2(n6284), .A3(n5812), .A4(n5787), .ZN(n5791)
         );
  INV_X1 U7236 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5815) );
  INV_X1 U7237 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5789) );
  INV_X1 U7238 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6262) );
  NAND4_X1 U7239 ( .A1(n5815), .A2(n5789), .A3(n6262), .A4(n6266), .ZN(n5790)
         );
  NAND2_X1 U7240 ( .A1(n5817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5794) );
  INV_X1 U7241 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5793) );
  MUX2_X1 U7242 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5796), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5797) );
  INV_X1 U7243 ( .A(n6385), .ZN(n5798) );
  NAND2_X1 U7244 ( .A1(n5862), .A2(n5798), .ZN(n5805) );
  NAND2_X1 U7245 ( .A1(n4400), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5804) );
  INV_X2 U7246 ( .A(n6482), .ZN(n6424) );
  NAND2_X1 U7247 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n9691), .ZN(n5799) );
  MUX2_X1 U7248 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5799), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5802) );
  INV_X1 U7249 ( .A(n5800), .ZN(n5801) );
  NAND2_X1 U7250 ( .A1(n5802), .A2(n5801), .ZN(n6627) );
  INV_X1 U7251 ( .A(n6627), .ZN(n6448) );
  NAND2_X1 U7252 ( .A1(n6424), .A2(n6448), .ZN(n5803) );
  INV_X1 U7253 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5807) );
  NOR2_X1 U7254 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5808) );
  NAND2_X1 U7255 ( .A1(n5811), .A2(n5808), .ZN(n5809) );
  OAI21_X2 U7256 ( .B1(n5809), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6263) );
  INV_X1 U7257 ( .A(n8235), .ZN(n7509) );
  NAND2_X1 U7258 ( .A1(n5809), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5810) );
  INV_X1 U7259 ( .A(n8223), .ZN(n7384) );
  NAND2_X2 U7260 ( .A1(n7509), .A2(n7384), .ZN(n6293) );
  NAND2_X1 U7261 ( .A1(n8235), .A2(n4394), .ZN(n8219) );
  NAND2_X1 U7262 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  NAND2_X1 U7263 ( .A1(n5814), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5816) );
  XNOR2_X2 U7264 ( .A(n5816), .B(n5815), .ZN(n8226) );
  INV_X1 U7265 ( .A(n8226), .ZN(n6292) );
  NAND2_X1 U7266 ( .A1(n8223), .A2(n6292), .ZN(n8038) );
  XNOR2_X1 U7267 ( .A(n6892), .B(n4398), .ZN(n5829) );
  NAND2_X1 U7268 ( .A1(n5819), .A2(n5818), .ZN(n8756) );
  NAND2_X1 U7269 ( .A1(n5857), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7270 ( .A1(n4396), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5821) );
  AND2_X1 U7271 ( .A1(n5822), .A2(n5821), .ZN(n5827) );
  AND2_X4 U7272 ( .A1(n5823), .A2(n5824), .ZN(n6238) );
  NAND2_X1 U7273 ( .A1(n6238), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5826) );
  AND2_X4 U7274 ( .A1(n8240), .A2(n5824), .ZN(n6505) );
  NAND2_X1 U7275 ( .A1(n6505), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5825) );
  NAND3_X2 U7276 ( .A1(n5827), .A2(n5826), .A3(n5825), .ZN(n6891) );
  OR2_X2 U7277 ( .A1(n6293), .A2(n6305), .ZN(n8039) );
  NAND2_X1 U7278 ( .A1(n6891), .A2(n8039), .ZN(n5828) );
  NAND2_X1 U7279 ( .A1(n5829), .A2(n5828), .ZN(n5840) );
  NAND2_X1 U7280 ( .A1(n6238), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7281 ( .A1(n5857), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7282 ( .A1(n6505), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7283 ( .A1(n4396), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5831) );
  INV_X1 U7284 ( .A(SI_0_), .ZN(n5835) );
  OR2_X1 U7285 ( .A1(n6384), .A2(n5835), .ZN(n5837) );
  INV_X1 U7286 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5836) );
  XNOR2_X1 U7287 ( .A(n5837), .B(n5836), .ZN(n8772) );
  MUX2_X1 U7288 ( .A(n4617), .B(n8772), .S(n6482), .Z(n6760) );
  INV_X1 U7289 ( .A(n6760), .ZN(n7003) );
  NAND2_X1 U7290 ( .A1(n6649), .A2(n7003), .ZN(n7002) );
  NAND2_X1 U7291 ( .A1(n4390), .A2(n6760), .ZN(n5838) );
  AND2_X1 U7292 ( .A1(n5839), .A2(n5838), .ZN(n6738) );
  NAND2_X1 U7293 ( .A1(n6737), .A2(n5840), .ZN(n6730) );
  NAND2_X1 U7294 ( .A1(n6119), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5845) );
  INV_X1 U7295 ( .A(n6395), .ZN(n5841) );
  NAND2_X1 U7296 ( .A1(n5862), .A2(n5841), .ZN(n5844) );
  OR2_X1 U7297 ( .A1(n5800), .A2(n5795), .ZN(n5842) );
  XNOR2_X1 U7298 ( .A(n5842), .B(P2_IR_REG_2__SCAN_IN), .ZN(n8378) );
  NAND2_X1 U7299 ( .A1(n6424), .A2(n8378), .ZN(n5843) );
  XNOR2_X1 U7301 ( .A(n9779), .B(n5846), .ZN(n5852) );
  NAND2_X1 U7302 ( .A1(n6505), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U7303 ( .A1(n4396), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7304 ( .A1(n5857), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U7305 ( .A1(n6238), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5847) );
  NAND4_X2 U7306 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n8372)
         );
  NAND2_X1 U7307 ( .A1(n8372), .A2(n8039), .ZN(n5851) );
  XNOR2_X1 U7308 ( .A(n5852), .B(n5851), .ZN(n6731) );
  NAND2_X1 U7309 ( .A1(n6119), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7310 ( .A1(n5853), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5854) );
  XNOR2_X1 U7311 ( .A(n5854), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6535) );
  NAND2_X1 U7312 ( .A1(n6424), .A2(n6535), .ZN(n5855) );
  XNOR2_X1 U7313 ( .A(n5846), .B(n9806), .ZN(n5876) );
  NAND2_X1 U7314 ( .A1(n6238), .A2(n6901), .ZN(n5861) );
  NAND2_X1 U7315 ( .A1(n5857), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U7316 ( .A1(n6505), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7317 ( .A1(n4399), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7318 ( .A1(n9772), .A2(n8039), .ZN(n5875) );
  XNOR2_X1 U7319 ( .A(n5876), .B(n5875), .ZN(n6745) );
  INV_X1 U7320 ( .A(n6393), .ZN(n5863) );
  NAND2_X1 U7321 ( .A1(n5862), .A2(n5863), .ZN(n5868) );
  NAND2_X1 U7322 ( .A1(n6205), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7323 ( .A1(n5864), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5865) );
  XNOR2_X1 U7324 ( .A(n5865), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U7325 ( .A1(n4402), .A2(n6520), .ZN(n5866) );
  AND3_X2 U7326 ( .A1(n5868), .A2(n5867), .A3(n5866), .ZN(n9756) );
  XNOR2_X1 U7327 ( .A(n9756), .B(n5846), .ZN(n5879) );
  NAND2_X1 U7328 ( .A1(n5857), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5873) );
  NAND2_X1 U7329 ( .A1(n6505), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5872) );
  INV_X1 U7330 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5869) );
  XNOR2_X1 U7331 ( .A(n5869), .B(P2_REG3_REG_3__SCAN_IN), .ZN(n9749) );
  NAND2_X1 U7332 ( .A1(n6238), .A2(n9749), .ZN(n5871) );
  INV_X2 U7333 ( .A(n6213), .ZN(n6506) );
  NAND2_X1 U7334 ( .A1(n6506), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5870) );
  NAND4_X1 U7335 ( .A1(n5873), .A2(n5872), .A3(n5871), .A4(n5870), .ZN(n8371)
         );
  NAND2_X1 U7336 ( .A1(n8371), .A2(n8039), .ZN(n5878) );
  NAND2_X1 U7337 ( .A1(n5879), .A2(n5878), .ZN(n6669) );
  AND2_X1 U7338 ( .A1(n6745), .A2(n6669), .ZN(n5874) );
  INV_X1 U7339 ( .A(n6669), .ZN(n5881) );
  INV_X1 U7340 ( .A(n5875), .ZN(n5877) );
  NAND2_X1 U7341 ( .A1(n5877), .A2(n5876), .ZN(n6671) );
  OR2_X1 U7342 ( .A1(n5879), .A2(n5878), .ZN(n6670) );
  AND2_X1 U7343 ( .A1(n6671), .A2(n6670), .ZN(n5880) );
  NAND2_X1 U7344 ( .A1(n5883), .A2(n5882), .ZN(n6751) );
  INV_X1 U7345 ( .A(n6391), .ZN(n5884) );
  NAND2_X1 U7346 ( .A1(n5862), .A2(n5884), .ZN(n5893) );
  NAND2_X1 U7347 ( .A1(n6205), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5892) );
  NOR2_X1 U7348 ( .A1(n5887), .A2(n5795), .ZN(n5885) );
  MUX2_X1 U7349 ( .A(n5795), .B(n5885), .S(P2_IR_REG_5__SCAN_IN), .Z(n5889) );
  INV_X1 U7350 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5886) );
  NAND2_X1 U7351 ( .A1(n5887), .A2(n5886), .ZN(n5923) );
  INV_X1 U7352 ( .A(n5923), .ZN(n5888) );
  OR2_X1 U7353 ( .A1(n5889), .A2(n5888), .ZN(n6618) );
  INV_X1 U7354 ( .A(n6618), .ZN(n5890) );
  NAND2_X1 U7355 ( .A1(n6424), .A2(n5890), .ZN(n5891) );
  XNOR2_X1 U7356 ( .A(n9821), .B(n5846), .ZN(n5903) );
  NAND2_X1 U7357 ( .A1(n5857), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7358 ( .A1(n6505), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5899) );
  NAND3_X1 U7359 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5912) );
  INV_X1 U7360 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U7361 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5894) );
  NAND2_X1 U7362 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  AND2_X1 U7363 ( .A1(n5912), .A2(n5896), .ZN(n7038) );
  NAND2_X1 U7364 ( .A1(n6238), .A2(n7038), .ZN(n5898) );
  NAND2_X1 U7365 ( .A1(n4399), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5897) );
  NAND4_X1 U7366 ( .A1(n5900), .A2(n5899), .A3(n5898), .A4(n5897), .ZN(n8370)
         );
  AND2_X1 U7367 ( .A1(n8370), .A2(n8039), .ZN(n5901) );
  XNOR2_X1 U7368 ( .A(n5903), .B(n5901), .ZN(n6752) );
  NAND2_X1 U7369 ( .A1(n6751), .A2(n6752), .ZN(n5905) );
  INV_X1 U7370 ( .A(n5901), .ZN(n5902) );
  OR2_X1 U7371 ( .A1(n5903), .A2(n5902), .ZN(n5904) );
  INV_X1 U7372 ( .A(n6769), .ZN(n5921) );
  NAND2_X1 U7373 ( .A1(n5923), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5907) );
  XNOR2_X1 U7374 ( .A(n5907), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6584) );
  INV_X1 U7375 ( .A(n6584), .ZN(n6397) );
  NAND2_X1 U7376 ( .A1(n6205), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5908) );
  XNOR2_X1 U7377 ( .A(n5906), .B(n7115), .ZN(n5919) );
  NAND2_X1 U7378 ( .A1(n4399), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7379 ( .A1(n8025), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5916) );
  INV_X1 U7380 ( .A(n5912), .ZN(n5911) );
  NAND2_X1 U7381 ( .A1(n5911), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5929) );
  INV_X1 U7382 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9934) );
  NAND2_X1 U7383 ( .A1(n5912), .A2(n9934), .ZN(n5913) );
  AND2_X1 U7384 ( .A1(n5929), .A2(n5913), .ZN(n8628) );
  NAND2_X1 U7385 ( .A1(n6238), .A2(n8628), .ZN(n5915) );
  NAND2_X1 U7386 ( .A1(n6505), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5914) );
  OR2_X1 U7387 ( .A1(n7117), .A2(n6759), .ZN(n5918) );
  NAND2_X1 U7388 ( .A1(n5919), .A2(n5918), .ZN(n5922) );
  OAI21_X1 U7389 ( .B1(n5919), .B2(n5918), .A(n5922), .ZN(n6770) );
  INV_X1 U7390 ( .A(n6770), .ZN(n5920) );
  NAND2_X1 U7391 ( .A1(n6400), .A2(n5862), .ZN(n5926) );
  NAND2_X1 U7392 ( .A1(n5942), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5924) );
  XNOR2_X1 U7393 ( .A(n5924), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6549) );
  AOI22_X1 U7394 ( .A1(n6205), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n4402), .B2(
        n6549), .ZN(n5925) );
  NAND2_X1 U7395 ( .A1(n5926), .A2(n5925), .ZN(n9727) );
  XNOR2_X1 U7396 ( .A(n9727), .B(n5906), .ZN(n5936) );
  NAND2_X1 U7397 ( .A1(n6506), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7398 ( .A1(n8025), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5933) );
  INV_X1 U7399 ( .A(n5929), .ZN(n5927) );
  NAND2_X1 U7400 ( .A1(n5927), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5948) );
  INV_X1 U7401 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7402 ( .A1(n5929), .A2(n5928), .ZN(n5930) );
  AND2_X1 U7403 ( .A1(n5948), .A2(n5930), .ZN(n9725) );
  NAND2_X1 U7404 ( .A1(n6238), .A2(n9725), .ZN(n5932) );
  NAND2_X1 U7405 ( .A1(n6505), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5931) );
  NAND4_X1 U7406 ( .A1(n5934), .A2(n5933), .A3(n5932), .A4(n5931), .ZN(n8368)
         );
  NAND2_X1 U7407 ( .A1(n8368), .A2(n8039), .ZN(n5937) );
  XNOR2_X1 U7408 ( .A(n5936), .B(n5937), .ZN(n6941) );
  INV_X1 U7409 ( .A(n6941), .ZN(n5935) );
  INV_X1 U7410 ( .A(n5936), .ZN(n5939) );
  INV_X1 U7411 ( .A(n5937), .ZN(n5938) );
  NAND2_X1 U7412 ( .A1(n5939), .A2(n5938), .ZN(n5940) );
  NAND2_X1 U7413 ( .A1(n6409), .A2(n6204), .ZN(n5945) );
  NOR2_X1 U7414 ( .A1(n5942), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5959) );
  OR2_X1 U7415 ( .A1(n5959), .A2(n5795), .ZN(n5943) );
  XNOR2_X1 U7416 ( .A(n5943), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9694) );
  AOI22_X1 U7417 ( .A1(n6205), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6424), .B2(
        n9694), .ZN(n5944) );
  NAND2_X1 U7418 ( .A1(n5945), .A2(n5944), .ZN(n7226) );
  XNOR2_X1 U7419 ( .A(n7226), .B(n5906), .ZN(n5954) );
  NAND2_X1 U7420 ( .A1(n6506), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7421 ( .A1(n8025), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5952) );
  INV_X1 U7422 ( .A(n5948), .ZN(n5946) );
  NAND2_X1 U7423 ( .A1(n5946), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5963) );
  INV_X1 U7424 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U7425 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  AND2_X1 U7426 ( .A1(n5963), .A2(n5949), .ZN(n7125) );
  NAND2_X1 U7427 ( .A1(n6238), .A2(n7125), .ZN(n5951) );
  NAND2_X1 U7428 ( .A1(n6505), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5950) );
  NOR2_X1 U7429 ( .A1(n7225), .A2(n6759), .ZN(n5955) );
  XNOR2_X1 U7430 ( .A(n5954), .B(n5955), .ZN(n6926) );
  INV_X1 U7431 ( .A(n5954), .ZN(n5956) );
  NAND2_X1 U7432 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  NAND2_X1 U7433 ( .A1(n6414), .A2(n6204), .ZN(n5961) );
  NAND2_X1 U7434 ( .A1(n5959), .A2(n5958), .ZN(n6009) );
  NAND2_X1 U7435 ( .A1(n6009), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5975) );
  XNOR2_X1 U7436 ( .A(n5975), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6561) );
  AOI22_X1 U7437 ( .A1(n6205), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6424), .B2(
        n6561), .ZN(n5960) );
  NAND2_X1 U7438 ( .A1(n5961), .A2(n5960), .ZN(n7346) );
  XNOR2_X1 U7439 ( .A(n7346), .B(n5906), .ZN(n5969) );
  NAND2_X1 U7440 ( .A1(n6506), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7441 ( .A1(n8025), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5967) );
  INV_X1 U7442 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7443 ( .A1(n5963), .A2(n5962), .ZN(n5964) );
  AND2_X1 U7444 ( .A1(n5983), .A2(n5964), .ZN(n7243) );
  NAND2_X1 U7445 ( .A1(n6238), .A2(n7243), .ZN(n5966) );
  NAND2_X1 U7446 ( .A1(n6505), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5965) );
  OR2_X1 U7447 ( .A1(n7224), .A2(n6759), .ZN(n5970) );
  NAND2_X1 U7448 ( .A1(n5969), .A2(n5970), .ZN(n5974) );
  INV_X1 U7449 ( .A(n5969), .ZN(n5972) );
  INV_X1 U7450 ( .A(n5970), .ZN(n5971) );
  NAND2_X1 U7451 ( .A1(n5972), .A2(n5971), .ZN(n5973) );
  NAND2_X1 U7452 ( .A1(n5974), .A2(n5973), .ZN(n7095) );
  NAND2_X1 U7453 ( .A1(n7093), .A2(n5974), .ZN(n7103) );
  NAND2_X1 U7454 ( .A1(n6418), .A2(n6204), .ZN(n5981) );
  INV_X1 U7455 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7456 ( .A1(n5975), .A2(n6006), .ZN(n5976) );
  NAND2_X1 U7457 ( .A1(n5976), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5978) );
  NAND2_X1 U7458 ( .A1(n5978), .A2(n5977), .ZN(n5993) );
  OR2_X1 U7459 ( .A1(n5978), .A2(n5977), .ZN(n5979) );
  NAND2_X1 U7460 ( .A1(n5993), .A2(n5979), .ZN(n6480) );
  INV_X1 U7461 ( .A(n6480), .ZN(n9708) );
  AOI22_X1 U7462 ( .A1(n6205), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4402), .B2(
        n9708), .ZN(n5980) );
  NAND2_X1 U7463 ( .A1(n5981), .A2(n5980), .ZN(n7451) );
  XNOR2_X1 U7464 ( .A(n7451), .B(n5846), .ZN(n5989) );
  NAND2_X1 U7465 ( .A1(n8025), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7466 ( .A1(n6505), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5987) );
  INV_X1 U7467 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7468 ( .A1(n5983), .A2(n5982), .ZN(n5984) );
  AND2_X1 U7469 ( .A1(n6017), .A2(n5984), .ZN(n7354) );
  NAND2_X1 U7470 ( .A1(n6238), .A2(n7354), .ZN(n5986) );
  NAND2_X1 U7471 ( .A1(n6506), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5985) );
  NOR2_X1 U7472 ( .A1(n7446), .A2(n6759), .ZN(n5990) );
  XNOR2_X1 U7473 ( .A(n5989), .B(n5990), .ZN(n7102) );
  INV_X1 U7474 ( .A(n5989), .ZN(n5992) );
  INV_X1 U7475 ( .A(n5990), .ZN(n5991) );
  OAI22_X2 U7476 ( .A1(n7103), .A2(n7102), .B1(n5992), .B2(n5991), .ZN(n7216)
         );
  NAND2_X1 U7477 ( .A1(n6428), .A2(n6204), .ZN(n5996) );
  NAND2_X1 U7478 ( .A1(n5993), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5994) );
  XNOR2_X1 U7479 ( .A(n5994), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6681) );
  AOI22_X1 U7480 ( .A1(n6205), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6681), .B2(
        n4402), .ZN(n5995) );
  XNOR2_X1 U7481 ( .A(n7450), .B(n5906), .ZN(n6003) );
  NAND2_X1 U7482 ( .A1(n6506), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7483 ( .A1(n8025), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5999) );
  XNOR2_X1 U7484 ( .A(n6017), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n7447) );
  NAND2_X1 U7485 ( .A1(n6238), .A2(n7447), .ZN(n5998) );
  NAND2_X1 U7486 ( .A1(n6505), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5997) );
  NAND4_X1 U7487 ( .A1(n6000), .A2(n5999), .A3(n5998), .A4(n5997), .ZN(n8364)
         );
  NAND2_X1 U7488 ( .A1(n8364), .A2(n8039), .ZN(n6001) );
  XNOR2_X1 U7489 ( .A(n6003), .B(n6001), .ZN(n7215) );
  NAND2_X1 U7490 ( .A1(n7216), .A2(n7215), .ZN(n6005) );
  INV_X1 U7491 ( .A(n6001), .ZN(n6002) );
  NAND2_X1 U7492 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  NAND2_X1 U7493 ( .A1(n6005), .A2(n6004), .ZN(n7408) );
  NAND2_X1 U7494 ( .A1(n6641), .A2(n6204), .ZN(n6012) );
  INV_X1 U7495 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7496 ( .A1(n6007), .A2(n6006), .ZN(n6008) );
  NAND2_X1 U7497 ( .A1(n6029), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6010) );
  XNOR2_X1 U7498 ( .A(n6010), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8394) );
  AOI22_X1 U7499 ( .A1(n6205), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6424), .B2(
        n8394), .ZN(n6011) );
  XNOR2_X1 U7500 ( .A(n7559), .B(n5906), .ZN(n6023) );
  NAND2_X1 U7501 ( .A1(n6506), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U7502 ( .A1(n5857), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6021) );
  AND2_X1 U7503 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_REG3_REG_11__SCAN_IN), 
        .ZN(n6013) );
  INV_X1 U7504 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n6016) );
  INV_X1 U7505 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6015) );
  OAI21_X1 U7506 ( .B1(n6017), .B2(n6016), .A(n6015), .ZN(n6018) );
  AND2_X1 U7507 ( .A1(n6033), .A2(n6018), .ZN(n7469) );
  NAND2_X1 U7508 ( .A1(n6238), .A2(n7469), .ZN(n6020) );
  NAND2_X1 U7509 ( .A1(n6505), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6019) );
  OR2_X1 U7510 ( .A1(n7461), .A2(n6759), .ZN(n6024) );
  NAND2_X1 U7511 ( .A1(n6023), .A2(n6024), .ZN(n6028) );
  INV_X1 U7512 ( .A(n6023), .ZN(n6026) );
  INV_X1 U7513 ( .A(n6024), .ZN(n6025) );
  NAND2_X1 U7514 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  NAND2_X1 U7515 ( .A1(n6028), .A2(n6027), .ZN(n7407) );
  OR2_X2 U7516 ( .A1(n7408), .A2(n7407), .ZN(n7405) );
  NAND2_X1 U7517 ( .A1(n6656), .A2(n5862), .ZN(n6031) );
  OAI21_X1 U7518 ( .B1(n6029), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6043) );
  XNOR2_X1 U7519 ( .A(n6043), .B(P2_IR_REG_13__SCAN_IN), .ZN(n6697) );
  AOI22_X1 U7520 ( .A1(n6205), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6424), .B2(
        n6697), .ZN(n6030) );
  XNOR2_X1 U7521 ( .A(n7602), .B(n5846), .ZN(n6040) );
  INV_X1 U7522 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7438) );
  NAND2_X1 U7523 ( .A1(n6033), .A2(n7438), .ZN(n6034) );
  AND2_X1 U7524 ( .A1(n6048), .A2(n6034), .ZN(n7566) );
  NAND2_X1 U7525 ( .A1(n6238), .A2(n7566), .ZN(n6038) );
  NAND2_X1 U7526 ( .A1(n5857), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7527 ( .A1(n6505), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7528 ( .A1(n6506), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6035) );
  NOR2_X1 U7529 ( .A1(n7596), .A2(n6759), .ZN(n6039) );
  XNOR2_X1 U7530 ( .A(n6040), .B(n6039), .ZN(n7434) );
  NAND2_X1 U7531 ( .A1(n6662), .A2(n6204), .ZN(n6046) );
  INV_X1 U7532 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6042) );
  NAND2_X1 U7533 ( .A1(n6043), .A2(n6042), .ZN(n6044) );
  NAND2_X1 U7534 ( .A1(n6044), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6061) );
  XNOR2_X1 U7535 ( .A(n6061), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7046) );
  AOI22_X1 U7536 ( .A1(n7046), .A2(n4402), .B1(n6205), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6045) );
  XNOR2_X1 U7537 ( .A(n7671), .B(n5906), .ZN(n6054) );
  NAND2_X1 U7538 ( .A1(n6506), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7539 ( .A1(n8025), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6052) );
  INV_X1 U7540 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7541 ( .A1(n6048), .A2(n6047), .ZN(n6049) );
  AND2_X1 U7542 ( .A1(n6067), .A2(n6049), .ZN(n7597) );
  NAND2_X1 U7543 ( .A1(n6238), .A2(n7597), .ZN(n6051) );
  NAND2_X1 U7544 ( .A1(n6505), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6050) );
  OR2_X1 U7545 ( .A1(n7670), .A2(n6759), .ZN(n6055) );
  NAND2_X1 U7546 ( .A1(n6054), .A2(n6055), .ZN(n6059) );
  INV_X1 U7547 ( .A(n6054), .ZN(n6057) );
  INV_X1 U7548 ( .A(n6055), .ZN(n6056) );
  NAND2_X1 U7549 ( .A1(n6057), .A2(n6056), .ZN(n6058) );
  AND2_X1 U7550 ( .A1(n6059), .A2(n6058), .ZN(n7593) );
  NAND2_X1 U7551 ( .A1(n7591), .A2(n6059), .ZN(n7623) );
  NAND2_X1 U7552 ( .A1(n6743), .A2(n6204), .ZN(n6065) );
  INV_X1 U7553 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7554 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  NAND2_X1 U7555 ( .A1(n6062), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6063) );
  XNOR2_X1 U7556 ( .A(n6063), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7174) );
  AOI22_X1 U7557 ( .A1(n7174), .A2(n6424), .B1(n6205), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6064) );
  XNOR2_X1 U7558 ( .A(n8141), .B(n5906), .ZN(n6073) );
  NAND2_X1 U7559 ( .A1(n5857), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7560 ( .A1(n6505), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6071) );
  INV_X1 U7561 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7626) );
  NAND2_X1 U7562 ( .A1(n6067), .A2(n7626), .ZN(n6068) );
  AND2_X1 U7563 ( .A1(n6081), .A2(n6068), .ZN(n7680) );
  NAND2_X1 U7564 ( .A1(n6238), .A2(n7680), .ZN(n6070) );
  NAND2_X1 U7565 ( .A1(n6506), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6069) );
  NAND4_X1 U7566 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .ZN(n8360)
         );
  AND2_X1 U7567 ( .A1(n8360), .A2(n8039), .ZN(n7620) );
  INV_X1 U7568 ( .A(n6073), .ZN(n7621) );
  NAND2_X1 U7569 ( .A1(n6932), .A2(n6204), .ZN(n6079) );
  NOR2_X1 U7570 ( .A1(n5806), .A2(n5795), .ZN(n6074) );
  MUX2_X1 U7571 ( .A(n5795), .B(n6074), .S(P2_IR_REG_16__SCAN_IN), .Z(n6077)
         );
  INV_X1 U7572 ( .A(n6075), .ZN(n6076) );
  OR2_X1 U7573 ( .A1(n6077), .A2(n6076), .ZN(n7337) );
  INV_X1 U7574 ( .A(n7337), .ZN(n7178) );
  AOI22_X1 U7575 ( .A1(n6205), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4402), .B2(
        n7178), .ZN(n6078) );
  XNOR2_X1 U7576 ( .A(n7798), .B(n5906), .ZN(n6087) );
  NAND2_X1 U7577 ( .A1(n4399), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7578 ( .A1(n8025), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6085) );
  INV_X1 U7579 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7580 ( .A1(n6081), .A2(n6080), .ZN(n6082) );
  AND2_X1 U7581 ( .A1(n6098), .A2(n6082), .ZN(n7792) );
  NAND2_X1 U7582 ( .A1(n6238), .A2(n7792), .ZN(n6084) );
  NAND2_X1 U7583 ( .A1(n6505), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6083) );
  OR2_X1 U7584 ( .A1(n8359), .A2(n6759), .ZN(n6088) );
  NAND2_X1 U7585 ( .A1(n6087), .A2(n6088), .ZN(n6092) );
  INV_X1 U7586 ( .A(n6087), .ZN(n6090) );
  INV_X1 U7587 ( .A(n6088), .ZN(n6089) );
  NAND2_X1 U7588 ( .A1(n6090), .A2(n6089), .ZN(n6091) );
  NAND2_X1 U7589 ( .A1(n6092), .A2(n6091), .ZN(n7791) );
  NAND2_X1 U7590 ( .A1(n6911), .A2(n6204), .ZN(n6095) );
  NAND2_X1 U7591 ( .A1(n6075), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6093) );
  XNOR2_X1 U7592 ( .A(n6093), .B(n4647), .ZN(n7580) );
  INV_X1 U7593 ( .A(n7580), .ZN(n7335) );
  AOI22_X1 U7594 ( .A1(n6205), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6424), .B2(
        n7335), .ZN(n6094) );
  XNOR2_X1 U7595 ( .A(n8706), .B(n5906), .ZN(n6105) );
  NAND2_X1 U7596 ( .A1(n6506), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7597 ( .A1(n5857), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6102) );
  INV_X1 U7598 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7599 ( .A1(n6098), .A2(n6097), .ZN(n6099) );
  AND2_X1 U7600 ( .A1(n6110), .A2(n6099), .ZN(n8623) );
  NAND2_X1 U7601 ( .A1(n6238), .A2(n8623), .ZN(n6101) );
  NAND2_X1 U7602 ( .A1(n6505), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6100) );
  NAND4_X1 U7603 ( .A1(n6103), .A2(n6102), .A3(n6101), .A4(n6100), .ZN(n8358)
         );
  NAND2_X1 U7604 ( .A1(n8358), .A2(n8039), .ZN(n6104) );
  XNOR2_X1 U7605 ( .A(n6105), .B(n6104), .ZN(n7812) );
  NAND2_X1 U7606 ( .A1(n7077), .A2(n6204), .ZN(n6109) );
  NAND2_X1 U7607 ( .A1(n6106), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6107) );
  XNOR2_X1 U7608 ( .A(n6107), .B(P2_IR_REG_18__SCAN_IN), .ZN(n7588) );
  AOI22_X1 U7609 ( .A1(n6205), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6424), .B2(
        n7588), .ZN(n6108) );
  XNOR2_X1 U7610 ( .A(n8604), .B(n5906), .ZN(n6116) );
  INV_X1 U7611 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U7612 ( .A1(n6110), .A2(n7830), .ZN(n6111) );
  AND2_X1 U7613 ( .A1(n6123), .A2(n6111), .ZN(n8605) );
  NAND2_X1 U7614 ( .A1(n8605), .A2(n6238), .ZN(n6115) );
  NAND2_X1 U7615 ( .A1(n8025), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7616 ( .A1(n6505), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7617 ( .A1(n6506), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6112) );
  NOR2_X1 U7618 ( .A1(n8591), .A2(n6759), .ZN(n6117) );
  XNOR2_X1 U7619 ( .A(n6116), .B(n6117), .ZN(n7828) );
  INV_X1 U7620 ( .A(n6116), .ZN(n6118) );
  NAND2_X1 U7621 ( .A1(n7186), .A2(n6204), .ZN(n6121) );
  AOI22_X1 U7622 ( .A1(n6205), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4402), .B2(
        n4394), .ZN(n6120) );
  XNOR2_X1 U7623 ( .A(n8696), .B(n5906), .ZN(n6128) );
  INV_X1 U7624 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U7625 ( .A1(n6123), .A2(n9965), .ZN(n6124) );
  NAND2_X1 U7626 ( .A1(n6137), .A2(n6124), .ZN(n8582) );
  OR2_X1 U7627 ( .A1(n8582), .A2(n6295), .ZN(n6127) );
  AOI22_X1 U7628 ( .A1(n8025), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n4399), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7629 ( .A1(n6505), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6125) );
  OR2_X1 U7630 ( .A1(n8602), .A2(n6759), .ZN(n6129) );
  NAND2_X1 U7631 ( .A1(n6128), .A2(n6129), .ZN(n6133) );
  INV_X1 U7632 ( .A(n6128), .ZN(n6131) );
  INV_X1 U7633 ( .A(n6129), .ZN(n6130) );
  NAND2_X1 U7634 ( .A1(n6131), .A2(n6130), .ZN(n6132) );
  NAND2_X1 U7635 ( .A1(n6133), .A2(n6132), .ZN(n8287) );
  NAND2_X2 U7636 ( .A1(n8285), .A2(n6133), .ZN(n8319) );
  NAND2_X1 U7637 ( .A1(n7359), .A2(n6204), .ZN(n6135) );
  NAND2_X1 U7638 ( .A1(n6205), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6134) );
  XNOR2_X1 U7639 ( .A(n8689), .B(n5846), .ZN(n6156) );
  INV_X1 U7640 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U7641 ( .A1(n6137), .A2(n8320), .ZN(n6138) );
  NAND2_X1 U7642 ( .A1(n6144), .A2(n6138), .ZN(n8573) );
  OR2_X1 U7643 ( .A1(n8573), .A2(n6295), .ZN(n6141) );
  AOI22_X1 U7644 ( .A1(n5857), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n4399), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7645 ( .A1(n6505), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6139) );
  NOR2_X1 U7646 ( .A1(n8592), .A2(n6759), .ZN(n6155) );
  XNOR2_X1 U7647 ( .A(n6156), .B(n6155), .ZN(n8318) );
  NAND2_X1 U7648 ( .A1(n7383), .A2(n6204), .ZN(n6143) );
  NAND2_X1 U7649 ( .A1(n6119), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6142) );
  XNOR2_X1 U7650 ( .A(n8559), .B(n5846), .ZN(n6153) );
  INV_X1 U7651 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U7652 ( .A1(n6144), .A2(n8297), .ZN(n6145) );
  NAND2_X1 U7653 ( .A1(n6164), .A2(n6145), .ZN(n8557) );
  OR2_X1 U7654 ( .A1(n8557), .A2(n6295), .ZN(n6150) );
  INV_X1 U7655 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n10178) );
  INV_X1 U7656 ( .A(n6505), .ZN(n8028) );
  NAND2_X1 U7657 ( .A1(n6506), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7658 ( .A1(n8025), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6146) );
  OAI211_X1 U7659 ( .C1(n10178), .C2(n8028), .A(n6147), .B(n6146), .ZN(n6148)
         );
  INV_X1 U7660 ( .A(n6148), .ZN(n6149) );
  NAND2_X1 U7661 ( .A1(n6150), .A2(n6149), .ZN(n8567) );
  NAND2_X1 U7662 ( .A1(n8567), .A2(n8039), .ZN(n6152) );
  INV_X1 U7663 ( .A(n6152), .ZN(n6151) );
  NAND2_X1 U7664 ( .A1(n6153), .A2(n6151), .ZN(n6157) );
  INV_X1 U7665 ( .A(n6157), .ZN(n6154) );
  XNOR2_X1 U7666 ( .A(n6153), .B(n6152), .ZN(n8295) );
  NAND2_X1 U7667 ( .A1(n6156), .A2(n6155), .ZN(n8293) );
  AND2_X1 U7668 ( .A1(n8293), .A2(n6157), .ZN(n6158) );
  OAI21_X4 U7669 ( .B1(n8319), .B2(n6161), .A(n6160), .ZN(n6178) );
  NAND2_X1 U7670 ( .A1(n7508), .A2(n6204), .ZN(n6163) );
  NAND2_X1 U7671 ( .A1(n6119), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6162) );
  XNOR2_X1 U7672 ( .A(n8537), .B(n5846), .ZN(n6171) );
  INV_X1 U7673 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8328) );
  NAND2_X1 U7674 ( .A1(n6164), .A2(n8328), .ZN(n6165) );
  AND2_X1 U7675 ( .A1(n6181), .A2(n6165), .ZN(n8538) );
  NAND2_X1 U7676 ( .A1(n8538), .A2(n6238), .ZN(n6170) );
  INV_X1 U7677 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9913) );
  NAND2_X1 U7678 ( .A1(n8025), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7679 ( .A1(n6506), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6166) );
  OAI211_X1 U7680 ( .C1(n8028), .C2(n9913), .A(n6167), .B(n6166), .ZN(n6168)
         );
  INV_X1 U7681 ( .A(n6168), .ZN(n6169) );
  NOR2_X1 U7682 ( .A1(n8551), .A2(n6759), .ZN(n8326) );
  NOR2_X1 U7683 ( .A1(n6178), .A2(n6171), .ZN(n6175) );
  NAND2_X1 U7684 ( .A1(n7542), .A2(n6204), .ZN(n6173) );
  NAND2_X1 U7685 ( .A1(n6205), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6172) );
  XNOR2_X1 U7686 ( .A(n8525), .B(n5846), .ZN(n6174) );
  MUX2_X1 U7687 ( .A(n5846), .B(n8739), .S(n8326), .Z(n6176) );
  MUX2_X1 U7688 ( .A(n8537), .B(n5846), .S(n8326), .Z(n6177) );
  XNOR2_X1 U7689 ( .A(n6177), .B(n8674), .ZN(n6179) );
  INV_X1 U7690 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8280) );
  NAND2_X1 U7691 ( .A1(n6181), .A2(n8280), .ZN(n6182) );
  NAND2_X1 U7692 ( .A1(n6195), .A2(n6182), .ZN(n8521) );
  OR2_X1 U7693 ( .A1(n8521), .A2(n6295), .ZN(n6188) );
  INV_X1 U7694 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7695 ( .A1(n4399), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U7696 ( .A1(n5857), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6183) );
  OAI211_X1 U7697 ( .C1(n6185), .C2(n8028), .A(n6184), .B(n6183), .ZN(n6186)
         );
  INV_X1 U7698 ( .A(n6186), .ZN(n6187) );
  NOR2_X1 U7699 ( .A1(n8535), .A2(n6759), .ZN(n8278) );
  INV_X1 U7700 ( .A(n8278), .ZN(n6189) );
  OAI22_X2 U7701 ( .A1(n8325), .A2(n6190), .B1(n8279), .B2(n6189), .ZN(n6202)
         );
  NAND2_X1 U7702 ( .A1(n7686), .A2(n6204), .ZN(n6192) );
  NAND2_X1 U7703 ( .A1(n6119), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6191) );
  XNOR2_X1 U7704 ( .A(n8505), .B(n5846), .ZN(n6203) );
  INV_X1 U7705 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8313) );
  NAND2_X1 U7706 ( .A1(n6195), .A2(n8313), .ZN(n6196) );
  NAND2_X1 U7707 ( .A1(n6208), .A2(n6196), .ZN(n8503) );
  OR2_X1 U7708 ( .A1(n8503), .A2(n6295), .ZN(n6201) );
  INV_X1 U7709 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10180) );
  NAND2_X1 U7710 ( .A1(n6506), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7711 ( .A1(n8025), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6197) );
  OAI211_X1 U7712 ( .C1(n10180), .C2(n8028), .A(n6198), .B(n6197), .ZN(n6199)
         );
  INV_X1 U7713 ( .A(n6199), .ZN(n6200) );
  NOR2_X1 U7714 ( .A1(n8518), .A2(n6759), .ZN(n8312) );
  NAND2_X1 U7715 ( .A1(n7738), .A2(n6204), .ZN(n6207) );
  NAND2_X1 U7716 ( .A1(n6119), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6206) );
  XOR2_X1 U7717 ( .A(n5846), .B(n8664), .Z(n8303) );
  INV_X1 U7718 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9935) );
  NAND2_X1 U7719 ( .A1(n6208), .A2(n9935), .ZN(n6209) );
  AND2_X1 U7720 ( .A1(n6219), .A2(n6209), .ZN(n8306) );
  INV_X1 U7721 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U7722 ( .A1(n6505), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7723 ( .A1(n8025), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6210) );
  OAI211_X1 U7724 ( .C1(n6213), .C2(n6212), .A(n6211), .B(n6210), .ZN(n6214)
         );
  AOI21_X1 U7725 ( .B1(n8306), .B2(n6238), .A(n6214), .ZN(n8501) );
  INV_X1 U7726 ( .A(n8501), .ZN(n8355) );
  NAND2_X1 U7727 ( .A1(n8355), .A2(n8039), .ZN(n8302) );
  NAND2_X1 U7728 ( .A1(n7819), .A2(n6204), .ZN(n6216) );
  NAND2_X1 U7729 ( .A1(n6119), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6215) );
  XNOR2_X1 U7730 ( .A(n8477), .B(n5846), .ZN(n6227) );
  INV_X1 U7731 ( .A(n6219), .ZN(n6217) );
  NAND2_X1 U7732 ( .A1(n6217), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6232) );
  INV_X1 U7733 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7734 ( .A1(n6219), .A2(n6218), .ZN(n6220) );
  NAND2_X1 U7735 ( .A1(n6232), .A2(n6220), .ZN(n8474) );
  OR2_X1 U7736 ( .A1(n8474), .A2(n6295), .ZN(n6225) );
  INV_X1 U7737 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U7738 ( .A1(n4399), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7739 ( .A1(n8025), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6221) );
  OAI211_X1 U7740 ( .C1(n8660), .C2(n8028), .A(n6222), .B(n6221), .ZN(n6223)
         );
  INV_X1 U7741 ( .A(n6223), .ZN(n6224) );
  NOR2_X1 U7742 ( .A1(n8487), .A2(n6759), .ZN(n6226) );
  NAND2_X1 U7743 ( .A1(n6227), .A2(n6226), .ZN(n6228) );
  OAI21_X1 U7744 ( .B1(n6227), .B2(n6226), .A(n6228), .ZN(n8342) );
  NAND2_X1 U7745 ( .A1(n6119), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6229) );
  XNOR2_X1 U7746 ( .A(n8652), .B(n5846), .ZN(n6240) );
  INV_X1 U7747 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6231) );
  NAND2_X1 U7748 ( .A1(n6232), .A2(n6231), .ZN(n6233) );
  INV_X1 U7749 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6236) );
  NAND2_X1 U7750 ( .A1(n5857), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U7751 ( .A1(n4399), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6234) );
  OAI211_X1 U7752 ( .C1(n6236), .C2(n8028), .A(n6235), .B(n6234), .ZN(n6237)
         );
  NOR2_X1 U7753 ( .A1(n8471), .A2(n6759), .ZN(n6239) );
  NAND2_X1 U7754 ( .A1(n6240), .A2(n6239), .ZN(n6289) );
  OAI21_X1 U7755 ( .B1(n6240), .B2(n6239), .A(n6289), .ZN(n8270) );
  NOR2_X1 U7756 ( .A1(n8271), .A2(n8270), .ZN(n6288) );
  INV_X1 U7757 ( .A(n6288), .ZN(n8273) );
  NAND2_X1 U7758 ( .A1(n6119), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6241) );
  INV_X1 U7759 ( .A(n6244), .ZN(n6243) );
  NAND2_X1 U7760 ( .A1(n6243), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8252) );
  INV_X1 U7761 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6303) );
  NAND2_X1 U7762 ( .A1(n6244), .A2(n6303), .ZN(n6245) );
  NAND2_X1 U7763 ( .A1(n8252), .A2(n6245), .ZN(n8443) );
  INV_X1 U7764 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n10132) );
  NAND2_X1 U7765 ( .A1(n8025), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7766 ( .A1(n6506), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6246) );
  OAI211_X1 U7767 ( .C1(n10132), .C2(n8028), .A(n6247), .B(n6246), .ZN(n6248)
         );
  INV_X1 U7768 ( .A(n6248), .ZN(n6249) );
  NOR2_X1 U7769 ( .A1(n8249), .A2(n6759), .ZN(n6251) );
  XNOR2_X1 U7770 ( .A(n6251), .B(n5846), .ZN(n6252) );
  XNOR2_X1 U7771 ( .A(n8442), .B(n6252), .ZN(n6290) );
  INV_X1 U7772 ( .A(n6290), .ZN(n6287) );
  NOR4_X1 U7773 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6261) );
  NOR4_X1 U7774 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6260) );
  INV_X1 U7775 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9980) );
  INV_X1 U7776 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9951) );
  INV_X1 U7777 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9979) );
  INV_X1 U7778 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9937) );
  NAND4_X1 U7779 ( .A1(n9980), .A2(n9951), .A3(n9979), .A4(n9937), .ZN(n6258)
         );
  NOR4_X1 U7780 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6256) );
  NOR4_X1 U7781 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6255) );
  NOR4_X1 U7782 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6254) );
  NOR4_X1 U7783 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6253) );
  NAND4_X1 U7784 ( .A1(n6256), .A2(n6255), .A3(n6254), .A4(n6253), .ZN(n6257)
         );
  NOR4_X1 U7785 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        n6258), .A4(n6257), .ZN(n6259) );
  AND3_X1 U7786 ( .A1(n6261), .A2(n6260), .A3(n6259), .ZN(n6278) );
  NAND2_X1 U7787 ( .A1(n6263), .A2(n6262), .ZN(n6264) );
  NAND2_X1 U7788 ( .A1(n6264), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7789 ( .A1(n6285), .A2(n6284), .ZN(n6265) );
  NAND2_X1 U7790 ( .A1(n6265), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6267) );
  XNOR2_X1 U7791 ( .A(n7687), .B(P2_B_REG_SCAN_IN), .ZN(n6272) );
  NAND2_X1 U7792 ( .A1(n6268), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6269) );
  MUX2_X1 U7793 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6269), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n6271) );
  NAND2_X1 U7794 ( .A1(n6271), .A2(n6270), .ZN(n7741) );
  NAND2_X1 U7795 ( .A1(n6272), .A2(n7741), .ZN(n6276) );
  NAND2_X1 U7796 ( .A1(n6270), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6274) );
  INV_X1 U7797 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6273) );
  XNOR2_X1 U7798 ( .A(n6274), .B(n6273), .ZN(n7821) );
  INV_X1 U7799 ( .A(n7821), .ZN(n6275) );
  INV_X1 U7800 ( .A(n9787), .ZN(n6277) );
  NOR2_X1 U7801 ( .A1(n6278), .A2(n6277), .ZN(n6646) );
  INV_X1 U7802 ( .A(n6646), .ZN(n6283) );
  INV_X1 U7803 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9790) );
  AND2_X1 U7804 ( .A1(n7687), .A2(n7821), .ZN(n9791) );
  AOI21_X1 U7805 ( .B1(n9787), .B2(n9790), .A(n9791), .ZN(n6806) );
  INV_X1 U7806 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7807 ( .A1(n9787), .A2(n6279), .ZN(n6281) );
  AND2_X1 U7808 ( .A1(n7821), .A2(n7741), .ZN(n9793) );
  INV_X1 U7809 ( .A(n9793), .ZN(n6280) );
  NAND2_X1 U7810 ( .A1(n6281), .A2(n6280), .ZN(n6802) );
  INV_X1 U7811 ( .A(n6802), .ZN(n6282) );
  NAND3_X1 U7812 ( .A1(n6283), .A2(n6806), .A3(n6282), .ZN(n6309) );
  XNOR2_X1 U7813 ( .A(n6285), .B(n6284), .ZN(n6423) );
  NAND2_X1 U7814 ( .A1(n6460), .A2(n9794), .ZN(n9788) );
  INV_X1 U7815 ( .A(n6293), .ZN(n6653) );
  AND2_X1 U7816 ( .A1(n8235), .A2(n8223), .ZN(n6462) );
  OR2_X1 U7817 ( .A1(n9844), .A2(n6462), .ZN(n6286) );
  NOR2_X1 U7818 ( .A1(n6301), .A2(n6286), .ZN(n7594) );
  NAND2_X1 U7819 ( .A1(n8273), .A2(n4970), .ZN(n6317) );
  NAND3_X1 U7820 ( .A1(n6288), .A2(n7594), .A3(n6290), .ZN(n6316) );
  INV_X1 U7821 ( .A(n6289), .ZN(n6291) );
  NAND3_X1 U7822 ( .A1(n6291), .A2(n7594), .A3(n6290), .ZN(n6315) );
  NOR2_X1 U7823 ( .A1(n6293), .A2(n8226), .ZN(n6809) );
  INV_X1 U7824 ( .A(n6809), .ZN(n6294) );
  OR2_X1 U7825 ( .A1(n9838), .A2(n4504), .ZN(n6647) );
  OAI21_X2 U7826 ( .B1(n6301), .B2(n6294), .A(n9750), .ZN(n8336) );
  OR2_X1 U7827 ( .A1(n8252), .A2(n6295), .ZN(n6300) );
  INV_X1 U7828 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9966) );
  NAND2_X1 U7829 ( .A1(n4399), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U7830 ( .A1(n6505), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6296) );
  OAI211_X1 U7831 ( .C1(n5910), .C2(n9966), .A(n6297), .B(n6296), .ZN(n6298)
         );
  INV_X1 U7832 ( .A(n6298), .ZN(n6299) );
  INV_X1 U7833 ( .A(n6301), .ZN(n6302) );
  INV_X1 U7834 ( .A(n6305), .ZN(n8232) );
  NAND2_X1 U7835 ( .A1(n6302), .A2(n8232), .ZN(n7627) );
  INV_X1 U7836 ( .A(n6462), .ZN(n6650) );
  INV_X1 U7837 ( .A(n8765), .ZN(n6304) );
  OAI22_X1 U7838 ( .A1(n8438), .A2(n8333), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6303), .ZN(n6313) );
  INV_X1 U7839 ( .A(n9844), .ZN(n9854) );
  AND2_X1 U7840 ( .A1(n6462), .A2(n6305), .ZN(n6644) );
  INV_X1 U7841 ( .A(n6644), .ZN(n6306) );
  NAND3_X1 U7842 ( .A1(n6460), .A2(n6423), .A3(n6306), .ZN(n6307) );
  AOI21_X1 U7843 ( .B1(n6309), .B2(n9854), .A(n6307), .ZN(n6308) );
  OR2_X1 U7844 ( .A1(n6308), .A2(P2_U3152), .ZN(n6311) );
  INV_X1 U7845 ( .A(n9788), .ZN(n8233) );
  NAND3_X1 U7846 ( .A1(n6309), .A2(n8233), .A3(n6809), .ZN(n6310) );
  OAI22_X1 U7847 ( .A1(n8471), .A2(n8330), .B1(n8332), .B2(n8443), .ZN(n6312)
         );
  AOI211_X1 U7848 ( .C1(n8442), .C2(n8336), .A(n6313), .B(n6312), .ZN(n6314)
         );
  NAND4_X1 U7849 ( .A1(n6317), .A2(n6316), .A3(n6315), .A4(n6314), .ZN(
        P2_U3222) );
  INV_X1 U7850 ( .A(n9794), .ZN(n6318) );
  INV_X2 U7851 ( .A(n8354), .ZN(P2_U3966) );
  INV_X1 U7852 ( .A(n6785), .ZN(n6788) );
  AND2_X1 U7853 ( .A1(n6319), .A2(n6788), .ZN(n6350) );
  NAND2_X1 U7854 ( .A1(n6981), .A2(n6785), .ZN(n6320) );
  NAND2_X1 U7855 ( .A1(n6320), .A2(n6319), .ZN(n8991) );
  NAND2_X1 U7856 ( .A1(n8991), .A2(n5408), .ZN(n6321) );
  NAND2_X1 U7857 ( .A1(n6321), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  AND2_X1 U7858 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n8880) );
  INV_X1 U7859 ( .A(n6344), .ZN(n6496) );
  AOI22_X1 U7860 ( .A1(n6344), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7428), .B2(
        n6496), .ZN(n6494) );
  INV_X1 U7861 ( .A(n6343), .ZN(n6440) );
  AOI22_X1 U7862 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6343), .B1(n6440), .B2(
        n7284), .ZN(n6435) );
  NOR2_X1 U7863 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6338), .ZN(n6322) );
  AOI21_X1 U7864 ( .B1(n6338), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6322), .ZN(
        n9572) );
  INV_X1 U7865 ( .A(n9562), .ZN(n6326) );
  INV_X1 U7866 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6325) );
  INV_X1 U7867 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6324) );
  INV_X1 U7868 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6323) );
  MUX2_X1 U7869 ( .A(n6323), .B(P1_REG2_REG_1__SCAN_IN), .S(n6590), .Z(n6596)
         );
  AND2_X1 U7870 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6851) );
  NAND2_X1 U7871 ( .A1(n6596), .A2(n6851), .ZN(n6595) );
  OAI21_X1 U7872 ( .B1(n6323), .B2(n6590), .A(n6595), .ZN(n6859) );
  MUX2_X1 U7873 ( .A(n6324), .B(P1_REG2_REG_2__SCAN_IN), .S(n6861), .Z(n6860)
         );
  NAND2_X1 U7874 ( .A1(n6859), .A2(n6860), .ZN(n6858) );
  OAI21_X1 U7875 ( .B1(n6324), .B2(n6861), .A(n6858), .ZN(n6571) );
  MUX2_X1 U7876 ( .A(n6325), .B(P1_REG2_REG_3__SCAN_IN), .S(n6567), .Z(n6572)
         );
  NAND2_X1 U7877 ( .A1(n6571), .A2(n6572), .ZN(n6570) );
  OAI21_X1 U7878 ( .B1(n6325), .B2(n6567), .A(n6570), .ZN(n9560) );
  MUX2_X1 U7879 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n5469), .S(n9562), .Z(n9561)
         );
  NOR2_X1 U7880 ( .A1(n9560), .A2(n9561), .ZN(n9559) );
  NAND2_X1 U7881 ( .A1(n6341), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6327) );
  OAI21_X1 U7882 ( .B1(n6341), .B2(P1_REG2_REG_6__SCAN_IN), .A(n6327), .ZN(
        n6629) );
  NOR2_X1 U7883 ( .A1(n6630), .A2(n6629), .ZN(n6628) );
  OAI21_X1 U7884 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6344), .A(n6492), .ZN(
        n6331) );
  NAND2_X1 U7885 ( .A1(n6369), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6328) );
  OAI21_X1 U7886 ( .B1(n6369), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6328), .ZN(
        n6330) );
  NOR2_X1 U7887 ( .A1(n6331), .A2(n6330), .ZN(n6360) );
  OR2_X1 U7888 ( .A1(n5766), .A2(P1_U3084), .ZN(n7822) );
  NOR2_X1 U7889 ( .A1(n4391), .A2(n7822), .ZN(n6329) );
  AND2_X1 U7890 ( .A1(n8991), .A2(n6329), .ZN(n9575) );
  INV_X1 U7891 ( .A(n9575), .ZN(n9591) );
  AOI211_X1 U7892 ( .C1(n6331), .C2(n6330), .A(n6360), .B(n9591), .ZN(n6355)
         );
  NOR2_X1 U7893 ( .A1(n6341), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U7894 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6338), .ZN(n6340) );
  MUX2_X1 U7895 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6332), .S(n9562), .Z(n9554)
         );
  MUX2_X1 U7896 ( .A(n6333), .B(P1_REG1_REG_3__SCAN_IN), .S(n6567), .Z(n6568)
         );
  MUX2_X1 U7897 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6591), .S(n6590), .Z(n6334)
         );
  INV_X1 U7898 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n8986) );
  NOR2_X1 U7899 ( .A1(n6590), .A2(n6591), .ZN(n6862) );
  MUX2_X1 U7900 ( .A(n6335), .B(P1_REG1_REG_2__SCAN_IN), .S(n6861), .Z(n6336)
         );
  OAI21_X1 U7901 ( .B1(n6867), .B2(n6862), .A(n6336), .ZN(n6865) );
  OAI21_X1 U7902 ( .B1(n6333), .B2(n6567), .A(n6337), .ZN(n9555) );
  NOR2_X1 U7903 ( .A1(n9554), .A2(n9555), .ZN(n9553) );
  MUX2_X1 U7904 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6339), .S(n6338), .Z(n9577)
         );
  NAND2_X1 U7905 ( .A1(n9578), .A2(n9577), .ZN(n9576) );
  NAND2_X1 U7906 ( .A1(n6340), .A2(n9576), .ZN(n6633) );
  AOI22_X1 U7907 ( .A1(n6341), .A2(n5442), .B1(P1_REG1_REG_6__SCAN_IN), .B2(
        n6635), .ZN(n6632) );
  NOR2_X1 U7908 ( .A1(n6633), .A2(n6632), .ZN(n6631) );
  AOI22_X1 U7909 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6440), .B1(n6343), .B2(
        n5489), .ZN(n6437) );
  NOR2_X1 U7910 ( .A1(n6438), .A2(n6437), .ZN(n6436) );
  INV_X1 U7911 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9681) );
  NAND2_X1 U7912 ( .A1(n6496), .A2(n9681), .ZN(n6495) );
  AOI22_X1 U7913 ( .A1(n6498), .A2(n6495), .B1(P1_REG1_REG_8__SCAN_IN), .B2(
        n6344), .ZN(n6347) );
  MUX2_X1 U7914 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6345), .S(n6369), .Z(n6346)
         );
  NAND2_X1 U7915 ( .A1(n6347), .A2(n6346), .ZN(n6368) );
  OAI21_X1 U7916 ( .B1(n6347), .B2(n6346), .A(n6368), .ZN(n6349) );
  OR2_X1 U7917 ( .A1(n4391), .A2(P1_U3084), .ZN(n9476) );
  NOR2_X1 U7918 ( .A1(n9476), .A2(n9075), .ZN(n6348) );
  NAND2_X1 U7919 ( .A1(n8991), .A2(n6348), .ZN(n9558) );
  INV_X1 U7920 ( .A(n9558), .ZN(n9597) );
  AND2_X1 U7921 ( .A1(n6349), .A2(n9597), .ZN(n6354) );
  INV_X1 U7922 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10227) );
  INV_X1 U7923 ( .A(n6369), .ZN(n6416) );
  INV_X1 U7924 ( .A(n7822), .ZN(n6351) );
  AND2_X1 U7925 ( .A1(n6351), .A2(n4391), .ZN(n6352) );
  NAND2_X1 U7926 ( .A1(n8991), .A2(n6352), .ZN(n9583) );
  OAI22_X1 U7927 ( .A1(n9586), .A2(n10227), .B1(n6416), .B2(n9583), .ZN(n6353)
         );
  OR4_X1 U7928 ( .A1(n8880), .A2(n6355), .A3(n6354), .A4(n6353), .ZN(P1_U3250)
         );
  INV_X1 U7929 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6356) );
  MUX2_X1 U7930 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n6356), .S(n7083), .Z(n6357)
         );
  INV_X1 U7931 ( .A(n6357), .ZN(n7086) );
  NAND2_X1 U7932 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6642), .ZN(n6358) );
  OAI21_X1 U7933 ( .B1(n6642), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6358), .ZN(
        n6920) );
  NOR2_X1 U7934 ( .A1(n6371), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6359) );
  AOI21_X1 U7935 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6371), .A(n6359), .ZN(
        n8998) );
  NAND2_X1 U7936 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6370), .ZN(n6361) );
  OAI21_X1 U7937 ( .B1(n6370), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6361), .ZN(
        n9593) );
  OAI21_X1 U7938 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6371), .A(n8996), .ZN(
        n6921) );
  INV_X1 U7939 ( .A(n6373), .ZN(n7397) );
  NOR2_X1 U7940 ( .A1(n6362), .A2(n7397), .ZN(n6363) );
  XNOR2_X1 U7941 ( .A(n6362), .B(n7397), .ZN(n7399) );
  NOR2_X1 U7942 ( .A1(n7707), .A2(n7399), .ZN(n7398) );
  NOR2_X1 U7943 ( .A1(n6363), .A2(n7398), .ZN(n9010) );
  XNOR2_X1 U7944 ( .A(n9010), .B(n9017), .ZN(n6364) );
  NOR2_X1 U7945 ( .A1(n7764), .A2(n6364), .ZN(n9011) );
  AOI211_X1 U7946 ( .C1(n6364), .C2(n7764), .A(n9011), .B(n9591), .ZN(n6379)
         );
  INV_X1 U7947 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n6365) );
  NOR2_X1 U7948 ( .A1(n9586), .A2(n6365), .ZN(n6378) );
  INV_X1 U7949 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6375) );
  MUX2_X1 U7950 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6366), .S(n7083), .Z(n7082)
         );
  MUX2_X1 U7951 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6367), .S(n6642), .Z(n6914)
         );
  INV_X1 U7952 ( .A(n6371), .ZN(n9000) );
  AOI22_X1 U7953 ( .A1(n6371), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n5310), .B2(
        n9000), .ZN(n9005) );
  INV_X1 U7954 ( .A(n6370), .ZN(n9584) );
  AOI22_X1 U7955 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6370), .B1(n9584), .B2(
        n5328), .ZN(n9590) );
  OAI21_X1 U7956 ( .B1(n6369), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6368), .ZN(
        n9589) );
  NAND2_X1 U7957 ( .A1(n9590), .A2(n9589), .ZN(n9588) );
  OAI21_X1 U7958 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6371), .A(n9003), .ZN(
        n6915) );
  NAND2_X1 U7959 ( .A1(n6914), .A2(n6915), .ZN(n6913) );
  OAI21_X1 U7960 ( .B1(n7083), .B2(P1_REG1_REG_13__SCAN_IN), .A(n7080), .ZN(
        n7395) );
  MUX2_X1 U7961 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n6372), .S(n6373), .Z(n7396)
         );
  NAND2_X1 U7962 ( .A1(n7395), .A2(n7396), .ZN(n7394) );
  OAI21_X1 U7963 ( .B1(n6373), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7394), .ZN(
        n9016) );
  NOR2_X1 U7964 ( .A1(n6375), .A2(n6374), .ZN(n9018) );
  AOI211_X1 U7965 ( .C1(n6375), .C2(n6374), .A(n9018), .B(n9558), .ZN(n6377)
         );
  NAND2_X1 U7966 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3084), .ZN(n8959) );
  OAI21_X1 U7967 ( .B1(n9583), .B2(n9017), .A(n8959), .ZN(n6376) );
  OR4_X1 U7968 ( .A1(n6379), .A2(n6378), .A3(n6377), .A4(n6376), .ZN(P1_U3256)
         );
  XNOR2_X1 U7969 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U7970 ( .A1(n6380), .A2(P2_U3152), .ZN(n8758) );
  INV_X2 U7971 ( .A(n8758), .ZN(n8771) );
  INV_X1 U7972 ( .A(n8378), .ZN(n6449) );
  OAI222_X1 U7973 ( .A1(n8771), .A2(n6381), .B1(n8769), .B2(n6395), .C1(
        P2_U3152), .C2(n6449), .ZN(P2_U3356) );
  INV_X1 U7974 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6382) );
  OAI222_X1 U7975 ( .A1(n8771), .A2(n6382), .B1(n8769), .B2(n6385), .C1(
        P2_U3152), .C2(n6627), .ZN(P2_U3357) );
  INV_X1 U7976 ( .A(n6535), .ZN(n6542) );
  OAI222_X1 U7977 ( .A1(n8771), .A2(n6383), .B1(n8769), .B2(n6389), .C1(
        P2_U3152), .C2(n6542), .ZN(P2_U3355) );
  OR2_X1 U7978 ( .A1(n6384), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9479) );
  NAND2_X1 U7979 ( .A1(n6384), .A2(P1_U3084), .ZN(n9466) );
  OAI222_X1 U7980 ( .A1(n9479), .A2(n6386), .B1(n9466), .B2(n6385), .C1(
        P1_U3084), .C2(n6590), .ZN(P1_U3352) );
  INV_X1 U7981 ( .A(n6520), .ZN(n6474) );
  OAI222_X1 U7982 ( .A1(n8771), .A2(n6387), .B1(n8769), .B2(n6393), .C1(
        P2_U3152), .C2(n6474), .ZN(P2_U3354) );
  INV_X1 U7983 ( .A(n9479), .ZN(n7078) );
  INV_X1 U7984 ( .A(n7078), .ZN(n9468) );
  OAI222_X1 U7985 ( .A1(P1_U3084), .A2(n6567), .B1(n9466), .B2(n6389), .C1(
        n6388), .C2(n9468), .ZN(P1_U3350) );
  OAI222_X1 U7986 ( .A1(n8771), .A2(n6390), .B1(n8769), .B2(n6391), .C1(
        P2_U3152), .C2(n6618), .ZN(P2_U3353) );
  INV_X1 U7987 ( .A(n9466), .ZN(n9474) );
  INV_X1 U7988 ( .A(n9474), .ZN(n9473) );
  OAI222_X1 U7989 ( .A1(n9468), .A2(n6392), .B1(n9473), .B2(n6391), .C1(
        P1_U3084), .C2(n9568), .ZN(P1_U3348) );
  OAI222_X1 U7990 ( .A1(n9468), .A2(n6394), .B1(n9473), .B2(n6393), .C1(
        P1_U3084), .C2(n9562), .ZN(P1_U3349) );
  OAI222_X1 U7991 ( .A1(n9479), .A2(n6396), .B1(n9473), .B2(n6395), .C1(
        P1_U3084), .C2(n6861), .ZN(P1_U3351) );
  OAI222_X1 U7992 ( .A1(n9468), .A2(n9989), .B1(n9473), .B2(n6398), .C1(
        P1_U3084), .C2(n6635), .ZN(P1_U3347) );
  INV_X1 U7993 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6399) );
  OAI222_X1 U7994 ( .A1(n8771), .A2(n6399), .B1(n8769), .B2(n6398), .C1(
        P2_U3152), .C2(n6397), .ZN(P2_U3352) );
  INV_X1 U7995 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6401) );
  INV_X1 U7996 ( .A(n6400), .ZN(n6402) );
  INV_X1 U7997 ( .A(n6549), .ZN(n6476) );
  OAI222_X1 U7998 ( .A1(n8771), .A2(n6401), .B1(n8769), .B2(n6402), .C1(
        P2_U3152), .C2(n6476), .ZN(P2_U3351) );
  INV_X1 U7999 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6403) );
  OAI222_X1 U8000 ( .A1(n9468), .A2(n6403), .B1(n9466), .B2(n6402), .C1(
        P1_U3084), .C2(n6440), .ZN(P1_U3346) );
  INV_X1 U8001 ( .A(n6795), .ZN(n9617) );
  NAND2_X1 U8002 ( .A1(n7739), .A2(P1_B_REG_SCAN_IN), .ZN(n6404) );
  INV_X1 U8003 ( .A(n7689), .ZN(n6406) );
  MUX2_X1 U8004 ( .A(n6404), .B(P1_B_REG_SCAN_IN), .S(n6406), .Z(n6405) );
  INV_X1 U8005 ( .A(n7826), .ZN(n6407) );
  INV_X1 U8006 ( .A(n9616), .ZN(n6713) );
  OAI22_X1 U8007 ( .A1(n6713), .A2(P1_D_REG_0__SCAN_IN), .B1(n6407), .B2(n6406), .ZN(n6725) );
  NAND2_X1 U8008 ( .A1(n9617), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6408) );
  OAI21_X1 U8009 ( .B1(n9617), .B2(n6725), .A(n6408), .ZN(P1_U3440) );
  INV_X1 U8010 ( .A(n6409), .ZN(n6410) );
  OAI222_X1 U8011 ( .A1(n9468), .A2(n10091), .B1(n9466), .B2(n6410), .C1(
        P1_U3084), .C2(n6496), .ZN(P1_U3345) );
  INV_X1 U8012 ( .A(n9694), .ZN(n6477) );
  OAI222_X1 U8013 ( .A1(n8771), .A2(n6411), .B1(n8769), .B2(n6410), .C1(
        P2_U3152), .C2(n6477), .ZN(P2_U3350) );
  INV_X1 U8014 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10152) );
  NAND2_X1 U8015 ( .A1(n9616), .A2(n10152), .ZN(n6413) );
  NAND2_X1 U8016 ( .A1(n7826), .A2(n7739), .ZN(n6412) );
  NAND2_X1 U8017 ( .A1(n6413), .A2(n6412), .ZN(n7147) );
  OR2_X1 U8018 ( .A1(n9617), .A2(n7147), .ZN(n6782) );
  OAI21_X1 U8019 ( .B1(n6795), .B2(n10152), .A(n6782), .ZN(P1_U3441) );
  INV_X1 U8020 ( .A(n6414), .ZN(n6417) );
  INV_X1 U8021 ( .A(n6561), .ZN(n6479) );
  OAI222_X1 U8022 ( .A1(n8771), .A2(n6415), .B1(n8769), .B2(n6417), .C1(n6479), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI222_X1 U8023 ( .A1(n9479), .A2(n9976), .B1(n9466), .B2(n6417), .C1(n6416), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8024 ( .A(n6418), .ZN(n6420) );
  OAI222_X1 U8025 ( .A1(n8771), .A2(n6419), .B1(n8769), .B2(n6420), .C1(
        P2_U3152), .C2(n6480), .ZN(P2_U3348) );
  OAI222_X1 U8026 ( .A1(n9479), .A2(n6421), .B1(n9466), .B2(n6420), .C1(
        P1_U3084), .C2(n9584), .ZN(P1_U3343) );
  NAND2_X1 U8027 ( .A1(n8354), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6422) );
  OAI21_X1 U8028 ( .B1(n8551), .B2(n8354), .A(n6422), .ZN(P2_U3574) );
  OR2_X1 U8029 ( .A1(n6423), .A2(P2_U3152), .ZN(n8237) );
  NAND2_X1 U8030 ( .A1(n9788), .A2(n8237), .ZN(n6425) );
  NAND2_X1 U8031 ( .A1(n6425), .A2(n4402), .ZN(n6427) );
  OR2_X1 U8032 ( .A1(n9788), .A2(n6650), .ZN(n6426) );
  INV_X1 U8033 ( .A(n8419), .ZN(n9707) );
  NOR2_X1 U8034 ( .A1(n9707), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8035 ( .A(n6428), .ZN(n6430) );
  INV_X1 U8036 ( .A(n6681), .ZN(n6688) );
  OAI222_X1 U8037 ( .A1(n8771), .A2(n6429), .B1(n8769), .B2(n6430), .C1(n6688), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  OAI222_X1 U8038 ( .A1(n9479), .A2(n6431), .B1(n9466), .B2(n6430), .C1(n9000), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  NAND2_X1 U8039 ( .A1(n6791), .A2(P1_U4006), .ZN(n6432) );
  OAI21_X1 U8040 ( .B1(P1_U4006), .B2(n5836), .A(n6432), .ZN(P1_U3555) );
  INV_X1 U8041 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10186) );
  OAI21_X1 U8042 ( .B1(n6435), .B2(n6434), .A(n6433), .ZN(n6443) );
  AOI21_X1 U8043 ( .B1(n6438), .B2(n6437), .A(n6436), .ZN(n6439) );
  NOR2_X1 U8044 ( .A1(n9558), .A2(n6439), .ZN(n6442) );
  NAND2_X1 U8045 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3084), .ZN(n7376) );
  OAI21_X1 U8046 ( .B1(n9583), .B2(n6440), .A(n7376), .ZN(n6441) );
  AOI211_X1 U8047 ( .C1(n9575), .C2(n6443), .A(n6442), .B(n6441), .ZN(n6444)
         );
  OAI21_X1 U8048 ( .B1(n10186), .B2(n9586), .A(n6444), .ZN(P1_U3248) );
  INV_X1 U8049 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6456) );
  MUX2_X1 U8050 ( .A(n6456), .B(P2_REG2_REG_10__SCAN_IN), .S(n6480), .Z(n9716)
         );
  NAND2_X1 U8051 ( .A1(n6561), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6455) );
  INV_X1 U8052 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6445) );
  MUX2_X1 U8053 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6445), .S(n6561), .Z(n6563)
         );
  NAND2_X1 U8054 ( .A1(n9694), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6454) );
  INV_X1 U8055 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7127) );
  MUX2_X1 U8056 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7127), .S(n9694), .Z(n9696)
         );
  INV_X1 U8057 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6453) );
  MUX2_X1 U8058 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6453), .S(n6549), .Z(n6551)
         );
  NAND2_X1 U8059 ( .A1(n6584), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6452) );
  INV_X1 U8060 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6446) );
  MUX2_X1 U8061 ( .A(n6446), .B(P2_REG2_REG_6__SCAN_IN), .S(n6584), .Z(n6447)
         );
  INV_X1 U8062 ( .A(n6447), .ZN(n6586) );
  INV_X1 U8063 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10153) );
  INV_X1 U8064 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7010) );
  MUX2_X1 U8065 ( .A(n7010), .B(P2_REG2_REG_1__SCAN_IN), .S(n6627), .Z(n6623)
         );
  NAND3_X1 U8066 ( .A1(n6623), .A2(P2_REG2_REG_0__SCAN_IN), .A3(n9691), .ZN(
        n8375) );
  NAND2_X1 U8067 ( .A1(n6448), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8374) );
  INV_X1 U8068 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9961) );
  MUX2_X1 U8069 ( .A(n9961), .B(P2_REG2_REG_2__SCAN_IN), .S(n8378), .Z(n8373)
         );
  NOR2_X1 U8070 ( .A1(n6449), .A2(n9961), .ZN(n6534) );
  INV_X1 U8071 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6908) );
  MUX2_X1 U8072 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6908), .S(n6535), .Z(n6450)
         );
  OAI21_X1 U8073 ( .B1(n6533), .B2(n6534), .A(n6450), .ZN(n6539) );
  NAND2_X1 U8074 ( .A1(n6535), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6522) );
  INV_X1 U8075 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10185) );
  MUX2_X1 U8076 ( .A(n10185), .B(P2_REG2_REG_4__SCAN_IN), .S(n6520), .Z(n6521)
         );
  NOR2_X1 U8077 ( .A1(n6474), .A2(n10185), .ZN(n6610) );
  MUX2_X1 U8078 ( .A(n10153), .B(P2_REG2_REG_5__SCAN_IN), .S(n6618), .Z(n6451)
         );
  OAI21_X1 U8079 ( .B1(n6615), .B2(n6610), .A(n6451), .ZN(n6613) );
  OAI21_X1 U8080 ( .B1(n10153), .B2(n6618), .A(n6613), .ZN(n6587) );
  NAND2_X1 U8081 ( .A1(n6586), .A2(n6587), .ZN(n6585) );
  NAND2_X1 U8082 ( .A1(n6452), .A2(n6585), .ZN(n6552) );
  NAND2_X1 U8083 ( .A1(n6551), .A2(n6552), .ZN(n6550) );
  OAI21_X1 U8084 ( .B1(n6476), .B2(n6453), .A(n6550), .ZN(n9697) );
  NAND2_X1 U8085 ( .A1(n9696), .A2(n9697), .ZN(n9695) );
  NAND2_X1 U8086 ( .A1(n6454), .A2(n9695), .ZN(n6564) );
  NAND2_X1 U8087 ( .A1(n6563), .A2(n6564), .ZN(n6562) );
  NAND2_X1 U8088 ( .A1(n6455), .A2(n6562), .ZN(n9717) );
  NAND2_X1 U8089 ( .A1(n9716), .A2(n9717), .ZN(n9714) );
  OAI21_X1 U8090 ( .B1(n6456), .B2(n6480), .A(n9714), .ZN(n6459) );
  INV_X1 U8091 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6457) );
  AOI22_X1 U8092 ( .A1(n6681), .A2(n6457), .B1(P2_REG2_REG_11__SCAN_IN), .B2(
        n6688), .ZN(n6458) );
  NOR2_X1 U8093 ( .A1(n6459), .A2(n6458), .ZN(n6682) );
  AOI21_X1 U8094 ( .B1(n6459), .B2(n6458), .A(n6682), .ZN(n6490) );
  OAI21_X1 U8095 ( .B1(n6460), .B2(P2_U3152), .A(n8237), .ZN(n6461) );
  INV_X1 U8096 ( .A(n6461), .ZN(n6464) );
  OR2_X1 U8097 ( .A1(n9788), .A2(n6462), .ZN(n6463) );
  NAND2_X1 U8098 ( .A1(n6464), .A2(n6463), .ZN(n6484) );
  NAND2_X1 U8099 ( .A1(n6484), .A2(n6482), .ZN(n6465) );
  NAND2_X1 U8100 ( .A1(n6465), .A2(n8354), .ZN(n6467) );
  NOR2_X1 U8101 ( .A1(n8765), .A2(n8767), .ZN(n6466) );
  NAND2_X1 U8102 ( .A1(n6467), .A2(n6466), .ZN(n9686) );
  AND2_X1 U8103 ( .A1(n6467), .A2(n8765), .ZN(n9709) );
  INV_X1 U8104 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10159) );
  INV_X1 U8105 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9874) );
  MUX2_X1 U8106 ( .A(n9874), .B(P2_REG1_REG_10__SCAN_IN), .S(n6480), .Z(n9712)
         );
  INV_X1 U8107 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6478) );
  MUX2_X1 U8108 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6478), .S(n6561), .Z(n6556)
         );
  INV_X1 U8109 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9872) );
  MUX2_X1 U8110 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9872), .S(n9694), .Z(n9699)
         );
  INV_X1 U8111 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9870) );
  MUX2_X1 U8112 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9870), .S(n6549), .Z(n6544)
         );
  NAND2_X1 U8113 ( .A1(n6584), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6475) );
  INV_X1 U8114 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6468) );
  MUX2_X1 U8115 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6468), .S(n6584), .Z(n6579)
         );
  INV_X1 U8116 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9868) );
  INV_X1 U8117 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9862) );
  MUX2_X1 U8118 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9862), .S(n6627), .Z(n6619)
         );
  NAND2_X1 U8119 ( .A1(n9691), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6620) );
  NOR2_X1 U8120 ( .A1(n6619), .A2(n6620), .ZN(n8384) );
  NOR2_X1 U8121 ( .A1(n6627), .A2(n9862), .ZN(n8379) );
  INV_X1 U8122 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6469) );
  MUX2_X1 U8123 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6469), .S(n8378), .Z(n6470)
         );
  OAI21_X1 U8124 ( .B1(n8384), .B2(n8379), .A(n6470), .ZN(n8382) );
  NAND2_X1 U8125 ( .A1(n8378), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U8126 ( .A1(n8382), .A2(n6528), .ZN(n6473) );
  INV_X1 U8127 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6471) );
  MUX2_X1 U8128 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6471), .S(n6535), .Z(n6472)
         );
  NAND2_X1 U8129 ( .A1(n6473), .A2(n6472), .ZN(n6530) );
  NAND2_X1 U8130 ( .A1(n6535), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6514) );
  INV_X1 U8131 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9866) );
  MUX2_X1 U8132 ( .A(n9866), .B(P2_REG1_REG_4__SCAN_IN), .S(n6520), .Z(n6513)
         );
  AOI21_X1 U8133 ( .B1(n6530), .B2(n6514), .A(n6513), .ZN(n6605) );
  NOR2_X1 U8134 ( .A1(n6474), .A2(n9866), .ZN(n6604) );
  MUX2_X1 U8135 ( .A(n9868), .B(P2_REG1_REG_5__SCAN_IN), .S(n6618), .Z(n6603)
         );
  OAI21_X1 U8136 ( .B1(n6605), .B2(n6604), .A(n6603), .ZN(n6602) );
  OAI21_X1 U8137 ( .B1(n9868), .B2(n6618), .A(n6602), .ZN(n6580) );
  NAND2_X1 U8138 ( .A1(n6579), .A2(n6580), .ZN(n6578) );
  NAND2_X1 U8139 ( .A1(n6475), .A2(n6578), .ZN(n6545) );
  NAND2_X1 U8140 ( .A1(n6544), .A2(n6545), .ZN(n6543) );
  OAI21_X1 U8141 ( .B1(n6476), .B2(n9870), .A(n6543), .ZN(n9700) );
  NAND2_X1 U8142 ( .A1(n9699), .A2(n9700), .ZN(n9698) );
  OAI21_X1 U8143 ( .B1(n6477), .B2(n9872), .A(n9698), .ZN(n6557) );
  NAND2_X1 U8144 ( .A1(n6556), .A2(n6557), .ZN(n6555) );
  OAI21_X1 U8145 ( .B1(n6479), .B2(n6478), .A(n6555), .ZN(n9713) );
  NAND2_X1 U8146 ( .A1(n9712), .A2(n9713), .ZN(n9710) );
  OAI21_X1 U8147 ( .B1(n6480), .B2(n9874), .A(n9710), .ZN(n6486) );
  INV_X1 U8148 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6481) );
  MUX2_X1 U8149 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6481), .S(n6681), .Z(n6485)
         );
  AND2_X1 U8150 ( .A1(n6482), .A2(n8767), .ZN(n6483) );
  NAND2_X1 U8151 ( .A1(n6485), .A2(n6486), .ZN(n6687) );
  OAI211_X1 U8152 ( .C1(n6486), .C2(n6485), .A(n9711), .B(n6687), .ZN(n6487)
         );
  NAND2_X1 U8153 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3152), .ZN(n7218) );
  OAI211_X1 U8154 ( .C1(n8419), .C2(n10159), .A(n6487), .B(n7218), .ZN(n6488)
         );
  AOI21_X1 U8155 ( .B1(n6681), .B2(n9709), .A(n6488), .ZN(n6489) );
  OAI21_X1 U8156 ( .B1(n6490), .B2(n9686), .A(n6489), .ZN(P2_U3256) );
  NAND2_X1 U8157 ( .A1(n8354), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6491) );
  OAI21_X1 U8158 ( .B1(n8535), .B2(n8354), .A(n6491), .ZN(P2_U3575) );
  INV_X1 U8159 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6504) );
  OAI21_X1 U8160 ( .B1(n6494), .B2(n6493), .A(n6492), .ZN(n6502) );
  NAND2_X1 U8161 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3084), .ZN(n7531) );
  OAI21_X1 U8162 ( .B1(n9583), .B2(n6496), .A(n7531), .ZN(n6501) );
  OAI21_X1 U8163 ( .B1(n9681), .B2(n6496), .A(n6495), .ZN(n6497) );
  XOR2_X1 U8164 ( .A(n6498), .B(n6497), .Z(n6499) );
  NOR2_X1 U8165 ( .A1(n6499), .A2(n9558), .ZN(n6500) );
  AOI211_X1 U8166 ( .C1(n9575), .C2(n6502), .A(n6501), .B(n6500), .ZN(n6503)
         );
  OAI21_X1 U8167 ( .B1(n9586), .B2(n6504), .A(n6503), .ZN(P1_U3249) );
  NAND2_X1 U8168 ( .A1(n6505), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U8169 ( .A1(n6506), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U8170 ( .A1(n8025), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6507) );
  AND3_X1 U8171 ( .A1(n6509), .A2(n6508), .A3(n6507), .ZN(n8423) );
  INV_X1 U8172 ( .A(n8423), .ZN(n6510) );
  NAND2_X1 U8173 ( .A1(P2_U3966), .A2(n6510), .ZN(n6511) );
  OAI21_X1 U8174 ( .B1(P2_U3966), .B2(n9461), .A(n6511), .ZN(P2_U3583) );
  NAND2_X1 U8175 ( .A1(n8567), .A2(P2_U3966), .ZN(n6512) );
  OAI21_X1 U8176 ( .B1(P2_U3966), .B2(n5183), .A(n6512), .ZN(P2_U3573) );
  INV_X1 U8177 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6518) );
  INV_X1 U8178 ( .A(n6605), .ZN(n6516) );
  NAND3_X1 U8179 ( .A1(n6530), .A2(n6514), .A3(n6513), .ZN(n6515) );
  NAND3_X1 U8180 ( .A1(n9711), .A2(n6516), .A3(n6515), .ZN(n6517) );
  NAND2_X1 U8181 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n6675) );
  OAI211_X1 U8182 ( .C1(n8419), .C2(n6518), .A(n6517), .B(n6675), .ZN(n6519)
         );
  AOI21_X1 U8183 ( .B1(n6520), .B2(n9709), .A(n6519), .ZN(n6526) );
  INV_X1 U8184 ( .A(n6615), .ZN(n6524) );
  NAND3_X1 U8185 ( .A1(n6539), .A2(n6522), .A3(n6521), .ZN(n6523) );
  NAND3_X1 U8186 ( .A1(n9715), .A2(n6524), .A3(n6523), .ZN(n6525) );
  NAND2_X1 U8187 ( .A1(n6526), .A2(n6525), .ZN(P2_U3249) );
  INV_X1 U8188 ( .A(n9709), .ZN(n9685) );
  NAND2_X1 U8189 ( .A1(P2_U3152), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6746) );
  INV_X1 U8190 ( .A(n6746), .ZN(n6532) );
  MUX2_X1 U8191 ( .A(n6471), .B(P2_REG1_REG_3__SCAN_IN), .S(n6535), .Z(n6527)
         );
  NAND3_X1 U8192 ( .A1(n8382), .A2(n6528), .A3(n6527), .ZN(n6529) );
  AND3_X1 U8193 ( .A1(n9711), .A2(n6530), .A3(n6529), .ZN(n6531) );
  AOI211_X1 U8194 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n9707), .A(n6532), .B(
        n6531), .ZN(n6541) );
  INV_X1 U8195 ( .A(n6533), .ZN(n8377) );
  INV_X1 U8196 ( .A(n6534), .ZN(n6537) );
  MUX2_X1 U8197 ( .A(n6908), .B(P2_REG2_REG_3__SCAN_IN), .S(n6535), .Z(n6536)
         );
  NAND3_X1 U8198 ( .A1(n8377), .A2(n6537), .A3(n6536), .ZN(n6538) );
  NAND3_X1 U8199 ( .A1(n9715), .A2(n6539), .A3(n6538), .ZN(n6540) );
  OAI211_X1 U8200 ( .C1(n9685), .C2(n6542), .A(n6541), .B(n6540), .ZN(P2_U3248) );
  INV_X1 U8201 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6547) );
  OAI211_X1 U8202 ( .C1(n6545), .C2(n6544), .A(n9711), .B(n6543), .ZN(n6546)
         );
  NAND2_X1 U8203 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3152), .ZN(n6938) );
  OAI211_X1 U8204 ( .C1(n8419), .C2(n6547), .A(n6546), .B(n6938), .ZN(n6548)
         );
  AOI21_X1 U8205 ( .B1(n6549), .B2(n9709), .A(n6548), .ZN(n6554) );
  OAI211_X1 U8206 ( .C1(n6552), .C2(n6551), .A(n9715), .B(n6550), .ZN(n6553)
         );
  NAND2_X1 U8207 ( .A1(n6554), .A2(n6553), .ZN(P2_U3252) );
  INV_X1 U8208 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6559) );
  OAI211_X1 U8209 ( .C1(n6557), .C2(n6556), .A(n9711), .B(n6555), .ZN(n6558)
         );
  NAND2_X1 U8210 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7097) );
  OAI211_X1 U8211 ( .C1(n8419), .C2(n6559), .A(n6558), .B(n7097), .ZN(n6560)
         );
  AOI21_X1 U8212 ( .B1(n6561), .B2(n9709), .A(n6560), .ZN(n6566) );
  OAI211_X1 U8213 ( .C1(n6564), .C2(n6563), .A(n9715), .B(n6562), .ZN(n6565)
         );
  NAND2_X1 U8214 ( .A1(n6566), .A2(n6565), .ZN(P2_U3254) );
  INV_X1 U8215 ( .A(n9586), .ZN(n9022) );
  OAI22_X1 U8216 ( .A1(n9583), .A2(n6567), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6844), .ZN(n6576) );
  XNOR2_X1 U8217 ( .A(n6569), .B(n6568), .ZN(n6574) );
  OAI211_X1 U8218 ( .C1(n6572), .C2(n6571), .A(n9575), .B(n6570), .ZN(n6573)
         );
  OAI21_X1 U8219 ( .B1(n9558), .B2(n6574), .A(n6573), .ZN(n6575) );
  AOI211_X1 U8220 ( .C1(n9022), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n6576), .B(
        n6575), .ZN(n6577) );
  INV_X1 U8221 ( .A(n6577), .ZN(P1_U3244) );
  INV_X1 U8222 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6582) );
  OAI211_X1 U8223 ( .C1(n6580), .C2(n6579), .A(n9711), .B(n6578), .ZN(n6581)
         );
  NAND2_X1 U8224 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n6771) );
  OAI211_X1 U8225 ( .C1(n8419), .C2(n6582), .A(n6581), .B(n6771), .ZN(n6583)
         );
  AOI21_X1 U8226 ( .B1(n6584), .B2(n9709), .A(n6583), .ZN(n6589) );
  OAI211_X1 U8227 ( .C1(n6587), .C2(n6586), .A(n9715), .B(n6585), .ZN(n6588)
         );
  NAND2_X1 U8228 ( .A1(n6589), .A2(n6588), .ZN(P2_U3251) );
  OAI22_X1 U8229 ( .A1(n9583), .A2(n6590), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7159), .ZN(n6600) );
  INV_X1 U8230 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n8988) );
  NOR2_X1 U8231 ( .A1(n8986), .A2(n8988), .ZN(n6594) );
  MUX2_X1 U8232 ( .A(n6591), .B(P1_REG1_REG_1__SCAN_IN), .S(n6590), .Z(n6593)
         );
  INV_X1 U8233 ( .A(n6867), .ZN(n6592) );
  OAI211_X1 U8234 ( .C1(n6594), .C2(n6593), .A(n9597), .B(n6592), .ZN(n6598)
         );
  OAI211_X1 U8235 ( .C1(n6596), .C2(n6851), .A(n9575), .B(n6595), .ZN(n6597)
         );
  NAND2_X1 U8236 ( .A1(n6598), .A2(n6597), .ZN(n6599) );
  AOI211_X1 U8237 ( .C1(n9022), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n6600), .B(
        n6599), .ZN(n6601) );
  INV_X1 U8238 ( .A(n6601), .ZN(P1_U3242) );
  NAND2_X1 U8239 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3152), .ZN(n6753) );
  INV_X1 U8240 ( .A(n6753), .ZN(n6609) );
  INV_X1 U8241 ( .A(n9711), .ZN(n7342) );
  INV_X1 U8242 ( .A(n6602), .ZN(n6607) );
  NOR3_X1 U8243 ( .A1(n6605), .A2(n6604), .A3(n6603), .ZN(n6606) );
  NOR3_X1 U8244 ( .A1(n7342), .A2(n6607), .A3(n6606), .ZN(n6608) );
  AOI211_X1 U8245 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n9707), .A(n6609), .B(
        n6608), .ZN(n6617) );
  MUX2_X1 U8246 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10153), .S(n6618), .Z(n6612)
         );
  INV_X1 U8247 ( .A(n6610), .ZN(n6611) );
  NAND2_X1 U8248 ( .A1(n6612), .A2(n6611), .ZN(n6614) );
  OAI211_X1 U8249 ( .C1(n6615), .C2(n6614), .A(n9715), .B(n6613), .ZN(n6616)
         );
  OAI211_X1 U8250 ( .C1(n9685), .C2(n6618), .A(n6617), .B(n6616), .ZN(P2_U3250) );
  INV_X1 U8251 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7005) );
  NOR2_X1 U8252 ( .A1(n7005), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6622) );
  AOI211_X1 U8253 ( .C1(n6620), .C2(n6619), .A(n8384), .B(n7342), .ZN(n6621)
         );
  AOI211_X1 U8254 ( .C1(P2_ADDR_REG_1__SCAN_IN), .C2(n9707), .A(n6622), .B(
        n6621), .ZN(n6626) );
  INV_X1 U8255 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6813) );
  NOR2_X1 U8256 ( .A1(n4617), .A2(n6813), .ZN(n6624) );
  OAI211_X1 U8257 ( .C1(n6624), .C2(n6623), .A(n9715), .B(n8375), .ZN(n6625)
         );
  OAI211_X1 U8258 ( .C1(n9685), .C2(n6627), .A(n6626), .B(n6625), .ZN(P2_U3246) );
  INV_X1 U8259 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6640) );
  AOI211_X1 U8260 ( .C1(n6630), .C2(n6629), .A(n6628), .B(n9591), .ZN(n6638)
         );
  AOI21_X1 U8261 ( .B1(n6633), .B2(n6632), .A(n6631), .ZN(n6634) );
  NOR2_X1 U8262 ( .A1(n9558), .A2(n6634), .ZN(n6637) );
  NAND2_X1 U8263 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3084), .ZN(n7199) );
  OAI21_X1 U8264 ( .B1(n9583), .B2(n6635), .A(n7199), .ZN(n6636) );
  NOR3_X1 U8265 ( .A1(n6638), .A2(n6637), .A3(n6636), .ZN(n6639) );
  OAI21_X1 U8266 ( .B1(n9586), .B2(n6640), .A(n6639), .ZN(P1_U3247) );
  INV_X1 U8267 ( .A(n6641), .ZN(n6643) );
  INV_X1 U8268 ( .A(n6642), .ZN(n6918) );
  OAI222_X1 U8269 ( .A1(n9479), .A2(n9953), .B1(n9466), .B2(n6643), .C1(
        P1_U3084), .C2(n6918), .ZN(P1_U3341) );
  INV_X1 U8270 ( .A(n8394), .ZN(n6690) );
  OAI222_X1 U8271 ( .A1(n8771), .A2(n10181), .B1(n8769), .B2(n6643), .C1(
        P2_U3152), .C2(n6690), .ZN(P2_U3346) );
  OR2_X1 U8272 ( .A1(n9788), .A2(n6644), .ZN(n6645) );
  NAND2_X1 U8273 ( .A1(n6802), .A2(n6647), .ZN(n6648) );
  NOR2_X1 U8274 ( .A1(n6803), .A2(n6648), .ZN(n6666) );
  INV_X1 U8275 ( .A(n6806), .ZN(n6804) );
  AND2_X2 U8276 ( .A1(n6666), .A2(n6804), .ZN(n9861) );
  NAND2_X1 U8277 ( .A1(n6649), .A2(n6760), .ZN(n8078) );
  NAND2_X1 U8278 ( .A1(n7007), .A2(n8078), .ZN(n8043) );
  NAND2_X1 U8279 ( .A1(n5846), .A2(n6650), .ZN(n9848) );
  NAND2_X1 U8280 ( .A1(n8219), .A2(n8038), .ZN(n9774) );
  NAND2_X1 U8281 ( .A1(n9848), .A2(n9740), .ZN(n6651) );
  NAND2_X1 U8282 ( .A1(n8043), .A2(n6651), .ZN(n6652) );
  INV_X1 U8283 ( .A(n9743), .ZN(n9771) );
  NAND2_X1 U8284 ( .A1(n6891), .A2(n9771), .ZN(n6758) );
  NAND2_X1 U8285 ( .A1(n6652), .A2(n6758), .ZN(n6810) );
  AOI21_X1 U8286 ( .B1(n6653), .B2(n7003), .A(n6810), .ZN(n6668) );
  INV_X1 U8287 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6654) );
  OR2_X1 U8288 ( .A1(n9861), .A2(n6654), .ZN(n6655) );
  OAI21_X1 U8289 ( .B1(n9860), .B2(n6668), .A(n6655), .ZN(P2_U3451) );
  INV_X1 U8290 ( .A(n6656), .ZN(n6660) );
  AOI22_X1 U8291 ( .A1(n7083), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7078), .ZN(n6657) );
  OAI21_X1 U8292 ( .B1(n6660), .B2(n9473), .A(n6657), .ZN(P1_U3340) );
  INV_X1 U8293 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U8294 ( .A1(n9076), .A2(P1_U4006), .ZN(n6658) );
  OAI21_X1 U8295 ( .B1(P1_U4006), .B2(n6659), .A(n6658), .ZN(P1_U3586) );
  INV_X1 U8296 ( .A(n6697), .ZN(n6955) );
  OAI222_X1 U8297 ( .A1(n8771), .A2(n6661), .B1(n8769), .B2(n6660), .C1(n6955), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8298 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6663) );
  INV_X1 U8299 ( .A(n6662), .ZN(n6664) );
  INV_X1 U8300 ( .A(n7046), .ZN(n7051) );
  OAI222_X1 U8301 ( .A1(n8771), .A2(n6663), .B1(n8769), .B2(n6664), .C1(n7051), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8302 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6665) );
  OAI222_X1 U8303 ( .A1(n9479), .A2(n6665), .B1(n9466), .B2(n6664), .C1(n7397), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  AND2_X2 U8304 ( .A1(n6666), .A2(n6806), .ZN(n9879) );
  NAND2_X1 U8305 ( .A1(n9877), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U8306 ( .B1(n9877), .B2(n6668), .A(n6667), .ZN(P2_U3520) );
  NAND2_X1 U8307 ( .A1(n6670), .A2(n6669), .ZN(n6674) );
  NAND2_X1 U8308 ( .A1(n6672), .A2(n6671), .ZN(n6673) );
  XOR2_X1 U8309 ( .A(n6674), .B(n6673), .Z(n6680) );
  INV_X1 U8310 ( .A(n9756), .ZN(n9813) );
  NAND2_X1 U8311 ( .A1(n8336), .A2(n9813), .ZN(n6676) );
  NAND2_X1 U8312 ( .A1(n6676), .A2(n6675), .ZN(n6678) );
  INV_X1 U8313 ( .A(n9772), .ZN(n9746) );
  INV_X1 U8314 ( .A(n8370), .ZN(n9744) );
  OAI22_X1 U8315 ( .A1(n9746), .A2(n8330), .B1(n8333), .B2(n9744), .ZN(n6677)
         );
  AOI211_X1 U8316 ( .C1(n9749), .C2(n8344), .A(n6678), .B(n6677), .ZN(n6679)
         );
  OAI21_X1 U8317 ( .B1(n6680), .B2(n8340), .A(n6679), .ZN(P2_U3232) );
  NAND2_X1 U8318 ( .A1(n8394), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6684) );
  INV_X1 U8319 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8389) );
  NOR2_X1 U8320 ( .A1(n6681), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6683) );
  OAI211_X1 U8321 ( .C1(n8394), .C2(P2_REG2_REG_12__SCAN_IN), .A(n8392), .B(
        n6684), .ZN(n8390) );
  NAND2_X1 U8322 ( .A1(n6684), .A2(n8390), .ZN(n6686) );
  INV_X1 U8323 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n6948) );
  AOI22_X1 U8324 ( .A1(P2_REG2_REG_13__SCAN_IN), .A2(n6955), .B1(n6697), .B2(
        n6948), .ZN(n6685) );
  NOR2_X1 U8325 ( .A1(n6686), .A2(n6685), .ZN(n6947) );
  AOI21_X1 U8326 ( .B1(n6686), .B2(n6685), .A(n6947), .ZN(n6699) );
  INV_X1 U8327 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9940) );
  MUX2_X1 U8328 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9940), .S(n8394), .Z(n8398)
         );
  OAI21_X1 U8329 ( .B1(n6481), .B2(n6688), .A(n6687), .ZN(n6689) );
  INV_X1 U8330 ( .A(n6689), .ZN(n8397) );
  AOI21_X1 U8331 ( .B1(n9940), .B2(n6690), .A(n8395), .ZN(n6692) );
  INV_X1 U8332 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U8333 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n6955), .B1(n6697), .B2(
        n10183), .ZN(n6691) );
  NOR2_X1 U8334 ( .A1(n6692), .A2(n6691), .ZN(n6954) );
  AOI21_X1 U8335 ( .B1(n6692), .B2(n6691), .A(n6954), .ZN(n6695) );
  NOR2_X1 U8336 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7438), .ZN(n6693) );
  AOI21_X1 U8337 ( .B1(n9707), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n6693), .ZN(
        n6694) );
  OAI21_X1 U8338 ( .B1(n7342), .B2(n6695), .A(n6694), .ZN(n6696) );
  AOI21_X1 U8339 ( .B1(n6697), .B2(n9709), .A(n6696), .ZN(n6698) );
  OAI21_X1 U8340 ( .B1(n6699), .B2(n9686), .A(n6698), .ZN(P2_U3258) );
  OR2_X1 U8341 ( .A1(n6981), .A2(n6985), .ZN(n6839) );
  OR2_X1 U8342 ( .A1(n7065), .A2(n5762), .ZN(n6702) );
  NAND2_X1 U8343 ( .A1(n7150), .A2(n6702), .ZN(n6780) );
  INV_X1 U8344 ( .A(n7147), .ZN(n6715) );
  NOR4_X1 U8345 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6711) );
  NOR4_X1 U8346 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6710) );
  INV_X1 U8347 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9921) );
  INV_X1 U8348 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10093) );
  INV_X1 U8349 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10102) );
  INV_X1 U8350 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10104) );
  NAND4_X1 U8351 ( .A1(n9921), .A2(n10093), .A3(n10102), .A4(n10104), .ZN(
        n6708) );
  NOR4_X1 U8352 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6706) );
  NOR4_X1 U8353 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6705) );
  NOR4_X1 U8354 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6704) );
  NOR4_X1 U8355 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6703) );
  NAND4_X1 U8356 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .ZN(n6707)
         );
  NOR4_X1 U8357 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        n6708), .A4(n6707), .ZN(n6709) );
  AND3_X1 U8358 ( .A1(n6711), .A2(n6710), .A3(n6709), .ZN(n6712) );
  NOR2_X1 U8359 ( .A1(n6713), .A2(n6712), .ZN(n6724) );
  INV_X1 U8360 ( .A(n6724), .ZN(n6714) );
  NAND2_X1 U8361 ( .A1(n6714), .A2(n6725), .ZN(n7148) );
  OR2_X1 U8362 ( .A1(n6715), .A2(n7148), .ZN(n6716) );
  INV_X2 U8363 ( .A(n9674), .ZN(n9675) );
  INV_X1 U8364 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6723) );
  INV_X1 U8365 ( .A(n7206), .ZN(n6717) );
  OR3_X1 U8366 ( .A1(n6718), .A2(n6717), .A3(n7283), .ZN(n6720) );
  INV_X1 U8367 ( .A(n6818), .ZN(n8985) );
  NAND2_X1 U8368 ( .A1(n9305), .A2(n8985), .ZN(n6719) );
  NAND2_X1 U8369 ( .A1(n6720), .A2(n6719), .ZN(n7211) );
  INV_X1 U8370 ( .A(n7211), .ZN(n6721) );
  OAI21_X1 U8371 ( .B1(n7158), .B2(n7206), .A(n6721), .ZN(n6728) );
  NAND2_X1 U8372 ( .A1(n6728), .A2(n9675), .ZN(n6722) );
  OAI21_X1 U8373 ( .B1(n9675), .B2(n6723), .A(n6722), .ZN(P1_U3454) );
  OR2_X1 U8374 ( .A1(n6725), .A2(n6724), .ZN(n6781) );
  INV_X1 U8375 ( .A(n6781), .ZN(n6726) );
  NAND2_X1 U8376 ( .A1(n6726), .A2(n7147), .ZN(n6727) );
  INV_X2 U8377 ( .A(n9680), .ZN(n9683) );
  NAND2_X1 U8378 ( .A1(n6728), .A2(n9683), .ZN(n6729) );
  OAI21_X1 U8379 ( .B1(n9683), .B2(n8988), .A(n6729), .ZN(P1_U3523) );
  NOR2_X1 U8380 ( .A1(n8344), .A2(P2_U3152), .ZN(n6766) );
  INV_X1 U8381 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6736) );
  INV_X1 U8382 ( .A(n8330), .ZN(n8343) );
  INV_X1 U8383 ( .A(n8333), .ZN(n8346) );
  AOI22_X1 U8384 ( .A1(n8343), .A2(n6891), .B1(n8346), .B2(n9772), .ZN(n6735)
         );
  INV_X1 U8385 ( .A(n9779), .ZN(n6733) );
  XOR2_X1 U8386 ( .A(n6731), .B(n6730), .Z(n6732) );
  AOI22_X1 U8387 ( .A1(n6733), .A2(n8336), .B1(n7594), .B2(n6732), .ZN(n6734)
         );
  OAI211_X1 U8388 ( .C1(n6766), .C2(n6736), .A(n6735), .B(n6734), .ZN(P2_U3239) );
  AOI22_X1 U8389 ( .A1(n8343), .A2(n6649), .B1(n8346), .B2(n8372), .ZN(n6742)
         );
  OAI21_X1 U8390 ( .B1(n6739), .B2(n6738), .A(n6737), .ZN(n6740) );
  AOI22_X1 U8391 ( .A1(n6890), .A2(n8336), .B1(n7594), .B2(n6740), .ZN(n6741)
         );
  OAI211_X1 U8392 ( .C1(n6766), .C2(n7005), .A(n6742), .B(n6741), .ZN(P2_U3224) );
  INV_X1 U8393 ( .A(n6743), .ZN(n6776) );
  AOI22_X1 U8394 ( .A1(n7174), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n8758), .ZN(n6744) );
  OAI21_X1 U8395 ( .B1(n6776), .B2(n8769), .A(n6744), .ZN(P2_U3343) );
  INV_X1 U8396 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6901) );
  INV_X1 U8397 ( .A(n9806), .ZN(n8093) );
  INV_X1 U8398 ( .A(n7627), .ZN(n7794) );
  INV_X1 U8399 ( .A(n8371), .ZN(n7036) );
  INV_X1 U8400 ( .A(n8372), .ZN(n6896) );
  OAI22_X1 U8401 ( .A1(n7036), .A2(n9743), .B1(n6896), .B2(n9745), .ZN(n6906)
         );
  NAND2_X1 U8402 ( .A1(n7794), .A2(n6906), .ZN(n6747) );
  OAI211_X1 U8403 ( .C1(n8349), .C2(n8093), .A(n6747), .B(n6746), .ZN(n6748)
         );
  AOI21_X1 U8404 ( .B1(n6901), .B2(n8344), .A(n6748), .ZN(n6749) );
  OAI21_X1 U8405 ( .B1(n6750), .B2(n8340), .A(n6749), .ZN(P2_U3220) );
  XNOR2_X1 U8406 ( .A(n6751), .B(n6752), .ZN(n6757) );
  OAI21_X1 U8407 ( .B1(n8349), .B2(n9821), .A(n6753), .ZN(n6755) );
  OAI22_X1 U8408 ( .A1(n7036), .A2(n8330), .B1(n8333), .B2(n7117), .ZN(n6754)
         );
  AOI211_X1 U8409 ( .C1(n7038), .C2(n8344), .A(n6755), .B(n6754), .ZN(n6756)
         );
  OAI21_X1 U8410 ( .B1(n6757), .B2(n8340), .A(n6756), .ZN(P2_U3229) );
  INV_X1 U8411 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6765) );
  NOR2_X1 U8412 ( .A1(n7627), .A2(n6758), .ZN(n6763) );
  MUX2_X1 U8413 ( .A(n8078), .B(n6760), .S(n6759), .Z(n6761) );
  AOI21_X1 U8414 ( .B1(n7007), .B2(n6761), .A(n8340), .ZN(n6762) );
  AOI211_X1 U8415 ( .C1(n7003), .C2(n8336), .A(n6763), .B(n6762), .ZN(n6764)
         );
  OAI21_X1 U8416 ( .B1(n6766), .B2(n6765), .A(n6764), .ZN(P2_U3234) );
  INV_X1 U8417 ( .A(n6767), .ZN(n6768) );
  AOI21_X1 U8418 ( .B1(n6770), .B2(n6769), .A(n6768), .ZN(n6775) );
  AOI22_X1 U8419 ( .A1(n8343), .A2(n8370), .B1(n8346), .B2(n8368), .ZN(n6774)
         );
  OAI21_X1 U8420 ( .B1(n8349), .B2(n8631), .A(n6771), .ZN(n6772) );
  AOI21_X1 U8421 ( .B1(n8628), .B2(n8344), .A(n6772), .ZN(n6773) );
  OAI211_X1 U8422 ( .C1(n6775), .C2(n8340), .A(n6774), .B(n6773), .ZN(P2_U3241) );
  OAI222_X1 U8423 ( .A1(n9468), .A2(n6777), .B1(n9466), .B2(n6776), .C1(
        P1_U3084), .C2(n9017), .ZN(P1_U3338) );
  NAND2_X1 U8424 ( .A1(n8354), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6778) );
  OAI21_X1 U8425 ( .B1(n8438), .B2(n8354), .A(n6778), .ZN(P2_U3581) );
  NOR2_X1 U8426 ( .A1(n6781), .A2(n7147), .ZN(n6779) );
  OR2_X1 U8427 ( .A1(n6780), .A2(n6779), .ZN(n6842) );
  AND2_X1 U8428 ( .A1(n6842), .A2(n7150), .ZN(n6885) );
  NOR2_X1 U8429 ( .A1(n6782), .A2(n6781), .ZN(n6797) );
  NAND3_X1 U8430 ( .A1(n6797), .A2(n9666), .A3(n6981), .ZN(n8969) );
  AND2_X2 U8431 ( .A1(n6784), .A2(n6785), .ZN(n6825) );
  AOI21_X1 U8432 ( .B1(n6791), .B2(n6828), .A(n6787), .ZN(n6794) );
  NAND2_X1 U8433 ( .A1(n6788), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6789) );
  OAI21_X1 U8434 ( .B1(n4397), .B2(n7158), .A(n6789), .ZN(n6790) );
  INV_X1 U8435 ( .A(n6790), .ZN(n6793) );
  NAND2_X1 U8436 ( .A1(n6791), .A2(n6825), .ZN(n6792) );
  NAND2_X1 U8437 ( .A1(n6793), .A2(n6792), .ZN(n6815) );
  NAND2_X1 U8438 ( .A1(n6815), .A2(n6794), .ZN(n6817) );
  OAI21_X1 U8439 ( .B1(n6794), .B2(n6815), .A(n6817), .ZN(n6849) );
  AND2_X1 U8440 ( .A1(n7283), .A2(n6797), .ZN(n6843) );
  NAND2_X1 U8441 ( .A1(n6795), .A2(n5619), .ZN(n6796) );
  INV_X1 U8442 ( .A(n6797), .ZN(n6798) );
  OR2_X1 U8443 ( .A1(n7206), .A2(n7362), .ZN(n9602) );
  OR2_X1 U8444 ( .A1(n6798), .A2(n9602), .ZN(n6799) );
  NAND2_X1 U8445 ( .A1(n9605), .A2(n6799), .ZN(n8967) );
  OAI22_X1 U8446 ( .A1(n8960), .A2(n6818), .B1(n8954), .B2(n7158), .ZN(n6800)
         );
  AOI21_X1 U8447 ( .B1(n8944), .B2(n6849), .A(n6800), .ZN(n6801) );
  OAI21_X1 U8448 ( .B1(n6885), .B2(n7209), .A(n6801), .ZN(P1_U3230) );
  NOR2_X1 U8449 ( .A1(n6803), .A2(n6802), .ZN(n6808) );
  NAND2_X1 U8450 ( .A1(n6808), .A2(n6804), .ZN(n6805) );
  NOR2_X1 U8451 ( .A1(n6806), .A2(n4394), .ZN(n6807) );
  AND2_X1 U8452 ( .A1(n6808), .A2(n6807), .ZN(n9734) );
  INV_X1 U8453 ( .A(n9761), .ZN(n8562) );
  NAND2_X1 U8454 ( .A1(n9785), .A2(n6809), .ZN(n9757) );
  NAND2_X1 U8455 ( .A1(n8562), .A2(n9757), .ZN(n9783) );
  NAND2_X1 U8456 ( .A1(n9783), .A2(n7003), .ZN(n6812) );
  INV_X1 U8457 ( .A(n9750), .ZN(n9776) );
  AOI22_X1 U8458 ( .A1(n9785), .A2(n6810), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n9776), .ZN(n6811) );
  OAI211_X1 U8459 ( .C1(n6813), .C2(n9785), .A(n6812), .B(n6811), .ZN(P2_U3296) );
  AND2_X4 U8460 ( .A1(n7151), .A2(n6984), .ZN(n7955) );
  NAND2_X1 U8461 ( .A1(n6817), .A2(n6816), .ZN(n6823) );
  INV_X1 U8462 ( .A(n6823), .ZN(n6821) );
  INV_X2 U8463 ( .A(n6825), .ZN(n7848) );
  XNOR2_X1 U8464 ( .A(n6819), .B(n7955), .ZN(n6822) );
  INV_X1 U8465 ( .A(n6822), .ZN(n6820) );
  NAND2_X1 U8466 ( .A1(n6821), .A2(n6820), .ZN(n6881) );
  AOI22_X1 U8467 ( .A1(n7994), .A2(n8985), .B1(n7990), .B2(n7162), .ZN(n6884)
         );
  NAND2_X1 U8468 ( .A1(n6881), .A2(n6884), .ZN(n6824) );
  NAND2_X1 U8469 ( .A1(n6823), .A2(n6822), .ZN(n6882) );
  NAND2_X1 U8470 ( .A1(n6824), .A2(n6882), .ZN(n6874) );
  OAI22_X1 U8471 ( .A1(n6826), .A2(n7848), .B1(n9649), .B2(n6832), .ZN(n6827)
         );
  XNOR2_X1 U8472 ( .A(n6827), .B(n7955), .ZN(n6830) );
  AOI22_X1 U8473 ( .A1(n6828), .A2(n8984), .B1(n7990), .B2(n7305), .ZN(n6829)
         );
  NAND2_X1 U8474 ( .A1(n6830), .A2(n6829), .ZN(n6831) );
  OAI22_X1 U8475 ( .A1(n7848), .A2(n7297), .B1(n7838), .B2(n6832), .ZN(n6833)
         );
  XNOR2_X1 U8476 ( .A(n6833), .B(n7955), .ZN(n6835) );
  INV_X1 U8477 ( .A(n7297), .ZN(n8983) );
  AOI22_X1 U8478 ( .A1(n7994), .A2(n8983), .B1(n7990), .B2(n6973), .ZN(n6834)
         );
  AND2_X1 U8479 ( .A1(n6835), .A2(n6834), .ZN(n6992) );
  INV_X1 U8480 ( .A(n6992), .ZN(n6836) );
  OR2_X1 U8481 ( .A1(n6835), .A2(n6834), .ZN(n6994) );
  NAND2_X1 U8482 ( .A1(n6836), .A2(n6994), .ZN(n6837) );
  XNOR2_X1 U8483 ( .A(n6993), .B(n6837), .ZN(n6848) );
  NAND2_X1 U8484 ( .A1(n6839), .A2(n6838), .ZN(n6840) );
  NAND2_X1 U8485 ( .A1(n6840), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6841) );
  INV_X1 U8486 ( .A(n8965), .ZN(n8951) );
  INV_X1 U8487 ( .A(n8962), .ZN(n8948) );
  OAI22_X1 U8488 ( .A1(n8948), .A2(n6826), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6844), .ZN(n6846) );
  OAI22_X1 U8489 ( .A1(n8960), .A2(n7068), .B1(n7838), .B2(n8954), .ZN(n6845)
         );
  AOI211_X1 U8490 ( .C1(n6844), .C2(n8951), .A(n6846), .B(n6845), .ZN(n6847)
         );
  OAI21_X1 U8491 ( .B1(n6848), .B2(n8969), .A(n6847), .ZN(P1_U3216) );
  INV_X1 U8492 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6873) );
  INV_X1 U8493 ( .A(n6849), .ZN(n6850) );
  MUX2_X1 U8494 ( .A(n6851), .B(n6850), .S(n5766), .Z(n6855) );
  NOR2_X1 U8495 ( .A1(n5766), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6852) );
  NOR2_X1 U8496 ( .A1(n6852), .A2(n4391), .ZN(n8987) );
  OAI21_X1 U8497 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n8987), .A(P1_U4006), .ZN(
        n6853) );
  AOI21_X1 U8498 ( .B1(n6855), .B2(n6854), .A(n6853), .ZN(n9566) );
  INV_X1 U8499 ( .A(n9566), .ZN(n6872) );
  INV_X1 U8500 ( .A(n9583), .ZN(n6857) );
  INV_X1 U8501 ( .A(n6861), .ZN(n6856) );
  INV_X1 U8502 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U8503 ( .A1(n6857), .A2(n6856), .B1(P1_U3084), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n6870) );
  OAI211_X1 U8504 ( .C1(n6860), .C2(n6859), .A(n9575), .B(n6858), .ZN(n6869)
         );
  MUX2_X1 U8505 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6335), .S(n6861), .Z(n6864)
         );
  INV_X1 U8506 ( .A(n6862), .ZN(n6863) );
  NAND2_X1 U8507 ( .A1(n6864), .A2(n6863), .ZN(n6866) );
  OAI211_X1 U8508 ( .C1(n6867), .C2(n6866), .A(n9597), .B(n6865), .ZN(n6868)
         );
  AND3_X1 U8509 ( .A1(n6870), .A2(n6869), .A3(n6868), .ZN(n6871) );
  OAI211_X1 U8510 ( .C1(n6873), .C2(n9586), .A(n6872), .B(n6871), .ZN(P1_U3243) );
  OAI21_X1 U8511 ( .B1(n6876), .B2(n6874), .A(n6875), .ZN(n6877) );
  NAND2_X1 U8512 ( .A1(n6877), .A2(n8944), .ZN(n6880) );
  OAI22_X1 U8513 ( .A1(n6818), .A2(n8948), .B1(n8960), .B2(n7297), .ZN(n6878)
         );
  AOI21_X1 U8514 ( .B1(n7305), .B2(n8967), .A(n6878), .ZN(n6879) );
  OAI211_X1 U8515 ( .C1(n6885), .C2(n10193), .A(n6880), .B(n6879), .ZN(
        P1_U3235) );
  NAND2_X1 U8516 ( .A1(n6881), .A2(n6882), .ZN(n6883) );
  XNOR2_X1 U8517 ( .A(n6884), .B(n6883), .ZN(n6889) );
  NOR2_X1 U8518 ( .A1(n6885), .A2(n7159), .ZN(n6887) );
  OAI22_X1 U8519 ( .A1(n4827), .A2(n8948), .B1(n8960), .B2(n6826), .ZN(n6886)
         );
  AOI211_X1 U8520 ( .C1(n7162), .C2(n8967), .A(n6887), .B(n6886), .ZN(n6888)
         );
  OAI21_X1 U8521 ( .B1(n6889), .B2(n8969), .A(n6888), .ZN(P1_U3220) );
  NAND2_X1 U8522 ( .A1(n9785), .A2(n9859), .ZN(n9755) );
  INV_X1 U8523 ( .A(n9755), .ZN(n9782) );
  INV_X1 U8524 ( .A(n8086), .ZN(n7013) );
  NAND2_X1 U8525 ( .A1(n7008), .A2(n7002), .ZN(n6895) );
  NAND2_X1 U8526 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  OR2_X1 U8527 ( .A1(n8372), .A2(n9779), .ZN(n8081) );
  NAND2_X1 U8528 ( .A1(n8372), .A2(n9779), .ZN(n8079) );
  NAND2_X1 U8529 ( .A1(n9781), .A2(n6904), .ZN(n6898) );
  NAND2_X1 U8530 ( .A1(n6896), .A2(n9779), .ZN(n6897) );
  NAND2_X1 U8531 ( .A1(n6898), .A2(n6897), .ZN(n7014) );
  XNOR2_X1 U8532 ( .A(n7013), .B(n7014), .ZN(n9811) );
  NAND2_X1 U8533 ( .A1(n6899), .A2(n9806), .ZN(n6900) );
  AND2_X1 U8534 ( .A1(n9758), .A2(n6900), .ZN(n9807) );
  AOI22_X1 U8535 ( .A1(n9761), .A2(n9807), .B1(n9776), .B2(n6901), .ZN(n6902)
         );
  OAI21_X1 U8536 ( .B1(n8093), .B2(n9757), .A(n6902), .ZN(n6903) );
  AOI21_X1 U8537 ( .B1(n9782), .B2(n9811), .A(n6903), .ZN(n6910) );
  NAND2_X1 U8538 ( .A1(n6905), .A2(n8086), .ZN(n7020) );
  OAI21_X1 U8539 ( .B1(n6905), .B2(n8086), .A(n7020), .ZN(n6907) );
  AOI21_X1 U8540 ( .B1(n6907), .B2(n9774), .A(n6906), .ZN(n9809) );
  MUX2_X1 U8541 ( .A(n6908), .B(n9809), .S(n9785), .Z(n6909) );
  NAND2_X1 U8542 ( .A1(n6910), .A2(n6909), .ZN(P2_U3293) );
  INV_X1 U8543 ( .A(n6911), .ZN(n6964) );
  AOI22_X1 U8544 ( .A1(n9050), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7078), .ZN(n6912) );
  OAI21_X1 U8545 ( .B1(n6964), .B2(n9466), .A(n6912), .ZN(P1_U3336) );
  OAI21_X1 U8546 ( .B1(n6915), .B2(n6914), .A(n6913), .ZN(n6924) );
  NAND2_X1 U8547 ( .A1(n9022), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U8548 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n6916) );
  OAI211_X1 U8549 ( .C1(n9583), .C2(n6918), .A(n6917), .B(n6916), .ZN(n6923)
         );
  AOI211_X1 U8550 ( .C1(n6921), .C2(n6920), .A(n6919), .B(n9591), .ZN(n6922)
         );
  AOI211_X1 U8551 ( .C1(n9597), .C2(n6924), .A(n6923), .B(n6922), .ZN(n6925)
         );
  INV_X1 U8552 ( .A(n6925), .ZN(P1_U3253) );
  XNOR2_X1 U8553 ( .A(n6927), .B(n6926), .ZN(n6931) );
  INV_X1 U8554 ( .A(n7224), .ZN(n8366) );
  AOI22_X1 U8555 ( .A1(n8343), .A2(n8368), .B1(n8346), .B2(n8366), .ZN(n6930)
         );
  INV_X1 U8556 ( .A(n7226), .ZN(n9832) );
  NAND2_X1 U8557 ( .A1(P2_U3152), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n9692) );
  OAI21_X1 U8558 ( .B1(n8349), .B2(n9832), .A(n9692), .ZN(n6928) );
  AOI21_X1 U8559 ( .B1(n7125), .B2(n8344), .A(n6928), .ZN(n6929) );
  OAI211_X1 U8560 ( .C1(n6931), .C2(n8340), .A(n6930), .B(n6929), .ZN(P2_U3223) );
  INV_X1 U8561 ( .A(n6932), .ZN(n6935) );
  INV_X1 U8562 ( .A(n9034), .ZN(n9025) );
  OAI222_X1 U8563 ( .A1(n9468), .A2(n6933), .B1(n9473), .B2(n6935), .C1(n9025), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  OAI222_X1 U8564 ( .A1(P2_U3152), .A2(n7337), .B1(n8769), .B2(n6935), .C1(
        n6934), .C2(n8771), .ZN(P2_U3342) );
  OR2_X1 U8565 ( .A1(n7117), .A2(n9745), .ZN(n6937) );
  OR2_X1 U8566 ( .A1(n7225), .A2(n9743), .ZN(n6936) );
  NAND2_X1 U8567 ( .A1(n6937), .A2(n6936), .ZN(n9722) );
  INV_X1 U8568 ( .A(n9722), .ZN(n6940) );
  NAND2_X1 U8569 ( .A1(n8336), .A2(n9727), .ZN(n6939) );
  OAI211_X1 U8570 ( .C1(n6940), .C2(n7627), .A(n6939), .B(n6938), .ZN(n6945)
         );
  XNOR2_X1 U8571 ( .A(n6942), .B(n6941), .ZN(n6943) );
  NOR2_X1 U8572 ( .A1(n6943), .A2(n8340), .ZN(n6944) );
  AOI211_X1 U8573 ( .C1(n9725), .C2(n8344), .A(n6945), .B(n6944), .ZN(n6946)
         );
  INV_X1 U8574 ( .A(n6946), .ZN(P2_U3215) );
  INV_X1 U8575 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6949) );
  AOI22_X1 U8576 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7051), .B1(n7046), .B2(
        n6949), .ZN(n6950) );
  NOR2_X1 U8577 ( .A1(n6951), .A2(n6950), .ZN(n7047) );
  AOI21_X1 U8578 ( .B1(n6951), .B2(n6950), .A(n7047), .ZN(n6962) );
  INV_X1 U8579 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6953) );
  NOR2_X1 U8580 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6047), .ZN(n7599) );
  INV_X1 U8581 ( .A(n7599), .ZN(n6952) );
  OAI21_X1 U8582 ( .B1(n8419), .B2(n6953), .A(n6952), .ZN(n6960) );
  AOI21_X1 U8583 ( .B1(n10183), .B2(n6955), .A(n6954), .ZN(n6957) );
  INV_X1 U8584 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9523) );
  AOI22_X1 U8585 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n7051), .B1(n7046), .B2(
        n9523), .ZN(n6956) );
  NOR2_X1 U8586 ( .A1(n6957), .A2(n6956), .ZN(n7050) );
  AOI21_X1 U8587 ( .B1(n6957), .B2(n6956), .A(n7050), .ZN(n6958) );
  NOR2_X1 U8588 ( .A1(n6958), .A2(n7342), .ZN(n6959) );
  AOI211_X1 U8589 ( .C1(n9709), .C2(n7046), .A(n6960), .B(n6959), .ZN(n6961)
         );
  OAI21_X1 U8590 ( .B1(n6962), .B2(n9686), .A(n6961), .ZN(P2_U3259) );
  OAI222_X1 U8591 ( .A1(P2_U3152), .A2(n7580), .B1(n8769), .B2(n6964), .C1(
        n6963), .C2(n8771), .ZN(P2_U3341) );
  INV_X1 U8592 ( .A(n7065), .ZN(n9673) );
  NAND2_X1 U8593 ( .A1(n7146), .A2(n6965), .ZN(n7145) );
  OR2_X1 U8594 ( .A1(n6818), .A2(n9645), .ZN(n6966) );
  NAND2_X1 U8595 ( .A1(n7145), .A2(n6966), .ZN(n7294) );
  INV_X1 U8596 ( .A(n7294), .ZN(n6968) );
  INV_X1 U8597 ( .A(n7293), .ZN(n6967) );
  NAND2_X1 U8598 ( .A1(n6968), .A2(n6967), .ZN(n7296) );
  NAND2_X1 U8599 ( .A1(n6826), .A2(n9649), .ZN(n6969) );
  NAND2_X1 U8600 ( .A1(n7296), .A2(n6969), .ZN(n6971) );
  NAND2_X1 U8601 ( .A1(n6971), .A2(n6970), .ZN(n7060) );
  OR2_X1 U8602 ( .A1(n6971), .A2(n6970), .ZN(n6972) );
  NAND2_X1 U8603 ( .A1(n7060), .A2(n6972), .ZN(n7837) );
  NAND2_X1 U8604 ( .A1(n7158), .A2(n9645), .ZN(n7301) );
  AND2_X1 U8605 ( .A1(n7303), .A2(n6973), .ZN(n6974) );
  OR2_X1 U8606 ( .A1(n6974), .A2(n7260), .ZN(n7842) );
  OR2_X1 U8607 ( .A1(n7206), .A2(n6700), .ZN(n9668) );
  OAI22_X1 U8608 ( .A1(n7842), .A2(n9668), .B1(n7838), .B2(n9666), .ZN(n6990)
         );
  OAI21_X1 U8609 ( .B1(n6977), .B2(n6976), .A(n6975), .ZN(n6983) );
  NAND2_X1 U8610 ( .A1(n5762), .A2(n6700), .ZN(n6979) );
  OAI22_X1 U8611 ( .A1(n7068), .A2(n9492), .B1(n9491), .B2(n6826), .ZN(n6982)
         );
  AOI21_X1 U8612 ( .B1(n6983), .B2(n9308), .A(n6982), .ZN(n6989) );
  OR2_X1 U8613 ( .A1(n6984), .A2(n6784), .ZN(n6987) );
  AND2_X1 U8614 ( .A1(n6987), .A2(n6986), .ZN(n7645) );
  INV_X1 U8615 ( .A(n7645), .ZN(n9496) );
  NAND2_X1 U8616 ( .A1(n7837), .A2(n9496), .ZN(n6988) );
  NAND2_X1 U8617 ( .A1(n6989), .A2(n6988), .ZN(n7836) );
  AOI211_X1 U8618 ( .C1(n9673), .C2(n7837), .A(n6990), .B(n7836), .ZN(n7044)
         );
  NAND2_X1 U8619 ( .A1(n9680), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6991) );
  OAI21_X1 U8620 ( .B1(n7044), .B2(n9680), .A(n6991), .ZN(P1_U3526) );
  OAI22_X1 U8621 ( .A1(n7068), .A2(n7848), .B1(n9654), .B2(n6832), .ZN(n6995)
         );
  XNOR2_X1 U8622 ( .A(n6995), .B(n7992), .ZN(n7131) );
  INV_X1 U8623 ( .A(n7068), .ZN(n8982) );
  AOI22_X1 U8624 ( .A1(n7994), .A2(n8982), .B1(n7990), .B2(n7265), .ZN(n7132)
         );
  XNOR2_X1 U8625 ( .A(n7131), .B(n7132), .ZN(n6997) );
  NAND2_X1 U8626 ( .A1(n6996), .A2(n6997), .ZN(n7135) );
  OAI211_X1 U8627 ( .C1(n6996), .C2(n6997), .A(n7135), .B(n8944), .ZN(n7001)
         );
  NAND2_X1 U8628 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n9556) );
  INV_X1 U8629 ( .A(n9556), .ZN(n6999) );
  OAI22_X1 U8630 ( .A1(n8960), .A2(n7315), .B1(n9654), .B2(n8954), .ZN(n6998)
         );
  AOI211_X1 U8631 ( .C1(n8962), .C2(n8983), .A(n6999), .B(n6998), .ZN(n7000)
         );
  OAI211_X1 U8632 ( .C1(n8965), .C2(n7263), .A(n7001), .B(n7000), .ZN(P1_U3228) );
  INV_X1 U8633 ( .A(n7008), .ZN(n8042) );
  XNOR2_X1 U8634 ( .A(n8042), .B(n7002), .ZN(n9799) );
  NAND2_X1 U8635 ( .A1(n6890), .A2(n7003), .ZN(n9795) );
  NAND3_X1 U8636 ( .A1(n9761), .A2(n4716), .A3(n9795), .ZN(n7004) );
  OAI21_X1 U8637 ( .B1(n9750), .B2(n7005), .A(n7004), .ZN(n7006) );
  AOI21_X1 U8638 ( .B1(n9726), .B2(n6890), .A(n7006), .ZN(n7012) );
  XNOR2_X1 U8639 ( .A(n7008), .B(n7007), .ZN(n7009) );
  AOI222_X1 U8640 ( .A1(n9774), .A2(n7009), .B1(n8372), .B2(n9771), .C1(n6649), 
        .C2(n9770), .ZN(n9798) );
  MUX2_X1 U8641 ( .A(n7010), .B(n9798), .S(n9785), .Z(n7011) );
  OAI211_X1 U8642 ( .C1(n9799), .C2(n9755), .A(n7012), .B(n7011), .ZN(P2_U3295) );
  INV_X1 U8643 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U8644 ( .A1(n7014), .A2(n7013), .ZN(n7016) );
  NAND2_X1 U8645 ( .A1(n9746), .A2(n8093), .ZN(n7015) );
  NAND2_X1 U8646 ( .A1(n7016), .A2(n7015), .ZN(n9754) );
  OR2_X1 U8647 ( .A1(n8371), .A2(n9756), .ZN(n8068) );
  NAND2_X1 U8648 ( .A1(n8371), .A2(n9756), .ZN(n8091) );
  NAND2_X1 U8649 ( .A1(n8068), .A2(n8091), .ZN(n9738) );
  NAND2_X1 U8650 ( .A1(n9754), .A2(n9738), .ZN(n7018) );
  NAND2_X1 U8651 ( .A1(n7036), .A2(n9756), .ZN(n7017) );
  OR2_X1 U8652 ( .A1(n8370), .A2(n9821), .ZN(n8069) );
  NAND2_X1 U8653 ( .A1(n8370), .A2(n9821), .ZN(n8094) );
  NAND2_X1 U8654 ( .A1(n8069), .A2(n8094), .ZN(n8045) );
  INV_X1 U8655 ( .A(n9821), .ZN(n7041) );
  NAND2_X1 U8656 ( .A1(n7117), .A2(n7115), .ZN(n8101) );
  INV_X1 U8657 ( .A(n7117), .ZN(n8369) );
  NAND2_X1 U8658 ( .A1(n8369), .A2(n8631), .ZN(n8098) );
  XNOR2_X1 U8659 ( .A(n7114), .B(n4804), .ZN(n8630) );
  NOR2_X1 U8660 ( .A1(n9772), .A2(n8093), .ZN(n8065) );
  NOR2_X1 U8661 ( .A1(n9738), .A2(n8065), .ZN(n7019) );
  NAND2_X1 U8662 ( .A1(n7020), .A2(n7019), .ZN(n9737) );
  NAND2_X1 U8663 ( .A1(n9737), .A2(n8091), .ZN(n7032) );
  INV_X1 U8664 ( .A(n7032), .ZN(n7022) );
  NAND2_X1 U8665 ( .A1(n7022), .A2(n7021), .ZN(n7033) );
  NAND2_X1 U8666 ( .A1(n7033), .A2(n8069), .ZN(n7023) );
  OAI21_X1 U8667 ( .B1(n8046), .B2(n7023), .A(n7110), .ZN(n7024) );
  AOI222_X1 U8668 ( .A1(n9774), .A2(n7024), .B1(n8368), .B2(n9771), .C1(n8370), 
        .C2(n9770), .ZN(n8627) );
  NOR2_X1 U8669 ( .A1(n9758), .A2(n9813), .ZN(n9760) );
  NAND2_X1 U8670 ( .A1(n7030), .A2(n8631), .ZN(n9730) );
  OR2_X1 U8671 ( .A1(n7030), .A2(n8631), .ZN(n7025) );
  AND2_X1 U8672 ( .A1(n9730), .A2(n7025), .ZN(n8629) );
  AOI22_X1 U8673 ( .A1(n8629), .A2(n9845), .B1(n9844), .B2(n7115), .ZN(n7026)
         );
  OAI211_X1 U8674 ( .C1(n9848), .C2(n8630), .A(n8627), .B(n7026), .ZN(n7028)
         );
  NAND2_X1 U8675 ( .A1(n7028), .A2(n9861), .ZN(n7027) );
  OAI21_X1 U8676 ( .B1(n9861), .B2(n9985), .A(n7027), .ZN(P2_U3469) );
  NAND2_X1 U8677 ( .A1(n7028), .A2(n9879), .ZN(n7029) );
  OAI21_X1 U8678 ( .B1(n9879), .B2(n6468), .A(n7029), .ZN(P2_U3526) );
  INV_X1 U8679 ( .A(n7030), .ZN(n7031) );
  OAI211_X1 U8680 ( .C1(n9821), .C2(n9760), .A(n7031), .B(n9845), .ZN(n9820)
         );
  NOR2_X1 U8681 ( .A1(n9820), .A2(n4394), .ZN(n7037) );
  INV_X1 U8682 ( .A(n7033), .ZN(n7034) );
  AOI21_X1 U8683 ( .B1(n8045), .B2(n7032), .A(n7034), .ZN(n7035) );
  OAI222_X1 U8684 ( .A1(n9743), .A2(n7117), .B1(n9745), .B2(n7036), .C1(n9740), 
        .C2(n7035), .ZN(n9822) );
  AOI211_X1 U8685 ( .C1(n9776), .C2(n7038), .A(n7037), .B(n9822), .ZN(n7039)
         );
  MUX2_X1 U8686 ( .A(n10153), .B(n7039), .S(n9785), .Z(n7043) );
  XNOR2_X1 U8687 ( .A(n7040), .B(n8045), .ZN(n9824) );
  AOI22_X1 U8688 ( .A1(n9782), .A2(n9824), .B1(n9726), .B2(n7041), .ZN(n7042)
         );
  NAND2_X1 U8689 ( .A1(n7043), .A2(n7042), .ZN(P2_U3291) );
  OR2_X1 U8690 ( .A1(n7044), .A2(n9674), .ZN(n7045) );
  OAI21_X1 U8691 ( .B1(n9675), .B2(n5455), .A(n7045), .ZN(P1_U3463) );
  NOR2_X1 U8692 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n7046), .ZN(n7048) );
  XNOR2_X1 U8693 ( .A(n7174), .B(n7173), .ZN(n7049) );
  NOR2_X1 U8694 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7049), .ZN(n7175) );
  AOI21_X1 U8695 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n7049), .A(n7175), .ZN(
        n7058) );
  AOI21_X1 U8696 ( .B1(n9523), .B2(n7051), .A(n7050), .ZN(n7166) );
  XOR2_X1 U8697 ( .A(n7174), .B(n7166), .Z(n7052) );
  NAND2_X1 U8698 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7052), .ZN(n7167) );
  OAI211_X1 U8699 ( .C1(n7052), .C2(P2_REG1_REG_15__SCAN_IN), .A(n9711), .B(
        n7167), .ZN(n7057) );
  INV_X1 U8700 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7054) );
  OR2_X1 U8701 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7626), .ZN(n7053) );
  OAI21_X1 U8702 ( .B1(n8419), .B2(n7054), .A(n7053), .ZN(n7055) );
  AOI21_X1 U8703 ( .B1(n9709), .B2(n7174), .A(n7055), .ZN(n7056) );
  OAI211_X1 U8704 ( .C1(n7058), .C2(n9686), .A(n7057), .B(n7056), .ZN(P2_U3260) );
  INV_X1 U8705 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7074) );
  NAND2_X1 U8706 ( .A1(n7297), .A2(n7838), .ZN(n7059) );
  NAND2_X1 U8707 ( .A1(n7060), .A2(n7059), .ZN(n7257) );
  NAND2_X1 U8708 ( .A1(n7068), .A2(n9654), .ZN(n7061) );
  NAND2_X1 U8709 ( .A1(n7063), .A2(n7066), .ZN(n7064) );
  NAND2_X1 U8710 ( .A1(n7278), .A2(n7064), .ZN(n9612) );
  NAND2_X1 U8711 ( .A1(n7645), .A2(n7065), .ZN(n9528) );
  XNOR2_X1 U8712 ( .A(n7067), .B(n7062), .ZN(n7070) );
  OAI22_X1 U8713 ( .A1(n7068), .A2(n9491), .B1(n9492), .B2(n7378), .ZN(n7069)
         );
  AOI21_X1 U8714 ( .B1(n7070), .B2(n9308), .A(n7069), .ZN(n9610) );
  INV_X1 U8715 ( .A(n9666), .ZN(n9432) );
  NAND2_X1 U8716 ( .A1(n7260), .A2(n9654), .ZN(n7262) );
  AOI21_X1 U8717 ( .B1(n7262), .B2(n7137), .A(n9668), .ZN(n7071) );
  AND2_X1 U8718 ( .A1(n7071), .A2(n7321), .ZN(n9608) );
  AOI21_X1 U8719 ( .B1(n9432), .B2(n7137), .A(n9608), .ZN(n7072) );
  OAI211_X1 U8720 ( .C1(n9612), .C2(n9434), .A(n9610), .B(n7072), .ZN(n7075)
         );
  NAND2_X1 U8721 ( .A1(n7075), .A2(n9675), .ZN(n7073) );
  OAI21_X1 U8722 ( .B1(n9675), .B2(n7074), .A(n7073), .ZN(P1_U3469) );
  NAND2_X1 U8723 ( .A1(n7075), .A2(n9683), .ZN(n7076) );
  OAI21_X1 U8724 ( .B1(n9683), .B2(n6339), .A(n7076), .ZN(P1_U3528) );
  INV_X1 U8725 ( .A(n7077), .ZN(n7109) );
  AOI22_X1 U8726 ( .A1(n9062), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7078), .ZN(n7079) );
  OAI21_X1 U8727 ( .B1(n7109), .B2(n9473), .A(n7079), .ZN(P1_U3335) );
  INV_X1 U8728 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7092) );
  OAI21_X1 U8729 ( .B1(n7082), .B2(n7081), .A(n7080), .ZN(n7090) );
  INV_X1 U8730 ( .A(n7083), .ZN(n7084) );
  NAND2_X1 U8731 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3084), .ZN(n8905) );
  OAI21_X1 U8732 ( .B1(n9583), .B2(n7084), .A(n8905), .ZN(n7089) );
  AOI211_X1 U8733 ( .C1(n7087), .C2(n7086), .A(n7085), .B(n9591), .ZN(n7088)
         );
  AOI211_X1 U8734 ( .C1(n9597), .C2(n7090), .A(n7089), .B(n7088), .ZN(n7091)
         );
  OAI21_X1 U8735 ( .B1(n9586), .B2(n7092), .A(n7091), .ZN(P1_U3254) );
  INV_X1 U8736 ( .A(n7093), .ZN(n7094) );
  AOI21_X1 U8737 ( .B1(n7096), .B2(n7095), .A(n7094), .ZN(n7101) );
  INV_X1 U8738 ( .A(n7346), .ZN(n7251) );
  OAI21_X1 U8739 ( .B1(n8349), .B2(n7251), .A(n7097), .ZN(n7099) );
  OAI22_X1 U8740 ( .A1(n7225), .A2(n8330), .B1(n8333), .B2(n7446), .ZN(n7098)
         );
  AOI211_X1 U8741 ( .C1(n7243), .C2(n8344), .A(n7099), .B(n7098), .ZN(n7100)
         );
  OAI21_X1 U8742 ( .B1(n7101), .B2(n8340), .A(n7100), .ZN(P2_U3233) );
  XNOR2_X1 U8743 ( .A(n7103), .B(n7102), .ZN(n7107) );
  INV_X1 U8744 ( .A(n7451), .ZN(n9837) );
  NAND2_X1 U8745 ( .A1(P2_U3152), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9705) );
  OAI21_X1 U8746 ( .B1(n8349), .B2(n9837), .A(n9705), .ZN(n7105) );
  INV_X1 U8747 ( .A(n8364), .ZN(n7444) );
  OAI22_X1 U8748 ( .A1(n7224), .A2(n8330), .B1(n8333), .B2(n7444), .ZN(n7104)
         );
  AOI211_X1 U8749 ( .C1(n7354), .C2(n8344), .A(n7105), .B(n7104), .ZN(n7106)
         );
  OAI21_X1 U8750 ( .B1(n7107), .B2(n8340), .A(n7106), .ZN(P2_U3219) );
  INV_X1 U8751 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10090) );
  INV_X1 U8752 ( .A(n7588), .ZN(n7108) );
  OAI222_X1 U8753 ( .A1(n8771), .A2(n10090), .B1(n8769), .B2(n7109), .C1(
        P2_U3152), .C2(n7108), .ZN(P2_U3340) );
  OR2_X1 U8754 ( .A1(n7226), .A2(n7225), .ZN(n8108) );
  NAND2_X1 U8755 ( .A1(n7226), .A2(n7225), .ZN(n8109) );
  NAND2_X1 U8756 ( .A1(n8108), .A2(n8109), .ZN(n8102) );
  XNOR2_X1 U8757 ( .A(n9727), .B(n8368), .ZN(n8100) );
  INV_X1 U8758 ( .A(n9727), .ZN(n9828) );
  INV_X1 U8759 ( .A(n7113), .ZN(n7112) );
  NAND2_X1 U8760 ( .A1(n7112), .A2(n7111), .ZN(n7234) );
  INV_X1 U8761 ( .A(n7234), .ZN(n7233) );
  AOI21_X1 U8762 ( .B1(n8102), .B2(n7113), .A(n7233), .ZN(n7124) );
  AOI22_X1 U8763 ( .A1(n8366), .A2(n9771), .B1(n9770), .B2(n8368), .ZN(n7123)
         );
  NAND2_X1 U8764 ( .A1(n7116), .A2(n4416), .ZN(n7119) );
  NAND2_X1 U8765 ( .A1(n7117), .A2(n8631), .ZN(n7118) );
  INV_X1 U8766 ( .A(n8100), .ZN(n9728) );
  NOR2_X1 U8767 ( .A1(n9727), .A2(n8368), .ZN(n7120) );
  OAI211_X1 U8768 ( .C1(n7121), .C2(n8102), .A(n7228), .B(n9859), .ZN(n7122)
         );
  OAI211_X1 U8769 ( .C1(n7124), .C2(n9740), .A(n7123), .B(n7122), .ZN(n9833)
         );
  NAND2_X1 U8770 ( .A1(n9833), .A2(n9785), .ZN(n7130) );
  AOI21_X1 U8771 ( .B1(n7226), .B2(n9731), .A(n7241), .ZN(n9835) );
  INV_X1 U8772 ( .A(n7125), .ZN(n7126) );
  OAI22_X1 U8773 ( .A1(n9785), .A2(n7127), .B1(n7126), .B2(n9750), .ZN(n7128)
         );
  AOI21_X1 U8774 ( .B1(n9835), .B2(n9761), .A(n7128), .ZN(n7129) );
  OAI211_X1 U8775 ( .C1(n9832), .C2(n9757), .A(n7130), .B(n7129), .ZN(P2_U3288) );
  INV_X1 U8776 ( .A(n7131), .ZN(n7133) );
  OR2_X1 U8777 ( .A1(n7133), .A2(n7132), .ZN(n7134) );
  NAND2_X1 U8778 ( .A1(n7135), .A2(n7134), .ZN(n7190) );
  OAI22_X1 U8779 ( .A1(n7315), .A2(n7848), .B1(n9603), .B2(n6832), .ZN(n7136)
         );
  XNOR2_X1 U8780 ( .A(n7136), .B(n7955), .ZN(n7191) );
  XNOR2_X1 U8781 ( .A(n7190), .B(n7191), .ZN(n7139) );
  INV_X1 U8782 ( .A(n7315), .ZN(n8981) );
  AOI22_X1 U8783 ( .A1(n7994), .A2(n8981), .B1(n7990), .B2(n7137), .ZN(n7138)
         );
  OAI21_X1 U8784 ( .B1(n7139), .B2(n7138), .A(n7194), .ZN(n7140) );
  NAND2_X1 U8785 ( .A1(n7140), .A2(n8944), .ZN(n7144) );
  NAND2_X1 U8786 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3084), .ZN(n9581) );
  INV_X1 U8787 ( .A(n9581), .ZN(n7142) );
  OAI22_X1 U8788 ( .A1(n8960), .A2(n7378), .B1(n9603), .B2(n8954), .ZN(n7141)
         );
  AOI211_X1 U8789 ( .C1(n8962), .C2(n8982), .A(n7142), .B(n7141), .ZN(n7143)
         );
  OAI211_X1 U8790 ( .C1(n8965), .C2(n9604), .A(n7144), .B(n7143), .ZN(P1_U3225) );
  OAI21_X1 U8791 ( .B1(n7154), .B2(n7146), .A(n7145), .ZN(n7165) );
  NOR2_X1 U8792 ( .A1(n7148), .A2(n7147), .ZN(n7149) );
  NAND2_X1 U8793 ( .A1(n7150), .A2(n7149), .ZN(n7287) );
  NOR2_X1 U8794 ( .A1(n7151), .A2(n9607), .ZN(n7152) );
  AND2_X1 U8795 ( .A1(n9614), .A2(n7152), .ZN(n9508) );
  INV_X1 U8796 ( .A(n9508), .ZN(n7653) );
  XNOR2_X1 U8797 ( .A(n7154), .B(n7153), .ZN(n7157) );
  INV_X1 U8798 ( .A(n7165), .ZN(n9648) );
  OAI22_X1 U8799 ( .A1(n4827), .A2(n9491), .B1(n9492), .B2(n6826), .ZN(n7155)
         );
  AOI21_X1 U8800 ( .B1(n9648), .B2(n9496), .A(n7155), .ZN(n7156) );
  OAI21_X1 U8801 ( .B1(n9488), .B2(n7157), .A(n7156), .ZN(n9646) );
  OAI211_X1 U8802 ( .C1(n9645), .C2(n7158), .A(n9503), .B(n7301), .ZN(n9644)
         );
  OAI22_X1 U8803 ( .A1(n9644), .A2(n9214), .B1(n9605), .B2(n7159), .ZN(n7160)
         );
  OAI21_X1 U8804 ( .B1(n9646), .B2(n7160), .A(n9614), .ZN(n7164) );
  INV_X1 U8805 ( .A(n9602), .ZN(n7161) );
  NAND2_X1 U8806 ( .A1(n9614), .A2(n7161), .ZN(n9338) );
  AOI22_X1 U8807 ( .A1(n9500), .A2(n7162), .B1(n4393), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7163) );
  OAI211_X1 U8808 ( .C1(n7165), .C2(n7653), .A(n7164), .B(n7163), .ZN(P1_U3290) );
  NAND2_X1 U8809 ( .A1(n7174), .A2(n7166), .ZN(n7168) );
  NAND2_X1 U8810 ( .A1(n7168), .A2(n7167), .ZN(n7170) );
  INV_X1 U8811 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8711) );
  NAND2_X1 U8812 ( .A1(n7337), .A2(n8711), .ZN(n7330) );
  OAI21_X1 U8813 ( .B1(n7337), .B2(n8711), .A(n7330), .ZN(n7169) );
  NOR2_X1 U8814 ( .A1(n7170), .A2(n7169), .ZN(n7332) );
  AOI21_X1 U8815 ( .B1(n7170), .B2(n7169), .A(n7332), .ZN(n7185) );
  AND2_X1 U8816 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7172) );
  NOR2_X1 U8817 ( .A1(n9685), .A2(n7337), .ZN(n7171) );
  AOI211_X1 U8818 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n9707), .A(n7172), .B(
        n7171), .ZN(n7184) );
  NOR2_X1 U8819 ( .A1(n7174), .A2(n7173), .ZN(n7176) );
  NOR2_X1 U8820 ( .A1(n7176), .A2(n7175), .ZN(n7182) );
  INV_X1 U8821 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U8822 ( .A1(n7178), .A2(n7179), .ZN(n7177) );
  OAI21_X1 U8823 ( .B1(n7178), .B2(n7179), .A(n7177), .ZN(n7181) );
  NAND2_X1 U8824 ( .A1(n7337), .A2(n7179), .ZN(n7180) );
  OAI211_X1 U8825 ( .C1(n7182), .C2(n7181), .A(n7336), .B(n9715), .ZN(n7183)
         );
  OAI211_X1 U8826 ( .C1(n7185), .C2(n7342), .A(n7184), .B(n7183), .ZN(P2_U3261) );
  INV_X1 U8827 ( .A(n7186), .ZN(n7188) );
  OAI222_X1 U8828 ( .A1(n8771), .A2(n7187), .B1(n8769), .B2(n7188), .C1(
        P2_U3152), .C2(n4504), .ZN(P2_U3339) );
  OAI222_X1 U8829 ( .A1(n9479), .A2(n7189), .B1(n9473), .B2(n7188), .C1(n9607), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  INV_X1 U8830 ( .A(n7190), .ZN(n7192) );
  NAND2_X1 U8831 ( .A1(n7192), .A2(n7191), .ZN(n7193) );
  OAI22_X1 U8832 ( .A1(n7378), .A2(n7848), .B1(n9660), .B2(n6832), .ZN(n7195)
         );
  XNOR2_X1 U8833 ( .A(n7195), .B(n7955), .ZN(n7367) );
  OR2_X1 U8834 ( .A1(n7963), .A2(n7378), .ZN(n7197) );
  INV_X2 U8835 ( .A(n7848), .ZN(n7995) );
  NAND2_X1 U8836 ( .A1(n7995), .A2(n7326), .ZN(n7196) );
  XNOR2_X1 U8837 ( .A(n7367), .B(n7368), .ZN(n7198) );
  XNOR2_X1 U8838 ( .A(n7373), .B(n7198), .ZN(n7204) );
  INV_X1 U8839 ( .A(n7319), .ZN(n7202) );
  INV_X1 U8840 ( .A(n7423), .ZN(n8979) );
  AOI22_X1 U8841 ( .A1(n8921), .A2(n8979), .B1(n7326), .B2(n8967), .ZN(n7200)
         );
  OAI211_X1 U8842 ( .C1(n8948), .C2(n7315), .A(n7200), .B(n7199), .ZN(n7201)
         );
  AOI21_X1 U8843 ( .B1(n7202), .B2(n8951), .A(n7201), .ZN(n7203) );
  OAI21_X1 U8844 ( .B1(n7204), .B2(n8969), .A(n7203), .ZN(P1_U3237) );
  INV_X1 U8845 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7214) );
  NOR2_X1 U8846 ( .A1(n7206), .A2(n7205), .ZN(n7207) );
  NAND2_X1 U8847 ( .A1(n9614), .A2(n7207), .ZN(n9138) );
  INV_X1 U8848 ( .A(n9138), .ZN(n9313) );
  OAI21_X1 U8849 ( .B1(n9313), .B2(n9500), .A(n7208), .ZN(n7213) );
  NOR2_X1 U8850 ( .A1(n9605), .A2(n7209), .ZN(n7210) );
  OAI21_X1 U8851 ( .B1(n7211), .B2(n7210), .A(n9614), .ZN(n7212) );
  OAI211_X1 U8852 ( .C1(n7214), .C2(n9614), .A(n7213), .B(n7212), .ZN(P1_U3291) );
  XNOR2_X1 U8853 ( .A(n7216), .B(n7215), .ZN(n7223) );
  INV_X1 U8854 ( .A(n7447), .ZN(n7217) );
  OAI22_X1 U8855 ( .A1(n8333), .A2(n7461), .B1(n8332), .B2(n7217), .ZN(n7220)
         );
  OAI21_X1 U8856 ( .B1(n8330), .B2(n7446), .A(n7218), .ZN(n7219) );
  NOR2_X1 U8857 ( .A1(n7220), .A2(n7219), .ZN(n7222) );
  NAND2_X1 U8858 ( .A1(n8336), .A2(n9843), .ZN(n7221) );
  OAI211_X1 U8859 ( .C1(n7223), .C2(n8340), .A(n7222), .B(n7221), .ZN(P2_U3238) );
  OR2_X1 U8860 ( .A1(n7346), .A2(n7224), .ZN(n8116) );
  NAND2_X1 U8861 ( .A1(n7346), .A2(n7224), .ZN(n8112) );
  INV_X1 U8862 ( .A(n7225), .ZN(n8367) );
  NAND2_X1 U8863 ( .A1(n7226), .A2(n8367), .ZN(n7227) );
  INV_X1 U8864 ( .A(n7349), .ZN(n7230) );
  AOI21_X1 U8865 ( .B1(n8052), .B2(n7231), .A(n7230), .ZN(n7240) );
  INV_X1 U8866 ( .A(n7446), .ZN(n8365) );
  AOI22_X1 U8867 ( .A1(n9770), .A2(n8367), .B1(n8365), .B2(n9771), .ZN(n7239)
         );
  INV_X1 U8868 ( .A(n8109), .ZN(n7232) );
  NOR3_X1 U8869 ( .A1(n7233), .A2(n8052), .A3(n7232), .ZN(n7237) );
  NAND2_X1 U8870 ( .A1(n7234), .A2(n8109), .ZN(n7235) );
  NAND2_X1 U8871 ( .A1(n7235), .A2(n8052), .ZN(n7345) );
  INV_X1 U8872 ( .A(n7345), .ZN(n7236) );
  OAI21_X1 U8873 ( .B1(n7237), .B2(n7236), .A(n9774), .ZN(n7238) );
  OAI211_X1 U8874 ( .C1(n7240), .C2(n9848), .A(n7239), .B(n7238), .ZN(n7249)
         );
  INV_X1 U8875 ( .A(n7249), .ZN(n7247) );
  INV_X1 U8876 ( .A(n7241), .ZN(n7242) );
  AOI211_X1 U8877 ( .C1(n7346), .C2(n7242), .A(n9838), .B(n7344), .ZN(n7248)
         );
  AOI22_X1 U8878 ( .A1(n4392), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7243), .B2(
        n9776), .ZN(n7244) );
  OAI21_X1 U8879 ( .B1(n7251), .B2(n9757), .A(n7244), .ZN(n7245) );
  AOI21_X1 U8880 ( .B1(n7248), .B2(n9734), .A(n7245), .ZN(n7246) );
  OAI21_X1 U8881 ( .B1(n7247), .B2(n4392), .A(n7246), .ZN(P2_U3287) );
  NOR2_X1 U8882 ( .A1(n7249), .A2(n7248), .ZN(n7256) );
  NAND2_X1 U8883 ( .A1(n9861), .A2(n9844), .ZN(n8754) );
  INV_X1 U8884 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7250) );
  OAI22_X1 U8885 ( .A1(n8754), .A2(n7251), .B1(n9861), .B2(n7250), .ZN(n7252)
         );
  INV_X1 U8886 ( .A(n7252), .ZN(n7253) );
  OAI21_X1 U8887 ( .B1(n7256), .B2(n9860), .A(n7253), .ZN(P2_U3478) );
  NAND2_X1 U8888 ( .A1(n9879), .A2(n9844), .ZN(n8713) );
  INV_X1 U8889 ( .A(n8713), .ZN(n7254) );
  AOI22_X1 U8890 ( .A1(n7254), .A2(n7346), .B1(n9877), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7255) );
  OAI21_X1 U8891 ( .B1(n7256), .B2(n9877), .A(n7255), .ZN(P2_U3529) );
  OR2_X1 U8892 ( .A1(n7257), .A2(n7267), .ZN(n7258) );
  NAND2_X1 U8893 ( .A1(n7259), .A2(n7258), .ZN(n9658) );
  OR2_X1 U8894 ( .A1(n7260), .A2(n9654), .ZN(n7261) );
  NAND2_X1 U8895 ( .A1(n7262), .A2(n7261), .ZN(n9655) );
  INV_X1 U8896 ( .A(n7263), .ZN(n7264) );
  INV_X1 U8897 ( .A(n9605), .ZN(n9499) );
  AOI22_X1 U8898 ( .A1(n9500), .A2(n7265), .B1(n7264), .B2(n9499), .ZN(n7266)
         );
  OAI21_X1 U8899 ( .B1(n9138), .B2(n9655), .A(n7266), .ZN(n7274) );
  XNOR2_X1 U8900 ( .A(n7268), .B(n7267), .ZN(n7272) );
  NAND2_X1 U8901 ( .A1(n9658), .A2(n9496), .ZN(n7271) );
  OAI22_X1 U8902 ( .A1(n7297), .A2(n9491), .B1(n9492), .B2(n7315), .ZN(n7269)
         );
  INV_X1 U8903 ( .A(n7269), .ZN(n7270) );
  OAI211_X1 U8904 ( .C1(n9488), .C2(n7272), .A(n7271), .B(n7270), .ZN(n9656)
         );
  MUX2_X1 U8905 ( .A(n9656), .B(P1_REG2_REG_4__SCAN_IN), .S(n4393), .Z(n7273)
         );
  AOI211_X1 U8906 ( .C1(n9508), .C2(n9658), .A(n7274), .B(n7273), .ZN(n7275)
         );
  INV_X1 U8907 ( .A(n7275), .ZN(P1_U3287) );
  XNOR2_X1 U8908 ( .A(n7418), .B(n4927), .ZN(n7276) );
  INV_X1 U8909 ( .A(n7527), .ZN(n8978) );
  INV_X1 U8910 ( .A(n7378), .ZN(n8980) );
  AOI222_X1 U8911 ( .A1(n9308), .A2(n7276), .B1(n8978), .B2(n9305), .C1(n8980), 
        .C2(n9303), .ZN(n7389) );
  OR2_X1 U8912 ( .A1(n7315), .A2(n9603), .ZN(n7277) );
  NAND2_X1 U8913 ( .A1(n7312), .A2(n7311), .ZN(n7310) );
  NAND2_X1 U8914 ( .A1(n7378), .A2(n9660), .ZN(n7279) );
  NAND2_X1 U8915 ( .A1(n7310), .A2(n7279), .ZN(n7281) );
  OAI21_X1 U8916 ( .B1(n7281), .B2(n7280), .A(n7417), .ZN(n7282) );
  INV_X1 U8917 ( .A(n7282), .ZN(n7390) );
  NOR2_X1 U8918 ( .A1(n7283), .A2(n7955), .ZN(n9601) );
  NAND2_X1 U8919 ( .A1(n9614), .A2(n9601), .ZN(n9351) );
  OAI22_X1 U8920 ( .A1(n9614), .A2(n7284), .B1(n7375), .B2(n9605), .ZN(n7285)
         );
  AOI21_X1 U8921 ( .B1(n9500), .B2(n7387), .A(n7285), .ZN(n7289) );
  OAI21_X1 U8922 ( .B1(n7322), .B2(n7415), .A(n9503), .ZN(n7286) );
  NOR2_X1 U8923 ( .A1(n7286), .A2(n7429), .ZN(n7386) );
  NOR2_X1 U8924 ( .A1(n7287), .A2(n9214), .ZN(n9507) );
  NAND2_X1 U8925 ( .A1(n7386), .A2(n9507), .ZN(n7288) );
  OAI211_X1 U8926 ( .C1(n7390), .C2(n9351), .A(n7289), .B(n7288), .ZN(n7290)
         );
  INV_X1 U8927 ( .A(n7290), .ZN(n7291) );
  OAI21_X1 U8928 ( .B1(n4393), .B2(n7389), .A(n7291), .ZN(P1_U3284) );
  XOR2_X1 U8929 ( .A(n7293), .B(n7292), .Z(n7300) );
  NAND2_X1 U8930 ( .A1(n7294), .A2(n7293), .ZN(n7295) );
  NAND2_X1 U8931 ( .A1(n7296), .A2(n7295), .ZN(n9653) );
  OAI22_X1 U8932 ( .A1(n6818), .A2(n9491), .B1(n9492), .B2(n7297), .ZN(n7298)
         );
  AOI21_X1 U8933 ( .B1(n9653), .B2(n9496), .A(n7298), .ZN(n7299) );
  OAI21_X1 U8934 ( .B1(n7300), .B2(n9488), .A(n7299), .ZN(n9651) );
  NAND2_X1 U8935 ( .A1(n7301), .A2(n7305), .ZN(n7302) );
  NAND2_X1 U8936 ( .A1(n7303), .A2(n7302), .ZN(n9650) );
  OAI22_X1 U8937 ( .A1(n9605), .A2(n10193), .B1(n6324), .B2(n9614), .ZN(n7304)
         );
  AOI21_X1 U8938 ( .B1(n9500), .B2(n7305), .A(n7304), .ZN(n7307) );
  NAND2_X1 U8939 ( .A1(n9653), .A2(n9508), .ZN(n7306) );
  OAI211_X1 U8940 ( .C1(n9138), .C2(n9650), .A(n7307), .B(n7306), .ZN(n7308)
         );
  AOI21_X1 U8941 ( .B1(n9614), .B2(n9651), .A(n7308), .ZN(n7309) );
  INV_X1 U8942 ( .A(n7309), .ZN(P1_U3289) );
  OAI21_X1 U8943 ( .B1(n7312), .B2(n7311), .A(n7310), .ZN(n9664) );
  INV_X1 U8944 ( .A(n9664), .ZN(n7329) );
  XNOR2_X1 U8945 ( .A(n7314), .B(n7313), .ZN(n7318) );
  OAI22_X1 U8946 ( .A1(n7315), .A2(n9491), .B1(n9492), .B2(n7423), .ZN(n7316)
         );
  AOI21_X1 U8947 ( .B1(n9664), .B2(n9496), .A(n7316), .ZN(n7317) );
  OAI21_X1 U8948 ( .B1(n9488), .B2(n7318), .A(n7317), .ZN(n9662) );
  NAND2_X1 U8949 ( .A1(n9662), .A2(n9614), .ZN(n7328) );
  OAI22_X1 U8950 ( .A1(n9614), .A2(n7320), .B1(n7319), .B2(n9605), .ZN(n7325)
         );
  INV_X1 U8951 ( .A(n7322), .ZN(n7323) );
  OAI21_X1 U8952 ( .B1(n9660), .B2(n4703), .A(n7323), .ZN(n9661) );
  NOR2_X1 U8953 ( .A1(n9661), .A2(n9138), .ZN(n7324) );
  AOI211_X1 U8954 ( .C1(n9500), .C2(n7326), .A(n7325), .B(n7324), .ZN(n7327)
         );
  OAI211_X1 U8955 ( .C1(n7329), .C2(n7653), .A(n7328), .B(n7327), .ZN(P1_U3285) );
  INV_X1 U8956 ( .A(n7330), .ZN(n7331) );
  NOR2_X1 U8957 ( .A1(n7332), .A2(n7331), .ZN(n7576) );
  XNOR2_X1 U8958 ( .A(n7580), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n7577) );
  XNOR2_X1 U8959 ( .A(n7576), .B(n7577), .ZN(n7343) );
  INV_X1 U8960 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7333) );
  NAND2_X1 U8961 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7814) );
  OAI21_X1 U8962 ( .B1(n8419), .B2(n7333), .A(n7814), .ZN(n7334) );
  AOI21_X1 U8963 ( .B1(n9709), .B2(n7335), .A(n7334), .ZN(n7341) );
  XNOR2_X1 U8964 ( .A(n7580), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n7338) );
  NAND2_X1 U8965 ( .A1(n7338), .A2(n7339), .ZN(n7571) );
  OAI211_X1 U8966 ( .C1(n7339), .C2(n7338), .A(n9715), .B(n7571), .ZN(n7340)
         );
  OAI211_X1 U8967 ( .C1(n7343), .C2(n7342), .A(n7341), .B(n7340), .ZN(P2_U3262) );
  OAI21_X1 U8968 ( .B1(n7344), .B2(n9837), .A(n7448), .ZN(n9839) );
  NAND2_X1 U8969 ( .A1(n7451), .A2(n7446), .ZN(n8118) );
  NAND2_X1 U8970 ( .A1(n8119), .A2(n8118), .ZN(n8048) );
  XNOR2_X1 U8971 ( .A(n7443), .B(n8048), .ZN(n7353) );
  AOI22_X1 U8972 ( .A1(n8366), .A2(n9770), .B1(n9771), .B2(n8364), .ZN(n7352)
         );
  OR2_X1 U8973 ( .A1(n7346), .A2(n8366), .ZN(n7347) );
  AND2_X1 U8974 ( .A1(n7349), .A2(n7347), .ZN(n7350) );
  AND2_X1 U8975 ( .A1(n8048), .A2(n7347), .ZN(n7348) );
  OAI211_X1 U8976 ( .C1(n7350), .C2(n8048), .A(n9859), .B(n7453), .ZN(n7351)
         );
  OAI211_X1 U8977 ( .C1(n7353), .C2(n9740), .A(n7352), .B(n7351), .ZN(n9841)
         );
  NAND2_X1 U8978 ( .A1(n9841), .A2(n9785), .ZN(n7358) );
  INV_X1 U8979 ( .A(n7354), .ZN(n7355) );
  OAI22_X1 U8980 ( .A1(n9785), .A2(n6456), .B1(n7355), .B2(n9750), .ZN(n7356)
         );
  AOI21_X1 U8981 ( .B1(n9726), .B2(n7451), .A(n7356), .ZN(n7357) );
  OAI211_X1 U8982 ( .C1(n8562), .C2(n9839), .A(n7358), .B(n7357), .ZN(P2_U3286) );
  INV_X1 U8983 ( .A(n7359), .ZN(n7361) );
  OAI222_X1 U8984 ( .A1(n8771), .A2(n7360), .B1(n8769), .B2(n7361), .C1(n8226), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  OAI222_X1 U8985 ( .A1(n9479), .A2(n7363), .B1(P1_U3084), .B2(n7362), .C1(
        n9473), .C2(n7361), .ZN(P1_U3333) );
  OAI22_X1 U8986 ( .A1(n7423), .A2(n7848), .B1(n7415), .B2(n6832), .ZN(n7364)
         );
  XNOR2_X1 U8987 ( .A(n7364), .B(n7955), .ZN(n7366) );
  AOI22_X1 U8988 ( .A1(n7994), .A2(n8979), .B1(n7990), .B2(n7387), .ZN(n7365)
         );
  OR2_X1 U8989 ( .A1(n7366), .A2(n7365), .ZN(n7526) );
  NAND2_X1 U8990 ( .A1(n7366), .A2(n7365), .ZN(n7524) );
  NAND2_X1 U8991 ( .A1(n7526), .A2(n7524), .ZN(n7374) );
  INV_X1 U8992 ( .A(n7367), .ZN(n7370) );
  INV_X1 U8993 ( .A(n7368), .ZN(n7369) );
  NAND2_X1 U8994 ( .A1(n7370), .A2(n7369), .ZN(n7371) );
  XOR2_X1 U8995 ( .A(n7374), .B(n7525), .Z(n7382) );
  INV_X1 U8996 ( .A(n7375), .ZN(n7380) );
  AOI22_X1 U8997 ( .A1(n8921), .A2(n8978), .B1(n7387), .B2(n8967), .ZN(n7377)
         );
  OAI211_X1 U8998 ( .C1(n8948), .C2(n7378), .A(n7377), .B(n7376), .ZN(n7379)
         );
  AOI21_X1 U8999 ( .B1(n7380), .B2(n8951), .A(n7379), .ZN(n7381) );
  OAI21_X1 U9000 ( .B1(n7382), .B2(n8969), .A(n7381), .ZN(P1_U3211) );
  INV_X1 U9001 ( .A(n7383), .ZN(n8269) );
  OAI222_X1 U9002 ( .A1(n8771), .A2(n7385), .B1(n8769), .B2(n8269), .C1(n7384), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  INV_X1 U9003 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10119) );
  AOI21_X1 U9004 ( .B1(n9432), .B2(n7387), .A(n7386), .ZN(n7388) );
  OAI211_X1 U9005 ( .C1(n7390), .C2(n9434), .A(n7389), .B(n7388), .ZN(n7392)
         );
  NAND2_X1 U9006 ( .A1(n7392), .A2(n9675), .ZN(n7391) );
  OAI21_X1 U9007 ( .B1(n9675), .B2(n10119), .A(n7391), .ZN(P1_U3475) );
  NAND2_X1 U9008 ( .A1(n7392), .A2(n9683), .ZN(n7393) );
  OAI21_X1 U9009 ( .B1(n9683), .B2(n5489), .A(n7393), .ZN(P1_U3530) );
  INV_X1 U9010 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7404) );
  OAI21_X1 U9011 ( .B1(n7396), .B2(n7395), .A(n7394), .ZN(n7402) );
  NAND2_X1 U9012 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n8787) );
  OAI21_X1 U9013 ( .B1(n9583), .B2(n7397), .A(n8787), .ZN(n7401) );
  AOI211_X1 U9014 ( .C1(n7399), .C2(n7707), .A(n7398), .B(n9591), .ZN(n7400)
         );
  AOI211_X1 U9015 ( .C1(n9597), .C2(n7402), .A(n7401), .B(n7400), .ZN(n7403)
         );
  OAI21_X1 U9016 ( .B1(n9586), .B2(n7404), .A(n7403), .ZN(P1_U3255) );
  INV_X1 U9017 ( .A(n7405), .ZN(n7406) );
  AOI21_X1 U9018 ( .B1(n7408), .B2(n7407), .A(n7406), .ZN(n7414) );
  AND2_X1 U9019 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8393) );
  OR2_X1 U9020 ( .A1(n7596), .A2(n9743), .ZN(n7410) );
  NAND2_X1 U9021 ( .A1(n8364), .A2(n9770), .ZN(n7409) );
  AND2_X1 U9022 ( .A1(n7410), .A2(n7409), .ZN(n7462) );
  NOR2_X1 U9023 ( .A1(n7627), .A2(n7462), .ZN(n7411) );
  AOI211_X1 U9024 ( .C1(n7469), .C2(n8344), .A(n8393), .B(n7411), .ZN(n7413)
         );
  NAND2_X1 U9025 ( .A1(n8336), .A2(n7559), .ZN(n7412) );
  OAI211_X1 U9026 ( .C1(n7414), .C2(n8340), .A(n7413), .B(n7412), .ZN(P2_U3226) );
  NAND2_X1 U9027 ( .A1(n7423), .A2(n7415), .ZN(n7416) );
  OAI21_X1 U9028 ( .B1(n4489), .B2(n7421), .A(n7511), .ZN(n9665) );
  OR2_X1 U9029 ( .A1(n9665), .A2(n7645), .ZN(n7427) );
  NAND2_X1 U9030 ( .A1(n7418), .A2(n4927), .ZN(n7420) );
  AOI21_X1 U9031 ( .B1(n7422), .B2(n7421), .A(n9488), .ZN(n7425) );
  OAI22_X1 U9032 ( .A1(n7423), .A2(n9491), .B1(n9492), .B2(n9490), .ZN(n7424)
         );
  AOI21_X1 U9033 ( .B1(n7425), .B2(n7513), .A(n7424), .ZN(n7426) );
  NAND2_X1 U9034 ( .A1(n7427), .A2(n7426), .ZN(n9670) );
  NAND2_X1 U9035 ( .A1(n9670), .A2(n9614), .ZN(n7433) );
  OAI22_X1 U9036 ( .A1(n9614), .A2(n7428), .B1(n7534), .B2(n9605), .ZN(n7431)
         );
  INV_X1 U9037 ( .A(n7537), .ZN(n9667) );
  OAI21_X1 U9038 ( .B1(n7429), .B2(n9667), .A(n7516), .ZN(n9669) );
  NOR2_X1 U9039 ( .A1(n9669), .A2(n9138), .ZN(n7430) );
  AOI211_X1 U9040 ( .C1(n9500), .C2(n7537), .A(n7431), .B(n7430), .ZN(n7432)
         );
  OAI211_X1 U9041 ( .C1(n9665), .C2(n7653), .A(n7433), .B(n7432), .ZN(P1_U3283) );
  XNOR2_X1 U9042 ( .A(n7435), .B(n7434), .ZN(n7442) );
  OR2_X1 U9043 ( .A1(n7670), .A2(n9743), .ZN(n7437) );
  OR2_X1 U9044 ( .A1(n7461), .A2(n9745), .ZN(n7436) );
  AND2_X1 U9045 ( .A1(n7437), .A2(n7436), .ZN(n7563) );
  OAI22_X1 U9046 ( .A1(n7627), .A2(n7563), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7438), .ZN(n7440) );
  INV_X1 U9047 ( .A(n7602), .ZN(n7737) );
  NOR2_X1 U9048 ( .A1(n7737), .A2(n8349), .ZN(n7439) );
  AOI211_X1 U9049 ( .C1(n7566), .C2(n8344), .A(n7440), .B(n7439), .ZN(n7441)
         );
  OAI21_X1 U9050 ( .B1(n7442), .B2(n8340), .A(n7441), .ZN(P2_U3236) );
  AND2_X1 U9051 ( .A1(n7450), .A2(n8364), .ZN(n8122) );
  NAND2_X1 U9052 ( .A1(n9843), .A2(n7444), .ZN(n8128) );
  NAND2_X1 U9053 ( .A1(n4395), .A2(n8128), .ZN(n7454) );
  INV_X1 U9054 ( .A(n7454), .ZN(n8051) );
  XNOR2_X1 U9055 ( .A(n7460), .B(n8051), .ZN(n7445) );
  OAI222_X1 U9056 ( .A1(n9743), .A2(n7461), .B1(n9745), .B2(n7446), .C1(n9740), 
        .C2(n7445), .ZN(n9851) );
  AOI21_X1 U9057 ( .B1(n7447), .B2(n9776), .A(n9851), .ZN(n7459) );
  NAND2_X1 U9058 ( .A1(n7448), .A2(n9843), .ZN(n7449) );
  AND2_X1 U9059 ( .A1(n7467), .A2(n7449), .ZN(n9846) );
  OAI22_X1 U9060 ( .A1(n9757), .A2(n7450), .B1(n9785), .B2(n6457), .ZN(n7457)
         );
  NAND2_X1 U9061 ( .A1(n7451), .A2(n8365), .ZN(n7452) );
  OAI21_X1 U9062 ( .B1(n7455), .B2(n7454), .A(n7465), .ZN(n9849) );
  NOR2_X1 U9063 ( .A1(n9849), .A2(n9755), .ZN(n7456) );
  AOI211_X1 U9064 ( .C1(n9761), .C2(n9846), .A(n7457), .B(n7456), .ZN(n7458)
         );
  OAI21_X1 U9065 ( .B1(n7459), .B2(n4392), .A(n7458), .ZN(P2_U3285) );
  INV_X1 U9066 ( .A(n7559), .ZN(n9855) );
  INV_X1 U9067 ( .A(n7461), .ZN(n8363) );
  INV_X1 U9068 ( .A(n8127), .ZN(n8130) );
  NAND2_X1 U9069 ( .A1(n7559), .A2(n7461), .ZN(n8129) );
  XNOR2_X1 U9070 ( .A(n7554), .B(n8053), .ZN(n7463) );
  OAI21_X1 U9071 ( .B1(n7463), .B2(n9740), .A(n7462), .ZN(n9856) );
  INV_X1 U9072 ( .A(n9856), .ZN(n7474) );
  NAND2_X1 U9073 ( .A1(n9843), .A2(n8364), .ZN(n7464) );
  INV_X1 U9074 ( .A(n8053), .ZN(n7466) );
  OAI21_X1 U9075 ( .B1(n4495), .B2(n7466), .A(n7561), .ZN(n9858) );
  INV_X1 U9076 ( .A(n7467), .ZN(n7468) );
  OAI211_X1 U9077 ( .C1(n7468), .C2(n9855), .A(n9845), .B(n7565), .ZN(n9853)
         );
  INV_X1 U9078 ( .A(n9734), .ZN(n8578) );
  AOI22_X1 U9079 ( .A1(n4392), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7469), .B2(
        n9776), .ZN(n7471) );
  NAND2_X1 U9080 ( .A1(n9726), .A2(n7559), .ZN(n7470) );
  OAI211_X1 U9081 ( .C1(n9853), .C2(n8578), .A(n7471), .B(n7470), .ZN(n7472)
         );
  AOI21_X1 U9082 ( .B1(n9858), .B2(n9782), .A(n7472), .ZN(n7473) );
  OAI21_X1 U9083 ( .B1(n7474), .B2(n4392), .A(n7473), .ZN(P2_U3284) );
  INV_X1 U9084 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U9085 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7475) );
  AOI21_X1 U9086 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7475), .ZN(n9886) );
  NOR2_X1 U9087 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7476) );
  AOI21_X1 U9088 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7476), .ZN(n9889) );
  NOR2_X1 U9089 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7477) );
  AOI21_X1 U9090 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7477), .ZN(n9892) );
  NOR2_X1 U9091 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7478) );
  AOI21_X1 U9092 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7478), .ZN(n9895) );
  NOR2_X1 U9093 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7479) );
  AOI21_X1 U9094 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7479), .ZN(n9898) );
  NOR2_X1 U9095 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7486) );
  XNOR2_X1 U9096 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10235) );
  NAND2_X1 U9097 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7484) );
  XOR2_X1 U9098 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10233) );
  NAND2_X1 U9099 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7482) );
  XOR2_X1 U9100 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10231) );
  AOI21_X1 U9101 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9880) );
  INV_X1 U9102 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7480) );
  NAND3_X1 U9103 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9882) );
  OAI21_X1 U9104 ( .B1(n9880), .B2(n7480), .A(n9882), .ZN(n10230) );
  NAND2_X1 U9105 ( .A1(n10231), .A2(n10230), .ZN(n7481) );
  NAND2_X1 U9106 ( .A1(n7482), .A2(n7481), .ZN(n10232) );
  NAND2_X1 U9107 ( .A1(n10233), .A2(n10232), .ZN(n7483) );
  NAND2_X1 U9108 ( .A1(n7484), .A2(n7483), .ZN(n10234) );
  NOR2_X1 U9109 ( .A1(n10235), .A2(n10234), .ZN(n7485) );
  NOR2_X1 U9110 ( .A1(n7486), .A2(n7485), .ZN(n7487) );
  NOR2_X1 U9111 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7487), .ZN(n10218) );
  AND2_X1 U9112 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7487), .ZN(n10219) );
  NOR2_X1 U9113 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10219), .ZN(n7488) );
  NOR2_X1 U9114 ( .A1(n10218), .A2(n7488), .ZN(n7489) );
  NAND2_X1 U9115 ( .A1(n7489), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7491) );
  XOR2_X1 U9116 ( .A(n7489), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10217) );
  NAND2_X1 U9117 ( .A1(n10217), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7490) );
  NAND2_X1 U9118 ( .A1(n7491), .A2(n7490), .ZN(n7492) );
  NAND2_X1 U9119 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7492), .ZN(n7494) );
  XOR2_X1 U9120 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7492), .Z(n10229) );
  NAND2_X1 U9121 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10229), .ZN(n7493) );
  NAND2_X1 U9122 ( .A1(n7494), .A2(n7493), .ZN(n7495) );
  NAND2_X1 U9123 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7495), .ZN(n7497) );
  XOR2_X1 U9124 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7495), .Z(n10228) );
  NAND2_X1 U9125 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10228), .ZN(n7496) );
  NAND2_X1 U9126 ( .A1(n7497), .A2(n7496), .ZN(n7498) );
  AND2_X1 U9127 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7498), .ZN(n7499) );
  XNOR2_X1 U9128 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7498), .ZN(n10226) );
  NOR2_X1 U9129 ( .A1(n10227), .A2(n10226), .ZN(n10225) );
  NOR2_X1 U9130 ( .A1(n7499), .A2(n10225), .ZN(n9907) );
  NAND2_X1 U9131 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7500) );
  OAI21_X1 U9132 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7500), .ZN(n9906) );
  NOR2_X1 U9133 ( .A1(n9907), .A2(n9906), .ZN(n9905) );
  AOI21_X1 U9134 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9905), .ZN(n9904) );
  NAND2_X1 U9135 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7501) );
  OAI21_X1 U9136 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7501), .ZN(n9903) );
  NOR2_X1 U9137 ( .A1(n9904), .A2(n9903), .ZN(n9902) );
  AOI21_X1 U9138 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9902), .ZN(n9901) );
  NOR2_X1 U9139 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7502) );
  AOI21_X1 U9140 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7502), .ZN(n9900) );
  NAND2_X1 U9141 ( .A1(n9901), .A2(n9900), .ZN(n9899) );
  OAI21_X1 U9142 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9899), .ZN(n9897) );
  NAND2_X1 U9143 ( .A1(n9898), .A2(n9897), .ZN(n9896) );
  OAI21_X1 U9144 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9896), .ZN(n9894) );
  NAND2_X1 U9145 ( .A1(n9895), .A2(n9894), .ZN(n9893) );
  OAI21_X1 U9146 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9893), .ZN(n9891) );
  NAND2_X1 U9147 ( .A1(n9892), .A2(n9891), .ZN(n9890) );
  OAI21_X1 U9148 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9890), .ZN(n9888) );
  NAND2_X1 U9149 ( .A1(n9889), .A2(n9888), .ZN(n9887) );
  OAI21_X1 U9150 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9887), .ZN(n9885) );
  NAND2_X1 U9151 ( .A1(n9886), .A2(n9885), .ZN(n9884) );
  OAI21_X1 U9152 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9884), .ZN(n10222) );
  NOR2_X1 U9153 ( .A1(n10223), .A2(n10222), .ZN(n7503) );
  NAND2_X1 U9154 ( .A1(n10223), .A2(n10222), .ZN(n10221) );
  OAI21_X1 U9155 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7503), .A(n10221), .ZN(
        n7507) );
  NOR2_X1 U9156 ( .A1(n7504), .A2(n7505), .ZN(n7506) );
  XNOR2_X1 U9157 ( .A(n7507), .B(n7506), .ZN(ADD_1071_U4) );
  INV_X1 U9158 ( .A(n7508), .ZN(n8007) );
  OAI222_X1 U9159 ( .A1(n8771), .A2(n7510), .B1(n8769), .B2(n8007), .C1(
        P2_U3152), .C2(n7509), .ZN(P2_U3336) );
  XNOR2_X1 U9160 ( .A(n7634), .B(n7514), .ZN(n7553) );
  XNOR2_X1 U9161 ( .A(n9485), .B(n7514), .ZN(n7515) );
  AOI222_X1 U9162 ( .A1(n9308), .A2(n7515), .B1(n8976), .B2(n9305), .C1(n8978), 
        .C2(n9303), .ZN(n7548) );
  INV_X1 U9163 ( .A(n7647), .ZN(n9505) );
  AOI21_X1 U9164 ( .B1(n8885), .B2(n7516), .A(n9505), .ZN(n7551) );
  AOI22_X1 U9165 ( .A1(n7551), .A2(n9503), .B1(n9432), .B2(n8885), .ZN(n7517)
         );
  OAI211_X1 U9166 ( .C1(n9434), .C2(n7553), .A(n7548), .B(n7517), .ZN(n7519)
         );
  NAND2_X1 U9167 ( .A1(n7519), .A2(n9675), .ZN(n7518) );
  OAI21_X1 U9168 ( .B1(n9675), .B2(n5342), .A(n7518), .ZN(P1_U3481) );
  NAND2_X1 U9169 ( .A1(n7519), .A2(n9683), .ZN(n7520) );
  OAI21_X1 U9170 ( .B1(n9683), .B2(n6345), .A(n7520), .ZN(P1_U3532) );
  NAND2_X1 U9171 ( .A1(n7537), .A2(n7991), .ZN(n7522) );
  OAI21_X1 U9172 ( .B1(n7527), .B2(n7848), .A(n7522), .ZN(n7523) );
  XNOR2_X1 U9173 ( .A(n7523), .B(n7992), .ZN(n7846) );
  OR2_X1 U9174 ( .A1(n7963), .A2(n7527), .ZN(n7529) );
  NAND2_X1 U9175 ( .A1(n7995), .A2(n7537), .ZN(n7528) );
  NAND2_X1 U9176 ( .A1(n7847), .A2(n7845), .ZN(n7530) );
  XOR2_X1 U9177 ( .A(n7846), .B(n7530), .Z(n7539) );
  NAND2_X1 U9178 ( .A1(n8921), .A2(n8977), .ZN(n7533) );
  NAND2_X1 U9179 ( .A1(n8962), .A2(n8979), .ZN(n7532) );
  NAND3_X1 U9180 ( .A1(n7533), .A2(n7532), .A3(n7531), .ZN(n7536) );
  NOR2_X1 U9181 ( .A1(n8965), .A2(n7534), .ZN(n7535) );
  AOI211_X1 U9182 ( .C1(n7537), .C2(n8967), .A(n7536), .B(n7535), .ZN(n7538)
         );
  OAI21_X1 U9183 ( .B1(n7539), .B2(n8969), .A(n7538), .ZN(P1_U3219) );
  INV_X1 U9184 ( .A(n7542), .ZN(n7541) );
  NAND2_X1 U9185 ( .A1(n8758), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7540) );
  OAI211_X1 U9186 ( .C1(n7541), .C2(n8769), .A(n8237), .B(n7540), .ZN(P2_U3335) );
  NAND2_X1 U9187 ( .A1(n7542), .A2(n9474), .ZN(n7544) );
  OAI211_X1 U9188 ( .C1(n7545), .C2(n9468), .A(n7544), .B(n7543), .ZN(P1_U3330) );
  INV_X1 U9189 ( .A(n8883), .ZN(n7546) );
  AOI22_X1 U9190 ( .A1(n4393), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7546), .B2(
        n9499), .ZN(n7547) );
  OAI21_X1 U9191 ( .B1(n4706), .B2(n9338), .A(n7547), .ZN(n7550) );
  NOR2_X1 U9192 ( .A1(n7548), .A2(n4393), .ZN(n7549) );
  AOI211_X1 U9193 ( .C1(n7551), .C2(n9313), .A(n7550), .B(n7549), .ZN(n7552)
         );
  OAI21_X1 U9194 ( .B1(n9351), .B2(n7553), .A(n7552), .ZN(P1_U3282) );
  OR2_X1 U9195 ( .A1(n7602), .A2(n7596), .ZN(n8132) );
  NAND2_X1 U9196 ( .A1(n7602), .A2(n7596), .ZN(n8131) );
  NAND2_X1 U9197 ( .A1(n8132), .A2(n8131), .ZN(n8135) );
  NAND2_X1 U9198 ( .A1(n7554), .A2(n8129), .ZN(n7556) );
  NAND2_X1 U9199 ( .A1(n7556), .A2(n8130), .ZN(n7558) );
  NOR2_X1 U9200 ( .A1(n8135), .A2(n8127), .ZN(n7555) );
  NAND2_X1 U9201 ( .A1(n7556), .A2(n7555), .ZN(n7607) );
  INV_X1 U9202 ( .A(n7607), .ZN(n7557) );
  AOI21_X1 U9203 ( .B1(n8135), .B2(n7558), .A(n7557), .ZN(n7564) );
  OR2_X1 U9204 ( .A1(n7559), .A2(n8363), .ZN(n7560) );
  OAI211_X1 U9205 ( .C1(n4490), .C2(n8135), .A(n7605), .B(n9859), .ZN(n7562)
         );
  OAI211_X1 U9206 ( .C1(n7564), .C2(n9740), .A(n7563), .B(n7562), .ZN(n7731)
         );
  INV_X1 U9207 ( .A(n7731), .ZN(n7570) );
  AOI21_X1 U9208 ( .B1(n7602), .B2(n7565), .A(n7612), .ZN(n7732) );
  AOI22_X1 U9209 ( .A1(n4392), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7566), .B2(
        n9776), .ZN(n7567) );
  OAI21_X1 U9210 ( .B1(n7737), .B2(n9757), .A(n7567), .ZN(n7568) );
  AOI21_X1 U9211 ( .B1(n7732), .B2(n9761), .A(n7568), .ZN(n7569) );
  OAI21_X1 U9212 ( .B1(n7570), .B2(n4392), .A(n7569), .ZN(P2_U3283) );
  INV_X1 U9213 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7572) );
  OAI21_X1 U9214 ( .B1(n7580), .B2(n7572), .A(n7571), .ZN(n7573) );
  NOR2_X1 U9215 ( .A1(n7573), .A2(n7588), .ZN(n8404) );
  NOR2_X1 U9216 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n7574), .ZN(n8405) );
  AOI21_X1 U9217 ( .B1(n7574), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8405), .ZN(
        n7590) );
  OR2_X1 U9218 ( .A1(n7588), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U9219 ( .A1(n7588), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7575) );
  AND2_X1 U9220 ( .A1(n8407), .A2(n7575), .ZN(n7583) );
  INV_X1 U9221 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7579) );
  NAND2_X1 U9222 ( .A1(n7577), .A2(n7576), .ZN(n7578) );
  OAI21_X1 U9223 ( .B1(n7580), .B2(n7579), .A(n7578), .ZN(n7581) );
  INV_X1 U9224 ( .A(n7581), .ZN(n7582) );
  NAND2_X1 U9225 ( .A1(n7583), .A2(n7582), .ZN(n8408) );
  OAI21_X1 U9226 ( .B1(n7583), .B2(n7582), .A(n8408), .ZN(n7584) );
  NAND2_X1 U9227 ( .A1(n9711), .A2(n7584), .ZN(n7586) );
  NAND2_X1 U9228 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3152), .ZN(n7585) );
  OAI211_X1 U9229 ( .C1(n8419), .C2(n10223), .A(n7586), .B(n7585), .ZN(n7587)
         );
  AOI21_X1 U9230 ( .B1(n7588), .B2(n9709), .A(n7587), .ZN(n7589) );
  OAI21_X1 U9231 ( .B1(n7590), .B2(n9686), .A(n7589), .ZN(P2_U3263) );
  INV_X1 U9232 ( .A(n7671), .ZN(n9518) );
  OAI21_X1 U9233 ( .B1(n7593), .B2(n7592), .A(n7591), .ZN(n7595) );
  NAND2_X1 U9234 ( .A1(n7595), .A2(n7594), .ZN(n7601) );
  INV_X1 U9235 ( .A(n7596), .ZN(n8362) );
  INV_X1 U9236 ( .A(n8360), .ZN(n7777) );
  INV_X1 U9237 ( .A(n7597), .ZN(n7614) );
  OAI22_X1 U9238 ( .A1(n8333), .A2(n7777), .B1(n8332), .B2(n7614), .ZN(n7598)
         );
  AOI211_X1 U9239 ( .C1(n8343), .C2(n8362), .A(n7599), .B(n7598), .ZN(n7600)
         );
  OAI211_X1 U9240 ( .C1(n9518), .C2(n8349), .A(n7601), .B(n7600), .ZN(P2_U3217) );
  NAND2_X1 U9241 ( .A1(n7602), .A2(n8362), .ZN(n7603) );
  AND2_X1 U9242 ( .A1(n7605), .A2(n7603), .ZN(n7606) );
  NAND2_X1 U9243 ( .A1(n7671), .A2(n7670), .ZN(n8137) );
  NAND2_X1 U9244 ( .A1(n8136), .A2(n8137), .ZN(n8055) );
  AND2_X1 U9245 ( .A1(n8055), .A2(n7603), .ZN(n7604) );
  OAI21_X1 U9246 ( .B1(n7606), .B2(n8055), .A(n7673), .ZN(n9522) );
  INV_X1 U9247 ( .A(n9522), .ZN(n7619) );
  INV_X1 U9248 ( .A(n8055), .ZN(n8134) );
  OAI211_X1 U9249 ( .C1(n7609), .C2(n8134), .A(n9774), .B(n7674), .ZN(n7611)
         );
  AOI22_X1 U9250 ( .A1(n8362), .A2(n9770), .B1(n9771), .B2(n8360), .ZN(n7610)
         );
  NAND2_X1 U9251 ( .A1(n7611), .A2(n7610), .ZN(n9520) );
  NOR2_X1 U9252 ( .A1(n7612), .A2(n9518), .ZN(n7613) );
  OR2_X1 U9253 ( .A1(n7678), .A2(n7613), .ZN(n9519) );
  OAI22_X1 U9254 ( .A1(n9785), .A2(n6949), .B1(n7614), .B2(n9750), .ZN(n7615)
         );
  AOI21_X1 U9255 ( .B1(n7671), .B2(n9726), .A(n7615), .ZN(n7616) );
  OAI21_X1 U9256 ( .B1(n9519), .B2(n8562), .A(n7616), .ZN(n7617) );
  AOI21_X1 U9257 ( .B1(n9520), .B2(n9785), .A(n7617), .ZN(n7618) );
  OAI21_X1 U9258 ( .B1(n7619), .B2(n9755), .A(n7618), .ZN(P2_U3282) );
  XNOR2_X1 U9259 ( .A(n7621), .B(n7620), .ZN(n7622) );
  XNOR2_X1 U9260 ( .A(n7623), .B(n7622), .ZN(n7631) );
  OR2_X1 U9261 ( .A1(n8359), .A2(n9743), .ZN(n7625) );
  OR2_X1 U9262 ( .A1(n7670), .A2(n9745), .ZN(n7624) );
  AND2_X1 U9263 ( .A1(n7625), .A2(n7624), .ZN(n7676) );
  OAI22_X1 U9264 ( .A1(n7627), .A2(n7676), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7626), .ZN(n7629) );
  INV_X1 U9265 ( .A(n8141), .ZN(n8142) );
  NOR2_X1 U9266 ( .A1(n8142), .A2(n8349), .ZN(n7628) );
  AOI211_X1 U9267 ( .C1(n7680), .C2(n8344), .A(n7629), .B(n7628), .ZN(n7630)
         );
  OAI21_X1 U9268 ( .B1(n7631), .B2(n8340), .A(n7630), .ZN(P2_U3243) );
  AND2_X1 U9269 ( .A1(n8885), .A2(n8977), .ZN(n7633) );
  OR2_X1 U9270 ( .A1(n8885), .A2(n8977), .ZN(n7632) );
  NOR2_X1 U9271 ( .A1(n9501), .A2(n8976), .ZN(n7635) );
  XNOR2_X1 U9272 ( .A(n7749), .B(n7636), .ZN(n9541) );
  XNOR2_X1 U9273 ( .A(n7692), .B(n7640), .ZN(n7643) );
  OAI22_X1 U9274 ( .A1(n7641), .A2(n9491), .B1(n9492), .B2(n8906), .ZN(n7642)
         );
  AOI21_X1 U9275 ( .B1(n7643), .B2(n9308), .A(n7642), .ZN(n7644) );
  OAI21_X1 U9276 ( .B1(n9541), .B2(n7645), .A(n7644), .ZN(n9544) );
  NAND2_X1 U9277 ( .A1(n9544), .A2(n9614), .ZN(n7652) );
  OAI22_X1 U9278 ( .A1(n9614), .A2(n7646), .B1(n8924), .B2(n9605), .ZN(n7650)
         );
  INV_X1 U9279 ( .A(n8930), .ZN(n9542) );
  NOR2_X1 U9280 ( .A1(n9502), .A2(n9542), .ZN(n7648) );
  OR2_X1 U9281 ( .A1(n7664), .A2(n7648), .ZN(n9543) );
  NOR2_X1 U9282 ( .A1(n9543), .A2(n9138), .ZN(n7649) );
  AOI211_X1 U9283 ( .C1(n9500), .C2(n8930), .A(n7650), .B(n7649), .ZN(n7651)
         );
  OAI211_X1 U9284 ( .C1(n9541), .C2(n7653), .A(n7652), .B(n7651), .ZN(P1_U3280) );
  OR2_X1 U9285 ( .A1(n8930), .A2(n8975), .ZN(n7698) );
  NAND2_X1 U9286 ( .A1(n7749), .A2(n7698), .ZN(n7654) );
  NAND2_X1 U9287 ( .A1(n8930), .A2(n8975), .ZN(n7702) );
  NAND2_X1 U9288 ( .A1(n7654), .A2(n7702), .ZN(n7655) );
  XNOR2_X1 U9289 ( .A(n7655), .B(n4457), .ZN(n9538) );
  INV_X1 U9290 ( .A(n7656), .ZN(n7658) );
  OAI21_X1 U9291 ( .B1(n7692), .B2(n7658), .A(n7657), .ZN(n7659) );
  XNOR2_X1 U9292 ( .A(n7659), .B(n4457), .ZN(n7662) );
  OAI22_X1 U9293 ( .A1(n9493), .A2(n9491), .B1(n9492), .B2(n8788), .ZN(n7660)
         );
  INV_X1 U9294 ( .A(n7660), .ZN(n7661) );
  OAI21_X1 U9295 ( .B1(n7662), .B2(n9488), .A(n7661), .ZN(n7663) );
  AOI21_X1 U9296 ( .B1(n9538), .B2(n9496), .A(n7663), .ZN(n9540) );
  INV_X1 U9297 ( .A(n8837), .ZN(n9536) );
  OAI211_X1 U9298 ( .C1(n7664), .C2(n9536), .A(n9503), .B(n7724), .ZN(n9535)
         );
  INV_X1 U9299 ( .A(n9507), .ZN(n7767) );
  INV_X1 U9300 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7665) );
  OAI22_X1 U9301 ( .A1(n9614), .A2(n7665), .B1(n8835), .B2(n9605), .ZN(n7666)
         );
  AOI21_X1 U9302 ( .B1(n8837), .B2(n9500), .A(n7666), .ZN(n7667) );
  OAI21_X1 U9303 ( .B1(n9535), .B2(n7767), .A(n7667), .ZN(n7668) );
  AOI21_X1 U9304 ( .B1(n9538), .B2(n9508), .A(n7668), .ZN(n7669) );
  OAI21_X1 U9305 ( .B1(n9540), .B2(n4393), .A(n7669), .ZN(P1_U3279) );
  INV_X1 U9306 ( .A(n7670), .ZN(n8361) );
  OR2_X1 U9307 ( .A1(n7671), .A2(n8361), .ZN(n7672) );
  NAND2_X1 U9308 ( .A1(n7673), .A2(n7672), .ZN(n7772) );
  XNOR2_X1 U9309 ( .A(n8141), .B(n8360), .ZN(n8139) );
  INV_X1 U9310 ( .A(n8139), .ZN(n7771) );
  XNOR2_X1 U9311 ( .A(n7772), .B(n7771), .ZN(n7804) );
  INV_X1 U9312 ( .A(n7804), .ZN(n7685) );
  NAND3_X1 U9313 ( .A1(n7674), .A2(n7771), .A3(n8136), .ZN(n7675) );
  NAND3_X1 U9314 ( .A1(n7776), .A2(n9774), .A3(n7675), .ZN(n7677) );
  NAND2_X1 U9315 ( .A1(n7677), .A2(n7676), .ZN(n7803) );
  OAI21_X1 U9316 ( .B1(n7678), .B2(n8142), .A(n9845), .ZN(n7679) );
  OR2_X1 U9317 ( .A1(n7781), .A2(n7679), .ZN(n7801) );
  AOI22_X1 U9318 ( .A1(n4392), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7680), .B2(
        n9776), .ZN(n7682) );
  NAND2_X1 U9319 ( .A1(n8141), .A2(n9726), .ZN(n7681) );
  OAI211_X1 U9320 ( .C1(n7801), .C2(n8578), .A(n7682), .B(n7681), .ZN(n7683)
         );
  AOI21_X1 U9321 ( .B1(n7803), .B2(n9785), .A(n7683), .ZN(n7684) );
  OAI21_X1 U9322 ( .B1(n7685), .B2(n9755), .A(n7684), .ZN(P2_U3281) );
  INV_X1 U9323 ( .A(n7686), .ZN(n7688) );
  OAI222_X1 U9324 ( .A1(P2_U3152), .A2(n7687), .B1(n8769), .B2(n7688), .C1(
        n9911), .C2(n8771), .ZN(P2_U3334) );
  OAI222_X1 U9325 ( .A1(n9479), .A2(n7690), .B1(P1_U3084), .B2(n7689), .C1(
        n9473), .C2(n7688), .ZN(P1_U3329) );
  INV_X1 U9326 ( .A(n7753), .ZN(n7695) );
  XNOR2_X1 U9327 ( .A(n7754), .B(n7695), .ZN(n7697) );
  OAI22_X1 U9328 ( .A1(n9348), .A2(n9492), .B1(n9491), .B2(n8788), .ZN(n7696)
         );
  AOI21_X1 U9329 ( .B1(n7697), .B2(n9308), .A(n7696), .ZN(n9526) );
  NAND2_X1 U9330 ( .A1(n8837), .A2(n8974), .ZN(n7701) );
  AND2_X1 U9331 ( .A1(n7698), .A2(n7700), .ZN(n7713) );
  OR2_X1 U9332 ( .A1(n8898), .A2(n8973), .ZN(n7699) );
  AND2_X1 U9333 ( .A1(n7713), .A2(n7699), .ZN(n7745) );
  NAND2_X1 U9334 ( .A1(n7749), .A2(n7745), .ZN(n7705) );
  INV_X1 U9335 ( .A(n7699), .ZN(n7704) );
  AND2_X1 U9336 ( .A1(n7705), .A2(n7746), .ZN(n7706) );
  XOR2_X1 U9337 ( .A(n7753), .B(n7706), .Z(n9529) );
  INV_X1 U9338 ( .A(n9351), .ZN(n9259) );
  NAND2_X1 U9339 ( .A1(n9529), .A2(n9259), .ZN(n7712) );
  OAI22_X1 U9340 ( .A1(n9614), .A2(n7707), .B1(n8791), .B2(n9605), .ZN(n7710)
         );
  INV_X1 U9341 ( .A(n7726), .ZN(n7708) );
  OAI211_X1 U9342 ( .C1(n7708), .C2(n4697), .A(n9503), .B(n7762), .ZN(n9525)
         );
  NOR2_X1 U9343 ( .A1(n9525), .A2(n7767), .ZN(n7709) );
  AOI211_X1 U9344 ( .C1(n9500), .C2(n8793), .A(n7710), .B(n7709), .ZN(n7711)
         );
  OAI211_X1 U9345 ( .C1(n4393), .C2(n9526), .A(n7712), .B(n7711), .ZN(P1_U3277) );
  NAND2_X1 U9346 ( .A1(n7749), .A2(n7713), .ZN(n7715) );
  NAND2_X1 U9347 ( .A1(n7715), .A2(n7714), .ZN(n7716) );
  XNOR2_X1 U9348 ( .A(n7716), .B(n7719), .ZN(n9532) );
  NAND2_X1 U9349 ( .A1(n9532), .A2(n9496), .ZN(n7723) );
  OAI21_X1 U9350 ( .B1(n7719), .B2(n7718), .A(n7717), .ZN(n7721) );
  OAI22_X1 U9351 ( .A1(n8906), .A2(n9491), .B1(n9492), .B2(n7757), .ZN(n7720)
         );
  AOI21_X1 U9352 ( .B1(n7721), .B2(n9308), .A(n7720), .ZN(n7722) );
  NAND2_X1 U9353 ( .A1(n7724), .A2(n8898), .ZN(n7725) );
  NAND2_X1 U9354 ( .A1(n7726), .A2(n7725), .ZN(n9530) );
  OAI22_X1 U9355 ( .A1(n9614), .A2(n6356), .B1(n8907), .B2(n9605), .ZN(n7727)
         );
  AOI21_X1 U9356 ( .B1(n8898), .B2(n9500), .A(n7727), .ZN(n7728) );
  OAI21_X1 U9357 ( .B1(n9530), .B2(n9138), .A(n7728), .ZN(n7729) );
  AOI21_X1 U9358 ( .B1(n9532), .B2(n9508), .A(n7729), .ZN(n7730) );
  OAI21_X1 U9359 ( .B1(n9534), .B2(n4393), .A(n7730), .ZN(P1_U3278) );
  INV_X1 U9360 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7733) );
  AOI21_X1 U9361 ( .B1(n9845), .B2(n7732), .A(n7731), .ZN(n7735) );
  MUX2_X1 U9362 ( .A(n7733), .B(n7735), .S(n9861), .Z(n7734) );
  OAI21_X1 U9363 ( .B1(n7737), .B2(n8754), .A(n7734), .ZN(P2_U3490) );
  MUX2_X1 U9364 ( .A(n10183), .B(n7735), .S(n9879), .Z(n7736) );
  OAI21_X1 U9365 ( .B1(n7737), .B2(n8713), .A(n7736), .ZN(P2_U3533) );
  INV_X1 U9366 ( .A(n7738), .ZN(n7742) );
  OAI222_X1 U9367 ( .A1(n9479), .A2(n7740), .B1(n9473), .B2(n7742), .C1(n7739), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U9368 ( .A1(n8771), .A2(n7743), .B1(n8769), .B2(n7742), .C1(
        P2_U3152), .C2(n7741), .ZN(P2_U3333) );
  NOR2_X1 U9369 ( .A1(n8793), .A2(n8972), .ZN(n7747) );
  INV_X1 U9370 ( .A(n7747), .ZN(n7744) );
  AND2_X1 U9371 ( .A1(n7745), .A2(n7744), .ZN(n7748) );
  AOI21_X1 U9372 ( .B1(n7749), .B2(n7748), .A(n4966), .ZN(n7751) );
  NAND2_X1 U9373 ( .A1(n8793), .A2(n8972), .ZN(n7750) );
  XNOR2_X1 U9374 ( .A(n9086), .B(n7755), .ZN(n9436) );
  INV_X1 U9375 ( .A(n9436), .ZN(n7770) );
  XNOR2_X1 U9376 ( .A(n9109), .B(n7755), .ZN(n7756) );
  NAND2_X1 U9377 ( .A1(n7756), .A2(n9308), .ZN(n7760) );
  OAI22_X1 U9378 ( .A1(n7757), .A2(n9491), .B1(n9492), .B2(n9327), .ZN(n7758)
         );
  INV_X1 U9379 ( .A(n7758), .ZN(n7759) );
  NAND2_X1 U9380 ( .A1(n7760), .A2(n7759), .ZN(n9440) );
  NAND2_X1 U9381 ( .A1(n7762), .A2(n9084), .ZN(n7761) );
  NAND2_X1 U9382 ( .A1(n7761), .A2(n9503), .ZN(n7763) );
  OR2_X1 U9383 ( .A1(n7763), .A2(n9334), .ZN(n9437) );
  OAI22_X1 U9384 ( .A1(n9614), .A2(n7764), .B1(n8964), .B2(n9605), .ZN(n7765)
         );
  AOI21_X1 U9385 ( .B1(n9084), .B2(n9500), .A(n7765), .ZN(n7766) );
  OAI21_X1 U9386 ( .B1(n9437), .B2(n7767), .A(n7766), .ZN(n7768) );
  AOI21_X1 U9387 ( .B1(n9440), .B2(n9614), .A(n7768), .ZN(n7769) );
  OAI21_X1 U9388 ( .B1(n7770), .B2(n9351), .A(n7769), .ZN(P1_U3276) );
  NAND2_X1 U9389 ( .A1(n7772), .A2(n7771), .ZN(n7774) );
  OR2_X1 U9390 ( .A1(n8141), .A2(n8360), .ZN(n7773) );
  NAND2_X1 U9391 ( .A1(n7798), .A2(n8359), .ZN(n8149) );
  XNOR2_X1 U9392 ( .A(n8242), .B(n8241), .ZN(n7780) );
  OR2_X1 U9393 ( .A1(n8141), .A2(n7777), .ZN(n7775) );
  NAND2_X1 U9394 ( .A1(n7776), .A2(n7775), .ZN(n8009) );
  INV_X1 U9395 ( .A(n8241), .ZN(n8056) );
  XNOR2_X1 U9396 ( .A(n8009), .B(n8056), .ZN(n7778) );
  INV_X1 U9397 ( .A(n8358), .ZN(n8601) );
  OAI22_X1 U9398 ( .A1(n7777), .A2(n9745), .B1(n8601), .B2(n9743), .ZN(n7793)
         );
  AOI21_X1 U9399 ( .B1(n7778), .B2(n9774), .A(n7793), .ZN(n7779) );
  OAI21_X1 U9400 ( .B1(n7780), .B2(n9848), .A(n7779), .ZN(n8709) );
  INV_X1 U9401 ( .A(n8709), .ZN(n7787) );
  INV_X1 U9402 ( .A(n7781), .ZN(n7783) );
  INV_X1 U9403 ( .A(n8613), .ZN(n7782) );
  AOI21_X1 U9404 ( .B1(n7798), .B2(n7783), .A(n7782), .ZN(n8710) );
  AOI22_X1 U9405 ( .A1(n4392), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n7792), .B2(
        n9776), .ZN(n7784) );
  OAI21_X1 U9406 ( .B1(n8755), .B2(n9757), .A(n7784), .ZN(n7785) );
  AOI21_X1 U9407 ( .B1(n8710), .B2(n9761), .A(n7785), .ZN(n7786) );
  OAI21_X1 U9408 ( .B1(n7787), .B2(n4392), .A(n7786), .ZN(P2_U3280) );
  INV_X1 U9409 ( .A(n7788), .ZN(n7789) );
  AOI21_X1 U9410 ( .B1(n7791), .B2(n7790), .A(n7789), .ZN(n7800) );
  INV_X1 U9411 ( .A(n7792), .ZN(n7796) );
  AOI22_X1 U9412 ( .A1(n7794), .A2(n7793), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n7795) );
  OAI21_X1 U9413 ( .B1(n8332), .B2(n7796), .A(n7795), .ZN(n7797) );
  AOI21_X1 U9414 ( .B1(n7798), .B2(n8336), .A(n7797), .ZN(n7799) );
  OAI21_X1 U9415 ( .B1(n7800), .B2(n8340), .A(n7799), .ZN(P2_U3228) );
  INV_X1 U9416 ( .A(n7801), .ZN(n7802) );
  NOR2_X1 U9417 ( .A1(n7803), .A2(n7802), .ZN(n7806) );
  NAND2_X1 U9418 ( .A1(n7804), .A2(n9859), .ZN(n7805) );
  NAND2_X1 U9419 ( .A1(n7806), .A2(n7805), .ZN(n7809) );
  MUX2_X1 U9420 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n7809), .S(n9861), .Z(n7807)
         );
  INV_X1 U9421 ( .A(n7807), .ZN(n7808) );
  OAI21_X1 U9422 ( .B1(n8142), .B2(n8754), .A(n7808), .ZN(P2_U3496) );
  MUX2_X1 U9423 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n7809), .S(n9879), .Z(n7810)
         );
  INV_X1 U9424 ( .A(n7810), .ZN(n7811) );
  OAI21_X1 U9425 ( .B1(n8142), .B2(n8713), .A(n7811), .ZN(P2_U3535) );
  XNOR2_X1 U9426 ( .A(n7813), .B(n7812), .ZN(n7818) );
  INV_X1 U9427 ( .A(n8591), .ZN(n8620) );
  AOI22_X1 U9428 ( .A1(n8346), .A2(n8620), .B1(n8344), .B2(n8623), .ZN(n7815)
         );
  OAI211_X1 U9429 ( .C1(n8359), .C2(n8330), .A(n7815), .B(n7814), .ZN(n7816)
         );
  AOI21_X1 U9430 ( .B1(n8706), .B2(n8336), .A(n7816), .ZN(n7817) );
  OAI21_X1 U9431 ( .B1(n7818), .B2(n8340), .A(n7817), .ZN(P2_U3230) );
  INV_X1 U9432 ( .A(n7819), .ZN(n7825) );
  OAI222_X1 U9433 ( .A1(P2_U3152), .A2(n7821), .B1(n8769), .B2(n7825), .C1(
        n7820), .C2(n8771), .ZN(P2_U3332) );
  NAND2_X1 U9434 ( .A1(n8766), .A2(n9474), .ZN(n7823) );
  OAI211_X1 U9435 ( .C1(n9479), .C2(n7824), .A(n7823), .B(n7822), .ZN(P1_U3326) );
  OAI222_X1 U9436 ( .A1(n9479), .A2(n7827), .B1(P1_U3084), .B2(n7826), .C1(
        n9473), .C2(n7825), .ZN(P1_U3327) );
  XNOR2_X1 U9437 ( .A(n7829), .B(n7828), .ZN(n7835) );
  OAI22_X1 U9438 ( .A1(n8330), .A2(n8601), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7830), .ZN(n7833) );
  INV_X1 U9439 ( .A(n8605), .ZN(n7831) );
  OAI22_X1 U9440 ( .A1(n8333), .A2(n8602), .B1(n8332), .B2(n7831), .ZN(n7832)
         );
  AOI211_X1 U9441 ( .C1(n8604), .C2(n8336), .A(n7833), .B(n7832), .ZN(n7834)
         );
  OAI21_X1 U9442 ( .B1(n7835), .B2(n8340), .A(n7834), .ZN(P2_U3240) );
  MUX2_X1 U9443 ( .A(n7836), .B(P1_REG2_REG_3__SCAN_IN), .S(n4393), .Z(n7844)
         );
  NAND2_X1 U9444 ( .A1(n7837), .A2(n9508), .ZN(n7841) );
  OAI22_X1 U9445 ( .A1(n9338), .A2(n7838), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9605), .ZN(n7839) );
  INV_X1 U9446 ( .A(n7839), .ZN(n7840) );
  OAI211_X1 U9447 ( .C1(n9138), .C2(n7842), .A(n7841), .B(n7840), .ZN(n7843)
         );
  OR2_X1 U9448 ( .A1(n7844), .A2(n7843), .ZN(P1_U3288) );
  NAND2_X1 U9449 ( .A1(n8885), .A2(n7991), .ZN(n7850) );
  NAND2_X1 U9450 ( .A1(n7995), .A2(n8977), .ZN(n7849) );
  NAND2_X1 U9451 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  XNOR2_X1 U9452 ( .A(n7851), .B(n7955), .ZN(n7856) );
  NAND2_X1 U9453 ( .A1(n8885), .A2(n7995), .ZN(n7853) );
  NAND2_X1 U9454 ( .A1(n7994), .A2(n8977), .ZN(n7852) );
  NAND2_X1 U9455 ( .A1(n7853), .A2(n7852), .ZN(n7854) );
  XNOR2_X1 U9456 ( .A(n7856), .B(n7854), .ZN(n8878) );
  INV_X1 U9457 ( .A(n7854), .ZN(n7855) );
  NAND2_X1 U9458 ( .A1(n7856), .A2(n7855), .ZN(n7857) );
  NAND2_X1 U9459 ( .A1(n9501), .A2(n7991), .ZN(n7859) );
  NAND2_X1 U9460 ( .A1(n7995), .A2(n8976), .ZN(n7858) );
  NAND2_X1 U9461 ( .A1(n7859), .A2(n7858), .ZN(n7860) );
  XNOR2_X1 U9462 ( .A(n7860), .B(n7955), .ZN(n8807) );
  NAND2_X1 U9463 ( .A1(n9501), .A2(n7995), .ZN(n7862) );
  NAND2_X1 U9464 ( .A1(n7994), .A2(n8976), .ZN(n7861) );
  AND2_X1 U9465 ( .A1(n8807), .A2(n8806), .ZN(n7863) );
  NAND2_X1 U9466 ( .A1(n8930), .A2(n7991), .ZN(n7865) );
  NAND2_X1 U9467 ( .A1(n7995), .A2(n8975), .ZN(n7864) );
  NAND2_X1 U9468 ( .A1(n7865), .A2(n7864), .ZN(n7866) );
  XNOR2_X1 U9469 ( .A(n7866), .B(n7992), .ZN(n7870) );
  NOR2_X1 U9470 ( .A1(n7963), .A2(n9493), .ZN(n7867) );
  AOI21_X1 U9471 ( .B1(n8930), .B2(n7995), .A(n7867), .ZN(n7868) );
  XNOR2_X1 U9472 ( .A(n7870), .B(n7868), .ZN(n8925) );
  INV_X1 U9473 ( .A(n7868), .ZN(n7869) );
  NAND2_X1 U9474 ( .A1(n7870), .A2(n7869), .ZN(n7871) );
  NAND2_X1 U9475 ( .A1(n8837), .A2(n7991), .ZN(n7873) );
  NAND2_X1 U9476 ( .A1(n7995), .A2(n8974), .ZN(n7872) );
  NAND2_X1 U9477 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  XNOR2_X1 U9478 ( .A(n7874), .B(n7955), .ZN(n7876) );
  NOR2_X1 U9479 ( .A1(n7963), .A2(n8906), .ZN(n7875) );
  AOI21_X1 U9480 ( .B1(n8837), .B2(n7995), .A(n7875), .ZN(n7877) );
  NAND2_X1 U9481 ( .A1(n7876), .A2(n7877), .ZN(n7882) );
  INV_X1 U9482 ( .A(n7876), .ZN(n7879) );
  INV_X1 U9483 ( .A(n7877), .ZN(n7878) );
  NAND2_X1 U9484 ( .A1(n7879), .A2(n7878), .ZN(n7880) );
  NAND2_X1 U9485 ( .A1(n7882), .A2(n7880), .ZN(n8832) );
  NAND2_X1 U9486 ( .A1(n8898), .A2(n7991), .ZN(n7884) );
  NAND2_X1 U9487 ( .A1(n7995), .A2(n8973), .ZN(n7883) );
  NAND2_X1 U9488 ( .A1(n7884), .A2(n7883), .ZN(n7885) );
  XNOR2_X1 U9489 ( .A(n7885), .B(n7955), .ZN(n7890) );
  NOR2_X1 U9490 ( .A1(n7963), .A2(n8788), .ZN(n7886) );
  AOI21_X1 U9491 ( .B1(n8898), .B2(n7995), .A(n7886), .ZN(n7891) );
  AND2_X1 U9492 ( .A1(n7890), .A2(n7891), .ZN(n8901) );
  NAND2_X1 U9493 ( .A1(n8793), .A2(n7991), .ZN(n7888) );
  NAND2_X1 U9494 ( .A1(n7995), .A2(n8972), .ZN(n7887) );
  NAND2_X1 U9495 ( .A1(n7888), .A2(n7887), .ZN(n7889) );
  XNOR2_X1 U9496 ( .A(n7889), .B(n7955), .ZN(n7897) );
  INV_X1 U9497 ( .A(n7890), .ZN(n7893) );
  INV_X1 U9498 ( .A(n7891), .ZN(n7892) );
  NAND2_X1 U9499 ( .A1(n7893), .A2(n7892), .ZN(n8899) );
  AND2_X1 U9500 ( .A1(n7897), .A2(n8899), .ZN(n7894) );
  NAND2_X1 U9501 ( .A1(n8904), .A2(n7894), .ZN(n8783) );
  NAND2_X1 U9502 ( .A1(n8793), .A2(n7995), .ZN(n7896) );
  NAND2_X1 U9503 ( .A1(n7994), .A2(n8972), .ZN(n7895) );
  NAND2_X1 U9504 ( .A1(n7896), .A2(n7895), .ZN(n8786) );
  NAND2_X1 U9505 ( .A1(n8783), .A2(n8786), .ZN(n7900) );
  NAND2_X1 U9506 ( .A1(n8904), .A2(n8899), .ZN(n7899) );
  INV_X1 U9507 ( .A(n7897), .ZN(n7898) );
  NAND2_X1 U9508 ( .A1(n7899), .A2(n7898), .ZN(n8784) );
  NAND2_X1 U9509 ( .A1(n7900), .A2(n8784), .ZN(n8958) );
  NAND2_X1 U9510 ( .A1(n9084), .A2(n7991), .ZN(n7902) );
  NAND2_X1 U9511 ( .A1(n7995), .A2(n10214), .ZN(n7901) );
  NAND2_X1 U9512 ( .A1(n7902), .A2(n7901), .ZN(n7903) );
  XNOR2_X1 U9513 ( .A(n7903), .B(n7955), .ZN(n8956) );
  NOR2_X1 U9514 ( .A1(n7963), .A2(n9348), .ZN(n7904) );
  AOI21_X1 U9515 ( .B1(n9084), .B2(n7995), .A(n7904), .ZN(n7906) );
  NAND2_X1 U9516 ( .A1(n8956), .A2(n7906), .ZN(n7905) );
  NAND2_X1 U9517 ( .A1(n8958), .A2(n7905), .ZN(n7909) );
  INV_X1 U9518 ( .A(n8956), .ZN(n7907) );
  INV_X1 U9519 ( .A(n7906), .ZN(n8955) );
  NAND2_X1 U9520 ( .A1(n7907), .A2(n8955), .ZN(n7908) );
  NAND2_X1 U9521 ( .A1(n9431), .A2(n7991), .ZN(n7911) );
  NAND2_X1 U9522 ( .A1(n7995), .A2(n9087), .ZN(n7910) );
  NAND2_X1 U9523 ( .A1(n7911), .A2(n7910), .ZN(n7912) );
  XNOR2_X1 U9524 ( .A(n7912), .B(n7992), .ZN(n7915) );
  NAND2_X1 U9525 ( .A1(n9431), .A2(n7995), .ZN(n7914) );
  NAND2_X1 U9526 ( .A1(n7994), .A2(n9087), .ZN(n7913) );
  NAND2_X1 U9527 ( .A1(n7914), .A2(n7913), .ZN(n7916) );
  INV_X1 U9528 ( .A(n7915), .ZN(n7918) );
  INV_X1 U9529 ( .A(n7916), .ZN(n7917) );
  NAND2_X1 U9530 ( .A1(n7918), .A2(n7917), .ZN(n8849) );
  NAND2_X1 U9531 ( .A1(n9426), .A2(n7991), .ZN(n7920) );
  NAND2_X1 U9532 ( .A1(n7995), .A2(n9304), .ZN(n7919) );
  NAND2_X1 U9533 ( .A1(n7920), .A2(n7919), .ZN(n7921) );
  XNOR2_X1 U9534 ( .A(n7921), .B(n7992), .ZN(n7923) );
  NOR2_X1 U9535 ( .A1(n7963), .A2(n9347), .ZN(n7922) );
  AOI21_X1 U9536 ( .B1(n9426), .B2(n7995), .A(n7922), .ZN(n7924) );
  XNOR2_X1 U9537 ( .A(n7923), .B(n7924), .ZN(n8858) );
  INV_X1 U9538 ( .A(n7923), .ZN(n7925) );
  NAND2_X1 U9539 ( .A1(n9419), .A2(n7991), .ZN(n7927) );
  NAND2_X1 U9540 ( .A1(n7995), .A2(n9288), .ZN(n7926) );
  NAND2_X1 U9541 ( .A1(n7927), .A2(n7926), .ZN(n7928) );
  NOR2_X1 U9542 ( .A1(n7963), .A2(n9328), .ZN(n7929) );
  AOI21_X1 U9543 ( .B1(n9419), .B2(n7995), .A(n7929), .ZN(n8933) );
  NAND2_X1 U9544 ( .A1(n9415), .A2(n7991), .ZN(n7931) );
  NAND2_X1 U9545 ( .A1(n7995), .A2(n9306), .ZN(n7930) );
  NAND2_X1 U9546 ( .A1(n7931), .A2(n7930), .ZN(n7932) );
  XNOR2_X1 U9547 ( .A(n7932), .B(n7992), .ZN(n7934) );
  NOR2_X1 U9548 ( .A1(n7963), .A2(n9276), .ZN(n7933) );
  AOI21_X1 U9549 ( .B1(n9415), .B2(n7995), .A(n7933), .ZN(n7935) );
  XNOR2_X1 U9550 ( .A(n7934), .B(n7935), .ZN(n8815) );
  INV_X1 U9551 ( .A(n7934), .ZN(n7936) );
  NAND2_X1 U9552 ( .A1(n9411), .A2(n7991), .ZN(n7938) );
  NAND2_X1 U9553 ( .A1(n7995), .A2(n9289), .ZN(n7937) );
  NAND2_X1 U9554 ( .A1(n7938), .A2(n7937), .ZN(n7939) );
  XNOR2_X1 U9555 ( .A(n7939), .B(n7955), .ZN(n7942) );
  NOR2_X1 U9556 ( .A1(n9254), .A2(n7963), .ZN(n7940) );
  AOI21_X1 U9557 ( .B1(n9411), .B2(n7995), .A(n7940), .ZN(n7941) );
  NOR2_X1 U9558 ( .A1(n7942), .A2(n7941), .ZN(n8890) );
  NAND2_X1 U9559 ( .A1(n7942), .A2(n7941), .ZN(n8888) );
  NAND2_X1 U9560 ( .A1(n9405), .A2(n7991), .ZN(n7944) );
  NAND2_X1 U9561 ( .A1(n9092), .A2(n7995), .ZN(n7943) );
  NAND2_X1 U9562 ( .A1(n7944), .A2(n7943), .ZN(n7945) );
  XNOR2_X1 U9563 ( .A(n7945), .B(n7992), .ZN(n7946) );
  AOI22_X1 U9564 ( .A1(n9405), .A2(n7995), .B1(n7994), .B2(n9092), .ZN(n7947)
         );
  XNOR2_X1 U9565 ( .A(n7946), .B(n7947), .ZN(n8822) );
  INV_X1 U9566 ( .A(n7946), .ZN(n7948) );
  OAI22_X1 U9567 ( .A1(n9244), .A2(n7848), .B1(n9255), .B2(n7963), .ZN(n7950)
         );
  AOI22_X1 U9568 ( .A1(n9399), .A2(n7991), .B1(n7990), .B2(n9228), .ZN(n7949)
         );
  XNOR2_X1 U9569 ( .A(n7949), .B(n7992), .ZN(n8913) );
  AOI22_X1 U9570 ( .A1(n9392), .A2(n7991), .B1(n7990), .B2(n8971), .ZN(n7952)
         );
  NAND2_X1 U9571 ( .A1(n9389), .A2(n7991), .ZN(n7954) );
  NAND2_X1 U9572 ( .A1(n9229), .A2(n7990), .ZN(n7953) );
  NAND2_X1 U9573 ( .A1(n7954), .A2(n7953), .ZN(n7956) );
  XNOR2_X1 U9574 ( .A(n7956), .B(n7955), .ZN(n7958) );
  AND2_X1 U9575 ( .A1(n9229), .A2(n7994), .ZN(n7957) );
  AOI21_X1 U9576 ( .B1(n9389), .B2(n7995), .A(n7957), .ZN(n7959) );
  NAND2_X1 U9577 ( .A1(n7958), .A2(n7959), .ZN(n7965) );
  INV_X1 U9578 ( .A(n7958), .ZN(n7961) );
  INV_X1 U9579 ( .A(n7959), .ZN(n7960) );
  NAND2_X1 U9580 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  AND2_X1 U9581 ( .A1(n8868), .A2(n8866), .ZN(n7964) );
  OAI22_X1 U9582 ( .A1(n9225), .A2(n7848), .B1(n9238), .B2(n7963), .ZN(n8798)
         );
  NAND2_X1 U9583 ( .A1(n8796), .A2(n8798), .ZN(n8867) );
  NAND2_X1 U9584 ( .A1(n7964), .A2(n8867), .ZN(n8865) );
  NAND2_X1 U9585 ( .A1(n9382), .A2(n7991), .ZN(n7967) );
  NAND2_X1 U9586 ( .A1(n9185), .A2(n7995), .ZN(n7966) );
  NAND2_X1 U9587 ( .A1(n7967), .A2(n7966), .ZN(n7968) );
  XNOR2_X1 U9588 ( .A(n7968), .B(n7992), .ZN(n7973) );
  AOI22_X1 U9589 ( .A1(n9382), .A2(n7995), .B1(n7994), .B2(n9185), .ZN(n7974)
         );
  XNOR2_X1 U9590 ( .A(n7973), .B(n7974), .ZN(n8842) );
  NAND2_X1 U9591 ( .A1(n9377), .A2(n7991), .ZN(n7970) );
  NAND2_X1 U9592 ( .A1(n9201), .A2(n7990), .ZN(n7969) );
  NAND2_X1 U9593 ( .A1(n7970), .A2(n7969), .ZN(n7971) );
  XNOR2_X1 U9594 ( .A(n7971), .B(n7992), .ZN(n7986) );
  AND2_X1 U9595 ( .A1(n9201), .A2(n7994), .ZN(n7972) );
  AOI21_X1 U9596 ( .B1(n9377), .B2(n7995), .A(n7972), .ZN(n7984) );
  XNOR2_X1 U9597 ( .A(n7986), .B(n7984), .ZN(n8945) );
  INV_X1 U9598 ( .A(n7973), .ZN(n7975) );
  NAND2_X1 U9599 ( .A1(n7975), .A2(n7974), .ZN(n8942) );
  NAND2_X1 U9600 ( .A1(n9373), .A2(n7991), .ZN(n7978) );
  NAND2_X1 U9601 ( .A1(n7990), .A2(n9186), .ZN(n7977) );
  NAND2_X1 U9602 ( .A1(n7978), .A2(n7977), .ZN(n7979) );
  XNOR2_X1 U9603 ( .A(n7979), .B(n7992), .ZN(n7983) );
  NAND2_X1 U9604 ( .A1(n9373), .A2(n6825), .ZN(n7981) );
  NAND2_X1 U9605 ( .A1(n7994), .A2(n9186), .ZN(n7980) );
  NAND2_X1 U9606 ( .A1(n7981), .A2(n7980), .ZN(n7982) );
  NOR2_X1 U9607 ( .A1(n7983), .A2(n7982), .ZN(n7988) );
  AOI21_X1 U9608 ( .B1(n7983), .B2(n7982), .A(n7988), .ZN(n8775) );
  INV_X1 U9609 ( .A(n7984), .ZN(n7985) );
  NAND2_X1 U9610 ( .A1(n7986), .A2(n7985), .ZN(n8776) );
  INV_X1 U9611 ( .A(n7988), .ZN(n7989) );
  NAND2_X1 U9612 ( .A1(n8774), .A2(n7989), .ZN(n7999) );
  AOI22_X1 U9613 ( .A1(n9367), .A2(n7991), .B1(n7990), .B2(n9132), .ZN(n7993)
         );
  XNOR2_X1 U9614 ( .A(n7993), .B(n7992), .ZN(n7997) );
  AOI22_X1 U9615 ( .A1(n9367), .A2(n7995), .B1(n7994), .B2(n9132), .ZN(n7996)
         );
  XNOR2_X1 U9616 ( .A(n7997), .B(n7996), .ZN(n7998) );
  XNOR2_X1 U9617 ( .A(n7999), .B(n7998), .ZN(n8004) );
  AOI22_X1 U9618 ( .A1(n8962), .A2(n9186), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8001) );
  NAND2_X1 U9619 ( .A1(n8921), .A2(n9155), .ZN(n8000) );
  OAI211_X1 U9620 ( .C1(n8965), .C2(n9149), .A(n8001), .B(n8000), .ZN(n8002)
         );
  AOI21_X1 U9621 ( .B1(n9367), .B2(n8967), .A(n8002), .ZN(n8003) );
  OAI21_X1 U9622 ( .B1(n8004), .B2(n8969), .A(n8003), .ZN(P1_U3218) );
  INV_X1 U9623 ( .A(n8022), .ZN(n8239) );
  OAI222_X1 U9624 ( .A1(n9468), .A2(n8006), .B1(n9473), .B2(n8239), .C1(n8005), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  NAND2_X1 U9625 ( .A1(n8009), .A2(n8149), .ZN(n8010) );
  NAND2_X1 U9626 ( .A1(n8010), .A2(n8147), .ZN(n8617) );
  NAND2_X1 U9627 ( .A1(n8617), .A2(n8618), .ZN(n8011) );
  OR2_X1 U9628 ( .A1(n8706), .A2(n8601), .ZN(n8148) );
  NAND2_X1 U9629 ( .A1(n8604), .A2(n8591), .ZN(n8164) );
  OR2_X1 U9630 ( .A1(n8696), .A2(n8602), .ZN(n8165) );
  NAND2_X1 U9631 ( .A1(n8696), .A2(n8602), .ZN(n8564) );
  NAND2_X1 U9632 ( .A1(n8165), .A2(n8564), .ZN(n8589) );
  NAND2_X1 U9633 ( .A1(n8689), .A2(n8592), .ZN(n8168) );
  NAND2_X1 U9634 ( .A1(n8013), .A2(n8168), .ZN(n8245) );
  INV_X1 U9635 ( .A(n8564), .ZN(n8012) );
  INV_X1 U9636 ( .A(n8013), .ZN(n8171) );
  XNOR2_X1 U9637 ( .A(n8559), .B(n8567), .ZN(n8547) );
  AND2_X2 U9638 ( .A1(n8545), .A2(n8547), .ZN(n8550) );
  INV_X1 U9639 ( .A(n8567), .ZN(n8329) );
  AND2_X1 U9640 ( .A1(n8559), .A2(n8329), .ZN(n8530) );
  NAND2_X1 U9641 ( .A1(n8537), .A2(n8551), .ZN(n8162) );
  NAND2_X1 U9642 ( .A1(n8515), .A2(n8162), .ZN(n8529) );
  INV_X1 U9643 ( .A(n8515), .ZN(n8179) );
  OR2_X1 U9644 ( .A1(n8674), .A2(n8535), .ZN(n8180) );
  NAND2_X1 U9645 ( .A1(n8674), .A2(n8535), .ZN(n8181) );
  NAND2_X1 U9646 ( .A1(n8180), .A2(n8181), .ZN(n8512) );
  INV_X1 U9647 ( .A(n8181), .ZN(n8497) );
  NAND2_X1 U9648 ( .A1(n8505), .A2(n8518), .ZN(n8185) );
  NAND2_X1 U9649 ( .A1(n8184), .A2(n8185), .ZN(n8041) );
  INV_X1 U9650 ( .A(n8184), .ZN(n8015) );
  NAND2_X1 U9651 ( .A1(n8664), .A2(n8501), .ZN(n8189) );
  NAND2_X1 U9652 ( .A1(n8477), .A2(n8487), .ZN(n8017) );
  NAND2_X1 U9653 ( .A1(n8652), .A2(n8471), .ZN(n8198) );
  INV_X1 U9654 ( .A(n8017), .ZN(n8457) );
  NAND2_X1 U9655 ( .A1(n8442), .A2(n8249), .ZN(n8199) );
  INV_X1 U9656 ( .A(n8435), .ZN(n8021) );
  NAND2_X1 U9657 ( .A1(n8760), .A2(n6204), .ZN(n8020) );
  NAND2_X1 U9658 ( .A1(n6119), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U9659 ( .A1(n8643), .A2(n8438), .ZN(n8205) );
  NAND3_X1 U9660 ( .A1(n8021), .A2(n4641), .A3(n8256), .ZN(n8259) );
  NAND2_X1 U9661 ( .A1(n8259), .A2(n8205), .ZN(n8029) );
  INV_X1 U9662 ( .A(n8029), .ZN(n8031) );
  NAND2_X1 U9663 ( .A1(n8022), .A2(n6204), .ZN(n8024) );
  NAND2_X1 U9664 ( .A1(n6119), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8023) );
  INV_X1 U9665 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U9666 ( .A1(n8025), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8027) );
  NAND2_X1 U9667 ( .A1(n6506), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8026) );
  OAI211_X1 U9668 ( .C1(n8028), .C2(n8641), .A(n8027), .B(n8026), .ZN(n8352)
         );
  OAI211_X1 U9669 ( .C1(n8029), .C2(n8429), .A(n8423), .B(n8223), .ZN(n8030)
         );
  OAI21_X1 U9670 ( .B1(n8031), .B2(n8211), .A(n8030), .ZN(n8036) );
  NAND2_X1 U9671 ( .A1(n8032), .A2(n6204), .ZN(n8034) );
  NAND2_X1 U9672 ( .A1(n6119), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8033) );
  INV_X1 U9673 ( .A(n8352), .ZN(n8035) );
  NAND2_X1 U9674 ( .A1(n8429), .A2(n8035), .ZN(n8210) );
  NAND2_X1 U9675 ( .A1(n8215), .A2(n8210), .ZN(n8213) );
  NAND2_X1 U9676 ( .A1(n8421), .A2(n8423), .ZN(n8216) );
  XNOR2_X1 U9677 ( .A(n8037), .B(n4394), .ZN(n8231) );
  NAND2_X1 U9678 ( .A1(n8039), .A2(n8038), .ZN(n8230) );
  INV_X1 U9679 ( .A(n8211), .ZN(n8040) );
  NAND2_X1 U9680 ( .A1(n8216), .A2(n8040), .ZN(n8212) );
  INV_X1 U9681 ( .A(n8436), .ZN(n8062) );
  NAND2_X1 U9682 ( .A1(n9769), .A2(n8042), .ZN(n8044) );
  NOR4_X1 U9683 ( .A1(n8044), .A2(n9738), .A3(n8043), .A4(n8226), .ZN(n8047)
         );
  NAND4_X1 U9684 ( .A1(n8047), .A2(n7021), .A3(n8046), .A4(n8086), .ZN(n8049)
         );
  NOR4_X1 U9685 ( .A1(n8049), .A2(n8048), .A3(n9728), .A4(n8102), .ZN(n8050)
         );
  NAND4_X1 U9686 ( .A1(n8053), .A2(n8052), .A3(n8051), .A4(n8050), .ZN(n8054)
         );
  NOR4_X1 U9687 ( .A1(n8056), .A2(n8055), .A3(n8135), .A4(n8054), .ZN(n8057)
         );
  NAND4_X1 U9688 ( .A1(n8599), .A2(n8057), .A3(n8618), .A4(n8139), .ZN(n8058)
         );
  NOR4_X1 U9689 ( .A1(n8529), .A2(n8589), .A3(n8245), .A4(n8058), .ZN(n8059)
         );
  NAND4_X1 U9690 ( .A1(n8498), .A2(n4942), .A3(n8059), .A4(n8547), .ZN(n8060)
         );
  NOR4_X1 U9691 ( .A1(n8458), .A2(n8469), .A3(n8484), .A4(n8060), .ZN(n8061)
         );
  NAND3_X1 U9692 ( .A1(n4641), .A2(n8062), .A3(n8061), .ZN(n8063) );
  NOR3_X1 U9693 ( .A1(n8213), .A2(n8212), .A3(n8063), .ZN(n8064) );
  XNOR2_X1 U9694 ( .A(n8064), .B(n4394), .ZN(n8222) );
  INV_X1 U9695 ( .A(n8204), .ZN(n8207) );
  INV_X1 U9696 ( .A(n8214), .ZN(n8197) );
  INV_X1 U9697 ( .A(n8065), .ZN(n9739) );
  NAND2_X1 U9698 ( .A1(n8069), .A2(n8068), .ZN(n8067) );
  NAND2_X1 U9699 ( .A1(n8091), .A2(n8094), .ZN(n8066) );
  MUX2_X1 U9700 ( .A(n8067), .B(n8066), .S(n8214), .Z(n8095) );
  AOI21_X1 U9701 ( .B1(n8068), .B2(n9739), .A(n8095), .ZN(n8072) );
  INV_X1 U9702 ( .A(n8101), .ZN(n8071) );
  INV_X1 U9703 ( .A(n8069), .ZN(n8070) );
  NOR3_X1 U9704 ( .A1(n8072), .A2(n8071), .A3(n8070), .ZN(n8090) );
  INV_X1 U9705 ( .A(n8080), .ZN(n8075) );
  INV_X1 U9706 ( .A(n8078), .ZN(n8074) );
  OAI211_X1 U9707 ( .C1(n8075), .C2(n8074), .A(n8081), .B(n8073), .ZN(n8076)
         );
  NAND2_X1 U9708 ( .A1(n8076), .A2(n8079), .ZN(n8085) );
  AOI21_X1 U9709 ( .B1(n8223), .B2(n8078), .A(n8077), .ZN(n8083) );
  NAND2_X1 U9710 ( .A1(n8080), .A2(n8079), .ZN(n8082) );
  OAI21_X1 U9711 ( .B1(n8083), .B2(n8082), .A(n8081), .ZN(n8084) );
  MUX2_X1 U9712 ( .A(n8085), .B(n8084), .S(n8214), .Z(n8088) );
  INV_X1 U9713 ( .A(n8095), .ZN(n8087) );
  NAND3_X1 U9714 ( .A1(n8088), .A2(n8087), .A3(n8086), .ZN(n8089) );
  OAI21_X1 U9715 ( .B1(n8090), .B2(n8197), .A(n8089), .ZN(n8099) );
  INV_X1 U9716 ( .A(n8091), .ZN(n8092) );
  AOI21_X1 U9717 ( .B1(n8093), .B2(n9772), .A(n8092), .ZN(n8096) );
  OAI211_X1 U9718 ( .C1(n8096), .C2(n8095), .A(n8094), .B(n8098), .ZN(n8097)
         );
  AOI22_X1 U9719 ( .A1(n8099), .A2(n8098), .B1(n8197), .B2(n8097), .ZN(n8107)
         );
  OAI21_X1 U9720 ( .B1(n8101), .B2(n8214), .A(n8100), .ZN(n8106) );
  NAND2_X1 U9721 ( .A1(n9727), .A2(n8214), .ZN(n8104) );
  NAND2_X1 U9722 ( .A1(n9828), .A2(n8197), .ZN(n8103) );
  MUX2_X1 U9723 ( .A(n8104), .B(n8103), .S(n8368), .Z(n8105) );
  OAI211_X1 U9724 ( .C1(n8107), .C2(n8106), .A(n7111), .B(n8105), .ZN(n8111)
         );
  MUX2_X1 U9725 ( .A(n8109), .B(n8108), .S(n8214), .Z(n8110) );
  NAND3_X1 U9726 ( .A1(n8111), .A2(n8112), .A3(n8110), .ZN(n8115) );
  INV_X1 U9727 ( .A(n8118), .ZN(n8113) );
  OAI21_X1 U9728 ( .B1(n8113), .B2(n4793), .A(n8214), .ZN(n8114) );
  NAND4_X1 U9729 ( .A1(n8115), .A2(n8119), .A3(n8116), .A4(n8114), .ZN(n8126)
         );
  AND2_X1 U9730 ( .A1(n8128), .A2(n8118), .ZN(n8124) );
  INV_X1 U9731 ( .A(n8116), .ZN(n8117) );
  NAND2_X1 U9732 ( .A1(n8118), .A2(n8117), .ZN(n8120) );
  NAND2_X1 U9733 ( .A1(n8120), .A2(n8119), .ZN(n8121) );
  NOR2_X1 U9734 ( .A1(n8122), .A2(n8121), .ZN(n8123) );
  MUX2_X1 U9735 ( .A(n8124), .B(n8123), .S(n8214), .Z(n8125) );
  MUX2_X1 U9736 ( .A(n8132), .B(n8131), .S(n8214), .Z(n8133) );
  MUX2_X1 U9737 ( .A(n8137), .B(n8136), .S(n8214), .Z(n8138) );
  NAND3_X1 U9738 ( .A1(n8140), .A2(n8139), .A3(n8138), .ZN(n8146) );
  NAND2_X1 U9739 ( .A1(n8141), .A2(n8214), .ZN(n8144) );
  NAND2_X1 U9740 ( .A1(n8142), .A2(n8197), .ZN(n8143) );
  MUX2_X1 U9741 ( .A(n8144), .B(n8143), .S(n8360), .Z(n8145) );
  INV_X1 U9742 ( .A(n8148), .ZN(n8154) );
  INV_X1 U9743 ( .A(n8706), .ZN(n8152) );
  INV_X1 U9744 ( .A(n8149), .ZN(n8150) );
  NAND2_X1 U9745 ( .A1(n8618), .A2(n8150), .ZN(n8151) );
  OAI211_X1 U9746 ( .C1(n8152), .C2(n8358), .A(n8151), .B(n8164), .ZN(n8153)
         );
  MUX2_X1 U9747 ( .A(n8154), .B(n8153), .S(n8197), .Z(n8155) );
  NAND3_X1 U9748 ( .A1(n8157), .A2(n8156), .A3(n8165), .ZN(n8158) );
  AOI21_X1 U9749 ( .B1(n8158), .B2(n8564), .A(n8171), .ZN(n8160) );
  INV_X1 U9750 ( .A(n8168), .ZN(n8159) );
  OR2_X1 U9751 ( .A1(n8559), .A2(n8329), .ZN(n8170) );
  OAI21_X1 U9752 ( .B1(n8160), .B2(n8159), .A(n8170), .ZN(n8163) );
  INV_X1 U9753 ( .A(n8530), .ZN(n8161) );
  AND2_X1 U9754 ( .A1(n8162), .A2(n8161), .ZN(n8173) );
  AOI21_X1 U9755 ( .B1(n8163), .B2(n8173), .A(n8179), .ZN(n8178) );
  INV_X1 U9756 ( .A(n8164), .ZN(n8166) );
  OAI21_X1 U9757 ( .B1(n8167), .B2(n8166), .A(n8165), .ZN(n8169) );
  NAND3_X1 U9758 ( .A1(n8169), .A2(n8564), .A3(n8168), .ZN(n8176) );
  INV_X1 U9759 ( .A(n8170), .ZN(n8172) );
  NOR2_X1 U9760 ( .A1(n8172), .A2(n8171), .ZN(n8175) );
  INV_X1 U9761 ( .A(n8173), .ZN(n8174) );
  AOI21_X1 U9762 ( .B1(n8176), .B2(n8175), .A(n8174), .ZN(n8177) );
  NAND2_X1 U9763 ( .A1(n8498), .A2(n8180), .ZN(n8183) );
  NAND2_X1 U9764 ( .A1(n8185), .A2(n8181), .ZN(n8182) );
  MUX2_X1 U9765 ( .A(n8183), .B(n8182), .S(n8214), .Z(n8188) );
  INV_X1 U9766 ( .A(n8484), .ZN(n8187) );
  MUX2_X1 U9767 ( .A(n8185), .B(n8184), .S(n8214), .Z(n8186) );
  INV_X1 U9768 ( .A(n8189), .ZN(n8190) );
  OAI21_X1 U9769 ( .B1(n8469), .B2(n8190), .A(n8214), .ZN(n8191) );
  AOI21_X1 U9770 ( .B1(n8194), .B2(n8192), .A(n8214), .ZN(n8193) );
  AOI21_X1 U9771 ( .B1(n8195), .B2(n8194), .A(n8193), .ZN(n8196) );
  AOI211_X1 U9772 ( .C1(n8457), .C2(n8197), .A(n8458), .B(n8196), .ZN(n8203)
         );
  NAND2_X1 U9773 ( .A1(n8199), .A2(n8198), .ZN(n8200) );
  MUX2_X1 U9774 ( .A(n8201), .B(n8200), .S(n8214), .Z(n8202) );
  NOR2_X1 U9775 ( .A1(n8203), .A2(n8202), .ZN(n8209) );
  NAND2_X1 U9776 ( .A1(n8204), .A2(n8249), .ZN(n8206) );
  MUX2_X1 U9777 ( .A(n8214), .B(n8249), .S(n8442), .Z(n8208) );
  MUX2_X1 U9778 ( .A(n8213), .B(n8212), .S(n8214), .Z(n8218) );
  MUX2_X1 U9779 ( .A(n8216), .B(n8215), .S(n8214), .Z(n8217) );
  INV_X1 U9780 ( .A(n8219), .ZN(n8220) );
  OAI21_X1 U9781 ( .B1(n8227), .B2(n8220), .A(n8226), .ZN(n8221) );
  OAI21_X1 U9782 ( .B1(n8223), .B2(n8222), .A(n8221), .ZN(n8229) );
  INV_X1 U9783 ( .A(n8224), .ZN(n8225) );
  NAND3_X1 U9784 ( .A1(n8227), .A2(n8226), .A3(n8225), .ZN(n8228) );
  AOI21_X1 U9785 ( .B1(n8231), .B2(n8230), .A(n4971), .ZN(n8238) );
  INV_X1 U9786 ( .A(n8767), .ZN(n8262) );
  NAND4_X1 U9787 ( .A1(n8233), .A2(n8262), .A3(n8232), .A4(n9770), .ZN(n8234)
         );
  OAI211_X1 U9788 ( .C1(n8235), .C2(n8237), .A(n8234), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8236) );
  OAI21_X1 U9789 ( .B1(n8238), .B2(n8237), .A(n8236), .ZN(P2_U3244) );
  INV_X1 U9790 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9960) );
  OAI222_X1 U9791 ( .A1(P2_U3152), .A2(n8240), .B1(n8769), .B2(n8239), .C1(
        n9960), .C2(n8771), .ZN(P2_U3328) );
  INV_X1 U9792 ( .A(n8471), .ZN(n8353) );
  INV_X1 U9793 ( .A(n8487), .ZN(n8461) );
  OR2_X1 U9794 ( .A1(n8706), .A2(n8358), .ZN(n8243) );
  NOR2_X1 U9795 ( .A1(n8604), .A2(n8620), .ZN(n8244) );
  INV_X1 U9796 ( .A(n8604), .ZN(n8749) );
  INV_X1 U9797 ( .A(n8602), .ZN(n8566) );
  OR2_X2 U9798 ( .A1(n8572), .A2(n8571), .ZN(n8688) );
  INV_X1 U9799 ( .A(n8592), .ZN(n8357) );
  NAND2_X1 U9800 ( .A1(n8689), .A2(n8357), .ZN(n8246) );
  NAND2_X2 U9801 ( .A1(n8688), .A2(n8246), .ZN(n8546) );
  INV_X1 U9802 ( .A(n8559), .ZN(n8743) );
  NAND2_X1 U9803 ( .A1(n8743), .A2(n8329), .ZN(n8247) );
  INV_X1 U9804 ( .A(n8518), .ZN(n8356) );
  NAND2_X1 U9805 ( .A1(n8482), .A2(n8484), .ZN(n8481) );
  NAND2_X1 U9806 ( .A1(n8481), .A2(n8248), .ZN(n8466) );
  NOR2_X1 U9807 ( .A1(n8611), .A2(n8604), .ZN(n8603) );
  INV_X1 U9808 ( .A(n8696), .ZN(n8250) );
  INV_X1 U9809 ( .A(n8689), .ZN(n8570) );
  INV_X1 U9810 ( .A(n8505), .ZN(n8734) );
  INV_X1 U9811 ( .A(n8441), .ZN(n8251) );
  INV_X1 U9812 ( .A(n8643), .ZN(n8255) );
  AOI21_X1 U9813 ( .B1(n8643), .B2(n8251), .A(n8428), .ZN(n8644) );
  INV_X1 U9814 ( .A(n8252), .ZN(n8253) );
  AOI22_X1 U9815 ( .A1(n8253), .A2(n9776), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n4392), .ZN(n8254) );
  OAI21_X1 U9816 ( .B1(n8255), .B2(n9757), .A(n8254), .ZN(n8267) );
  INV_X1 U9817 ( .A(n8256), .ZN(n8258) );
  OAI21_X1 U9818 ( .B1(n8435), .B2(n8258), .A(n8257), .ZN(n8260) );
  NAND2_X1 U9819 ( .A1(n8260), .A2(n8259), .ZN(n8261) );
  AOI21_X1 U9820 ( .B1(n8262), .B2(P2_B_REG_SCAN_IN), .A(n9743), .ZN(n8422) );
  AND2_X1 U9821 ( .A1(n8352), .A2(n8422), .ZN(n8263) );
  OAI21_X1 U9822 ( .B1(n8647), .B2(n9755), .A(n8268), .ZN(P2_U3267) );
  OAI222_X1 U9823 ( .A1(n9473), .A2(n8269), .B1(n9468), .B2(n5183), .C1(n5619), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  AOI21_X1 U9824 ( .B1(n8271), .B2(n8270), .A(n8340), .ZN(n8272) );
  NAND2_X1 U9825 ( .A1(n8273), .A2(n8272), .ZN(n8277) );
  AOI22_X1 U9826 ( .A1(n8343), .A2(n8461), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8276) );
  AOI22_X1 U9827 ( .A1(n8460), .A2(n8346), .B1(n8455), .B2(n8344), .ZN(n8275)
         );
  NAND2_X1 U9828 ( .A1(n8652), .A2(n8336), .ZN(n8274) );
  NAND4_X1 U9829 ( .A1(n8277), .A2(n8276), .A3(n8275), .A4(n8274), .ZN(
        P2_U3216) );
  XOR2_X1 U9830 ( .A(n8279), .B(n8278), .Z(n8284) );
  OAI22_X1 U9831 ( .A1(n8330), .A2(n8551), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8280), .ZN(n8282) );
  OAI22_X1 U9832 ( .A1(n8333), .A2(n8518), .B1(n8332), .B2(n8521), .ZN(n8281)
         );
  AOI211_X1 U9833 ( .C1(n8674), .C2(n8336), .A(n8282), .B(n8281), .ZN(n8283)
         );
  OAI21_X1 U9834 ( .B1(n8284), .B2(n8340), .A(n8283), .ZN(P2_U3218) );
  INV_X1 U9835 ( .A(n8285), .ZN(n8286) );
  AOI21_X1 U9836 ( .B1(n8288), .B2(n8287), .A(n8286), .ZN(n8292) );
  NAND2_X1 U9837 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8416) );
  OAI21_X1 U9838 ( .B1(n8330), .B2(n8591), .A(n8416), .ZN(n8290) );
  OAI22_X1 U9839 ( .A1(n8333), .A2(n8592), .B1(n8332), .B2(n8582), .ZN(n8289)
         );
  AOI211_X1 U9840 ( .C1(n8696), .C2(n8336), .A(n8290), .B(n8289), .ZN(n8291)
         );
  OAI21_X1 U9841 ( .B1(n8292), .B2(n8340), .A(n8291), .ZN(P2_U3221) );
  OR2_X1 U9842 ( .A1(n8319), .A2(n8318), .ZN(n8294) );
  NAND2_X1 U9843 ( .A1(n8294), .A2(n8293), .ZN(n8296) );
  XNOR2_X1 U9844 ( .A(n8296), .B(n8295), .ZN(n8301) );
  OAI22_X1 U9845 ( .A1(n8330), .A2(n8592), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8297), .ZN(n8299) );
  OAI22_X1 U9846 ( .A1(n8333), .A2(n8551), .B1(n8332), .B2(n8557), .ZN(n8298)
         );
  AOI211_X1 U9847 ( .C1(n8559), .C2(n8336), .A(n8299), .B(n8298), .ZN(n8300)
         );
  OAI21_X1 U9848 ( .B1(n8301), .B2(n8340), .A(n8300), .ZN(P2_U3225) );
  XNOR2_X1 U9849 ( .A(n8303), .B(n8302), .ZN(n8304) );
  XNOR2_X1 U9850 ( .A(n8305), .B(n8304), .ZN(n8310) );
  OAI22_X1 U9851 ( .A1(n8333), .A2(n8487), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9935), .ZN(n8308) );
  INV_X1 U9852 ( .A(n8306), .ZN(n8489) );
  OAI22_X1 U9853 ( .A1(n8330), .A2(n8518), .B1(n8332), .B2(n8489), .ZN(n8307)
         );
  AOI211_X1 U9854 ( .C1(n8664), .C2(n8336), .A(n8308), .B(n8307), .ZN(n8309)
         );
  OAI21_X1 U9855 ( .B1(n8310), .B2(n8340), .A(n8309), .ZN(P2_U3227) );
  XNOR2_X1 U9856 ( .A(n8311), .B(n8312), .ZN(n8317) );
  OAI22_X1 U9857 ( .A1(n8330), .A2(n8535), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8313), .ZN(n8315) );
  OAI22_X1 U9858 ( .A1(n8333), .A2(n8501), .B1(n8332), .B2(n8503), .ZN(n8314)
         );
  AOI211_X1 U9859 ( .C1(n8505), .C2(n8336), .A(n8315), .B(n8314), .ZN(n8316)
         );
  OAI21_X1 U9860 ( .B1(n8317), .B2(n8340), .A(n8316), .ZN(P2_U3231) );
  XNOR2_X1 U9861 ( .A(n8319), .B(n8318), .ZN(n8324) );
  OAI22_X1 U9862 ( .A1(n8330), .A2(n8602), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8320), .ZN(n8322) );
  OAI22_X1 U9863 ( .A1(n8333), .A2(n8329), .B1(n8332), .B2(n8573), .ZN(n8321)
         );
  AOI211_X1 U9864 ( .C1(n8689), .C2(n8336), .A(n8322), .B(n8321), .ZN(n8323)
         );
  OAI21_X1 U9865 ( .B1(n8324), .B2(n8340), .A(n8323), .ZN(P2_U3235) );
  AOI21_X1 U9866 ( .B1(n8327), .B2(n8326), .A(n8325), .ZN(n8338) );
  OAI22_X1 U9867 ( .A1(n8330), .A2(n8329), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8328), .ZN(n8335) );
  INV_X1 U9868 ( .A(n8538), .ZN(n8331) );
  OAI22_X1 U9869 ( .A1(n8333), .A2(n8535), .B1(n8332), .B2(n8331), .ZN(n8334)
         );
  AOI211_X1 U9870 ( .C1(n8537), .C2(n8336), .A(n8335), .B(n8334), .ZN(n8337)
         );
  OAI21_X1 U9871 ( .B1(n8338), .B2(n8340), .A(n8337), .ZN(P2_U3237) );
  AOI22_X1 U9872 ( .A1(n8343), .A2(n8355), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8348) );
  INV_X1 U9873 ( .A(n8474), .ZN(n8345) );
  AOI22_X1 U9874 ( .A1(n8353), .A2(n8346), .B1(n8345), .B2(n8344), .ZN(n8347)
         );
  OAI211_X1 U9875 ( .C1(n8729), .C2(n8349), .A(n8348), .B(n8347), .ZN(n8350)
         );
  OR2_X1 U9876 ( .A1(n8351), .A2(n8350), .ZN(P2_U3242) );
  MUX2_X1 U9877 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8352), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9878 ( .A(n8460), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8354), .Z(
        P2_U3580) );
  MUX2_X1 U9879 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8353), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9880 ( .A(n8461), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8354), .Z(
        P2_U3578) );
  MUX2_X1 U9881 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8355), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9882 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8356), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9883 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8357), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9884 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8566), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9885 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8620), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9886 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8358), .S(P2_U3966), .Z(
        P2_U3569) );
  INV_X1 U9887 ( .A(n8359), .ZN(n8619) );
  MUX2_X1 U9888 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8619), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9889 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8360), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9890 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8361), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9891 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8362), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9892 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8363), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9893 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8364), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9894 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8365), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9895 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8366), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9896 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8367), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9897 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8368), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9898 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8369), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9899 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8370), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9900 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8371), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9901 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n9772), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9902 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8372), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9903 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6891), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9904 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6649), .S(P2_U3966), .Z(
        P2_U3552) );
  NAND3_X1 U9905 ( .A1(n8375), .A2(n8374), .A3(n8373), .ZN(n8376) );
  NAND3_X1 U9906 ( .A1(n9715), .A2(n8377), .A3(n8376), .ZN(n8388) );
  AOI22_X1 U9907 ( .A1(n9707), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n8387) );
  NAND2_X1 U9908 ( .A1(n9709), .A2(n8378), .ZN(n8386) );
  MUX2_X1 U9909 ( .A(n6469), .B(P2_REG1_REG_2__SCAN_IN), .S(n8378), .Z(n8381)
         );
  INV_X1 U9910 ( .A(n8379), .ZN(n8380) );
  NAND2_X1 U9911 ( .A1(n8381), .A2(n8380), .ZN(n8383) );
  OAI211_X1 U9912 ( .C1(n8384), .C2(n8383), .A(n9711), .B(n8382), .ZN(n8385)
         );
  NAND4_X1 U9913 ( .A1(n8388), .A2(n8387), .A3(n8386), .A4(n8385), .ZN(
        P2_U3247) );
  MUX2_X1 U9914 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8389), .S(n8394), .Z(n8391)
         );
  OAI211_X1 U9915 ( .C1(n8392), .C2(n8391), .A(n8390), .B(n9715), .ZN(n8403)
         );
  AOI21_X1 U9916 ( .B1(n9707), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8393), .ZN(
        n8402) );
  NAND2_X1 U9917 ( .A1(n9709), .A2(n8394), .ZN(n8401) );
  INV_X1 U9918 ( .A(n8395), .ZN(n8396) );
  OAI21_X1 U9919 ( .B1(n8398), .B2(n8397), .A(n8396), .ZN(n8399) );
  NAND2_X1 U9920 ( .A1(n9711), .A2(n8399), .ZN(n8400) );
  NAND4_X1 U9921 ( .A1(n8403), .A2(n8402), .A3(n8401), .A4(n8400), .ZN(
        P2_U3257) );
  INV_X1 U9922 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8418) );
  NOR2_X1 U9923 ( .A1(n8405), .A2(n8404), .ZN(n8406) );
  XOR2_X1 U9924 ( .A(n8406), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8412) );
  NAND2_X1 U9925 ( .A1(n8408), .A2(n8407), .ZN(n8410) );
  INV_X1 U9926 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8409) );
  XNOR2_X1 U9927 ( .A(n8410), .B(n8409), .ZN(n8414) );
  INV_X1 U9928 ( .A(n8414), .ZN(n8411) );
  AOI22_X1 U9929 ( .A1(n8412), .A2(n9715), .B1(n8411), .B2(n9711), .ZN(n8415)
         );
  NOR2_X1 U9930 ( .A1(n8412), .A2(n9686), .ZN(n8413) );
  OAI211_X1 U9931 ( .C1(n8419), .C2(n8418), .A(n8417), .B(n8416), .ZN(P2_U3264) );
  NAND2_X1 U9932 ( .A1(n8719), .A2(n8428), .ZN(n8420) );
  NAND2_X1 U9933 ( .A1(n8636), .A2(n9761), .ZN(n8427) );
  INV_X1 U9934 ( .A(n8422), .ZN(n8424) );
  NOR2_X1 U9935 ( .A1(n8424), .A2(n8423), .ZN(n8639) );
  INV_X1 U9936 ( .A(n8639), .ZN(n8425) );
  NOR2_X1 U9937 ( .A1(n4392), .A2(n8425), .ZN(n8430) );
  AOI21_X1 U9938 ( .B1(n4392), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8430), .ZN(
        n8426) );
  OAI211_X1 U9939 ( .C1(n4714), .C2(n9757), .A(n8427), .B(n8426), .ZN(P2_U3265) );
  XNOR2_X1 U9940 ( .A(n8429), .B(n8428), .ZN(n8640) );
  NAND2_X1 U9941 ( .A1(n8640), .A2(n9761), .ZN(n8432) );
  AOI21_X1 U9942 ( .B1(n4392), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8430), .ZN(
        n8431) );
  OAI211_X1 U9943 ( .C1(n8719), .C2(n9757), .A(n8432), .B(n8431), .ZN(P2_U3266) );
  OAI21_X1 U9944 ( .B1(n8434), .B2(n8436), .A(n8433), .ZN(n8650) );
  INV_X1 U9945 ( .A(n8650), .ZN(n8449) );
  AOI211_X1 U9946 ( .C1(n8437), .C2(n8436), .A(n9740), .B(n8435), .ZN(n8440)
         );
  OAI22_X1 U9947 ( .A1(n8438), .A2(n9743), .B1(n8471), .B2(n9745), .ZN(n8439)
         );
  OR2_X1 U9948 ( .A1(n8440), .A2(n8439), .ZN(n8648) );
  INV_X1 U9949 ( .A(n8442), .ZN(n8724) );
  AOI211_X1 U9950 ( .C1(n8442), .C2(n8453), .A(n9838), .B(n8441), .ZN(n8649)
         );
  NAND2_X1 U9951 ( .A1(n8649), .A2(n9734), .ZN(n8446) );
  INV_X1 U9952 ( .A(n8443), .ZN(n8444) );
  AOI22_X1 U9953 ( .A1(n8444), .A2(n9776), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n4392), .ZN(n8445) );
  OAI211_X1 U9954 ( .C1(n8724), .C2(n9757), .A(n8446), .B(n8445), .ZN(n8447)
         );
  AOI21_X1 U9955 ( .B1(n8648), .B2(n9785), .A(n8447), .ZN(n8448) );
  OAI21_X1 U9956 ( .B1(n8449), .B2(n9755), .A(n8448), .ZN(P2_U3268) );
  OAI21_X1 U9957 ( .B1(n8451), .B2(n8458), .A(n8450), .ZN(n8452) );
  INV_X1 U9958 ( .A(n8452), .ZN(n8656) );
  INV_X1 U9959 ( .A(n8453), .ZN(n8454) );
  AOI21_X1 U9960 ( .B1(n8652), .B2(n8472), .A(n8454), .ZN(n8653) );
  AOI22_X1 U9961 ( .A1(n8455), .A2(n9776), .B1(n4392), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8456) );
  OAI21_X1 U9962 ( .B1(n4723), .B2(n9757), .A(n8456), .ZN(n8463) );
  NOR2_X1 U9963 ( .A1(n8467), .A2(n8457), .ZN(n8459) );
  NOR2_X1 U9964 ( .A1(n8655), .A2(n4392), .ZN(n8462) );
  AOI211_X1 U9965 ( .C1(n8653), .C2(n9761), .A(n8463), .B(n8462), .ZN(n8464)
         );
  OAI21_X1 U9966 ( .B1(n8656), .B2(n9755), .A(n8464), .ZN(P2_U3269) );
  OAI21_X1 U9967 ( .B1(n8466), .B2(n8469), .A(n8465), .ZN(n8659) );
  INV_X1 U9968 ( .A(n8659), .ZN(n8480) );
  OAI222_X1 U9969 ( .A1(n9743), .A2(n8471), .B1(n9745), .B2(n8501), .C1(n9740), 
        .C2(n8470), .ZN(n8657) );
  INV_X1 U9970 ( .A(n8472), .ZN(n8473) );
  AOI211_X1 U9971 ( .C1(n8477), .C2(n4727), .A(n9838), .B(n8473), .ZN(n8658)
         );
  INV_X1 U9972 ( .A(n8658), .ZN(n8475) );
  OAI22_X1 U9973 ( .A1(n8475), .A2(n4394), .B1(n9750), .B2(n8474), .ZN(n8476)
         );
  OAI21_X1 U9974 ( .B1(n8657), .B2(n8476), .A(n9785), .ZN(n8479) );
  AOI22_X1 U9975 ( .A1(n8477), .A2(n9726), .B1(n4392), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8478) );
  OAI211_X1 U9976 ( .C1(n8480), .C2(n9755), .A(n8479), .B(n8478), .ZN(P2_U3270) );
  OAI21_X1 U9977 ( .B1(n8482), .B2(n8484), .A(n8481), .ZN(n8483) );
  INV_X1 U9978 ( .A(n8483), .ZN(n8666) );
  XNOR2_X1 U9979 ( .A(n8485), .B(n8484), .ZN(n8486) );
  OAI222_X1 U9980 ( .A1(n9743), .A2(n8487), .B1(n9745), .B2(n8518), .C1(n9740), 
        .C2(n8486), .ZN(n8662) );
  AOI211_X1 U9981 ( .C1(n8664), .C2(n8502), .A(n9838), .B(n8488), .ZN(n8663)
         );
  INV_X1 U9982 ( .A(n8663), .ZN(n8491) );
  OAI22_X1 U9983 ( .A1(n8491), .A2(n4394), .B1(n9750), .B2(n8489), .ZN(n8492)
         );
  OAI21_X1 U9984 ( .B1(n8662), .B2(n8492), .A(n9785), .ZN(n8494) );
  AOI22_X1 U9985 ( .A1(n8664), .A2(n9726), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n4392), .ZN(n8493) );
  OAI211_X1 U9986 ( .C1(n8666), .C2(n9755), .A(n8494), .B(n8493), .ZN(P2_U3271) );
  XNOR2_X1 U9987 ( .A(n8495), .B(n8498), .ZN(n8670) );
  INV_X1 U9988 ( .A(n8670), .ZN(n8510) );
  NOR2_X1 U9989 ( .A1(n8496), .A2(n8497), .ZN(n8499) );
  XNOR2_X1 U9990 ( .A(n8499), .B(n8498), .ZN(n8500) );
  OAI222_X1 U9991 ( .A1(n9743), .A2(n8501), .B1(n9745), .B2(n8535), .C1(n8500), 
        .C2(n9740), .ZN(n8668) );
  OAI21_X1 U9992 ( .B1(n8734), .B2(n8519), .A(n8502), .ZN(n8667) );
  INV_X1 U9993 ( .A(n8503), .ZN(n8504) );
  AOI22_X1 U9994 ( .A1(n4392), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8504), .B2(
        n9776), .ZN(n8507) );
  NAND2_X1 U9995 ( .A1(n8505), .A2(n9726), .ZN(n8506) );
  OAI211_X1 U9996 ( .C1(n8667), .C2(n8562), .A(n8507), .B(n8506), .ZN(n8508)
         );
  AOI21_X1 U9997 ( .B1(n8668), .B2(n9785), .A(n8508), .ZN(n8509) );
  OAI21_X1 U9998 ( .B1(n9755), .B2(n8510), .A(n8509), .ZN(P2_U3272) );
  OAI21_X1 U9999 ( .B1(n8513), .B2(n8512), .A(n8511), .ZN(n8676) );
  INV_X1 U10000 ( .A(n8514), .ZN(n8532) );
  AOI21_X1 U10001 ( .B1(n8532), .B2(n8515), .A(n4942), .ZN(n8516) );
  NOR2_X1 U10002 ( .A1(n8496), .A2(n8516), .ZN(n8517) );
  OAI222_X1 U10003 ( .A1(n9745), .A2(n8551), .B1(n9743), .B2(n8518), .C1(n9740), .C2(n8517), .ZN(n8672) );
  INV_X1 U10004 ( .A(n8536), .ZN(n8520) );
  AOI211_X1 U10005 ( .C1(n8674), .C2(n8520), .A(n9838), .B(n8519), .ZN(n8673)
         );
  NAND2_X1 U10006 ( .A1(n8673), .A2(n9734), .ZN(n8524) );
  INV_X1 U10007 ( .A(n8521), .ZN(n8522) );
  AOI22_X1 U10008 ( .A1(n4392), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8522), .B2(
        n9776), .ZN(n8523) );
  OAI211_X1 U10009 ( .C1(n8525), .C2(n9757), .A(n8524), .B(n8523), .ZN(n8526)
         );
  AOI21_X1 U10010 ( .B1(n8672), .B2(n9785), .A(n8526), .ZN(n8527) );
  OAI21_X1 U10011 ( .B1(n9755), .B2(n8676), .A(n8527), .ZN(P2_U3273) );
  XOR2_X1 U10012 ( .A(n8529), .B(n8528), .Z(n8677) );
  OAI21_X1 U10013 ( .B1(n8550), .B2(n8530), .A(n8529), .ZN(n8531) );
  NAND3_X1 U10014 ( .A1(n8532), .A2(n9774), .A3(n8531), .ZN(n8534) );
  NAND2_X1 U10015 ( .A1(n8567), .A2(n9770), .ZN(n8533) );
  OAI211_X1 U10016 ( .C1(n8535), .C2(n9743), .A(n8534), .B(n8533), .ZN(n8679)
         );
  AOI21_X1 U10017 ( .B1(n8537), .B2(n8544), .A(n8536), .ZN(n8680) );
  NAND2_X1 U10018 ( .A1(n8680), .A2(n9761), .ZN(n8540) );
  AOI22_X1 U10019 ( .A1(n4392), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8538), .B2(
        n9776), .ZN(n8539) );
  OAI211_X1 U10020 ( .C1(n8739), .C2(n9757), .A(n8540), .B(n8539), .ZN(n8541)
         );
  AOI21_X1 U10021 ( .B1(n8679), .B2(n9785), .A(n8541), .ZN(n8542) );
  OAI21_X1 U10022 ( .B1(n8677), .B2(n9755), .A(n8542), .ZN(P2_U3274) );
  NAND2_X1 U10023 ( .A1(n8569), .A2(n8559), .ZN(n8543) );
  AND2_X1 U10024 ( .A1(n8544), .A2(n8543), .ZN(n8682) );
  INV_X1 U10025 ( .A(n8682), .ZN(n8563) );
  OAI22_X1 U10026 ( .A1(n8546), .A2(n9848), .B1(n8545), .B2(n9740), .ZN(n8549)
         );
  AND2_X1 U10027 ( .A1(n8546), .A2(n9859), .ZN(n8548) );
  MUX2_X1 U10028 ( .A(n8549), .B(n8548), .S(n8547), .Z(n8556) );
  NAND2_X1 U10029 ( .A1(n8550), .A2(n9774), .ZN(n8554) );
  OAI22_X1 U10030 ( .A1(n8551), .A2(n9743), .B1(n8592), .B2(n9745), .ZN(n8552)
         );
  INV_X1 U10031 ( .A(n8552), .ZN(n8553) );
  NAND2_X1 U10032 ( .A1(n8554), .A2(n8553), .ZN(n8555) );
  NOR2_X1 U10033 ( .A1(n8556), .A2(n8555), .ZN(n8684) );
  OAI21_X1 U10034 ( .B1(n8557), .B2(n9750), .A(n8684), .ZN(n8558) );
  NAND2_X1 U10035 ( .A1(n8558), .A2(n9785), .ZN(n8561) );
  AOI22_X1 U10036 ( .A1(n8559), .A2(n9726), .B1(n4392), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n8560) );
  OAI211_X1 U10037 ( .C1(n8563), .C2(n8562), .A(n8561), .B(n8560), .ZN(
        P2_U3275) );
  NAND2_X1 U10038 ( .A1(n8587), .A2(n8564), .ZN(n8565) );
  XNOR2_X1 U10039 ( .A(n8565), .B(n8571), .ZN(n8568) );
  AOI222_X1 U10040 ( .A1(n9774), .A2(n8568), .B1(n8567), .B2(n9771), .C1(n8566), .C2(n9770), .ZN(n8693) );
  OAI211_X1 U10041 ( .C1(n8584), .C2(n8570), .A(n9845), .B(n8569), .ZN(n8692)
         );
  NAND2_X1 U10042 ( .A1(n8572), .A2(n8571), .ZN(n8687) );
  NAND3_X1 U10043 ( .A1(n8688), .A2(n8687), .A3(n9782), .ZN(n8577) );
  INV_X1 U10044 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8574) );
  OAI22_X1 U10045 ( .A1(n9785), .A2(n8574), .B1(n8573), .B2(n9750), .ZN(n8575)
         );
  AOI21_X1 U10046 ( .B1(n8689), .B2(n9726), .A(n8575), .ZN(n8576) );
  OAI211_X1 U10047 ( .C1(n8692), .C2(n8578), .A(n8577), .B(n8576), .ZN(n8579)
         );
  INV_X1 U10048 ( .A(n8579), .ZN(n8580) );
  OAI21_X1 U10049 ( .B1(n8693), .B2(n4392), .A(n8580), .ZN(P2_U3276) );
  XNOR2_X1 U10050 ( .A(n8581), .B(n8589), .ZN(n8698) );
  INV_X1 U10051 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8583) );
  OAI22_X1 U10052 ( .A1(n9785), .A2(n8583), .B1(n8582), .B2(n9750), .ZN(n8595)
         );
  INV_X1 U10053 ( .A(n8603), .ZN(n8585) );
  AOI211_X1 U10054 ( .C1(n8696), .C2(n8585), .A(n9838), .B(n8584), .ZN(n8695)
         );
  INV_X1 U10055 ( .A(n8587), .ZN(n8588) );
  AOI21_X1 U10056 ( .B1(n8586), .B2(n8589), .A(n8588), .ZN(n8590) );
  OAI222_X1 U10057 ( .A1(n9743), .A2(n8592), .B1(n9745), .B2(n8591), .C1(n9740), .C2(n8590), .ZN(n8694) );
  AOI21_X1 U10058 ( .B1(n8695), .B2(n4504), .A(n8694), .ZN(n8593) );
  NOR2_X1 U10059 ( .A1(n8593), .A2(n4392), .ZN(n8594) );
  AOI211_X1 U10060 ( .C1(n9726), .C2(n8696), .A(n8595), .B(n8594), .ZN(n8596)
         );
  OAI21_X1 U10061 ( .B1(n9755), .B2(n8698), .A(n8596), .ZN(P2_U3277) );
  XOR2_X1 U10062 ( .A(n8599), .B(n8597), .Z(n8701) );
  INV_X1 U10063 ( .A(n8701), .ZN(n8610) );
  XNOR2_X1 U10064 ( .A(n8598), .B(n8599), .ZN(n8600) );
  OAI222_X1 U10065 ( .A1(n9743), .A2(n8602), .B1(n9745), .B2(n8601), .C1(n9740), .C2(n8600), .ZN(n8699) );
  AOI211_X1 U10066 ( .C1(n8604), .C2(n8611), .A(n9838), .B(n8603), .ZN(n8700)
         );
  NAND2_X1 U10067 ( .A1(n8700), .A2(n9734), .ZN(n8607) );
  AOI22_X1 U10068 ( .A1(n4392), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8605), .B2(
        n9776), .ZN(n8606) );
  OAI211_X1 U10069 ( .C1(n8749), .C2(n9757), .A(n8607), .B(n8606), .ZN(n8608)
         );
  AOI21_X1 U10070 ( .B1(n8699), .B2(n9785), .A(n8608), .ZN(n8609) );
  OAI21_X1 U10071 ( .B1(n8610), .B2(n9755), .A(n8609), .ZN(P2_U3278) );
  INV_X1 U10072 ( .A(n8611), .ZN(n8612) );
  AOI211_X1 U10073 ( .C1(n8706), .C2(n8613), .A(n9838), .B(n8612), .ZN(n8705)
         );
  NAND2_X1 U10074 ( .A1(n8614), .A2(n8618), .ZN(n8615) );
  AOI21_X1 U10075 ( .B1(n8616), .B2(n8615), .A(n9848), .ZN(n8704) );
  XOR2_X1 U10076 ( .A(n8617), .B(n8618), .Z(n8621) );
  AOI222_X1 U10077 ( .A1(n9774), .A2(n8621), .B1(n8620), .B2(n9771), .C1(n8619), .C2(n9770), .ZN(n8707) );
  INV_X1 U10078 ( .A(n8707), .ZN(n8622) );
  AOI211_X1 U10079 ( .C1(n8705), .C2(n4504), .A(n8704), .B(n8622), .ZN(n8626)
         );
  AOI22_X1 U10080 ( .A1(n4392), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8623), .B2(
        n9776), .ZN(n8625) );
  NAND2_X1 U10081 ( .A1(n8706), .A2(n9726), .ZN(n8624) );
  OAI211_X1 U10082 ( .C1(n8626), .C2(n4392), .A(n8625), .B(n8624), .ZN(
        P2_U3279) );
  MUX2_X1 U10083 ( .A(n6446), .B(n8627), .S(n9785), .Z(n8635) );
  AOI22_X1 U10084 ( .A1(n9761), .A2(n8629), .B1(n8628), .B2(n9776), .ZN(n8634)
         );
  OR2_X1 U10085 ( .A1(n8630), .A2(n9755), .ZN(n8633) );
  OR2_X1 U10086 ( .A1(n9757), .A2(n8631), .ZN(n8632) );
  NAND4_X1 U10087 ( .A1(n8635), .A2(n8634), .A3(n8633), .A4(n8632), .ZN(
        P2_U3290) );
  INV_X1 U10088 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8637) );
  MUX2_X1 U10089 ( .A(n8637), .B(n8714), .S(n9879), .Z(n8638) );
  OAI21_X1 U10090 ( .B1(n4714), .B2(n8713), .A(n8638), .ZN(P2_U3551) );
  AOI21_X1 U10091 ( .B1(n8640), .B2(n9845), .A(n8639), .ZN(n8716) );
  MUX2_X1 U10092 ( .A(n8641), .B(n8716), .S(n9879), .Z(n8642) );
  OAI21_X1 U10093 ( .B1(n8719), .B2(n8713), .A(n8642), .ZN(P2_U3550) );
  AOI22_X1 U10094 ( .A1(n8644), .A2(n9845), .B1(n9844), .B2(n8643), .ZN(n8645)
         );
  OAI211_X1 U10095 ( .C1(n8647), .C2(n9848), .A(n8646), .B(n8645), .ZN(n8720)
         );
  MUX2_X1 U10096 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8720), .S(n9879), .Z(
        P2_U3549) );
  AOI211_X1 U10097 ( .C1(n9859), .C2(n8650), .A(n8649), .B(n8648), .ZN(n8721)
         );
  MUX2_X1 U10098 ( .A(n10132), .B(n8721), .S(n9879), .Z(n8651) );
  OAI21_X1 U10099 ( .B1(n8724), .B2(n8713), .A(n8651), .ZN(P2_U3548) );
  AOI22_X1 U10100 ( .A1(n8653), .A2(n9845), .B1(n9844), .B2(n8652), .ZN(n8654)
         );
  OAI211_X1 U10101 ( .C1(n8656), .C2(n9848), .A(n8655), .B(n8654), .ZN(n8725)
         );
  MUX2_X1 U10102 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8725), .S(n9879), .Z(
        P2_U3547) );
  AOI211_X1 U10103 ( .C1(n9859), .C2(n8659), .A(n8658), .B(n8657), .ZN(n8726)
         );
  MUX2_X1 U10104 ( .A(n8660), .B(n8726), .S(n9879), .Z(n8661) );
  OAI21_X1 U10105 ( .B1(n8729), .B2(n8713), .A(n8661), .ZN(P2_U3546) );
  AOI211_X1 U10106 ( .C1(n9844), .C2(n8664), .A(n8663), .B(n8662), .ZN(n8665)
         );
  OAI21_X1 U10107 ( .B1(n8666), .B2(n9848), .A(n8665), .ZN(n8730) );
  MUX2_X1 U10108 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8730), .S(n9879), .Z(
        P2_U3545) );
  NOR2_X1 U10109 ( .A1(n8667), .A2(n9838), .ZN(n8669) );
  AOI211_X1 U10110 ( .C1(n8670), .C2(n9859), .A(n8669), .B(n8668), .ZN(n8731)
         );
  MUX2_X1 U10111 ( .A(n10180), .B(n8731), .S(n9879), .Z(n8671) );
  OAI21_X1 U10112 ( .B1(n8734), .B2(n8713), .A(n8671), .ZN(P2_U3544) );
  AOI211_X1 U10113 ( .C1(n9844), .C2(n8674), .A(n8673), .B(n8672), .ZN(n8675)
         );
  OAI21_X1 U10114 ( .B1(n9848), .B2(n8676), .A(n8675), .ZN(n8735) );
  MUX2_X1 U10115 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8735), .S(n9879), .Z(
        P2_U3543) );
  NOR2_X1 U10116 ( .A1(n8677), .A2(n9848), .ZN(n8678) );
  AOI211_X1 U10117 ( .C1(n9845), .C2(n8680), .A(n8679), .B(n8678), .ZN(n8736)
         );
  MUX2_X1 U10118 ( .A(n9913), .B(n8736), .S(n9879), .Z(n8681) );
  OAI21_X1 U10119 ( .B1(n8739), .B2(n8713), .A(n8681), .ZN(P2_U3542) );
  NAND2_X1 U10120 ( .A1(n8682), .A2(n9845), .ZN(n8683) );
  NAND2_X1 U10121 ( .A1(n8684), .A2(n8683), .ZN(n8740) );
  MUX2_X1 U10122 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8740), .S(n9879), .Z(n8685) );
  INV_X1 U10123 ( .A(n8685), .ZN(n8686) );
  OAI21_X1 U10124 ( .B1(n8743), .B2(n8713), .A(n8686), .ZN(P2_U3541) );
  NAND3_X1 U10125 ( .A1(n8688), .A2(n9859), .A3(n8687), .ZN(n8691) );
  NAND2_X1 U10126 ( .A1(n8689), .A2(n9844), .ZN(n8690) );
  NAND4_X1 U10127 ( .A1(n8693), .A2(n8692), .A3(n8691), .A4(n8690), .ZN(n8744)
         );
  MUX2_X1 U10128 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8744), .S(n9879), .Z(
        P2_U3540) );
  AOI211_X1 U10129 ( .C1(n9844), .C2(n8696), .A(n8695), .B(n8694), .ZN(n8697)
         );
  OAI21_X1 U10130 ( .B1(n9848), .B2(n8698), .A(n8697), .ZN(n8745) );
  MUX2_X1 U10131 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8745), .S(n9879), .Z(
        P2_U3539) );
  INV_X1 U10132 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8702) );
  AOI211_X1 U10133 ( .C1(n9859), .C2(n8701), .A(n8700), .B(n8699), .ZN(n8746)
         );
  MUX2_X1 U10134 ( .A(n8702), .B(n8746), .S(n9879), .Z(n8703) );
  OAI21_X1 U10135 ( .B1(n8749), .B2(n8713), .A(n8703), .ZN(P2_U3538) );
  AOI211_X1 U10136 ( .C1(n9844), .C2(n8706), .A(n8705), .B(n8704), .ZN(n8708)
         );
  NAND2_X1 U10137 ( .A1(n8708), .A2(n8707), .ZN(n8750) );
  MUX2_X1 U10138 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8750), .S(n9879), .Z(
        P2_U3537) );
  AOI21_X1 U10139 ( .B1(n9845), .B2(n8710), .A(n8709), .ZN(n8751) );
  MUX2_X1 U10140 ( .A(n8711), .B(n8751), .S(n9879), .Z(n8712) );
  OAI21_X1 U10141 ( .B1(n8755), .B2(n8713), .A(n8712), .ZN(P2_U3536) );
  INV_X1 U10142 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8715) );
  INV_X1 U10143 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8717) );
  MUX2_X1 U10144 ( .A(n8717), .B(n8716), .S(n9861), .Z(n8718) );
  OAI21_X1 U10145 ( .B1(n8719), .B2(n8754), .A(n8718), .ZN(P2_U3518) );
  MUX2_X1 U10146 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8720), .S(n9861), .Z(
        P2_U3517) );
  INV_X1 U10147 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8722) );
  MUX2_X1 U10148 ( .A(n8722), .B(n8721), .S(n9861), .Z(n8723) );
  OAI21_X1 U10149 ( .B1(n8724), .B2(n8754), .A(n8723), .ZN(P2_U3516) );
  MUX2_X1 U10150 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8725), .S(n9861), .Z(
        P2_U3515) );
  INV_X1 U10151 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8727) );
  MUX2_X1 U10152 ( .A(n8727), .B(n8726), .S(n9861), .Z(n8728) );
  OAI21_X1 U10153 ( .B1(n8729), .B2(n8754), .A(n8728), .ZN(P2_U3514) );
  MUX2_X1 U10154 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8730), .S(n9861), .Z(
        P2_U3513) );
  INV_X1 U10155 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8732) );
  MUX2_X1 U10156 ( .A(n8732), .B(n8731), .S(n9861), .Z(n8733) );
  OAI21_X1 U10157 ( .B1(n8734), .B2(n8754), .A(n8733), .ZN(P2_U3512) );
  MUX2_X1 U10158 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8735), .S(n9861), .Z(
        P2_U3511) );
  INV_X1 U10159 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8737) );
  MUX2_X1 U10160 ( .A(n8737), .B(n8736), .S(n9861), .Z(n8738) );
  OAI21_X1 U10161 ( .B1(n8739), .B2(n8754), .A(n8738), .ZN(P2_U3510) );
  MUX2_X1 U10162 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8740), .S(n9861), .Z(n8741) );
  INV_X1 U10163 ( .A(n8741), .ZN(n8742) );
  OAI21_X1 U10164 ( .B1(n8743), .B2(n8754), .A(n8742), .ZN(P2_U3509) );
  MUX2_X1 U10165 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8744), .S(n9861), .Z(
        P2_U3508) );
  MUX2_X1 U10166 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8745), .S(n9861), .Z(
        P2_U3507) );
  INV_X1 U10167 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8747) );
  MUX2_X1 U10168 ( .A(n8747), .B(n8746), .S(n9861), .Z(n8748) );
  OAI21_X1 U10169 ( .B1(n8749), .B2(n8754), .A(n8748), .ZN(P2_U3505) );
  MUX2_X1 U10170 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8750), .S(n9861), .Z(
        P2_U3502) );
  INV_X1 U10171 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8752) );
  MUX2_X1 U10172 ( .A(n8752), .B(n8751), .S(n9861), .Z(n8753) );
  OAI21_X1 U10173 ( .B1(n8755), .B2(n8754), .A(n8753), .ZN(P2_U3499) );
  INV_X1 U10174 ( .A(n8032), .ZN(n9467) );
  NOR4_X1 U10175 ( .A1(n8756), .A2(P2_IR_REG_30__SCAN_IN), .A3(n5795), .A4(
        P2_U3152), .ZN(n8757) );
  AOI21_X1 U10176 ( .B1(n8758), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8757), .ZN(
        n8759) );
  OAI21_X1 U10177 ( .B1(n9467), .B2(n8769), .A(n8759), .ZN(P2_U3327) );
  INV_X1 U10178 ( .A(n8760), .ZN(n9472) );
  OAI222_X1 U10179 ( .A1(n8762), .A2(P2_U3152), .B1(n8769), .B2(n9472), .C1(
        n8761), .C2(n8771), .ZN(P2_U3329) );
  INV_X1 U10180 ( .A(n9475), .ZN(n8764) );
  OAI222_X1 U10181 ( .A1(n8765), .A2(P2_U3152), .B1(n8769), .B2(n8764), .C1(
        n8763), .C2(n8771), .ZN(P2_U3330) );
  INV_X1 U10182 ( .A(n8766), .ZN(n8768) );
  OAI222_X1 U10183 ( .A1(n8771), .A2(n8770), .B1(n8769), .B2(n8768), .C1(n8767), .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U10184 ( .A(n8772), .ZN(n8773) );
  MUX2_X1 U10185 ( .A(n8773), .B(n9691), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10186 ( .A(n8774), .ZN(n8778) );
  AOI21_X1 U10187 ( .B1(n8943), .B2(n8776), .A(n8775), .ZN(n8777) );
  AOI22_X1 U10188 ( .A1(n8921), .A2(n9132), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8779) );
  OAI21_X1 U10189 ( .B1(n8965), .B2(n9162), .A(n8779), .ZN(n8780) );
  AOI21_X1 U10190 ( .B1(n8962), .B2(n9201), .A(n8780), .ZN(n8781) );
  OAI211_X1 U10191 ( .C1(n9165), .C2(n8954), .A(n8782), .B(n8781), .ZN(
        P1_U3212) );
  NAND2_X1 U10192 ( .A1(n8784), .A2(n8783), .ZN(n8785) );
  XOR2_X1 U10193 ( .A(n8786), .B(n8785), .Z(n8795) );
  OAI21_X1 U10194 ( .B1(n8948), .B2(n8788), .A(n8787), .ZN(n8789) );
  AOI21_X1 U10195 ( .B1(n8921), .B2(n10214), .A(n8789), .ZN(n8790) );
  OAI21_X1 U10196 ( .B1(n8965), .B2(n8791), .A(n8790), .ZN(n8792) );
  AOI21_X1 U10197 ( .B1(n8793), .B2(n8967), .A(n8792), .ZN(n8794) );
  OAI21_X1 U10198 ( .B1(n8795), .B2(n8969), .A(n8794), .ZN(P1_U3213) );
  NAND2_X1 U10199 ( .A1(n8868), .A2(n8796), .ZN(n8797) );
  XOR2_X1 U10200 ( .A(n8798), .B(n8797), .Z(n8803) );
  AOI22_X1 U10201 ( .A1(n8962), .A2(n9228), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8800) );
  NAND2_X1 U10202 ( .A1(n8921), .A2(n9229), .ZN(n8799) );
  OAI211_X1 U10203 ( .C1(n8965), .C2(n9222), .A(n8800), .B(n8799), .ZN(n8801)
         );
  AOI21_X1 U10204 ( .B1(n9392), .B2(n8967), .A(n8801), .ZN(n8802) );
  OAI21_X1 U10205 ( .B1(n8803), .B2(n8969), .A(n8802), .ZN(P1_U3214) );
  AND2_X1 U10206 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3084), .ZN(n9596) );
  AOI21_X1 U10207 ( .B1(n8962), .B2(n8977), .A(n9596), .ZN(n8805) );
  NAND2_X1 U10208 ( .A1(n8921), .A2(n8975), .ZN(n8804) );
  OAI211_X1 U10209 ( .C1(n8965), .C2(n9497), .A(n8805), .B(n8804), .ZN(n8812)
         );
  XNOR2_X1 U10210 ( .A(n8807), .B(n8806), .ZN(n8808) );
  XNOR2_X1 U10211 ( .A(n8809), .B(n8808), .ZN(n8810) );
  NOR2_X1 U10212 ( .A1(n8810), .A2(n8969), .ZN(n8811) );
  AOI211_X1 U10213 ( .C1(n9501), .C2(n8967), .A(n8812), .B(n8811), .ZN(n8813)
         );
  INV_X1 U10214 ( .A(n8813), .ZN(P1_U3215) );
  XOR2_X1 U10215 ( .A(n8815), .B(n8814), .Z(n8820) );
  NAND2_X1 U10216 ( .A1(n8951), .A2(n9282), .ZN(n8817) );
  INV_X1 U10217 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10171) );
  NOR2_X1 U10218 ( .A1(n10171), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9070) );
  AOI21_X1 U10219 ( .B1(n8921), .B2(n9289), .A(n9070), .ZN(n8816) );
  OAI211_X1 U10220 ( .C1(n9328), .C2(n8948), .A(n8817), .B(n8816), .ZN(n8818)
         );
  AOI21_X1 U10221 ( .B1(n9415), .B2(n8967), .A(n8818), .ZN(n8819) );
  OAI21_X1 U10222 ( .B1(n8820), .B2(n8969), .A(n8819), .ZN(P1_U3217) );
  XOR2_X1 U10223 ( .A(n8822), .B(n8821), .Z(n8828) );
  OAI22_X1 U10224 ( .A1(n8960), .A2(n9255), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8823), .ZN(n8824) );
  AOI21_X1 U10225 ( .B1(n8962), .B2(n9289), .A(n8824), .ZN(n8825) );
  OAI21_X1 U10226 ( .B1(n8965), .B2(n9249), .A(n8825), .ZN(n8826) );
  AOI21_X1 U10227 ( .B1(n9405), .B2(n8967), .A(n8826), .ZN(n8827) );
  OAI21_X1 U10228 ( .B1(n8828), .B2(n8969), .A(n8827), .ZN(P1_U3221) );
  INV_X1 U10229 ( .A(n8829), .ZN(n8830) );
  AOI21_X1 U10230 ( .B1(n8832), .B2(n8831), .A(n8830), .ZN(n8839) );
  OAI22_X1 U10231 ( .A1(n8948), .A2(n9493), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5298), .ZN(n8833) );
  AOI21_X1 U10232 ( .B1(n8921), .B2(n8973), .A(n8833), .ZN(n8834) );
  OAI21_X1 U10233 ( .B1(n8965), .B2(n8835), .A(n8834), .ZN(n8836) );
  AOI21_X1 U10234 ( .B1(n8837), .B2(n8967), .A(n8836), .ZN(n8838) );
  OAI21_X1 U10235 ( .B1(n8839), .B2(n8969), .A(n8838), .ZN(P1_U3222) );
  OAI21_X1 U10236 ( .B1(n8842), .B2(n8841), .A(n8840), .ZN(n8843) );
  NAND2_X1 U10237 ( .A1(n8843), .A2(n8944), .ZN(n8847) );
  AOI22_X1 U10238 ( .A1(n8962), .A2(n9229), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8844) );
  OAI21_X1 U10239 ( .B1(n8965), .B2(n9195), .A(n8844), .ZN(n8845) );
  AOI21_X1 U10240 ( .B1(n8921), .B2(n9201), .A(n8845), .ZN(n8846) );
  OAI211_X1 U10241 ( .C1(n9198), .C2(n8954), .A(n8847), .B(n8846), .ZN(
        P1_U3223) );
  INV_X1 U10242 ( .A(n8849), .ZN(n8851) );
  NOR2_X1 U10243 ( .A1(n8851), .A2(n8850), .ZN(n8852) );
  XNOR2_X1 U10244 ( .A(n8848), .B(n8852), .ZN(n8857) );
  NAND2_X1 U10245 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n9023) );
  OAI21_X1 U10246 ( .B1(n8948), .B2(n9348), .A(n9023), .ZN(n8853) );
  AOI21_X1 U10247 ( .B1(n8921), .B2(n9304), .A(n8853), .ZN(n8854) );
  OAI21_X1 U10248 ( .B1(n8965), .B2(n9340), .A(n8854), .ZN(n8855) );
  AOI21_X1 U10249 ( .B1(n9431), .B2(n8967), .A(n8855), .ZN(n8856) );
  OAI21_X1 U10250 ( .B1(n8857), .B2(n8969), .A(n8856), .ZN(P1_U3224) );
  XOR2_X1 U10251 ( .A(n8859), .B(n8858), .Z(n8864) );
  NAND2_X1 U10252 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9037) );
  OAI21_X1 U10253 ( .B1(n8960), .B2(n9328), .A(n9037), .ZN(n8860) );
  AOI21_X1 U10254 ( .B1(n8962), .B2(n9087), .A(n8860), .ZN(n8861) );
  OAI21_X1 U10255 ( .B1(n8965), .B2(n9320), .A(n8861), .ZN(n8862) );
  AOI21_X1 U10256 ( .B1(n9426), .B2(n8967), .A(n8862), .ZN(n8863) );
  OAI21_X1 U10257 ( .B1(n8864), .B2(n8969), .A(n8863), .ZN(P1_U3226) );
  INV_X1 U10258 ( .A(n8865), .ZN(n8870) );
  AOI21_X1 U10259 ( .B1(n8868), .B2(n8867), .A(n8866), .ZN(n8869) );
  OAI21_X1 U10260 ( .B1(n8870), .B2(n8869), .A(n8944), .ZN(n8875) );
  OAI22_X1 U10261 ( .A1(n8948), .A2(n9238), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8871), .ZN(n8873) );
  NOR2_X1 U10262 ( .A1(n9210), .A2(n8960), .ZN(n8872) );
  AOI211_X1 U10263 ( .C1(n9212), .C2(n8951), .A(n8873), .B(n8872), .ZN(n8874)
         );
  OAI211_X1 U10264 ( .C1(n9096), .C2(n8954), .A(n8875), .B(n8874), .ZN(
        P1_U3227) );
  OAI21_X1 U10265 ( .B1(n8878), .B2(n8877), .A(n8876), .ZN(n8879) );
  NAND2_X1 U10266 ( .A1(n8879), .A2(n8944), .ZN(n8887) );
  AOI21_X1 U10267 ( .B1(n8962), .B2(n8978), .A(n8880), .ZN(n8882) );
  NAND2_X1 U10268 ( .A1(n8921), .A2(n8976), .ZN(n8881) );
  OAI211_X1 U10269 ( .C1(n8965), .C2(n8883), .A(n8882), .B(n8881), .ZN(n8884)
         );
  AOI21_X1 U10270 ( .B1(n8885), .B2(n8967), .A(n8884), .ZN(n8886) );
  NAND2_X1 U10271 ( .A1(n8887), .A2(n8886), .ZN(P1_U3229) );
  INV_X1 U10272 ( .A(n8888), .ZN(n8889) );
  NOR2_X1 U10273 ( .A1(n8890), .A2(n8889), .ZN(n8891) );
  XNOR2_X1 U10274 ( .A(n8892), .B(n8891), .ZN(n8897) );
  OAI22_X1 U10275 ( .A1(n8960), .A2(n9275), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9992), .ZN(n8893) );
  AOI21_X1 U10276 ( .B1(n8962), .B2(n9306), .A(n8893), .ZN(n8894) );
  OAI21_X1 U10277 ( .B1(n8965), .B2(n9268), .A(n8894), .ZN(n8895) );
  AOI21_X1 U10278 ( .B1(n9411), .B2(n8967), .A(n8895), .ZN(n8896) );
  OAI21_X1 U10279 ( .B1(n8897), .B2(n8969), .A(n8896), .ZN(P1_U3231) );
  INV_X1 U10280 ( .A(n8899), .ZN(n8903) );
  OAI21_X1 U10281 ( .B1(n8901), .B2(n8903), .A(n8900), .ZN(n8902) );
  OAI211_X1 U10282 ( .C1(n8904), .C2(n8903), .A(n8944), .B(n8902), .ZN(n8911)
         );
  OAI21_X1 U10283 ( .B1(n8948), .B2(n8906), .A(n8905), .ZN(n8909) );
  NOR2_X1 U10284 ( .A1(n8965), .A2(n8907), .ZN(n8908) );
  AOI211_X1 U10285 ( .C1(n8921), .C2(n8972), .A(n8909), .B(n8908), .ZN(n8910)
         );
  OAI211_X1 U10286 ( .C1(n4698), .C2(n8954), .A(n8911), .B(n8910), .ZN(
        P1_U3232) );
  NAND2_X1 U10287 ( .A1(n4429), .A2(n8912), .ZN(n8914) );
  XNOR2_X1 U10288 ( .A(n8914), .B(n8913), .ZN(n8919) );
  AOI22_X1 U10289 ( .A1(n8962), .A2(n9092), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8916) );
  NAND2_X1 U10290 ( .A1(n8921), .A2(n8971), .ZN(n8915) );
  OAI211_X1 U10291 ( .C1(n8965), .C2(n9240), .A(n8916), .B(n8915), .ZN(n8917)
         );
  AOI21_X1 U10292 ( .B1(n9399), .B2(n8967), .A(n8917), .ZN(n8918) );
  OAI21_X1 U10293 ( .B1(n8919), .B2(n8969), .A(n8918), .ZN(P1_U3233) );
  INV_X1 U10294 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n8920) );
  NOR2_X1 U10295 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8920), .ZN(n9002) );
  AOI21_X1 U10296 ( .B1(n8962), .B2(n8976), .A(n9002), .ZN(n8923) );
  NAND2_X1 U10297 ( .A1(n8921), .A2(n8974), .ZN(n8922) );
  OAI211_X1 U10298 ( .C1(n8965), .C2(n8924), .A(n8923), .B(n8922), .ZN(n8929)
         );
  XNOR2_X1 U10299 ( .A(n8926), .B(n8925), .ZN(n8927) );
  NOR2_X1 U10300 ( .A1(n8927), .A2(n8969), .ZN(n8928) );
  AOI211_X1 U10301 ( .C1(n8930), .C2(n8967), .A(n8929), .B(n8928), .ZN(n8931)
         );
  INV_X1 U10302 ( .A(n8931), .ZN(P1_U3234) );
  INV_X1 U10303 ( .A(n9419), .ZN(n9298) );
  INV_X1 U10304 ( .A(n8932), .ZN(n8937) );
  OAI21_X1 U10305 ( .B1(n8934), .B2(n8936), .A(n8933), .ZN(n8935) );
  OAI211_X1 U10306 ( .C1(n8937), .C2(n8936), .A(n8944), .B(n8935), .ZN(n8941)
         );
  NAND2_X1 U10307 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9047) );
  NAND2_X1 U10308 ( .A1(n8962), .A2(n9304), .ZN(n8938) );
  OAI211_X1 U10309 ( .C1(n8960), .C2(n9276), .A(n9047), .B(n8938), .ZN(n8939)
         );
  AOI21_X1 U10310 ( .B1(n9309), .B2(n8951), .A(n8939), .ZN(n8940) );
  OAI211_X1 U10311 ( .C1(n9298), .C2(n8954), .A(n8941), .B(n8940), .ZN(
        P1_U3236) );
  INV_X1 U10312 ( .A(n9377), .ZN(n9179) );
  AND2_X1 U10313 ( .A1(n8840), .A2(n8942), .ZN(n8946) );
  OAI211_X1 U10314 ( .C1(n8946), .C2(n8945), .A(n8944), .B(n8943), .ZN(n8953)
         );
  OAI22_X1 U10315 ( .A1(n8960), .A2(n9103), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8947), .ZN(n8950) );
  NOR2_X1 U10316 ( .A1(n9210), .A2(n8948), .ZN(n8949) );
  AOI211_X1 U10317 ( .C1(n9177), .C2(n8951), .A(n8950), .B(n8949), .ZN(n8952)
         );
  OAI211_X1 U10318 ( .C1(n9179), .C2(n8954), .A(n8953), .B(n8952), .ZN(
        P1_U3238) );
  XNOR2_X1 U10319 ( .A(n8956), .B(n8955), .ZN(n8957) );
  XNOR2_X1 U10320 ( .A(n8958), .B(n8957), .ZN(n8970) );
  OAI21_X1 U10321 ( .B1(n8960), .B2(n9327), .A(n8959), .ZN(n8961) );
  AOI21_X1 U10322 ( .B1(n8962), .B2(n8972), .A(n8961), .ZN(n8963) );
  OAI21_X1 U10323 ( .B1(n8965), .B2(n8964), .A(n8963), .ZN(n8966) );
  AOI21_X1 U10324 ( .B1(n9084), .B2(n8967), .A(n8966), .ZN(n8968) );
  OAI21_X1 U10325 ( .B1(n8970), .B2(n8969), .A(n8968), .ZN(P1_U3239) );
  MUX2_X1 U10326 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9133), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10327 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9155), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10328 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9132), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10329 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9186), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10330 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9201), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10331 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9185), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10332 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9229), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10333 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n8971), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10334 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9228), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10335 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9092), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10336 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9289), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10337 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9306), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10338 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9288), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10339 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9304), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10340 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9087), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10341 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8972), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10342 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8973), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10343 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8974), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10344 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8975), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10345 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8976), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10346 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8977), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10347 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8978), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10348 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8979), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10349 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8980), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10350 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8981), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10351 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8982), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10352 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8983), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10353 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8984), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10354 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n8985), .S(P1_U4006), .Z(
        P1_U3556) );
  NAND2_X1 U10355 ( .A1(n9022), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n8995) );
  OR3_X1 U10356 ( .A1(n9558), .A2(n8986), .A3(P1_REG1_REG_0__SCAN_IN), .ZN(
        n8994) );
  XNOR2_X1 U10357 ( .A(n8987), .B(n8986), .ZN(n8990) );
  AOI21_X1 U10358 ( .B1(n5766), .B2(n8988), .A(P1_U3084), .ZN(n8989) );
  NAND4_X1 U10359 ( .A1(n8991), .A2(n8990), .A3(n8989), .A4(n5408), .ZN(n8993)
         );
  NAND2_X1 U10360 ( .A1(P1_U3084), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n8992) );
  NAND4_X1 U10361 ( .A1(n8995), .A2(n8994), .A3(n8993), .A4(n8992), .ZN(
        P1_U3241) );
  OAI21_X1 U10362 ( .B1(n8998), .B2(n8997), .A(n8996), .ZN(n8999) );
  NAND2_X1 U10363 ( .A1(n8999), .A2(n9575), .ZN(n9009) );
  NOR2_X1 U10364 ( .A1(n9583), .A2(n9000), .ZN(n9001) );
  AOI211_X1 U10365 ( .C1(n9022), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9002), .B(
        n9001), .ZN(n9008) );
  OAI21_X1 U10366 ( .B1(n9005), .B2(n9004), .A(n9003), .ZN(n9006) );
  NAND2_X1 U10367 ( .A1(n9006), .A2(n9597), .ZN(n9007) );
  NAND3_X1 U10368 ( .A1(n9009), .A2(n9008), .A3(n9007), .ZN(P1_U3252) );
  NOR2_X1 U10369 ( .A1(n9010), .A2(n9017), .ZN(n9012) );
  NAND2_X1 U10370 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9034), .ZN(n9013) );
  OAI21_X1 U10371 ( .B1(n9034), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9013), .ZN(
        n9014) );
  AOI211_X1 U10372 ( .C1(n9015), .C2(n9014), .A(n9029), .B(n9591), .ZN(n9028)
         );
  NOR2_X1 U10373 ( .A1(n9017), .A2(n9016), .ZN(n9019) );
  NOR2_X1 U10374 ( .A1(n9019), .A2(n9018), .ZN(n9021) );
  XNOR2_X1 U10375 ( .A(n9034), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9020) );
  NOR2_X1 U10376 ( .A1(n9021), .A2(n9020), .ZN(n9033) );
  AOI211_X1 U10377 ( .C1(n9021), .C2(n9020), .A(n9033), .B(n9558), .ZN(n9027)
         );
  NAND2_X1 U10378 ( .A1(n9022), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9024) );
  OAI211_X1 U10379 ( .C1(n9025), .C2(n9583), .A(n9024), .B(n9023), .ZN(n9026)
         );
  OR3_X1 U10380 ( .A1(n9028), .A2(n9027), .A3(n9026), .ZN(P1_U3257) );
  INV_X1 U10381 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U10382 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9050), .ZN(n9030) );
  OAI21_X1 U10383 ( .B1(n9050), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9030), .ZN(
        n9031) );
  AOI211_X1 U10384 ( .C1(n9032), .C2(n9031), .A(n9049), .B(n9591), .ZN(n9041)
         );
  XNOR2_X1 U10385 ( .A(n9050), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9035) );
  NOR2_X1 U10386 ( .A1(n9036), .A2(n9035), .ZN(n9044) );
  AOI211_X1 U10387 ( .C1(n9036), .C2(n9035), .A(n9044), .B(n9558), .ZN(n9040)
         );
  INV_X1 U10388 ( .A(n9050), .ZN(n9038) );
  OAI21_X1 U10389 ( .B1(n9583), .B2(n9038), .A(n9037), .ZN(n9039) );
  NOR3_X1 U10390 ( .A1(n9041), .A2(n9040), .A3(n9039), .ZN(n9042) );
  OAI21_X1 U10391 ( .B1(n9586), .B2(n9043), .A(n9042), .ZN(P1_U3258) );
  INV_X1 U10392 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9058) );
  XOR2_X1 U10393 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9062), .Z(n9046) );
  NAND2_X1 U10394 ( .A1(n9046), .A2(n9045), .ZN(n9061) );
  OAI21_X1 U10395 ( .B1(n9046), .B2(n9045), .A(n9061), .ZN(n9056) );
  INV_X1 U10396 ( .A(n9062), .ZN(n9048) );
  OAI21_X1 U10397 ( .B1(n9583), .B2(n9048), .A(n9047), .ZN(n9055) );
  AOI21_X1 U10398 ( .B1(n9050), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9049), .ZN(
        n9053) );
  NAND2_X1 U10399 ( .A1(n9062), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9051) );
  OAI21_X1 U10400 ( .B1(n9062), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9051), .ZN(
        n9052) );
  NOR2_X1 U10401 ( .A1(n9053), .A2(n9052), .ZN(n9059) );
  AOI211_X1 U10402 ( .C1(n9053), .C2(n9052), .A(n9059), .B(n9591), .ZN(n9054)
         );
  AOI211_X1 U10403 ( .C1(n9597), .C2(n9056), .A(n9055), .B(n9054), .ZN(n9057)
         );
  OAI21_X1 U10404 ( .B1(n9586), .B2(n9058), .A(n9057), .ZN(P1_U3259) );
  INV_X1 U10405 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9073) );
  AOI21_X1 U10406 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9062), .A(n9059), .ZN(
        n9060) );
  XNOR2_X1 U10407 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9060), .ZN(n9067) );
  INV_X1 U10408 ( .A(n9067), .ZN(n9065) );
  OAI21_X1 U10409 ( .B1(n9062), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9061), .ZN(
        n9063) );
  XNOR2_X1 U10410 ( .A(n9063), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9066) );
  OAI21_X1 U10411 ( .B1(n9066), .B2(n9558), .A(n9583), .ZN(n9064) );
  AOI21_X1 U10412 ( .B1(n9065), .B2(n9575), .A(n9064), .ZN(n9069) );
  AOI22_X1 U10413 ( .A1(n9067), .A2(n9575), .B1(n9597), .B2(n9066), .ZN(n9068)
         );
  MUX2_X1 U10414 ( .A(n9069), .B(n9068), .S(n9607), .Z(n9072) );
  INV_X1 U10415 ( .A(n9070), .ZN(n9071) );
  OAI211_X1 U10416 ( .C1(n9073), .C2(n9586), .A(n9072), .B(n9071), .ZN(
        P1_U3260) );
  INV_X1 U10417 ( .A(n9431), .ZN(n9339) );
  NAND2_X1 U10418 ( .A1(n9334), .A2(n9339), .ZN(n9335) );
  NOR2_X1 U10419 ( .A1(n9317), .A2(n9419), .ZN(n9296) );
  INV_X1 U10420 ( .A(n9415), .ZN(n9284) );
  INV_X1 U10421 ( .A(n9411), .ZN(n9267) );
  XNOR2_X1 U10422 ( .A(n9079), .B(n9074), .ZN(n9352) );
  NAND2_X1 U10423 ( .A1(n9352), .A2(n9313), .ZN(n9078) );
  AOI21_X1 U10424 ( .B1(n9075), .B2(P1_B_REG_SCAN_IN), .A(n9492), .ZN(n9134)
         );
  NAND2_X1 U10425 ( .A1(n9134), .A2(n9076), .ZN(n9357) );
  NOR2_X1 U10426 ( .A1(n4393), .A2(n9357), .ZN(n9081) );
  AOI21_X1 U10427 ( .B1(n4393), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9081), .ZN(
        n9077) );
  OAI211_X1 U10428 ( .C1(n9354), .C2(n9338), .A(n9078), .B(n9077), .ZN(
        P1_U3261) );
  INV_X1 U10429 ( .A(n9079), .ZN(n9356) );
  NAND2_X1 U10430 ( .A1(n9080), .A2(n9137), .ZN(n9355) );
  NAND3_X1 U10431 ( .A1(n9356), .A2(n9313), .A3(n9355), .ZN(n9083) );
  AOI21_X1 U10432 ( .B1(n4393), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9081), .ZN(
        n9082) );
  OAI211_X1 U10433 ( .C1(n9359), .C2(n9338), .A(n9083), .B(n9082), .ZN(
        P1_U3262) );
  INV_X1 U10434 ( .A(n9084), .ZN(n9438) );
  NOR2_X1 U10435 ( .A1(n9438), .A2(n9348), .ZN(n9085) );
  NOR2_X1 U10436 ( .A1(n9426), .A2(n9304), .ZN(n9088) );
  INV_X1 U10437 ( .A(n9426), .ZN(n9319) );
  OAI21_X1 U10438 ( .B1(n9254), .B2(n9267), .A(n9263), .ZN(n9091) );
  NAND2_X1 U10439 ( .A1(n9225), .A2(n9238), .ZN(n9094) );
  NOR2_X1 U10440 ( .A1(n9225), .A2(n9238), .ZN(n9093) );
  OAI21_X1 U10441 ( .B1(n9095), .B2(n9096), .A(n9206), .ZN(n9098) );
  NAND2_X1 U10442 ( .A1(n9096), .A2(n9095), .ZN(n9097) );
  NAND2_X1 U10443 ( .A1(n9098), .A2(n9097), .ZN(n9191) );
  NAND2_X1 U10444 ( .A1(n9198), .A2(n9210), .ZN(n9099) );
  NAND2_X1 U10445 ( .A1(n9165), .A2(n9103), .ZN(n9104) );
  OAI21_X1 U10446 ( .B1(n4710), .B2(n9168), .A(n9146), .ZN(n9106) );
  XNOR2_X1 U10447 ( .A(n9106), .B(n9131), .ZN(n9360) );
  INV_X1 U10448 ( .A(n9360), .ZN(n9145) );
  INV_X1 U10449 ( .A(n9110), .ZN(n9112) );
  NAND2_X1 U10450 ( .A1(n9286), .A2(n9287), .ZN(n9285) );
  NAND2_X1 U10451 ( .A1(n9285), .A2(n9116), .ZN(n9272) );
  OAI21_X1 U10452 ( .B1(n9272), .B2(n9118), .A(n9117), .ZN(n9251) );
  INV_X1 U10453 ( .A(n9257), .ZN(n9252) );
  NAND2_X1 U10454 ( .A1(n9153), .A2(n9154), .ZN(n9152) );
  NAND2_X1 U10455 ( .A1(n9152), .A2(n9129), .ZN(n9130) );
  XOR2_X1 U10456 ( .A(n9131), .B(n9130), .Z(n9136) );
  AOI22_X1 U10457 ( .A1(n9134), .A2(n9133), .B1(n9303), .B2(n9132), .ZN(n9135)
         );
  OAI21_X1 U10458 ( .B1(n9136), .B2(n9488), .A(n9135), .ZN(n9364) );
  OAI21_X1 U10459 ( .B1(n9148), .B2(n9361), .A(n9137), .ZN(n9362) );
  NOR2_X1 U10460 ( .A1(n9362), .A2(n9138), .ZN(n9143) );
  INV_X1 U10461 ( .A(n9139), .ZN(n9140) );
  AOI22_X1 U10462 ( .A1(n4393), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9140), .B2(
        n9499), .ZN(n9141) );
  OAI21_X1 U10463 ( .B1(n9361), .B2(n9338), .A(n9141), .ZN(n9142) );
  AOI211_X1 U10464 ( .C1(n9364), .C2(n9614), .A(n9143), .B(n9142), .ZN(n9144)
         );
  OAI21_X1 U10465 ( .B1(n9145), .B2(n9351), .A(n9144), .ZN(P1_U3355) );
  AOI21_X1 U10466 ( .B1(n9367), .B2(n9159), .A(n9148), .ZN(n9368) );
  INV_X1 U10467 ( .A(n9149), .ZN(n9150) );
  AOI22_X1 U10468 ( .A1(n4393), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9150), .B2(
        n9499), .ZN(n9151) );
  OAI21_X1 U10469 ( .B1(n4710), .B2(n9338), .A(n9151), .ZN(n9157) );
  OAI21_X1 U10470 ( .B1(n9154), .B2(n9153), .A(n9152), .ZN(n9156) );
  XNOR2_X1 U10471 ( .A(n9158), .B(n9167), .ZN(n9376) );
  INV_X1 U10472 ( .A(n9176), .ZN(n9161) );
  INV_X1 U10473 ( .A(n9159), .ZN(n9160) );
  AOI211_X1 U10474 ( .C1(n9373), .C2(n9161), .A(n9668), .B(n9160), .ZN(n9372)
         );
  INV_X1 U10475 ( .A(n9162), .ZN(n9163) );
  AOI22_X1 U10476 ( .A1(n4393), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9163), .B2(
        n9499), .ZN(n9164) );
  OAI21_X1 U10477 ( .B1(n9165), .B2(n9338), .A(n9164), .ZN(n9173) );
  AOI211_X1 U10478 ( .C1(n9167), .C2(n9166), .A(n9488), .B(n4444), .ZN(n9171)
         );
  OAI22_X1 U10479 ( .A1(n9169), .A2(n9491), .B1(n9168), .B2(n9492), .ZN(n9170)
         );
  NOR2_X1 U10480 ( .A1(n9171), .A2(n9170), .ZN(n9375) );
  NOR2_X1 U10481 ( .A1(n9375), .A2(n4393), .ZN(n9172) );
  AOI211_X1 U10482 ( .C1(n9372), .C2(n9507), .A(n9173), .B(n9172), .ZN(n9174)
         );
  OAI21_X1 U10483 ( .B1(n9376), .B2(n9351), .A(n9174), .ZN(P1_U3264) );
  XNOR2_X1 U10484 ( .A(n9175), .B(n9183), .ZN(n9381) );
  AOI21_X1 U10485 ( .B1(n9377), .B2(n9192), .A(n9176), .ZN(n9378) );
  AOI22_X1 U10486 ( .A1(n4393), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9177), .B2(
        n9499), .ZN(n9178) );
  OAI21_X1 U10487 ( .B1(n9179), .B2(n9338), .A(n9178), .ZN(n9189) );
  INV_X1 U10488 ( .A(n9180), .ZN(n9181) );
  NOR2_X1 U10489 ( .A1(n9182), .A2(n9181), .ZN(n9184) );
  XNOR2_X1 U10490 ( .A(n9184), .B(n9183), .ZN(n9187) );
  AOI222_X1 U10491 ( .A1(n9308), .A2(n9187), .B1(n9186), .B2(n9305), .C1(n9185), .C2(n9303), .ZN(n9380) );
  NOR2_X1 U10492 ( .A1(n9380), .A2(n4393), .ZN(n9188) );
  AOI211_X1 U10493 ( .C1(n9378), .C2(n9313), .A(n9189), .B(n9188), .ZN(n9190)
         );
  OAI21_X1 U10494 ( .B1(n9381), .B2(n9351), .A(n9190), .ZN(P1_U3265) );
  XOR2_X1 U10495 ( .A(n9200), .B(n9191), .Z(n9386) );
  INV_X1 U10496 ( .A(n9211), .ZN(n9194) );
  INV_X1 U10497 ( .A(n9192), .ZN(n9193) );
  AOI21_X1 U10498 ( .B1(n9382), .B2(n9194), .A(n9193), .ZN(n9383) );
  INV_X1 U10499 ( .A(n9195), .ZN(n9196) );
  AOI22_X1 U10500 ( .A1(n4393), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9196), .B2(
        n9499), .ZN(n9197) );
  OAI21_X1 U10501 ( .B1(n9198), .B2(n9338), .A(n9197), .ZN(n9204) );
  XOR2_X1 U10502 ( .A(n9200), .B(n9199), .Z(n9202) );
  AOI222_X1 U10503 ( .A1(n9308), .A2(n9202), .B1(n9229), .B2(n9303), .C1(n9201), .C2(n9305), .ZN(n9385) );
  NOR2_X1 U10504 ( .A1(n9385), .A2(n4393), .ZN(n9203) );
  AOI211_X1 U10505 ( .C1(n9383), .C2(n9313), .A(n9204), .B(n9203), .ZN(n9205)
         );
  OAI21_X1 U10506 ( .B1(n9386), .B2(n9351), .A(n9205), .ZN(P1_U3266) );
  XNOR2_X1 U10507 ( .A(n9206), .B(n9207), .ZN(n9391) );
  AOI22_X1 U10508 ( .A1(n9389), .A2(n9500), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4393), .ZN(n9218) );
  XNOR2_X1 U10509 ( .A(n9208), .B(n9207), .ZN(n9209) );
  OAI222_X1 U10510 ( .A1(n9491), .A2(n9238), .B1(n9492), .B2(n9210), .C1(n9209), .C2(n9488), .ZN(n9387) );
  AOI211_X1 U10511 ( .C1(n9389), .C2(n9220), .A(n9668), .B(n9211), .ZN(n9388)
         );
  INV_X1 U10512 ( .A(n9388), .ZN(n9215) );
  INV_X1 U10513 ( .A(n9212), .ZN(n9213) );
  OAI22_X1 U10514 ( .A1(n9215), .A2(n9214), .B1(n9605), .B2(n9213), .ZN(n9216)
         );
  OAI21_X1 U10515 ( .B1(n9387), .B2(n9216), .A(n9614), .ZN(n9217) );
  OAI211_X1 U10516 ( .C1(n9391), .C2(n9351), .A(n9218), .B(n9217), .ZN(
        P1_U3267) );
  XNOR2_X1 U10517 ( .A(n9219), .B(n9227), .ZN(n9396) );
  INV_X1 U10518 ( .A(n9220), .ZN(n9221) );
  AOI21_X1 U10519 ( .B1(n9392), .B2(n4702), .A(n9221), .ZN(n9393) );
  INV_X1 U10520 ( .A(n9222), .ZN(n9223) );
  AOI22_X1 U10521 ( .A1(n4393), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9223), .B2(
        n9499), .ZN(n9224) );
  OAI21_X1 U10522 ( .B1(n9225), .B2(n9338), .A(n9224), .ZN(n9232) );
  XOR2_X1 U10523 ( .A(n9227), .B(n9226), .Z(n9230) );
  AOI222_X1 U10524 ( .A1(n9308), .A2(n9230), .B1(n9229), .B2(n9305), .C1(n9228), .C2(n9303), .ZN(n9395) );
  NOR2_X1 U10525 ( .A1(n9395), .A2(n4393), .ZN(n9231) );
  AOI211_X1 U10526 ( .C1(n9393), .C2(n9313), .A(n9232), .B(n9231), .ZN(n9233)
         );
  OAI21_X1 U10527 ( .B1(n9396), .B2(n9351), .A(n9233), .ZN(P1_U3268) );
  XOR2_X1 U10528 ( .A(n9236), .B(n9234), .Z(n9401) );
  XOR2_X1 U10529 ( .A(n9236), .B(n9235), .Z(n9237) );
  OAI222_X1 U10530 ( .A1(n9492), .A2(n9238), .B1(n9491), .B2(n9275), .C1(n9237), .C2(n9488), .ZN(n9397) );
  AOI211_X1 U10531 ( .C1(n9399), .C2(n9247), .A(n9668), .B(n9239), .ZN(n9398)
         );
  NAND2_X1 U10532 ( .A1(n9398), .A2(n9507), .ZN(n9243) );
  INV_X1 U10533 ( .A(n9240), .ZN(n9241) );
  AOI22_X1 U10534 ( .A1(n4393), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9499), .B2(
        n9241), .ZN(n9242) );
  OAI211_X1 U10535 ( .C1(n9244), .C2(n9338), .A(n9243), .B(n9242), .ZN(n9245)
         );
  AOI21_X1 U10536 ( .B1(n9397), .B2(n9614), .A(n9245), .ZN(n9246) );
  OAI21_X1 U10537 ( .B1(n9401), .B2(n9351), .A(n9246), .ZN(P1_U3269) );
  AOI21_X1 U10538 ( .B1(n9264), .B2(n9405), .A(n9668), .ZN(n9248) );
  AND2_X1 U10539 ( .A1(n9248), .A2(n9247), .ZN(n9404) );
  NOR2_X1 U10540 ( .A1(n9605), .A2(n9249), .ZN(n9256) );
  AOI21_X1 U10541 ( .B1(n9252), .B2(n9251), .A(n9250), .ZN(n9253) );
  OAI222_X1 U10542 ( .A1(n9492), .A2(n9255), .B1(n9491), .B2(n9254), .C1(n9488), .C2(n9253), .ZN(n9403) );
  AOI211_X1 U10543 ( .C1(n9404), .C2(n9607), .A(n9256), .B(n9403), .ZN(n9262)
         );
  NAND2_X1 U10544 ( .A1(n9258), .A2(n9257), .ZN(n9402) );
  NAND3_X1 U10545 ( .A1(n4664), .A2(n9259), .A3(n9402), .ZN(n9261) );
  AOI22_X1 U10546 ( .A1(n9405), .A2(n9500), .B1(n4393), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n9260) );
  OAI211_X1 U10547 ( .C1(n4393), .C2(n9262), .A(n9261), .B(n9260), .ZN(
        P1_U3270) );
  XNOR2_X1 U10548 ( .A(n9263), .B(n9273), .ZN(n9413) );
  INV_X1 U10549 ( .A(n9280), .ZN(n9266) );
  INV_X1 U10550 ( .A(n9264), .ZN(n9265) );
  AOI211_X1 U10551 ( .C1(n9411), .C2(n9266), .A(n9668), .B(n9265), .ZN(n9410)
         );
  NOR2_X1 U10552 ( .A1(n9267), .A2(n9338), .ZN(n9271) );
  OAI22_X1 U10553 ( .A1(n9614), .A2(n9269), .B1(n9268), .B2(n9605), .ZN(n9270)
         );
  AOI211_X1 U10554 ( .C1(n9410), .C2(n9507), .A(n9271), .B(n9270), .ZN(n9278)
         );
  XOR2_X1 U10555 ( .A(n9273), .B(n9272), .Z(n9274) );
  OAI222_X1 U10556 ( .A1(n9491), .A2(n9276), .B1(n9492), .B2(n9275), .C1(n9274), .C2(n9488), .ZN(n9409) );
  NAND2_X1 U10557 ( .A1(n9409), .A2(n9614), .ZN(n9277) );
  OAI211_X1 U10558 ( .C1(n9413), .C2(n9351), .A(n9278), .B(n9277), .ZN(
        P1_U3271) );
  XNOR2_X1 U10559 ( .A(n9279), .B(n9287), .ZN(n9418) );
  INV_X1 U10560 ( .A(n9296), .ZN(n9281) );
  AOI211_X1 U10561 ( .C1(n9415), .C2(n9281), .A(n9668), .B(n9280), .ZN(n9414)
         );
  AOI22_X1 U10562 ( .A1(n4393), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9282), .B2(
        n9499), .ZN(n9283) );
  OAI21_X1 U10563 ( .B1(n9284), .B2(n9338), .A(n9283), .ZN(n9292) );
  OAI21_X1 U10564 ( .B1(n9287), .B2(n9286), .A(n9285), .ZN(n9290) );
  AOI222_X1 U10565 ( .A1(n9308), .A2(n9290), .B1(n9289), .B2(n9305), .C1(n9288), .C2(n9303), .ZN(n9417) );
  NOR2_X1 U10566 ( .A1(n9417), .A2(n4393), .ZN(n9291) );
  AOI211_X1 U10567 ( .C1(n9414), .C2(n9507), .A(n9292), .B(n9291), .ZN(n9293)
         );
  OAI21_X1 U10568 ( .B1(n9351), .B2(n9418), .A(n9293), .ZN(P1_U3272) );
  XNOR2_X1 U10569 ( .A(n9294), .B(n9302), .ZN(n9423) );
  AND2_X1 U10570 ( .A1(n9317), .A2(n9419), .ZN(n9295) );
  NOR2_X1 U10571 ( .A1(n9296), .A2(n9295), .ZN(n9420) );
  OAI22_X1 U10572 ( .A1(n9298), .A2(n9338), .B1(n9297), .B2(n9614), .ZN(n9312)
         );
  INV_X1 U10573 ( .A(n9299), .ZN(n9300) );
  NOR2_X1 U10574 ( .A1(n4482), .A2(n9300), .ZN(n9301) );
  XOR2_X1 U10575 ( .A(n9302), .B(n9301), .Z(n9307) );
  AOI222_X1 U10576 ( .A1(n9308), .A2(n9307), .B1(n9306), .B2(n9305), .C1(n9304), .C2(n9303), .ZN(n9422) );
  NAND2_X1 U10577 ( .A1(n9499), .A2(n9309), .ZN(n9310) );
  AOI21_X1 U10578 ( .B1(n9422), .B2(n9310), .A(n4393), .ZN(n9311) );
  AOI211_X1 U10579 ( .C1(n9420), .C2(n9313), .A(n9312), .B(n9311), .ZN(n9314)
         );
  OAI21_X1 U10580 ( .B1(n9351), .B2(n9423), .A(n9314), .ZN(P1_U3273) );
  XNOR2_X1 U10581 ( .A(n9316), .B(n9315), .ZN(n9428) );
  INV_X1 U10582 ( .A(n9317), .ZN(n9318) );
  AOI211_X1 U10583 ( .C1(n9426), .C2(n9335), .A(n9668), .B(n9318), .ZN(n9425)
         );
  NOR2_X1 U10584 ( .A1(n9319), .A2(n9338), .ZN(n9323) );
  INV_X1 U10585 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9321) );
  OAI22_X1 U10586 ( .A1(n9614), .A2(n9321), .B1(n9320), .B2(n9605), .ZN(n9322)
         );
  AOI211_X1 U10587 ( .C1(n9425), .C2(n9507), .A(n9323), .B(n9322), .ZN(n9330)
         );
  XNOR2_X1 U10588 ( .A(n9325), .B(n9324), .ZN(n9326) );
  OAI222_X1 U10589 ( .A1(n9492), .A2(n9328), .B1(n9491), .B2(n9327), .C1(n9326), .C2(n9488), .ZN(n9424) );
  NAND2_X1 U10590 ( .A1(n9424), .A2(n9614), .ZN(n9329) );
  OAI211_X1 U10591 ( .C1(n9428), .C2(n9351), .A(n9330), .B(n9329), .ZN(
        P1_U3274) );
  AOI21_X1 U10592 ( .B1(n9344), .B2(n9332), .A(n9331), .ZN(n9333) );
  INV_X1 U10593 ( .A(n9333), .ZN(n9435) );
  INV_X1 U10594 ( .A(n9334), .ZN(n9337) );
  INV_X1 U10595 ( .A(n9335), .ZN(n9336) );
  AOI211_X1 U10596 ( .C1(n9431), .C2(n9337), .A(n9668), .B(n9336), .ZN(n9430)
         );
  NOR2_X1 U10597 ( .A1(n9339), .A2(n9338), .ZN(n9343) );
  INV_X1 U10598 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9341) );
  OAI22_X1 U10599 ( .A1(n9614), .A2(n9341), .B1(n9340), .B2(n9605), .ZN(n9342)
         );
  AOI211_X1 U10600 ( .C1(n9430), .C2(n9507), .A(n9343), .B(n9342), .ZN(n9350)
         );
  XNOR2_X1 U10601 ( .A(n9345), .B(n9344), .ZN(n9346) );
  OAI222_X1 U10602 ( .A1(n9491), .A2(n9348), .B1(n9492), .B2(n9347), .C1(n9488), .C2(n9346), .ZN(n9429) );
  NAND2_X1 U10603 ( .A1(n9429), .A2(n9614), .ZN(n9349) );
  OAI211_X1 U10604 ( .C1(n9435), .C2(n9351), .A(n9350), .B(n9349), .ZN(
        P1_U3275) );
  NAND2_X1 U10605 ( .A1(n9352), .A2(n9503), .ZN(n9353) );
  OAI211_X1 U10606 ( .C1(n9354), .C2(n9666), .A(n9353), .B(n9357), .ZN(n9443)
         );
  MUX2_X1 U10607 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9443), .S(n9683), .Z(
        P1_U3554) );
  NAND3_X1 U10608 ( .A1(n9356), .A2(n9503), .A3(n9355), .ZN(n9358) );
  OAI211_X1 U10609 ( .C1(n9359), .C2(n9666), .A(n9358), .B(n9357), .ZN(n9444)
         );
  MUX2_X1 U10610 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9444), .S(n9683), .Z(
        P1_U3553) );
  NAND2_X1 U10611 ( .A1(n9360), .A2(n9528), .ZN(n9366) );
  OAI22_X1 U10612 ( .A1(n9362), .A2(n9668), .B1(n9361), .B2(n9666), .ZN(n9363)
         );
  NOR2_X1 U10613 ( .A1(n9364), .A2(n9363), .ZN(n9365) );
  NAND2_X1 U10614 ( .A1(n9366), .A2(n9365), .ZN(n9445) );
  MUX2_X1 U10615 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9445), .S(n9683), .Z(
        P1_U3552) );
  AOI22_X1 U10616 ( .A1(n9368), .A2(n9503), .B1(n9432), .B2(n9367), .ZN(n9369)
         );
  OAI211_X1 U10617 ( .C1(n9371), .C2(n9434), .A(n9370), .B(n9369), .ZN(n9446)
         );
  MUX2_X1 U10618 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9446), .S(n9683), .Z(
        P1_U3551) );
  AOI21_X1 U10619 ( .B1(n9432), .B2(n9373), .A(n9372), .ZN(n9374) );
  OAI211_X1 U10620 ( .C1(n9376), .C2(n9434), .A(n9375), .B(n9374), .ZN(n9447)
         );
  MUX2_X1 U10621 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9447), .S(n9683), .Z(
        P1_U3550) );
  AOI22_X1 U10622 ( .A1(n9378), .A2(n9503), .B1(n9432), .B2(n9377), .ZN(n9379)
         );
  OAI211_X1 U10623 ( .C1(n9381), .C2(n9434), .A(n9380), .B(n9379), .ZN(n9448)
         );
  MUX2_X1 U10624 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9448), .S(n9683), .Z(
        P1_U3549) );
  AOI22_X1 U10625 ( .A1(n9383), .A2(n9503), .B1(n9432), .B2(n9382), .ZN(n9384)
         );
  OAI211_X1 U10626 ( .C1(n9386), .C2(n9434), .A(n9385), .B(n9384), .ZN(n9449)
         );
  MUX2_X1 U10627 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9449), .S(n9683), .Z(
        P1_U3548) );
  AOI211_X1 U10628 ( .C1(n9432), .C2(n9389), .A(n9388), .B(n9387), .ZN(n9390)
         );
  OAI21_X1 U10629 ( .B1(n9391), .B2(n9434), .A(n9390), .ZN(n9450) );
  MUX2_X1 U10630 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9450), .S(n9683), .Z(
        P1_U3547) );
  AOI22_X1 U10631 ( .A1(n9393), .A2(n9503), .B1(n9432), .B2(n9392), .ZN(n9394)
         );
  OAI211_X1 U10632 ( .C1(n9396), .C2(n9434), .A(n9395), .B(n9394), .ZN(n9451)
         );
  MUX2_X1 U10633 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9451), .S(n9683), .Z(
        P1_U3546) );
  AOI211_X1 U10634 ( .C1(n9432), .C2(n9399), .A(n9398), .B(n9397), .ZN(n9400)
         );
  OAI21_X1 U10635 ( .B1(n9401), .B2(n9434), .A(n9400), .ZN(n9452) );
  MUX2_X1 U10636 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9452), .S(n9683), .Z(
        P1_U3545) );
  NAND2_X1 U10637 ( .A1(n9402), .A2(n9528), .ZN(n9407) );
  AOI211_X1 U10638 ( .C1(n9432), .C2(n9405), .A(n9404), .B(n9403), .ZN(n9406)
         );
  OAI21_X1 U10639 ( .B1(n9408), .B2(n9407), .A(n9406), .ZN(n9453) );
  MUX2_X1 U10640 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9453), .S(n9683), .Z(
        P1_U3544) );
  AOI211_X1 U10641 ( .C1(n9432), .C2(n9411), .A(n9410), .B(n9409), .ZN(n9412)
         );
  OAI21_X1 U10642 ( .B1(n9413), .B2(n9434), .A(n9412), .ZN(n9454) );
  MUX2_X1 U10643 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9454), .S(n9683), .Z(
        P1_U3543) );
  AOI21_X1 U10644 ( .B1(n9432), .B2(n9415), .A(n9414), .ZN(n9416) );
  OAI211_X1 U10645 ( .C1(n9418), .C2(n9434), .A(n9417), .B(n9416), .ZN(n9455)
         );
  MUX2_X1 U10646 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9455), .S(n9683), .Z(
        P1_U3542) );
  AOI22_X1 U10647 ( .A1(n9420), .A2(n9503), .B1(n9432), .B2(n9419), .ZN(n9421)
         );
  OAI211_X1 U10648 ( .C1(n9423), .C2(n9434), .A(n9422), .B(n9421), .ZN(n9456)
         );
  MUX2_X1 U10649 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9456), .S(n9683), .Z(
        P1_U3541) );
  AOI211_X1 U10650 ( .C1(n9432), .C2(n9426), .A(n9425), .B(n9424), .ZN(n9427)
         );
  OAI21_X1 U10651 ( .B1(n9428), .B2(n9434), .A(n9427), .ZN(n9457) );
  MUX2_X1 U10652 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9457), .S(n9683), .Z(
        P1_U3540) );
  AOI211_X1 U10653 ( .C1(n9432), .C2(n9431), .A(n9430), .B(n9429), .ZN(n9433)
         );
  OAI21_X1 U10654 ( .B1(n9435), .B2(n9434), .A(n9433), .ZN(n9458) );
  MUX2_X1 U10655 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9458), .S(n9683), .Z(
        P1_U3539) );
  NAND2_X1 U10656 ( .A1(n9436), .A2(n9528), .ZN(n9442) );
  OAI21_X1 U10657 ( .B1(n9438), .B2(n9666), .A(n9437), .ZN(n9439) );
  NOR2_X1 U10658 ( .A1(n9440), .A2(n9439), .ZN(n9441) );
  NAND2_X1 U10659 ( .A1(n9442), .A2(n9441), .ZN(n9459) );
  MUX2_X1 U10660 ( .A(n9459), .B(P1_REG1_REG_15__SCAN_IN), .S(n9680), .Z(
        P1_U3538) );
  MUX2_X1 U10661 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9443), .S(n9675), .Z(
        P1_U3522) );
  MUX2_X1 U10662 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9444), .S(n9675), .Z(
        P1_U3521) );
  MUX2_X1 U10663 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9445), .S(n9675), .Z(
        P1_U3520) );
  MUX2_X1 U10664 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9446), .S(n9675), .Z(
        P1_U3519) );
  MUX2_X1 U10665 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9447), .S(n9675), .Z(
        P1_U3518) );
  MUX2_X1 U10666 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9448), .S(n9675), .Z(
        P1_U3517) );
  MUX2_X1 U10667 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9449), .S(n9675), .Z(
        P1_U3516) );
  MUX2_X1 U10668 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9450), .S(n9675), .Z(
        P1_U3515) );
  MUX2_X1 U10669 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9451), .S(n9675), .Z(
        P1_U3514) );
  MUX2_X1 U10670 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9452), .S(n9675), .Z(
        P1_U3513) );
  MUX2_X1 U10671 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9453), .S(n9675), .Z(
        P1_U3512) );
  MUX2_X1 U10672 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9454), .S(n9675), .Z(
        P1_U3511) );
  MUX2_X1 U10673 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9455), .S(n9675), .Z(
        P1_U3510) );
  MUX2_X1 U10674 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9456), .S(n9675), .Z(
        P1_U3508) );
  MUX2_X1 U10675 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9457), .S(n9675), .Z(
        P1_U3505) );
  MUX2_X1 U10676 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9458), .S(n9675), .Z(
        P1_U3502) );
  MUX2_X1 U10677 ( .A(n9459), .B(P1_REG0_REG_15__SCAN_IN), .S(n9674), .Z(
        P1_U3499) );
  NAND3_X1 U10678 ( .A1(n9460), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9462) );
  OAI22_X1 U10679 ( .A1(n9463), .A2(n9462), .B1(n9461), .B2(n9468), .ZN(n9464)
         );
  INV_X1 U10680 ( .A(n9464), .ZN(n9465) );
  OAI21_X1 U10681 ( .B1(n9467), .B2(n9466), .A(n9465), .ZN(P1_U3322) );
  OAI222_X1 U10682 ( .A1(n9473), .A2(n9472), .B1(P1_U3084), .B2(n9470), .C1(
        n9469), .C2(n9468), .ZN(P1_U3324) );
  NAND2_X1 U10683 ( .A1(n9475), .A2(n9474), .ZN(n9477) );
  OAI211_X1 U10684 ( .C1(n9479), .C2(n9478), .A(n9477), .B(n9476), .ZN(
        P1_U3325) );
  MUX2_X1 U10685 ( .A(n9480), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  XNOR2_X1 U10686 ( .A(n9481), .B(n9486), .ZN(n9516) );
  INV_X1 U10687 ( .A(n9482), .ZN(n9483) );
  AOI21_X1 U10688 ( .B1(n9485), .B2(n9484), .A(n9483), .ZN(n9487) );
  XNOR2_X1 U10689 ( .A(n9487), .B(n9486), .ZN(n9489) );
  NOR2_X1 U10690 ( .A1(n9489), .A2(n9488), .ZN(n9495) );
  OAI22_X1 U10691 ( .A1(n9493), .A2(n9492), .B1(n9491), .B2(n9490), .ZN(n9494)
         );
  AOI211_X1 U10692 ( .C1(n9516), .C2(n9496), .A(n9495), .B(n9494), .ZN(n9513)
         );
  INV_X1 U10693 ( .A(n9497), .ZN(n9498) );
  AOI222_X1 U10694 ( .A1(n9501), .A2(n9500), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n4393), .C1(n9499), .C2(n9498), .ZN(n9510) );
  INV_X1 U10695 ( .A(n9501), .ZN(n9512) );
  INV_X1 U10696 ( .A(n9502), .ZN(n9504) );
  OAI211_X1 U10697 ( .C1(n9512), .C2(n9505), .A(n9504), .B(n9503), .ZN(n9511)
         );
  INV_X1 U10698 ( .A(n9511), .ZN(n9506) );
  AOI22_X1 U10699 ( .A1(n9516), .A2(n9508), .B1(n9507), .B2(n9506), .ZN(n9509)
         );
  OAI211_X1 U10700 ( .C1(n4393), .C2(n9513), .A(n9510), .B(n9509), .ZN(
        P1_U3281) );
  OAI21_X1 U10701 ( .B1(n9512), .B2(n9666), .A(n9511), .ZN(n9515) );
  INV_X1 U10702 ( .A(n9513), .ZN(n9514) );
  AOI211_X1 U10703 ( .C1(n9673), .C2(n9516), .A(n9515), .B(n9514), .ZN(n9517)
         );
  AOI22_X1 U10704 ( .A1(n9675), .A2(n9517), .B1(n5325), .B2(n9674), .ZN(
        P1_U3484) );
  AOI22_X1 U10705 ( .A1(n9683), .A2(n9517), .B1(n5328), .B2(n9680), .ZN(
        P1_U3533) );
  OAI22_X1 U10706 ( .A1(n9519), .A2(n9838), .B1(n9518), .B2(n9854), .ZN(n9521)
         );
  AOI211_X1 U10707 ( .C1(n9859), .C2(n9522), .A(n9521), .B(n9520), .ZN(n9524)
         );
  AOI22_X1 U10708 ( .A1(n9879), .A2(n9524), .B1(n9523), .B2(n9877), .ZN(
        P2_U3534) );
  INV_X1 U10709 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9922) );
  AOI22_X1 U10710 ( .A1(n9861), .A2(n9524), .B1(n9922), .B2(n9860), .ZN(
        P2_U3493) );
  OAI211_X1 U10711 ( .C1(n4697), .C2(n9666), .A(n9526), .B(n9525), .ZN(n9527)
         );
  AOI21_X1 U10712 ( .B1(n9529), .B2(n9528), .A(n9527), .ZN(n9548) );
  AOI22_X1 U10713 ( .A1(n9683), .A2(n9548), .B1(n6372), .B2(n9680), .ZN(
        P1_U3537) );
  OAI22_X1 U10714 ( .A1(n9530), .A2(n9668), .B1(n4698), .B2(n9666), .ZN(n9531)
         );
  AOI21_X1 U10715 ( .B1(n9532), .B2(n9673), .A(n9531), .ZN(n9533) );
  AOI22_X1 U10716 ( .A1(n9683), .A2(n9549), .B1(n6366), .B2(n9680), .ZN(
        P1_U3536) );
  OAI21_X1 U10717 ( .B1(n9536), .B2(n9666), .A(n9535), .ZN(n9537) );
  AOI21_X1 U10718 ( .B1(n9538), .B2(n9673), .A(n9537), .ZN(n9539) );
  AND2_X1 U10719 ( .A1(n9540), .A2(n9539), .ZN(n9550) );
  AOI22_X1 U10720 ( .A1(n9683), .A2(n9550), .B1(n6367), .B2(n9680), .ZN(
        P1_U3535) );
  INV_X1 U10721 ( .A(n9541), .ZN(n9546) );
  OAI22_X1 U10722 ( .A1(n9543), .A2(n9668), .B1(n9542), .B2(n9666), .ZN(n9545)
         );
  AOI211_X1 U10723 ( .C1(n9673), .C2(n9546), .A(n9545), .B(n9544), .ZN(n9552)
         );
  AOI22_X1 U10724 ( .A1(n9683), .A2(n9552), .B1(n5310), .B2(n9680), .ZN(
        P1_U3534) );
  INV_X1 U10725 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9547) );
  AOI22_X1 U10726 ( .A1(n9675), .A2(n9548), .B1(n9547), .B2(n9674), .ZN(
        P1_U3496) );
  AOI22_X1 U10727 ( .A1(n9675), .A2(n9549), .B1(n5283), .B2(n9674), .ZN(
        P1_U3493) );
  AOI22_X1 U10728 ( .A1(n9675), .A2(n9550), .B1(n5297), .B2(n9674), .ZN(
        P1_U3490) );
  INV_X1 U10729 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9551) );
  AOI22_X1 U10730 ( .A1(n9675), .A2(n9552), .B1(n9551), .B2(n9674), .ZN(
        P1_U3487) );
  XNOR2_X1 U10731 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X1 U10732 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10160) );
  AOI21_X1 U10733 ( .B1(n9555), .B2(n9554), .A(n9553), .ZN(n9557) );
  OAI21_X1 U10734 ( .B1(n9558), .B2(n9557), .A(n9556), .ZN(n9565) );
  AOI21_X1 U10735 ( .B1(n9561), .B2(n9560), .A(n9559), .ZN(n9563) );
  OAI22_X1 U10736 ( .A1(n9591), .A2(n9563), .B1(n9562), .B2(n9583), .ZN(n9564)
         );
  NOR3_X1 U10737 ( .A1(n9566), .A2(n9565), .A3(n9564), .ZN(n9567) );
  OAI21_X1 U10738 ( .B1(n9586), .B2(n10160), .A(n9567), .ZN(P1_U3245) );
  INV_X1 U10739 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9569) );
  OAI22_X1 U10740 ( .A1(n9586), .A2(n9569), .B1(n9568), .B2(n9583), .ZN(n9570)
         );
  INV_X1 U10741 ( .A(n9570), .ZN(n9582) );
  OAI21_X1 U10742 ( .B1(n9573), .B2(n9572), .A(n9571), .ZN(n9574) );
  NAND2_X1 U10743 ( .A1(n9575), .A2(n9574), .ZN(n9580) );
  OAI211_X1 U10744 ( .C1(n9578), .C2(n9577), .A(n9597), .B(n9576), .ZN(n9579)
         );
  NAND4_X1 U10745 ( .A1(n9582), .A2(n9581), .A3(n9580), .A4(n9579), .ZN(
        P1_U3246) );
  INV_X1 U10746 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9585) );
  OAI22_X1 U10747 ( .A1(n9586), .A2(n9585), .B1(n9584), .B2(n9583), .ZN(n9587)
         );
  INV_X1 U10748 ( .A(n9587), .ZN(n9600) );
  OAI21_X1 U10749 ( .B1(n9590), .B2(n9589), .A(n9588), .ZN(n9598) );
  AOI211_X1 U10750 ( .C1(n9594), .C2(n9593), .A(n9592), .B(n9591), .ZN(n9595)
         );
  AOI211_X1 U10751 ( .C1(n9598), .C2(n9597), .A(n9596), .B(n9595), .ZN(n9599)
         );
  NAND2_X1 U10752 ( .A1(n9600), .A2(n9599), .ZN(P1_U3251) );
  INV_X1 U10753 ( .A(n9601), .ZN(n9611) );
  OAI22_X1 U10754 ( .A1(n9605), .A2(n9604), .B1(n9603), .B2(n9602), .ZN(n9606)
         );
  AOI21_X1 U10755 ( .B1(n9608), .B2(n9607), .A(n9606), .ZN(n9609) );
  OAI211_X1 U10756 ( .C1(n9612), .C2(n9611), .A(n9610), .B(n9609), .ZN(n9613)
         );
  INV_X1 U10757 ( .A(n9613), .ZN(n9615) );
  AOI22_X1 U10758 ( .A1(n4393), .A2(n5428), .B1(n9615), .B2(n9614), .ZN(
        P1_U3286) );
  NOR2_X1 U10759 ( .A1(n9617), .A2(n9616), .ZN(n9643) );
  INV_X1 U10760 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10114) );
  NOR2_X1 U10761 ( .A1(n9633), .A2(n10114), .ZN(P1_U3292) );
  INV_X1 U10762 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9618) );
  NOR2_X1 U10763 ( .A1(n9633), .A2(n9618), .ZN(P1_U3293) );
  INV_X1 U10764 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9619) );
  NOR2_X1 U10765 ( .A1(n9633), .A2(n9619), .ZN(P1_U3294) );
  INV_X1 U10766 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9620) );
  NOR2_X1 U10767 ( .A1(n9633), .A2(n9620), .ZN(P1_U3295) );
  INV_X1 U10768 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9621) );
  NOR2_X1 U10769 ( .A1(n9633), .A2(n9621), .ZN(P1_U3296) );
  INV_X1 U10770 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9622) );
  NOR2_X1 U10771 ( .A1(n9633), .A2(n9622), .ZN(P1_U3297) );
  INV_X1 U10772 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n9623) );
  NOR2_X1 U10773 ( .A1(n9633), .A2(n9623), .ZN(P1_U3298) );
  INV_X1 U10774 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9624) );
  NOR2_X1 U10775 ( .A1(n9633), .A2(n9624), .ZN(P1_U3299) );
  INV_X1 U10776 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9625) );
  NOR2_X1 U10777 ( .A1(n9633), .A2(n9625), .ZN(P1_U3300) );
  INV_X1 U10778 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9626) );
  NOR2_X1 U10779 ( .A1(n9633), .A2(n9626), .ZN(P1_U3301) );
  INV_X1 U10780 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n9627) );
  NOR2_X1 U10781 ( .A1(n9633), .A2(n9627), .ZN(P1_U3302) );
  INV_X1 U10782 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U10783 ( .A1(n9633), .A2(n10198), .ZN(P1_U3303) );
  INV_X1 U10784 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9628) );
  NOR2_X1 U10785 ( .A1(n9633), .A2(n9628), .ZN(P1_U3304) );
  INV_X1 U10786 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9629) );
  NOR2_X1 U10787 ( .A1(n9633), .A2(n9629), .ZN(P1_U3305) );
  NOR2_X1 U10788 ( .A1(n9633), .A2(n9921), .ZN(P1_U3306) );
  NOR2_X1 U10789 ( .A1(n9633), .A2(n10102), .ZN(P1_U3307) );
  INV_X1 U10790 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9630) );
  NOR2_X1 U10791 ( .A1(n9633), .A2(n9630), .ZN(P1_U3308) );
  INV_X1 U10792 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n9631) );
  NOR2_X1 U10793 ( .A1(n9633), .A2(n9631), .ZN(P1_U3309) );
  INV_X1 U10794 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9632) );
  NOR2_X1 U10795 ( .A1(n9633), .A2(n9632), .ZN(P1_U3310) );
  NOR2_X1 U10796 ( .A1(n9643), .A2(n10104), .ZN(P1_U3311) );
  INV_X1 U10797 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9634) );
  NOR2_X1 U10798 ( .A1(n9643), .A2(n9634), .ZN(P1_U3312) );
  INV_X1 U10799 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n9635) );
  NOR2_X1 U10800 ( .A1(n9643), .A2(n9635), .ZN(P1_U3313) );
  INV_X1 U10801 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9636) );
  NOR2_X1 U10802 ( .A1(n9643), .A2(n9636), .ZN(P1_U3314) );
  INV_X1 U10803 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9637) );
  NOR2_X1 U10804 ( .A1(n9643), .A2(n9637), .ZN(P1_U3315) );
  NOR2_X1 U10805 ( .A1(n9643), .A2(n10093), .ZN(P1_U3316) );
  INV_X1 U10806 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n9638) );
  NOR2_X1 U10807 ( .A1(n9643), .A2(n9638), .ZN(P1_U3317) );
  INV_X1 U10808 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n9639) );
  NOR2_X1 U10809 ( .A1(n9643), .A2(n9639), .ZN(P1_U3318) );
  INV_X1 U10810 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9640) );
  NOR2_X1 U10811 ( .A1(n9643), .A2(n9640), .ZN(P1_U3319) );
  INV_X1 U10812 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9641) );
  NOR2_X1 U10813 ( .A1(n9643), .A2(n9641), .ZN(P1_U3320) );
  INV_X1 U10814 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9642) );
  NOR2_X1 U10815 ( .A1(n9643), .A2(n9642), .ZN(P1_U3321) );
  OAI21_X1 U10816 ( .B1(n9645), .B2(n9666), .A(n9644), .ZN(n9647) );
  AOI211_X1 U10817 ( .C1(n9673), .C2(n9648), .A(n9647), .B(n9646), .ZN(n9676)
         );
  INV_X1 U10818 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9975) );
  AOI22_X1 U10819 ( .A1(n9675), .A2(n9676), .B1(n9975), .B2(n9674), .ZN(
        P1_U3457) );
  OAI22_X1 U10820 ( .A1(n9650), .A2(n9668), .B1(n9666), .B2(n9649), .ZN(n9652)
         );
  AOI211_X1 U10821 ( .C1(n9673), .C2(n9653), .A(n9652), .B(n9651), .ZN(n9677)
         );
  INV_X1 U10822 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U10823 ( .A1(n9675), .A2(n9677), .B1(n10128), .B2(n9674), .ZN(
        P1_U3460) );
  OAI22_X1 U10824 ( .A1(n9655), .A2(n9668), .B1(n9654), .B2(n9666), .ZN(n9657)
         );
  AOI211_X1 U10825 ( .C1(n9673), .C2(n9658), .A(n9657), .B(n9656), .ZN(n9678)
         );
  INV_X1 U10826 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9659) );
  AOI22_X1 U10827 ( .A1(n9675), .A2(n9678), .B1(n9659), .B2(n9674), .ZN(
        P1_U3466) );
  OAI22_X1 U10828 ( .A1(n9661), .A2(n9668), .B1(n9660), .B2(n9666), .ZN(n9663)
         );
  AOI211_X1 U10829 ( .C1(n9673), .C2(n9664), .A(n9663), .B(n9662), .ZN(n9679)
         );
  INV_X1 U10830 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U10831 ( .A1(n9675), .A2(n9679), .B1(n10116), .B2(n9674), .ZN(
        P1_U3472) );
  INV_X1 U10832 ( .A(n9665), .ZN(n9672) );
  OAI22_X1 U10833 ( .A1(n9669), .A2(n9668), .B1(n9667), .B2(n9666), .ZN(n9671)
         );
  AOI211_X1 U10834 ( .C1(n9673), .C2(n9672), .A(n9671), .B(n9670), .ZN(n9682)
         );
  AOI22_X1 U10835 ( .A1(n9675), .A2(n9682), .B1(n5352), .B2(n9674), .ZN(
        P1_U3478) );
  AOI22_X1 U10836 ( .A1(n9683), .A2(n9676), .B1(n6591), .B2(n9680), .ZN(
        P1_U3524) );
  AOI22_X1 U10837 ( .A1(n9683), .A2(n9677), .B1(n6335), .B2(n9680), .ZN(
        P1_U3525) );
  AOI22_X1 U10838 ( .A1(n9683), .A2(n9678), .B1(n6332), .B2(n9680), .ZN(
        P1_U3527) );
  AOI22_X1 U10839 ( .A1(n9683), .A2(n9679), .B1(n5442), .B2(n9680), .ZN(
        P1_U3529) );
  AOI22_X1 U10840 ( .A1(n9683), .A2(n9682), .B1(n9681), .B2(n9680), .ZN(
        P1_U3531) );
  AOI22_X1 U10841 ( .A1(n9715), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9711), .ZN(n9690) );
  INV_X1 U10842 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10149) );
  NAND2_X1 U10843 ( .A1(n9711), .A2(n10149), .ZN(n9684) );
  OAI211_X1 U10844 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n9686), .A(n9685), .B(
        n9684), .ZN(n9687) );
  INV_X1 U10845 ( .A(n9687), .ZN(n9689) );
  AOI22_X1 U10846 ( .A1(n9707), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9688) );
  OAI221_X1 U10847 ( .B1(n9691), .B2(n9690), .C1(n4617), .C2(n9689), .A(n9688), 
        .ZN(P2_U3245) );
  INV_X1 U10848 ( .A(n9692), .ZN(n9693) );
  AOI21_X1 U10849 ( .B1(n9707), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n9693), .ZN(
        n9704) );
  NAND2_X1 U10850 ( .A1(n9709), .A2(n9694), .ZN(n9703) );
  OAI211_X1 U10851 ( .C1(n9697), .C2(n9696), .A(n9715), .B(n9695), .ZN(n9702)
         );
  OAI211_X1 U10852 ( .C1(n9700), .C2(n9699), .A(n9711), .B(n9698), .ZN(n9701)
         );
  NAND4_X1 U10853 ( .A1(n9704), .A2(n9703), .A3(n9702), .A4(n9701), .ZN(
        P2_U3253) );
  INV_X1 U10854 ( .A(n9705), .ZN(n9706) );
  AOI21_X1 U10855 ( .B1(n9707), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9706), .ZN(
        n9721) );
  NAND2_X1 U10856 ( .A1(n9709), .A2(n9708), .ZN(n9720) );
  OAI211_X1 U10857 ( .C1(n9713), .C2(n9712), .A(n9711), .B(n9710), .ZN(n9719)
         );
  OAI211_X1 U10858 ( .C1(n9717), .C2(n9716), .A(n9715), .B(n9714), .ZN(n9718)
         );
  NAND4_X1 U10859 ( .A1(n9721), .A2(n9720), .A3(n9719), .A4(n9718), .ZN(
        P2_U3255) );
  AOI21_X1 U10860 ( .B1(n4493), .B2(n9728), .A(n9740), .ZN(n9724) );
  AOI21_X1 U10861 ( .B1(n9724), .B2(n9723), .A(n9722), .ZN(n9827) );
  AOI222_X1 U10862 ( .A1(n9727), .A2(n9726), .B1(P2_REG2_REG_7__SCAN_IN), .B2(
        n4392), .C1(n9776), .C2(n9725), .ZN(n9736) );
  XNOR2_X1 U10863 ( .A(n9729), .B(n9728), .ZN(n9830) );
  INV_X1 U10864 ( .A(n9730), .ZN(n9732) );
  OAI211_X1 U10865 ( .C1(n9732), .C2(n9828), .A(n9845), .B(n9731), .ZN(n9826)
         );
  INV_X1 U10866 ( .A(n9826), .ZN(n9733) );
  AOI22_X1 U10867 ( .A1(n9830), .A2(n9782), .B1(n9734), .B2(n9733), .ZN(n9735)
         );
  OAI211_X1 U10868 ( .C1(n4392), .C2(n9827), .A(n9736), .B(n9735), .ZN(
        P2_U3289) );
  INV_X1 U10869 ( .A(n9737), .ZN(n9742) );
  INV_X1 U10870 ( .A(n9738), .ZN(n9753) );
  AOI21_X1 U10871 ( .B1(n7020), .B2(n9739), .A(n9753), .ZN(n9741) );
  NOR3_X1 U10872 ( .A1(n9742), .A2(n9741), .A3(n9740), .ZN(n9748) );
  OAI22_X1 U10873 ( .A1(n9746), .A2(n9745), .B1(n9744), .B2(n9743), .ZN(n9747)
         );
  NOR2_X1 U10874 ( .A1(n9748), .A2(n9747), .ZN(n9816) );
  INV_X1 U10875 ( .A(n9749), .ZN(n9751) );
  OAI22_X1 U10876 ( .A1(n9785), .A2(n10185), .B1(n9751), .B2(n9750), .ZN(n9752) );
  INV_X1 U10877 ( .A(n9752), .ZN(n9765) );
  XNOR2_X1 U10878 ( .A(n9754), .B(n9753), .ZN(n9817) );
  OR2_X1 U10879 ( .A1(n9755), .A2(n9817), .ZN(n9764) );
  OR2_X1 U10880 ( .A1(n9757), .A2(n9756), .ZN(n9763) );
  AND2_X1 U10881 ( .A1(n9758), .A2(n9813), .ZN(n9759) );
  NOR2_X1 U10882 ( .A1(n9760), .A2(n9759), .ZN(n9814) );
  NAND2_X1 U10883 ( .A1(n9761), .A2(n9814), .ZN(n9762) );
  AND4_X1 U10884 ( .A1(n9765), .A2(n9764), .A3(n9763), .A4(n9762), .ZN(n9766)
         );
  OAI21_X1 U10885 ( .B1(n4392), .B2(n9816), .A(n9766), .ZN(P2_U3292) );
  OAI21_X1 U10886 ( .B1(n9769), .B2(n9768), .A(n9767), .ZN(n9773) );
  AOI222_X1 U10887 ( .A1(n9774), .A2(n9773), .B1(n9772), .B2(n9771), .C1(n6891), .C2(n9770), .ZN(n9775) );
  INV_X1 U10888 ( .A(n9775), .ZN(n9802) );
  AOI21_X1 U10889 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n9776), .A(n9802), .ZN(
        n9786) );
  NAND2_X1 U10890 ( .A1(n9778), .A2(n9845), .ZN(n9777) );
  NAND2_X1 U10891 ( .A1(n9777), .A2(n9854), .ZN(n9780) );
  NOR2_X1 U10892 ( .A1(n9778), .A2(n9838), .ZN(n9796) );
  MUX2_X1 U10893 ( .A(n9780), .B(n9796), .S(n9779), .Z(n9803) );
  XNOR2_X1 U10894 ( .A(n9781), .B(n6904), .ZN(n9804) );
  AOI22_X1 U10895 ( .A1(n9783), .A2(n9803), .B1(n9782), .B2(n9804), .ZN(n9784)
         );
  OAI221_X1 U10896 ( .B1(n4392), .B2(n9786), .C1(n9785), .C2(n9961), .A(n9784), 
        .ZN(P2_U3294) );
  NOR2_X1 U10897 ( .A1(n9788), .A2(n9787), .ZN(n9789) );
  NOR2_X1 U10898 ( .A1(n9789), .A2(n9951), .ZN(P2_U3297) );
  AND2_X1 U10899 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n9792), .ZN(P2_U3298) );
  AND2_X1 U10900 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9792), .ZN(P2_U3299) );
  AND2_X1 U10901 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9792), .ZN(P2_U3300) );
  AND2_X1 U10902 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9792), .ZN(P2_U3301) );
  AND2_X1 U10903 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9792), .ZN(P2_U3302) );
  NOR2_X1 U10904 ( .A1(n9789), .A2(n9979), .ZN(P2_U3303) );
  AND2_X1 U10905 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9792), .ZN(P2_U3304) );
  AND2_X1 U10906 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9792), .ZN(P2_U3305) );
  AND2_X1 U10907 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9792), .ZN(P2_U3306) );
  AND2_X1 U10908 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9792), .ZN(P2_U3307) );
  AND2_X1 U10909 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9792), .ZN(P2_U3308) );
  AND2_X1 U10910 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9792), .ZN(P2_U3309) );
  AND2_X1 U10911 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9792), .ZN(P2_U3310) );
  NOR2_X1 U10912 ( .A1(n9789), .A2(n9980), .ZN(P2_U3311) );
  AND2_X1 U10913 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n9792), .ZN(P2_U3312) );
  AND2_X1 U10914 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9792), .ZN(P2_U3313) );
  AND2_X1 U10915 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9792), .ZN(P2_U3314) );
  INV_X1 U10916 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10169) );
  NOR2_X1 U10917 ( .A1(n9789), .A2(n10169), .ZN(P2_U3315) );
  AND2_X1 U10918 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9792), .ZN(P2_U3316) );
  AND2_X1 U10919 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9792), .ZN(P2_U3317) );
  AND2_X1 U10920 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9792), .ZN(P2_U3318) );
  AND2_X1 U10921 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9792), .ZN(P2_U3319) );
  AND2_X1 U10922 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9792), .ZN(P2_U3320) );
  AND2_X1 U10923 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9792), .ZN(P2_U3321) );
  AND2_X1 U10924 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9792), .ZN(P2_U3322) );
  INV_X1 U10925 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10105) );
  NOR2_X1 U10926 ( .A1(n9789), .A2(n10105), .ZN(P2_U3323) );
  AND2_X1 U10927 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9792), .ZN(P2_U3324) );
  AND2_X1 U10928 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9792), .ZN(P2_U3325) );
  NOR2_X1 U10929 ( .A1(n9789), .A2(n9937), .ZN(P2_U3326) );
  AOI22_X1 U10930 ( .A1(n9794), .A2(n9791), .B1(n9790), .B2(n9792), .ZN(
        P2_U3437) );
  AOI22_X1 U10931 ( .A1(n9794), .A2(n9793), .B1(n6279), .B2(n9792), .ZN(
        P2_U3438) );
  AOI22_X1 U10932 ( .A1(n9796), .A2(n9795), .B1(n9844), .B2(n6890), .ZN(n9797)
         );
  OAI211_X1 U10933 ( .C1(n9799), .C2(n9848), .A(n9798), .B(n9797), .ZN(n9800)
         );
  INV_X1 U10934 ( .A(n9800), .ZN(n9863) );
  INV_X1 U10935 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9801) );
  AOI22_X1 U10936 ( .A1(n9861), .A2(n9863), .B1(n9801), .B2(n9860), .ZN(
        P2_U3454) );
  AOI211_X1 U10937 ( .C1(n9859), .C2(n9804), .A(n9803), .B(n9802), .ZN(n9864)
         );
  INV_X1 U10938 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9805) );
  AOI22_X1 U10939 ( .A1(n9861), .A2(n9864), .B1(n9805), .B2(n9860), .ZN(
        P2_U3457) );
  AOI22_X1 U10940 ( .A1(n9807), .A2(n9845), .B1(n9844), .B2(n9806), .ZN(n9808)
         );
  NAND2_X1 U10941 ( .A1(n9809), .A2(n9808), .ZN(n9810) );
  AOI21_X1 U10942 ( .B1(n9859), .B2(n9811), .A(n9810), .ZN(n9865) );
  INV_X1 U10943 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9812) );
  AOI22_X1 U10944 ( .A1(n9861), .A2(n9865), .B1(n9812), .B2(n9860), .ZN(
        P2_U3460) );
  AOI22_X1 U10945 ( .A1(n9814), .A2(n9845), .B1(n9844), .B2(n9813), .ZN(n9815)
         );
  OAI211_X1 U10946 ( .C1(n9817), .C2(n9848), .A(n9816), .B(n9815), .ZN(n9818)
         );
  INV_X1 U10947 ( .A(n9818), .ZN(n9867) );
  INV_X1 U10948 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9819) );
  AOI22_X1 U10949 ( .A1(n9861), .A2(n9867), .B1(n9819), .B2(n9860), .ZN(
        P2_U3463) );
  OAI21_X1 U10950 ( .B1(n9821), .B2(n9854), .A(n9820), .ZN(n9823) );
  AOI211_X1 U10951 ( .C1(n9859), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9869)
         );
  INV_X1 U10952 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9825) );
  AOI22_X1 U10953 ( .A1(n9861), .A2(n9869), .B1(n9825), .B2(n9860), .ZN(
        P2_U3466) );
  OAI211_X1 U10954 ( .C1(n9828), .C2(n9854), .A(n9827), .B(n9826), .ZN(n9829)
         );
  AOI21_X1 U10955 ( .B1(n9859), .B2(n9830), .A(n9829), .ZN(n9871) );
  INV_X1 U10956 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U10957 ( .A1(n9861), .A2(n9871), .B1(n9831), .B2(n9860), .ZN(
        P2_U3472) );
  NOR2_X1 U10958 ( .A1(n9832), .A2(n9854), .ZN(n9834) );
  AOI211_X1 U10959 ( .C1(n9845), .C2(n9835), .A(n9834), .B(n9833), .ZN(n9873)
         );
  INV_X1 U10960 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9836) );
  AOI22_X1 U10961 ( .A1(n9861), .A2(n9873), .B1(n9836), .B2(n9860), .ZN(
        P2_U3475) );
  OAI22_X1 U10962 ( .A1(n9839), .A2(n9838), .B1(n9837), .B2(n9854), .ZN(n9840)
         );
  NOR2_X1 U10963 ( .A1(n9841), .A2(n9840), .ZN(n9875) );
  INV_X1 U10964 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9842) );
  AOI22_X1 U10965 ( .A1(n9861), .A2(n9875), .B1(n9842), .B2(n9860), .ZN(
        P2_U3481) );
  AOI22_X1 U10966 ( .A1(n9846), .A2(n9845), .B1(n9844), .B2(n9843), .ZN(n9847)
         );
  OAI21_X1 U10967 ( .B1(n9849), .B2(n9848), .A(n9847), .ZN(n9850) );
  NOR2_X1 U10968 ( .A1(n9851), .A2(n9850), .ZN(n9876) );
  INV_X1 U10969 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9852) );
  AOI22_X1 U10970 ( .A1(n9861), .A2(n9876), .B1(n9852), .B2(n9860), .ZN(
        P2_U3484) );
  OAI21_X1 U10971 ( .B1(n9855), .B2(n9854), .A(n9853), .ZN(n9857) );
  AOI211_X1 U10972 ( .C1(n9859), .C2(n9858), .A(n9857), .B(n9856), .ZN(n9878)
         );
  INV_X1 U10973 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U10974 ( .A1(n9861), .A2(n9878), .B1(n10130), .B2(n9860), .ZN(
        P2_U3487) );
  AOI22_X1 U10975 ( .A1(n9879), .A2(n9863), .B1(n9862), .B2(n9877), .ZN(
        P2_U3521) );
  AOI22_X1 U10976 ( .A1(n9879), .A2(n9864), .B1(n6469), .B2(n9877), .ZN(
        P2_U3522) );
  AOI22_X1 U10977 ( .A1(n9879), .A2(n9865), .B1(n6471), .B2(n9877), .ZN(
        P2_U3523) );
  AOI22_X1 U10978 ( .A1(n9879), .A2(n9867), .B1(n9866), .B2(n9877), .ZN(
        P2_U3524) );
  AOI22_X1 U10979 ( .A1(n9879), .A2(n9869), .B1(n9868), .B2(n9877), .ZN(
        P2_U3525) );
  AOI22_X1 U10980 ( .A1(n9879), .A2(n9871), .B1(n9870), .B2(n9877), .ZN(
        P2_U3527) );
  AOI22_X1 U10981 ( .A1(n9879), .A2(n9873), .B1(n9872), .B2(n9877), .ZN(
        P2_U3528) );
  AOI22_X1 U10982 ( .A1(n9879), .A2(n9875), .B1(n9874), .B2(n9877), .ZN(
        P2_U3530) );
  AOI22_X1 U10983 ( .A1(n9879), .A2(n9876), .B1(n6481), .B2(n9877), .ZN(
        P2_U3531) );
  AOI22_X1 U10984 ( .A1(n9879), .A2(n9878), .B1(n9940), .B2(n9877), .ZN(
        P2_U3532) );
  INV_X1 U10985 ( .A(n9880), .ZN(n9881) );
  NAND2_X1 U10986 ( .A1(n9882), .A2(n9881), .ZN(n9883) );
  XNOR2_X1 U10987 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9883), .ZN(ADD_1071_U5) );
  XOR2_X1 U10988 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10989 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(ADD_1071_U56) );
  OAI21_X1 U10990 ( .B1(n9889), .B2(n9888), .A(n9887), .ZN(ADD_1071_U57) );
  OAI21_X1 U10991 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(ADD_1071_U58) );
  OAI21_X1 U10992 ( .B1(n9895), .B2(n9894), .A(n9893), .ZN(ADD_1071_U59) );
  OAI21_X1 U10993 ( .B1(n9898), .B2(n9897), .A(n9896), .ZN(ADD_1071_U60) );
  OAI21_X1 U10994 ( .B1(n9901), .B2(n9900), .A(n9899), .ZN(ADD_1071_U61) );
  AOI21_X1 U10995 ( .B1(n9904), .B2(n9903), .A(n9902), .ZN(ADD_1071_U62) );
  AOI21_X1 U10996 ( .B1(n9907), .B2(n9906), .A(n9905), .ZN(ADD_1071_U63) );
  INV_X1 U10997 ( .A(SI_21_), .ZN(n9909) );
  AOI22_X1 U10998 ( .A1(n9909), .A2(keyinput8), .B1(keyinput19), .B2(n9569), 
        .ZN(n9908) );
  OAI221_X1 U10999 ( .B1(n9909), .B2(keyinput8), .C1(n9569), .C2(keyinput19), 
        .A(n9908), .ZN(n9919) );
  AOI22_X1 U11000 ( .A1(n9911), .A2(keyinput57), .B1(keyinput30), .B2(n9585), 
        .ZN(n9910) );
  OAI221_X1 U11001 ( .B1(n9911), .B2(keyinput57), .C1(n9585), .C2(keyinput30), 
        .A(n9910), .ZN(n9918) );
  AOI22_X1 U11002 ( .A1(n6007), .A2(keyinput36), .B1(keyinput10), .B2(n9913), 
        .ZN(n9912) );
  OAI221_X1 U11003 ( .B1(n6007), .B2(keyinput36), .C1(n9913), .C2(keyinput10), 
        .A(n9912), .ZN(n9917) );
  XNOR2_X1 U11004 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(keyinput62), .ZN(n9915)
         );
  XNOR2_X1 U11005 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput1), .ZN(n9914) );
  NAND2_X1 U11006 ( .A1(n9915), .A2(n9914), .ZN(n9916) );
  NOR4_X1 U11007 ( .A1(n9919), .A2(n9918), .A3(n9917), .A4(n9916), .ZN(n10213)
         );
  AOI22_X1 U11008 ( .A1(n9922), .A2(keyinput12), .B1(n9921), .B2(keyinput43), 
        .ZN(n9920) );
  OAI221_X1 U11009 ( .B1(n9922), .B2(keyinput12), .C1(n9921), .C2(keyinput43), 
        .A(n9920), .ZN(n9931) );
  XNOR2_X1 U11010 ( .A(n9923), .B(keyinput78), .ZN(n9930) );
  XNOR2_X1 U11011 ( .A(keyinput34), .B(n6367), .ZN(n9929) );
  XNOR2_X1 U11012 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput54), .ZN(n9927) );
  XNOR2_X1 U11013 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(keyinput91), .ZN(n9926)
         );
  XNOR2_X1 U11014 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput121), .ZN(n9925)
         );
  XNOR2_X1 U11015 ( .A(SI_6_), .B(keyinput81), .ZN(n9924) );
  NAND4_X1 U11016 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n9928)
         );
  NOR4_X1 U11017 ( .A1(n9931), .A2(n9930), .A3(n9929), .A4(n9928), .ZN(n10212)
         );
  AOI22_X1 U11018 ( .A1(n9341), .A2(keyinput80), .B1(keyinput68), .B2(n5818), 
        .ZN(n9932) );
  OAI221_X1 U11019 ( .B1(n9341), .B2(keyinput80), .C1(n5818), .C2(keyinput68), 
        .A(n9932), .ZN(n9944) );
  AOI22_X1 U11020 ( .A1(n9935), .A2(keyinput15), .B1(keyinput106), .B2(n9934), 
        .ZN(n9933) );
  OAI221_X1 U11021 ( .B1(n9935), .B2(keyinput15), .C1(n9934), .C2(keyinput106), 
        .A(n9933), .ZN(n9943) );
  AOI22_X1 U11022 ( .A1(n9938), .A2(keyinput65), .B1(keyinput122), .B2(n9937), 
        .ZN(n9936) );
  OAI221_X1 U11023 ( .B1(n9938), .B2(keyinput65), .C1(n9937), .C2(keyinput122), 
        .A(n9936), .ZN(n9942) );
  AOI22_X1 U11024 ( .A1(n6006), .A2(keyinput113), .B1(keyinput46), .B2(n9940), 
        .ZN(n9939) );
  OAI221_X1 U11025 ( .B1(n6006), .B2(keyinput113), .C1(n9940), .C2(keyinput46), 
        .A(n9939), .ZN(n9941) );
  NOR4_X1 U11026 ( .A1(n9944), .A2(n9943), .A3(n9942), .A4(n9941), .ZN(n10024)
         );
  INV_X1 U11027 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9947) );
  AOI22_X1 U11028 ( .A1(n9947), .A2(keyinput59), .B1(n9946), .B2(keyinput75), 
        .ZN(n9945) );
  OAI221_X1 U11029 ( .B1(n9947), .B2(keyinput59), .C1(n9946), .C2(keyinput75), 
        .A(n9945), .ZN(n9958) );
  AOI22_X1 U11030 ( .A1(n5537), .A2(keyinput52), .B1(keyinput21), .B2(n6736), 
        .ZN(n9948) );
  OAI221_X1 U11031 ( .B1(n5537), .B2(keyinput52), .C1(n6736), .C2(keyinput21), 
        .A(n9948), .ZN(n9957) );
  AOI22_X1 U11032 ( .A1(n9951), .A2(keyinput20), .B1(n9950), .B2(keyinput99), 
        .ZN(n9949) );
  OAI221_X1 U11033 ( .B1(n9951), .B2(keyinput20), .C1(n9950), .C2(keyinput99), 
        .A(n9949), .ZN(n9956) );
  INV_X1 U11034 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9954) );
  AOI22_X1 U11035 ( .A1(n9954), .A2(keyinput127), .B1(n9953), .B2(keyinput73), 
        .ZN(n9952) );
  OAI221_X1 U11036 ( .B1(n9954), .B2(keyinput127), .C1(n9953), .C2(keyinput73), 
        .A(n9952), .ZN(n9955) );
  NOR4_X1 U11037 ( .A1(n9958), .A2(n9957), .A3(n9956), .A4(n9955), .ZN(n10023)
         );
  AOI22_X1 U11038 ( .A1(n9961), .A2(keyinput44), .B1(n9960), .B2(keyinput7), 
        .ZN(n9959) );
  OAI221_X1 U11039 ( .B1(n9961), .B2(keyinput44), .C1(n9960), .C2(keyinput7), 
        .A(n9959), .ZN(n9973) );
  INV_X1 U11040 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9963) );
  AOI22_X1 U11041 ( .A1(n6047), .A2(keyinput22), .B1(keyinput107), .B2(n9963), 
        .ZN(n9962) );
  OAI221_X1 U11042 ( .B1(n6047), .B2(keyinput22), .C1(n9963), .C2(keyinput107), 
        .A(n9962), .ZN(n9972) );
  AOI22_X1 U11043 ( .A1(n9966), .A2(keyinput32), .B1(n9965), .B2(keyinput66), 
        .ZN(n9964) );
  OAI221_X1 U11044 ( .B1(n9966), .B2(keyinput32), .C1(n9965), .C2(keyinput66), 
        .A(n9964), .ZN(n9971) );
  INV_X1 U11045 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U11046 ( .A1(n9969), .A2(keyinput50), .B1(keyinput96), .B2(n9968), 
        .ZN(n9967) );
  OAI221_X1 U11047 ( .B1(n9969), .B2(keyinput50), .C1(n9968), .C2(keyinput96), 
        .A(n9967), .ZN(n9970) );
  NOR4_X1 U11048 ( .A1(n9973), .A2(n9972), .A3(n9971), .A4(n9970), .ZN(n10022)
         );
  AOI22_X1 U11049 ( .A1(n9976), .A2(keyinput103), .B1(keyinput39), .B2(n9975), 
        .ZN(n9974) );
  OAI221_X1 U11050 ( .B1(n9976), .B2(keyinput103), .C1(n9975), .C2(keyinput39), 
        .A(n9974), .ZN(n9983) );
  INV_X1 U11051 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U11052 ( .A1(n9979), .A2(keyinput67), .B1(keyinput90), .B2(n9978), 
        .ZN(n9977) );
  OAI221_X1 U11053 ( .B1(n9979), .B2(keyinput67), .C1(n9978), .C2(keyinput90), 
        .A(n9977), .ZN(n9982) );
  XNOR2_X1 U11054 ( .A(n9980), .B(keyinput63), .ZN(n9981) );
  NOR3_X1 U11055 ( .A1(n9983), .A2(n9982), .A3(n9981), .ZN(n10020) );
  INV_X1 U11056 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9986) );
  AOI22_X1 U11057 ( .A1(n9986), .A2(keyinput56), .B1(keyinput6), .B2(n9985), 
        .ZN(n9984) );
  OAI221_X1 U11058 ( .B1(n9986), .B2(keyinput56), .C1(n9985), .C2(keyinput6), 
        .A(n9984), .ZN(n9995) );
  INV_X1 U11059 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9988) );
  AOI22_X1 U11060 ( .A1(n9989), .A2(keyinput17), .B1(keyinput64), .B2(n9988), 
        .ZN(n9987) );
  OAI221_X1 U11061 ( .B1(n9989), .B2(keyinput17), .C1(n9988), .C2(keyinput64), 
        .A(n9987), .ZN(n9994) );
  INV_X1 U11062 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9991) );
  AOI22_X1 U11063 ( .A1(n9992), .A2(keyinput27), .B1(keyinput11), .B2(n9991), 
        .ZN(n9990) );
  OAI221_X1 U11064 ( .B1(n9992), .B2(keyinput27), .C1(n9991), .C2(keyinput11), 
        .A(n9990), .ZN(n9993) );
  NOR3_X1 U11065 ( .A1(n9995), .A2(n9994), .A3(n9993), .ZN(n10019) );
  AOI22_X1 U11066 ( .A1(n7646), .A2(keyinput4), .B1(n9997), .B2(keyinput29), 
        .ZN(n9996) );
  OAI221_X1 U11067 ( .B1(n7646), .B2(keyinput4), .C1(n9997), .C2(keyinput29), 
        .A(n9996), .ZN(n10002) );
  INV_X1 U11068 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n10000) );
  AOI22_X1 U11069 ( .A1(n10000), .A2(keyinput42), .B1(n9999), .B2(keyinput41), 
        .ZN(n9998) );
  OAI221_X1 U11070 ( .B1(n10000), .B2(keyinput42), .C1(n9999), .C2(keyinput41), 
        .A(n9998), .ZN(n10001) );
  NOR2_X1 U11071 ( .A1(n10002), .A2(n10001), .ZN(n10018) );
  INV_X1 U11072 ( .A(keyinput115), .ZN(n10044) );
  NAND2_X1 U11073 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n10044), .ZN(n10004) );
  NAND2_X1 U11074 ( .A1(keyinput115), .A2(n7127), .ZN(n10003) );
  OAI211_X1 U11075 ( .C1(n10005), .C2(keyinput126), .A(n10004), .B(n10003), 
        .ZN(n10006) );
  INV_X1 U11076 ( .A(n10006), .ZN(n10010) );
  XNOR2_X1 U11077 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput94), .ZN(n10009) );
  XNOR2_X1 U11078 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput55), .ZN(n10008) );
  XNOR2_X1 U11079 ( .A(P2_STATE_REG_SCAN_IN), .B(keyinput2), .ZN(n10007) );
  NAND4_X1 U11080 ( .A1(n10010), .A2(n10009), .A3(n10008), .A4(n10007), .ZN(
        n10016) );
  XNOR2_X1 U11081 ( .A(P2_REG1_REG_27__SCAN_IN), .B(keyinput48), .ZN(n10014)
         );
  XNOR2_X1 U11082 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput86), .ZN(n10013) );
  XNOR2_X1 U11083 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput109), .ZN(n10012) );
  XNOR2_X1 U11084 ( .A(keyinput13), .B(SI_30_), .ZN(n10011) );
  NAND4_X1 U11085 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10015) );
  NOR2_X1 U11086 ( .A1(n10016), .A2(n10015), .ZN(n10017) );
  AND4_X1 U11087 ( .A1(n10020), .A2(n10019), .A3(n10018), .A4(n10017), .ZN(
        n10021) );
  AND4_X1 U11088 ( .A1(n10024), .A2(n10023), .A3(n10022), .A4(n10021), .ZN(
        n10211) );
  NOR2_X1 U11089 ( .A1(keyinput75), .A2(keyinput52), .ZN(n10025) );
  NAND3_X1 U11090 ( .A1(keyinput10), .A2(keyinput127), .A3(n10025), .ZN(n10026) );
  NOR3_X1 U11091 ( .A1(keyinput73), .A2(keyinput20), .A3(n10026), .ZN(n10038)
         );
  NAND2_X1 U11092 ( .A1(keyinput42), .A2(keyinput122), .ZN(n10027) );
  NOR3_X1 U11093 ( .A1(keyinput29), .A2(keyinput4), .A3(n10027), .ZN(n10028)
         );
  NAND3_X1 U11094 ( .A1(keyinput41), .A2(keyinput56), .A3(n10028), .ZN(n10036)
         );
  NAND2_X1 U11095 ( .A1(keyinput48), .A2(keyinput27), .ZN(n10029) );
  NOR3_X1 U11096 ( .A1(keyinput64), .A2(keyinput11), .A3(n10029), .ZN(n10034)
         );
  NOR4_X1 U11097 ( .A1(keyinput99), .A2(keyinput17), .A3(keyinput86), .A4(
        keyinput67), .ZN(n10033) );
  NAND2_X1 U11098 ( .A1(keyinput68), .A2(keyinput106), .ZN(n10030) );
  NOR3_X1 U11099 ( .A1(keyinput80), .A2(keyinput113), .A3(n10030), .ZN(n10032)
         );
  NOR4_X1 U11100 ( .A1(keyinput90), .A2(keyinput15), .A3(keyinput46), .A4(
        keyinput65), .ZN(n10031) );
  NAND4_X1 U11101 ( .A1(n10034), .A2(n10033), .A3(n10032), .A4(n10031), .ZN(
        n10035) );
  NOR4_X1 U11102 ( .A1(keyinput6), .A2(keyinput109), .A3(n10036), .A4(n10035), 
        .ZN(n10037) );
  NAND4_X1 U11103 ( .A1(keyinput21), .A2(keyinput59), .A3(n10038), .A4(n10037), 
        .ZN(n10087) );
  NAND2_X1 U11104 ( .A1(keyinput36), .A2(keyinput30), .ZN(n10039) );
  NOR3_X1 U11105 ( .A1(keyinput1), .A2(keyinput62), .A3(n10039), .ZN(n10085)
         );
  NOR4_X1 U11106 ( .A1(keyinput43), .A2(keyinput8), .A3(keyinput19), .A4(
        keyinput57), .ZN(n10084) );
  INV_X1 U11107 ( .A(keyinput78), .ZN(n10040) );
  NOR4_X1 U11108 ( .A1(keyinput91), .A2(keyinput34), .A3(keyinput12), .A4(
        n10040), .ZN(n10041) );
  NAND3_X1 U11109 ( .A1(keyinput66), .A2(keyinput81), .A3(n10041), .ZN(n10049)
         );
  INV_X1 U11110 ( .A(keyinput63), .ZN(n10042) );
  NAND4_X1 U11111 ( .A1(keyinput55), .A2(keyinput2), .A3(keyinput103), .A4(
        n10042), .ZN(n10043) );
  NOR4_X1 U11112 ( .A1(keyinput58), .A2(keyinput94), .A3(n10044), .A4(n10043), 
        .ZN(n10047) );
  NAND4_X1 U11113 ( .A1(keyinput107), .A2(keyinput44), .A3(keyinput96), .A4(
        keyinput32), .ZN(n10045) );
  NOR3_X1 U11114 ( .A1(keyinput7), .A2(keyinput50), .A3(n10045), .ZN(n10046)
         );
  NAND4_X1 U11115 ( .A1(n10047), .A2(keyinput39), .A3(keyinput22), .A4(n10046), 
        .ZN(n10048) );
  NOR4_X1 U11116 ( .A1(keyinput121), .A2(keyinput54), .A3(n10049), .A4(n10048), 
        .ZN(n10083) );
  NOR2_X1 U11117 ( .A1(keyinput13), .A2(keyinput102), .ZN(n10050) );
  NAND3_X1 U11118 ( .A1(keyinput123), .A2(keyinput38), .A3(n10050), .ZN(n10051) );
  NOR3_X1 U11119 ( .A1(keyinput110), .A2(keyinput60), .A3(n10051), .ZN(n10065)
         );
  NAND2_X1 U11120 ( .A1(keyinput40), .A2(keyinput95), .ZN(n10052) );
  NOR3_X1 U11121 ( .A1(keyinput61), .A2(keyinput26), .A3(n10052), .ZN(n10053)
         );
  NAND3_X1 U11122 ( .A1(keyinput70), .A2(keyinput74), .A3(n10053), .ZN(n10063)
         );
  INV_X1 U11123 ( .A(keyinput76), .ZN(n10054) );
  NOR4_X1 U11124 ( .A1(keyinput35), .A2(keyinput31), .A3(keyinput116), .A4(
        n10054), .ZN(n10061) );
  NAND2_X1 U11125 ( .A1(keyinput49), .A2(keyinput14), .ZN(n10055) );
  NOR3_X1 U11126 ( .A1(keyinput28), .A2(keyinput79), .A3(n10055), .ZN(n10060)
         );
  INV_X1 U11127 ( .A(keyinput72), .ZN(n10056) );
  NOR4_X1 U11128 ( .A1(keyinput47), .A2(keyinput105), .A3(keyinput125), .A4(
        n10056), .ZN(n10059) );
  NAND2_X1 U11129 ( .A1(keyinput87), .A2(keyinput82), .ZN(n10057) );
  NOR3_X1 U11130 ( .A1(keyinput119), .A2(keyinput88), .A3(n10057), .ZN(n10058)
         );
  NAND4_X1 U11131 ( .A1(n10061), .A2(n10060), .A3(n10059), .A4(n10058), .ZN(
        n10062) );
  NOR4_X1 U11132 ( .A1(keyinput37), .A2(keyinput114), .A3(n10063), .A4(n10062), 
        .ZN(n10064) );
  NAND4_X1 U11133 ( .A1(keyinput45), .A2(keyinput24), .A3(n10065), .A4(n10064), 
        .ZN(n10081) );
  NAND4_X1 U11134 ( .A1(keyinput111), .A2(keyinput118), .A3(keyinput53), .A4(
        keyinput93), .ZN(n10080) );
  NOR2_X1 U11135 ( .A1(keyinput83), .A2(keyinput98), .ZN(n10066) );
  NAND3_X1 U11136 ( .A1(keyinput97), .A2(keyinput104), .A3(n10066), .ZN(n10079) );
  NOR2_X1 U11137 ( .A1(keyinput3), .A2(keyinput85), .ZN(n10067) );
  NAND3_X1 U11138 ( .A1(keyinput77), .A2(keyinput112), .A3(n10067), .ZN(n10068) );
  NOR3_X1 U11139 ( .A1(keyinput5), .A2(keyinput92), .A3(n10068), .ZN(n10077)
         );
  NAND4_X1 U11140 ( .A1(keyinput120), .A2(keyinput100), .A3(keyinput89), .A4(
        keyinput71), .ZN(n10075) );
  NOR2_X1 U11141 ( .A1(keyinput0), .A2(keyinput33), .ZN(n10069) );
  NAND3_X1 U11142 ( .A1(keyinput18), .A2(keyinput23), .A3(n10069), .ZN(n10074)
         );
  NOR2_X1 U11143 ( .A1(keyinput69), .A2(keyinput117), .ZN(n10070) );
  NAND3_X1 U11144 ( .A1(keyinput51), .A2(keyinput16), .A3(n10070), .ZN(n10073)
         );
  INV_X1 U11145 ( .A(keyinput101), .ZN(n10071) );
  NAND4_X1 U11146 ( .A1(keyinput25), .A2(keyinput84), .A3(keyinput108), .A4(
        n10071), .ZN(n10072) );
  NOR4_X1 U11147 ( .A1(n10075), .A2(n10074), .A3(n10073), .A4(n10072), .ZN(
        n10076) );
  NAND4_X1 U11148 ( .A1(keyinput124), .A2(keyinput9), .A3(n10077), .A4(n10076), 
        .ZN(n10078) );
  NOR4_X1 U11149 ( .A1(n10081), .A2(n10080), .A3(n10079), .A4(n10078), .ZN(
        n10082) );
  NAND4_X1 U11150 ( .A1(n10085), .A2(n10084), .A3(n10083), .A4(n10082), .ZN(
        n10086) );
  OAI21_X1 U11151 ( .B1(n10087), .B2(n10086), .A(P1_IR_REG_16__SCAN_IN), .ZN(
        n10209) );
  AOI22_X1 U11152 ( .A1(n8574), .A2(keyinput123), .B1(n6218), .B2(keyinput102), 
        .ZN(n10088) );
  OAI221_X1 U11153 ( .B1(n8574), .B2(keyinput123), .C1(n6218), .C2(keyinput102), .A(n10088), .ZN(n10100) );
  AOI22_X1 U11154 ( .A1(n10091), .A2(keyinput38), .B1(n10090), .B2(keyinput45), 
        .ZN(n10089) );
  OAI221_X1 U11155 ( .B1(n10091), .B2(keyinput38), .C1(n10090), .C2(keyinput45), .A(n10089), .ZN(n10099) );
  AOI22_X1 U11156 ( .A1(n10094), .A2(keyinput24), .B1(n10093), .B2(keyinput110), .ZN(n10092) );
  OAI221_X1 U11157 ( .B1(n10094), .B2(keyinput24), .C1(n10093), .C2(
        keyinput110), .A(n10092), .ZN(n10098) );
  AOI22_X1 U11158 ( .A1(n6445), .A2(keyinput60), .B1(n10096), .B2(keyinput28), 
        .ZN(n10095) );
  OAI221_X1 U11159 ( .B1(n6445), .B2(keyinput60), .C1(n10096), .C2(keyinput28), 
        .A(n10095), .ZN(n10097) );
  NOR4_X1 U11160 ( .A1(n10100), .A2(n10099), .A3(n10098), .A4(n10097), .ZN(
        n10144) );
  AOI22_X1 U11161 ( .A1(n5836), .A2(keyinput14), .B1(n10102), .B2(keyinput49), 
        .ZN(n10101) );
  OAI221_X1 U11162 ( .B1(n5836), .B2(keyinput14), .C1(n10102), .C2(keyinput49), 
        .A(n10101), .ZN(n10112) );
  AOI22_X1 U11163 ( .A1(n10105), .A2(keyinput79), .B1(n10104), .B2(keyinput35), 
        .ZN(n10103) );
  OAI221_X1 U11164 ( .B1(n10105), .B2(keyinput79), .C1(n10104), .C2(keyinput35), .A(n10103), .ZN(n10111) );
  XOR2_X1 U11165 ( .A(n6284), .B(keyinput31), .Z(n10109) );
  XOR2_X1 U11166 ( .A(n6765), .B(keyinput82), .Z(n10108) );
  XNOR2_X1 U11167 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput116), .ZN(n10107) );
  XNOR2_X1 U11168 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput76), .ZN(n10106) );
  NAND4_X1 U11169 ( .A1(n10109), .A2(n10108), .A3(n10107), .A4(n10106), .ZN(
        n10110) );
  NOR3_X1 U11170 ( .A1(n10112), .A2(n10111), .A3(n10110), .ZN(n10143) );
  AOI22_X1 U11171 ( .A1(n10114), .A2(keyinput105), .B1(keyinput125), .B2(n7764), .ZN(n10113) );
  OAI221_X1 U11172 ( .B1(n10114), .B2(keyinput105), .C1(n7764), .C2(
        keyinput125), .A(n10113), .ZN(n10125) );
  AOI22_X1 U11173 ( .A1(n10116), .A2(keyinput87), .B1(n6345), .B2(keyinput47), 
        .ZN(n10115) );
  OAI221_X1 U11174 ( .B1(n10116), .B2(keyinput87), .C1(n6345), .C2(keyinput47), 
        .A(n10115), .ZN(n10124) );
  AOI22_X1 U11175 ( .A1(n10119), .A2(keyinput88), .B1(n10118), .B2(keyinput119), .ZN(n10117) );
  OAI221_X1 U11176 ( .B1(n10119), .B2(keyinput88), .C1(n10118), .C2(
        keyinput119), .A(n10117), .ZN(n10123) );
  XOR2_X1 U11177 ( .A(n7428), .B(keyinput72), .Z(n10121) );
  XNOR2_X1 U11178 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput70), .ZN(n10120)
         );
  NAND2_X1 U11179 ( .A1(n10121), .A2(n10120), .ZN(n10122) );
  NOR4_X1 U11180 ( .A1(n10125), .A2(n10124), .A3(n10123), .A4(n10122), .ZN(
        n10142) );
  AOI22_X1 U11181 ( .A1(n10128), .A2(keyinput74), .B1(n10127), .B2(keyinput95), 
        .ZN(n10126) );
  OAI221_X1 U11182 ( .B1(n10128), .B2(keyinput74), .C1(n10127), .C2(keyinput95), .A(n10126), .ZN(n10140) );
  AOI22_X1 U11183 ( .A1(n4616), .A2(keyinput26), .B1(keyinput61), .B2(n10130), 
        .ZN(n10129) );
  OAI221_X1 U11184 ( .B1(n4616), .B2(keyinput26), .C1(n10130), .C2(keyinput61), 
        .A(n10129), .ZN(n10139) );
  INV_X1 U11185 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U11186 ( .A1(n10133), .A2(keyinput40), .B1(n10132), .B2(keyinput37), 
        .ZN(n10131) );
  OAI221_X1 U11187 ( .B1(n10133), .B2(keyinput40), .C1(n10132), .C2(keyinput37), .A(n10131), .ZN(n10138) );
  INV_X1 U11188 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n10136) );
  INV_X1 U11189 ( .A(SI_7_), .ZN(n10135) );
  AOI22_X1 U11190 ( .A1(n10136), .A2(keyinput114), .B1(n10135), .B2(keyinput97), .ZN(n10134) );
  OAI221_X1 U11191 ( .B1(n10136), .B2(keyinput114), .C1(n10135), .C2(
        keyinput97), .A(n10134), .ZN(n10137) );
  NOR4_X1 U11192 ( .A1(n10140), .A2(n10139), .A3(n10138), .A4(n10137), .ZN(
        n10141) );
  NAND4_X1 U11193 ( .A1(n10144), .A2(n10143), .A3(n10142), .A4(n10141), .ZN(
        n10208) );
  INV_X1 U11194 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U11195 ( .A1(n10146), .A2(keyinput98), .B1(keyinput83), .B2(n6212), 
        .ZN(n10145) );
  OAI221_X1 U11196 ( .B1(n10146), .B2(keyinput98), .C1(n6212), .C2(keyinput83), 
        .A(n10145), .ZN(n10157) );
  AOI22_X1 U11197 ( .A1(n10149), .A2(keyinput104), .B1(n10148), .B2(
        keyinput111), .ZN(n10147) );
  OAI221_X1 U11198 ( .B1(n10149), .B2(keyinput104), .C1(n10148), .C2(
        keyinput111), .A(n10147), .ZN(n10156) );
  AOI22_X1 U11199 ( .A1(n6042), .A2(keyinput118), .B1(keyinput53), .B2(n6582), 
        .ZN(n10150) );
  OAI221_X1 U11200 ( .B1(n6042), .B2(keyinput118), .C1(n6582), .C2(keyinput53), 
        .A(n10150), .ZN(n10155) );
  AOI22_X1 U11201 ( .A1(n10153), .A2(keyinput93), .B1(n10152), .B2(keyinput18), 
        .ZN(n10151) );
  OAI221_X1 U11202 ( .B1(n10153), .B2(keyinput93), .C1(n10152), .C2(keyinput18), .A(n10151), .ZN(n10154) );
  NOR4_X1 U11203 ( .A1(n10157), .A2(n10156), .A3(n10155), .A4(n10154), .ZN(
        n10206) );
  AOI22_X1 U11204 ( .A1(n10160), .A2(keyinput33), .B1(n10159), .B2(keyinput89), 
        .ZN(n10158) );
  OAI221_X1 U11205 ( .B1(n10160), .B2(keyinput33), .C1(n10159), .C2(keyinput89), .A(n10158), .ZN(n10161) );
  INV_X1 U11206 ( .A(n10161), .ZN(n10176) );
  AOI22_X1 U11207 ( .A1(n10164), .A2(keyinput100), .B1(n10163), .B2(keyinput23), .ZN(n10162) );
  OAI221_X1 U11208 ( .B1(n10164), .B2(keyinput100), .C1(n10163), .C2(
        keyinput23), .A(n10162), .ZN(n10167) );
  INV_X1 U11209 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n10165) );
  XNOR2_X1 U11210 ( .A(n10165), .B(keyinput120), .ZN(n10166) );
  NOR2_X1 U11211 ( .A1(n10167), .A2(n10166), .ZN(n10175) );
  INV_X1 U11212 ( .A(keyinput0), .ZN(n10168) );
  XNOR2_X1 U11213 ( .A(n10169), .B(n10168), .ZN(n10174) );
  AOI22_X1 U11214 ( .A1(n9058), .A2(keyinput71), .B1(n10171), .B2(keyinput3), 
        .ZN(n10170) );
  OAI221_X1 U11215 ( .B1(n9058), .B2(keyinput71), .C1(n10171), .C2(keyinput3), 
        .A(n10170), .ZN(n10172) );
  INV_X1 U11216 ( .A(n10172), .ZN(n10173) );
  AND4_X1 U11217 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10205) );
  AOI22_X1 U11218 ( .A1(n10178), .A2(keyinput77), .B1(n6323), .B2(keyinput124), 
        .ZN(n10177) );
  OAI221_X1 U11219 ( .B1(n10178), .B2(keyinput77), .C1(n6323), .C2(keyinput124), .A(n10177), .ZN(n10190) );
  AOI22_X1 U11220 ( .A1(n10181), .A2(keyinput9), .B1(keyinput5), .B2(n10180), 
        .ZN(n10179) );
  OAI221_X1 U11221 ( .B1(n10181), .B2(keyinput9), .C1(n10180), .C2(keyinput5), 
        .A(n10179), .ZN(n10189) );
  AOI22_X1 U11222 ( .A1(n6468), .A2(keyinput92), .B1(n10183), .B2(keyinput85), 
        .ZN(n10182) );
  OAI221_X1 U11223 ( .B1(n6468), .B2(keyinput92), .C1(n10183), .C2(keyinput85), 
        .A(n10182), .ZN(n10188) );
  AOI22_X1 U11224 ( .A1(n10186), .A2(keyinput112), .B1(n10185), .B2(keyinput25), .ZN(n10184) );
  OAI221_X1 U11225 ( .B1(n10186), .B2(keyinput112), .C1(n10185), .C2(
        keyinput25), .A(n10184), .ZN(n10187) );
  NOR4_X1 U11226 ( .A1(n10190), .A2(n10189), .A3(n10188), .A4(n10187), .ZN(
        n10204) );
  AOI22_X1 U11227 ( .A1(n5033), .A2(keyinput101), .B1(keyinput84), .B2(n5134), 
        .ZN(n10191) );
  OAI221_X1 U11228 ( .B1(n5033), .B2(keyinput101), .C1(n5134), .C2(keyinput84), 
        .A(n10191), .ZN(n10202) );
  INV_X1 U11229 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U11230 ( .A1(n10194), .A2(keyinput108), .B1(n10193), .B2(keyinput51), .ZN(n10192) );
  OAI221_X1 U11231 ( .B1(n10194), .B2(keyinput108), .C1(n10193), .C2(
        keyinput51), .A(n10192), .ZN(n10201) );
  AOI22_X1 U11232 ( .A1(n10196), .A2(keyinput69), .B1(P1_U3084), .B2(
        keyinput16), .ZN(n10195) );
  OAI221_X1 U11233 ( .B1(n10196), .B2(keyinput69), .C1(P1_U3084), .C2(
        keyinput16), .A(n10195), .ZN(n10200) );
  AOI22_X1 U11234 ( .A1(n4618), .A2(keyinput58), .B1(n10198), .B2(keyinput117), 
        .ZN(n10197) );
  OAI221_X1 U11235 ( .B1(n4618), .B2(keyinput58), .C1(n10198), .C2(keyinput117), .A(n10197), .ZN(n10199) );
  NOR4_X1 U11236 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10203) );
  NAND4_X1 U11237 ( .A1(n10206), .A2(n10205), .A3(n10204), .A4(n10203), .ZN(
        n10207) );
  AOI211_X1 U11238 ( .C1(keyinput126), .C2(n10209), .A(n10208), .B(n10207), 
        .ZN(n10210) );
  NAND4_X1 U11239 ( .A1(n10213), .A2(n10212), .A3(n10211), .A4(n10210), .ZN(
        n10216) );
  MUX2_X1 U11240 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n10214), .S(P1_U4006), .Z(
        n10215) );
  XNOR2_X1 U11241 ( .A(n10216), .B(n10215), .ZN(P1_U3570) );
  XNOR2_X1 U11242 ( .A(n10217), .B(n6582), .ZN(ADD_1071_U50) );
  NOR2_X1 U11243 ( .A1(n10219), .A2(n10218), .ZN(n10220) );
  XNOR2_X1 U11244 ( .A(n10220), .B(n9569), .ZN(ADD_1071_U51) );
  OAI21_X1 U11245 ( .B1(n10223), .B2(n10222), .A(n10221), .ZN(n10224) );
  XNOR2_X1 U11246 ( .A(n10224), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11247 ( .B1(n10227), .B2(n10226), .A(n10225), .ZN(ADD_1071_U47) );
  XOR2_X1 U11248 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10228), .Z(ADD_1071_U48) );
  XOR2_X1 U11249 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10229), .Z(ADD_1071_U49) );
  XOR2_X1 U11250 ( .A(n10231), .B(n10230), .Z(ADD_1071_U54) );
  XOR2_X1 U11251 ( .A(n10233), .B(n10232), .Z(ADD_1071_U53) );
  XNOR2_X1 U11252 ( .A(n10235), .B(n10234), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4907 ( .A(n7521), .Z(n7991) );
  AND3_X1 U4923 ( .A1(n5845), .A2(n5844), .A3(n5843), .ZN(n9779) );
  CLKBUF_X1 U5062 ( .A(n5411), .Z(n5558) );
  CLKBUF_X2 U5063 ( .A(n5765), .Z(n4391) );
endmodule

