

module b15_C_AntiSAT_k_256_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        keyinput128, keyinput129, keyinput130, keyinput131, keyinput132, 
        keyinput133, keyinput134, keyinput135, keyinput136, keyinput137, 
        keyinput138, keyinput139, keyinput140, keyinput141, keyinput142, 
        keyinput143, keyinput144, keyinput145, keyinput146, keyinput147, 
        keyinput148, keyinput149, keyinput150, keyinput151, keyinput152, 
        keyinput153, keyinput154, keyinput155, keyinput156, keyinput157, 
        keyinput158, keyinput159, keyinput160, keyinput161, keyinput162, 
        keyinput163, keyinput164, keyinput165, keyinput166, keyinput167, 
        keyinput168, keyinput169, keyinput170, keyinput171, keyinput172, 
        keyinput173, keyinput174, keyinput175, keyinput176, keyinput177, 
        keyinput178, keyinput179, keyinput180, keyinput181, keyinput182, 
        keyinput183, keyinput184, keyinput185, keyinput186, keyinput187, 
        keyinput188, keyinput189, keyinput190, keyinput191, keyinput192, 
        keyinput193, keyinput194, keyinput195, keyinput196, keyinput197, 
        keyinput198, keyinput199, keyinput200, keyinput201, keyinput202, 
        keyinput203, keyinput204, keyinput205, keyinput206, keyinput207, 
        keyinput208, keyinput209, keyinput210, keyinput211, keyinput212, 
        keyinput213, keyinput214, keyinput215, keyinput216, keyinput217, 
        keyinput218, keyinput219, keyinput220, keyinput221, keyinput222, 
        keyinput223, keyinput224, keyinput225, keyinput226, keyinput227, 
        keyinput228, keyinput229, keyinput230, keyinput231, keyinput232, 
        keyinput233, keyinput234, keyinput235, keyinput236, keyinput237, 
        keyinput238, keyinput239, keyinput240, keyinput241, keyinput242, 
        keyinput243, keyinput244, keyinput245, keyinput246, keyinput247, 
        keyinput248, keyinput249, keyinput250, keyinput251, keyinput252, 
        keyinput253, keyinput254, keyinput255, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127, keyinput128,
         keyinput129, keyinput130, keyinput131, keyinput132, keyinput133,
         keyinput134, keyinput135, keyinput136, keyinput137, keyinput138,
         keyinput139, keyinput140, keyinput141, keyinput142, keyinput143,
         keyinput144, keyinput145, keyinput146, keyinput147, keyinput148,
         keyinput149, keyinput150, keyinput151, keyinput152, keyinput153,
         keyinput154, keyinput155, keyinput156, keyinput157, keyinput158,
         keyinput159, keyinput160, keyinput161, keyinput162, keyinput163,
         keyinput164, keyinput165, keyinput166, keyinput167, keyinput168,
         keyinput169, keyinput170, keyinput171, keyinput172, keyinput173,
         keyinput174, keyinput175, keyinput176, keyinput177, keyinput178,
         keyinput179, keyinput180, keyinput181, keyinput182, keyinput183,
         keyinput184, keyinput185, keyinput186, keyinput187, keyinput188,
         keyinput189, keyinput190, keyinput191, keyinput192, keyinput193,
         keyinput194, keyinput195, keyinput196, keyinput197, keyinput198,
         keyinput199, keyinput200, keyinput201, keyinput202, keyinput203,
         keyinput204, keyinput205, keyinput206, keyinput207, keyinput208,
         keyinput209, keyinput210, keyinput211, keyinput212, keyinput213,
         keyinput214, keyinput215, keyinput216, keyinput217, keyinput218,
         keyinput219, keyinput220, keyinput221, keyinput222, keyinput223,
         keyinput224, keyinput225, keyinput226, keyinput227, keyinput228,
         keyinput229, keyinput230, keyinput231, keyinput232, keyinput233,
         keyinput234, keyinput235, keyinput236, keyinput237, keyinput238,
         keyinput239, keyinput240, keyinput241, keyinput242, keyinput243,
         keyinput244, keyinput245, keyinput246, keyinput247, keyinput248,
         keyinput249, keyinput250, keyinput251, keyinput252, keyinput253,
         keyinput254, keyinput255;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150;

  NAND2_X1 U3619 ( .A1(n5570), .A2(n5572), .ZN(n5571) );
  AND2_X1 U3620 ( .A1(n3761), .A2(n3760), .ZN(n4612) );
  CLKBUF_X2 U3621 ( .A(n3429), .Z(n4099) );
  CLKBUF_X1 U3622 ( .A(n3589), .Z(n3841) );
  CLKBUF_X2 U3623 ( .A(n3428), .Z(n4271) );
  CLKBUF_X1 U3624 ( .A(n3407), .Z(n4864) );
  AND4_X1 U3625 ( .A1(n3319), .A2(n3318), .A3(n3317), .A4(n3316), .ZN(n3341)
         );
  CLKBUF_X2 U3626 ( .A(n3427), .Z(n4264) );
  AND4_X1 U3627 ( .A1(n3327), .A2(n3326), .A3(n3325), .A4(n3324), .ZN(n3340)
         );
  INV_X1 U3628 ( .A(n3728), .ZN(n3749) );
  NOR2_X1 U3629 ( .A1(n5370), .A2(n5369), .ZN(n5408) );
  INV_X1 U3630 ( .A(n4857), .ZN(n4845) );
  NAND2_X1 U3631 ( .A1(n4461), .A2(n4462), .ZN(n4430) );
  INV_X1 U3632 ( .A(n6207), .ZN(n6188) );
  OR2_X1 U3633 ( .A1(n5459), .A2(n6292), .ZN(n4298) );
  AND2_X2 U3634 ( .A1(n4486), .A2(n3886), .ZN(n4461) );
  INV_X2 U3635 ( .A(n3240), .ZN(n5526) );
  AND2_X4 U3636 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4530) );
  AOI21_X2 U3637 ( .B1(n5715), .B2(n5707), .A(n5714), .ZN(n5858) );
  AND2_X4 U3638 ( .A1(n3406), .A2(n3475), .ZN(n5662) );
  OR2_X4 U3639 ( .A1(n3353), .A2(n3352), .ZN(n3475) );
  OR2_X1 U3640 ( .A1(n3210), .A2(n5728), .ZN(n5721) );
  INV_X4 U3641 ( .A(n6271), .ZN(n3171) );
  NAND2_X1 U3642 ( .A1(n3599), .A2(n3598), .ZN(n3629) );
  NAND2_X1 U3644 ( .A1(n6221), .A2(n5460), .ZN(n5678) );
  CLKBUF_X2 U3645 ( .A(n4371), .Z(n4417) );
  NAND2_X1 U3646 ( .A1(n3223), .A2(n3471), .ZN(n3533) );
  NAND3_X1 U3647 ( .A1(n3479), .A2(n3195), .A3(n3481), .ZN(n4615) );
  NAND2_X1 U3648 ( .A1(n3311), .A2(n3310), .ZN(n3763) );
  INV_X2 U3649 ( .A(n4434), .ZN(n5473) );
  AND2_X1 U3650 ( .A1(n4424), .A2(n4864), .ZN(n3195) );
  BUF_X2 U3651 ( .A(n3391), .Z(n4270) );
  CLKBUF_X2 U3652 ( .A(n3451), .Z(n4272) );
  NAND2_X1 U3653 ( .A1(n4243), .A2(n6530), .ZN(n6292) );
  BUF_X2 U3654 ( .A(n3612), .Z(n4263) );
  AND2_X1 U3655 ( .A1(n3730), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3273)
         );
  AND2_X2 U3656 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4520) );
  AOI21_X1 U3657 ( .B1(n5749), .B2(n5889), .A(n3242), .ZN(n5743) );
  INV_X1 U3658 ( .A(n5684), .ZN(n5705) );
  AND2_X2 U3659 ( .A1(n5428), .A2(n5429), .ZN(n5403) );
  NAND2_X1 U3660 ( .A1(n4014), .A2(n4013), .ZN(n4029) );
  AOI21_X1 U3661 ( .B1(n3198), .B2(n3200), .A(n3180), .ZN(n3197) );
  OAI21_X1 U3662 ( .B1(n3251), .B2(n3194), .A(n3171), .ZN(n3247) );
  XNOR2_X1 U3663 ( .A(n3692), .B(n3681), .ZN(n3930) );
  NAND2_X2 U3664 ( .A1(n3692), .A2(n3691), .ZN(n6271) );
  NAND2_X1 U3665 ( .A1(n3669), .A2(n3668), .ZN(n3692) );
  AOI21_X1 U3666 ( .B1(n3894), .B2(n4043), .A(n3905), .ZN(n4431) );
  OAI211_X1 U3667 ( .C1(n3887), .C2(n4059), .A(n3893), .B(n3892), .ZN(n4462)
         );
  AOI21_X1 U3668 ( .B1(n4522), .B2(n6743), .A(n3597), .ZN(n4587) );
  AND2_X1 U3669 ( .A1(n3531), .A2(n3530), .ZN(n3560) );
  OAI21_X1 U3670 ( .B1(n4819), .B2(n3728), .A(n3467), .ZN(n4357) );
  AND2_X1 U3671 ( .A1(n3513), .A2(n3512), .ZN(n3524) );
  NAND2_X1 U3672 ( .A1(n3241), .A2(n3503), .ZN(n3526) );
  NAND2_X1 U3673 ( .A1(n4838), .A2(n4837), .ZN(n5326) );
  CLKBUF_X1 U3674 ( .A(n3874), .Z(n6597) );
  XNOR2_X1 U3675 ( .A(n3533), .B(n3532), .ZN(n4664) );
  NAND2_X1 U3676 ( .A1(n3582), .A2(n3581), .ZN(n4975) );
  NAND2_X1 U3677 ( .A1(n3259), .A2(n3423), .ZN(n4326) );
  AND3_X1 U3678 ( .A1(n3263), .A2(n3420), .A3(n4327), .ZN(n3424) );
  OAI211_X1 U3679 ( .C1(n4313), .C2(n3483), .A(n4615), .B(n4524), .ZN(n3484)
         );
  CLKBUF_X1 U3680 ( .A(n4524), .Z(n6081) );
  AND2_X1 U3681 ( .A1(n3403), .A2(n4527), .ZN(n4327) );
  NOR2_X1 U3682 ( .A1(n3461), .A2(n6743), .ZN(n3690) );
  OR2_X1 U3683 ( .A1(n3507), .A2(n3584), .ZN(n3503) );
  INV_X2 U3684 ( .A(n4854), .ZN(n6739) );
  NAND2_X1 U3685 ( .A1(n4873), .A2(n4857), .ZN(n4839) );
  NAND2_X1 U3686 ( .A1(n3764), .A2(n4603), .ZN(n3728) );
  OR2_X2 U3687 ( .A1(n4857), .A2(n3406), .ZN(n4854) );
  AND2_X1 U3689 ( .A1(n3860), .A2(n3764), .ZN(n3417) );
  OR2_X1 U3690 ( .A1(n3457), .A2(n3456), .ZN(n3693) );
  OR2_X1 U3691 ( .A1(n3406), .A2(n3192), .ZN(n3478) );
  OR2_X1 U3692 ( .A1(n3441), .A2(n3440), .ZN(n3565) );
  INV_X1 U3693 ( .A(n4880), .ZN(n4607) );
  NAND4_X2 U3694 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(n3406)
         );
  AND2_X1 U3695 ( .A1(n4673), .A2(n3400), .ZN(n3401) );
  AND2_X2 U3696 ( .A1(n3337), .A2(n3336), .ZN(n4880) );
  AND4_X1 U3697 ( .A1(n3359), .A2(n3358), .A3(n3357), .A4(n3356), .ZN(n3375)
         );
  AND4_X1 U3698 ( .A1(n3343), .A2(n3341), .A3(n3342), .A4(n3340), .ZN(n3407)
         );
  NAND4_X2 U3699 ( .A1(n3343), .A2(n3342), .A3(n3341), .A4(n3340), .ZN(n3764)
         );
  AND4_X1 U3700 ( .A1(n3283), .A2(n3282), .A3(n3281), .A4(n3280), .ZN(n3289)
         );
  AND4_X1 U3701 ( .A1(n3386), .A2(n3385), .A3(n3384), .A4(n3383), .ZN(n3398)
         );
  AND4_X1 U3702 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3288)
         );
  AND4_X1 U3703 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(n3399)
         );
  AND4_X1 U3704 ( .A1(n3297), .A2(n3296), .A3(n3295), .A4(n3294), .ZN(n3308)
         );
  AND4_X1 U3705 ( .A1(n3367), .A2(n3366), .A3(n3365), .A4(n3364), .ZN(n3373)
         );
  AND4_X1 U3706 ( .A1(n3293), .A2(n3292), .A3(n3291), .A4(n3290), .ZN(n3309)
         );
  AND4_X1 U3707 ( .A1(n3301), .A2(n3300), .A3(n3299), .A4(n3298), .ZN(n3307)
         );
  AND4_X1 U3708 ( .A1(n3363), .A2(n3362), .A3(n3361), .A4(n3360), .ZN(n3374)
         );
  AND4_X1 U3709 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3278)
         );
  AND4_X1 U3710 ( .A1(n3305), .A2(n3304), .A3(n3303), .A4(n3302), .ZN(n3306)
         );
  AND4_X1 U3711 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3396)
         );
  AND4_X1 U3712 ( .A1(n3271), .A2(n3270), .A3(n3269), .A4(n3268), .ZN(n3279)
         );
  AND4_X1 U3713 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3397)
         );
  AND4_X1 U3714 ( .A1(n3323), .A2(n3322), .A3(n3321), .A4(n3320), .ZN(n3342)
         );
  AND4_X1 U3715 ( .A1(n3315), .A2(n3314), .A3(n3313), .A4(n3312), .ZN(n3343)
         );
  AND4_X1 U3716 ( .A1(n3335), .A2(n3334), .A3(n3333), .A4(n3332), .ZN(n3336)
         );
  AND4_X1 U3717 ( .A1(n3331), .A2(n3330), .A3(n3329), .A4(n3328), .ZN(n3337)
         );
  BUF_X2 U3718 ( .A(n3444), .Z(n4262) );
  CLKBUF_X2 U3719 ( .A(n3378), .Z(n3428) );
  AOI22_X1 U3720 ( .A1(n3496), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3451), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3269) );
  BUF_X2 U3721 ( .A(n3549), .Z(n4273) );
  BUF_X2 U3722 ( .A(n3377), .Z(n4261) );
  BUF_X2 U3723 ( .A(n3496), .Z(n3443) );
  AND2_X2 U3724 ( .A1(n4535), .A2(n5444), .ZN(n3496) );
  AND2_X2 U3725 ( .A1(n5444), .A2(n4520), .ZN(n3451) );
  AND2_X2 U3726 ( .A1(n4520), .A2(n3273), .ZN(n3612) );
  AND2_X2 U3727 ( .A1(n5444), .A2(n4531), .ZN(n3427) );
  AND2_X2 U3728 ( .A1(n5444), .A2(n3272), .ZN(n3444) );
  AND2_X2 U3729 ( .A1(n3273), .A2(n4535), .ZN(n3549) );
  AND2_X2 U3730 ( .A1(n3273), .A2(n4531), .ZN(n3378) );
  AND2_X2 U3731 ( .A1(n6743), .A2(n4591), .ZN(n6747) );
  CLKBUF_X1 U3732 ( .A(n6486), .Z(n6530) );
  AND2_X2 U3733 ( .A1(n4558), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4535)
         );
  AND2_X2 U3734 ( .A1(n4534), .A2(n3267), .ZN(n3589) );
  AND2_X2 U3735 ( .A1(n3266), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5444)
         );
  INV_X2 U3736 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4558) );
  INV_X2 U3737 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4521) );
  AND2_X1 U3738 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4534) );
  INV_X1 U3739 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5452) );
  INV_X2 U3740 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6743) );
  NAND2_X2 U3741 ( .A1(n3923), .A2(n3922), .ZN(n4655) );
  AND2_X2 U3742 ( .A1(n4740), .A2(n3226), .ZN(n5229) );
  NOR2_X4 U3743 ( .A1(n4655), .A2(n4654), .ZN(n4740) );
  AND2_X2 U3744 ( .A1(n4530), .A2(n4531), .ZN(n4265) );
  NAND2_X2 U3745 ( .A1(n3629), .A2(n3601), .ZN(n3887) );
  AND2_X2 U3746 ( .A1(n4520), .A2(n4581), .ZN(n3429) );
  AND2_X2 U3747 ( .A1(n3272), .A2(n4581), .ZN(n3391) );
  AND2_X2 U3748 ( .A1(n4535), .A2(n4581), .ZN(n3377) );
  NOR3_X4 U3749 ( .A1(n5731), .A2(n5728), .A3(n3713), .ZN(n5709) );
  AND2_X2 U3750 ( .A1(n3210), .A2(n3188), .ZN(n5731) );
  XNOR2_X1 U3751 ( .A(n4572), .B(n4975), .ZN(n4522) );
  AND2_X2 U3752 ( .A1(n5599), .A2(n5648), .ZN(n5587) );
  NOR2_X2 U3753 ( .A1(n5600), .A2(n5601), .ZN(n5599) );
  NAND2_X2 U3754 ( .A1(n3563), .A2(n3600), .ZN(n4585) );
  XNOR2_X2 U3755 ( .A(n3515), .B(n3514), .ZN(n3868) );
  XNOR2_X2 U3756 ( .A(n5526), .B(n4293), .ZN(n5459) );
  NOR2_X4 U3757 ( .A1(n5571), .A2(n5558), .ZN(n4241) );
  NAND2_X1 U3758 ( .A1(n3631), .A2(n3630), .ZN(n3652) );
  OR2_X1 U3759 ( .A1(n3758), .A2(n3665), .ZN(n3667) );
  INV_X1 U3760 ( .A(n4059), .ZN(n4043) );
  INV_X1 U3761 ( .A(n3908), .ZN(n4289) );
  INV_X1 U3762 ( .A(n5484), .ZN(n5502) );
  NAND2_X1 U3763 ( .A1(n5575), .A2(n5559), .ZN(n5549) );
  INV_X1 U3764 ( .A(n3925), .ZN(n4290) );
  OR2_X1 U3765 ( .A1(n4233), .A2(n6958), .ZN(n4260) );
  NOR2_X1 U3766 ( .A1(n5632), .A2(n3237), .ZN(n3235) );
  NOR2_X2 U3767 ( .A1(n5707), .A2(n5845), .ZN(n5698) );
  OR2_X1 U3768 ( .A1(n3759), .A2(n4306), .ZN(n3760) );
  OAI21_X1 U3769 ( .B1(n4306), .B2(n3758), .A(n3757), .ZN(n3761) );
  AOI21_X1 U3770 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6743), .A(n3756), 
        .ZN(n3757) );
  AOI22_X1 U3771 ( .A1(n3612), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3274) );
  NAND2_X1 U3772 ( .A1(n3620), .A2(n3619), .ZN(n3630) );
  OR2_X1 U3773 ( .A1(n3758), .A2(n3645), .ZN(n3620) );
  OR2_X1 U3774 ( .A1(n3502), .A2(n3501), .ZN(n3564) );
  INV_X1 U3775 ( .A(n3564), .ZN(n3507) );
  INV_X1 U3776 ( .A(n3769), .ZN(n3540) );
  INV_X1 U3777 ( .A(n4250), .ZN(n3541) );
  AND2_X2 U3778 ( .A1(n4521), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3272)
         );
  INV_X1 U3779 ( .A(n5670), .ZN(n3230) );
  NOR2_X1 U3780 ( .A1(n5674), .A2(n3232), .ZN(n3231) );
  NOR2_X1 U3781 ( .A1(n4737), .A2(n3229), .ZN(n3228) );
  INV_X1 U3782 ( .A(n4741), .ZN(n3229) );
  XNOR2_X1 U3783 ( .A(n3629), .B(n3630), .ZN(n3894) );
  NAND2_X1 U3784 ( .A1(n3220), .A2(n5492), .ZN(n3219) );
  INV_X1 U3785 ( .A(n5650), .ZN(n3220) );
  NOR2_X1 U3786 ( .A1(n5793), .A2(n3254), .ZN(n3253) );
  NAND2_X1 U3787 ( .A1(n5783), .A2(n3707), .ZN(n3254) );
  INV_X1 U3788 ( .A(n3705), .ZN(n3204) );
  INV_X1 U3789 ( .A(n5675), .ZN(n3213) );
  AND2_X1 U3790 ( .A1(n3215), .A2(n5407), .ZN(n3214) );
  INV_X1 U3791 ( .A(n5412), .ZN(n3215) );
  INV_X1 U3792 ( .A(n3671), .ZN(n3669) );
  INV_X1 U3793 ( .A(n3199), .ZN(n3198) );
  OAI21_X1 U3794 ( .B1(n3698), .B2(n3200), .A(n4940), .ZN(n3199) );
  INV_X1 U3795 ( .A(n4939), .ZN(n3200) );
  AND2_X1 U3796 ( .A1(n5473), .A2(n5662), .ZN(n5484) );
  OR2_X1 U3797 ( .A1(n3604), .A2(n4854), .ZN(n3605) );
  NAND2_X1 U3798 ( .A1(n4438), .A2(n5473), .ZN(n3221) );
  NOR2_X1 U3799 ( .A1(n3516), .A2(n3764), .ZN(n3476) );
  NAND2_X1 U3800 ( .A1(n5326), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5518) );
  OR2_X1 U3801 ( .A1(n5604), .A2(n5477), .ZN(n5651) );
  INV_X1 U3802 ( .A(n5528), .ZN(n3238) );
  INV_X1 U3803 ( .A(n4229), .ZN(n3856) );
  NAND2_X1 U3804 ( .A1(n4200), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4219)
         );
  NOR2_X1 U3805 ( .A1(n3234), .A2(n5628), .ZN(n3233) );
  INV_X1 U3806 ( .A(n3235), .ZN(n3234) );
  AND3_X1 U3807 ( .A1(n3993), .A2(n3992), .A3(n3991), .ZN(n5228) );
  NAND2_X1 U3808 ( .A1(n3912), .A2(n3911), .ZN(n4502) );
  NOR2_X1 U3809 ( .A1(n3217), .A2(n3179), .ZN(n5551) );
  NOR2_X1 U3810 ( .A1(n5536), .A2(n5662), .ZN(n3217) );
  NOR2_X1 U3811 ( .A1(n3176), .A2(n5573), .ZN(n5575) );
  AND2_X1 U3812 ( .A1(n5730), .A2(n3188), .ZN(n3209) );
  NAND2_X1 U3813 ( .A1(n5763), .A2(n3245), .ZN(n5756) );
  NAND2_X1 U3814 ( .A1(n6271), .A2(n5913), .ZN(n3245) );
  NAND2_X1 U3815 ( .A1(n5765), .A2(n5764), .ZN(n5763) );
  NAND2_X1 U3816 ( .A1(n6067), .A2(n5665), .ZN(n5604) );
  INV_X1 U3817 ( .A(n5662), .ZN(n5605) );
  NAND2_X1 U3818 ( .A1(n5408), .A2(n3214), .ZN(n5676) );
  NAND2_X1 U3819 ( .A1(n5361), .A2(n5360), .ZN(n5359) );
  OR2_X1 U3820 ( .A1(n6161), .A2(n5242), .ZN(n5370) );
  AOI21_X1 U3821 ( .B1(n4559), .B2(n6743), .A(n3556), .ZN(n3558) );
  OAI21_X1 U3822 ( .B1(n4242), .B2(n4241), .A(n5527), .ZN(n5687) );
  INV_X1 U3823 ( .A(n6308), .ZN(n6276) );
  NAND2_X1 U3824 ( .A1(n4602), .A2(n3770), .ZN(n6294) );
  INV_X1 U3825 ( .A(n3623), .ZN(n3645) );
  CLKBUF_X2 U3826 ( .A(n3434), .Z(n3442) );
  OR2_X1 U3827 ( .A1(n3555), .A2(n3554), .ZN(n3566) );
  OR2_X1 U3828 ( .A1(n3751), .A2(n3750), .ZN(n4307) );
  OAI211_X1 U3829 ( .C1(n3485), .C2(n5440), .A(n3486), .B(n3487), .ZN(n3535)
         );
  AOI22_X1 U3830 ( .A1(n3549), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3444), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3277) );
  NOR2_X1 U3831 ( .A1(n3854), .A2(n6116), .ZN(n4110) );
  INV_X1 U3832 ( .A(n4078), .ZN(n3854) );
  NOR2_X1 U3833 ( .A1(n6816), .A2(n3888), .ZN(n3889) );
  NOR2_X1 U3834 ( .A1(n4434), .A2(n5662), .ZN(n5495) );
  NAND2_X1 U3835 ( .A1(n4436), .A2(n4437), .ZN(n3222) );
  NAND2_X1 U3836 ( .A1(n3415), .A2(n3414), .ZN(n3223) );
  NAND2_X1 U3837 ( .A1(n4664), .A2(n6743), .ZN(n3241) );
  NOR2_X1 U3838 ( .A1(n4857), .A2(n6743), .ZN(n3426) );
  NAND2_X1 U3839 ( .A1(n4857), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3583) );
  NAND2_X1 U3840 ( .A1(n4673), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3584) );
  NAND2_X1 U3841 ( .A1(n3511), .A2(n3510), .ZN(n3513) );
  OR2_X1 U3842 ( .A1(n3595), .A2(n3594), .ZN(n3621) );
  INV_X1 U3843 ( .A(n3758), .ZN(n3736) );
  INV_X1 U3844 ( .A(n3729), .ZN(n3752) );
  OR2_X1 U3845 ( .A1(n3729), .A2(n3728), .ZN(n3759) );
  AND2_X1 U3846 ( .A1(n3584), .A2(n3583), .ZN(n3758) );
  AND2_X2 U3847 ( .A1(n4535), .A2(n4530), .ZN(n3434) );
  INV_X1 U3848 ( .A(n3480), .ZN(n3860) );
  INV_X1 U3849 ( .A(n4877), .ZN(n4749) );
  OAI21_X1 U3850 ( .B1(n4833), .B2(n4591), .A(n6629), .ZN(n4672) );
  INV_X1 U3851 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6607) );
  AND2_X1 U3852 ( .A1(n4570), .A2(n4569), .ZN(n6606) );
  AND2_X1 U3853 ( .A1(n5605), .A2(n5153), .ZN(n5497) );
  NOR2_X1 U3854 ( .A1(n4612), .A2(n4314), .ZN(n4364) );
  OR2_X1 U3855 ( .A1(n4313), .A2(n6638), .ZN(n4314) );
  OAI21_X1 U3856 ( .B1(n4289), .B2(n5717), .A(n4240), .ZN(n5558) );
  AND2_X1 U3857 ( .A1(n4195), .A2(n4194), .ZN(n5637) );
  NOR2_X1 U3858 ( .A1(n4165), .A2(n5766), .ZN(n4183) );
  AND2_X1 U3859 ( .A1(n4183), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4193)
         );
  NAND2_X1 U3860 ( .A1(n4149), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4165)
         );
  AND2_X1 U3861 ( .A1(n4130), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4149)
         );
  AND2_X1 U3862 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n4110), .ZN(n4130)
         );
  OR2_X1 U3863 ( .A1(n6111), .A2(n4289), .ZN(n4115) );
  INV_X1 U3864 ( .A(n5657), .ZN(n5672) );
  OR2_X1 U3866 ( .A1(n6118), .A2(n4289), .ZN(n4094) );
  AND2_X1 U3867 ( .A1(n4077), .A2(n4076), .ZN(n5674) );
  AND2_X1 U3868 ( .A1(n4004), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4008)
         );
  INV_X1 U3869 ( .A(n5377), .ZN(n4027) );
  AND2_X1 U3870 ( .A1(n3227), .A2(n3187), .ZN(n3226) );
  INV_X1 U3871 ( .A(n5228), .ZN(n3227) );
  NOR2_X1 U3872 ( .A1(n6975), .A2(n3962), .ZN(n3990) );
  INV_X1 U3873 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6975) );
  NAND2_X1 U3874 ( .A1(n3941), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3946)
         );
  AND2_X1 U3875 ( .A1(n3924), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3941)
         );
  NAND2_X1 U3876 ( .A1(n3907), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3915)
         );
  INV_X1 U3877 ( .A(n4431), .ZN(n3225) );
  AND2_X1 U3878 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3889), .ZN(n3907)
         );
  NOR2_X1 U3879 ( .A1(n4430), .A2(n4431), .ZN(n4432) );
  NAND2_X1 U3880 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3888) );
  OR2_X1 U3881 ( .A1(n5549), .A2(n5545), .ZN(n5536) );
  OR2_X1 U3882 ( .A1(n3191), .A2(n5621), .ZN(n3218) );
  NOR2_X1 U3883 ( .A1(n5889), .A2(n6985), .ZN(n3244) );
  NOR3_X1 U3884 ( .A1(n5651), .A2(n3191), .A3(n5650), .ZN(n5642) );
  NOR2_X1 U3885 ( .A1(n5651), .A2(n5650), .ZN(n5652) );
  NAND2_X1 U3886 ( .A1(n3256), .A2(n3255), .ZN(n5770) );
  NAND2_X1 U3887 ( .A1(n3171), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3255) );
  NAND2_X1 U3888 ( .A1(n5777), .A2(n3257), .ZN(n3256) );
  NAND2_X1 U3889 ( .A1(n6271), .A2(n3258), .ZN(n3257) );
  AND2_X1 U3890 ( .A1(n5408), .A2(n3190), .ZN(n6067) );
  INV_X1 U3891 ( .A(n3193), .ZN(n3212) );
  NAND2_X1 U3892 ( .A1(n3708), .A2(n3249), .ZN(n3248) );
  NOR2_X1 U3893 ( .A1(n5793), .A2(n3250), .ZN(n3249) );
  INV_X1 U3894 ( .A(n3707), .ZN(n3250) );
  AND2_X1 U3895 ( .A1(n3253), .A2(n3203), .ZN(n3202) );
  NAND2_X1 U3896 ( .A1(n3205), .A2(n3706), .ZN(n3201) );
  NAND2_X1 U3897 ( .A1(n3706), .A2(n3204), .ZN(n3203) );
  NAND2_X1 U3898 ( .A1(n5385), .A2(n3706), .ZN(n3708) );
  NAND2_X1 U3899 ( .A1(n3171), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5794) );
  OR2_X1 U3900 ( .A1(n6159), .A2(n6158), .ZN(n6161) );
  AND2_X1 U3901 ( .A1(n4704), .A2(n4703), .ZN(n4745) );
  NAND2_X1 U3902 ( .A1(n4745), .A2(n4744), .ZN(n6159) );
  AND2_X1 U3903 ( .A1(n4622), .A2(n5962), .ZN(n6348) );
  AND2_X1 U3904 ( .A1(n4636), .A2(n4635), .ZN(n4637) );
  NOR2_X1 U3905 ( .A1(n4638), .A2(n4637), .ZN(n4704) );
  OR2_X1 U3906 ( .A1(n4513), .A2(n4512), .ZN(n4638) );
  OR2_X1 U3907 ( .A1(n6727), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4250) );
  OR2_X1 U3908 ( .A1(n4489), .A2(n4488), .ZN(n4518) );
  NOR2_X1 U3909 ( .A1(n4518), .A2(n4517), .ZN(n4516) );
  OR2_X1 U3910 ( .A1(n6348), .A2(n4957), .ZN(n5815) );
  XNOR2_X1 U3911 ( .A(n3222), .B(n4438), .ZN(n4494) );
  AOI21_X1 U3912 ( .B1(n4614), .B2(n4613), .A(n6638), .ZN(n4627) );
  INV_X1 U3913 ( .A(n3763), .ZN(n3765) );
  INV_X1 U3914 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U3915 ( .A1(n3479), .A2(n3195), .ZN(n4526) );
  INV_X1 U3916 ( .A(n5094), .ZN(n4773) );
  CLKBUF_X1 U3917 ( .A(n3860), .Z(n3861) );
  NAND2_X1 U3918 ( .A1(n6718), .A2(n4672), .ZN(n4881) );
  AOI21_X1 U3919 ( .B1(n5177), .B2(STATE2_REG_3__SCAN_IN), .A(n4877), .ZN(
        n6488) );
  CLKBUF_X1 U3920 ( .A(n3908), .Z(n4834) );
  INV_X1 U3921 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n5263) );
  OR2_X1 U3922 ( .A1(n4364), .A2(n4336), .ZN(n6745) );
  NOR2_X1 U3923 ( .A1(n6001), .A2(n5510), .ZN(n5987) );
  NAND2_X1 U3924 ( .A1(n5418), .A2(n5417), .ZN(n6139) );
  INV_X1 U3925 ( .A(n6177), .ZN(n6167) );
  OR2_X1 U3926 ( .A1(n5518), .A2(n4859), .ZN(n6172) );
  INV_X1 U3927 ( .A(n6186), .ZN(n6175) );
  CLKBUF_X1 U3928 ( .A(n4664), .Z(n4665) );
  OR2_X1 U3929 ( .A1(n5518), .A2(n4847), .ZN(n5516) );
  OR2_X1 U3930 ( .A1(n5518), .A2(n4848), .ZN(n5131) );
  NAND2_X1 U3931 ( .A1(n4494), .A2(n5473), .ZN(n4849) );
  AND2_X1 U3932 ( .A1(n5326), .A2(n4843), .ZN(n6207) );
  INV_X1 U3933 ( .A(n6202), .ZN(n6193) );
  AND2_X1 U3934 ( .A1(n5551), .A2(n5550), .ZN(n5844) );
  AND2_X1 U3935 ( .A1(n4427), .A2(n4426), .ZN(n5634) );
  INV_X1 U3936 ( .A(n5678), .ZN(n6217) );
  INV_X2 U3937 ( .A(n5634), .ZN(n6221) );
  NAND2_X1 U3938 ( .A1(n3240), .A2(n3239), .ZN(n5684) );
  NAND2_X1 U3939 ( .A1(n5527), .A2(n5528), .ZN(n3239) );
  INV_X1 U3940 ( .A(n6240), .ZN(n6230) );
  OR2_X1 U3941 ( .A1(n6228), .A2(n6231), .ZN(n6236) );
  INV_X1 U3942 ( .A(n6236), .ZN(n5235) );
  CLKBUF_X1 U3943 ( .A(n6266), .Z(n6262) );
  CLKBUF_X1 U3944 ( .A(n4420), .Z(n4415) );
  INV_X1 U3945 ( .A(n4645), .ZN(n4418) );
  AND2_X1 U3946 ( .A1(n4233), .A2(n4230), .ZN(n5726) );
  INV_X1 U3947 ( .A(n5733), .ZN(n6029) );
  OR2_X1 U3948 ( .A1(n5629), .A2(n5618), .ZN(n6032) );
  INV_X1 U3949 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6816) );
  INV_X1 U3950 ( .A(n6063), .ZN(n6299) );
  NAND2_X1 U3951 ( .A1(n5698), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5700) );
  NOR2_X1 U3952 ( .A1(n5756), .A2(n3243), .ZN(n3242) );
  NAND2_X1 U3953 ( .A1(n6271), .A2(n3244), .ZN(n3243) );
  NAND2_X1 U3954 ( .A1(n5408), .A2(n5407), .ZN(n5413) );
  CLKBUF_X1 U3955 ( .A(n5385), .Z(n5387) );
  OR2_X1 U3956 ( .A1(n5803), .A2(n5940), .ZN(n6311) );
  NAND2_X1 U3957 ( .A1(n5159), .A2(n5160), .ZN(n6270) );
  CLKBUF_X1 U3958 ( .A(n4465), .Z(n4466) );
  INV_X1 U3959 ( .A(n5814), .ZN(n6392) );
  INV_X1 U3960 ( .A(n4819), .ZN(n4968) );
  INV_X1 U3961 ( .A(n3560), .ZN(n3561) );
  CLKBUF_X1 U3962 ( .A(n4559), .Z(n4560) );
  NOR2_X1 U3963 ( .A1(n5263), .A2(n4612), .ZN(n5448) );
  INV_X1 U3964 ( .A(n5448), .ZN(n6629) );
  INV_X1 U3965 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6978) );
  OR2_X1 U3966 ( .A1(n4969), .A2(n4968), .ZN(n5149) );
  AND2_X1 U3967 ( .A1(n6622), .A2(n6621), .ZN(n6639) );
  AND2_X1 U3968 ( .A1(n3769), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U3969 ( .A1(n4245), .A2(n4244), .ZN(n4254) );
  AND2_X1 U3970 ( .A1(n5403), .A2(n3231), .ZN(n3173) );
  OAI22_X1 U3971 ( .A1(n5359), .A2(n3201), .B1(n3202), .B2(n3251), .ZN(n5782)
         );
  NAND2_X1 U3972 ( .A1(n3208), .A2(n5739), .ZN(n3210) );
  OR2_X1 U3973 ( .A1(n5782), .A2(n5915), .ZN(n3174) );
  NAND2_X1 U3974 ( .A1(n4740), .A2(n4741), .ZN(n4736) );
  NAND2_X1 U3975 ( .A1(n4740), .A2(n3187), .ZN(n4996) );
  OR3_X1 U3976 ( .A1(n5651), .A2(n3219), .A3(n3191), .ZN(n3175) );
  OR3_X1 U3977 ( .A1(n5651), .A2(n3219), .A3(n3218), .ZN(n3176) );
  BUF_X1 U3978 ( .A(n3435), .Z(n4062) );
  NAND2_X1 U3979 ( .A1(n3210), .A2(n3209), .ZN(n5707) );
  NAND2_X1 U3980 ( .A1(n3248), .A2(n5794), .ZN(n5784) );
  NAND2_X1 U3981 ( .A1(n5587), .A2(n3236), .ZN(n5631) );
  AND2_X1 U3982 ( .A1(n5618), .A2(n5619), .ZN(n5570) );
  AND2_X1 U3983 ( .A1(n3246), .A2(n3247), .ZN(n3177) );
  NAND2_X1 U3984 ( .A1(n6271), .A2(n3700), .ZN(n3178) );
  AND2_X1 U3985 ( .A1(n5587), .A2(n5588), .ZN(n5586) );
  OAI21_X1 U3986 ( .B1(n3887), .B2(n3728), .A(n3605), .ZN(n3606) );
  AND2_X1 U3987 ( .A1(n5560), .A2(n5546), .ZN(n3179) );
  INV_X1 U3988 ( .A(n3251), .ZN(n3205) );
  NOR2_X1 U3989 ( .A1(n5794), .A2(n3252), .ZN(n3251) );
  NAND2_X1 U3990 ( .A1(n3543), .A2(n3542), .ZN(n3576) );
  AND2_X1 U3991 ( .A1(n5587), .A2(n3233), .ZN(n5618) );
  NAND2_X1 U3992 ( .A1(n3207), .A2(n3206), .ZN(n3208) );
  NAND2_X1 U3993 ( .A1(n3178), .A2(n5160), .ZN(n3180) );
  AND2_X1 U3994 ( .A1(n3238), .A2(n4242), .ZN(n3181) );
  AND2_X1 U3995 ( .A1(n3253), .A2(n3171), .ZN(n3182) );
  NAND2_X1 U3996 ( .A1(n5587), .A2(n3235), .ZN(n3183) );
  OR2_X1 U3997 ( .A1(n3400), .A2(n6737), .ZN(n3184) );
  AND2_X1 U3998 ( .A1(n4740), .A2(n3228), .ZN(n4735) );
  AND2_X2 U3999 ( .A1(n3477), .A2(n3476), .ZN(n4342) );
  AND2_X1 U4000 ( .A1(n3231), .A2(n6056), .ZN(n3185) );
  AND2_X1 U4001 ( .A1(n3214), .A2(n3213), .ZN(n3186) );
  NAND2_X1 U4002 ( .A1(n5403), .A2(n5404), .ZN(n5402) );
  AND2_X1 U4003 ( .A1(n3228), .A2(n3979), .ZN(n3187) );
  OAI21_X1 U4004 ( .B1(n4793), .B2(n3200), .A(n3198), .ZN(n5159) );
  NAND2_X1 U4005 ( .A1(n4793), .A2(n3698), .ZN(n4938) );
  INV_X1 U4006 ( .A(n5783), .ZN(n3252) );
  NAND2_X1 U4007 ( .A1(n3708), .A2(n3707), .ZN(n5792) );
  NAND2_X1 U4008 ( .A1(n5403), .A2(n3185), .ZN(n5669) );
  INV_X1 U4009 ( .A(n3237), .ZN(n3236) );
  NAND2_X1 U4010 ( .A1(n5637), .A2(n5588), .ZN(n3237) );
  NAND2_X1 U4011 ( .A1(n6271), .A2(n6887), .ZN(n3188) );
  AND2_X1 U4012 ( .A1(n3185), .A2(n3230), .ZN(n3189) );
  AND2_X1 U4013 ( .A1(n3186), .A2(n3212), .ZN(n3190) );
  NAND2_X1 U4014 ( .A1(n5639), .A2(n5640), .ZN(n3191) );
  XOR2_X1 U4015 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .Z(n3192) );
  OR2_X2 U4016 ( .A1(n3475), .A2(n4857), .ZN(n5153) );
  NAND2_X1 U4017 ( .A1(n5408), .A2(n3186), .ZN(n3216) );
  INV_X1 U4018 ( .A(n5404), .ZN(n3232) );
  NAND2_X1 U4019 ( .A1(n5469), .A2(n5468), .ZN(n3193) );
  INV_X1 U4020 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3258) );
  NAND3_X1 U4021 ( .A1(n6078), .A2(n5943), .A3(n6054), .ZN(n3194) );
  NAND2_X1 U4022 ( .A1(n4793), .A2(n3198), .ZN(n3196) );
  NAND2_X1 U4023 ( .A1(n3196), .A2(n3197), .ZN(n3703) );
  NAND2_X1 U4024 ( .A1(n5359), .A2(n3705), .ZN(n5385) );
  INV_X1 U4025 ( .A(n3711), .ZN(n3206) );
  INV_X1 U4026 ( .A(n3712), .ZN(n3207) );
  NAND2_X1 U4027 ( .A1(n3211), .A2(n3576), .ZN(n4572) );
  INV_X1 U4028 ( .A(n3575), .ZN(n3211) );
  NAND2_X1 U4029 ( .A1(n3534), .A2(n3535), .ZN(n3575) );
  INV_X2 U4030 ( .A(n3406), .ZN(n4873) );
  INV_X1 U4031 ( .A(n3216), .ZN(n6066) );
  NAND2_X1 U4032 ( .A1(n3222), .A2(n3221), .ZN(n4489) );
  XNOR2_X1 U4033 ( .A(n3223), .B(n3425), .ZN(n3874) );
  INV_X1 U4034 ( .A(n4430), .ZN(n3224) );
  NAND3_X1 U4035 ( .A1(n3224), .A2(n3225), .A3(n4502), .ZN(n4501) );
  AND2_X2 U4036 ( .A1(n5403), .A2(n3189), .ZN(n5657) );
  NAND2_X1 U4037 ( .A1(n4241), .A2(n4242), .ZN(n5527) );
  NAND2_X1 U4038 ( .A1(n4241), .A2(n3181), .ZN(n3240) );
  NAND2_X1 U4039 ( .A1(n3884), .A2(n3883), .ZN(n3885) );
  OAI21_X2 U4040 ( .B1(n4585), .B2(n4059), .A(n3925), .ZN(n3884) );
  NAND2_X1 U4041 ( .A1(n3708), .A2(n3182), .ZN(n3246) );
  NAND2_X2 U4042 ( .A1(n3177), .A2(n3174), .ZN(n5777) );
  INV_X1 U4043 ( .A(n5687), .ZN(n4245) );
  NOR2_X1 U4044 ( .A1(n3887), .A2(n4663), .ZN(n6528) );
  NAND2_X1 U4045 ( .A1(n3405), .A2(n3475), .ZN(n3762) );
  INV_X1 U4046 ( .A(n4319), .ZN(n3405) );
  NAND2_X1 U4047 ( .A1(n4299), .A2(n3482), .ZN(n4524) );
  OAI21_X1 U4048 ( .B1(n4585), .B2(n3728), .A(n3570), .ZN(n3571) );
  OR2_X2 U4049 ( .A1(n4873), .A2(n4857), .ZN(n4434) );
  XNOR2_X1 U4050 ( .A(n3526), .B(n3527), .ZN(n3515) );
  INV_X1 U4051 ( .A(n3629), .ZN(n3631) );
  CLKBUF_X1 U4052 ( .A(n5340), .Z(n5342) );
  AOI22_X1 U4053 ( .A1(n3391), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3429), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3276) );
  INV_X1 U4054 ( .A(n3559), .ZN(n3562) );
  OAI22_X1 U4055 ( .A1(n5770), .A2(n5771), .B1(n3171), .B2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5765) );
  AND2_X1 U4056 ( .A1(n3422), .A2(n3421), .ZN(n3259) );
  INV_X1 U4057 ( .A(n3475), .ZN(n4688) );
  AND2_X1 U4058 ( .A1(n4253), .A2(n4252), .ZN(n3260) );
  NOR2_X1 U4059 ( .A1(n4560), .A2(n4665), .ZN(n3261) );
  NOR2_X1 U4060 ( .A1(n4560), .A2(n5969), .ZN(n3262) );
  AOI21_X1 U4061 ( .B1(n3921), .B2(n4043), .A(n3920), .ZN(n4633) );
  INV_X1 U4062 ( .A(n4633), .ZN(n3922) );
  AND4_X1 U4063 ( .A1(n4563), .A2(n4320), .A3(n6641), .A4(n5153), .ZN(n3263)
         );
  INV_X1 U4064 ( .A(n3690), .ZN(n3512) );
  INV_X1 U4065 ( .A(n4647), .ZN(n3481) );
  INV_X1 U4066 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3914) );
  INV_X1 U4067 ( .A(n4995), .ZN(n3979) );
  NAND2_X1 U4068 ( .A1(n5379), .A2(n4029), .ZN(n5428) );
  OR2_X1 U4069 ( .A1(n5503), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3264)
         );
  INV_X1 U4070 ( .A(n6292), .ZN(n4244) );
  INV_X1 U4071 ( .A(n4735), .ZN(n4994) );
  AND2_X1 U4072 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3265) );
  INV_X1 U4073 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6435) );
  INV_X1 U4074 ( .A(n5697), .ZN(n6237) );
  AND2_X1 U4075 ( .A1(n5177), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3732)
         );
  OR2_X1 U4076 ( .A1(n3618), .A2(n3617), .ZN(n3623) );
  OR2_X1 U4077 ( .A1(n3641), .A2(n3640), .ZN(n3673) );
  AND2_X1 U4078 ( .A1(n3540), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3473)
         );
  INV_X1 U4079 ( .A(n4673), .ZN(n3310) );
  INV_X1 U4080 ( .A(n3566), .ZN(n3602) );
  NAND2_X1 U4081 ( .A1(n3474), .A2(n3402), .ZN(n3403) );
  INV_X1 U4082 ( .A(n5660), .ZN(n4134) );
  OR2_X1 U4083 ( .A1(n3729), .A2(n6978), .ZN(n3619) );
  NAND2_X1 U4084 ( .A1(n4845), .A2(n4880), .ZN(n3423) );
  INV_X1 U4085 ( .A(n3652), .ZN(n3654) );
  OR2_X1 U4086 ( .A1(n3758), .A2(n3642), .ZN(n3644) );
  OR2_X1 U4087 ( .A1(n3664), .A2(n3663), .ZN(n3683) );
  INV_X1 U4088 ( .A(n3569), .ZN(n3570) );
  NAND2_X1 U4089 ( .A1(n3533), .A2(n3532), .ZN(n3534) );
  OR2_X1 U4090 ( .A1(n3751), .A2(n3721), .ZN(n3722) );
  NAND2_X1 U4091 ( .A1(n3426), .A2(n3310), .ZN(n3729) );
  AND2_X1 U4092 ( .A1(n3667), .A2(n3666), .ZN(n3670) );
  OR2_X1 U4093 ( .A1(n6594), .A2(n6743), .ZN(n4286) );
  NAND2_X1 U4094 ( .A1(n3644), .A2(n3643), .ZN(n3653) );
  INV_X1 U4095 ( .A(n3762), .ZN(n3767) );
  INV_X1 U4096 ( .A(n3670), .ZN(n3668) );
  INV_X1 U4097 ( .A(n3524), .ZN(n3514) );
  NAND2_X1 U4098 ( .A1(n3562), .A2(n3561), .ZN(n3563) );
  INV_X1 U4099 ( .A(n3596), .ZN(n3597) );
  AND4_X1 U4100 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3372)
         );
  INV_X1 U4101 ( .A(n5516), .ZN(n5418) );
  NOR2_X1 U4102 ( .A1(n4260), .A2(n4259), .ZN(n4294) );
  NOR2_X1 U4103 ( .A1(n4030), .A2(n4031), .ZN(n4056) );
  OR2_X1 U4104 ( .A1(n3946), .A2(n4942), .ZN(n3962) );
  AND2_X1 U4105 ( .A1(n3481), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3895) );
  AND2_X1 U4106 ( .A1(n6269), .A2(n3701), .ZN(n3702) );
  INV_X1 U4107 ( .A(n3571), .ZN(n6300) );
  XNOR2_X1 U4108 ( .A(n3575), .B(n3576), .ZN(n4559) );
  INV_X1 U4109 ( .A(n3508), .ZN(n3462) );
  AND2_X1 U4110 ( .A1(n3472), .A2(n3538), .ZN(n5258) );
  INV_X1 U4111 ( .A(n5180), .ZN(n5217) );
  INV_X1 U4112 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6601) );
  AND2_X1 U4113 ( .A1(n4193), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4200)
         );
  NAND2_X1 U4114 ( .A1(n4056), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4061)
         );
  AND2_X1 U4115 ( .A1(n3990), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4004)
         );
  AND2_X1 U4116 ( .A1(n4187), .A2(n4186), .ZN(n5588) );
  INV_X1 U4117 ( .A(n5497), .ZN(n5503) );
  INV_X1 U4118 ( .A(n4292), .ZN(n4293) );
  NAND2_X1 U4119 ( .A1(n3856), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4233)
         );
  AND2_X1 U4120 ( .A1(n4167), .A2(n4166), .ZN(n5648) );
  NOR2_X1 U4121 ( .A1(n7050), .A2(n4061), .ZN(n4078) );
  NAND2_X1 U4122 ( .A1(n5709), .A2(n6910), .ZN(n5699) );
  NOR2_X1 U4123 ( .A1(n5343), .A2(n5345), .ZN(n5803) );
  NAND2_X1 U4124 ( .A1(n3508), .A2(n3510), .ZN(n3464) );
  OR2_X1 U4125 ( .A1(n4585), .A2(n3598), .ZN(n5094) );
  INV_X1 U4126 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n5177) );
  INV_X1 U4127 ( .A(n4671), .ZN(n5078) );
  AND2_X1 U4128 ( .A1(n5452), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3769) );
  INV_X1 U4129 ( .A(n6745), .ZN(n4838) );
  AND2_X1 U4130 ( .A1(n4312), .A2(n6640), .ZN(n4336) );
  OR2_X1 U4131 ( .A1(n4219), .A2(n3855), .ZN(n4229) );
  NAND2_X1 U4132 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n4008), .ZN(n4030)
         );
  AND2_X1 U4133 ( .A1(n4842), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4840) );
  AND2_X1 U4134 ( .A1(n5326), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6197) );
  INV_X1 U4135 ( .A(n5680), .ZN(n6218) );
  AND2_X1 U4136 ( .A1(n6240), .A2(n4650), .ZN(n6231) );
  NOR2_X1 U4137 ( .A1(n6747), .A2(n6241), .ZN(n6266) );
  NOR2_X1 U4138 ( .A1(n3915), .A2(n3914), .ZN(n3924) );
  INV_X1 U4139 ( .A(n4612), .ZN(n4602) );
  INV_X1 U4140 ( .A(n5815), .ZN(n6399) );
  INV_X1 U4141 ( .A(n6390), .ZN(n6383) );
  INV_X1 U4142 ( .A(n6370), .ZN(n6396) );
  NAND2_X1 U4143 ( .A1(n6743), .A2(n4672), .ZN(n4877) );
  INV_X1 U4144 ( .A(n4886), .ZN(n5080) );
  INV_X1 U4145 ( .A(n6459), .ZN(n6468) );
  INV_X1 U4146 ( .A(n5149), .ZN(n5120) );
  NOR2_X1 U4147 ( .A1(n4969), .A2(n4819), .ZN(n6477) );
  INV_X1 U4148 ( .A(n6514), .ZN(n6517) );
  AND2_X1 U4149 ( .A1(n4806), .A2(n4968), .ZN(n5297) );
  INV_X1 U4150 ( .A(n6581), .ZN(n6586) );
  AND2_X1 U4151 ( .A1(n3868), .A2(n4968), .ZN(n5175) );
  OR3_X1 U4152 ( .A1(n5566), .A2(n6704), .A3(n6705), .ZN(n5544) );
  INV_X1 U4153 ( .A(n6197), .ZN(n6171) );
  NAND2_X1 U4154 ( .A1(n5326), .A2(n4840), .ZN(n6177) );
  AND2_X1 U4155 ( .A1(n4841), .A2(n6177), .ZN(n6205) );
  NAND2_X1 U4156 ( .A1(n6240), .A2(n4649), .ZN(n5697) );
  AOI21_X1 U4157 ( .B1(n4842), .B2(n6276), .A(n4296), .ZN(n4297) );
  NAND2_X1 U4158 ( .A1(n6294), .A2(n4246), .ZN(n6063) );
  NAND2_X1 U4159 ( .A1(n6063), .A2(n4249), .ZN(n6308) );
  NAND2_X1 U4160 ( .A1(n4627), .A2(n4619), .ZN(n6370) );
  AND2_X1 U4161 ( .A1(n4668), .A2(n4667), .ZN(n5083) );
  NAND2_X1 U4162 ( .A1(n6406), .A2(n3887), .ZN(n6474) );
  INV_X1 U4163 ( .A(n6477), .ZN(n5123) );
  INV_X1 U4164 ( .A(n6478), .ZN(n5067) );
  OR2_X1 U4165 ( .A1(n4710), .A2(n4968), .ZN(n5014) );
  NAND2_X1 U4166 ( .A1(n6528), .A2(n5175), .ZN(n6592) );
  NAND2_X1 U4167 ( .A1(n4750), .A2(n4968), .ZN(n5087) );
  INV_X1 U4168 ( .A(n4755), .ZN(n5092) );
  INV_X1 U4169 ( .A(n6640), .ZN(n6638) );
  AND2_X1 U4170 ( .A1(n6628), .A2(n6627), .ZN(n6719) );
  INV_X1 U4171 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3266) );
  NOR2_X4 U4172 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4531) );
  AOI22_X1 U4173 ( .A1(n3427), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3271) );
  AND2_X4 U4174 ( .A1(n3272), .A2(n4530), .ZN(n3495) );
  NOR2_X1 U4175 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4176 ( .A1(n3495), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3270) );
  NOR2_X4 U4177 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4581) );
  AND2_X4 U4178 ( .A1(n4581), .A2(n4531), .ZN(n3435) );
  AND2_X4 U4179 ( .A1(n4530), .A2(n4520), .ZN(n3544) );
  AOI22_X1 U4180 ( .A1(n3435), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3268) );
  INV_X1 U4181 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4182 ( .A1(n3377), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4265), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3275) );
  NAND2_X2 U4183 ( .A1(n3279), .A2(n3278), .ZN(n3480) );
  AOI22_X1 U4184 ( .A1(n3549), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3377), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U4185 ( .A1(n3444), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3451), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4186 ( .A1(n3495), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        INSTQUEUE_REG_0__7__SCAN_IN), .B2(n3435), .ZN(n3281) );
  AOI22_X1 U4187 ( .A1(n3378), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4188 ( .A1(n3427), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4189 ( .A1(n3391), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4265), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4190 ( .A1(n3612), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4191 ( .A1(n3496), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3429), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3284) );
  NAND2_X2 U4192 ( .A1(n3289), .A2(n3288), .ZN(n3400) );
  NAND2_X1 U4193 ( .A1(n3860), .A2(n3400), .ZN(n3416) );
  INV_X1 U4194 ( .A(n3416), .ZN(n3311) );
  NAND2_X1 U4195 ( .A1(n3377), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3293) );
  NAND2_X1 U4196 ( .A1(n3451), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3292)
         );
  NAND2_X1 U4197 ( .A1(n3434), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3291)
         );
  NAND2_X1 U4198 ( .A1(n3495), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U4199 ( .A1(n3549), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3297)
         );
  NAND2_X1 U4200 ( .A1(n3444), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3296) );
  NAND2_X1 U4201 ( .A1(n3391), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3295) );
  NAND2_X1 U4202 ( .A1(n3429), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3294)
         );
  NAND2_X1 U4203 ( .A1(n3427), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3301) );
  NAND2_X1 U4204 ( .A1(n3612), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3300)
         );
  NAND2_X1 U4205 ( .A1(n3435), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3299) );
  NAND2_X1 U4206 ( .A1(n3589), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3298) );
  NAND2_X1 U4207 ( .A1(n3496), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3305) );
  NAND2_X1 U4208 ( .A1(n3378), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3304) );
  NAND2_X1 U4209 ( .A1(n4265), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3303) );
  NAND2_X1 U4210 ( .A1(n3544), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3302)
         );
  AND4_X4 U4211 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n4673)
         );
  NAND2_X1 U4212 ( .A1(n3434), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3315)
         );
  NAND2_X1 U4213 ( .A1(n3496), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3314) );
  NAND2_X1 U4214 ( .A1(n3377), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3313) );
  NAND2_X1 U4215 ( .A1(n3378), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U4216 ( .A1(n3427), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U4217 ( .A1(n3612), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3318)
         );
  NAND2_X1 U4218 ( .A1(n3495), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U4219 ( .A1(n3589), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4220 ( .A1(n3549), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3323)
         );
  NAND2_X1 U4221 ( .A1(n3451), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3322)
         );
  NAND2_X1 U4222 ( .A1(n3435), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U4223 ( .A1(n4265), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4224 ( .A1(n3444), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3327) );
  NAND2_X1 U4225 ( .A1(n3391), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3326) );
  NAND2_X1 U4226 ( .A1(n3429), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3325)
         );
  NAND2_X1 U4227 ( .A1(n3544), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3324)
         );
  NAND2_X2 U4228 ( .A1(n3480), .A2(n3407), .ZN(n4422) );
  AOI22_X1 U4229 ( .A1(n3444), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3331) );
  AOI22_X1 U4230 ( .A1(n3377), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3330) );
  AOI22_X1 U4231 ( .A1(n3496), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3329) );
  AOI22_X1 U4232 ( .A1(n3429), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3328) );
  AOI22_X1 U4233 ( .A1(n3427), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3495), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4234 ( .A1(n3451), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4235 ( .A1(n3549), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4265), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4236 ( .A1(n3612), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4237 ( .A1(n4422), .A2(n4880), .ZN(n3338) );
  NAND2_X1 U4238 ( .A1(n3338), .A2(n3400), .ZN(n3339) );
  NAND2_X1 U4239 ( .A1(n3763), .A2(n3339), .ZN(n3355) );
  INV_X1 U4240 ( .A(n3417), .ZN(n3418) );
  AOI22_X1 U4241 ( .A1(n3549), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3347) );
  AOI22_X1 U4242 ( .A1(n3444), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3434), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3346) );
  AOI22_X1 U4243 ( .A1(n3496), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3495), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4244 ( .A1(n3377), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3344) );
  NAND4_X1 U4245 ( .A1(n3347), .A2(n3346), .A3(n3345), .A4(n3344), .ZN(n3353)
         );
  AOI22_X1 U4246 ( .A1(n3428), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4265), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4247 ( .A1(n3427), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3451), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4248 ( .A1(n3435), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3429), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4249 ( .A1(n3612), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3348) );
  NAND4_X1 U4250 ( .A1(n3351), .A2(n3350), .A3(n3349), .A4(n3348), .ZN(n3352)
         );
  NAND2_X1 U4251 ( .A1(n3418), .A2(n3475), .ZN(n3354) );
  AND2_X2 U4252 ( .A1(n3355), .A2(n3354), .ZN(n4299) );
  NAND3_X1 U4253 ( .A1(n3416), .A2(n4422), .A3(n4673), .ZN(n4300) );
  NAND2_X1 U4254 ( .A1(n3549), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3359)
         );
  NAND2_X1 U4255 ( .A1(n3496), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3358) );
  NAND2_X1 U4256 ( .A1(n3428), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3357) );
  NAND2_X1 U4257 ( .A1(n3391), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4258 ( .A1(n3434), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3363)
         );
  NAND2_X1 U4259 ( .A1(n3451), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3362)
         );
  NAND2_X1 U4260 ( .A1(n3495), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3361) );
  NAND2_X1 U4261 ( .A1(n4265), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3360) );
  NAND2_X1 U4262 ( .A1(n3444), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3367) );
  NAND2_X1 U4263 ( .A1(n3377), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3366) );
  NAND2_X1 U4264 ( .A1(n3429), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3365)
         );
  NAND2_X1 U4265 ( .A1(n3544), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3364)
         );
  NAND2_X1 U4266 ( .A1(n3427), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3371) );
  NAND2_X1 U4267 ( .A1(n3612), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3370)
         );
  NAND2_X1 U4268 ( .A1(n3435), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3369) );
  NAND2_X1 U4269 ( .A1(n3589), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3368) );
  AOI21_X1 U4270 ( .B1(n4300), .B2(n4607), .A(n4603), .ZN(n3376) );
  NAND2_X1 U4271 ( .A1(n4299), .A2(n3376), .ZN(n3421) );
  NAND2_X1 U4272 ( .A1(n3434), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3382)
         );
  NAND2_X1 U4273 ( .A1(n3496), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3381) );
  NAND2_X1 U4274 ( .A1(n3377), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3380) );
  NAND2_X1 U4275 ( .A1(n3378), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3379) );
  NAND2_X1 U4276 ( .A1(n3549), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3386)
         );
  NAND2_X1 U4277 ( .A1(n3451), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3385)
         );
  NAND2_X1 U4278 ( .A1(n3435), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3384) );
  NAND2_X1 U4279 ( .A1(n4265), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4280 ( .A1(n3427), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4281 ( .A1(n3612), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3389)
         );
  NAND2_X1 U4282 ( .A1(n3495), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3388) );
  NAND2_X1 U4283 ( .A1(n3589), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U4284 ( .A1(n3444), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3395) );
  NAND2_X1 U4285 ( .A1(n3391), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3394) );
  NAND2_X1 U4286 ( .A1(n3429), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3393)
         );
  NAND2_X1 U4287 ( .A1(n3544), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3392)
         );
  AND4_X4 U4288 ( .A1(n3399), .A2(n3398), .A3(n3397), .A4(n3396), .ZN(n4857)
         );
  NAND2_X1 U4289 ( .A1(n3421), .A2(n4857), .ZN(n3411) );
  NAND2_X1 U4290 ( .A1(n4422), .A2(n3401), .ZN(n3474) );
  INV_X1 U4291 ( .A(n4854), .ZN(n3402) );
  NAND2_X1 U4292 ( .A1(n4673), .A2(n3764), .ZN(n3768) );
  INV_X1 U4293 ( .A(n3768), .ZN(n3734) );
  NAND2_X1 U4294 ( .A1(n3734), .A2(n5662), .ZN(n4527) );
  NAND2_X1 U4295 ( .A1(n3417), .A2(n4673), .ZN(n3404) );
  NAND3_X1 U4296 ( .A1(n3404), .A2(n3400), .A3(n4422), .ZN(n4319) );
  NAND3_X1 U4297 ( .A1(n3474), .A2(n4845), .A3(n3418), .ZN(n4321) );
  AOI21_X1 U4298 ( .B1(n3478), .B2(n4864), .A(n4607), .ZN(n3408) );
  NAND2_X1 U4299 ( .A1(n4321), .A2(n3408), .ZN(n3409) );
  NOR2_X1 U4300 ( .A1(n3762), .A2(n3409), .ZN(n3410) );
  NAND3_X1 U4301 ( .A1(n3411), .A2(n4327), .A3(n3410), .ZN(n3412) );
  NAND2_X1 U4302 ( .A1(n3412), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3485) );
  INV_X1 U4303 ( .A(n3485), .ZN(n3536) );
  NAND2_X1 U4304 ( .A1(n3536), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3415) );
  NAND2_X1 U4305 ( .A1(n5263), .A2(n5452), .ZN(n6727) );
  MUX2_X1 U4306 ( .A(n3540), .B(n3541), .S(n5177), .Z(n3413) );
  INV_X1 U4307 ( .A(n3413), .ZN(n3414) );
  INV_X1 U4308 ( .A(n3416), .ZN(n3873) );
  NOR2_X2 U4309 ( .A1(n3475), .A2(n4607), .ZN(n4424) );
  NAND3_X1 U4310 ( .A1(n3873), .A2(n4424), .A3(n3310), .ZN(n4563) );
  NAND2_X1 U4311 ( .A1(n6739), .A2(n3417), .ZN(n4320) );
  NOR2_X1 U4312 ( .A1(n6727), .A2(n6743), .ZN(n6641) );
  AND2_X1 U4313 ( .A1(n3418), .A2(n3310), .ZN(n3419) );
  OAI21_X1 U4314 ( .B1(n3762), .B2(n3419), .A(n4603), .ZN(n3420) );
  NAND2_X1 U4315 ( .A1(n3749), .A2(n4673), .ZN(n3422) );
  NAND2_X1 U4316 ( .A1(n3424), .A2(n4326), .ZN(n3471) );
  INV_X1 U4317 ( .A(n3471), .ZN(n3425) );
  NAND2_X1 U4318 ( .A1(n3874), .A2(n6743), .ZN(n3509) );
  INV_X1 U4319 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4699) );
  OR2_X1 U4320 ( .A1(n3729), .A2(n4699), .ZN(n3460) );
  AOI22_X1 U4321 ( .A1(n3450), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4322 ( .A1(n4261), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3451), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4323 ( .A1(n4264), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4324 ( .A1(n4099), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3430) );
  NAND4_X1 U4325 ( .A1(n3433), .A2(n3432), .A3(n3431), .A4(n3430), .ZN(n3441)
         );
  AOI22_X1 U4326 ( .A1(n3443), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4327 ( .A1(n3442), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4263), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4328 ( .A1(n4262), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3437) );
  BUF_X2 U4329 ( .A(n4265), .Z(n4172) );
  AOI22_X1 U4330 ( .A1(n4172), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3436) );
  NAND4_X1 U4331 ( .A1(n3439), .A2(n3438), .A3(n3437), .A4(n3436), .ZN(n3440)
         );
  AOI21_X1 U4332 ( .B1(n4857), .B2(n3565), .A(n6743), .ZN(n3458) );
  AOI22_X1 U4333 ( .A1(n3443), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4334 ( .A1(n4261), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4335 ( .A1(n4262), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3447) );
  BUF_X1 U4336 ( .A(n3544), .Z(n3445) );
  AOI22_X1 U4337 ( .A1(n4099), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3446) );
  NAND4_X1 U4338 ( .A1(n3449), .A2(n3448), .A3(n3447), .A4(n3446), .ZN(n3457)
         );
  BUF_X1 U4339 ( .A(n3495), .Z(n3450) );
  AOI22_X1 U4340 ( .A1(n4264), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3450), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4341 ( .A1(n3451), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4342 ( .A1(n4273), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4343 ( .A1(n4263), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3452) );
  NAND4_X1 U4344 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(n3456)
         );
  NAND2_X1 U4345 ( .A1(n4673), .A2(n3693), .ZN(n3461) );
  AND2_X1 U4346 ( .A1(n3458), .A2(n3461), .ZN(n3459) );
  NAND2_X1 U4347 ( .A1(n3460), .A2(n3459), .ZN(n3510) );
  NAND2_X1 U4348 ( .A1(n3509), .A2(n3510), .ZN(n3463) );
  NOR2_X1 U4349 ( .A1(n3584), .A2(n3693), .ZN(n3504) );
  MUX2_X1 U4350 ( .A(n3690), .B(n3504), .S(n3565), .Z(n3508) );
  NAND2_X1 U4351 ( .A1(n3463), .A2(n3462), .ZN(n3465) );
  NAND2_X2 U4352 ( .A1(n3465), .A2(n3464), .ZN(n4819) );
  NAND2_X1 U4353 ( .A1(n4857), .A2(n3475), .ZN(n3567) );
  OAI21_X1 U4354 ( .B1(n4854), .B2(n3565), .A(n3567), .ZN(n3466) );
  INV_X1 U4355 ( .A(n3466), .ZN(n3467) );
  NAND2_X1 U4356 ( .A1(n4357), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3468)
         );
  INV_X1 U4357 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U4358 ( .A1(n3468), .A2(n6852), .ZN(n3470) );
  AND2_X1 U4359 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3469) );
  NAND2_X1 U4360 ( .A1(n4357), .A2(n3469), .ZN(n3522) );
  AND2_X1 U4361 ( .A1(n3470), .A2(n3522), .ZN(n4453) );
  NAND2_X1 U4362 ( .A1(n5177), .A2(n6601), .ZN(n3472) );
  NAND2_X1 U4363 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3538) );
  AOI21_X1 U4364 ( .B1(n3541), .B2(n5258), .A(n3473), .ZN(n3486) );
  INV_X1 U4365 ( .A(n3474), .ZN(n3477) );
  NAND2_X1 U4366 ( .A1(n3475), .A2(n4880), .ZN(n3516) );
  NAND2_X1 U4367 ( .A1(n4342), .A2(n4845), .ZN(n4313) );
  INV_X1 U4368 ( .A(n3478), .ZN(n3483) );
  INV_X1 U4369 ( .A(n4839), .ZN(n3479) );
  NAND2_X1 U4370 ( .A1(n3480), .A2(n3400), .ZN(n4647) );
  NOR2_X1 U4371 ( .A1(n4300), .A2(n4839), .ZN(n3482) );
  NAND2_X1 U4372 ( .A1(n3484), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3487) );
  INV_X1 U4373 ( .A(n3486), .ZN(n3489) );
  INV_X1 U4374 ( .A(n3487), .ZN(n3488) );
  OAI21_X1 U4375 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3489), .A(n3488), 
        .ZN(n3490) );
  AND2_X2 U4376 ( .A1(n3535), .A2(n3490), .ZN(n3532) );
  AOI22_X1 U4377 ( .A1(n4272), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4378 ( .A1(n4261), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4379 ( .A1(n4273), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4380 ( .A1(n4262), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3491) );
  NAND4_X1 U4381 ( .A1(n3494), .A2(n3493), .A3(n3492), .A4(n3491), .ZN(n3502)
         );
  AOI22_X1 U4382 ( .A1(n4264), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4383 ( .A1(n3450), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4384 ( .A1(n4263), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4385 ( .A1(n3443), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3497) );
  NAND4_X1 U4386 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3501)
         );
  INV_X1 U4387 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5025) );
  OR2_X1 U4388 ( .A1(n3729), .A2(n5025), .ZN(n3506) );
  INV_X1 U4389 ( .A(n3504), .ZN(n3505) );
  OAI211_X1 U4390 ( .C1(n3507), .C2(n3583), .A(n3506), .B(n3505), .ZN(n3527)
         );
  NAND2_X1 U4391 ( .A1(n3509), .A2(n3462), .ZN(n3511) );
  NAND2_X1 U4392 ( .A1(n3868), .A2(n3749), .ZN(n3521) );
  XNOR2_X1 U4393 ( .A(n3565), .B(n3564), .ZN(n3518) );
  INV_X1 U4394 ( .A(n3516), .ZN(n3517) );
  OAI211_X1 U4395 ( .C1(n3518), .C2(n4854), .A(n3517), .B(n3764), .ZN(n3519)
         );
  INV_X1 U4396 ( .A(n3519), .ZN(n3520) );
  NAND2_X1 U4397 ( .A1(n3521), .A2(n3520), .ZN(n4452) );
  NAND2_X1 U4398 ( .A1(n4453), .A2(n4452), .ZN(n3523) );
  NAND2_X1 U4399 ( .A1(n3523), .A2(n3522), .ZN(n6302) );
  NAND2_X1 U4400 ( .A1(n6302), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3572)
         );
  NAND2_X1 U4401 ( .A1(n3526), .A2(n3527), .ZN(n3525) );
  NAND2_X1 U4402 ( .A1(n3525), .A2(n3524), .ZN(n3531) );
  INV_X1 U4403 ( .A(n3526), .ZN(n3529) );
  INV_X1 U4404 ( .A(n3527), .ZN(n3528) );
  NAND2_X1 U4405 ( .A1(n3529), .A2(n3528), .ZN(n3530) );
  NAND2_X1 U4407 ( .A1(n3577), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3543) );
  INV_X1 U4408 ( .A(n3538), .ZN(n3537) );
  NAND2_X1 U4409 ( .A1(n3537), .A2(n6607), .ZN(n6525) );
  NAND2_X1 U4410 ( .A1(n3538), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3539) );
  NAND2_X1 U4411 ( .A1(n6525), .A2(n3539), .ZN(n4675) );
  AOI22_X1 U4412 ( .A1(n3541), .A2(n4675), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3540), .ZN(n3542) );
  AOI22_X1 U4413 ( .A1(n3443), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4414 ( .A1(n4261), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3547) );
  INV_X1 U4415 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6948) );
  AOI22_X1 U4416 ( .A1(n4262), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4417 ( .A1(n4099), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3545) );
  NAND4_X1 U4418 ( .A1(n3548), .A2(n3547), .A3(n3546), .A4(n3545), .ZN(n3555)
         );
  AOI22_X1 U4419 ( .A1(n4264), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3450), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4420 ( .A1(n4272), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4421 ( .A1(n4273), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4422 ( .A1(n4263), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3550) );
  NAND4_X1 U4423 ( .A1(n3553), .A2(n3552), .A3(n3551), .A4(n3550), .ZN(n3554)
         );
  NOR2_X1 U4424 ( .A1(n3584), .A2(n3602), .ZN(n3556) );
  INV_X1 U4425 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5032) );
  OAI22_X1 U4426 ( .A1(n3729), .A2(n5032), .B1(n3602), .B2(n3583), .ZN(n3557)
         );
  XNOR2_X1 U4427 ( .A(n3558), .B(n3557), .ZN(n3559) );
  NAND2_X1 U4428 ( .A1(n3560), .A2(n3559), .ZN(n3600) );
  NAND2_X1 U4429 ( .A1(n3565), .A2(n3564), .ZN(n3603) );
  XNOR2_X1 U4430 ( .A(n3603), .B(n3566), .ZN(n3568) );
  OAI21_X1 U4431 ( .B1(n3568), .B2(n4854), .A(n3567), .ZN(n3569) );
  NAND2_X1 U4432 ( .A1(n3572), .A2(n6300), .ZN(n3574) );
  OR2_X1 U4433 ( .A1(n6302), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3573)
         );
  AND2_X1 U4434 ( .A1(n3574), .A2(n3573), .ZN(n4464) );
  INV_X1 U4435 ( .A(n3600), .ZN(n3599) );
  NAND2_X1 U4436 ( .A1(n3577), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3582) );
  NAND3_X1 U4437 ( .A1(n6435), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6490) );
  INV_X1 U4438 ( .A(n6490), .ZN(n3578) );
  NAND2_X1 U4439 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3578), .ZN(n6481) );
  NAND2_X1 U4440 ( .A1(n6435), .A2(n6481), .ZN(n3579) );
  NOR3_X1 U4441 ( .A1(n6435), .A2(n6607), .A3(n6601), .ZN(n4917) );
  NAND2_X1 U4442 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4917), .ZN(n4915) );
  NAND2_X1 U4443 ( .A1(n3579), .A2(n4915), .ZN(n4708) );
  OAI22_X1 U4444 ( .A1(n4250), .A2(n4708), .B1(n3769), .B2(n6435), .ZN(n3580)
         );
  INV_X1 U4445 ( .A(n3580), .ZN(n3581) );
  AOI22_X1 U4446 ( .A1(n4273), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4263), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4447 ( .A1(n4261), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4448 ( .A1(n3442), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4449 ( .A1(n4262), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3585) );
  NAND4_X1 U4450 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3595)
         );
  AOI22_X1 U4451 ( .A1(n4264), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4452 ( .A1(n3450), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4453 ( .A1(n4172), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3591) );
  AOI22_X1 U4454 ( .A1(n3443), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3590) );
  NAND4_X1 U4455 ( .A1(n3593), .A2(n3592), .A3(n3591), .A4(n3590), .ZN(n3594)
         );
  AOI22_X1 U4456 ( .A1(n3736), .A2(n3621), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3752), .ZN(n3596) );
  INV_X1 U4457 ( .A(n4587), .ZN(n3598) );
  NAND2_X1 U4458 ( .A1(n3600), .A2(n4587), .ZN(n3601) );
  NAND2_X1 U4459 ( .A1(n3603), .A2(n3602), .ZN(n3622) );
  XNOR2_X1 U4460 ( .A(n3622), .B(n3621), .ZN(n3604) );
  INV_X1 U4461 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6386) );
  XNOR2_X1 U4462 ( .A(n3606), .B(n6386), .ZN(n4463) );
  NAND2_X1 U4463 ( .A1(n4464), .A2(n4463), .ZN(n4465) );
  NAND2_X1 U4464 ( .A1(n3606), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3607)
         );
  NAND2_X1 U4465 ( .A1(n4465), .A2(n3607), .ZN(n6289) );
  AOI22_X1 U4466 ( .A1(n3443), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4467 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4261), .B1(n4271), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4468 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4262), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4469 ( .A1(n4099), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3608) );
  NAND4_X1 U4470 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3618)
         );
  AOI22_X1 U4471 ( .A1(n4264), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3450), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4472 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4272), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4473 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4273), .B1(n4172), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4474 ( .A1(n4263), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3613) );
  NAND4_X1 U4475 ( .A1(n3616), .A2(n3615), .A3(n3614), .A4(n3613), .ZN(n3617)
         );
  NAND2_X1 U4476 ( .A1(n3894), .A2(n3749), .ZN(n3626) );
  NAND2_X1 U4477 ( .A1(n3622), .A2(n3621), .ZN(n3646) );
  XNOR2_X1 U4478 ( .A(n3646), .B(n3623), .ZN(n3624) );
  NAND2_X1 U4479 ( .A1(n3624), .A2(n6739), .ZN(n3625) );
  NAND2_X1 U4480 ( .A1(n3626), .A2(n3625), .ZN(n3627) );
  INV_X1 U4481 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6377) );
  XNOR2_X1 U4482 ( .A(n3627), .B(n6377), .ZN(n6288) );
  NAND2_X1 U4483 ( .A1(n6289), .A2(n6288), .ZN(n6291) );
  NAND2_X1 U4484 ( .A1(n3627), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3628)
         );
  NAND2_X1 U4485 ( .A1(n6291), .A2(n3628), .ZN(n4505) );
  AOI22_X1 U4486 ( .A1(n4264), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4487 ( .A1(n3443), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4261), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4488 ( .A1(n3442), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4489 ( .A1(n3450), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3632) );
  NAND4_X1 U4490 ( .A1(n3635), .A2(n3634), .A3(n3633), .A4(n3632), .ZN(n3641)
         );
  AOI22_X1 U4491 ( .A1(n4273), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4492 ( .A1(n4262), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4493 ( .A1(n4263), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4494 ( .A1(n4099), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3636) );
  NAND4_X1 U4495 ( .A1(n3639), .A2(n3638), .A3(n3637), .A4(n3636), .ZN(n3640)
         );
  INV_X1 U4496 ( .A(n3673), .ZN(n3642) );
  INV_X1 U4497 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5082) );
  OR2_X1 U4498 ( .A1(n3729), .A2(n5082), .ZN(n3643) );
  XNOR2_X1 U4499 ( .A(n3652), .B(n3653), .ZN(n3906) );
  NAND2_X1 U4500 ( .A1(n3906), .A2(n3749), .ZN(n3649) );
  OR2_X1 U4501 ( .A1(n3646), .A2(n3645), .ZN(n3672) );
  XNOR2_X1 U4502 ( .A(n3672), .B(n3673), .ZN(n3647) );
  NAND2_X1 U4503 ( .A1(n3647), .A2(n6739), .ZN(n3648) );
  NAND2_X1 U4504 ( .A1(n3649), .A2(n3648), .ZN(n3650) );
  INV_X1 U4505 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6813) );
  XNOR2_X1 U4506 ( .A(n3650), .B(n6813), .ZN(n4504) );
  NAND2_X1 U4507 ( .A1(n4505), .A2(n4504), .ZN(n4503) );
  NAND2_X1 U4508 ( .A1(n3650), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3651)
         );
  NAND2_X1 U4509 ( .A1(n4503), .A2(n3651), .ZN(n6282) );
  NAND2_X1 U4510 ( .A1(n3654), .A2(n3653), .ZN(n3671) );
  AOI22_X1 U4511 ( .A1(n3443), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4512 ( .A1(n4261), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4513 ( .A1(n4262), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4514 ( .A1(n4099), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3655) );
  NAND4_X1 U4515 ( .A1(n3658), .A2(n3657), .A3(n3656), .A4(n3655), .ZN(n3664)
         );
  AOI22_X1 U4516 ( .A1(n4264), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3450), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4517 ( .A1(n4272), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4518 ( .A1(n4273), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4519 ( .A1(n4263), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3659) );
  NAND4_X1 U4520 ( .A1(n3662), .A2(n3661), .A3(n3660), .A4(n3659), .ZN(n3663)
         );
  INV_X1 U4521 ( .A(n3683), .ZN(n3665) );
  INV_X1 U4522 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5040) );
  OR2_X1 U4523 ( .A1(n3729), .A2(n5040), .ZN(n3666) );
  NAND2_X1 U4524 ( .A1(n3671), .A2(n3670), .ZN(n3921) );
  NAND3_X1 U4525 ( .A1(n3692), .A2(n3921), .A3(n3749), .ZN(n3677) );
  INV_X1 U4526 ( .A(n3672), .ZN(n3674) );
  NAND2_X1 U4527 ( .A1(n3674), .A2(n3673), .ZN(n3682) );
  XNOR2_X1 U4528 ( .A(n3682), .B(n3683), .ZN(n3675) );
  NAND2_X1 U4529 ( .A1(n3675), .A2(n6739), .ZN(n3676) );
  NAND2_X1 U4530 ( .A1(n3677), .A2(n3676), .ZN(n3678) );
  INV_X1 U4531 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6355) );
  XNOR2_X1 U4532 ( .A(n3678), .B(n6355), .ZN(n6281) );
  NAND2_X1 U4533 ( .A1(n6282), .A2(n6281), .ZN(n6280) );
  NAND2_X1 U4534 ( .A1(n3678), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3679)
         );
  NAND2_X1 U4535 ( .A1(n6280), .A2(n3679), .ZN(n4653) );
  INV_X1 U4536 ( .A(n3693), .ZN(n3680) );
  INV_X1 U4537 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4685) );
  OAI22_X1 U4538 ( .A1(n3758), .A2(n3680), .B1(n3729), .B2(n4685), .ZN(n3681)
         );
  NAND2_X1 U4539 ( .A1(n3930), .A2(n3749), .ZN(n3687) );
  INV_X1 U4540 ( .A(n3682), .ZN(n3684) );
  NAND2_X1 U4541 ( .A1(n3684), .A2(n3683), .ZN(n3695) );
  XNOR2_X1 U4542 ( .A(n3695), .B(n3693), .ZN(n3685) );
  NAND2_X1 U4543 ( .A1(n3685), .A2(n6739), .ZN(n3686) );
  NAND2_X1 U4544 ( .A1(n3687), .A2(n3686), .ZN(n3688) );
  INV_X1 U4545 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6342) );
  XNOR2_X1 U4546 ( .A(n3688), .B(n6342), .ZN(n4652) );
  NAND2_X1 U4547 ( .A1(n4653), .A2(n4652), .ZN(n4651) );
  NAND2_X1 U4548 ( .A1(n3688), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3689)
         );
  NAND2_X1 U4549 ( .A1(n4651), .A2(n3689), .ZN(n4795) );
  NOR2_X1 U4550 ( .A1(n3512), .A2(n3728), .ZN(n3691) );
  NAND2_X1 U4551 ( .A1(n6739), .A2(n3693), .ZN(n3694) );
  OR2_X1 U4552 ( .A1(n3695), .A2(n3694), .ZN(n3696) );
  NAND2_X1 U4553 ( .A1(n6271), .A2(n3696), .ZN(n3697) );
  INV_X1 U4554 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4961) );
  XNOR2_X1 U4555 ( .A(n3697), .B(n4961), .ZN(n4794) );
  NAND2_X1 U4556 ( .A1(n4795), .A2(n4794), .ZN(n4793) );
  NAND2_X1 U4557 ( .A1(n3697), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3698)
         );
  INV_X1 U4558 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U4559 ( .A1(n6271), .A2(n6316), .ZN(n4939) );
  NAND2_X1 U4560 ( .A1(n3171), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4940)
         );
  INV_X1 U4561 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U4562 ( .A1(n6271), .A2(n3699), .ZN(n5160) );
  INV_X1 U4563 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U4564 ( .A1(n3171), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U4565 ( .A1(n3171), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3701) );
  NAND2_X1 U4566 ( .A1(n3703), .A2(n3702), .ZN(n5340) );
  INV_X1 U4567 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6885) );
  XNOR2_X1 U4568 ( .A(n6271), .B(n6885), .ZN(n5341) );
  NAND2_X1 U4569 ( .A1(n6271), .A2(n6885), .ZN(n3704) );
  OAI21_X2 U4570 ( .B1(n5340), .B2(n5341), .A(n3704), .ZN(n5361) );
  XNOR2_X1 U4571 ( .A(n6271), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5360)
         );
  INV_X1 U4572 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U4573 ( .A1(n6271), .A2(n5375), .ZN(n3705) );
  NAND2_X1 U4574 ( .A1(n3171), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3706) );
  INV_X1 U4575 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U4576 ( .A1(n6271), .A2(n5392), .ZN(n3707) );
  INV_X1 U4577 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6073) );
  AND2_X1 U4578 ( .A1(n6271), .A2(n6073), .ZN(n5793) );
  NAND2_X1 U4579 ( .A1(n6271), .A2(n6078), .ZN(n5783) );
  INV_X1 U4580 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5943) );
  INV_X1 U4581 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U4582 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5915) );
  AND2_X1 U4583 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5897) );
  AND2_X1 U4584 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5923) );
  AND2_X1 U4585 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5824) );
  AND3_X1 U4586 ( .A1(n5897), .A2(n5923), .A3(n5824), .ZN(n3709) );
  AOI21_X1 U4587 ( .B1(n5777), .B2(n3709), .A(n3171), .ZN(n3712) );
  NOR2_X1 U4588 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5924) );
  NOR2_X1 U4589 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5898) );
  INV_X1 U4590 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5742) );
  INV_X1 U4591 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5889) );
  NAND4_X1 U4592 ( .A1(n5924), .A2(n5898), .A3(n5742), .A4(n5889), .ZN(n3710)
         );
  NOR2_X1 U4593 ( .A1(n5777), .A2(n3710), .ZN(n3711) );
  XNOR2_X1 U4594 ( .A(n6271), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5739)
         );
  INV_X1 U4595 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6887) );
  INV_X1 U4596 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U4597 ( .A1(n3171), .A2(n5867), .ZN(n5728) );
  INV_X1 U4598 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5710) );
  INV_X1 U4599 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U4600 ( .A1(n5710), .A2(n5708), .ZN(n3713) );
  NOR2_X1 U4601 ( .A1(n3171), .A2(n5867), .ZN(n5730) );
  NAND2_X1 U4602 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5845) );
  NOR2_X1 U4603 ( .A1(n5709), .A2(n5698), .ZN(n3714) );
  INV_X1 U4604 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6910) );
  XNOR2_X1 U4605 ( .A(n3714), .B(n6910), .ZN(n5851) );
  XNOR2_X1 U4606 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3727) );
  NAND2_X1 U4607 ( .A1(n3732), .A2(n3727), .ZN(n3716) );
  NAND2_X1 U4608 ( .A1(n6601), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4609 ( .A1(n3716), .A2(n3715), .ZN(n3726) );
  XNOR2_X1 U4610 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3725) );
  NAND2_X1 U4611 ( .A1(n3726), .A2(n3725), .ZN(n3718) );
  NAND2_X1 U4612 ( .A1(n6607), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3717) );
  NAND2_X1 U4613 ( .A1(n3718), .A2(n3717), .ZN(n3724) );
  MUX2_X1 U4614 ( .A(n6435), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n3723) );
  NAND2_X1 U4615 ( .A1(n3724), .A2(n3723), .ZN(n3720) );
  NAND2_X1 U4616 ( .A1(n6435), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3719) );
  NAND2_X1 U4617 ( .A1(n3720), .A2(n3719), .ZN(n3751) );
  INV_X1 U4618 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6611) );
  AND2_X1 U4619 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6611), .ZN(n3721)
         );
  INV_X1 U4620 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U4621 ( .A1(n4575), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3750) );
  NAND2_X1 U4622 ( .A1(n3722), .A2(n3750), .ZN(n4306) );
  XNOR2_X1 U4623 ( .A(n3724), .B(n3723), .ZN(n4302) );
  OAI21_X1 U4624 ( .B1(n4857), .B2(n3764), .A(n4873), .ZN(n3743) );
  XNOR2_X1 U4625 ( .A(n3726), .B(n3725), .ZN(n4303) );
  NOR3_X1 U4626 ( .A1(n3758), .A2(n3743), .A3(n4303), .ZN(n3748) );
  XNOR2_X1 U4627 ( .A(n3727), .B(n3732), .ZN(n4304) );
  INV_X1 U4628 ( .A(n3759), .ZN(n3742) );
  AOI21_X1 U4629 ( .B1(n3736), .B2(n4603), .A(n4864), .ZN(n3738) );
  NOR3_X1 U4630 ( .A1(n3738), .A2(n4304), .A3(n6743), .ZN(n3741) );
  AND2_X1 U4631 ( .A1(n3730), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3731)
         );
  NOR2_X1 U4632 ( .A1(n3732), .A2(n3731), .ZN(n3735) );
  INV_X1 U4633 ( .A(n3735), .ZN(n3733) );
  OAI21_X1 U4634 ( .B1(n3734), .B2(n3733), .A(n4845), .ZN(n3739) );
  NAND2_X1 U4635 ( .A1(n3736), .A2(n3735), .ZN(n3737) );
  AOI222_X1 U4636 ( .A1(n3739), .A2(n3743), .B1(n4304), .B2(n3738), .C1(n3737), 
        .C2(n3759), .ZN(n3740) );
  AOI211_X1 U4637 ( .C1(n4304), .C2(n3742), .A(n3741), .B(n3740), .ZN(n3746)
         );
  OAI21_X1 U4638 ( .B1(n3758), .B2(n4303), .A(n3743), .ZN(n3744) );
  AOI21_X1 U4639 ( .B1(n3752), .B2(n4303), .A(n3744), .ZN(n3745) );
  NOR2_X1 U4640 ( .A1(n3746), .A2(n3745), .ZN(n3747) );
  AOI211_X1 U4641 ( .C1(n3749), .C2(n4302), .A(n3748), .B(n3747), .ZN(n3755)
         );
  INV_X1 U4642 ( .A(n4302), .ZN(n3753) );
  AOI21_X1 U4643 ( .B1(n3753), .B2(n4307), .A(n3752), .ZN(n3754) );
  OAI22_X1 U4644 ( .A1(n3755), .A2(n3754), .B1(n3759), .B2(n4307), .ZN(n3756)
         );
  NAND2_X1 U4645 ( .A1(n3765), .A2(n3764), .ZN(n6594) );
  NAND2_X1 U4646 ( .A1(n6594), .A2(n4857), .ZN(n3766) );
  NAND3_X1 U4647 ( .A1(n3767), .A2(n4880), .A3(n3766), .ZN(n4547) );
  OR2_X1 U4648 ( .A1(n4547), .A2(n3768), .ZN(n6615) );
  NOR2_X1 U4649 ( .A1(n6615), .A2(n6638), .ZN(n3770) );
  AOI22_X1 U4650 ( .A1(n3443), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4651 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3442), .B1(n4270), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4652 ( .A1(n4273), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4653 ( .A1(n4099), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3771) );
  NAND4_X1 U4654 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3780)
         );
  AOI22_X1 U4655 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4262), .B1(n4261), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4656 ( .A1(n4264), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4263), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4657 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4271), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4658 ( .A1(n3450), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3775) );
  NAND4_X1 U4659 ( .A1(n3778), .A2(n3777), .A3(n3776), .A4(n3775), .ZN(n3779)
         );
  NOR2_X1 U4660 ( .A1(n3780), .A2(n3779), .ZN(n4224) );
  AOI22_X1 U4661 ( .A1(n4273), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4662 ( .A1(n4264), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4263), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4663 ( .A1(n3442), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4664 ( .A1(n3450), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3781) );
  NAND4_X1 U4665 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3790)
         );
  AOI22_X1 U4666 ( .A1(n4261), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4667 ( .A1(n4262), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4668 ( .A1(n3443), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4669 ( .A1(n4099), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4670 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3789)
         );
  NOR2_X1 U4671 ( .A1(n3790), .A2(n3789), .ZN(n4205) );
  AOI22_X1 U4672 ( .A1(n4263), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4673 ( .A1(n4261), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3793) );
  AOI22_X1 U4674 ( .A1(n3442), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4675 ( .A1(n4099), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3791) );
  NAND4_X1 U4676 ( .A1(n3794), .A2(n3793), .A3(n3792), .A4(n3791), .ZN(n3800)
         );
  AOI22_X1 U4677 ( .A1(n4272), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3450), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4678 ( .A1(n3443), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4273), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4679 ( .A1(n4262), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4680 ( .A1(n4264), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3795) );
  NAND4_X1 U4681 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3799)
         );
  NOR2_X1 U4682 ( .A1(n3800), .A2(n3799), .ZN(n4188) );
  AOI22_X1 U4683 ( .A1(n4262), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4684 ( .A1(n4271), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4685 ( .A1(n3443), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4686 ( .A1(n3495), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3801) );
  NAND4_X1 U4687 ( .A1(n3804), .A2(n3803), .A3(n3802), .A4(n3801), .ZN(n3810)
         );
  AOI22_X1 U4688 ( .A1(n4273), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4689 ( .A1(n4264), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4263), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4690 ( .A1(n4270), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4691 ( .A1(n4261), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3805) );
  NAND4_X1 U4692 ( .A1(n3808), .A2(n3807), .A3(n3806), .A4(n3805), .ZN(n3809)
         );
  NOR2_X1 U4693 ( .A1(n3810), .A2(n3809), .ZN(n4189) );
  OR2_X1 U4694 ( .A1(n4188), .A2(n4189), .ZN(n4198) );
  AOI22_X1 U4695 ( .A1(n4261), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4696 ( .A1(n4262), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4697 ( .A1(n4263), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3812) );
  INV_X1 U4698 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n7037) );
  AOI22_X1 U4699 ( .A1(n3442), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3811) );
  NAND4_X1 U4700 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(n3820)
         );
  AOI22_X1 U4701 ( .A1(n3443), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4702 ( .A1(n4273), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4703 ( .A1(n3450), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4704 ( .A1(n3445), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3815) );
  NAND4_X1 U4705 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3819)
         );
  NOR2_X1 U4706 ( .A1(n3820), .A2(n3819), .ZN(n4196) );
  OR2_X1 U4707 ( .A1(n4198), .A2(n4196), .ZN(n4204) );
  NOR2_X1 U4708 ( .A1(n4205), .A2(n4204), .ZN(n4214) );
  AOI22_X1 U4709 ( .A1(n3443), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4710 ( .A1(n4261), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4711 ( .A1(n4262), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4712 ( .A1(n4099), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3821) );
  NAND4_X1 U4713 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3830)
         );
  AOI22_X1 U4714 ( .A1(n4264), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3450), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4715 ( .A1(n4272), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4716 ( .A1(n4273), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4717 ( .A1(n4263), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3825) );
  NAND4_X1 U4718 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3829)
         );
  OR2_X1 U4719 ( .A1(n3830), .A2(n3829), .ZN(n4212) );
  NAND2_X1 U4720 ( .A1(n4214), .A2(n4212), .ZN(n4225) );
  NOR2_X1 U4721 ( .A1(n4224), .A2(n4225), .ZN(n4236) );
  AOI22_X1 U4722 ( .A1(n3443), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4723 ( .A1(n4261), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4724 ( .A1(n4262), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4725 ( .A1(n4099), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3831) );
  NAND4_X1 U4726 ( .A1(n3834), .A2(n3833), .A3(n3832), .A4(n3831), .ZN(n3840)
         );
  AOI22_X1 U4727 ( .A1(n4264), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3450), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3838) );
  AOI22_X1 U4728 ( .A1(n4272), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4729 ( .A1(n4273), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4730 ( .A1(n4263), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3835) );
  NAND4_X1 U4731 ( .A1(n3838), .A2(n3837), .A3(n3836), .A4(n3835), .ZN(n3839)
         );
  OR2_X1 U4732 ( .A1(n3840), .A2(n3839), .ZN(n4235) );
  NAND2_X1 U4733 ( .A1(n4236), .A2(n4235), .ZN(n4280) );
  AOI22_X1 U4734 ( .A1(n3442), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4735 ( .A1(n4264), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4736 ( .A1(n4273), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4737 ( .A1(n4099), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4738 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3851)
         );
  AOI22_X1 U4739 ( .A1(n4272), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3450), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4740 ( .A1(n4262), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4261), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4741 ( .A1(n3443), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4742 ( .A1(n4263), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4265), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3846) );
  NAND4_X1 U4743 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3850)
         );
  NOR2_X1 U4744 ( .A1(n3851), .A2(n3850), .ZN(n4281) );
  XOR2_X1 U4745 ( .A(n4280), .B(n4281), .Z(n3852) );
  INV_X1 U4746 ( .A(n4286), .ZN(n4226) );
  NAND2_X1 U4747 ( .A1(n3852), .A2(n4226), .ZN(n3859) );
  INV_X2 U4748 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6737) );
  INV_X1 U4749 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4259) );
  AOI21_X1 U4750 ( .B1(n4259), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3853) );
  AOI21_X1 U4751 ( .B1(n4291), .B2(EAX_REG_29__SCAN_IN), .A(n3853), .ZN(n3858)
         );
  NOR2_X1 U4752 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3908) );
  INV_X1 U4753 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n7050) );
  INV_X1 U4754 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4031) );
  INV_X1 U4755 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6116) );
  INV_X1 U4756 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U4757 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3855) );
  INV_X1 U4758 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6958) );
  INV_X1 U4759 ( .A(n4260), .ZN(n3857) );
  XOR2_X1 U4760 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .B(n3857), .Z(n5552) );
  AOI22_X1 U4761 ( .A1(n3859), .A2(n3858), .B1(n4834), .B2(n5552), .ZN(n4242)
         );
  NAND2_X1 U4762 ( .A1(n3861), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4059) );
  NAND2_X1 U4763 ( .A1(n6737), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3925) );
  INV_X1 U4764 ( .A(n3884), .ZN(n3867) );
  NAND2_X1 U4765 ( .A1(n3895), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3866) );
  OAI21_X1 U4766 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3888), .ZN(n6307) );
  NAND2_X1 U4767 ( .A1(n3908), .A2(n6307), .ZN(n3863) );
  NAND2_X1 U4768 ( .A1(n4290), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3862)
         );
  NAND2_X1 U4769 ( .A1(n3863), .A2(n3862), .ZN(n3864) );
  AOI21_X1 U4770 ( .B1(n4291), .B2(EAX_REG_2__SCAN_IN), .A(n3864), .ZN(n3865)
         );
  AND2_X1 U4771 ( .A1(n3866), .A2(n3865), .ZN(n3882) );
  NAND2_X1 U4772 ( .A1(n3867), .A2(n3882), .ZN(n4486) );
  NAND2_X1 U4773 ( .A1(n3868), .A2(n4043), .ZN(n3872) );
  INV_X2 U4774 ( .A(n3184), .ZN(n4291) );
  AOI22_X1 U4775 ( .A1(n4291), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6737), .ZN(n3870) );
  NAND2_X1 U4776 ( .A1(n3895), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3869) );
  AND2_X1 U4777 ( .A1(n3870), .A2(n3869), .ZN(n3871) );
  NAND2_X1 U4778 ( .A1(n3872), .A2(n3871), .ZN(n4456) );
  NAND2_X1 U4779 ( .A1(n4819), .A2(n3873), .ZN(n4352) );
  NAND2_X1 U4780 ( .A1(n6597), .A2(n4043), .ZN(n3878) );
  AOI22_X1 U4781 ( .A1(n4291), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6737), .ZN(n3876) );
  NAND2_X1 U4782 ( .A1(n3895), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3875) );
  AND2_X1 U4783 ( .A1(n3876), .A2(n3875), .ZN(n3877) );
  NAND2_X1 U4784 ( .A1(n3878), .A2(n3877), .ZN(n3880) );
  AND2_X1 U4785 ( .A1(n3880), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3879) );
  NAND2_X1 U4786 ( .A1(n4352), .A2(n3879), .ZN(n4355) );
  INV_X1 U4787 ( .A(n3880), .ZN(n4353) );
  NAND2_X1 U4788 ( .A1(n4353), .A2(n3908), .ZN(n3881) );
  NAND2_X1 U4789 ( .A1(n4355), .A2(n3881), .ZN(n4455) );
  NAND2_X1 U4790 ( .A1(n4456), .A2(n4455), .ZN(n4454) );
  INV_X1 U4791 ( .A(n3882), .ZN(n3883) );
  NAND2_X1 U4792 ( .A1(n4454), .A2(n3885), .ZN(n3886) );
  NAND2_X1 U4793 ( .A1(n6816), .A2(n3888), .ZN(n3890) );
  INV_X1 U4794 ( .A(n3889), .ZN(n3900) );
  AND2_X1 U4795 ( .A1(n3890), .A2(n3900), .ZN(n6208) );
  OAI22_X1 U4796 ( .A1(n4289), .A2(n6208), .B1(n3925), .B2(n6816), .ZN(n3891)
         );
  AOI21_X1 U4797 ( .B1(n4291), .B2(EAX_REG_3__SCAN_IN), .A(n3891), .ZN(n3893)
         );
  NAND2_X1 U4798 ( .A1(n3895), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3892) );
  INV_X1 U4799 ( .A(n3895), .ZN(n3898) );
  NAND2_X1 U4800 ( .A1(n6737), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3897)
         );
  NAND2_X1 U4801 ( .A1(n4291), .A2(EAX_REG_4__SCAN_IN), .ZN(n3896) );
  OAI211_X1 U4802 ( .C1(n3898), .C2(n4575), .A(n3897), .B(n3896), .ZN(n3899)
         );
  NAND2_X1 U4803 ( .A1(n3899), .A2(n4289), .ZN(n3904) );
  INV_X1 U4804 ( .A(n3907), .ZN(n3902) );
  NAND2_X1 U4805 ( .A1(n6911), .A2(n3900), .ZN(n3901) );
  NAND2_X1 U4806 ( .A1(n3902), .A2(n3901), .ZN(n6298) );
  NAND2_X1 U4807 ( .A1(n6298), .A2(n4834), .ZN(n3903) );
  NAND2_X1 U4808 ( .A1(n3904), .A2(n3903), .ZN(n3905) );
  NAND2_X1 U4809 ( .A1(n3906), .A2(n4043), .ZN(n3912) );
  INV_X1 U4810 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5167) );
  OAI21_X1 U4811 ( .B1(n3907), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3915), 
        .ZN(n5170) );
  NAND2_X1 U4812 ( .A1(n5170), .A2(n4834), .ZN(n3909) );
  OAI21_X1 U4813 ( .B1(n5167), .B2(n3925), .A(n3909), .ZN(n3910) );
  AOI21_X1 U4814 ( .B1(n4291), .B2(EAX_REG_5__SCAN_IN), .A(n3910), .ZN(n3911)
         );
  INV_X1 U4815 ( .A(n4501), .ZN(n3923) );
  NAND2_X1 U4816 ( .A1(n4291), .A2(EAX_REG_6__SCAN_IN), .ZN(n3919) );
  AOI21_X1 U4817 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3914), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3913) );
  INV_X1 U4818 ( .A(n3913), .ZN(n3918) );
  AND2_X1 U4819 ( .A1(n3915), .A2(n3914), .ZN(n3916) );
  OR2_X1 U4820 ( .A1(n3916), .A2(n3924), .ZN(n6287) );
  NOR2_X1 U4821 ( .A1(n6287), .A2(n4289), .ZN(n3917) );
  AOI21_X1 U4822 ( .B1(n3919), .B2(n3918), .A(n3917), .ZN(n3920) );
  INV_X1 U4823 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3928) );
  XNOR2_X1 U4824 ( .A(n3924), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5252) );
  INV_X1 U4825 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5248) );
  NOR2_X1 U4826 ( .A1(n3925), .A2(n5248), .ZN(n3926) );
  AOI21_X1 U4827 ( .B1(n5252), .B2(n4834), .A(n3926), .ZN(n3927) );
  OAI21_X1 U4828 ( .B1(n3184), .B2(n3928), .A(n3927), .ZN(n3929) );
  AOI21_X2 U4829 ( .B1(n3930), .B2(n4043), .A(n3929), .ZN(n4654) );
  AOI22_X1 U4830 ( .A1(n4273), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4831 ( .A1(n4270), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4832 ( .A1(n4263), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4833 ( .A1(n4271), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3931) );
  NAND4_X1 U4834 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3940)
         );
  AOI22_X1 U4835 ( .A1(n4261), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4836 ( .A1(n4262), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4837 ( .A1(n3450), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4838 ( .A1(n3443), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3935) );
  NAND4_X1 U4839 ( .A1(n3938), .A2(n3937), .A3(n3936), .A4(n3935), .ZN(n3939)
         );
  OAI21_X1 U4840 ( .B1(n3940), .B2(n3939), .A(n4043), .ZN(n3945) );
  NAND2_X1 U4841 ( .A1(n4291), .A2(EAX_REG_8__SCAN_IN), .ZN(n3944) );
  XNOR2_X1 U4842 ( .A(n3941), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U4843 ( .A1(n5309), .A2(n4834), .ZN(n3943) );
  NAND2_X1 U4844 ( .A1(n4290), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3942)
         );
  NAND4_X1 U4845 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n4741)
         );
  XOR2_X1 U4846 ( .A(n4942), .B(n3946), .Z(n6166) );
  INV_X1 U4847 ( .A(n6166), .ZN(n3961) );
  AOI22_X1 U4848 ( .A1(n4273), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4849 ( .A1(n3442), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4850 ( .A1(n4271), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4851 ( .A1(n4263), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3947) );
  NAND4_X1 U4852 ( .A1(n3950), .A2(n3949), .A3(n3948), .A4(n3947), .ZN(n3956)
         );
  AOI22_X1 U4853 ( .A1(n4262), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4261), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4854 ( .A1(n4272), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3450), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4855 ( .A1(n3443), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4856 ( .A1(n4099), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3951) );
  NAND4_X1 U4857 ( .A1(n3954), .A2(n3953), .A3(n3952), .A4(n3951), .ZN(n3955)
         );
  OAI21_X1 U4858 ( .B1(n3956), .B2(n3955), .A(n4043), .ZN(n3959) );
  NAND2_X1 U4859 ( .A1(n4291), .A2(EAX_REG_9__SCAN_IN), .ZN(n3958) );
  NAND2_X1 U4860 ( .A1(n4290), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3957)
         );
  NAND3_X1 U4861 ( .A1(n3959), .A2(n3958), .A3(n3957), .ZN(n3960) );
  AOI21_X1 U4862 ( .B1(n3961), .B2(n4834), .A(n3960), .ZN(n4737) );
  NAND2_X1 U4863 ( .A1(n3962), .A2(n6975), .ZN(n3964) );
  INV_X1 U4864 ( .A(n3990), .ZN(n3963) );
  NAND2_X1 U4865 ( .A1(n3964), .A2(n3963), .ZN(n5317) );
  AOI22_X1 U4866 ( .A1(n4273), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4867 ( .A1(n4272), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4868 ( .A1(n4261), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4869 ( .A1(n4172), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3965) );
  NAND4_X1 U4870 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(n3974)
         );
  AOI22_X1 U4871 ( .A1(n3450), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4872 ( .A1(n4262), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4873 ( .A1(n3443), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4263), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4874 ( .A1(n4099), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3969) );
  NAND4_X1 U4875 ( .A1(n3972), .A2(n3971), .A3(n3970), .A4(n3969), .ZN(n3973)
         );
  OAI21_X1 U4876 ( .B1(n3974), .B2(n3973), .A(n4043), .ZN(n3977) );
  NAND2_X1 U4877 ( .A1(n4291), .A2(EAX_REG_10__SCAN_IN), .ZN(n3976) );
  NAND2_X1 U4878 ( .A1(n4290), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3975)
         );
  NAND3_X1 U4879 ( .A1(n3977), .A2(n3976), .A3(n3975), .ZN(n3978) );
  AOI21_X1 U4880 ( .B1(n5317), .B2(n4834), .A(n3978), .ZN(n4995) );
  AOI22_X1 U4881 ( .A1(n4273), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4882 ( .A1(n4261), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4883 ( .A1(n4272), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4884 ( .A1(n4263), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3980) );
  NAND4_X1 U4885 ( .A1(n3983), .A2(n3982), .A3(n3981), .A4(n3980), .ZN(n3989)
         );
  AOI22_X1 U4886 ( .A1(n3450), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4887 ( .A1(n4262), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4888 ( .A1(n3443), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4889 ( .A1(n4099), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3984) );
  NAND4_X1 U4890 ( .A1(n3987), .A2(n3986), .A3(n3985), .A4(n3984), .ZN(n3988)
         );
  OAI21_X1 U4891 ( .B1(n3989), .B2(n3988), .A(n4043), .ZN(n3993) );
  XOR2_X1 U4892 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3990), .Z(n6275) );
  INV_X1 U4893 ( .A(n6275), .ZN(n5329) );
  AOI22_X1 U4894 ( .A1(n4834), .A2(n5329), .B1(n4290), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3992) );
  NAND2_X1 U4895 ( .A1(n4291), .A2(EAX_REG_11__SCAN_IN), .ZN(n3991) );
  AOI22_X1 U4896 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4262), .B1(n4272), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4897 ( .A1(n4273), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4263), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4898 ( .A1(n3443), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4899 ( .A1(n3450), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3994) );
  NAND4_X1 U4900 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), .ZN(n4003)
         );
  AOI22_X1 U4901 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3442), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4902 ( .A1(n4261), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4903 ( .A1(n4264), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4904 ( .A1(n4172), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3998) );
  NAND4_X1 U4905 ( .A1(n4001), .A2(n4000), .A3(n3999), .A4(n3998), .ZN(n4002)
         );
  NOR2_X1 U4906 ( .A1(n4003), .A2(n4002), .ZN(n4007) );
  XNOR2_X1 U4907 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n4004), .ZN(n6152)
         );
  AOI22_X1 U4908 ( .A1(n4834), .A2(n6152), .B1(n4290), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n4006) );
  NAND2_X1 U4909 ( .A1(n4291), .A2(EAX_REG_12__SCAN_IN), .ZN(n4005) );
  OAI211_X1 U4910 ( .C1(n4059), .C2(n4007), .A(n4006), .B(n4005), .ZN(n5334)
         );
  NAND2_X1 U4911 ( .A1(n5229), .A2(n5334), .ZN(n4012) );
  NAND2_X1 U4912 ( .A1(n4291), .A2(EAX_REG_13__SCAN_IN), .ZN(n4010) );
  OAI21_X1 U4913 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n4008), .A(n4030), 
        .ZN(n6148) );
  AOI22_X1 U4914 ( .A1(n4834), .A2(n6148), .B1(n4290), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n4009) );
  NAND2_X1 U4915 ( .A1(n4010), .A2(n4009), .ZN(n4013) );
  INV_X1 U4916 ( .A(n4013), .ZN(n4011) );
  NAND2_X1 U4917 ( .A1(n4012), .A2(n4011), .ZN(n4015) );
  INV_X1 U4918 ( .A(n4012), .ZN(n4014) );
  NAND2_X1 U4919 ( .A1(n4015), .A2(n4029), .ZN(n5376) );
  INV_X1 U4920 ( .A(n5376), .ZN(n4028) );
  AOI22_X1 U4921 ( .A1(n3443), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4922 ( .A1(n4262), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4923 ( .A1(n4264), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4924 ( .A1(n4273), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U4925 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4025)
         );
  AOI22_X1 U4926 ( .A1(n4272), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3495), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4927 ( .A1(n4261), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4928 ( .A1(n4263), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4929 ( .A1(n4099), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4020) );
  NAND4_X1 U4930 ( .A1(n4023), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(n4024)
         );
  OR2_X1 U4931 ( .A1(n4025), .A2(n4024), .ZN(n4026) );
  NAND2_X1 U4932 ( .A1(n4043), .A2(n4026), .ZN(n5377) );
  NAND2_X1 U4933 ( .A1(n4028), .A2(n4027), .ZN(n5379) );
  XOR2_X1 U4934 ( .A(n4031), .B(n4030), .Z(n6131) );
  AOI22_X1 U4935 ( .A1(n4273), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4936 ( .A1(n3442), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U4937 ( .A1(n3495), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4938 ( .A1(n4263), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4032) );
  NAND4_X1 U4939 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(n4041)
         );
  AOI22_X1 U4940 ( .A1(n3443), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4262), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4941 ( .A1(n4272), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4942 ( .A1(n4261), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4943 ( .A1(n4099), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4036) );
  NAND4_X1 U4944 ( .A1(n4039), .A2(n4038), .A3(n4037), .A4(n4036), .ZN(n4040)
         );
  OR2_X1 U4945 ( .A1(n4041), .A2(n4040), .ZN(n4042) );
  AOI22_X1 U4946 ( .A1(n4043), .A2(n4042), .B1(n4290), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U4947 ( .A1(n4291), .A2(EAX_REG_14__SCAN_IN), .ZN(n4044) );
  OAI211_X1 U4948 ( .C1(n6131), .C2(n4289), .A(n4045), .B(n4044), .ZN(n5429)
         );
  AOI22_X1 U4949 ( .A1(n4262), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4950 ( .A1(n4273), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4261), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U4951 ( .A1(n4062), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U4952 ( .A1(n4270), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4046) );
  NAND4_X1 U4953 ( .A1(n4049), .A2(n4048), .A3(n4047), .A4(n4046), .ZN(n4055)
         );
  AOI22_X1 U4954 ( .A1(n4264), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U4955 ( .A1(n3443), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3495), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4052) );
  AOI22_X1 U4956 ( .A1(n4271), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4957 ( .A1(n4263), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4050) );
  NAND4_X1 U4958 ( .A1(n4053), .A2(n4052), .A3(n4051), .A4(n4050), .ZN(n4054)
         );
  NOR2_X1 U4959 ( .A1(n4055), .A2(n4054), .ZN(n4060) );
  XNOR2_X1 U4960 ( .A(n4056), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5798)
         );
  NAND2_X1 U4961 ( .A1(n5798), .A2(n4834), .ZN(n4058) );
  AOI22_X1 U4962 ( .A1(n4291), .A2(EAX_REG_15__SCAN_IN), .B1(n4290), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4057) );
  OAI211_X1 U4963 ( .C1(n4060), .C2(n4059), .A(n4058), .B(n4057), .ZN(n5404)
         );
  AOI21_X1 U4964 ( .B1(n7050), .B2(n4061), .A(n4078), .ZN(n6127) );
  OR2_X1 U4965 ( .A1(n6127), .A2(n4289), .ZN(n4077) );
  AOI22_X1 U4966 ( .A1(n4273), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U4967 ( .A1(n4272), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U4968 ( .A1(n4261), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U4969 ( .A1(n4263), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4063) );
  NAND4_X1 U4970 ( .A1(n4066), .A2(n4065), .A3(n4064), .A4(n4063), .ZN(n4072)
         );
  AOI22_X1 U4971 ( .A1(n4262), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U4972 ( .A1(n4271), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4069) );
  AOI22_X1 U4973 ( .A1(n3443), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U4974 ( .A1(n3495), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4067) );
  NAND4_X1 U4975 ( .A1(n4070), .A2(n4069), .A3(n4068), .A4(n4067), .ZN(n4071)
         );
  NOR2_X1 U4976 ( .A1(n4072), .A2(n4071), .ZN(n4074) );
  AOI22_X1 U4977 ( .A1(n4291), .A2(EAX_REG_16__SCAN_IN), .B1(n4290), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4073) );
  OAI21_X1 U4978 ( .B1(n4286), .B2(n4074), .A(n4073), .ZN(n4075) );
  INV_X1 U4979 ( .A(n4075), .ZN(n4076) );
  XNOR2_X1 U4980 ( .A(n4078), .B(n6116), .ZN(n6118) );
  AOI22_X1 U4981 ( .A1(n4264), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U4982 ( .A1(n3443), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3495), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U4983 ( .A1(n4261), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U4984 ( .A1(n4172), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4079) );
  NAND4_X1 U4985 ( .A1(n4082), .A2(n4081), .A3(n4080), .A4(n4079), .ZN(n4088)
         );
  AOI22_X1 U4986 ( .A1(n4273), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4262), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U4987 ( .A1(n4263), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U4988 ( .A1(n4270), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U4989 ( .A1(n4272), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4083) );
  NAND4_X1 U4990 ( .A1(n4086), .A2(n4085), .A3(n4084), .A4(n4083), .ZN(n4087)
         );
  NOR2_X1 U4991 ( .A1(n4088), .A2(n4087), .ZN(n4091) );
  NOR2_X1 U4992 ( .A1(n6116), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4089) );
  AOI21_X1 U4993 ( .B1(n4291), .B2(EAX_REG_17__SCAN_IN), .A(n4089), .ZN(n4090)
         );
  OAI21_X1 U4994 ( .B1(n4286), .B2(n4091), .A(n4090), .ZN(n4092) );
  NAND2_X1 U4995 ( .A1(n4092), .A2(n4289), .ZN(n4093) );
  NAND2_X1 U4996 ( .A1(n4094), .A2(n4093), .ZN(n6056) );
  AOI22_X1 U4997 ( .A1(n4273), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4263), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U4998 ( .A1(n3443), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U4999 ( .A1(n4262), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5000 ( .A1(n3450), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3841), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4095) );
  NAND4_X1 U5001 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(n4105)
         );
  AOI22_X1 U5002 ( .A1(n4261), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5003 ( .A1(n3442), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5004 ( .A1(n4264), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5005 ( .A1(n4099), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4100) );
  NAND4_X1 U5006 ( .A1(n4103), .A2(n4102), .A3(n4101), .A4(n4100), .ZN(n4104)
         );
  NOR2_X1 U5007 ( .A1(n4105), .A2(n4104), .ZN(n4109) );
  NAND2_X1 U5008 ( .A1(n6737), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4106)
         );
  NAND2_X1 U5009 ( .A1(n4289), .A2(n4106), .ZN(n4107) );
  AOI21_X1 U5010 ( .B1(n4291), .B2(EAX_REG_18__SCAN_IN), .A(n4107), .ZN(n4108)
         );
  OAI21_X1 U5011 ( .B1(n4286), .B2(n4109), .A(n4108), .ZN(n4116) );
  INV_X1 U5012 ( .A(n4130), .ZN(n4114) );
  INV_X1 U5013 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4112) );
  INV_X1 U5014 ( .A(n4110), .ZN(n4111) );
  NAND2_X1 U5015 ( .A1(n4112), .A2(n4111), .ZN(n4113) );
  NAND2_X1 U5016 ( .A1(n4114), .A2(n4113), .ZN(n6111) );
  NAND2_X1 U5017 ( .A1(n4116), .A2(n4115), .ZN(n5670) );
  AOI22_X1 U5018 ( .A1(n4273), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5019 ( .A1(n4262), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5020 ( .A1(n4272), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4062), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4118) );
  AOI22_X1 U5021 ( .A1(n4263), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4117) );
  NAND4_X1 U5022 ( .A1(n4120), .A2(n4119), .A3(n4118), .A4(n4117), .ZN(n4126)
         );
  AOI22_X1 U5023 ( .A1(n4261), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3450), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5024 ( .A1(n4271), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5025 ( .A1(n3443), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5026 ( .A1(n4099), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4121) );
  NAND4_X1 U5027 ( .A1(n4124), .A2(n4123), .A3(n4122), .A4(n4121), .ZN(n4125)
         );
  NOR2_X1 U5028 ( .A1(n4126), .A2(n4125), .ZN(n4129) );
  INV_X1 U5029 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n6957) );
  OAI21_X1 U5030 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6957), .A(n4289), .ZN(
        n4127) );
  AOI21_X1 U5031 ( .B1(n4291), .B2(EAX_REG_19__SCAN_IN), .A(n4127), .ZN(n4128)
         );
  OAI21_X1 U5032 ( .B1(n4286), .B2(n4129), .A(n4128), .ZN(n4133) );
  NOR2_X1 U5033 ( .A1(n4130), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4131)
         );
  NOR2_X1 U5034 ( .A1(n4149), .A2(n4131), .ZN(n6022) );
  NAND2_X1 U5035 ( .A1(n6022), .A2(n4834), .ZN(n4132) );
  NAND2_X1 U5036 ( .A1(n4133), .A2(n4132), .ZN(n5660) );
  NAND2_X1 U5037 ( .A1(n5657), .A2(n4134), .ZN(n5600) );
  AOI22_X1 U5038 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4262), .B1(n4272), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U5039 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4273), .B1(n4261), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5040 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3442), .B1(n3495), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5041 ( .A1(n3435), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4135) );
  NAND4_X1 U5042 ( .A1(n4138), .A2(n4137), .A3(n4136), .A4(n4135), .ZN(n4144)
         );
  AOI22_X1 U5043 ( .A1(n4264), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5044 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4270), .B1(n4172), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U5045 ( .A1(n3443), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5046 ( .A1(n4263), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4139) );
  NAND4_X1 U5047 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(n4143)
         );
  NOR2_X1 U5048 ( .A1(n4144), .A2(n4143), .ZN(n4148) );
  INV_X1 U5049 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6738) );
  OAI21_X1 U5050 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6738), .A(n6737), 
        .ZN(n4145) );
  INV_X1 U5051 ( .A(n4145), .ZN(n4146) );
  AOI21_X1 U5052 ( .B1(n4291), .B2(EAX_REG_20__SCAN_IN), .A(n4146), .ZN(n4147)
         );
  OAI21_X1 U5053 ( .B1(n4286), .B2(n4148), .A(n4147), .ZN(n4151) );
  OAI21_X1 U5054 ( .B1(n4149), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n4165), 
        .ZN(n5773) );
  OR2_X1 U5055 ( .A1(n5773), .A2(n4289), .ZN(n4150) );
  NAND2_X1 U5056 ( .A1(n4151), .A2(n4150), .ZN(n5601) );
  AOI22_X1 U5057 ( .A1(n3443), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5058 ( .A1(n4261), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U5059 ( .A1(n4262), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5060 ( .A1(n4099), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4152) );
  NAND4_X1 U5061 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4161)
         );
  AOI22_X1 U5062 ( .A1(n4264), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3450), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5063 ( .A1(n4272), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5064 ( .A1(n4273), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U5065 ( .A1(n4263), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4156) );
  NAND4_X1 U5066 ( .A1(n4159), .A2(n4158), .A3(n4157), .A4(n4156), .ZN(n4160)
         );
  NOR2_X1 U5067 ( .A1(n4161), .A2(n4160), .ZN(n4164) );
  AOI21_X1 U5068 ( .B1(n5766), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4162) );
  AOI21_X1 U5069 ( .B1(n4291), .B2(EAX_REG_21__SCAN_IN), .A(n4162), .ZN(n4163)
         );
  OAI21_X1 U5070 ( .B1(n4286), .B2(n4164), .A(n4163), .ZN(n4167) );
  XNOR2_X1 U5071 ( .A(n4165), .B(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6011)
         );
  NAND2_X1 U5072 ( .A1(n6011), .A2(n4834), .ZN(n4166) );
  AOI22_X1 U5073 ( .A1(n3443), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4272), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U5074 ( .A1(n4262), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4271), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5075 ( .A1(n4261), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5076 ( .A1(n3442), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4168) );
  NAND4_X1 U5077 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4178)
         );
  AOI22_X1 U5078 ( .A1(n4264), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3495), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5079 ( .A1(n4273), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5080 ( .A1(n3435), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4172), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5081 ( .A1(n4263), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3544), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4173) );
  NAND4_X1 U5082 ( .A1(n4176), .A2(n4175), .A3(n4174), .A4(n4173), .ZN(n4177)
         );
  NOR2_X1 U5083 ( .A1(n4178), .A2(n4177), .ZN(n4182) );
  OAI21_X1 U5084 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6738), .A(n6737), 
        .ZN(n4179) );
  INV_X1 U5085 ( .A(n4179), .ZN(n4180) );
  AOI21_X1 U5086 ( .B1(n4291), .B2(EAX_REG_22__SCAN_IN), .A(n4180), .ZN(n4181)
         );
  OAI21_X1 U5087 ( .B1(n4286), .B2(n4182), .A(n4181), .ZN(n4187) );
  NOR2_X1 U5088 ( .A1(n4183), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4184)
         );
  OR2_X1 U5089 ( .A1(n4193), .A2(n4184), .ZN(n5760) );
  INV_X1 U5090 ( .A(n5760), .ZN(n4185) );
  NAND2_X1 U5091 ( .A1(n4185), .A2(n4834), .ZN(n4186) );
  XNOR2_X1 U5092 ( .A(n4189), .B(n4188), .ZN(n4192) );
  INV_X1 U5093 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6009) );
  OAI21_X1 U5094 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6009), .A(n4289), .ZN(
        n4190) );
  AOI21_X1 U5095 ( .B1(n4291), .B2(EAX_REG_23__SCAN_IN), .A(n4190), .ZN(n4191)
         );
  OAI21_X1 U5096 ( .B1(n4286), .B2(n4192), .A(n4191), .ZN(n4195) );
  XNOR2_X1 U5097 ( .A(n4193), .B(n6009), .ZN(n6000) );
  NAND2_X1 U5098 ( .A1(n6000), .A2(n4834), .ZN(n4194) );
  INV_X1 U5099 ( .A(n4196), .ZN(n4197) );
  XNOR2_X1 U5100 ( .A(n4198), .B(n4197), .ZN(n4203) );
  INV_X1 U5101 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4199) );
  XNOR2_X1 U5102 ( .A(n4200), .B(n4199), .ZN(n5994) );
  AOI22_X1 U5103 ( .A1(n4291), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n4290), .ZN(n4201) );
  OAI21_X1 U5104 ( .B1(n5994), .B2(n4289), .A(n4201), .ZN(n4202) );
  AOI21_X1 U5105 ( .B1(n4226), .B2(n4203), .A(n4202), .ZN(n5632) );
  XOR2_X1 U5106 ( .A(n4205), .B(n4204), .Z(n4208) );
  INV_X1 U5107 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U5108 ( .A1(n4291), .A2(EAX_REG_25__SCAN_IN), .ZN(n4206) );
  OAI211_X1 U5109 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n5737), .A(n4206), .B(
        n4289), .ZN(n4207) );
  AOI21_X1 U5110 ( .B1(n4208), .B2(n4226), .A(n4207), .ZN(n4209) );
  INV_X1 U5111 ( .A(n4209), .ZN(n4211) );
  XNOR2_X1 U5112 ( .A(n4219), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5983)
         );
  NAND2_X1 U5113 ( .A1(n5983), .A2(n4834), .ZN(n4210) );
  NAND2_X1 U5114 ( .A1(n4211), .A2(n4210), .ZN(n5628) );
  INV_X1 U5115 ( .A(n4212), .ZN(n4213) );
  XNOR2_X1 U5116 ( .A(n4214), .B(n4213), .ZN(n4215) );
  NAND2_X1 U5117 ( .A1(n4215), .A2(n4226), .ZN(n4223) );
  NAND2_X1 U5118 ( .A1(n6737), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4216)
         );
  NAND2_X1 U5119 ( .A1(n4289), .A2(n4216), .ZN(n4217) );
  AOI21_X1 U5120 ( .B1(n4291), .B2(EAX_REG_26__SCAN_IN), .A(n4217), .ZN(n4222)
         );
  INV_X1 U5121 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4218) );
  OAI21_X1 U5122 ( .B1(n4219), .B2(n5737), .A(n4218), .ZN(n4220) );
  NAND2_X1 U5123 ( .A1(n4220), .A2(n4229), .ZN(n5981) );
  NOR2_X1 U5124 ( .A1(n5981), .A2(n4289), .ZN(n4221) );
  AOI21_X1 U5125 ( .B1(n4223), .B2(n4222), .A(n4221), .ZN(n5619) );
  XOR2_X1 U5126 ( .A(n4225), .B(n4224), .Z(n4227) );
  NAND2_X1 U5127 ( .A1(n4227), .A2(n4226), .ZN(n4232) );
  INV_X1 U5128 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n7026) );
  NOR2_X1 U5129 ( .A1(n7026), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4228) );
  AOI211_X1 U5130 ( .C1(n4291), .C2(EAX_REG_27__SCAN_IN), .A(n4834), .B(n4228), 
        .ZN(n4231) );
  NAND2_X1 U5131 ( .A1(n4229), .A2(n7026), .ZN(n4230) );
  AOI22_X1 U5132 ( .A1(n4232), .A2(n4231), .B1(n4834), .B2(n5726), .ZN(n5572)
         );
  NAND2_X1 U5133 ( .A1(n4233), .A2(n6958), .ZN(n4234) );
  NAND2_X1 U5134 ( .A1(n4260), .A2(n4234), .ZN(n5717) );
  XNOR2_X1 U5135 ( .A(n4236), .B(n4235), .ZN(n4239) );
  OAI21_X1 U5136 ( .B1(n6738), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n6737), 
        .ZN(n4238) );
  NAND2_X1 U5137 ( .A1(n4291), .A2(EAX_REG_28__SCAN_IN), .ZN(n4237) );
  OAI211_X1 U5138 ( .C1(n4239), .C2(n4286), .A(n4238), .B(n4237), .ZN(n4240)
         );
  NAND3_X1 U5139 ( .A1(n6743), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6647) );
  INV_X1 U5140 ( .A(n6647), .ZN(n4243) );
  NOR2_X1 U5141 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6486) );
  INV_X1 U5142 ( .A(n6486), .ZN(n6535) );
  NAND2_X1 U5143 ( .A1(n6535), .A2(n4250), .ZN(n6746) );
  NAND2_X1 U5144 ( .A1(n6746), .A2(n6743), .ZN(n4246) );
  NAND2_X1 U5145 ( .A1(n6743), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4248) );
  NAND2_X1 U5146 ( .A1(n6738), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4247) );
  AND2_X1 U5147 ( .A1(n4248), .A2(n4247), .ZN(n4358) );
  INV_X1 U5148 ( .A(n4358), .ZN(n4249) );
  NAND2_X1 U5149 ( .A1(n6276), .A2(n5552), .ZN(n4253) );
  OR2_X1 U5150 ( .A1(n4250), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6388) );
  INV_X2 U5151 ( .A(n6388), .ZN(n6353) );
  NAND2_X1 U5152 ( .A1(n6353), .A2(REIP_REG_29__SCAN_IN), .ZN(n5842) );
  OAI21_X1 U5153 ( .B1(n6063), .B2(n4259), .A(n5842), .ZN(n4251) );
  INV_X1 U5154 ( .A(n4251), .ZN(n4252) );
  OAI211_X1 U5155 ( .C1(n5851), .C2(n6294), .A(n4254), .B(n3260), .ZN(U2957)
         );
  INV_X1 U5156 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5827) );
  AND2_X1 U5157 ( .A1(n6910), .A2(n5827), .ZN(n4255) );
  NAND2_X1 U5158 ( .A1(n5709), .A2(n4255), .ZN(n4257) );
  NAND2_X1 U5159 ( .A1(n5698), .A2(n3265), .ZN(n4256) );
  NAND2_X1 U5160 ( .A1(n4257), .A2(n4256), .ZN(n4258) );
  XNOR2_X1 U5161 ( .A(n4258), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5833)
         );
  XNOR2_X1 U5162 ( .A(n4294), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5703)
         );
  AOI22_X1 U5163 ( .A1(n4262), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4261), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4269) );
  AOI22_X1 U5164 ( .A1(n4264), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4263), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4268) );
  AOI22_X1 U5165 ( .A1(n3495), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4265), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U5166 ( .A1(n4099), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4266) );
  NAND4_X1 U5167 ( .A1(n4269), .A2(n4268), .A3(n4267), .A4(n4266), .ZN(n4279)
         );
  AOI22_X1 U5168 ( .A1(n3443), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3442), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4277) );
  AOI22_X1 U5169 ( .A1(n4271), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4270), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4276) );
  AOI22_X1 U5170 ( .A1(n4272), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3435), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4275) );
  AOI22_X1 U5171 ( .A1(n4273), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3589), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4274) );
  NAND4_X1 U5172 ( .A1(n4277), .A2(n4276), .A3(n4275), .A4(n4274), .ZN(n4278)
         );
  NOR2_X1 U5173 ( .A1(n4279), .A2(n4278), .ZN(n4283) );
  NOR2_X1 U5174 ( .A1(n4281), .A2(n4280), .ZN(n4282) );
  XOR2_X1 U5175 ( .A(n4283), .B(n4282), .Z(n4287) );
  AOI21_X1 U5176 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6737), .A(n4834), 
        .ZN(n4285) );
  NAND2_X1 U5177 ( .A1(n4291), .A2(EAX_REG_30__SCAN_IN), .ZN(n4284) );
  OAI211_X1 U5178 ( .C1(n4287), .C2(n4286), .A(n4285), .B(n4284), .ZN(n4288)
         );
  OAI21_X1 U5179 ( .B1(n4289), .B2(n5703), .A(n4288), .ZN(n5528) );
  AOI22_X1 U5180 ( .A1(n4291), .A2(EAX_REG_31__SCAN_IN), .B1(n4290), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4292) );
  NAND2_X1 U5181 ( .A1(n4294), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4295)
         );
  XNOR2_X1 U5182 ( .A(n4295), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4842)
         );
  INV_X1 U5183 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U5184 ( .A1(n6353), .A2(REIP_REG_31__SCAN_IN), .ZN(n5818) );
  OAI21_X1 U5185 ( .B1(n6063), .B2(n6832), .A(n5818), .ZN(n4296) );
  OAI211_X1 U5186 ( .C1(n5833), .C2(n6294), .A(n4298), .B(n4297), .ZN(U2955)
         );
  NOR2_X1 U5187 ( .A1(n4300), .A2(n4845), .ZN(n4301) );
  NAND2_X1 U5188 ( .A1(n4299), .A2(n4301), .ZN(n4548) );
  OR3_X1 U5189 ( .A1(n4304), .A2(n4303), .A3(n4302), .ZN(n4305) );
  NAND2_X1 U5190 ( .A1(n4306), .A2(n4305), .ZN(n4308) );
  NAND2_X1 U5191 ( .A1(n4308), .A2(n4307), .ZN(n4555) );
  INV_X1 U5192 ( .A(n4555), .ZN(n4330) );
  NOR2_X1 U5193 ( .A1(n4548), .A2(n4330), .ZN(n4312) );
  INV_X1 U5194 ( .A(n4313), .ZN(n4329) );
  NOR2_X1 U5195 ( .A1(n4312), .A2(n4329), .ZN(n4309) );
  AOI21_X1 U5196 ( .B1(n4612), .B2(n4839), .A(n4309), .ZN(n4318) );
  AND2_X1 U5197 ( .A1(n4318), .A2(n6640), .ZN(n4311) );
  INV_X1 U5198 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6969) );
  AND2_X1 U5199 ( .A1(n6530), .A2(n5452), .ZN(n5166) );
  NAND2_X1 U5200 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5166), .ZN(n4310) );
  OAI21_X1 U5201 ( .B1(n4311), .B2(n6969), .A(n4310), .ZN(U2790) );
  INV_X1 U5202 ( .A(n4336), .ZN(n4340) );
  OR2_X1 U5203 ( .A1(n4364), .A2(n5166), .ZN(n4337) );
  AOI21_X1 U5204 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n4340), .A(n4337), .ZN(
        n4315) );
  INV_X1 U5205 ( .A(n4315), .ZN(U2788) );
  NAND2_X1 U5206 ( .A1(n4857), .A2(n4603), .ZN(n4853) );
  NAND2_X1 U5207 ( .A1(n4854), .A2(n4853), .ZN(n4341) );
  INV_X1 U5208 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4316) );
  NAND2_X1 U5209 ( .A1(n3192), .A2(n4316), .ZN(n6655) );
  NAND2_X1 U5210 ( .A1(n4341), .A2(n6655), .ZN(n6740) );
  INV_X1 U5211 ( .A(READY_N), .ZN(n4599) );
  NAND2_X1 U5212 ( .A1(n6740), .A2(n4599), .ZN(n4317) );
  NAND2_X1 U5213 ( .A1(n4318), .A2(n4317), .ZN(n6618) );
  AND2_X1 U5214 ( .A1(n6618), .A2(n6640), .ZN(n6091) );
  INV_X1 U5215 ( .A(MORE_REG_SCAN_IN), .ZN(n4335) );
  AOI22_X1 U5216 ( .A1(n4319), .A2(n5662), .B1(n4607), .B2(n4647), .ZN(n4324)
         );
  AND2_X1 U5217 ( .A1(n4321), .A2(n4320), .ZN(n4545) );
  OR2_X1 U5218 ( .A1(n4853), .A2(n4607), .ZN(n4550) );
  NAND2_X1 U5219 ( .A1(n5497), .A2(n4550), .ZN(n4322) );
  NAND2_X1 U5220 ( .A1(n4322), .A2(n3516), .ZN(n4323) );
  AND3_X1 U5221 ( .A1(n4324), .A2(n4545), .A3(n4323), .ZN(n4325) );
  NAND2_X1 U5222 ( .A1(n4326), .A2(n4325), .ZN(n4523) );
  AOI21_X1 U5223 ( .B1(n4327), .B2(n4563), .A(n4845), .ZN(n4328) );
  NOR2_X1 U5224 ( .A1(n4523), .A2(n4328), .ZN(n4620) );
  NOR2_X1 U5225 ( .A1(n6594), .A2(n4873), .ZN(n4611) );
  NAND2_X1 U5226 ( .A1(n4620), .A2(n4611), .ZN(n4544) );
  OR2_X1 U5227 ( .A1(n4547), .A2(n4839), .ZN(n4556) );
  NAND2_X1 U5228 ( .A1(n6615), .A2(n4556), .ZN(n4618) );
  OAI21_X1 U5229 ( .B1(n4329), .B2(n4618), .A(n4612), .ZN(n4333) );
  INV_X1 U5230 ( .A(n4548), .ZN(n4331) );
  NAND2_X1 U5231 ( .A1(n4331), .A2(n4330), .ZN(n4332) );
  OAI211_X1 U5232 ( .C1(n4612), .C2(n4544), .A(n4333), .B(n4332), .ZN(n6614)
         );
  NAND2_X1 U5233 ( .A1(n6091), .A2(n6614), .ZN(n4334) );
  OAI21_X1 U5234 ( .B1(n6091), .B2(n4335), .A(n4334), .ZN(U3471) );
  INV_X1 U5235 ( .A(n4341), .ZN(n4338) );
  OAI22_X1 U5236 ( .A1(n4838), .A2(n4338), .B1(READREQUEST_REG_SCAN_IN), .B2(
        n4337), .ZN(n4339) );
  OAI21_X1 U5237 ( .B1(n4341), .B2(n4340), .A(n4339), .ZN(U3474) );
  INV_X1 U5238 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4405) );
  NOR2_X1 U5239 ( .A1(n4548), .A2(n4873), .ZN(n6598) );
  NAND2_X1 U5240 ( .A1(n4342), .A2(n6739), .ZN(n4625) );
  INV_X1 U5241 ( .A(n4625), .ZN(n6626) );
  INV_X1 U5242 ( .A(n6655), .ZN(n4343) );
  OAI211_X1 U5243 ( .C1(n6598), .C2(n6626), .A(n4343), .B(n6640), .ZN(n4344)
         );
  NOR2_X1 U5244 ( .A1(n4612), .A2(n4344), .ZN(n6241) );
  NAND2_X1 U5245 ( .A1(n6241), .A2(n4845), .ZN(n4484) );
  NOR2_X1 U5246 ( .A1(n5452), .A2(n6737), .ZN(n4591) );
  AOI22_X1 U5247 ( .A1(n6747), .A2(UWORD_REG_9__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4345) );
  OAI21_X1 U5248 ( .B1(n4405), .B2(n4484), .A(n4345), .ZN(U2898) );
  INV_X1 U5249 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4401) );
  AOI22_X1 U5250 ( .A1(n6747), .A2(UWORD_REG_10__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4346) );
  OAI21_X1 U5251 ( .B1(n4401), .B2(n4484), .A(n4346), .ZN(U2897) );
  INV_X1 U5252 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6972) );
  AOI22_X1 U5253 ( .A1(n6747), .A2(UWORD_REG_8__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4347) );
  OAI21_X1 U5254 ( .B1(n6972), .B2(n4484), .A(n4347), .ZN(U2899) );
  INV_X1 U5255 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4377) );
  AOI22_X1 U5256 ( .A1(n6747), .A2(UWORD_REG_12__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4348) );
  OAI21_X1 U5257 ( .B1(n4377), .B2(n4484), .A(n4348), .ZN(U2895) );
  INV_X1 U5258 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4373) );
  AOI22_X1 U5259 ( .A1(n6747), .A2(UWORD_REG_13__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4349) );
  OAI21_X1 U5260 ( .B1(n4373), .B2(n4484), .A(n4349), .ZN(U2894) );
  INV_X1 U5261 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6925) );
  AOI22_X1 U5262 ( .A1(n6747), .A2(UWORD_REG_11__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4350) );
  OAI21_X1 U5263 ( .B1(n6925), .B2(n4484), .A(n4350), .ZN(U2896) );
  INV_X1 U5264 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4416) );
  AOI22_X1 U5265 ( .A1(n6747), .A2(UWORD_REG_14__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4351) );
  OAI21_X1 U5266 ( .B1(n4416), .B2(n4484), .A(n4351), .ZN(U2893) );
  NAND2_X1 U5267 ( .A1(n4352), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4354) );
  NAND2_X1 U5268 ( .A1(n4354), .A2(n4353), .ZN(n4356) );
  NAND2_X1 U5269 ( .A1(n4356), .A2(n4355), .ZN(n5236) );
  INV_X1 U5270 ( .A(n6294), .ZN(n6303) );
  XNOR2_X1 U5271 ( .A(n4357), .B(n5451), .ZN(n5961) );
  NAND2_X1 U5272 ( .A1(n6303), .A2(n5961), .ZN(n4362) );
  NAND2_X1 U5273 ( .A1(n4358), .A2(n6063), .ZN(n4360) );
  NAND2_X1 U5274 ( .A1(n6353), .A2(REIP_REG_0__SCAN_IN), .ZN(n5958) );
  INV_X1 U5275 ( .A(n5958), .ZN(n4359) );
  AOI21_X1 U5276 ( .B1(PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4360), .A(n4359), 
        .ZN(n4361) );
  OAI211_X1 U5277 ( .C1(n5236), .C2(n6292), .A(n4362), .B(n4361), .ZN(U2986)
         );
  NAND2_X1 U5278 ( .A1(n4364), .A2(n4873), .ZN(n4420) );
  INV_X1 U5279 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4473) );
  AND2_X1 U5280 ( .A1(n4603), .A2(n4599), .ZN(n4363) );
  NAND2_X1 U5281 ( .A1(n4364), .A2(n4363), .ZN(n4645) );
  NAND2_X1 U5282 ( .A1(n4418), .A2(DATAI_4_), .ZN(n4410) );
  OAI21_X1 U5283 ( .B1(n6739), .B2(n4599), .A(n4364), .ZN(n4371) );
  NAND2_X1 U5284 ( .A1(n4371), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4365) );
  OAI211_X1 U5285 ( .C1(n4415), .C2(n4473), .A(n4410), .B(n4365), .ZN(U2928)
         );
  INV_X1 U5286 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4475) );
  NAND2_X1 U5287 ( .A1(n4418), .A2(DATAI_6_), .ZN(n4398) );
  NAND2_X1 U5288 ( .A1(n4371), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4366) );
  OAI211_X1 U5289 ( .C1(n4415), .C2(n4475), .A(n4398), .B(n4366), .ZN(U2930)
         );
  INV_X1 U5290 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4479) );
  NAND2_X1 U5291 ( .A1(n4418), .A2(DATAI_3_), .ZN(n4394) );
  NAND2_X1 U5292 ( .A1(n4371), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4367) );
  OAI211_X1 U5293 ( .C1(n4479), .C2(n4415), .A(n4394), .B(n4367), .ZN(U2927)
         );
  INV_X1 U5294 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U5295 ( .A1(n4418), .A2(DATAI_5_), .ZN(n4381) );
  NAND2_X1 U5296 ( .A1(n4371), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4368) );
  OAI211_X1 U5297 ( .C1(n4471), .C2(n4415), .A(n4381), .B(n4368), .ZN(U2929)
         );
  INV_X1 U5298 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4477) );
  NAND2_X1 U5299 ( .A1(n4418), .A2(DATAI_7_), .ZN(n4396) );
  NAND2_X1 U5300 ( .A1(n4371), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4369) );
  OAI211_X1 U5301 ( .C1(n4477), .C2(n4415), .A(n4396), .B(n4369), .ZN(U2931)
         );
  INV_X1 U5302 ( .A(EAX_REG_18__SCAN_IN), .ZN(n7029) );
  NAND2_X1 U5303 ( .A1(n4418), .A2(DATAI_2_), .ZN(n4386) );
  NAND2_X1 U5304 ( .A1(n4371), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4370) );
  OAI211_X1 U5305 ( .C1(n7029), .C2(n4415), .A(n4386), .B(n4370), .ZN(U2926)
         );
  NAND2_X1 U5306 ( .A1(n4418), .A2(DATAI_13_), .ZN(n4384) );
  NAND2_X1 U5307 ( .A1(n4417), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4372) );
  OAI211_X1 U5308 ( .C1(n4373), .C2(n4415), .A(n4384), .B(n4372), .ZN(U2937)
         );
  INV_X1 U5309 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U5310 ( .A1(n4418), .A2(DATAI_11_), .ZN(n4379) );
  NAND2_X1 U5311 ( .A1(n4417), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4374) );
  OAI211_X1 U5312 ( .C1(n6248), .C2(n4420), .A(n4379), .B(n4374), .ZN(U2950)
         );
  INV_X1 U5313 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U5314 ( .A1(n4418), .A2(DATAI_8_), .ZN(n4392) );
  NAND2_X1 U5315 ( .A1(n4417), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4375) );
  OAI211_X1 U5316 ( .C1(n6253), .C2(n4420), .A(n4392), .B(n4375), .ZN(U2947)
         );
  NAND2_X1 U5317 ( .A1(n4418), .A2(DATAI_12_), .ZN(n4388) );
  NAND2_X1 U5318 ( .A1(n4417), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4376) );
  OAI211_X1 U5319 ( .C1(n4415), .C2(n4377), .A(n4388), .B(n4376), .ZN(U2936)
         );
  NAND2_X1 U5320 ( .A1(n4417), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4378) );
  OAI211_X1 U5321 ( .C1(n6925), .C2(n4415), .A(n4379), .B(n4378), .ZN(U2935)
         );
  INV_X1 U5322 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U5323 ( .A1(n4417), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4380) );
  OAI211_X1 U5324 ( .C1(n6258), .C2(n4420), .A(n4381), .B(n4380), .ZN(U2944)
         );
  INV_X1 U5325 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U5326 ( .A1(n4418), .A2(DATAI_9_), .ZN(n4404) );
  NAND2_X1 U5327 ( .A1(n4417), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4382) );
  OAI211_X1 U5328 ( .C1(n6251), .C2(n4420), .A(n4404), .B(n4382), .ZN(U2948)
         );
  INV_X1 U5329 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U5330 ( .A1(n4417), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4383) );
  OAI211_X1 U5331 ( .C1(n6860), .C2(n4420), .A(n4384), .B(n4383), .ZN(U2952)
         );
  INV_X1 U5332 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6973) );
  NAND2_X1 U5333 ( .A1(n4417), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4385) );
  OAI211_X1 U5334 ( .C1(n6973), .C2(n4415), .A(n4386), .B(n4385), .ZN(U2941)
         );
  INV_X1 U5335 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6841) );
  NAND2_X1 U5336 ( .A1(n4417), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4387) );
  OAI211_X1 U5337 ( .C1(n6841), .C2(n4420), .A(n4388), .B(n4387), .ZN(U2951)
         );
  INV_X1 U5338 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6988) );
  NAND2_X1 U5339 ( .A1(n4418), .A2(DATAI_0_), .ZN(n4412) );
  NAND2_X1 U5340 ( .A1(n4417), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4389) );
  OAI211_X1 U5341 ( .C1(n6988), .C2(n4415), .A(n4412), .B(n4389), .ZN(U2939)
         );
  INV_X1 U5342 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U5343 ( .A1(n4418), .A2(DATAI_10_), .ZN(n4400) );
  NAND2_X1 U5344 ( .A1(n4417), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4390) );
  OAI211_X1 U5345 ( .C1(n6859), .C2(n4420), .A(n4400), .B(n4390), .ZN(U2949)
         );
  NAND2_X1 U5346 ( .A1(n4417), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4391) );
  OAI211_X1 U5347 ( .C1(n4415), .C2(n6972), .A(n4392), .B(n4391), .ZN(U2932)
         );
  INV_X1 U5348 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U5349 ( .A1(n4417), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4393) );
  OAI211_X1 U5350 ( .C1(n4415), .C2(n6827), .A(n4394), .B(n4393), .ZN(U2942)
         );
  NAND2_X1 U5351 ( .A1(n4417), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4395) );
  OAI211_X1 U5352 ( .C1(n3928), .C2(n4420), .A(n4396), .B(n4395), .ZN(U2946)
         );
  INV_X1 U5353 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U5354 ( .A1(n4417), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4397) );
  OAI211_X1 U5355 ( .C1(n6256), .C2(n4420), .A(n4398), .B(n4397), .ZN(U2945)
         );
  NAND2_X1 U5356 ( .A1(n4417), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4399) );
  OAI211_X1 U5357 ( .C1(n4401), .C2(n4415), .A(n4400), .B(n4399), .ZN(U2934)
         );
  INV_X1 U5358 ( .A(EAX_REG_14__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U5359 ( .A1(n4418), .A2(DATAI_14_), .ZN(n4414) );
  NAND2_X1 U5360 ( .A1(n4417), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4402) );
  OAI211_X1 U5361 ( .C1(n7058), .C2(n4420), .A(n4414), .B(n4402), .ZN(U2953)
         );
  NAND2_X1 U5362 ( .A1(n4417), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4403) );
  OAI211_X1 U5363 ( .C1(n4405), .C2(n4415), .A(n4404), .B(n4403), .ZN(U2933)
         );
  INV_X1 U5364 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6829) );
  NAND2_X1 U5365 ( .A1(n4418), .A2(DATAI_1_), .ZN(n4408) );
  NAND2_X1 U5366 ( .A1(n4417), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4406) );
  OAI211_X1 U5367 ( .C1(n6829), .C2(n4415), .A(n4408), .B(n4406), .ZN(U2925)
         );
  INV_X1 U5368 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U5369 ( .A1(n4417), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4407) );
  OAI211_X1 U5370 ( .C1(n6265), .C2(n4415), .A(n4408), .B(n4407), .ZN(U2940)
         );
  INV_X1 U5371 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U5372 ( .A1(n4417), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4409) );
  OAI211_X1 U5373 ( .C1(n6260), .C2(n4420), .A(n4410), .B(n4409), .ZN(U2943)
         );
  INV_X1 U5374 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4482) );
  NAND2_X1 U5375 ( .A1(n4417), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4411) );
  OAI211_X1 U5376 ( .C1(n4482), .C2(n4420), .A(n4412), .B(n4411), .ZN(U2924)
         );
  NAND2_X1 U5377 ( .A1(n4417), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4413) );
  OAI211_X1 U5378 ( .C1(n4416), .C2(n4415), .A(n4414), .B(n4413), .ZN(U2938)
         );
  INV_X1 U5379 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6243) );
  AOI22_X1 U5380 ( .A1(n4418), .A2(DATAI_15_), .B1(n4417), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n4419) );
  OAI21_X1 U5381 ( .B1(n6243), .B2(n4420), .A(n4419), .ZN(U2954) );
  NOR2_X1 U5382 ( .A1(n4544), .A2(n6638), .ZN(n4421) );
  NAND2_X1 U5383 ( .A1(n4612), .A2(n4421), .ZN(n4427) );
  INV_X1 U5384 ( .A(n4422), .ZN(n4425) );
  INV_X1 U5385 ( .A(n3400), .ZN(n5460) );
  AND3_X1 U5386 ( .A1(n5460), .A2(n4673), .A3(n6640), .ZN(n4423) );
  NAND3_X1 U5387 ( .A1(n4425), .A2(n4424), .A3(n4423), .ZN(n4646) );
  OR2_X1 U5388 ( .A1(n4646), .A2(n4434), .ZN(n4426) );
  NAND2_X1 U5389 ( .A1(n6221), .A2(n3400), .ZN(n5680) );
  INV_X1 U5390 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6960) );
  NAND2_X1 U5391 ( .A1(n5497), .A2(n5451), .ZN(n4429) );
  NAND2_X1 U5392 ( .A1(n5153), .A2(EBX_REG_0__SCAN_IN), .ZN(n4428) );
  OAI21_X1 U5393 ( .B1(n5662), .B2(EBX_REG_0__SCAN_IN), .A(n4428), .ZN(n4438)
         );
  NAND2_X1 U5394 ( .A1(n4429), .A2(n4438), .ZN(n5959) );
  OAI222_X1 U5395 ( .A1(n5236), .A2(n5680), .B1(n6221), .B2(n6960), .C1(n5959), 
        .C2(n5678), .ZN(U2859) );
  AND2_X1 U5396 ( .A1(n4430), .A2(n4431), .ZN(n4433) );
  OR2_X1 U5397 ( .A1(n4433), .A2(n4432), .ZN(n6293) );
  INV_X1 U5398 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4496) );
  NAND2_X1 U5399 ( .A1(n5484), .A2(n4496), .ZN(n4437) );
  NAND2_X1 U5400 ( .A1(n5153), .A2(n6852), .ZN(n4435) );
  OAI211_X1 U5401 ( .C1(n4434), .C2(EBX_REG_1__SCAN_IN), .A(n4435), .B(n5605), 
        .ZN(n4436) );
  INV_X1 U5402 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4491) );
  NAND2_X1 U5403 ( .A1(n5484), .A2(n4491), .ZN(n4441) );
  INV_X1 U5404 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U5405 ( .A1(n5153), .A2(n6398), .ZN(n4439) );
  OAI211_X1 U5406 ( .C1(n4434), .C2(EBX_REG_2__SCAN_IN), .A(n4439), .B(n5605), 
        .ZN(n4440) );
  AND2_X1 U5407 ( .A1(n4441), .A2(n4440), .ZN(n4488) );
  MUX2_X1 U5408 ( .A(n5495), .B(n5662), .S(EBX_REG_3__SCAN_IN), .Z(n4442) );
  INV_X1 U5409 ( .A(n4442), .ZN(n4444) );
  NAND2_X1 U5410 ( .A1(n5497), .A2(n6386), .ZN(n4443) );
  NAND2_X1 U5411 ( .A1(n4444), .A2(n4443), .ZN(n4517) );
  NAND2_X1 U5412 ( .A1(n5153), .A2(n6377), .ZN(n4445) );
  OAI211_X1 U5413 ( .C1(n4434), .C2(EBX_REG_4__SCAN_IN), .A(n4445), .B(n5605), 
        .ZN(n4446) );
  OAI21_X1 U5414 ( .B1(n5502), .B2(EBX_REG_4__SCAN_IN), .A(n4446), .ZN(n4447)
         );
  NAND2_X1 U5415 ( .A1(n4516), .A2(n4447), .ZN(n4513) );
  OR2_X1 U5416 ( .A1(n4516), .A2(n4447), .ZN(n4448) );
  NAND2_X1 U5417 ( .A1(n4513), .A2(n4448), .ZN(n6372) );
  INV_X1 U5418 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4449) );
  OAI22_X1 U5419 ( .A1(n5678), .A2(n6372), .B1(n4449), .B2(n6221), .ZN(n4450)
         );
  INV_X1 U5420 ( .A(n4450), .ZN(n4451) );
  OAI21_X1 U5421 ( .B1(n6293), .B2(n5680), .A(n4451), .ZN(U2855) );
  XNOR2_X1 U5422 ( .A(n4453), .B(n4452), .ZN(n4632) );
  OR2_X1 U5423 ( .A1(n4456), .A2(n4455), .ZN(n4457) );
  NAND2_X1 U5424 ( .A1(n4454), .A2(n4457), .ZN(n5233) );
  INV_X1 U5425 ( .A(n5233), .ZN(n4499) );
  INV_X1 U5426 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6104) );
  NOR2_X1 U5427 ( .A1(n6388), .A2(n6104), .ZN(n4628) );
  AOI21_X1 U5428 ( .B1(n6299), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4628), 
        .ZN(n4458) );
  OAI21_X1 U5429 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6308), .A(n4458), 
        .ZN(n4459) );
  AOI21_X1 U5430 ( .B1(n4244), .B2(n4499), .A(n4459), .ZN(n4460) );
  OAI21_X1 U5431 ( .B1(n4632), .B2(n6294), .A(n4460), .ZN(U2985) );
  OAI21_X1 U5432 ( .B1(n4461), .B2(n4462), .A(n4430), .ZN(n6204) );
  OR2_X1 U5433 ( .A1(n4464), .A2(n4463), .ZN(n6379) );
  NAND3_X1 U5434 ( .A1(n6379), .A2(n4466), .A3(n6303), .ZN(n4469) );
  NAND2_X1 U5435 ( .A1(n6353), .A2(REIP_REG_3__SCAN_IN), .ZN(n6378) );
  OAI21_X1 U5436 ( .B1(n6063), .B2(n6816), .A(n6378), .ZN(n4467) );
  AOI21_X1 U5437 ( .B1(n6276), .B2(n6208), .A(n4467), .ZN(n4468) );
  OAI211_X1 U5438 ( .C1(n6204), .C2(n6292), .A(n4469), .B(n4468), .ZN(U2983)
         );
  AOI22_X1 U5439 ( .A1(n6747), .A2(UWORD_REG_5__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4470) );
  OAI21_X1 U5440 ( .B1(n4471), .B2(n4484), .A(n4470), .ZN(U2902) );
  AOI22_X1 U5441 ( .A1(n6747), .A2(UWORD_REG_4__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4472) );
  OAI21_X1 U5442 ( .B1(n4473), .B2(n4484), .A(n4472), .ZN(U2903) );
  AOI22_X1 U5443 ( .A1(n6747), .A2(UWORD_REG_6__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4474) );
  OAI21_X1 U5444 ( .B1(n4475), .B2(n4484), .A(n4474), .ZN(U2901) );
  AOI22_X1 U5445 ( .A1(n6747), .A2(UWORD_REG_7__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4476) );
  OAI21_X1 U5446 ( .B1(n4477), .B2(n4484), .A(n4476), .ZN(U2900) );
  AOI22_X1 U5447 ( .A1(n6747), .A2(UWORD_REG_3__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4478) );
  OAI21_X1 U5448 ( .B1(n4479), .B2(n4484), .A(n4478), .ZN(U2904) );
  AOI22_X1 U5449 ( .A1(n6747), .A2(UWORD_REG_2__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4480) );
  OAI21_X1 U5450 ( .B1(n7029), .B2(n4484), .A(n4480), .ZN(U2905) );
  AOI22_X1 U5451 ( .A1(n6747), .A2(UWORD_REG_0__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4481) );
  OAI21_X1 U5452 ( .B1(n4482), .B2(n4484), .A(n4481), .ZN(U2907) );
  AOI22_X1 U5453 ( .A1(n6747), .A2(UWORD_REG_1__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4483) );
  OAI21_X1 U5454 ( .B1(n6829), .B2(n4484), .A(n4483), .ZN(U2906) );
  INV_X1 U5455 ( .A(n4454), .ZN(n4487) );
  INV_X1 U5456 ( .A(n4461), .ZN(n4485) );
  OAI21_X1 U5457 ( .B1(n4487), .B2(n4486), .A(n4485), .ZN(n5139) );
  INV_X1 U5458 ( .A(n5139), .ZN(n6304) );
  NAND2_X1 U5459 ( .A1(n4489), .A2(n4488), .ZN(n4490) );
  AND2_X1 U5460 ( .A1(n4518), .A2(n4490), .ZN(n5132) );
  INV_X1 U5461 ( .A(n5132), .ZN(n6389) );
  OAI22_X1 U5462 ( .A1(n5678), .A2(n6389), .B1(n4491), .B2(n6221), .ZN(n4492)
         );
  AOI21_X1 U5463 ( .B1(n6304), .B2(n6218), .A(n4492), .ZN(n4493) );
  INV_X1 U5464 ( .A(n4493), .ZN(U2857) );
  OR2_X1 U5465 ( .A1(n4494), .A2(n5473), .ZN(n4495) );
  NAND2_X1 U5466 ( .A1(n4849), .A2(n4495), .ZN(n4629) );
  INV_X1 U5467 ( .A(n4629), .ZN(n4497) );
  OAI22_X1 U5468 ( .A1(n5678), .A2(n4497), .B1(n4496), .B2(n6221), .ZN(n4498)
         );
  AOI21_X1 U5469 ( .B1(n4499), .B2(n6218), .A(n4498), .ZN(n4500) );
  INV_X1 U5470 ( .A(n4500), .ZN(U2858) );
  OAI21_X1 U5471 ( .B1(n4432), .B2(n4502), .A(n4501), .ZN(n5174) );
  OAI21_X1 U5472 ( .B1(n4505), .B2(n4504), .A(n4503), .ZN(n4506) );
  INV_X1 U5473 ( .A(n4506), .ZN(n6364) );
  NAND2_X1 U5474 ( .A1(n6364), .A2(n6303), .ZN(n4509) );
  AND2_X1 U5475 ( .A1(n6353), .A2(REIP_REG_5__SCAN_IN), .ZN(n6359) );
  NOR2_X1 U5476 ( .A1(n6308), .A2(n5170), .ZN(n4507) );
  AOI211_X1 U5477 ( .C1(n6299), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n6359), 
        .B(n4507), .ZN(n4508) );
  OAI211_X1 U5478 ( .C1(n6292), .C2(n5174), .A(n4509), .B(n4508), .ZN(U2981)
         );
  MUX2_X1 U5479 ( .A(n5495), .B(n5662), .S(EBX_REG_5__SCAN_IN), .Z(n4510) );
  INV_X1 U5480 ( .A(n4510), .ZN(n4511) );
  NAND2_X1 U5481 ( .A1(n4511), .A2(n3264), .ZN(n4512) );
  NAND2_X1 U5482 ( .A1(n4513), .A2(n4512), .ZN(n4514) );
  NAND2_X1 U5483 ( .A1(n4638), .A2(n4514), .ZN(n6358) );
  INV_X1 U5484 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4515) );
  OAI222_X1 U5485 ( .A1(n6358), .A2(n5678), .B1(n6221), .B2(n4515), .C1(n5680), 
        .C2(n5174), .ZN(U2854) );
  AOI21_X1 U5486 ( .B1(n4518), .B2(n4517), .A(n4516), .ZN(n6382) );
  AOI22_X1 U5487 ( .A1(n6217), .A2(n6382), .B1(n5634), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4519) );
  OAI21_X1 U5488 ( .B1(n6204), .B2(n5680), .A(n4519), .ZN(U2856) );
  INV_X1 U5489 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6090) );
  NAND2_X1 U5490 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6090), .ZN(n4580) );
  INV_X1 U5491 ( .A(n4520), .ZN(n4579) );
  INV_X1 U5492 ( .A(n4523), .ZN(n4529) );
  INV_X1 U5493 ( .A(n4342), .ZN(n4525) );
  AND4_X1 U5494 ( .A1(n6081), .A2(n4527), .A3(n4526), .A4(n4525), .ZN(n4528)
         );
  NAND2_X1 U5495 ( .A1(n4529), .A2(n4528), .ZN(n6596) );
  NAND2_X1 U5496 ( .A1(n4544), .A2(n4556), .ZN(n4561) );
  INV_X1 U5497 ( .A(n4530), .ZN(n5453) );
  MUX2_X1 U5498 ( .A(n4531), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4530), 
        .Z(n4532) );
  NOR2_X1 U5499 ( .A1(n4532), .A2(n4520), .ZN(n4533) );
  NAND2_X1 U5500 ( .A1(n4561), .A2(n4533), .ZN(n4541) );
  XNOR2_X1 U5501 ( .A(n4534), .B(n4521), .ZN(n4539) );
  INV_X1 U5502 ( .A(n4535), .ZN(n4536) );
  OAI21_X1 U5503 ( .B1(n4530), .B2(n4521), .A(n4536), .ZN(n4537) );
  NOR2_X1 U5504 ( .A1(n4537), .A2(n3450), .ZN(n5972) );
  NOR2_X1 U5505 ( .A1(n4563), .A2(n5972), .ZN(n4538) );
  AOI21_X1 U5506 ( .B1(n6598), .B2(n4539), .A(n4538), .ZN(n4540) );
  NAND2_X1 U5507 ( .A1(n4541), .A2(n4540), .ZN(n4542) );
  AOI21_X1 U5508 ( .B1(n3172), .B2(n6596), .A(n4542), .ZN(n5973) );
  NAND2_X1 U5509 ( .A1(n4342), .A2(n5473), .ZN(n4616) );
  AOI21_X1 U5510 ( .B1(n4616), .B2(n6655), .A(READY_N), .ZN(n4543) );
  OAI21_X1 U5511 ( .B1(n6598), .B2(n4342), .A(n4543), .ZN(n4554) );
  INV_X1 U5512 ( .A(n4544), .ZN(n4623) );
  NAND2_X1 U5513 ( .A1(n4612), .A2(n4623), .ZN(n4553) );
  INV_X1 U5514 ( .A(n4545), .ZN(n4546) );
  OR2_X1 U5515 ( .A1(n4547), .A2(n4546), .ZN(n4549) );
  AND2_X1 U5516 ( .A1(n4549), .A2(n4548), .ZN(n4610) );
  INV_X1 U5517 ( .A(n4550), .ZN(n4551) );
  NOR2_X1 U5518 ( .A1(n4610), .A2(n4551), .ZN(n4552) );
  OAI211_X1 U5519 ( .C1(n4612), .C2(n4554), .A(n4553), .B(n4552), .ZN(n4557)
         );
  NAND2_X1 U5520 ( .A1(n4599), .A2(n4555), .ZN(n4604) );
  OAI22_X1 U5521 ( .A1(n4612), .A2(n4556), .B1(n4604), .B2(n6081), .ZN(n4643)
         );
  OR2_X1 U5522 ( .A1(n4557), .A2(n4643), .ZN(n6600) );
  MUX2_X1 U5523 ( .A(n4521), .B(n5973), .S(n6600), .Z(n6608) );
  INV_X1 U5524 ( .A(n6608), .ZN(n4571) );
  INV_X1 U5525 ( .A(n6600), .ZN(n5438) );
  NAND2_X1 U5526 ( .A1(n5438), .A2(n4558), .ZN(n4570) );
  XNOR2_X1 U5527 ( .A(n4530), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4562)
         );
  NAND2_X1 U5528 ( .A1(n4561), .A2(n4562), .ZN(n4567) );
  XNOR2_X1 U5529 ( .A(n4558), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4565)
         );
  NOR2_X1 U5530 ( .A1(n4563), .A2(n4562), .ZN(n4564) );
  AOI21_X1 U5531 ( .B1(n6598), .B2(n4565), .A(n4564), .ZN(n4566) );
  NAND2_X1 U5532 ( .A1(n4567), .A2(n4566), .ZN(n4568) );
  AOI21_X1 U5533 ( .B1(n4560), .B2(n6596), .A(n4568), .ZN(n5449) );
  NAND2_X1 U5534 ( .A1(n6600), .A2(n5449), .ZN(n4569) );
  NAND3_X1 U5535 ( .A1(n4571), .A2(n6606), .A3(n5452), .ZN(n4578) );
  INV_X1 U5536 ( .A(n4975), .ZN(n5095) );
  NOR2_X1 U5537 ( .A1(n4572), .A2(n5095), .ZN(n4573) );
  XNOR2_X1 U5538 ( .A(n4573), .B(n4575), .ZN(n6183) );
  INV_X1 U5539 ( .A(n6183), .ZN(n4574) );
  OAI22_X1 U5540 ( .A1(n6600), .A2(n4575), .B1(n4574), .B2(n6081), .ZN(n4577)
         );
  NOR2_X1 U5541 ( .A1(n4575), .A2(n4580), .ZN(n4576) );
  AOI21_X1 U5542 ( .B1(n4577), .B2(n5452), .A(n4576), .ZN(n4582) );
  OAI211_X1 U5543 ( .C1(n4580), .C2(n4579), .A(n4578), .B(n4582), .ZN(n6620)
         );
  NAND2_X1 U5544 ( .A1(n4582), .A2(n4581), .ZN(n4583) );
  NAND2_X1 U5545 ( .A1(n6620), .A2(n4583), .ZN(n6632) );
  AND2_X1 U5546 ( .A1(n6632), .A2(n6090), .ZN(n4584) );
  NAND2_X1 U5547 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4591), .ZN(n6645) );
  NOR2_X1 U5548 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n4833) );
  OAI21_X1 U5549 ( .B1(n4584), .B2(n6645), .A(n4877), .ZN(n6404) );
  OR3_X1 U5550 ( .A1(n4585), .A2(n4587), .A3(n3868), .ZN(n4893) );
  INV_X1 U5551 ( .A(n4893), .ZN(n4750) );
  NAND2_X1 U5552 ( .A1(n4750), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4889) );
  INV_X1 U5553 ( .A(n4889), .ZN(n4586) );
  INV_X1 U5554 ( .A(n4585), .ZN(n4663) );
  NOR2_X1 U5555 ( .A1(n4586), .A2(n6528), .ZN(n6437) );
  AND2_X1 U5556 ( .A1(n3868), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6529) );
  NAND2_X1 U5557 ( .A1(n4773), .A2(n6529), .ZN(n6489) );
  AOI21_X1 U5558 ( .B1(n6437), .B2(n6489), .A(n6535), .ZN(n4589) );
  NOR2_X1 U5559 ( .A1(n6535), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4712) );
  INV_X1 U5560 ( .A(n4712), .ZN(n6409) );
  INV_X1 U5561 ( .A(n3172), .ZN(n6407) );
  NAND2_X1 U5562 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5263), .ZN(n4594) );
  INV_X1 U5563 ( .A(n4594), .ZN(n5968) );
  OAI22_X1 U5564 ( .A1(n3887), .A2(n6409), .B1(n6407), .B2(n5968), .ZN(n4588)
         );
  OAI21_X1 U5565 ( .B1(n4589), .B2(n4588), .A(n6404), .ZN(n4590) );
  OAI21_X1 U5566 ( .B1(n6435), .B2(n6404), .A(n4590), .ZN(U3462) );
  INV_X1 U5567 ( .A(n6404), .ZN(n4598) );
  AOI222_X1 U5568 ( .A1(n6632), .A2(n4591), .B1(n4968), .B2(n6486), .C1(n6597), 
        .C2(n4594), .ZN(n4593) );
  NAND2_X1 U5569 ( .A1(n4598), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4592) );
  OAI21_X1 U5570 ( .B1(n4598), .B2(n4593), .A(n4592), .ZN(U3465) );
  XNOR2_X1 U5571 ( .A(n4585), .B(n6529), .ZN(n4595) );
  AOI22_X1 U5572 ( .A1(n4595), .A2(n6486), .B1(n4594), .B2(n4560), .ZN(n4597)
         );
  NAND2_X1 U5573 ( .A1(n4598), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4596) );
  OAI21_X1 U5574 ( .B1(n4598), .B2(n4597), .A(n4596), .ZN(U3463) );
  NAND2_X1 U5575 ( .A1(n4873), .A2(n6655), .ZN(n4846) );
  NAND3_X1 U5576 ( .A1(n4342), .A2(n4846), .A3(n4599), .ZN(n4600) );
  NAND3_X1 U5577 ( .A1(n4600), .A2(n4845), .A3(n4647), .ZN(n4601) );
  NAND2_X1 U5578 ( .A1(n4602), .A2(n4601), .ZN(n4609) );
  NAND2_X1 U5579 ( .A1(n4603), .A2(n6655), .ZN(n4606) );
  INV_X1 U5580 ( .A(n4604), .ZN(n4605) );
  NAND2_X1 U5581 ( .A1(n4606), .A2(n4605), .ZN(n4608) );
  MUX2_X1 U5582 ( .A(n4609), .B(n4608), .S(n4607), .Z(n4614) );
  AOI21_X1 U5583 ( .B1(n4612), .B2(n4611), .A(n4610), .ZN(n4613) );
  OAI211_X1 U5584 ( .C1(n4673), .C2(n4615), .A(n6081), .B(n4616), .ZN(n4617)
         );
  OR2_X1 U5585 ( .A1(n4618), .A2(n4617), .ZN(n4619) );
  INV_X1 U5586 ( .A(n4620), .ZN(n4621) );
  AND2_X1 U5587 ( .A1(n4627), .A2(n4621), .ZN(n5389) );
  INV_X1 U5588 ( .A(n5389), .ZN(n4622) );
  NAND2_X1 U5589 ( .A1(n4627), .A2(n6598), .ZN(n5962) );
  NAND2_X1 U5590 ( .A1(n4627), .A2(n4623), .ZN(n5814) );
  NAND2_X1 U5591 ( .A1(n6348), .A2(n5814), .ZN(n6350) );
  INV_X1 U5592 ( .A(n6350), .ZN(n6321) );
  AND2_X1 U5593 ( .A1(n5962), .A2(n5451), .ZN(n4957) );
  OR2_X1 U5594 ( .A1(n6321), .A2(n4957), .ZN(n4624) );
  NOR2_X1 U5595 ( .A1(n6353), .A2(n4627), .ZN(n5963) );
  NOR2_X1 U5596 ( .A1(n6392), .A2(n5389), .ZN(n5357) );
  NOR2_X1 U5597 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5357), .ZN(n5957)
         );
  NOR2_X1 U5598 ( .A1(n5963), .A2(n5957), .ZN(n6347) );
  MUX2_X1 U5599 ( .A(n4624), .B(n6347), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4631) );
  OAI21_X1 U5600 ( .B1(n4615), .B2(n3310), .A(n4625), .ZN(n4626) );
  NAND2_X1 U5601 ( .A1(n4627), .A2(n4626), .ZN(n6390) );
  AOI21_X1 U5602 ( .B1(n6383), .B2(n4629), .A(n4628), .ZN(n4630) );
  OAI211_X1 U5603 ( .C1(n4632), .C2(n6370), .A(n4631), .B(n4630), .ZN(U3017)
         );
  OAI21_X1 U5604 ( .B1(n3923), .B2(n3922), .A(n4655), .ZN(n6178) );
  INV_X1 U5605 ( .A(n6178), .ZN(n6284) );
  INV_X1 U5606 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U5607 ( .A1(n5484), .A2(n6173), .ZN(n4636) );
  NAND2_X1 U5608 ( .A1(n5153), .A2(n6355), .ZN(n4634) );
  OAI211_X1 U5609 ( .C1(n4434), .C2(EBX_REG_6__SCAN_IN), .A(n4634), .B(n5605), 
        .ZN(n4635) );
  AND2_X1 U5610 ( .A1(n4638), .A2(n4637), .ZN(n4639) );
  NOR2_X1 U5611 ( .A1(n4704), .A2(n4639), .ZN(n6352) );
  INV_X1 U5612 ( .A(n6352), .ZN(n4640) );
  OAI22_X1 U5613 ( .A1(n5678), .A2(n4640), .B1(n6173), .B2(n6221), .ZN(n4641)
         );
  AOI21_X1 U5614 ( .B1(n6284), .B2(n6218), .A(n4641), .ZN(n4642) );
  INV_X1 U5615 ( .A(n4642), .ZN(U2853) );
  NAND2_X1 U5616 ( .A1(n4643), .A2(n6640), .ZN(n4644) );
  OAI211_X2 U5617 ( .C1(n4839), .C2(n4646), .A(n4645), .B(n4644), .ZN(n6240)
         );
  AND2_X1 U5618 ( .A1(n4864), .A2(n3400), .ZN(n4650) );
  INV_X1 U5619 ( .A(n4650), .ZN(n4648) );
  AND2_X1 U5620 ( .A1(n4648), .A2(n4647), .ZN(n4649) );
  AND2_X1 U5621 ( .A1(n6240), .A2(n3481), .ZN(n6228) );
  INV_X1 U5622 ( .A(DATAI_5_), .ZN(n4863) );
  OAI222_X1 U5623 ( .A1(n5174), .A2(n5697), .B1(n5235), .B2(n4863), .C1(n6240), 
        .C2(n6258), .ZN(U2886) );
  INV_X1 U5624 ( .A(DATAI_2_), .ZN(n7055) );
  OAI222_X1 U5625 ( .A1(n5139), .A2(n5697), .B1(n5235), .B2(n7055), .C1(n6240), 
        .C2(n6973), .ZN(U2889) );
  INV_X1 U5626 ( .A(DATAI_4_), .ZN(n4674) );
  OAI222_X1 U5627 ( .A1(n6293), .A2(n5697), .B1(n5235), .B2(n4674), .C1(n6240), 
        .C2(n6260), .ZN(U2887) );
  INV_X1 U5628 ( .A(DATAI_3_), .ZN(n4689) );
  OAI222_X1 U5629 ( .A1(n6204), .A2(n5697), .B1(n5235), .B2(n4689), .C1(n6827), 
        .C2(n6240), .ZN(U2888) );
  OAI21_X1 U5630 ( .B1(n4653), .B2(n4652), .A(n4651), .ZN(n6337) );
  XOR2_X1 U5631 ( .A(n4655), .B(n4654), .Z(n5255) );
  NAND2_X1 U5632 ( .A1(n6353), .A2(REIP_REG_7__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U5633 ( .A1(n6299), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4656)
         );
  OAI211_X1 U5634 ( .C1(n6308), .C2(n5252), .A(n6334), .B(n4656), .ZN(n4657)
         );
  AOI21_X1 U5635 ( .B1(n5255), .B2(n4244), .A(n4657), .ZN(n4658) );
  OAI21_X1 U5636 ( .B1(n6337), .B2(n6294), .A(n4658), .ZN(U2979) );
  NAND3_X1 U5637 ( .A1(n6435), .A2(n6607), .A3(n6601), .ZN(n4816) );
  NOR2_X1 U5638 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4816), .ZN(n5076)
         );
  INV_X1 U5639 ( .A(n5076), .ZN(n4661) );
  INV_X1 U5640 ( .A(n4675), .ZN(n4659) );
  NOR2_X1 U5641 ( .A1(n4659), .A2(n6737), .ZN(n5261) );
  INV_X1 U5642 ( .A(n4708), .ZN(n4660) );
  NOR2_X1 U5643 ( .A1(n4660), .A2(n5258), .ZN(n4676) );
  OAI21_X1 U5644 ( .B1(n4676), .B2(n6737), .A(n4749), .ZN(n4979) );
  AOI211_X1 U5645 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4661), .A(n5261), .B(
        n4979), .ZN(n4668) );
  INV_X1 U5646 ( .A(n3868), .ZN(n4772) );
  AND2_X1 U5647 ( .A1(n4585), .A2(n4772), .ZN(n4662) );
  NAND2_X1 U5648 ( .A1(n4662), .A2(n3887), .ZN(n4820) );
  INV_X1 U5649 ( .A(n4820), .ZN(n4813) );
  NAND2_X1 U5650 ( .A1(n4813), .A2(n4819), .ZN(n4886) );
  NAND3_X1 U5651 ( .A1(n4663), .A2(n3598), .A3(n3868), .ZN(n4913) );
  NOR2_X1 U5652 ( .A1(n4913), .A2(n4819), .ZN(n4671) );
  NOR3_X1 U5653 ( .A1(n5080), .A2(n4671), .A3(n6535), .ZN(n4666) );
  NAND2_X1 U5654 ( .A1(n6407), .A2(n3261), .ZN(n4811) );
  OAI21_X1 U5655 ( .B1(n4666), .B2(n4712), .A(n4811), .ZN(n4667) );
  INV_X1 U5656 ( .A(DATAI_20_), .ZN(n4669) );
  OR2_X1 U5657 ( .A1(n6292), .A2(n4669), .ZN(n6568) );
  INV_X1 U5658 ( .A(n6568), .ZN(n6460) );
  INV_X1 U5659 ( .A(DATAI_28_), .ZN(n4670) );
  OR2_X1 U5660 ( .A1(n6292), .A2(n4670), .ZN(n6463) );
  NOR2_X1 U5661 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n5263), .ZN(n6718) );
  NOR2_X2 U5662 ( .A1(n4881), .A2(n4673), .ZN(n6563) );
  NOR2_X2 U5663 ( .A1(n4674), .A2(n4877), .ZN(n6565) );
  NOR2_X1 U5664 ( .A1(n4675), .A2(n6737), .ZN(n5259) );
  INV_X1 U5665 ( .A(n5259), .ZN(n5186) );
  INV_X1 U5666 ( .A(n4676), .ZN(n4972) );
  OAI22_X1 U5667 ( .A1(n4811), .A2(n6535), .B1(n5186), .B2(n4972), .ZN(n5075)
         );
  AOI22_X1 U5668 ( .A1(n6563), .A2(n5076), .B1(n6565), .B2(n5075), .ZN(n4677)
         );
  OAI21_X1 U5669 ( .B1(n6463), .B2(n5078), .A(n4677), .ZN(n4678) );
  AOI21_X1 U5670 ( .B1(n6460), .B2(n5080), .A(n4678), .ZN(n4679) );
  OAI21_X1 U5671 ( .B1(n5083), .B2(n6978), .A(n4679), .ZN(U3024) );
  INV_X1 U5672 ( .A(DATAI_23_), .ZN(n4680) );
  OR2_X1 U5673 ( .A1(n6292), .A2(n4680), .ZN(n6593) );
  INV_X1 U5674 ( .A(n6593), .ZN(n6516) );
  INV_X1 U5675 ( .A(DATAI_31_), .ZN(n4681) );
  OR2_X1 U5676 ( .A1(n6292), .A2(n4681), .ZN(n6524) );
  NOR2_X2 U5677 ( .A1(n4881), .A2(n5460), .ZN(n6584) );
  INV_X1 U5678 ( .A(DATAI_7_), .ZN(n4700) );
  NOR2_X2 U5679 ( .A1(n4700), .A2(n4877), .ZN(n6588) );
  AOI22_X1 U5680 ( .A1(n6584), .A2(n5076), .B1(n6588), .B2(n5075), .ZN(n4682)
         );
  OAI21_X1 U5681 ( .B1(n6524), .B2(n5078), .A(n4682), .ZN(n4683) );
  AOI21_X1 U5682 ( .B1(n6516), .B2(n5080), .A(n4683), .ZN(n4684) );
  OAI21_X1 U5683 ( .B1(n5083), .B2(n4685), .A(n4684), .ZN(U3027) );
  INV_X1 U5684 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4693) );
  INV_X1 U5685 ( .A(DATAI_19_), .ZN(n4686) );
  OR2_X1 U5686 ( .A1(n6292), .A2(n4686), .ZN(n6562) );
  INV_X1 U5687 ( .A(n6562), .ZN(n6500) );
  INV_X1 U5688 ( .A(DATAI_27_), .ZN(n4687) );
  OR2_X1 U5689 ( .A1(n6292), .A2(n4687), .ZN(n6503) );
  NOR2_X2 U5690 ( .A1(n4881), .A2(n4688), .ZN(n6557) );
  NOR2_X2 U5691 ( .A1(n4689), .A2(n4877), .ZN(n6559) );
  AOI22_X1 U5692 ( .A1(n6557), .A2(n5076), .B1(n6559), .B2(n5075), .ZN(n4690)
         );
  OAI21_X1 U5693 ( .B1(n6503), .B2(n5078), .A(n4690), .ZN(n4691) );
  AOI21_X1 U5694 ( .B1(n6500), .B2(n5080), .A(n4691), .ZN(n4692) );
  OAI21_X1 U5695 ( .B1(n5083), .B2(n4693), .A(n4692), .ZN(U3023) );
  INV_X1 U5696 ( .A(DATAI_16_), .ZN(n4694) );
  OR2_X1 U5697 ( .A1(n6292), .A2(n4694), .ZN(n6544) );
  INV_X1 U5698 ( .A(n6544), .ZN(n6482) );
  INV_X1 U5699 ( .A(DATAI_24_), .ZN(n4695) );
  OR2_X1 U5700 ( .A1(n6292), .A2(n4695), .ZN(n6495) );
  NOR2_X2 U5701 ( .A1(n4881), .A2(n4857), .ZN(n6526) );
  INV_X1 U5702 ( .A(DATAI_0_), .ZN(n5234) );
  NOR2_X2 U5703 ( .A1(n5234), .A2(n4877), .ZN(n6541) );
  AOI22_X1 U5704 ( .A1(n6526), .A2(n5076), .B1(n6541), .B2(n5075), .ZN(n4696)
         );
  OAI21_X1 U5705 ( .B1(n6495), .B2(n5078), .A(n4696), .ZN(n4697) );
  AOI21_X1 U5706 ( .B1(n6482), .B2(n5080), .A(n4697), .ZN(n4698) );
  OAI21_X1 U5707 ( .B1(n5083), .B2(n4699), .A(n4698), .ZN(U3020) );
  INV_X1 U5708 ( .A(n5255), .ZN(n4707) );
  OAI222_X1 U5709 ( .A1(n5697), .A2(n4707), .B1(n6240), .B2(n3928), .C1(n4700), 
        .C2(n5235), .ZN(U2884) );
  MUX2_X1 U5710 ( .A(n5495), .B(n5662), .S(EBX_REG_7__SCAN_IN), .Z(n4702) );
  NOR2_X1 U5711 ( .A1(n5503), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4701)
         );
  NOR2_X1 U5712 ( .A1(n4702), .A2(n4701), .ZN(n4703) );
  NOR2_X1 U5713 ( .A1(n4704), .A2(n4703), .ZN(n4705) );
  OR2_X1 U5714 ( .A1(n4745), .A2(n4705), .ZN(n5246) );
  INV_X1 U5715 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4706) );
  OAI222_X1 U5716 ( .A1(n5246), .A2(n5678), .B1(n5680), .B2(n4707), .C1(n4706), 
        .C2(n6221), .ZN(U2852) );
  NAND3_X1 U5717 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6607), .A3(n6601), .ZN(n4803) );
  NOR2_X1 U5718 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4803), .ZN(n5011)
         );
  INV_X1 U5719 ( .A(n5011), .ZN(n4709) );
  NOR2_X1 U5720 ( .A1(n5258), .A2(n4708), .ZN(n5179) );
  OAI21_X1 U5721 ( .B1(n5179), .B2(n6737), .A(n4749), .ZN(n5185) );
  AOI211_X1 U5722 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4709), .A(n5261), .B(
        n5185), .ZN(n4715) );
  AND2_X1 U5723 ( .A1(n6528), .A2(n4772), .ZN(n4806) );
  INV_X1 U5724 ( .A(n4806), .ZN(n4710) );
  INV_X1 U5725 ( .A(n5014), .ZN(n4711) );
  NAND2_X1 U5726 ( .A1(n4773), .A2(n5175), .ZN(n6514) );
  NOR3_X1 U5727 ( .A1(n4711), .A2(n6517), .A3(n6535), .ZN(n4713) );
  NAND2_X1 U5728 ( .A1(n3261), .A2(n3172), .ZN(n4716) );
  OAI21_X1 U5729 ( .B1(n4713), .B2(n4712), .A(n4716), .ZN(n4714) );
  NAND2_X1 U5730 ( .A1(n4715), .A2(n4714), .ZN(n5016) );
  OR2_X1 U5731 ( .A1(n4716), .A2(n6535), .ZN(n4718) );
  NAND2_X1 U5732 ( .A1(n5259), .A2(n5179), .ZN(n4717) );
  NAND2_X1 U5733 ( .A1(n4718), .A2(n4717), .ZN(n5010) );
  AOI22_X1 U5734 ( .A1(n6563), .A2(n5011), .B1(n6565), .B2(n5010), .ZN(n4720)
         );
  OR2_X1 U5735 ( .A1(n6514), .A2(n6463), .ZN(n4719) );
  OAI211_X1 U5736 ( .C1(n6568), .C2(n5014), .A(n4720), .B(n4719), .ZN(n4721)
         );
  AOI21_X1 U5737 ( .B1(n5016), .B2(INSTQUEUE_REG_8__4__SCAN_IN), .A(n4721), 
        .ZN(n4722) );
  INV_X1 U5738 ( .A(n4722), .ZN(U3088) );
  AOI22_X1 U5739 ( .A1(n6584), .A2(n5011), .B1(n6588), .B2(n5010), .ZN(n4724)
         );
  OR2_X1 U5740 ( .A1(n6514), .A2(n6524), .ZN(n4723) );
  OAI211_X1 U5741 ( .C1(n6593), .C2(n5014), .A(n4724), .B(n4723), .ZN(n4725)
         );
  AOI21_X1 U5742 ( .B1(n5016), .B2(INSTQUEUE_REG_8__7__SCAN_IN), .A(n4725), 
        .ZN(n4726) );
  INV_X1 U5743 ( .A(n4726), .ZN(U3091) );
  AOI22_X1 U5744 ( .A1(n6526), .A2(n5011), .B1(n6541), .B2(n5010), .ZN(n4728)
         );
  OR2_X1 U5745 ( .A1(n5014), .A2(n6544), .ZN(n4727) );
  OAI211_X1 U5746 ( .C1(n6514), .C2(n6495), .A(n4728), .B(n4727), .ZN(n4729)
         );
  AOI21_X1 U5747 ( .B1(n5016), .B2(INSTQUEUE_REG_8__0__SCAN_IN), .A(n4729), 
        .ZN(n4730) );
  INV_X1 U5748 ( .A(n4730), .ZN(U3084) );
  AOI22_X1 U5749 ( .A1(n6557), .A2(n5011), .B1(n6559), .B2(n5010), .ZN(n4732)
         );
  OR2_X1 U5750 ( .A1(n6514), .A2(n6503), .ZN(n4731) );
  OAI211_X1 U5751 ( .C1(n6562), .C2(n5014), .A(n4732), .B(n4731), .ZN(n4733)
         );
  AOI21_X1 U5752 ( .B1(n5016), .B2(INSTQUEUE_REG_8__3__SCAN_IN), .A(n4733), 
        .ZN(n4734) );
  INV_X1 U5753 ( .A(n4734), .ZN(U3087) );
  NAND2_X1 U5754 ( .A1(n4736), .A2(n4737), .ZN(n4738) );
  NAND2_X1 U5755 ( .A1(n4994), .A2(n4738), .ZN(n6165) );
  AOI22_X1 U5756 ( .A1(n6236), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6230), .ZN(n4739) );
  OAI21_X1 U5757 ( .B1(n6165), .B2(n5697), .A(n4739), .ZN(U2882) );
  OAI21_X1 U5758 ( .B1(n4740), .B2(n4741), .A(n4736), .ZN(n5316) );
  INV_X1 U5759 ( .A(n5316), .ZN(n4798) );
  NAND2_X1 U5760 ( .A1(n5153), .A2(n4961), .ZN(n4742) );
  OAI211_X1 U5761 ( .C1(n4434), .C2(EBX_REG_8__SCAN_IN), .A(n4742), .B(n5605), 
        .ZN(n4743) );
  OAI21_X1 U5762 ( .B1(n5502), .B2(EBX_REG_8__SCAN_IN), .A(n4743), .ZN(n4744)
         );
  OR2_X1 U5763 ( .A1(n4745), .A2(n4744), .ZN(n4746) );
  NAND2_X1 U5764 ( .A1(n6159), .A2(n4746), .ZN(n5311) );
  INV_X1 U5765 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6946) );
  OAI22_X1 U5766 ( .A1(n5678), .A2(n5311), .B1(n6946), .B2(n6221), .ZN(n4747)
         );
  AOI21_X1 U5767 ( .B1(n4798), .B2(n6218), .A(n4747), .ZN(n4748) );
  INV_X1 U5768 ( .A(n4748), .ZN(U2851) );
  INV_X1 U5769 ( .A(n4917), .ZN(n4920) );
  NOR2_X1 U5770 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4920), .ZN(n5085)
         );
  OAI21_X1 U5771 ( .B1(n5258), .B2(n6737), .A(n4749), .ZN(n5260) );
  NOR3_X1 U5772 ( .A1(n5260), .A2(n6435), .A3(n5259), .ZN(n4754) );
  NAND2_X1 U5773 ( .A1(n4560), .A2(n4665), .ZN(n4775) );
  NOR2_X2 U5774 ( .A1(n4913), .A2(n4968), .ZN(n5089) );
  INV_X1 U5775 ( .A(n5087), .ZN(n4751) );
  OAI21_X1 U5776 ( .B1(n5089), .B2(n4751), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4752) );
  NAND3_X1 U5777 ( .A1(n4775), .A2(n6486), .A3(n4752), .ZN(n4753) );
  OAI211_X1 U5778 ( .C1(n5085), .C2(n5263), .A(n4754), .B(n4753), .ZN(n4755)
         );
  INV_X1 U5779 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4759) );
  INV_X1 U5780 ( .A(n4775), .ZN(n6485) );
  NAND2_X1 U5781 ( .A1(n6485), .A2(n6530), .ZN(n4780) );
  NAND2_X1 U5782 ( .A1(n5261), .A2(n5258), .ZN(n4779) );
  OAI22_X1 U5783 ( .A1(n4780), .A2(n6407), .B1(n6435), .B2(n4779), .ZN(n5084)
         );
  AOI22_X1 U5784 ( .A1(n6584), .A2(n5085), .B1(n6588), .B2(n5084), .ZN(n4756)
         );
  OAI21_X1 U5785 ( .B1(n6524), .B2(n5087), .A(n4756), .ZN(n4757) );
  AOI21_X1 U5786 ( .B1(n6516), .B2(n5089), .A(n4757), .ZN(n4758) );
  OAI21_X1 U5787 ( .B1(n5092), .B2(n4759), .A(n4758), .ZN(U3139) );
  INV_X1 U5788 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4763) );
  AOI22_X1 U5789 ( .A1(n6563), .A2(n5085), .B1(n6565), .B2(n5084), .ZN(n4760)
         );
  OAI21_X1 U5790 ( .B1(n6463), .B2(n5087), .A(n4760), .ZN(n4761) );
  AOI21_X1 U5791 ( .B1(n6460), .B2(n5089), .A(n4761), .ZN(n4762) );
  OAI21_X1 U5792 ( .B1(n5092), .B2(n4763), .A(n4762), .ZN(U3136) );
  INV_X1 U5793 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4767) );
  AOI22_X1 U5794 ( .A1(n6526), .A2(n5085), .B1(n6541), .B2(n5084), .ZN(n4764)
         );
  OAI21_X1 U5795 ( .B1(n6495), .B2(n5087), .A(n4764), .ZN(n4765) );
  AOI21_X1 U5796 ( .B1(n6482), .B2(n5089), .A(n4765), .ZN(n4766) );
  OAI21_X1 U5797 ( .B1(n5092), .B2(n4767), .A(n4766), .ZN(U3132) );
  INV_X1 U5798 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4771) );
  AOI22_X1 U5799 ( .A1(n6557), .A2(n5085), .B1(n6559), .B2(n5084), .ZN(n4768)
         );
  OAI21_X1 U5800 ( .B1(n6503), .B2(n5087), .A(n4768), .ZN(n4769) );
  AOI21_X1 U5801 ( .B1(n6500), .B2(n5089), .A(n4769), .ZN(n4770) );
  OAI21_X1 U5802 ( .B1(n5092), .B2(n4771), .A(n4770), .ZN(U3135) );
  NAND2_X1 U5803 ( .A1(n4773), .A2(n4772), .ZN(n4969) );
  AND2_X1 U5804 ( .A1(n3868), .A2(n4819), .ZN(n6405) );
  NAND2_X1 U5805 ( .A1(n4773), .A2(n6405), .ZN(n6523) );
  INV_X1 U5806 ( .A(n6523), .ZN(n6511) );
  OAI21_X1 U5807 ( .B1(n6477), .B2(n6511), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4774) );
  NAND3_X1 U5808 ( .A1(n4775), .A2(n6486), .A3(n4774), .ZN(n4777) );
  NAND2_X1 U5809 ( .A1(n5177), .A2(n3578), .ZN(n4778) );
  AOI211_X1 U5810 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4778), .A(n5259), .B(
        n5260), .ZN(n4776) );
  NAND3_X1 U5811 ( .A1(n6435), .A2(n4777), .A3(n4776), .ZN(n6478) );
  INV_X1 U5812 ( .A(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4784) );
  INV_X1 U5813 ( .A(n6503), .ZN(n6558) );
  INV_X1 U5814 ( .A(n4778), .ZN(n6476) );
  OAI22_X1 U5815 ( .A1(n4780), .A2(n3172), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4779), .ZN(n6475) );
  AOI22_X1 U5816 ( .A1(n6557), .A2(n6476), .B1(n6559), .B2(n6475), .ZN(n4781)
         );
  OAI21_X1 U5817 ( .B1(n6562), .B2(n6523), .A(n4781), .ZN(n4782) );
  AOI21_X1 U5818 ( .B1(n6558), .B2(n6477), .A(n4782), .ZN(n4783) );
  OAI21_X1 U5819 ( .B1(n5067), .B2(n4784), .A(n4783), .ZN(U3071) );
  INV_X1 U5820 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4788) );
  INV_X1 U5821 ( .A(n6524), .ZN(n6585) );
  AOI22_X1 U5822 ( .A1(n6584), .A2(n6476), .B1(n6588), .B2(n6475), .ZN(n4785)
         );
  OAI21_X1 U5823 ( .B1(n6593), .B2(n6523), .A(n4785), .ZN(n4786) );
  AOI21_X1 U5824 ( .B1(n6585), .B2(n6477), .A(n4786), .ZN(n4787) );
  OAI21_X1 U5825 ( .B1(n5067), .B2(n4788), .A(n4787), .ZN(U3075) );
  INV_X1 U5826 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4792) );
  INV_X1 U5827 ( .A(n6463), .ZN(n6564) );
  AOI22_X1 U5828 ( .A1(n6563), .A2(n6476), .B1(n6565), .B2(n6475), .ZN(n4789)
         );
  OAI21_X1 U5829 ( .B1(n6568), .B2(n6523), .A(n4789), .ZN(n4790) );
  AOI21_X1 U5830 ( .B1(n6564), .B2(n6477), .A(n4790), .ZN(n4791) );
  OAI21_X1 U5831 ( .B1(n5067), .B2(n4792), .A(n4791), .ZN(U3072) );
  OAI21_X1 U5832 ( .B1(n4795), .B2(n4794), .A(n4793), .ZN(n4967) );
  INV_X1 U5833 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5303) );
  NOR2_X1 U5834 ( .A1(n6388), .A2(n5303), .ZN(n4964) );
  AOI21_X1 U5835 ( .B1(n6299), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n4964), 
        .ZN(n4796) );
  OAI21_X1 U5836 ( .B1(n5309), .B2(n6308), .A(n4796), .ZN(n4797) );
  AOI21_X1 U5837 ( .B1(n4798), .B2(n4244), .A(n4797), .ZN(n4799) );
  OAI21_X1 U5838 ( .B1(n4967), .B2(n6294), .A(n4799), .ZN(U2978) );
  AND2_X1 U5839 ( .A1(n3172), .A2(n6597), .ZN(n4916) );
  NOR2_X1 U5840 ( .A1(n5177), .A2(n4803), .ZN(n4954) );
  AOI21_X1 U5841 ( .B1(n4916), .B2(n3261), .A(n4954), .ZN(n4805) );
  OR2_X1 U5842 ( .A1(n3868), .A2(n6738), .ZN(n5093) );
  INV_X1 U5843 ( .A(n5093), .ZN(n4800) );
  AOI21_X1 U5844 ( .B1(n6528), .B2(n4800), .A(n6535), .ZN(n4802) );
  AOI22_X1 U5845 ( .A1(n4805), .A2(n4802), .B1(n6535), .B2(n4803), .ZN(n4801)
         );
  NAND2_X1 U5846 ( .A1(n6488), .A2(n4801), .ZN(n4953) );
  INV_X1 U5847 ( .A(n4802), .ZN(n4804) );
  OAI22_X1 U5848 ( .A1(n4805), .A2(n4804), .B1(n6737), .B2(n4803), .ZN(n4952)
         );
  AOI22_X1 U5849 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4953), .B1(n6565), 
        .B2(n4952), .ZN(n4808) );
  AOI22_X1 U5850 ( .A1(n5297), .A2(n6460), .B1(n4954), .B2(n6563), .ZN(n4807)
         );
  OAI211_X1 U5851 ( .C1(n5014), .C2(n6463), .A(n4808), .B(n4807), .ZN(U3096)
         );
  AOI22_X1 U5852 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4953), .B1(n6559), 
        .B2(n4952), .ZN(n4810) );
  AOI22_X1 U5853 ( .A1(n5297), .A2(n6500), .B1(n4954), .B2(n6557), .ZN(n4809)
         );
  OAI211_X1 U5854 ( .C1(n5014), .C2(n6503), .A(n4810), .B(n4809), .ZN(U3095)
         );
  INV_X1 U5855 ( .A(n4811), .ZN(n4812) );
  NOR2_X1 U5856 ( .A1(n5177), .A2(n4816), .ZN(n4883) );
  AOI21_X1 U5857 ( .B1(n4812), .B2(n6597), .A(n4883), .ZN(n4818) );
  AOI21_X1 U5858 ( .B1(n4813), .B2(STATEBS16_REG_SCAN_IN), .A(n6535), .ZN(
        n4815) );
  AOI22_X1 U5859 ( .A1(n4818), .A2(n4815), .B1(n6535), .B2(n4816), .ZN(n4814)
         );
  NAND2_X1 U5860 ( .A1(n6488), .A2(n4814), .ZN(n4879) );
  INV_X1 U5861 ( .A(n4815), .ZN(n4817) );
  OAI22_X1 U5862 ( .A1(n4818), .A2(n4817), .B1(n6737), .B2(n4816), .ZN(n4878)
         );
  AOI22_X1 U5863 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4879), .B1(n6541), 
        .B2(n4878), .ZN(n4822) );
  NOR2_X2 U5864 ( .A1(n4820), .A2(n4819), .ZN(n6431) );
  AOI22_X1 U5865 ( .A1(n6526), .A2(n4883), .B1(n6431), .B2(n6482), .ZN(n4821)
         );
  OAI211_X1 U5866 ( .C1(n6495), .C2(n4886), .A(n4822), .B(n4821), .ZN(U3028)
         );
  AOI22_X1 U5867 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4953), .B1(n6588), 
        .B2(n4952), .ZN(n4824) );
  AOI22_X1 U5868 ( .A1(n5297), .A2(n6516), .B1(n4954), .B2(n6584), .ZN(n4823)
         );
  OAI211_X1 U5869 ( .C1(n5014), .C2(n6524), .A(n4824), .B(n4823), .ZN(U3099)
         );
  AOI22_X1 U5870 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4879), .B1(n6588), 
        .B2(n4878), .ZN(n4826) );
  AOI22_X1 U5871 ( .A1(n6584), .A2(n4883), .B1(n6431), .B2(n6516), .ZN(n4825)
         );
  OAI211_X1 U5872 ( .C1(n6524), .C2(n4886), .A(n4826), .B(n4825), .ZN(U3035)
         );
  AOI22_X1 U5873 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4879), .B1(n6559), 
        .B2(n4878), .ZN(n4828) );
  AOI22_X1 U5874 ( .A1(n6557), .A2(n4883), .B1(n6431), .B2(n6500), .ZN(n4827)
         );
  OAI211_X1 U5875 ( .C1(n6503), .C2(n4886), .A(n4828), .B(n4827), .ZN(U3031)
         );
  AOI22_X1 U5876 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4879), .B1(n6565), 
        .B2(n4878), .ZN(n4830) );
  AOI22_X1 U5877 ( .A1(n6563), .A2(n4883), .B1(n6431), .B2(n6460), .ZN(n4829)
         );
  OAI211_X1 U5878 ( .C1(n6463), .C2(n4886), .A(n4830), .B(n4829), .ZN(U3032)
         );
  AOI22_X1 U5879 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4953), .B1(n6541), 
        .B2(n4952), .ZN(n4832) );
  AOI22_X1 U5880 ( .A1(n5297), .A2(n6482), .B1(n6526), .B2(n4954), .ZN(n4831)
         );
  OAI211_X1 U5881 ( .C1(n5014), .C2(n6495), .A(n4832), .B(n4831), .ZN(U3092)
         );
  INV_X1 U5882 ( .A(n4833), .ZN(n6742) );
  NOR3_X1 U5883 ( .A1(n6743), .A2(n5263), .A3(n6742), .ZN(n6631) );
  INV_X1 U5884 ( .A(n6631), .ZN(n4835) );
  NAND3_X1 U5885 ( .A1(n6743), .A2(STATE2_REG_1__SCAN_IN), .A3(n4834), .ZN(
        n6643) );
  NAND2_X1 U5886 ( .A1(n4835), .A2(n6643), .ZN(n4836) );
  NOR2_X1 U5887 ( .A1(n6353), .A2(n4836), .ZN(n4837) );
  OR2_X1 U5888 ( .A1(n5518), .A2(n4839), .ZN(n4841) );
  NOR2_X1 U5889 ( .A1(n4842), .A2(n5452), .ZN(n4843) );
  INV_X1 U5890 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4852) );
  OAI22_X1 U5891 ( .A1(n6171), .A2(n4852), .B1(n6104), .B2(n5326), .ZN(n4851)
         );
  NAND2_X1 U5892 ( .A1(n4599), .A2(n6738), .ZN(n4855) );
  INV_X1 U5893 ( .A(n4855), .ZN(n4844) );
  NAND3_X1 U5894 ( .A1(n4846), .A2(n4845), .A3(n4844), .ZN(n4847) );
  NAND2_X1 U5895 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4855), .ZN(n4848) );
  OAI22_X1 U5896 ( .A1(n5516), .A2(REIP_REG_1__SCAN_IN), .B1(n5131), .B2(n4849), .ZN(n4850) );
  AOI211_X1 U5897 ( .C1(n6207), .C2(n4852), .A(n4851), .B(n4850), .ZN(n4861)
         );
  NOR2_X1 U5898 ( .A1(n5518), .A2(n4853), .ZN(n6196) );
  NOR2_X1 U5899 ( .A1(n6655), .A2(n4855), .ZN(n6625) );
  NOR2_X1 U5900 ( .A1(n4854), .A2(n6625), .ZN(n5519) );
  INV_X1 U5901 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U5902 ( .A1(n5613), .A2(n4855), .ZN(n4856) );
  NOR2_X1 U5903 ( .A1(n4857), .A2(n4856), .ZN(n4858) );
  NOR2_X1 U5904 ( .A1(n5519), .A2(n4858), .ZN(n4859) );
  INV_X2 U5905 ( .A(n6172), .ZN(n6198) );
  AOI22_X1 U5906 ( .A1(n4665), .A2(n6196), .B1(n6198), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4860) );
  OAI211_X1 U5907 ( .C1(n6205), .C2(n5233), .A(n4861), .B(n4860), .ZN(U2826)
         );
  INV_X1 U5908 ( .A(DATAI_29_), .ZN(n4862) );
  OR2_X1 U5909 ( .A1(n6292), .A2(n4862), .ZN(n6509) );
  NOR2_X2 U5910 ( .A1(n4863), .A2(n4877), .ZN(n6571) );
  AOI22_X1 U5911 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4879), .B1(n6571), 
        .B2(n4878), .ZN(n4867) );
  NOR2_X2 U5912 ( .A1(n4881), .A2(n4864), .ZN(n6569) );
  INV_X1 U5913 ( .A(DATAI_21_), .ZN(n4865) );
  OR2_X1 U5914 ( .A1(n6292), .A2(n4865), .ZN(n6574) );
  INV_X1 U5915 ( .A(n6574), .ZN(n6506) );
  AOI22_X1 U5916 ( .A1(n6569), .A2(n4883), .B1(n6431), .B2(n6506), .ZN(n4866)
         );
  OAI211_X1 U5917 ( .C1(n6509), .C2(n4886), .A(n4867), .B(n4866), .ZN(U3033)
         );
  INV_X1 U5918 ( .A(DATAI_30_), .ZN(n4868) );
  OR2_X1 U5919 ( .A1(n6292), .A2(n4868), .ZN(n6582) );
  INV_X1 U5920 ( .A(DATAI_6_), .ZN(n6868) );
  NOR2_X2 U5921 ( .A1(n6868), .A2(n4877), .ZN(n6578) );
  AOI22_X1 U5922 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4879), .B1(n6578), 
        .B2(n4878), .ZN(n4871) );
  NOR2_X2 U5923 ( .A1(n4881), .A2(n3861), .ZN(n6575) );
  INV_X1 U5924 ( .A(DATAI_22_), .ZN(n4869) );
  OR2_X1 U5925 ( .A1(n6292), .A2(n4869), .ZN(n6515) );
  INV_X1 U5926 ( .A(n6515), .ZN(n6576) );
  AOI22_X1 U5927 ( .A1(n6575), .A2(n4883), .B1(n6431), .B2(n6576), .ZN(n4870)
         );
  OAI211_X1 U5928 ( .C1(n6582), .C2(n4886), .A(n4871), .B(n4870), .ZN(U3034)
         );
  INV_X1 U5929 ( .A(DATAI_25_), .ZN(n4872) );
  OR2_X1 U5930 ( .A1(n6292), .A2(n4872), .ZN(n6550) );
  INV_X1 U5931 ( .A(DATAI_1_), .ZN(n7004) );
  NOR2_X2 U5932 ( .A1(n7004), .A2(n4877), .ZN(n6547) );
  AOI22_X1 U5933 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4879), .B1(n6547), 
        .B2(n4878), .ZN(n4875) );
  NOR2_X2 U5934 ( .A1(n4881), .A2(n4873), .ZN(n6545) );
  INV_X1 U5935 ( .A(DATAI_17_), .ZN(n7024) );
  OR2_X1 U5936 ( .A1(n6292), .A2(n7024), .ZN(n6418) );
  INV_X1 U5937 ( .A(n6418), .ZN(n6546) );
  AOI22_X1 U5938 ( .A1(n6545), .A2(n4883), .B1(n6431), .B2(n6546), .ZN(n4874)
         );
  OAI211_X1 U5939 ( .C1(n6550), .C2(n4886), .A(n4875), .B(n4874), .ZN(U3029)
         );
  INV_X1 U5940 ( .A(DATAI_26_), .ZN(n4876) );
  OR2_X1 U5941 ( .A1(n6292), .A2(n4876), .ZN(n6455) );
  NOR2_X2 U5942 ( .A1(n7055), .A2(n4877), .ZN(n6553) );
  AOI22_X1 U5943 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4879), .B1(n6553), 
        .B2(n4878), .ZN(n4885) );
  NOR2_X2 U5944 ( .A1(n4881), .A2(n4880), .ZN(n6551) );
  INV_X1 U5945 ( .A(DATAI_18_), .ZN(n4882) );
  OR2_X1 U5946 ( .A1(n6292), .A2(n4882), .ZN(n6556) );
  INV_X1 U5947 ( .A(n6556), .ZN(n6452) );
  AOI22_X1 U5948 ( .A1(n6551), .A2(n4883), .B1(n6431), .B2(n6452), .ZN(n4884)
         );
  OAI211_X1 U5949 ( .C1(n6455), .C2(n4886), .A(n4885), .B(n4884), .ZN(U3030)
         );
  NAND2_X1 U5950 ( .A1(n6601), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4971) );
  NOR2_X1 U5951 ( .A1(n6435), .A2(n4971), .ZN(n5176) );
  INV_X1 U5952 ( .A(n4665), .ZN(n5969) );
  NAND2_X1 U5953 ( .A1(n4560), .A2(n5969), .ZN(n5178) );
  INV_X1 U5954 ( .A(n5178), .ZN(n4887) );
  AND2_X1 U5955 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5176), .ZN(n4910)
         );
  AOI21_X1 U5956 ( .B1(n4916), .B2(n4887), .A(n4910), .ZN(n4892) );
  NAND3_X1 U5957 ( .A1(n6486), .A2(n4892), .A3(n4889), .ZN(n4888) );
  OAI211_X1 U5958 ( .C1(n6530), .C2(n5176), .A(n6488), .B(n4888), .ZN(n4909)
         );
  NAND2_X1 U5959 ( .A1(n6530), .A2(n4889), .ZN(n4891) );
  NAND2_X1 U5960 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4890) );
  OAI22_X1 U5961 ( .A1(n4892), .A2(n4891), .B1(n4971), .B2(n4890), .ZN(n4908)
         );
  AOI22_X1 U5962 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4909), .B1(n6588), 
        .B2(n4908), .ZN(n4895) );
  NOR2_X2 U5963 ( .A1(n4893), .A2(n4968), .ZN(n5222) );
  AOI22_X1 U5964 ( .A1(n6584), .A2(n4910), .B1(n6585), .B2(n5222), .ZN(n4894)
         );
  OAI211_X1 U5965 ( .C1(n6593), .C2(n5087), .A(n4895), .B(n4894), .ZN(U3131)
         );
  AOI22_X1 U5966 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4909), .B1(n6578), 
        .B2(n4908), .ZN(n4897) );
  INV_X1 U5967 ( .A(n6582), .ZN(n6510) );
  AOI22_X1 U5968 ( .A1(n6575), .A2(n4910), .B1(n6510), .B2(n5222), .ZN(n4896)
         );
  OAI211_X1 U5969 ( .C1(n6515), .C2(n5087), .A(n4897), .B(n4896), .ZN(U3130)
         );
  AOI22_X1 U5970 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4909), .B1(n6571), 
        .B2(n4908), .ZN(n4899) );
  INV_X1 U5971 ( .A(n6509), .ZN(n6570) );
  AOI22_X1 U5972 ( .A1(n6569), .A2(n4910), .B1(n6570), .B2(n5222), .ZN(n4898)
         );
  OAI211_X1 U5973 ( .C1(n6574), .C2(n5087), .A(n4899), .B(n4898), .ZN(U3129)
         );
  AOI22_X1 U5974 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4909), .B1(n6565), 
        .B2(n4908), .ZN(n4901) );
  AOI22_X1 U5975 ( .A1(n6563), .A2(n4910), .B1(n6564), .B2(n5222), .ZN(n4900)
         );
  OAI211_X1 U5976 ( .C1(n6568), .C2(n5087), .A(n4901), .B(n4900), .ZN(U3128)
         );
  AOI22_X1 U5977 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4909), .B1(n6559), 
        .B2(n4908), .ZN(n4903) );
  AOI22_X1 U5978 ( .A1(n6557), .A2(n4910), .B1(n6558), .B2(n5222), .ZN(n4902)
         );
  OAI211_X1 U5979 ( .C1(n6562), .C2(n5087), .A(n4903), .B(n4902), .ZN(U3127)
         );
  AOI22_X1 U5980 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4909), .B1(n6547), 
        .B2(n4908), .ZN(n4905) );
  INV_X1 U5981 ( .A(n6550), .ZN(n6415) );
  AOI22_X1 U5982 ( .A1(n6545), .A2(n4910), .B1(n6415), .B2(n5222), .ZN(n4904)
         );
  OAI211_X1 U5983 ( .C1(n6418), .C2(n5087), .A(n4905), .B(n4904), .ZN(U3125)
         );
  AOI22_X1 U5984 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4909), .B1(n6541), 
        .B2(n4908), .ZN(n4907) );
  INV_X1 U5985 ( .A(n6495), .ZN(n6527) );
  AOI22_X1 U5986 ( .A1(n6526), .A2(n4910), .B1(n6527), .B2(n5222), .ZN(n4906)
         );
  OAI211_X1 U5987 ( .C1(n6544), .C2(n5087), .A(n4907), .B(n4906), .ZN(U3124)
         );
  AOI22_X1 U5988 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4909), .B1(n6553), 
        .B2(n4908), .ZN(n4912) );
  INV_X1 U5989 ( .A(n6455), .ZN(n6552) );
  AOI22_X1 U5990 ( .A1(n6551), .A2(n4910), .B1(n6552), .B2(n5222), .ZN(n4911)
         );
  OAI211_X1 U5991 ( .C1(n6556), .C2(n5087), .A(n4912), .B(n4911), .ZN(U3126)
         );
  INV_X1 U5992 ( .A(n4913), .ZN(n4914) );
  OAI21_X1 U5993 ( .B1(n4914), .B2(n6292), .A(n6409), .ZN(n4919) );
  INV_X1 U5994 ( .A(n4915), .ZN(n5069) );
  AOI21_X1 U5995 ( .B1(n4916), .B2(n6485), .A(n5069), .ZN(n4921) );
  OAI21_X1 U5996 ( .B1(n6486), .B2(n4917), .A(n6488), .ZN(n4918) );
  AOI21_X1 U5997 ( .B1(n4919), .B2(n4921), .A(n4918), .ZN(n5074) );
  INV_X1 U5998 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4925) );
  OAI22_X1 U5999 ( .A1(n4921), .A2(n6535), .B1(n4920), .B2(n6737), .ZN(n5068)
         );
  AOI22_X1 U6000 ( .A1(n6526), .A2(n5069), .B1(n6541), .B2(n5068), .ZN(n4922)
         );
  OAI21_X1 U6001 ( .B1(n6544), .B2(n5078), .A(n4922), .ZN(n4923) );
  AOI21_X1 U6002 ( .B1(n6527), .B2(n5089), .A(n4923), .ZN(n4924) );
  OAI21_X1 U6003 ( .B1(n5074), .B2(n4925), .A(n4924), .ZN(U3140) );
  INV_X1 U6004 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4929) );
  AOI22_X1 U6005 ( .A1(n6563), .A2(n5069), .B1(n6565), .B2(n5068), .ZN(n4926)
         );
  OAI21_X1 U6006 ( .B1(n6568), .B2(n5078), .A(n4926), .ZN(n4927) );
  AOI21_X1 U6007 ( .B1(n6564), .B2(n5089), .A(n4927), .ZN(n4928) );
  OAI21_X1 U6008 ( .B1(n5074), .B2(n4929), .A(n4928), .ZN(U3144) );
  INV_X1 U6009 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4933) );
  AOI22_X1 U6010 ( .A1(n6584), .A2(n5069), .B1(n6588), .B2(n5068), .ZN(n4930)
         );
  OAI21_X1 U6011 ( .B1(n6593), .B2(n5078), .A(n4930), .ZN(n4931) );
  AOI21_X1 U6012 ( .B1(n6585), .B2(n5089), .A(n4931), .ZN(n4932) );
  OAI21_X1 U6013 ( .B1(n5074), .B2(n4933), .A(n4932), .ZN(U3147) );
  INV_X1 U6014 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4937) );
  AOI22_X1 U6015 ( .A1(n6557), .A2(n5069), .B1(n6559), .B2(n5068), .ZN(n4934)
         );
  OAI21_X1 U6016 ( .B1(n6562), .B2(n5078), .A(n4934), .ZN(n4935) );
  AOI21_X1 U6017 ( .B1(n6558), .B2(n5089), .A(n4935), .ZN(n4936) );
  OAI21_X1 U6018 ( .B1(n5074), .B2(n4937), .A(n4936), .ZN(U3143) );
  NAND2_X1 U6019 ( .A1(n4940), .A2(n4939), .ZN(n4941) );
  XNOR2_X1 U6020 ( .A(n4938), .B(n4941), .ZN(n6330) );
  NAND2_X1 U6021 ( .A1(n6330), .A2(n6303), .ZN(n4945) );
  INV_X1 U6022 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4942) );
  NAND2_X1 U6023 ( .A1(n6353), .A2(REIP_REG_9__SCAN_IN), .ZN(n6326) );
  OAI21_X1 U6024 ( .B1(n6063), .B2(n4942), .A(n6326), .ZN(n4943) );
  AOI21_X1 U6025 ( .B1(n6276), .B2(n6166), .A(n4943), .ZN(n4944) );
  OAI211_X1 U6026 ( .C1(n6292), .C2(n6165), .A(n4945), .B(n4944), .ZN(U2977)
         );
  AOI22_X1 U6027 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4953), .B1(n6553), 
        .B2(n4952), .ZN(n4947) );
  AOI22_X1 U6028 ( .A1(n5297), .A2(n6452), .B1(n4954), .B2(n6551), .ZN(n4946)
         );
  OAI211_X1 U6029 ( .C1(n5014), .C2(n6455), .A(n4947), .B(n4946), .ZN(U3094)
         );
  AOI22_X1 U6030 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4953), .B1(n6571), 
        .B2(n4952), .ZN(n4949) );
  AOI22_X1 U6031 ( .A1(n5297), .A2(n6506), .B1(n4954), .B2(n6569), .ZN(n4948)
         );
  OAI211_X1 U6032 ( .C1(n5014), .C2(n6509), .A(n4949), .B(n4948), .ZN(U3097)
         );
  AOI22_X1 U6033 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4953), .B1(n6578), 
        .B2(n4952), .ZN(n4951) );
  AOI22_X1 U6034 ( .A1(n5297), .A2(n6576), .B1(n4954), .B2(n6575), .ZN(n4950)
         );
  OAI211_X1 U6035 ( .C1(n5014), .C2(n6582), .A(n4951), .B(n4950), .ZN(U3098)
         );
  AOI22_X1 U6036 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4953), .B1(n6547), 
        .B2(n4952), .ZN(n4956) );
  AOI22_X1 U6037 ( .A1(n5297), .A2(n6546), .B1(n4954), .B2(n6545), .ZN(n4955)
         );
  OAI211_X1 U6038 ( .C1(n5014), .C2(n6550), .A(n4956), .B(n4955), .ZN(U3093)
         );
  INV_X1 U6039 ( .A(n5311), .ZN(n4965) );
  NOR2_X1 U6040 ( .A1(n6342), .A2(n4961), .ZN(n6320) );
  NOR2_X1 U6041 ( .A1(n6386), .A2(n6377), .ZN(n6369) );
  NAND3_X1 U6042 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6369), .ZN(n4958) );
  AOI21_X1 U6043 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6394) );
  INV_X1 U6044 ( .A(n6394), .ZN(n6344) );
  NOR2_X1 U6045 ( .A1(n6398), .A2(n6852), .ZN(n6393) );
  NAND2_X1 U6046 ( .A1(n6393), .A2(n6399), .ZN(n6361) );
  NAND2_X1 U6047 ( .A1(n5814), .A2(n6361), .ZN(n6345) );
  NAND2_X1 U6048 ( .A1(n6344), .A2(n6345), .ZN(n6387) );
  NOR2_X1 U6049 ( .A1(n4958), .A2(n6387), .ZN(n6338) );
  OAI21_X1 U6050 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6338), .ZN(n4962) );
  NAND2_X1 U6051 ( .A1(n5814), .A2(n6347), .ZN(n5804) );
  INV_X1 U6052 ( .A(n4958), .ZN(n4959) );
  NAND3_X1 U6053 ( .A1(n6392), .A2(n4959), .A3(n6344), .ZN(n5343) );
  INV_X1 U6054 ( .A(n6348), .ZN(n4960) );
  NAND2_X1 U6055 ( .A1(n4959), .A2(n6393), .ZN(n5344) );
  AOI22_X1 U6056 ( .A1(n5804), .A2(n5343), .B1(n4960), .B2(n5344), .ZN(n6343)
         );
  OAI22_X1 U6057 ( .A1(n6320), .A2(n4962), .B1(n6343), .B2(n4961), .ZN(n4963)
         );
  AOI211_X1 U6058 ( .C1(n6383), .C2(n4965), .A(n4964), .B(n4963), .ZN(n4966)
         );
  OAI21_X1 U6059 ( .B1(n6370), .B2(n4967), .A(n4966), .ZN(U3010) );
  AND2_X1 U6060 ( .A1(n4585), .A2(n5175), .ZN(n4970) );
  NAND2_X1 U6061 ( .A1(n4970), .A2(n3887), .ZN(n6459) );
  INV_X1 U6062 ( .A(n6557), .ZN(n5189) );
  OR2_X1 U6063 ( .A1(n4971), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5099)
         );
  NOR2_X1 U6064 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5099), .ZN(n4981)
         );
  INV_X1 U6065 ( .A(n4981), .ZN(n5146) );
  NAND2_X1 U6066 ( .A1(n6407), .A2(n6486), .ZN(n4974) );
  INV_X1 U6067 ( .A(n5261), .ZN(n4973) );
  OAI22_X1 U6068 ( .A1(n4974), .A2(n5178), .B1(n4973), .B2(n4972), .ZN(n5144)
         );
  NAND2_X1 U6069 ( .A1(n5149), .A2(n6459), .ZN(n4977) );
  OAI21_X1 U6070 ( .B1(n5178), .B2(n4975), .A(n6530), .ZN(n4976) );
  AOI21_X1 U6071 ( .B1(n4977), .B2(STATEBS16_REG_SCAN_IN), .A(n4976), .ZN(
        n4978) );
  NOR3_X1 U6072 ( .A1(n4979), .A2(n5259), .A3(n4978), .ZN(n4980) );
  OAI21_X1 U6073 ( .B1(n4981), .B2(n5263), .A(n4980), .ZN(n5143) );
  AOI22_X1 U6074 ( .A1(n5144), .A2(n6559), .B1(INSTQUEUE_REG_4__3__SCAN_IN), 
        .B2(n5143), .ZN(n4982) );
  OAI21_X1 U6075 ( .B1(n5189), .B2(n5146), .A(n4982), .ZN(n4983) );
  AOI21_X1 U6076 ( .B1(n6558), .B2(n6468), .A(n4983), .ZN(n4984) );
  OAI21_X1 U6077 ( .B1(n6562), .B2(n5149), .A(n4984), .ZN(U3055) );
  INV_X1 U6078 ( .A(n6526), .ZN(n5201) );
  AOI22_X1 U6079 ( .A1(n5144), .A2(n6541), .B1(INSTQUEUE_REG_4__0__SCAN_IN), 
        .B2(n5143), .ZN(n4985) );
  OAI21_X1 U6080 ( .B1(n5201), .B2(n5146), .A(n4985), .ZN(n4986) );
  AOI21_X1 U6081 ( .B1(n6527), .B2(n6468), .A(n4986), .ZN(n4987) );
  OAI21_X1 U6082 ( .B1(n6544), .B2(n5149), .A(n4987), .ZN(U3052) );
  INV_X1 U6083 ( .A(n6563), .ZN(n5193) );
  AOI22_X1 U6084 ( .A1(n5144), .A2(n6565), .B1(INSTQUEUE_REG_4__4__SCAN_IN), 
        .B2(n5143), .ZN(n4988) );
  OAI21_X1 U6085 ( .B1(n5193), .B2(n5146), .A(n4988), .ZN(n4989) );
  AOI21_X1 U6086 ( .B1(n6564), .B2(n6468), .A(n4989), .ZN(n4990) );
  OAI21_X1 U6087 ( .B1(n6568), .B2(n5149), .A(n4990), .ZN(U3056) );
  INV_X1 U6088 ( .A(n6584), .ZN(n5197) );
  AOI22_X1 U6089 ( .A1(n5144), .A2(n6588), .B1(INSTQUEUE_REG_4__7__SCAN_IN), 
        .B2(n5143), .ZN(n4991) );
  OAI21_X1 U6090 ( .B1(n5197), .B2(n5146), .A(n4991), .ZN(n4992) );
  AOI21_X1 U6091 ( .B1(n6585), .B2(n6468), .A(n4992), .ZN(n4993) );
  OAI21_X1 U6092 ( .B1(n6593), .B2(n5149), .A(n4993), .ZN(U3059) );
  OAI21_X1 U6093 ( .B1(n4735), .B2(n3979), .A(n4996), .ZN(n5324) );
  AOI22_X1 U6094 ( .A1(n6236), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6230), .ZN(n4997) );
  OAI21_X1 U6095 ( .B1(n5324), .B2(n5697), .A(n4997), .ZN(U2881) );
  AOI22_X1 U6096 ( .A1(n6569), .A2(n5011), .B1(n6571), .B2(n5010), .ZN(n4999)
         );
  OR2_X1 U6097 ( .A1(n6514), .A2(n6509), .ZN(n4998) );
  OAI211_X1 U6098 ( .C1(n6574), .C2(n5014), .A(n4999), .B(n4998), .ZN(n5000)
         );
  AOI21_X1 U6099 ( .B1(n5016), .B2(INSTQUEUE_REG_8__5__SCAN_IN), .A(n5000), 
        .ZN(n5001) );
  INV_X1 U6100 ( .A(n5001), .ZN(U3089) );
  AOI22_X1 U6101 ( .A1(n6575), .A2(n5011), .B1(n6578), .B2(n5010), .ZN(n5003)
         );
  OR2_X1 U6102 ( .A1(n6514), .A2(n6582), .ZN(n5002) );
  OAI211_X1 U6103 ( .C1(n6515), .C2(n5014), .A(n5003), .B(n5002), .ZN(n5004)
         );
  AOI21_X1 U6104 ( .B1(n5016), .B2(INSTQUEUE_REG_8__6__SCAN_IN), .A(n5004), 
        .ZN(n5005) );
  INV_X1 U6105 ( .A(n5005), .ZN(U3090) );
  AOI22_X1 U6106 ( .A1(n6545), .A2(n5011), .B1(n6547), .B2(n5010), .ZN(n5007)
         );
  OR2_X1 U6107 ( .A1(n6514), .A2(n6550), .ZN(n5006) );
  OAI211_X1 U6108 ( .C1(n6418), .C2(n5014), .A(n5007), .B(n5006), .ZN(n5008)
         );
  AOI21_X1 U6109 ( .B1(n5016), .B2(INSTQUEUE_REG_8__1__SCAN_IN), .A(n5008), 
        .ZN(n5009) );
  INV_X1 U6110 ( .A(n5009), .ZN(U3085) );
  AOI22_X1 U6111 ( .A1(n6551), .A2(n5011), .B1(n6553), .B2(n5010), .ZN(n5013)
         );
  OR2_X1 U6112 ( .A1(n6514), .A2(n6455), .ZN(n5012) );
  OAI211_X1 U6113 ( .C1(n6556), .C2(n5014), .A(n5013), .B(n5012), .ZN(n5015)
         );
  AOI21_X1 U6114 ( .B1(n5016), .B2(INSTQUEUE_REG_8__2__SCAN_IN), .A(n5015), 
        .ZN(n5017) );
  INV_X1 U6115 ( .A(n5017), .ZN(U3086) );
  INV_X1 U6116 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5021) );
  AOI22_X1 U6117 ( .A1(n6575), .A2(n6476), .B1(n6578), .B2(n6475), .ZN(n5018)
         );
  OAI21_X1 U6118 ( .B1(n6515), .B2(n6523), .A(n5018), .ZN(n5019) );
  AOI21_X1 U6119 ( .B1(n6510), .B2(n6477), .A(n5019), .ZN(n5020) );
  OAI21_X1 U6120 ( .B1(n5067), .B2(n5021), .A(n5020), .ZN(U3074) );
  AOI22_X1 U6121 ( .A1(n6545), .A2(n5076), .B1(n6547), .B2(n5075), .ZN(n5022)
         );
  OAI21_X1 U6122 ( .B1(n6550), .B2(n5078), .A(n5022), .ZN(n5023) );
  AOI21_X1 U6123 ( .B1(n6546), .B2(n5080), .A(n5023), .ZN(n5024) );
  OAI21_X1 U6124 ( .B1(n5083), .B2(n5025), .A(n5024), .ZN(U3021) );
  AOI22_X1 U6125 ( .A1(n6551), .A2(n6476), .B1(n6553), .B2(n6475), .ZN(n5026)
         );
  OAI21_X1 U6126 ( .B1(n6556), .B2(n6523), .A(n5026), .ZN(n5027) );
  AOI21_X1 U6127 ( .B1(n6552), .B2(n6477), .A(n5027), .ZN(n5028) );
  OAI21_X1 U6128 ( .B1(n5067), .B2(n6948), .A(n5028), .ZN(U3070) );
  AOI22_X1 U6129 ( .A1(n6551), .A2(n5076), .B1(n6553), .B2(n5075), .ZN(n5029)
         );
  OAI21_X1 U6130 ( .B1(n6455), .B2(n5078), .A(n5029), .ZN(n5030) );
  AOI21_X1 U6131 ( .B1(n6452), .B2(n5080), .A(n5030), .ZN(n5031) );
  OAI21_X1 U6132 ( .B1(n5083), .B2(n5032), .A(n5031), .ZN(U3022) );
  INV_X1 U6133 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5036) );
  AOI22_X1 U6134 ( .A1(n6545), .A2(n6476), .B1(n6547), .B2(n6475), .ZN(n5033)
         );
  OAI21_X1 U6135 ( .B1(n6418), .B2(n6523), .A(n5033), .ZN(n5034) );
  AOI21_X1 U6136 ( .B1(n6415), .B2(n6477), .A(n5034), .ZN(n5035) );
  OAI21_X1 U6137 ( .B1(n5067), .B2(n5036), .A(n5035), .ZN(U3069) );
  AOI22_X1 U6138 ( .A1(n6575), .A2(n5076), .B1(n6578), .B2(n5075), .ZN(n5037)
         );
  OAI21_X1 U6139 ( .B1(n6582), .B2(n5078), .A(n5037), .ZN(n5038) );
  AOI21_X1 U6140 ( .B1(n6576), .B2(n5080), .A(n5038), .ZN(n5039) );
  OAI21_X1 U6141 ( .B1(n5083), .B2(n5040), .A(n5039), .ZN(U3026) );
  INV_X1 U6142 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5044) );
  AOI22_X1 U6143 ( .A1(n6551), .A2(n5069), .B1(n6553), .B2(n5068), .ZN(n5041)
         );
  OAI21_X1 U6144 ( .B1(n6556), .B2(n5078), .A(n5041), .ZN(n5042) );
  AOI21_X1 U6145 ( .B1(n6552), .B2(n5089), .A(n5042), .ZN(n5043) );
  OAI21_X1 U6146 ( .B1(n5074), .B2(n5044), .A(n5043), .ZN(U3142) );
  INV_X1 U6147 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5048) );
  AOI22_X1 U6148 ( .A1(n6551), .A2(n5085), .B1(n6553), .B2(n5084), .ZN(n5045)
         );
  OAI21_X1 U6149 ( .B1(n6455), .B2(n5087), .A(n5045), .ZN(n5046) );
  AOI21_X1 U6150 ( .B1(n6452), .B2(n5089), .A(n5046), .ZN(n5047) );
  OAI21_X1 U6151 ( .B1(n5092), .B2(n5048), .A(n5047), .ZN(U3134) );
  INV_X1 U6152 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5052) );
  AOI22_X1 U6153 ( .A1(n6575), .A2(n5069), .B1(n6578), .B2(n5068), .ZN(n5049)
         );
  OAI21_X1 U6154 ( .B1(n6515), .B2(n5078), .A(n5049), .ZN(n5050) );
  AOI21_X1 U6155 ( .B1(n6510), .B2(n5089), .A(n5050), .ZN(n5051) );
  OAI21_X1 U6156 ( .B1(n5074), .B2(n5052), .A(n5051), .ZN(U3146) );
  AOI22_X1 U6157 ( .A1(n6575), .A2(n5085), .B1(n6578), .B2(n5084), .ZN(n5053)
         );
  OAI21_X1 U6158 ( .B1(n6582), .B2(n5087), .A(n5053), .ZN(n5054) );
  AOI21_X1 U6159 ( .B1(n6576), .B2(n5089), .A(n5054), .ZN(n5055) );
  OAI21_X1 U6160 ( .B1(n5092), .B2(n7005), .A(n5055), .ZN(U3138) );
  AOI22_X1 U6161 ( .A1(n6545), .A2(n5069), .B1(n6547), .B2(n5068), .ZN(n5056)
         );
  OAI21_X1 U6162 ( .B1(n6418), .B2(n5078), .A(n5056), .ZN(n5057) );
  AOI21_X1 U6163 ( .B1(n6415), .B2(n5089), .A(n5057), .ZN(n5058) );
  OAI21_X1 U6164 ( .B1(n5074), .B2(n7037), .A(n5058), .ZN(U3141) );
  INV_X1 U6165 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5062) );
  AOI22_X1 U6166 ( .A1(n6545), .A2(n5085), .B1(n6547), .B2(n5084), .ZN(n5059)
         );
  OAI21_X1 U6167 ( .B1(n6550), .B2(n5087), .A(n5059), .ZN(n5060) );
  AOI21_X1 U6168 ( .B1(n6546), .B2(n5089), .A(n5060), .ZN(n5061) );
  OAI21_X1 U6169 ( .B1(n5092), .B2(n5062), .A(n5061), .ZN(U3133) );
  INV_X1 U6170 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5066) );
  AOI22_X1 U6171 ( .A1(n6569), .A2(n6476), .B1(n6571), .B2(n6475), .ZN(n5063)
         );
  OAI21_X1 U6172 ( .B1(n6574), .B2(n6523), .A(n5063), .ZN(n5064) );
  AOI21_X1 U6173 ( .B1(n6570), .B2(n6477), .A(n5064), .ZN(n5065) );
  OAI21_X1 U6174 ( .B1(n5067), .B2(n5066), .A(n5065), .ZN(U3073) );
  INV_X1 U6175 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5073) );
  AOI22_X1 U6176 ( .A1(n6569), .A2(n5069), .B1(n6571), .B2(n5068), .ZN(n5070)
         );
  OAI21_X1 U6177 ( .B1(n6574), .B2(n5078), .A(n5070), .ZN(n5071) );
  AOI21_X1 U6178 ( .B1(n6570), .B2(n5089), .A(n5071), .ZN(n5072) );
  OAI21_X1 U6179 ( .B1(n5074), .B2(n5073), .A(n5072), .ZN(U3145) );
  AOI22_X1 U6180 ( .A1(n6569), .A2(n5076), .B1(n6571), .B2(n5075), .ZN(n5077)
         );
  OAI21_X1 U6181 ( .B1(n6509), .B2(n5078), .A(n5077), .ZN(n5079) );
  AOI21_X1 U6182 ( .B1(n6506), .B2(n5080), .A(n5079), .ZN(n5081) );
  OAI21_X1 U6183 ( .B1(n5083), .B2(n5082), .A(n5081), .ZN(U3025) );
  INV_X1 U6184 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5091) );
  AOI22_X1 U6185 ( .A1(n6569), .A2(n5085), .B1(n6571), .B2(n5084), .ZN(n5086)
         );
  OAI21_X1 U6186 ( .B1(n6509), .B2(n5087), .A(n5086), .ZN(n5088) );
  AOI21_X1 U6187 ( .B1(n6506), .B2(n5089), .A(n5088), .ZN(n5090) );
  OAI21_X1 U6188 ( .B1(n5092), .B2(n5091), .A(n5090), .ZN(U3137) );
  OAI21_X1 U6189 ( .B1(n5094), .B2(n5093), .A(n6530), .ZN(n5102) );
  NAND2_X1 U6190 ( .A1(n6597), .A2(n5095), .ZN(n6483) );
  OR2_X1 U6191 ( .A1(n5178), .A2(n6483), .ZN(n5097) );
  NOR2_X1 U6192 ( .A1(n5177), .A2(n5099), .ZN(n5119) );
  INV_X1 U6193 ( .A(n5119), .ZN(n5096) );
  AND2_X1 U6194 ( .A1(n5097), .A2(n5096), .ZN(n5098) );
  OAI22_X1 U6195 ( .A1(n5102), .A2(n5098), .B1(n5099), .B2(n6737), .ZN(n5118)
         );
  INV_X1 U6196 ( .A(n5098), .ZN(n5101) );
  INV_X1 U6197 ( .A(n6488), .ZN(n6534) );
  AOI21_X1 U6198 ( .B1(n5099), .B2(n6535), .A(n6534), .ZN(n5100) );
  OAI21_X1 U6199 ( .B1(n5102), .B2(n5101), .A(n5100), .ZN(n5117) );
  AOI22_X1 U6200 ( .A1(n6565), .A2(n5118), .B1(n5117), .B2(
        INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5104) );
  AOI22_X1 U6201 ( .A1(n6564), .A2(n5120), .B1(n6563), .B2(n5119), .ZN(n5103)
         );
  OAI211_X1 U6202 ( .C1(n6568), .C2(n5123), .A(n5104), .B(n5103), .ZN(U3064)
         );
  AOI22_X1 U6203 ( .A1(n6547), .A2(n5118), .B1(n5117), .B2(
        INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n5106) );
  AOI22_X1 U6204 ( .A1(n6415), .A2(n5120), .B1(n6545), .B2(n5119), .ZN(n5105)
         );
  OAI211_X1 U6205 ( .C1(n6418), .C2(n5123), .A(n5106), .B(n5105), .ZN(U3061)
         );
  AOI22_X1 U6206 ( .A1(n6571), .A2(n5118), .B1(n5117), .B2(
        INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5108) );
  AOI22_X1 U6207 ( .A1(n6570), .A2(n5120), .B1(n6569), .B2(n5119), .ZN(n5107)
         );
  OAI211_X1 U6208 ( .C1(n6574), .C2(n5123), .A(n5108), .B(n5107), .ZN(U3065)
         );
  AOI22_X1 U6209 ( .A1(n6578), .A2(n5118), .B1(n5117), .B2(
        INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5110) );
  AOI22_X1 U6210 ( .A1(n6510), .A2(n5120), .B1(n6575), .B2(n5119), .ZN(n5109)
         );
  OAI211_X1 U6211 ( .C1(n6515), .C2(n5123), .A(n5110), .B(n5109), .ZN(U3066)
         );
  AOI22_X1 U6212 ( .A1(n6588), .A2(n5118), .B1(n5117), .B2(
        INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5112) );
  AOI22_X1 U6213 ( .A1(n6585), .A2(n5120), .B1(n6584), .B2(n5119), .ZN(n5111)
         );
  OAI211_X1 U6214 ( .C1(n6593), .C2(n5123), .A(n5112), .B(n5111), .ZN(U3067)
         );
  AOI22_X1 U6215 ( .A1(n6553), .A2(n5118), .B1(n5117), .B2(
        INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5114) );
  AOI22_X1 U6216 ( .A1(n6552), .A2(n5120), .B1(n6551), .B2(n5119), .ZN(n5113)
         );
  OAI211_X1 U6217 ( .C1(n6556), .C2(n5123), .A(n5114), .B(n5113), .ZN(U3062)
         );
  AOI22_X1 U6218 ( .A1(n6559), .A2(n5118), .B1(n5117), .B2(
        INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5116) );
  AOI22_X1 U6219 ( .A1(n6558), .A2(n5120), .B1(n6557), .B2(n5119), .ZN(n5115)
         );
  OAI211_X1 U6220 ( .C1(n6562), .C2(n5123), .A(n5116), .B(n5115), .ZN(U3063)
         );
  AOI22_X1 U6221 ( .A1(n6541), .A2(n5118), .B1(n5117), .B2(
        INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5122) );
  AOI22_X1 U6222 ( .A1(n6527), .A2(n5120), .B1(n6526), .B2(n5119), .ZN(n5121)
         );
  OAI211_X1 U6223 ( .C1(n6544), .C2(n5123), .A(n5122), .B(n5121), .ZN(U3060)
         );
  INV_X1 U6224 ( .A(n6551), .ZN(n5220) );
  AOI22_X1 U6225 ( .A1(n5144), .A2(n6553), .B1(INSTQUEUE_REG_4__2__SCAN_IN), 
        .B2(n5143), .ZN(n5124) );
  OAI21_X1 U6226 ( .B1(n5220), .B2(n5146), .A(n5124), .ZN(n5125) );
  AOI21_X1 U6227 ( .B1(n6552), .B2(n6468), .A(n5125), .ZN(n5126) );
  OAI21_X1 U6228 ( .B1(n6556), .B2(n5149), .A(n5126), .ZN(U3054) );
  INV_X1 U6229 ( .A(n6575), .ZN(n5213) );
  AOI22_X1 U6230 ( .A1(n5144), .A2(n6578), .B1(INSTQUEUE_REG_4__6__SCAN_IN), 
        .B2(n5143), .ZN(n5127) );
  OAI21_X1 U6231 ( .B1(n5213), .B2(n5146), .A(n5127), .ZN(n5128) );
  AOI21_X1 U6232 ( .B1(n6510), .B2(n6468), .A(n5128), .ZN(n5129) );
  OAI21_X1 U6233 ( .B1(n6515), .B2(n5149), .A(n5129), .ZN(U3058) );
  OAI21_X1 U6234 ( .B1(n5516), .B2(REIP_REG_1__SCAN_IN), .A(n5326), .ZN(n6195)
         );
  AOI22_X1 U6235 ( .A1(n6196), .A2(n4560), .B1(n6198), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n5136) );
  INV_X1 U6236 ( .A(n6307), .ZN(n5130) );
  AOI22_X1 U6237 ( .A1(n6197), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6207), 
        .B2(n5130), .ZN(n5135) );
  NOR2_X2 U6238 ( .A1(n5131), .A2(n4434), .ZN(n6202) );
  NAND2_X1 U6239 ( .A1(n6202), .A2(n5132), .ZN(n5134) );
  INV_X1 U6240 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6194) );
  NAND3_X1 U6241 ( .A1(n5418), .A2(REIP_REG_1__SCAN_IN), .A3(n6194), .ZN(n5133) );
  NAND4_X1 U6242 ( .A1(n5136), .A2(n5135), .A3(n5134), .A4(n5133), .ZN(n5137)
         );
  AOI21_X1 U6243 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6195), .A(n5137), .ZN(n5138)
         );
  OAI21_X1 U6244 ( .B1(n6205), .B2(n5139), .A(n5138), .ZN(U2825) );
  INV_X1 U6245 ( .A(n6545), .ZN(n5205) );
  AOI22_X1 U6246 ( .A1(n5144), .A2(n6547), .B1(INSTQUEUE_REG_4__1__SCAN_IN), 
        .B2(n5143), .ZN(n5140) );
  OAI21_X1 U6247 ( .B1(n5205), .B2(n5146), .A(n5140), .ZN(n5141) );
  AOI21_X1 U6248 ( .B1(n6415), .B2(n6468), .A(n5141), .ZN(n5142) );
  OAI21_X1 U6249 ( .B1(n6418), .B2(n5149), .A(n5142), .ZN(U3053) );
  INV_X1 U6250 ( .A(n6569), .ZN(n5209) );
  AOI22_X1 U6251 ( .A1(n5144), .A2(n6571), .B1(INSTQUEUE_REG_4__5__SCAN_IN), 
        .B2(n5143), .ZN(n5145) );
  OAI21_X1 U6252 ( .B1(n5209), .B2(n5146), .A(n5145), .ZN(n5147) );
  AOI21_X1 U6253 ( .B1(n6570), .B2(n6468), .A(n5147), .ZN(n5148) );
  OAI21_X1 U6254 ( .B1(n6574), .B2(n5149), .A(n5148), .ZN(U3057) );
  INV_X1 U6255 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6883) );
  NAND2_X1 U6256 ( .A1(n5495), .A2(n6883), .ZN(n5152) );
  NAND2_X1 U6257 ( .A1(n5605), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5150)
         );
  OAI211_X1 U6258 ( .C1(n4434), .C2(EBX_REG_9__SCAN_IN), .A(n5150), .B(n5153), 
        .ZN(n5151) );
  NAND2_X1 U6259 ( .A1(n5152), .A2(n5151), .ZN(n6158) );
  MUX2_X1 U6260 ( .A(n5502), .B(n5153), .S(EBX_REG_10__SCAN_IN), .Z(n5157) );
  INV_X1 U6261 ( .A(n5153), .ZN(n5154) );
  NAND2_X1 U6262 ( .A1(n5154), .A2(n4434), .ZN(n5464) );
  NAND2_X1 U6263 ( .A1(n4434), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5155) );
  AND2_X1 U6264 ( .A1(n5464), .A2(n5155), .ZN(n5156) );
  NAND2_X1 U6265 ( .A1(n5157), .A2(n5156), .ZN(n5241) );
  INV_X1 U6266 ( .A(n5241), .ZN(n5237) );
  XNOR2_X1 U6267 ( .A(n6161), .B(n5237), .ZN(n6317) );
  INV_X1 U6268 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5158) );
  OAI222_X1 U6269 ( .A1(n5324), .A2(n5680), .B1(n5678), .B2(n6317), .C1(n5158), 
        .C2(n6221), .ZN(U2849) );
  NAND2_X1 U6270 ( .A1(n6269), .A2(n5160), .ZN(n5161) );
  XNOR2_X1 U6271 ( .A(n5159), .B(n5161), .ZN(n6322) );
  NAND2_X1 U6272 ( .A1(n6322), .A2(n6303), .ZN(n5164) );
  AND2_X1 U6273 ( .A1(n6353), .A2(REIP_REG_10__SCAN_IN), .ZN(n6318) );
  NOR2_X1 U6274 ( .A1(n6308), .A2(n5317), .ZN(n5162) );
  AOI211_X1 U6275 ( .C1(n6299), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6318), 
        .B(n5162), .ZN(n5163) );
  OAI211_X1 U6276 ( .C1(n6292), .C2(n5324), .A(n5164), .B(n5163), .ZN(U2976)
         );
  NAND2_X1 U6277 ( .A1(REIP_REG_5__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .ZN(
        n5249) );
  INV_X1 U6278 ( .A(n5249), .ZN(n5307) );
  INV_X1 U6279 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6667) );
  NOR3_X1 U6280 ( .A1(n6104), .A2(n6667), .A3(n6194), .ZN(n5308) );
  AND2_X1 U6281 ( .A1(n5326), .A2(n5308), .ZN(n6184) );
  NAND2_X1 U6282 ( .A1(n5516), .A2(n5326), .ZN(n6132) );
  INV_X1 U6283 ( .A(n6132), .ZN(n6185) );
  AOI21_X1 U6284 ( .B1(n5307), .B2(n6184), .A(n6185), .ZN(n6176) );
  INV_X1 U6285 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6669) );
  NAND2_X1 U6286 ( .A1(n5418), .A2(n5308), .ZN(n6187) );
  INV_X1 U6287 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6671) );
  OAI21_X1 U6288 ( .B1(n6669), .B2(n6187), .A(n6671), .ZN(n5165) );
  NAND2_X1 U6289 ( .A1(n6176), .A2(n5165), .ZN(n5173) );
  NAND2_X1 U6290 ( .A1(n5166), .A2(n5326), .ZN(n6186) );
  OAI22_X1 U6291 ( .A1(n5167), .A2(n6171), .B1(n6193), .B2(n6358), .ZN(n5168)
         );
  NOR2_X1 U6292 ( .A1(n6175), .A2(n5168), .ZN(n5169) );
  OAI21_X1 U6293 ( .B1(n6188), .B2(n5170), .A(n5169), .ZN(n5171) );
  AOI21_X1 U6294 ( .B1(EBX_REG_5__SCAN_IN), .B2(n6198), .A(n5171), .ZN(n5172)
         );
  OAI211_X1 U6295 ( .C1(n6205), .C2(n5174), .A(n5173), .B(n5172), .ZN(U2822)
         );
  NAND2_X1 U6296 ( .A1(n5177), .A2(n5176), .ZN(n5219) );
  NOR2_X1 U6297 ( .A1(n6407), .A2(n5178), .ZN(n5182) );
  AOI22_X1 U6298 ( .A1(n5182), .A2(n6530), .B1(n5261), .B2(n5179), .ZN(n5180)
         );
  INV_X1 U6299 ( .A(n5222), .ZN(n5181) );
  AOI21_X1 U6300 ( .B1(n5181), .B2(n6592), .A(n6738), .ZN(n5183) );
  NOR3_X1 U6301 ( .A1(n5183), .A2(n5182), .A3(n6535), .ZN(n5184) );
  AOI211_X1 U6302 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5219), .A(n5185), .B(
        n5184), .ZN(n5187) );
  NAND2_X1 U6303 ( .A1(n5187), .A2(n5186), .ZN(n5216) );
  AOI22_X1 U6304 ( .A1(n5217), .A2(n6559), .B1(INSTQUEUE_REG_12__3__SCAN_IN), 
        .B2(n5216), .ZN(n5188) );
  OAI21_X1 U6305 ( .B1(n5189), .B2(n5219), .A(n5188), .ZN(n5190) );
  AOI21_X1 U6306 ( .B1(n6500), .B2(n5222), .A(n5190), .ZN(n5191) );
  OAI21_X1 U6307 ( .B1(n6503), .B2(n6592), .A(n5191), .ZN(U3119) );
  AOI22_X1 U6308 ( .A1(n5217), .A2(n6565), .B1(INSTQUEUE_REG_12__4__SCAN_IN), 
        .B2(n5216), .ZN(n5192) );
  OAI21_X1 U6309 ( .B1(n5193), .B2(n5219), .A(n5192), .ZN(n5194) );
  AOI21_X1 U6310 ( .B1(n6460), .B2(n5222), .A(n5194), .ZN(n5195) );
  OAI21_X1 U6311 ( .B1(n6463), .B2(n6592), .A(n5195), .ZN(U3120) );
  AOI22_X1 U6312 ( .A1(n5217), .A2(n6588), .B1(INSTQUEUE_REG_12__7__SCAN_IN), 
        .B2(n5216), .ZN(n5196) );
  OAI21_X1 U6313 ( .B1(n5197), .B2(n5219), .A(n5196), .ZN(n5198) );
  AOI21_X1 U6314 ( .B1(n6516), .B2(n5222), .A(n5198), .ZN(n5199) );
  OAI21_X1 U6315 ( .B1(n6524), .B2(n6592), .A(n5199), .ZN(U3123) );
  AOI22_X1 U6316 ( .A1(n5217), .A2(n6541), .B1(INSTQUEUE_REG_12__0__SCAN_IN), 
        .B2(n5216), .ZN(n5200) );
  OAI21_X1 U6317 ( .B1(n5201), .B2(n5219), .A(n5200), .ZN(n5202) );
  AOI21_X1 U6318 ( .B1(n6482), .B2(n5222), .A(n5202), .ZN(n5203) );
  OAI21_X1 U6319 ( .B1(n6495), .B2(n6592), .A(n5203), .ZN(U3116) );
  AOI22_X1 U6320 ( .A1(n5217), .A2(n6547), .B1(INSTQUEUE_REG_12__1__SCAN_IN), 
        .B2(n5216), .ZN(n5204) );
  OAI21_X1 U6321 ( .B1(n5205), .B2(n5219), .A(n5204), .ZN(n5206) );
  AOI21_X1 U6322 ( .B1(n6546), .B2(n5222), .A(n5206), .ZN(n5207) );
  OAI21_X1 U6323 ( .B1(n6550), .B2(n6592), .A(n5207), .ZN(U3117) );
  AOI22_X1 U6324 ( .A1(n5217), .A2(n6571), .B1(INSTQUEUE_REG_12__5__SCAN_IN), 
        .B2(n5216), .ZN(n5208) );
  OAI21_X1 U6325 ( .B1(n5209), .B2(n5219), .A(n5208), .ZN(n5210) );
  AOI21_X1 U6326 ( .B1(n6506), .B2(n5222), .A(n5210), .ZN(n5211) );
  OAI21_X1 U6327 ( .B1(n6509), .B2(n6592), .A(n5211), .ZN(U3121) );
  AOI22_X1 U6328 ( .A1(n5217), .A2(n6578), .B1(INSTQUEUE_REG_12__6__SCAN_IN), 
        .B2(n5216), .ZN(n5212) );
  OAI21_X1 U6329 ( .B1(n5213), .B2(n5219), .A(n5212), .ZN(n5214) );
  AOI21_X1 U6330 ( .B1(n6576), .B2(n5222), .A(n5214), .ZN(n5215) );
  OAI21_X1 U6331 ( .B1(n6582), .B2(n6592), .A(n5215), .ZN(U3122) );
  AOI22_X1 U6332 ( .A1(n5217), .A2(n6553), .B1(INSTQUEUE_REG_12__2__SCAN_IN), 
        .B2(n5216), .ZN(n5218) );
  OAI21_X1 U6333 ( .B1(n5220), .B2(n5219), .A(n5218), .ZN(n5221) );
  AOI21_X1 U6334 ( .B1(n6452), .B2(n5222), .A(n5221), .ZN(n5223) );
  OAI21_X1 U6335 ( .B1(n6455), .B2(n6592), .A(n5223), .ZN(U3118) );
  OAI22_X1 U6336 ( .A1(n6205), .A2(n5236), .B1(n6960), .B2(n6172), .ZN(n5224)
         );
  AOI21_X1 U6337 ( .B1(REIP_REG_0__SCAN_IN), .B2(n6132), .A(n5224), .ZN(n5227)
         );
  NAND2_X1 U6338 ( .A1(n6171), .A2(n6188), .ZN(n5225) );
  AOI22_X1 U6339 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n5225), .B1(n6196), 
        .B2(n6597), .ZN(n5226) );
  OAI211_X1 U6340 ( .C1(n6193), .C2(n5959), .A(n5227), .B(n5226), .ZN(U2827)
         );
  AND2_X1 U6341 ( .A1(n4996), .A2(n5228), .ZN(n5230) );
  OR2_X1 U6342 ( .A1(n5230), .A2(n5229), .ZN(n6274) );
  AOI22_X1 U6343 ( .A1(n6236), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6230), .ZN(n5231) );
  OAI21_X1 U6344 ( .B1(n6274), .B2(n5697), .A(n5231), .ZN(U2880) );
  AOI22_X1 U6345 ( .A1(n6236), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6230), .ZN(n5232) );
  OAI21_X1 U6346 ( .B1(n5316), .B2(n5697), .A(n5232), .ZN(U2883) );
  OAI222_X1 U6347 ( .A1(n5233), .A2(n5697), .B1(n5235), .B2(n7004), .C1(n6240), 
        .C2(n6265), .ZN(U2890) );
  OAI222_X1 U6348 ( .A1(n6178), .A2(n5697), .B1(n5235), .B2(n6868), .C1(n6240), 
        .C2(n6256), .ZN(U2885) );
  OAI222_X1 U6349 ( .A1(n5236), .A2(n5697), .B1(n5235), .B2(n5234), .C1(n6240), 
        .C2(n6988), .ZN(U2891) );
  INV_X1 U6350 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5245) );
  NOR2_X1 U6351 ( .A1(n6161), .A2(n5237), .ZN(n5244) );
  NAND2_X1 U6352 ( .A1(n5495), .A2(n5245), .ZN(n5240) );
  NAND2_X1 U6353 ( .A1(n5605), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5238) );
  OAI211_X1 U6354 ( .C1(EBX_REG_11__SCAN_IN), .C2(n4434), .A(n5238), .B(n5153), 
        .ZN(n5239) );
  AND2_X1 U6355 ( .A1(n5240), .A2(n5239), .ZN(n5243) );
  NAND2_X1 U6356 ( .A1(n5241), .A2(n5243), .ZN(n5242) );
  OAI21_X1 U6357 ( .B1(n5244), .B2(n5243), .A(n5370), .ZN(n6309) );
  OAI222_X1 U6358 ( .A1(n6274), .A2(n5680), .B1(n6221), .B2(n5245), .C1(n5678), 
        .C2(n6309), .ZN(U2848) );
  INV_X1 U6359 ( .A(n5246), .ZN(n6336) );
  AOI22_X1 U6360 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6198), .B1(n6202), .B2(n6336), 
        .ZN(n5247) );
  OAI211_X1 U6361 ( .C1(n6171), .C2(n5248), .A(n5247), .B(n6186), .ZN(n5254)
         );
  OR2_X1 U6362 ( .A1(n5249), .A2(n6187), .ZN(n5305) );
  NOR2_X1 U6363 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5305), .ZN(n6179) );
  OAI21_X1 U6364 ( .B1(n6176), .B2(n6179), .A(REIP_REG_7__SCAN_IN), .ZN(n5251)
         );
  INV_X1 U6365 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6673) );
  OR3_X1 U6366 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6673), .A3(n5305), .ZN(n5250)
         );
  OAI211_X1 U6367 ( .C1(n6188), .C2(n5252), .A(n5251), .B(n5250), .ZN(n5253)
         );
  AOI211_X1 U6368 ( .C1(n5255), .C2(n6167), .A(n5254), .B(n5253), .ZN(n5256)
         );
  INV_X1 U6369 ( .A(n5256), .ZN(U2820) );
  NAND2_X1 U6370 ( .A1(n6528), .A2(n6405), .ZN(n6581) );
  OAI21_X1 U6371 ( .B1(n5297), .B2(n6586), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5257) );
  NAND2_X1 U6372 ( .A1(n5257), .A2(n6530), .ZN(n5264) );
  NAND2_X1 U6373 ( .A1(n3262), .A2(n3172), .ZN(n5262) );
  NAND2_X1 U6374 ( .A1(n5259), .A2(n5258), .ZN(n6408) );
  OAI22_X1 U6375 ( .A1(n5264), .A2(n5262), .B1(n6435), .B2(n6408), .ZN(n5301)
         );
  NAND3_X1 U6376 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6607), .ZN(n6538) );
  NOR2_X1 U6377 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6538), .ZN(n5296)
         );
  NOR2_X1 U6378 ( .A1(n5261), .A2(n5260), .ZN(n6411) );
  INV_X1 U6379 ( .A(n5262), .ZN(n6533) );
  OAI22_X1 U6380 ( .A1(n5264), .A2(n6533), .B1(n5296), .B2(n5263), .ZN(n5265)
         );
  INV_X1 U6381 ( .A(n5265), .ZN(n5266) );
  OAI211_X1 U6382 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6737), .A(n6411), .B(n5266), .ZN(n5295) );
  AOI22_X1 U6383 ( .A1(n6557), .A2(n5296), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5295), .ZN(n5268) );
  NAND2_X1 U6384 ( .A1(n5297), .A2(n6558), .ZN(n5267) );
  OAI211_X1 U6385 ( .C1(n6581), .C2(n6562), .A(n5268), .B(n5267), .ZN(n5269)
         );
  AOI21_X1 U6386 ( .B1(n5301), .B2(n6559), .A(n5269), .ZN(n5270) );
  INV_X1 U6387 ( .A(n5270), .ZN(U3103) );
  AOI22_X1 U6388 ( .A1(n6584), .A2(n5296), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5295), .ZN(n5272) );
  NAND2_X1 U6389 ( .A1(n5297), .A2(n6585), .ZN(n5271) );
  OAI211_X1 U6390 ( .C1(n6581), .C2(n6593), .A(n5272), .B(n5271), .ZN(n5273)
         );
  AOI21_X1 U6391 ( .B1(n5301), .B2(n6588), .A(n5273), .ZN(n5274) );
  INV_X1 U6392 ( .A(n5274), .ZN(U3107) );
  AOI22_X1 U6393 ( .A1(n6526), .A2(n5296), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5295), .ZN(n5276) );
  NAND2_X1 U6394 ( .A1(n5297), .A2(n6527), .ZN(n5275) );
  OAI211_X1 U6395 ( .C1(n6581), .C2(n6544), .A(n5276), .B(n5275), .ZN(n5277)
         );
  AOI21_X1 U6396 ( .B1(n5301), .B2(n6541), .A(n5277), .ZN(n5278) );
  INV_X1 U6397 ( .A(n5278), .ZN(U3100) );
  AOI22_X1 U6398 ( .A1(n6563), .A2(n5296), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5295), .ZN(n5280) );
  NAND2_X1 U6399 ( .A1(n5297), .A2(n6564), .ZN(n5279) );
  OAI211_X1 U6400 ( .C1(n6581), .C2(n6568), .A(n5280), .B(n5279), .ZN(n5281)
         );
  AOI21_X1 U6401 ( .B1(n5301), .B2(n6565), .A(n5281), .ZN(n5282) );
  INV_X1 U6402 ( .A(n5282), .ZN(U3104) );
  AOI22_X1 U6403 ( .A1(n6545), .A2(n5296), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5295), .ZN(n5284) );
  NAND2_X1 U6404 ( .A1(n5297), .A2(n6415), .ZN(n5283) );
  OAI211_X1 U6405 ( .C1(n6581), .C2(n6418), .A(n5284), .B(n5283), .ZN(n5285)
         );
  AOI21_X1 U6406 ( .B1(n5301), .B2(n6547), .A(n5285), .ZN(n5286) );
  INV_X1 U6407 ( .A(n5286), .ZN(U3101) );
  AOI22_X1 U6408 ( .A1(n6551), .A2(n5296), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5295), .ZN(n5288) );
  NAND2_X1 U6409 ( .A1(n5297), .A2(n6552), .ZN(n5287) );
  OAI211_X1 U6410 ( .C1(n6581), .C2(n6556), .A(n5288), .B(n5287), .ZN(n5289)
         );
  AOI21_X1 U6411 ( .B1(n5301), .B2(n6553), .A(n5289), .ZN(n5290) );
  INV_X1 U6412 ( .A(n5290), .ZN(U3102) );
  AOI22_X1 U6413 ( .A1(n6575), .A2(n5296), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5295), .ZN(n5292) );
  NAND2_X1 U6414 ( .A1(n5297), .A2(n6510), .ZN(n5291) );
  OAI211_X1 U6415 ( .C1(n6581), .C2(n6515), .A(n5292), .B(n5291), .ZN(n5293)
         );
  AOI21_X1 U6416 ( .B1(n5301), .B2(n6578), .A(n5293), .ZN(n5294) );
  INV_X1 U6417 ( .A(n5294), .ZN(U3106) );
  AOI22_X1 U6418 ( .A1(n6569), .A2(n5296), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5295), .ZN(n5299) );
  NAND2_X1 U6419 ( .A1(n5297), .A2(n6570), .ZN(n5298) );
  OAI211_X1 U6420 ( .C1(n6581), .C2(n6574), .A(n5299), .B(n5298), .ZN(n5300)
         );
  AOI21_X1 U6421 ( .B1(n5301), .B2(n6571), .A(n5300), .ZN(n5302) );
  INV_X1 U6422 ( .A(n5302), .ZN(U3105) );
  INV_X1 U6423 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6993) );
  NOR2_X1 U6424 ( .A1(n6993), .A2(n6673), .ZN(n5306) );
  INV_X1 U6425 ( .A(n5306), .ZN(n5304) );
  OAI21_X1 U6426 ( .B1(n5305), .B2(n5304), .A(n5303), .ZN(n5314) );
  NAND4_X1 U6427 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5308), .A3(n5307), .A4(n5306), .ZN(n5325) );
  INV_X1 U6428 ( .A(n5325), .ZN(n5318) );
  OAI21_X1 U6429 ( .B1(n5516), .B2(n5318), .A(n5326), .ZN(n6162) );
  NOR2_X1 U6430 ( .A1(n6188), .A2(n5309), .ZN(n5313) );
  AOI22_X1 U6431 ( .A1(EBX_REG_8__SCAN_IN), .A2(n6198), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n6197), .ZN(n5310) );
  OAI211_X1 U6432 ( .C1(n6193), .C2(n5311), .A(n5310), .B(n6186), .ZN(n5312)
         );
  AOI211_X1 U6433 ( .C1(n5314), .C2(n6162), .A(n5313), .B(n5312), .ZN(n5315)
         );
  OAI21_X1 U6434 ( .B1(n6177), .B2(n5316), .A(n5315), .ZN(U2819) );
  OAI22_X1 U6435 ( .A1(n6193), .A2(n6317), .B1(n5317), .B2(n6188), .ZN(n5322)
         );
  NAND2_X1 U6436 ( .A1(n5418), .A2(n5318), .ZN(n6163) );
  NAND2_X1 U6437 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5327) );
  OAI21_X1 U6438 ( .B1(REIP_REG_10__SCAN_IN), .B2(REIP_REG_9__SCAN_IN), .A(
        n5327), .ZN(n5320) );
  AOI22_X1 U6439 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6198), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n6197), .ZN(n5319) );
  OAI211_X1 U6440 ( .C1(n6163), .C2(n5320), .A(n5319), .B(n6186), .ZN(n5321)
         );
  AOI211_X1 U6441 ( .C1(REIP_REG_10__SCAN_IN), .C2(n6162), .A(n5322), .B(n5321), .ZN(n5323) );
  OAI21_X1 U6442 ( .B1(n5324), .B2(n6177), .A(n5323), .ZN(U2817) );
  INV_X1 U6443 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6679) );
  NOR3_X1 U6444 ( .A1(n6679), .A2(n5325), .A3(n5327), .ZN(n5417) );
  AND2_X1 U6445 ( .A1(n5326), .A2(n5417), .ZN(n5420) );
  NOR2_X1 U6446 ( .A1(n6185), .A2(n5420), .ZN(n6149) );
  OAI21_X1 U6447 ( .B1(n5327), .B2(n6163), .A(n6679), .ZN(n5332) );
  NOR2_X1 U6448 ( .A1(n6193), .A2(n6309), .ZN(n5331) );
  AOI22_X1 U6449 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6198), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n6197), .ZN(n5328) );
  OAI211_X1 U6450 ( .C1(n6188), .C2(n5329), .A(n5328), .B(n6186), .ZN(n5330)
         );
  AOI211_X1 U6451 ( .C1(n6149), .C2(n5332), .A(n5331), .B(n5330), .ZN(n5333)
         );
  OAI21_X1 U6452 ( .B1(n6274), .B2(n6177), .A(n5333), .ZN(U2816) );
  XOR2_X1 U6453 ( .A(n5229), .B(n5334), .Z(n6238) );
  INV_X1 U6454 ( .A(n6238), .ZN(n5339) );
  MUX2_X1 U6455 ( .A(n5502), .B(n5153), .S(EBX_REG_12__SCAN_IN), .Z(n5337) );
  NAND2_X1 U6456 ( .A1(n4434), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5335) );
  AND2_X1 U6457 ( .A1(n5464), .A2(n5335), .ZN(n5336) );
  NAND2_X1 U6458 ( .A1(n5337), .A2(n5336), .ZN(n5368) );
  XNOR2_X1 U6459 ( .A(n5370), .B(n5368), .ZN(n6150) );
  AOI22_X1 U6460 ( .A1(n6150), .A2(n6217), .B1(EBX_REG_12__SCAN_IN), .B2(n5634), .ZN(n5338) );
  OAI21_X1 U6461 ( .B1(n5339), .B2(n5680), .A(n5338), .ZN(U2847) );
  XOR2_X1 U6462 ( .A(n5342), .B(n5341), .Z(n5355) );
  INV_X1 U6463 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6902) );
  NAND3_X1 U6464 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6320), .ZN(n5345) );
  NOR2_X1 U6465 ( .A1(n5345), .A2(n5344), .ZN(n5805) );
  NAND2_X1 U6466 ( .A1(n5805), .A2(n6399), .ZN(n5348) );
  INV_X1 U6467 ( .A(n5348), .ZN(n5940) );
  NAND3_X1 U6468 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6885), .A3(n6311), .ZN(n5346) );
  OAI21_X1 U6469 ( .B1(n6388), .B2(n6902), .A(n5346), .ZN(n5347) );
  AOI21_X1 U6470 ( .B1(n6383), .B2(n6150), .A(n5347), .ZN(n5351) );
  INV_X1 U6471 ( .A(n5804), .ZN(n5917) );
  OAI22_X1 U6472 ( .A1(n5917), .A2(n5803), .B1(n6348), .B2(n5805), .ZN(n6312)
         );
  AOI21_X1 U6473 ( .B1(n5814), .B2(n5348), .A(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n5349) );
  OAI21_X1 U6474 ( .B1(n6312), .B2(n5349), .A(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n5350) );
  OAI211_X1 U6475 ( .C1(n5355), .C2(n6370), .A(n5351), .B(n5350), .ZN(U3006)
         );
  AOI22_X1 U6476 ( .A1(n6299), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6353), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5352) );
  OAI21_X1 U6477 ( .B1(n6152), .B2(n6308), .A(n5352), .ZN(n5353) );
  AOI21_X1 U6478 ( .B1(n6238), .B2(n4244), .A(n5353), .ZN(n5354) );
  OAI21_X1 U6479 ( .B1(n5355), .B2(n6294), .A(n5354), .ZN(U2974) );
  NOR2_X1 U6480 ( .A1(n3700), .A2(n6885), .ZN(n5356) );
  INV_X1 U6481 ( .A(n5356), .ZN(n5362) );
  NOR2_X1 U6482 ( .A1(n5375), .A2(n5362), .ZN(n5802) );
  OAI22_X1 U6483 ( .A1(n5802), .A2(n5962), .B1(n5357), .B2(n5356), .ZN(n5358)
         );
  NOR2_X1 U6484 ( .A1(n6312), .A2(n5358), .ZN(n5391) );
  OAI21_X1 U6485 ( .B1(n5361), .B2(n5360), .A(n5359), .ZN(n6060) );
  NAND2_X1 U6486 ( .A1(n6060), .A2(n6396), .ZN(n5374) );
  NOR2_X1 U6487 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5362), .ZN(n5388)
         );
  INV_X1 U6488 ( .A(n5370), .ZN(n5366) );
  INV_X1 U6489 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6490 ( .A1(n5495), .A2(n5382), .ZN(n5365) );
  NAND2_X1 U6491 ( .A1(n5605), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5363) );
  OAI211_X1 U6492 ( .C1(n4434), .C2(EBX_REG_13__SCAN_IN), .A(n5363), .B(n5153), 
        .ZN(n5364) );
  AND2_X1 U6493 ( .A1(n5365), .A2(n5364), .ZN(n5367) );
  AOI21_X1 U6494 ( .B1(n5366), .B2(n5368), .A(n5367), .ZN(n5371) );
  NAND2_X1 U6495 ( .A1(n5368), .A2(n5367), .ZN(n5369) );
  OR2_X1 U6496 ( .A1(n5371), .A2(n5408), .ZN(n6143) );
  NAND2_X1 U6497 ( .A1(n6353), .A2(REIP_REG_13__SCAN_IN), .ZN(n6061) );
  OAI21_X1 U6498 ( .B1(n6390), .B2(n6143), .A(n6061), .ZN(n5372) );
  AOI21_X1 U6499 ( .B1(n6311), .B2(n5388), .A(n5372), .ZN(n5373) );
  OAI211_X1 U6500 ( .C1(n5391), .C2(n5375), .A(n5374), .B(n5373), .ZN(U3005)
         );
  NAND2_X1 U6501 ( .A1(n5376), .A2(n5377), .ZN(n5378) );
  AND2_X1 U6502 ( .A1(n5379), .A2(n5378), .ZN(n6145) );
  INV_X1 U6503 ( .A(n6145), .ZN(n5381) );
  AOI22_X1 U6504 ( .A1(n6236), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n6230), .ZN(n5380) );
  OAI21_X1 U6505 ( .B1(n5381), .B2(n5697), .A(n5380), .ZN(U2878) );
  OAI22_X1 U6506 ( .A1(n6143), .A2(n5678), .B1(n5382), .B2(n6221), .ZN(n5383)
         );
  AOI21_X1 U6507 ( .B1(n6145), .B2(n6218), .A(n5383), .ZN(n5384) );
  INV_X1 U6508 ( .A(n5384), .ZN(U2846) );
  XNOR2_X1 U6509 ( .A(n6271), .B(n5392), .ZN(n5386) );
  XNOR2_X1 U6510 ( .A(n5387), .B(n5386), .ZN(n5435) );
  OAI21_X1 U6511 ( .B1(n5389), .B2(n5803), .A(n5388), .ZN(n5390) );
  AOI21_X1 U6512 ( .B1(n5391), .B2(n5390), .A(n5392), .ZN(n5400) );
  INV_X1 U6513 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6684) );
  NAND3_X1 U6514 ( .A1(n5802), .A2(n5392), .A3(n6311), .ZN(n5398) );
  MUX2_X1 U6515 ( .A(n5502), .B(n5153), .S(EBX_REG_14__SCAN_IN), .Z(n5395) );
  NAND2_X1 U6516 ( .A1(n4434), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5393) );
  AND2_X1 U6517 ( .A1(n5464), .A2(n5393), .ZN(n5394) );
  NAND2_X1 U6518 ( .A1(n5395), .A2(n5394), .ZN(n5407) );
  INV_X1 U6519 ( .A(n5407), .ZN(n5396) );
  XNOR2_X1 U6520 ( .A(n5408), .B(n5396), .ZN(n6215) );
  NAND2_X1 U6521 ( .A1(n6383), .A2(n6215), .ZN(n5397) );
  OAI211_X1 U6522 ( .C1(n6684), .C2(n6388), .A(n5398), .B(n5397), .ZN(n5399)
         );
  NOR2_X1 U6523 ( .A1(n5400), .A2(n5399), .ZN(n5401) );
  OAI21_X1 U6524 ( .B1(n5435), .B2(n6370), .A(n5401), .ZN(U3004) );
  INV_X1 U6525 ( .A(n5403), .ZN(n5405) );
  NAND2_X1 U6526 ( .A1(n5405), .A2(n3232), .ZN(n5406) );
  AND2_X1 U6527 ( .A1(n5402), .A2(n5406), .ZN(n5800) );
  INV_X1 U6528 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6529 ( .A1(n5495), .A2(n5425), .ZN(n5411) );
  NAND2_X1 U6530 ( .A1(n5605), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5409) );
  OAI211_X1 U6531 ( .C1(n4434), .C2(EBX_REG_15__SCAN_IN), .A(n5409), .B(n5153), 
        .ZN(n5410) );
  NAND2_X1 U6532 ( .A1(n5411), .A2(n5410), .ZN(n5412) );
  NAND2_X1 U6533 ( .A1(n5413), .A2(n5412), .ZN(n5414) );
  NAND2_X1 U6534 ( .A1(n5676), .A2(n5414), .ZN(n5952) );
  AOI22_X1 U6535 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6198), .B1(
        PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n6197), .ZN(n5415) );
  OAI211_X1 U6536 ( .C1(n5952), .C2(n6193), .A(n5415), .B(n6186), .ZN(n5416)
         );
  INV_X1 U6537 ( .A(n5416), .ZN(n5422) );
  NAND3_X1 U6538 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_14__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .ZN(n5419) );
  NOR2_X1 U6539 ( .A1(n6139), .A2(n5419), .ZN(n5508) );
  INV_X1 U6540 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6686) );
  NAND4_X1 U6541 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_14__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .A4(n5420), .ZN(n6133) );
  NOR2_X1 U6542 ( .A1(n6686), .A2(n6133), .ZN(n5512) );
  NOR2_X1 U6543 ( .A1(n6185), .A2(n5512), .ZN(n6123) );
  OAI21_X1 U6544 ( .B1(REIP_REG_15__SCAN_IN), .B2(n5508), .A(n6123), .ZN(n5421) );
  OAI211_X1 U6545 ( .C1(n6188), .C2(n5798), .A(n5422), .B(n5421), .ZN(n5423)
         );
  AOI21_X1 U6546 ( .B1(n5800), .B2(n6167), .A(n5423), .ZN(n5424) );
  INV_X1 U6547 ( .A(n5424), .ZN(U2812) );
  OAI22_X1 U6548 ( .A1(n5952), .A2(n5678), .B1(n5425), .B2(n6221), .ZN(n5426)
         );
  AOI21_X1 U6549 ( .B1(n5800), .B2(n6218), .A(n5426), .ZN(n5427) );
  INV_X1 U6550 ( .A(n5427), .ZN(U2844) );
  NOR2_X1 U6551 ( .A1(n5428), .A2(n5429), .ZN(n5430) );
  NOR2_X1 U6552 ( .A1(n5403), .A2(n5430), .ZN(n6234) );
  INV_X1 U6553 ( .A(n6131), .ZN(n5432) );
  AOI22_X1 U6554 ( .A1(n6299), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6353), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5431) );
  OAI21_X1 U6555 ( .B1(n6308), .B2(n5432), .A(n5431), .ZN(n5433) );
  AOI21_X1 U6556 ( .B1(n6234), .B2(n4244), .A(n5433), .ZN(n5434) );
  OAI21_X1 U6557 ( .B1(n5435), .B2(n6294), .A(n5434), .ZN(U2972) );
  INV_X1 U6558 ( .A(n5800), .ZN(n5437) );
  AOI22_X1 U6559 ( .A1(n6236), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6230), .ZN(n5436) );
  OAI21_X1 U6560 ( .B1(n5437), .B2(n5697), .A(n5436), .ZN(U2876) );
  OAI22_X1 U6561 ( .A1(n5438), .A2(n6638), .B1(n6645), .B2(n6090), .ZN(n6084)
         );
  NOR2_X1 U6562 ( .A1(n6084), .A2(n6718), .ZN(n6080) );
  INV_X1 U6563 ( .A(n6596), .ZN(n5442) );
  NOR3_X1 U6564 ( .A1(n6594), .A2(n4581), .A3(n4530), .ZN(n5439) );
  AOI21_X1 U6565 ( .B1(n6598), .B2(n5440), .A(n5439), .ZN(n5441) );
  OAI21_X1 U6566 ( .B1(n5969), .B2(n5442), .A(n5441), .ZN(n6599) );
  INV_X1 U6567 ( .A(n6727), .ZN(n6082) );
  INV_X1 U6568 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5443) );
  AOI22_X1 U6569 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5443), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6852), .ZN(n5450) );
  INV_X1 U6570 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5451) );
  NOR2_X1 U6571 ( .A1(n5452), .A2(n5451), .ZN(n5445) );
  AOI222_X1 U6572 ( .A1(n6599), .A2(n6082), .B1(n5450), .B2(n5445), .C1(n5444), 
        .C2(n5448), .ZN(n5447) );
  NOR2_X1 U6573 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6629), .ZN(n6721)
         );
  OAI21_X1 U6574 ( .B1(n6080), .B2(n6721), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n5446) );
  OAI21_X1 U6575 ( .B1(n6080), .B2(n5447), .A(n5446), .ZN(U3460) );
  AOI21_X1 U6576 ( .B1(n5448), .B2(n5453), .A(n6080), .ZN(n5458) );
  INV_X1 U6577 ( .A(n5449), .ZN(n5456) );
  NOR3_X1 U6578 ( .A1(n5452), .A2(n5451), .A3(n5450), .ZN(n5455) );
  NOR3_X1 U6579 ( .A1(n5453), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6629), 
        .ZN(n5454) );
  AOI211_X1 U6580 ( .C1(n5456), .C2(n6082), .A(n5455), .B(n5454), .ZN(n5457)
         );
  OAI22_X1 U6581 ( .A1(n5458), .A2(n4558), .B1(n6080), .B2(n5457), .ZN(U3459)
         );
  NAND2_X1 U6582 ( .A1(n6240), .A2(n5460), .ZN(n5462) );
  AOI22_X1 U6583 ( .A1(n6228), .A2(DATAI_31_), .B1(n6230), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5461) );
  OAI21_X1 U6584 ( .B1(n5459), .B2(n5462), .A(n5461), .ZN(U2860) );
  OAI22_X1 U6585 ( .A1(n5503), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4434), .ZN(n5507) );
  MUX2_X1 U6586 ( .A(n5502), .B(n5153), .S(EBX_REG_16__SCAN_IN), .Z(n5466) );
  NAND2_X1 U6587 ( .A1(n4434), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5463) );
  AND2_X1 U6588 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  AND2_X1 U6589 ( .A1(n5466), .A2(n5465), .ZN(n5675) );
  INV_X1 U6590 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U6591 ( .A1(n5495), .A2(n6214), .ZN(n5469) );
  NAND2_X1 U6592 ( .A1(n5605), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5467) );
  OAI211_X1 U6593 ( .C1(n4434), .C2(EBX_REG_17__SCAN_IN), .A(n5467), .B(n5153), 
        .ZN(n5468) );
  MUX2_X1 U6594 ( .A(n5502), .B(n5153), .S(EBX_REG_19__SCAN_IN), .Z(n5471) );
  NAND2_X1 U6595 ( .A1(n4434), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6596 ( .A1(n5471), .A2(n5470), .ZN(n5665) );
  NAND2_X1 U6597 ( .A1(n5497), .A2(n5943), .ZN(n5474) );
  INV_X1 U6598 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6599 ( .A1(n5473), .A2(n5472), .ZN(n5661) );
  AND2_X1 U6600 ( .A1(n5474), .A2(n5661), .ZN(n5664) );
  OAI22_X1 U6601 ( .A1(n5503), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n4434), .ZN(n5607) );
  NAND2_X1 U6602 ( .A1(n5664), .A2(n5607), .ZN(n5476) );
  NAND2_X1 U6603 ( .A1(n5662), .A2(EBX_REG_20__SCAN_IN), .ZN(n5475) );
  OAI211_X1 U6604 ( .C1(n5664), .C2(n5662), .A(n5476), .B(n5475), .ZN(n5477)
         );
  MUX2_X1 U6605 ( .A(n5495), .B(n5662), .S(EBX_REG_21__SCAN_IN), .Z(n5478) );
  INV_X1 U6606 ( .A(n5478), .ZN(n5480) );
  INV_X1 U6607 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U6608 ( .A1(n5497), .A2(n5913), .ZN(n5479) );
  NAND2_X1 U6609 ( .A1(n5480), .A2(n5479), .ZN(n5650) );
  INV_X1 U6610 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6888) );
  NAND2_X1 U6611 ( .A1(n5495), .A2(n6888), .ZN(n5483) );
  NAND2_X1 U6612 ( .A1(n5605), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5481) );
  OAI211_X1 U6613 ( .C1(n4434), .C2(EBX_REG_23__SCAN_IN), .A(n5481), .B(n5153), 
        .ZN(n5482) );
  AND2_X1 U6614 ( .A1(n5483), .A2(n5482), .ZN(n5639) );
  INV_X1 U6615 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U6616 ( .A1(n5484), .A2(n5645), .ZN(n5487) );
  INV_X1 U6617 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6985) );
  NAND2_X1 U6618 ( .A1(n5153), .A2(n6985), .ZN(n5485) );
  OAI211_X1 U6619 ( .C1(n4434), .C2(EBX_REG_22__SCAN_IN), .A(n5485), .B(n5605), 
        .ZN(n5486) );
  NAND2_X1 U6620 ( .A1(n5487), .A2(n5486), .ZN(n5640) );
  MUX2_X1 U6621 ( .A(n5502), .B(n5153), .S(EBX_REG_24__SCAN_IN), .Z(n5489) );
  NAND2_X1 U6622 ( .A1(n4434), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U6623 ( .A1(n5489), .A2(n5488), .ZN(n5633) );
  MUX2_X1 U6624 ( .A(n5495), .B(n5662), .S(EBX_REG_25__SCAN_IN), .Z(n5491) );
  NOR2_X1 U6625 ( .A1(n5503), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5490)
         );
  NOR2_X1 U6626 ( .A1(n5491), .A2(n5490), .ZN(n5624) );
  AND2_X1 U6627 ( .A1(n5633), .A2(n5624), .ZN(n5492) );
  MUX2_X1 U6628 ( .A(n5502), .B(n5153), .S(EBX_REG_26__SCAN_IN), .Z(n5494) );
  NAND2_X1 U6629 ( .A1(n4434), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5493) );
  AND2_X1 U6630 ( .A1(n5494), .A2(n5493), .ZN(n5621) );
  MUX2_X1 U6631 ( .A(n5495), .B(n5662), .S(EBX_REG_27__SCAN_IN), .Z(n5496) );
  INV_X1 U6632 ( .A(n5496), .ZN(n5499) );
  NAND2_X1 U6633 ( .A1(n5497), .A2(n5710), .ZN(n5498) );
  NAND2_X1 U6634 ( .A1(n5499), .A2(n5498), .ZN(n5573) );
  NAND2_X1 U6635 ( .A1(n5153), .A2(n5708), .ZN(n5500) );
  OAI211_X1 U6636 ( .C1(n4434), .C2(EBX_REG_28__SCAN_IN), .A(n5500), .B(n5605), 
        .ZN(n5501) );
  OAI21_X1 U6637 ( .B1(n5502), .B2(EBX_REG_28__SCAN_IN), .A(n5501), .ZN(n5559)
         );
  OAI22_X1 U6638 ( .A1(n5503), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n4434), .ZN(n5545) );
  INV_X1 U6639 ( .A(n5549), .ZN(n5560) );
  NOR2_X1 U6640 ( .A1(n5502), .A2(EBX_REG_29__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U6641 ( .A1(n5503), .A2(EBX_REG_30__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U6642 ( .A1(n4434), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U6643 ( .A1(n5505), .A2(n5504), .ZN(n5533) );
  NAND2_X1 U6644 ( .A1(n5536), .A2(n5605), .ZN(n5532) );
  OAI21_X1 U6645 ( .B1(n5551), .B2(n5533), .A(n5532), .ZN(n5506) );
  XOR2_X1 U6646 ( .A(n5507), .B(n5506), .Z(n5830) );
  NAND2_X1 U6647 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5508), .ZN(n6125) );
  NAND2_X1 U6648 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .ZN(
        n5509) );
  NOR2_X1 U6649 ( .A1(n6125), .A2(n5509), .ZN(n6019) );
  NAND2_X1 U6650 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6019), .ZN(n6020) );
  NAND2_X1 U6651 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n5513) );
  NOR2_X1 U6652 ( .A1(n6020), .A2(n5513), .ZN(n5591) );
  NAND2_X1 U6653 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5591), .ZN(n6001) );
  NAND2_X1 U6654 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .ZN(
        n5510) );
  NAND3_X1 U6655 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5579) );
  INV_X1 U6656 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5583) );
  NOR2_X1 U6657 ( .A1(n5579), .A2(n5583), .ZN(n5511) );
  NAND2_X1 U6658 ( .A1(n5987), .A2(n5511), .ZN(n5566) );
  INV_X1 U6659 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6704) );
  INV_X1 U6660 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6705) );
  INV_X1 U6661 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6708) );
  NOR3_X1 U6662 ( .A1(n5544), .A2(REIP_REG_31__SCAN_IN), .A3(n6708), .ZN(n5524) );
  INV_X1 U6663 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6690) );
  NAND3_X1 U6664 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        n5512), .ZN(n6018) );
  NOR3_X1 U6665 ( .A1(n6690), .A2(n5513), .A3(n6018), .ZN(n5590) );
  NAND4_X1 U6666 ( .A1(n5590), .A2(REIP_REG_23__SCAN_IN), .A3(
        REIP_REG_22__SCAN_IN), .A4(REIP_REG_21__SCAN_IN), .ZN(n5986) );
  OR2_X1 U6667 ( .A1(n5986), .A2(n5579), .ZN(n5514) );
  NAND2_X1 U6668 ( .A1(n5514), .A2(n6132), .ZN(n5976) );
  NAND2_X1 U6669 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5976), .ZN(n5515) );
  OAI21_X1 U6670 ( .B1(n5515), .B2(n6705), .A(n6132), .ZN(n5565) );
  OAI21_X1 U6671 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5516), .A(n5565), .ZN(n5541) );
  NOR2_X1 U6672 ( .A1(n5516), .A2(REIP_REG_30__SCAN_IN), .ZN(n5517) );
  OAI21_X1 U6673 ( .B1(n5541), .B2(n5517), .A(REIP_REG_31__SCAN_IN), .ZN(n5522) );
  INV_X1 U6674 ( .A(n5518), .ZN(n5520) );
  NAND3_X1 U6675 ( .A1(n5520), .A2(EBX_REG_31__SCAN_IN), .A3(n5519), .ZN(n5521) );
  OAI211_X1 U6676 ( .C1(n6832), .C2(n6171), .A(n5522), .B(n5521), .ZN(n5523)
         );
  AOI211_X1 U6677 ( .C1(n5830), .C2(n6202), .A(n5524), .B(n5523), .ZN(n5525)
         );
  OAI21_X1 U6678 ( .B1(n5459), .B2(n6177), .A(n5525), .ZN(U2796) );
  NAND2_X1 U6679 ( .A1(n5705), .A2(n6167), .ZN(n5543) );
  INV_X1 U6680 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6843) );
  INV_X1 U6681 ( .A(n5703), .ZN(n5529) );
  AOI22_X1 U6682 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6197), .B1(n6207), 
        .B2(n5529), .ZN(n5530) );
  OAI21_X1 U6683 ( .B1(n6843), .B2(n6172), .A(n5530), .ZN(n5540) );
  NAND2_X1 U6684 ( .A1(n5536), .A2(n5560), .ZN(n5531) );
  NAND3_X1 U6685 ( .A1(n5532), .A2(n5531), .A3(n5533), .ZN(n5538) );
  INV_X1 U6686 ( .A(n5533), .ZN(n5535) );
  NAND2_X1 U6687 ( .A1(n5549), .A2(n5662), .ZN(n5534) );
  NAND3_X1 U6688 ( .A1(n5536), .A2(n5535), .A3(n5534), .ZN(n5537) );
  NAND2_X1 U6689 ( .A1(n5538), .A2(n5537), .ZN(n5836) );
  NOR2_X1 U6690 ( .A1(n5836), .A2(n6193), .ZN(n5539) );
  AOI211_X1 U6691 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5541), .A(n5540), .B(n5539), .ZN(n5542) );
  OAI211_X1 U6692 ( .C1(REIP_REG_30__SCAN_IN), .C2(n5544), .A(n5543), .B(n5542), .ZN(U2797) );
  INV_X1 U6693 ( .A(n5545), .ZN(n5547) );
  AOI21_X1 U6694 ( .B1(n5547), .B2(n5605), .A(n5546), .ZN(n5548) );
  NAND2_X1 U6695 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  AOI22_X1 U6696 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6197), .B1(n6207), 
        .B2(n5552), .ZN(n5554) );
  NAND2_X1 U6697 ( .A1(n6198), .A2(EBX_REG_29__SCAN_IN), .ZN(n5553) );
  OAI211_X1 U6698 ( .C1(n5565), .C2(n6704), .A(n5554), .B(n5553), .ZN(n5556)
         );
  NOR3_X1 U6699 ( .A1(n5566), .A2(REIP_REG_29__SCAN_IN), .A3(n6705), .ZN(n5555) );
  AOI211_X1 U6700 ( .C1(n6202), .C2(n5844), .A(n5556), .B(n5555), .ZN(n5557)
         );
  OAI21_X1 U6701 ( .B1(n5687), .B2(n6177), .A(n5557), .ZN(U2798) );
  AOI21_X1 U6702 ( .B1(n5558), .B2(n5571), .A(n4241), .ZN(n5719) );
  INV_X1 U6703 ( .A(n5719), .ZN(n5690) );
  INV_X1 U6704 ( .A(n5559), .ZN(n5562) );
  INV_X1 U6705 ( .A(n5575), .ZN(n5561) );
  AOI21_X1 U6706 ( .B1(n5562), .B2(n5561), .A(n5560), .ZN(n5852) );
  OAI22_X1 U6707 ( .A1(n6958), .A2(n6171), .B1(n6188), .B2(n5717), .ZN(n5563)
         );
  AOI21_X1 U6708 ( .B1(n6198), .B2(EBX_REG_28__SCAN_IN), .A(n5563), .ZN(n5564)
         );
  OAI21_X1 U6709 ( .B1(n6705), .B2(n5565), .A(n5564), .ZN(n5568) );
  NOR2_X1 U6710 ( .A1(n5566), .A2(REIP_REG_28__SCAN_IN), .ZN(n5567) );
  AOI211_X1 U6711 ( .C1(n6202), .C2(n5852), .A(n5568), .B(n5567), .ZN(n5569)
         );
  OAI21_X1 U6712 ( .B1(n5690), .B2(n6177), .A(n5569), .ZN(U2799) );
  OAI21_X1 U6713 ( .B1(n5570), .B2(n5572), .A(n5571), .ZN(n5723) );
  AND2_X1 U6714 ( .A1(n3176), .A2(n5573), .ZN(n5574) );
  OR2_X1 U6715 ( .A1(n5575), .A2(n5574), .ZN(n5861) );
  AOI22_X1 U6716 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6197), .B1(n6207), 
        .B2(n5726), .ZN(n5577) );
  NAND2_X1 U6717 ( .A1(n6198), .A2(EBX_REG_27__SCAN_IN), .ZN(n5576) );
  OAI211_X1 U6718 ( .C1(n5861), .C2(n6193), .A(n5577), .B(n5576), .ZN(n5578)
         );
  INV_X1 U6719 ( .A(n5578), .ZN(n5582) );
  INV_X1 U6720 ( .A(n5579), .ZN(n5580) );
  NAND3_X1 U6721 ( .A1(n5987), .A2(n5580), .A3(n5583), .ZN(n5581) );
  OAI211_X1 U6722 ( .C1(n5976), .C2(n5583), .A(n5582), .B(n5581), .ZN(n5584)
         );
  INV_X1 U6723 ( .A(n5584), .ZN(n5585) );
  OAI21_X1 U6724 ( .B1(n5723), .B2(n6177), .A(n5585), .ZN(U2800) );
  NOR2_X1 U6725 ( .A1(n5587), .A2(n5588), .ZN(n5589) );
  OR2_X1 U6726 ( .A1(n5586), .A2(n5589), .ZN(n5758) );
  NOR2_X1 U6727 ( .A1(n6185), .A2(n5590), .ZN(n6010) );
  INV_X1 U6728 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U6729 ( .A1(n6692), .A2(n5591), .ZN(n6014) );
  INV_X1 U6730 ( .A(n6014), .ZN(n5592) );
  OAI21_X1 U6731 ( .B1(n6010), .B2(n5592), .A(REIP_REG_22__SCAN_IN), .ZN(n5598) );
  XNOR2_X1 U6732 ( .A(n5652), .B(n5640), .ZN(n5902) );
  INV_X1 U6733 ( .A(n5902), .ZN(n5596) );
  OAI22_X1 U6734 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6001), .B1(n5645), .B2(
        n6172), .ZN(n5595) );
  INV_X1 U6735 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5593) );
  OAI22_X1 U6736 ( .A1(n5593), .A2(n6171), .B1(n5760), .B2(n6188), .ZN(n5594)
         );
  AOI211_X1 U6737 ( .C1(n6202), .C2(n5596), .A(n5595), .B(n5594), .ZN(n5597)
         );
  OAI211_X1 U6738 ( .C1(n5758), .C2(n6177), .A(n5598), .B(n5597), .ZN(U2805)
         );
  AND2_X1 U6739 ( .A1(n5600), .A2(n5601), .ZN(n5602) );
  NOR2_X1 U6740 ( .A1(n5599), .A2(n5602), .ZN(n6046) );
  INV_X1 U6741 ( .A(n6046), .ZN(n5655) );
  INV_X1 U6742 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6691) );
  INV_X1 U6743 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6693) );
  OAI21_X1 U6744 ( .B1(n6020), .B2(n6691), .A(n6693), .ZN(n5611) );
  INV_X1 U6745 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5603) );
  OAI22_X1 U6746 ( .A1(n5603), .A2(n6171), .B1(n5773), .B2(n6188), .ZN(n5610)
         );
  INV_X1 U6747 ( .A(n5664), .ZN(n5606) );
  MUX2_X1 U6748 ( .A(n5606), .B(n5605), .S(n5604), .Z(n5608) );
  XNOR2_X1 U6749 ( .A(n5608), .B(n5607), .ZN(n5922) );
  INV_X1 U6750 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5656) );
  OAI22_X1 U6751 ( .A1(n5922), .A2(n6193), .B1(n5656), .B2(n6172), .ZN(n5609)
         );
  AOI211_X1 U6752 ( .C1(n6010), .C2(n5611), .A(n5610), .B(n5609), .ZN(n5612)
         );
  OAI21_X1 U6753 ( .B1(n5655), .B2(n6177), .A(n5612), .ZN(U2807) );
  INV_X1 U6754 ( .A(n5830), .ZN(n5614) );
  OAI22_X1 U6755 ( .A1(n5614), .A2(n5678), .B1(n5613), .B2(n6221), .ZN(U2828)
         );
  OAI222_X1 U6756 ( .A1(n5680), .A2(n5684), .B1(n6221), .B2(n6843), .C1(n5836), 
        .C2(n5678), .ZN(U2829) );
  AOI22_X1 U6757 ( .A1(n5844), .A2(n6217), .B1(n5634), .B2(EBX_REG_29__SCAN_IN), .ZN(n5615) );
  OAI21_X1 U6758 ( .B1(n5687), .B2(n5680), .A(n5615), .ZN(U2830) );
  AOI22_X1 U6759 ( .A1(n5852), .A2(n6217), .B1(n5634), .B2(EBX_REG_28__SCAN_IN), .ZN(n5616) );
  OAI21_X1 U6760 ( .B1(n5690), .B2(n5680), .A(n5616), .ZN(U2831) );
  INV_X1 U6761 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5617) );
  OAI222_X1 U6762 ( .A1(n5680), .A2(n5723), .B1(n6221), .B2(n5617), .C1(n5861), 
        .C2(n5678), .ZN(U2832) );
  NOR2_X1 U6763 ( .A1(n5618), .A2(n5619), .ZN(n5620) );
  OR2_X1 U6764 ( .A1(n5570), .A2(n5620), .ZN(n5733) );
  INV_X1 U6765 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U6766 ( .A1(n3175), .A2(n5621), .ZN(n5622) );
  NAND2_X1 U6767 ( .A1(n3176), .A2(n5622), .ZN(n5975) );
  OAI222_X1 U6768 ( .A1(n5680), .A2(n5733), .B1(n6221), .B2(n5623), .C1(n5975), 
        .C2(n5678), .ZN(U2833) );
  NAND2_X1 U6769 ( .A1(n5642), .A2(n5633), .ZN(n5626) );
  INV_X1 U6770 ( .A(n5624), .ZN(n5625) );
  NAND2_X1 U6771 ( .A1(n5626), .A2(n5625), .ZN(n5627) );
  NAND2_X1 U6772 ( .A1(n5627), .A2(n3175), .ZN(n5984) );
  INV_X1 U6773 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5630) );
  AND2_X1 U6774 ( .A1(n3183), .A2(n5628), .ZN(n5629) );
  OAI222_X1 U6775 ( .A1(n5678), .A2(n5984), .B1(n6221), .B2(n5630), .C1(n5680), 
        .C2(n6032), .ZN(U2834) );
  XOR2_X1 U6776 ( .A(n5632), .B(n5631), .Z(n6036) );
  INV_X1 U6777 ( .A(n6036), .ZN(n5636) );
  XOR2_X1 U6778 ( .A(n5633), .B(n5642), .Z(n5995) );
  AOI22_X1 U6779 ( .A1(n5995), .A2(n6217), .B1(EBX_REG_24__SCAN_IN), .B2(n5634), .ZN(n5635) );
  OAI21_X1 U6780 ( .B1(n5636), .B2(n5680), .A(n5635), .ZN(U2835) );
  OR2_X1 U6781 ( .A1(n5586), .A2(n5637), .ZN(n5638) );
  NAND2_X1 U6782 ( .A1(n5631), .A2(n5638), .ZN(n6003) );
  AOI21_X1 U6783 ( .B1(n5652), .B2(n5640), .A(n5639), .ZN(n5641) );
  OR2_X1 U6784 ( .A1(n5642), .A2(n5641), .ZN(n6002) );
  OAI22_X1 U6785 ( .A1(n6002), .A2(n5678), .B1(n6888), .B2(n6221), .ZN(n5643)
         );
  INV_X1 U6786 ( .A(n5643), .ZN(n5644) );
  OAI21_X1 U6787 ( .B1(n6003), .B2(n5680), .A(n5644), .ZN(U2836) );
  OAI22_X1 U6788 ( .A1(n5902), .A2(n5678), .B1(n5645), .B2(n6221), .ZN(n5646)
         );
  INV_X1 U6789 ( .A(n5646), .ZN(n5647) );
  OAI21_X1 U6790 ( .B1(n5758), .B2(n5680), .A(n5647), .ZN(U2837) );
  NOR2_X1 U6791 ( .A1(n5599), .A2(n5648), .ZN(n5649) );
  OR2_X1 U6792 ( .A1(n5587), .A2(n5649), .ZN(n6042) );
  INV_X1 U6793 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5654) );
  AND2_X1 U6794 ( .A1(n5651), .A2(n5650), .ZN(n5653) );
  OR2_X1 U6795 ( .A1(n5653), .A2(n5652), .ZN(n6012) );
  OAI222_X1 U6796 ( .A1(n5680), .A2(n6042), .B1(n6221), .B2(n5654), .C1(n6012), 
        .C2(n5678), .ZN(U2838) );
  OAI222_X1 U6797 ( .A1(n5678), .A2(n5922), .B1(n6221), .B2(n5656), .C1(n5680), 
        .C2(n5655), .ZN(U2839) );
  INV_X1 U6798 ( .A(n5600), .ZN(n5659) );
  AOI21_X1 U6799 ( .B1(n5660), .B2(n5672), .A(n5659), .ZN(n5780) );
  INV_X1 U6800 ( .A(n5780), .ZN(n6025) );
  INV_X1 U6801 ( .A(n5661), .ZN(n5663) );
  MUX2_X1 U6802 ( .A(n5664), .B(n5663), .S(n5662), .Z(n5666) );
  NAND2_X1 U6803 ( .A1(n6067), .A2(n5666), .ZN(n5668) );
  XOR2_X1 U6804 ( .A(n5665), .B(n5668), .Z(n6024) );
  INV_X1 U6805 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6955) );
  OAI222_X1 U6806 ( .A1(n6025), .A2(n5680), .B1(n5678), .B2(n6024), .C1(n6221), 
        .C2(n6955), .ZN(U2840) );
  OR2_X1 U6807 ( .A1(n6067), .A2(n5666), .ZN(n5667) );
  NAND2_X1 U6808 ( .A1(n5668), .A2(n5667), .ZN(n6114) );
  NAND2_X1 U6809 ( .A1(n5669), .A2(n5670), .ZN(n5671) );
  AND2_X1 U6810 ( .A1(n5672), .A2(n5671), .ZN(n6222) );
  INV_X1 U6811 ( .A(n6222), .ZN(n5673) );
  OAI222_X1 U6812 ( .A1(n5678), .A2(n6114), .B1(n6221), .B2(n5472), .C1(n5673), 
        .C2(n5680), .ZN(U2841) );
  AOI21_X1 U6813 ( .B1(n5674), .B2(n5402), .A(n3173), .ZN(n6229) );
  INV_X1 U6814 ( .A(n6229), .ZN(n5681) );
  INV_X1 U6815 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5679) );
  AND2_X1 U6816 ( .A1(n5676), .A2(n5675), .ZN(n5677) );
  OR2_X1 U6817 ( .A1(n5677), .A2(n6066), .ZN(n6130) );
  OAI222_X1 U6818 ( .A1(n5681), .A2(n5680), .B1(n6221), .B2(n5679), .C1(n6130), 
        .C2(n5678), .ZN(U2843) );
  AOI22_X1 U6819 ( .A1(n6228), .A2(DATAI_30_), .B1(n6230), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U6820 ( .A1(n6231), .A2(DATAI_14_), .ZN(n5682) );
  OAI211_X1 U6821 ( .C1(n5684), .C2(n5697), .A(n5683), .B(n5682), .ZN(U2861)
         );
  AOI22_X1 U6822 ( .A1(n6228), .A2(DATAI_29_), .B1(n6230), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U6823 ( .A1(n6231), .A2(DATAI_13_), .ZN(n5685) );
  OAI211_X1 U6824 ( .C1(n5687), .C2(n5697), .A(n5686), .B(n5685), .ZN(U2862)
         );
  AOI22_X1 U6825 ( .A1(n6228), .A2(DATAI_28_), .B1(n6230), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U6826 ( .A1(n6231), .A2(DATAI_12_), .ZN(n5688) );
  OAI211_X1 U6827 ( .C1(n5690), .C2(n5697), .A(n5689), .B(n5688), .ZN(U2863)
         );
  AOI22_X1 U6828 ( .A1(n6228), .A2(DATAI_27_), .B1(n6230), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U6829 ( .A1(n6231), .A2(DATAI_11_), .ZN(n5691) );
  OAI211_X1 U6830 ( .C1(n5723), .C2(n5697), .A(n5692), .B(n5691), .ZN(U2864)
         );
  AOI22_X1 U6831 ( .A1(n6231), .A2(DATAI_7_), .B1(n6230), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U6832 ( .A1(n6228), .A2(DATAI_23_), .ZN(n5693) );
  OAI211_X1 U6833 ( .C1(n6003), .C2(n5697), .A(n5694), .B(n5693), .ZN(U2868)
         );
  AOI22_X1 U6834 ( .A1(n6231), .A2(DATAI_3_), .B1(n6230), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U6835 ( .A1(n6228), .A2(DATAI_19_), .ZN(n5695) );
  OAI211_X1 U6836 ( .C1(n6025), .C2(n5697), .A(n5696), .B(n5695), .ZN(U2872)
         );
  NAND2_X1 U6837 ( .A1(n5700), .A2(n5699), .ZN(n5701) );
  XNOR2_X1 U6838 ( .A(n5701), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5841)
         );
  NAND2_X1 U6839 ( .A1(n6353), .A2(REIP_REG_30__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U6840 ( .A1(n6299), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5702)
         );
  OAI211_X1 U6841 ( .C1(n6308), .C2(n5703), .A(n5835), .B(n5702), .ZN(n5704)
         );
  AOI21_X1 U6842 ( .B1(n5705), .B2(n4244), .A(n5704), .ZN(n5706) );
  OAI21_X1 U6843 ( .B1(n5841), .B2(n6294), .A(n5706), .ZN(U2956) );
  INV_X1 U6844 ( .A(n5845), .ZN(n5715) );
  NAND2_X1 U6845 ( .A1(n5708), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5713) );
  INV_X1 U6846 ( .A(n5709), .ZN(n5712) );
  NAND3_X1 U6847 ( .A1(n5721), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(n5710), .ZN(n5711) );
  OAI211_X1 U6848 ( .C1(n5707), .C2(n5713), .A(n5712), .B(n5711), .ZN(n5714)
         );
  NAND2_X1 U6849 ( .A1(n6353), .A2(REIP_REG_28__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U6850 ( .A1(n6299), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5716)
         );
  OAI211_X1 U6851 ( .C1(n6308), .C2(n5717), .A(n5853), .B(n5716), .ZN(n5718)
         );
  AOI21_X1 U6852 ( .B1(n5719), .B2(n4244), .A(n5718), .ZN(n5720) );
  OAI21_X1 U6853 ( .B1(n5858), .B2(n6294), .A(n5720), .ZN(U2958) );
  NAND2_X1 U6854 ( .A1(n5707), .A2(n5721), .ZN(n5722) );
  XNOR2_X1 U6855 ( .A(n5722), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5866)
         );
  NAND2_X1 U6856 ( .A1(n6353), .A2(REIP_REG_27__SCAN_IN), .ZN(n5860) );
  OAI21_X1 U6857 ( .B1(n6063), .B2(n7026), .A(n5860), .ZN(n5725) );
  NOR2_X1 U6858 ( .A1(n5723), .A2(n6292), .ZN(n5724) );
  AOI211_X1 U6859 ( .C1(n6276), .C2(n5726), .A(n5725), .B(n5724), .ZN(n5727)
         );
  OAI21_X1 U6860 ( .B1(n5866), .B2(n6294), .A(n5727), .ZN(U2959) );
  INV_X1 U6861 ( .A(n5728), .ZN(n5729) );
  NOR2_X1 U6862 ( .A1(n5730), .A2(n5729), .ZN(n5732) );
  XOR2_X1 U6863 ( .A(n5732), .B(n5731), .Z(n5874) );
  NAND2_X1 U6864 ( .A1(n6353), .A2(REIP_REG_26__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U6865 ( .A1(n6299), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5734)
         );
  OAI211_X1 U6866 ( .C1(n6308), .C2(n5981), .A(n5870), .B(n5734), .ZN(n5735)
         );
  AOI21_X1 U6867 ( .B1(n6029), .B2(n4244), .A(n5735), .ZN(n5736) );
  OAI21_X1 U6868 ( .B1(n5874), .B2(n6294), .A(n5736), .ZN(U2960) );
  NAND2_X1 U6869 ( .A1(n6353), .A2(REIP_REG_25__SCAN_IN), .ZN(n5876) );
  OAI21_X1 U6870 ( .B1(n6063), .B2(n5737), .A(n5876), .ZN(n5738) );
  AOI21_X1 U6871 ( .B1(n6276), .B2(n5983), .A(n5738), .ZN(n5741) );
  OAI21_X1 U6872 ( .B1(n5739), .B2(n3208), .A(n3210), .ZN(n5875) );
  NAND2_X1 U6873 ( .A1(n5875), .A2(n6303), .ZN(n5740) );
  OAI211_X1 U6874 ( .C1(n6032), .C2(n6292), .A(n5741), .B(n5740), .ZN(U2961)
         );
  XNOR2_X1 U6875 ( .A(n3171), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5771)
         );
  XNOR2_X1 U6876 ( .A(n6271), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5764)
         );
  NAND2_X1 U6877 ( .A1(n3171), .A2(n6985), .ZN(n5755) );
  NOR2_X1 U6878 ( .A1(n5763), .A2(n5755), .ZN(n5749) );
  XNOR2_X1 U6879 ( .A(n5743), .B(n5742), .ZN(n5888) );
  INV_X1 U6880 ( .A(n5994), .ZN(n5745) );
  AND2_X1 U6881 ( .A1(n6353), .A2(REIP_REG_24__SCAN_IN), .ZN(n5886) );
  AOI21_X1 U6882 ( .B1(n6299), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5886), 
        .ZN(n5744) );
  OAI21_X1 U6883 ( .B1(n5745), .B2(n6308), .A(n5744), .ZN(n5746) );
  AOI21_X1 U6884 ( .B1(n6036), .B2(n4244), .A(n5746), .ZN(n5747) );
  OAI21_X1 U6885 ( .B1(n5888), .B2(n6294), .A(n5747), .ZN(U2962) );
  INV_X1 U6886 ( .A(n5897), .ZN(n5812) );
  INV_X1 U6887 ( .A(n5923), .ZN(n5748) );
  NOR3_X1 U6888 ( .A1(n3171), .A2(n5812), .A3(n5748), .ZN(n5750) );
  AOI21_X1 U6889 ( .B1(n5750), .B2(n5777), .A(n5749), .ZN(n5751) );
  XNOR2_X1 U6890 ( .A(n5751), .B(n5889), .ZN(n5896) );
  NAND2_X1 U6891 ( .A1(n6353), .A2(REIP_REG_23__SCAN_IN), .ZN(n5891) );
  OAI21_X1 U6892 ( .B1(n6063), .B2(n6009), .A(n5891), .ZN(n5753) );
  NOR2_X1 U6893 ( .A1(n6003), .A2(n6292), .ZN(n5752) );
  AOI211_X1 U6894 ( .C1(n6276), .C2(n6000), .A(n5753), .B(n5752), .ZN(n5754)
         );
  OAI21_X1 U6895 ( .B1(n5896), .B2(n6294), .A(n5754), .ZN(U2963) );
  OAI21_X1 U6896 ( .B1(n3171), .B2(n6985), .A(n5755), .ZN(n5757) );
  XOR2_X1 U6897 ( .A(n5757), .B(n5756), .Z(n5905) );
  INV_X1 U6898 ( .A(n5758), .ZN(n6039) );
  NAND2_X1 U6899 ( .A1(n6353), .A2(REIP_REG_22__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U6900 ( .A1(n6299), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5759)
         );
  OAI211_X1 U6901 ( .C1(n6308), .C2(n5760), .A(n5901), .B(n5759), .ZN(n5761)
         );
  AOI21_X1 U6902 ( .B1(n6039), .B2(n4244), .A(n5761), .ZN(n5762) );
  OAI21_X1 U6903 ( .B1(n5905), .B2(n6294), .A(n5762), .ZN(U2964) );
  OAI21_X1 U6904 ( .B1(n5765), .B2(n5764), .A(n5763), .ZN(n5907) );
  NAND2_X1 U6905 ( .A1(n5907), .A2(n6303), .ZN(n5769) );
  NAND2_X1 U6906 ( .A1(n6353), .A2(REIP_REG_21__SCAN_IN), .ZN(n5908) );
  OAI21_X1 U6907 ( .B1(n6063), .B2(n5766), .A(n5908), .ZN(n5767) );
  AOI21_X1 U6908 ( .B1(n6276), .B2(n6011), .A(n5767), .ZN(n5768) );
  OAI211_X1 U6909 ( .C1(n6292), .C2(n6042), .A(n5769), .B(n5768), .ZN(U2965)
         );
  XOR2_X1 U6910 ( .A(n5771), .B(n5770), .Z(n5928) );
  NAND2_X1 U6911 ( .A1(n6353), .A2(REIP_REG_20__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U6912 ( .A1(n6299), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5772)
         );
  OAI211_X1 U6913 ( .C1(n6308), .C2(n5773), .A(n5921), .B(n5772), .ZN(n5774)
         );
  AOI21_X1 U6914 ( .B1(n6046), .B2(n4244), .A(n5774), .ZN(n5775) );
  OAI21_X1 U6915 ( .B1(n5928), .B2(n6294), .A(n5775), .ZN(U2966) );
  XNOR2_X1 U6916 ( .A(n6271), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5776)
         );
  XNOR2_X1 U6917 ( .A(n5777), .B(n5776), .ZN(n5935) );
  NAND2_X1 U6918 ( .A1(n6276), .A2(n6022), .ZN(n5778) );
  NAND2_X1 U6919 ( .A1(n6353), .A2(REIP_REG_19__SCAN_IN), .ZN(n5929) );
  OAI211_X1 U6920 ( .C1(n6063), .C2(n6957), .A(n5778), .B(n5929), .ZN(n5779)
         );
  AOI21_X1 U6921 ( .B1(n5780), .B2(n4244), .A(n5779), .ZN(n5781) );
  OAI21_X1 U6922 ( .B1(n5935), .B2(n6294), .A(n5781), .ZN(U2967) );
  INV_X1 U6923 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6078) );
  NOR2_X1 U6924 ( .A1(n6271), .A2(n6078), .ZN(n5787) );
  INV_X1 U6925 ( .A(n5784), .ZN(n5785) );
  OAI21_X1 U6926 ( .B1(n3252), .B2(n5787), .A(n5785), .ZN(n5786) );
  OAI21_X1 U6927 ( .B1(n5782), .B2(n5787), .A(n5786), .ZN(n6074) );
  INV_X1 U6928 ( .A(n6127), .ZN(n5789) );
  AOI22_X1 U6929 ( .A1(n6299), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6353), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5788) );
  OAI21_X1 U6930 ( .B1(n6308), .B2(n5789), .A(n5788), .ZN(n5790) );
  AOI21_X1 U6931 ( .B1(n6229), .B2(n4244), .A(n5790), .ZN(n5791) );
  OAI21_X1 U6932 ( .B1(n6074), .B2(n6294), .A(n5791), .ZN(U2970) );
  INV_X1 U6933 ( .A(n5793), .ZN(n5795) );
  NAND2_X1 U6934 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  XNOR2_X1 U6935 ( .A(n5792), .B(n5796), .ZN(n5956) );
  AOI22_X1 U6936 ( .A1(n6299), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6353), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5797) );
  OAI21_X1 U6937 ( .B1(n5798), .B2(n6308), .A(n5797), .ZN(n5799) );
  AOI21_X1 U6938 ( .B1(n5800), .B2(n4244), .A(n5799), .ZN(n5801) );
  OAI21_X1 U6939 ( .B1(n5956), .B2(n6294), .A(n5801), .ZN(U2971) );
  AND2_X1 U6940 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U6941 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5802), .ZN(n5951) );
  INV_X1 U6942 ( .A(n5951), .ZN(n5949) );
  NAND3_X1 U6943 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5949), .ZN(n5939) );
  NOR2_X1 U6944 ( .A1(n6054), .A2(n5939), .ZN(n5938) );
  AND2_X1 U6945 ( .A1(n5803), .A2(n5938), .ZN(n5918) );
  NAND4_X1 U6946 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(INSTADDRPOINTER_REG_19__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5819) );
  INV_X1 U6947 ( .A(n5819), .ZN(n5808) );
  NAND2_X1 U6948 ( .A1(n5918), .A2(n5808), .ZN(n5823) );
  NAND2_X1 U6949 ( .A1(n5823), .A2(n5804), .ZN(n5811) );
  INV_X1 U6950 ( .A(n5939), .ZN(n5806) );
  NAND2_X1 U6951 ( .A1(n5806), .A2(n5805), .ZN(n5820) );
  INV_X1 U6952 ( .A(n5820), .ZN(n5807) );
  OR2_X1 U6953 ( .A1(n6348), .A2(n5807), .ZN(n5916) );
  OR2_X1 U6954 ( .A1(n6348), .A2(n5808), .ZN(n5809) );
  AND2_X1 U6955 ( .A1(n5916), .A2(n5809), .ZN(n5810) );
  NAND2_X1 U6956 ( .A1(n5811), .A2(n5810), .ZN(n5906) );
  AND2_X1 U6957 ( .A1(n6350), .A2(n5812), .ZN(n5813) );
  OR2_X1 U6958 ( .A1(n5906), .A2(n5813), .ZN(n5894) );
  AOI21_X1 U6959 ( .B1(n5815), .B2(n5814), .A(n5824), .ZN(n5816) );
  NOR2_X1 U6960 ( .A1(n5894), .A2(n5816), .ZN(n5884) );
  OAI21_X1 U6961 ( .B1(n6321), .B2(n5826), .A(n5884), .ZN(n5864) );
  AOI21_X1 U6962 ( .B1(n5845), .B2(n6350), .A(n5864), .ZN(n5848) );
  OAI21_X1 U6963 ( .B1(n5827), .B2(n6910), .A(n6350), .ZN(n5817) );
  NAND2_X1 U6964 ( .A1(n5848), .A2(n5817), .ZN(n5839) );
  INV_X1 U6965 ( .A(n5818), .ZN(n5829) );
  NOR2_X1 U6966 ( .A1(n5820), .A2(n5819), .ZN(n5821) );
  NAND2_X1 U6967 ( .A1(n6399), .A2(n5821), .ZN(n5822) );
  NAND2_X1 U6968 ( .A1(n5823), .A2(n5822), .ZN(n5910) );
  NAND2_X1 U6969 ( .A1(n5910), .A2(n5897), .ZN(n5882) );
  INV_X1 U6970 ( .A(n5824), .ZN(n5825) );
  NOR2_X1 U6971 ( .A1(n5882), .A2(n5825), .ZN(n5868) );
  NAND2_X1 U6972 ( .A1(n5868), .A2(n5826), .ZN(n5859) );
  OR3_X1 U6973 ( .A1(n5859), .A2(n5845), .A3(n6910), .ZN(n5834) );
  NOR3_X1 U6974 ( .A1(n5834), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5827), 
        .ZN(n5828) );
  AOI211_X1 U6975 ( .C1(n5839), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5829), .B(n5828), .ZN(n5832) );
  NAND2_X1 U6976 ( .A1(n5830), .A2(n6383), .ZN(n5831) );
  OAI211_X1 U6977 ( .C1(n5833), .C2(n6370), .A(n5832), .B(n5831), .ZN(U2987)
         );
  NOR2_X1 U6978 ( .A1(n5834), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5838)
         );
  OAI21_X1 U6979 ( .B1(n5836), .B2(n6390), .A(n5835), .ZN(n5837) );
  AOI211_X1 U6980 ( .C1(INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n5839), .A(n5838), .B(n5837), .ZN(n5840) );
  OAI21_X1 U6981 ( .B1(n5841), .B2(n6370), .A(n5840), .ZN(U2988) );
  INV_X1 U6982 ( .A(n5842), .ZN(n5843) );
  AOI21_X1 U6983 ( .B1(n5844), .B2(n6383), .A(n5843), .ZN(n5847) );
  OR3_X1 U6984 ( .A1(n5859), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5845), 
        .ZN(n5846) );
  OAI211_X1 U6985 ( .C1(n5848), .C2(n6910), .A(n5847), .B(n5846), .ZN(n5849)
         );
  INV_X1 U6986 ( .A(n5849), .ZN(n5850) );
  OAI21_X1 U6987 ( .B1(n5851), .B2(n6370), .A(n5850), .ZN(U2989) );
  XNOR2_X1 U6988 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U6989 ( .A1(n5852), .A2(n6383), .ZN(n5854) );
  OAI211_X1 U6990 ( .C1(n5855), .C2(n5859), .A(n5854), .B(n5853), .ZN(n5856)
         );
  AOI21_X1 U6991 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5864), .A(n5856), 
        .ZN(n5857) );
  OAI21_X1 U6992 ( .B1(n5858), .B2(n6370), .A(n5857), .ZN(U2990) );
  NOR2_X1 U6993 ( .A1(n5859), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5863)
         );
  OAI21_X1 U6994 ( .B1(n5861), .B2(n6390), .A(n5860), .ZN(n5862) );
  AOI211_X1 U6995 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5864), .A(n5863), .B(n5862), .ZN(n5865) );
  OAI21_X1 U6996 ( .B1(n5866), .B2(n6370), .A(n5865), .ZN(U2991) );
  NAND2_X1 U6997 ( .A1(n5868), .A2(n6887), .ZN(n5877) );
  AOI21_X1 U6998 ( .B1(n5877), .B2(n5884), .A(n5867), .ZN(n5872) );
  NAND3_X1 U6999 ( .A1(n5868), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n5867), .ZN(n5869) );
  OAI211_X1 U7000 ( .C1(n5975), .C2(n6390), .A(n5870), .B(n5869), .ZN(n5871)
         );
  NOR2_X1 U7001 ( .A1(n5872), .A2(n5871), .ZN(n5873) );
  OAI21_X1 U7002 ( .B1(n5874), .B2(n6370), .A(n5873), .ZN(U2992) );
  INV_X1 U7003 ( .A(n5875), .ZN(n5881) );
  INV_X1 U7004 ( .A(n5884), .ZN(n5879) );
  OAI211_X1 U7005 ( .C1(n6390), .C2(n5984), .A(n5877), .B(n5876), .ZN(n5878)
         );
  AOI21_X1 U7006 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5879), .A(n5878), 
        .ZN(n5880) );
  OAI21_X1 U7007 ( .B1(n5881), .B2(n6370), .A(n5880), .ZN(U2993) );
  INV_X1 U7008 ( .A(n5882), .ZN(n5890) );
  AOI21_X1 U7009 ( .B1(n5890), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5883) );
  NOR2_X1 U7010 ( .A1(n5884), .A2(n5883), .ZN(n5885) );
  AOI211_X1 U7011 ( .C1(n6383), .C2(n5995), .A(n5886), .B(n5885), .ZN(n5887)
         );
  OAI21_X1 U7012 ( .B1(n5888), .B2(n6370), .A(n5887), .ZN(U2994) );
  NAND2_X1 U7013 ( .A1(n5890), .A2(n5889), .ZN(n5892) );
  OAI211_X1 U7014 ( .C1(n6390), .C2(n6002), .A(n5892), .B(n5891), .ZN(n5893)
         );
  AOI21_X1 U7015 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5894), .A(n5893), 
        .ZN(n5895) );
  OAI21_X1 U7016 ( .B1(n5896), .B2(n6370), .A(n5895), .ZN(U2995) );
  NOR2_X1 U7017 ( .A1(n5898), .A2(n5897), .ZN(n5899) );
  NAND2_X1 U7018 ( .A1(n5910), .A2(n5899), .ZN(n5900) );
  OAI211_X1 U7019 ( .C1(n5902), .C2(n6390), .A(n5901), .B(n5900), .ZN(n5903)
         );
  AOI21_X1 U7020 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5906), .A(n5903), 
        .ZN(n5904) );
  OAI21_X1 U7021 ( .B1(n5905), .B2(n6370), .A(n5904), .ZN(U2996) );
  INV_X1 U7022 ( .A(n5906), .ZN(n5914) );
  NAND2_X1 U7023 ( .A1(n5907), .A2(n6396), .ZN(n5912) );
  OAI21_X1 U7024 ( .B1(n6012), .B2(n6390), .A(n5908), .ZN(n5909) );
  AOI21_X1 U7025 ( .B1(n5913), .B2(n5910), .A(n5909), .ZN(n5911) );
  OAI211_X1 U7026 ( .C1(n5914), .C2(n5913), .A(n5912), .B(n5911), .ZN(U2997)
         );
  INV_X1 U7027 ( .A(n5915), .ZN(n5920) );
  OAI21_X1 U7028 ( .B1(n5918), .B2(n5917), .A(n5916), .ZN(n6068) );
  INV_X1 U7029 ( .A(n6068), .ZN(n5919) );
  OAI21_X1 U7030 ( .B1(n5920), .B2(n6321), .A(n5919), .ZN(n5933) );
  OAI21_X1 U7031 ( .B1(n5922), .B2(n6390), .A(n5921), .ZN(n5926) );
  NAND3_X1 U7032 ( .A1(n6311), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5938), .ZN(n5930) );
  NOR3_X1 U7033 ( .A1(n5930), .A2(n5924), .A3(n5923), .ZN(n5925) );
  AOI211_X1 U7034 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n5933), .A(n5926), .B(n5925), .ZN(n5927) );
  OAI21_X1 U7035 ( .B1(n5928), .B2(n6370), .A(n5927), .ZN(U2998) );
  OAI21_X1 U7036 ( .B1(n6024), .B2(n6390), .A(n5929), .ZN(n5932) );
  NOR2_X1 U7037 ( .A1(n5930), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5931)
         );
  AOI211_X1 U7038 ( .C1(n5933), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5932), .B(n5931), .ZN(n5934) );
  OAI21_X1 U7039 ( .B1(n5935), .B2(n6370), .A(n5934), .ZN(U2999) );
  NOR3_X1 U7040 ( .A1(n5784), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6271), 
        .ZN(n6053) );
  NOR3_X1 U7041 ( .A1(n5782), .A2(n3171), .A3(n6054), .ZN(n5936) );
  AOI21_X1 U7042 ( .B1(n6053), .B2(n6054), .A(n5936), .ZN(n5937) );
  XNOR2_X1 U7043 ( .A(n5937), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6049)
         );
  INV_X1 U7044 ( .A(n6049), .ZN(n5948) );
  INV_X1 U7045 ( .A(n6114), .ZN(n5946) );
  NAND2_X1 U7046 ( .A1(n5938), .A2(n6311), .ZN(n5944) );
  NOR2_X1 U7047 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5939), .ZN(n6065)
         );
  AOI21_X1 U7048 ( .B1(n5940), .B2(n6065), .A(n6068), .ZN(n5942) );
  NAND2_X1 U7049 ( .A1(n6353), .A2(REIP_REG_18__SCAN_IN), .ZN(n5941) );
  OAI221_X1 U7050 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5944), .C1(
        n5943), .C2(n5942), .A(n5941), .ZN(n5945) );
  AOI21_X1 U7051 ( .B1(n5946), .B2(n6383), .A(n5945), .ZN(n5947) );
  OAI21_X1 U7052 ( .B1(n5948), .B2(n6370), .A(n5947), .ZN(U3000) );
  NAND2_X1 U7053 ( .A1(n5949), .A2(n6311), .ZN(n6072) );
  NOR2_X1 U7054 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n6072), .ZN(n5950)
         );
  AOI211_X1 U7055 ( .C1(n5951), .C2(n6350), .A(n5950), .B(n6312), .ZN(n6079)
         );
  AOI21_X1 U7056 ( .B1(n6073), .B2(n6072), .A(n6079), .ZN(n5954) );
  OAI22_X1 U7057 ( .A1(n5952), .A2(n6390), .B1(n6686), .B2(n6388), .ZN(n5953)
         );
  NOR2_X1 U7058 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  OAI21_X1 U7059 ( .B1(n5956), .B2(n6370), .A(n5955), .ZN(U3003) );
  INV_X1 U7060 ( .A(n5957), .ZN(n5967) );
  OAI21_X1 U7061 ( .B1(n6390), .B2(n5959), .A(n5958), .ZN(n5960) );
  AOI21_X1 U7062 ( .B1(n6396), .B2(n5961), .A(n5960), .ZN(n5966) );
  INV_X1 U7063 ( .A(n5962), .ZN(n5964) );
  OAI21_X1 U7064 ( .B1(n5964), .B2(n5963), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5965) );
  NAND3_X1 U7065 ( .A1(n5967), .A2(n5966), .A3(n5965), .ZN(U3018) );
  OAI21_X1 U7066 ( .B1(n3868), .B2(STATEBS16_REG_SCAN_IN), .A(n6530), .ZN(
        n5970) );
  OAI22_X1 U7067 ( .A1(n5970), .A2(n6529), .B1(n5969), .B2(n5968), .ZN(n5971)
         );
  MUX2_X1 U7068 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5971), .S(n6404), 
        .Z(U3464) );
  OAI22_X1 U7069 ( .A1(n5973), .A2(n6727), .B1(n5972), .B2(n6629), .ZN(n5974)
         );
  MUX2_X1 U7070 ( .A(n5974), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6080), 
        .Z(U3456) );
  AND2_X1 U7071 ( .A1(n6262), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U7072 ( .A1(EBX_REG_26__SCAN_IN), .A2(n6198), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6197), .ZN(n5980) );
  AND2_X1 U7073 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5987), .ZN(n5982) );
  AOI21_X1 U7074 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5982), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5977) );
  OAI22_X1 U7075 ( .A1(n5977), .A2(n5976), .B1(n5975), .B2(n6193), .ZN(n5978)
         );
  AOI21_X1 U7076 ( .B1(n6029), .B2(n6167), .A(n5978), .ZN(n5979) );
  OAI211_X1 U7077 ( .C1(n5981), .C2(n6188), .A(n5980), .B(n5979), .ZN(U2801)
         );
  INV_X1 U7078 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6701) );
  AOI22_X1 U7079 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n6197), .B1(n5982), 
        .B2(n6701), .ZN(n5993) );
  AOI22_X1 U7080 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6198), .B1(n5983), .B2(n6207), .ZN(n5992) );
  OAI22_X1 U7081 ( .A1(n6032), .A2(n6177), .B1(n6193), .B2(n5984), .ZN(n5985)
         );
  INV_X1 U7082 ( .A(n5985), .ZN(n5991) );
  AND2_X1 U7083 ( .A1(n6132), .A2(n5986), .ZN(n6006) );
  INV_X1 U7084 ( .A(REIP_REG_24__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7085 ( .A1(n5988), .A2(n5987), .ZN(n5996) );
  INV_X1 U7086 ( .A(n5996), .ZN(n5989) );
  OAI21_X1 U7087 ( .B1(n6006), .B2(n5989), .A(REIP_REG_25__SCAN_IN), .ZN(n5990) );
  NAND4_X1 U7088 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(U2802)
         );
  AOI22_X1 U7089 ( .A1(EBX_REG_24__SCAN_IN), .A2(n6198), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6197), .ZN(n5999) );
  AOI22_X1 U7090 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6006), .B1(n5994), .B2(
        n6207), .ZN(n5998) );
  AOI22_X1 U7091 ( .A1(n6036), .A2(n6167), .B1(n6202), .B2(n5995), .ZN(n5997)
         );
  NAND4_X1 U7092 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), .ZN(U2803)
         );
  AOI22_X1 U7093 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6198), .B1(n6000), .B2(n6207), .ZN(n6008) );
  INV_X1 U7094 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6695) );
  INV_X1 U7095 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6698) );
  OAI21_X1 U7096 ( .B1(n6695), .B2(n6001), .A(n6698), .ZN(n6005) );
  OAI22_X1 U7097 ( .A1(n6003), .A2(n6177), .B1(n6002), .B2(n6193), .ZN(n6004)
         );
  AOI21_X1 U7098 ( .B1(n6006), .B2(n6005), .A(n6004), .ZN(n6007) );
  OAI211_X1 U7099 ( .C1(n6009), .C2(n6171), .A(n6008), .B(n6007), .ZN(U2804)
         );
  AOI22_X1 U7100 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6198), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6197), .ZN(n6017) );
  AOI22_X1 U7101 ( .A1(n6011), .A2(n6207), .B1(REIP_REG_21__SCAN_IN), .B2(
        n6010), .ZN(n6016) );
  OAI22_X1 U7102 ( .A1(n6042), .A2(n6177), .B1(n6012), .B2(n6193), .ZN(n6013)
         );
  INV_X1 U7103 ( .A(n6013), .ZN(n6015) );
  NAND4_X1 U7104 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(U2806)
         );
  NAND2_X1 U7105 ( .A1(n6132), .A2(n6018), .ZN(n6121) );
  NAND2_X1 U7106 ( .A1(n6019), .A2(n6690), .ZN(n6110) );
  INV_X1 U7107 ( .A(n6020), .ZN(n6021) );
  AOI22_X1 U7108 ( .A1(n6022), .A2(n6207), .B1(n6021), .B2(n6691), .ZN(n6023)
         );
  OAI211_X1 U7109 ( .C1(n6171), .C2(n6957), .A(n6023), .B(n6186), .ZN(n6027)
         );
  OAI22_X1 U7110 ( .A1(n6025), .A2(n6177), .B1(n6024), .B2(n6193), .ZN(n6026)
         );
  AOI211_X1 U7111 ( .C1(EBX_REG_19__SCAN_IN), .C2(n6198), .A(n6027), .B(n6026), 
        .ZN(n6028) );
  OAI221_X1 U7112 ( .B1(n6691), .B2(n6121), .C1(n6691), .C2(n6110), .A(n6028), 
        .ZN(U2808) );
  AOI22_X1 U7113 ( .A1(n6029), .A2(n6237), .B1(n6228), .B2(DATAI_26_), .ZN(
        n6031) );
  AOI22_X1 U7114 ( .A1(n6231), .A2(DATAI_10_), .B1(n6230), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6030) );
  NAND2_X1 U7115 ( .A1(n6031), .A2(n6030), .ZN(U2865) );
  INV_X1 U7116 ( .A(n6032), .ZN(n6033) );
  AOI22_X1 U7117 ( .A1(n6033), .A2(n6237), .B1(n6228), .B2(DATAI_25_), .ZN(
        n6035) );
  AOI22_X1 U7118 ( .A1(n6231), .A2(DATAI_9_), .B1(n6230), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7119 ( .A1(n6035), .A2(n6034), .ZN(U2866) );
  AOI22_X1 U7120 ( .A1(n6036), .A2(n6237), .B1(DATAI_24_), .B2(n6228), .ZN(
        n6038) );
  AOI22_X1 U7121 ( .A1(n6231), .A2(DATAI_8_), .B1(n6230), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7122 ( .A1(n6038), .A2(n6037), .ZN(U2867) );
  AOI22_X1 U7123 ( .A1(n6039), .A2(n6237), .B1(n6228), .B2(DATAI_22_), .ZN(
        n6041) );
  AOI22_X1 U7124 ( .A1(n6231), .A2(DATAI_6_), .B1(n6230), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7125 ( .A1(n6041), .A2(n6040), .ZN(U2869) );
  INV_X1 U7126 ( .A(n6042), .ZN(n6043) );
  AOI22_X1 U7127 ( .A1(n6043), .A2(n6237), .B1(n6228), .B2(DATAI_21_), .ZN(
        n6045) );
  AOI22_X1 U7128 ( .A1(n6231), .A2(DATAI_5_), .B1(n6230), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6044) );
  NAND2_X1 U7129 ( .A1(n6045), .A2(n6044), .ZN(U2870) );
  AOI22_X1 U7130 ( .A1(n6046), .A2(n6237), .B1(n6228), .B2(DATAI_20_), .ZN(
        n6048) );
  AOI22_X1 U7131 ( .A1(n6231), .A2(DATAI_4_), .B1(n6230), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6047) );
  NAND2_X1 U7132 ( .A1(n6048), .A2(n6047), .ZN(U2871) );
  AOI22_X1 U7133 ( .A1(n6353), .A2(REIP_REG_18__SCAN_IN), .B1(n6299), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6051) );
  AOI22_X1 U7134 ( .A1(n6049), .A2(n6303), .B1(n4244), .B2(n6222), .ZN(n6050)
         );
  OAI211_X1 U7135 ( .C1(n6308), .C2(n6111), .A(n6051), .B(n6050), .ZN(U2968)
         );
  AND3_X1 U7136 ( .A1(n5784), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6271), 
        .ZN(n6052) );
  NOR2_X1 U7137 ( .A1(n6053), .A2(n6052), .ZN(n6055) );
  XNOR2_X1 U7138 ( .A(n6055), .B(n6054), .ZN(n6071) );
  AOI22_X1 U7139 ( .A1(n6353), .A2(REIP_REG_17__SCAN_IN), .B1(n6299), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6058) );
  XOR2_X1 U7140 ( .A(n6056), .B(n3173), .Z(n6225) );
  AOI22_X1 U7141 ( .A1(n6225), .A2(n4244), .B1(n6118), .B2(n6276), .ZN(n6057)
         );
  OAI211_X1 U7142 ( .C1(n6071), .C2(n6294), .A(n6058), .B(n6057), .ZN(U2969)
         );
  INV_X1 U7143 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6064) );
  INV_X1 U7144 ( .A(n6148), .ZN(n6059) );
  AOI222_X1 U7145 ( .A1(n6060), .A2(n6303), .B1(n6059), .B2(n6276), .C1(n4244), 
        .C2(n6145), .ZN(n6062) );
  OAI211_X1 U7146 ( .C1(n6064), .C2(n6063), .A(n6062), .B(n6061), .ZN(U2973)
         );
  AOI22_X1 U7147 ( .A1(n6353), .A2(REIP_REG_17__SCAN_IN), .B1(n6065), .B2(
        n6311), .ZN(n6070) );
  AOI21_X1 U7148 ( .B1(n3216), .B2(n3193), .A(n6067), .ZN(n6212) );
  AOI22_X1 U7149 ( .A1(n6068), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n6383), .B2(n6212), .ZN(n6069) );
  OAI211_X1 U7150 ( .C1(n6071), .C2(n6370), .A(n6070), .B(n6069), .ZN(U3001)
         );
  NOR3_X1 U7151 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n6073), .A3(n6072), 
        .ZN(n6076) );
  OAI22_X1 U7152 ( .A1(n6074), .A2(n6370), .B1(n6390), .B2(n6130), .ZN(n6075)
         );
  AOI211_X1 U7153 ( .C1(REIP_REG_16__SCAN_IN), .C2(n6353), .A(n6076), .B(n6075), .ZN(n6077) );
  OAI21_X1 U7154 ( .B1(n6079), .B2(n6078), .A(n6077), .ZN(U3002) );
  INV_X1 U7155 ( .A(n6080), .ZN(n6725) );
  INV_X1 U7156 ( .A(n6081), .ZN(n6083) );
  NAND4_X1 U7157 ( .A1(n6084), .A2(n6083), .A3(n6082), .A4(n6183), .ZN(n6085)
         );
  OAI21_X1 U7158 ( .B1(n6725), .B2(n4575), .A(n6085), .ZN(U3455) );
  INV_X1 U7159 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6664) );
  AOI21_X1 U7160 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6664), .A(n4316), .ZN(n6088) );
  INV_X1 U7161 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6086) );
  AND2_X1 U7162 ( .A1(STATE_REG_1__SCAN_IN), .A2(n4316), .ZN(n6712) );
  AOI21_X1 U7163 ( .B1(n6088), .B2(n6086), .A(n6712), .ZN(U2789) );
  INV_X2 U7164 ( .A(n6712), .ZN(n7148) );
  NOR2_X1 U7165 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6089) );
  OAI21_X1 U7166 ( .B1(n6089), .B2(D_C_N_REG_SCAN_IN), .A(n7148), .ZN(n6087)
         );
  OAI21_X1 U7167 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n7148), .A(n6087), .ZN(
        U2791) );
  NOR2_X1 U7168 ( .A1(n6712), .A2(n6088), .ZN(n6716) );
  OAI21_X1 U7169 ( .B1(BS16_N), .B2(n6089), .A(n6716), .ZN(n6714) );
  OAI21_X1 U7170 ( .B1(n6716), .B2(n6738), .A(n6714), .ZN(U2792) );
  OAI21_X1 U7171 ( .B1(n6091), .B2(n6090), .A(n6294), .ZN(U2793) );
  NOR4_X1 U7172 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6095) );
  NOR4_X1 U7173 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6094) );
  NOR4_X1 U7174 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6093) );
  NOR4_X1 U7175 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_22__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6092) );
  NAND4_X1 U7176 ( .A1(n6095), .A2(n6094), .A3(n6093), .A4(n6092), .ZN(n6101)
         );
  NOR4_X1 U7177 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(DATAWIDTH_REG_23__SCAN_IN), .ZN(
        n6099) );
  AOI211_X1 U7178 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_5__SCAN_IN), .B(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6098) );
  NOR4_X1 U7179 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n6097) );
  NOR4_X1 U7180 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6096) );
  NAND4_X1 U7181 ( .A1(n6099), .A2(n6098), .A3(n6097), .A4(n6096), .ZN(n6100)
         );
  NOR2_X1 U7182 ( .A1(n6101), .A2(n6100), .ZN(n6735) );
  INV_X1 U7183 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7039) );
  NOR3_X1 U7184 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6103) );
  OAI21_X1 U7185 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6103), .A(n6735), .ZN(n6102)
         );
  OAI21_X1 U7186 ( .B1(n6735), .B2(n7039), .A(n6102), .ZN(U2794) );
  INV_X1 U7187 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6715) );
  AOI21_X1 U7188 ( .B1(n6104), .B2(n6715), .A(n6103), .ZN(n6106) );
  INV_X1 U7189 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6105) );
  INV_X1 U7190 ( .A(n6735), .ZN(n6732) );
  AOI22_X1 U7191 ( .A1(n6735), .A2(n6106), .B1(n6105), .B2(n6732), .ZN(U2795)
         );
  AOI22_X1 U7192 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6198), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6197), .ZN(n6107) );
  OAI211_X1 U7193 ( .C1(n6121), .C2(n6690), .A(n6107), .B(n6186), .ZN(n6108)
         );
  INV_X1 U7194 ( .A(n6108), .ZN(n6109) );
  OAI211_X1 U7195 ( .C1(n6188), .C2(n6111), .A(n6110), .B(n6109), .ZN(n6112)
         );
  AOI21_X1 U7196 ( .B1(n6222), .B2(n6167), .A(n6112), .ZN(n6113) );
  OAI21_X1 U7197 ( .B1(n6193), .B2(n6114), .A(n6113), .ZN(U2809) );
  INV_X1 U7198 ( .A(n6125), .ZN(n6115) );
  AOI21_X1 U7199 ( .B1(n6115), .B2(REIP_REG_16__SCAN_IN), .A(
        REIP_REG_17__SCAN_IN), .ZN(n6122) );
  OAI22_X1 U7200 ( .A1(n6214), .A2(n6172), .B1(n6116), .B2(n6171), .ZN(n6117)
         );
  AOI211_X1 U7201 ( .C1(n6207), .C2(n6118), .A(n6175), .B(n6117), .ZN(n6120)
         );
  AOI22_X1 U7202 ( .A1(n6225), .A2(n6167), .B1(n6202), .B2(n6212), .ZN(n6119)
         );
  OAI211_X1 U7203 ( .C1(n6122), .C2(n6121), .A(n6120), .B(n6119), .ZN(U2810)
         );
  AOI22_X1 U7204 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6198), .B1(
        REIP_REG_16__SCAN_IN), .B2(n6123), .ZN(n6124) );
  OAI21_X1 U7205 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6125), .A(n6124), .ZN(n6126) );
  AOI211_X1 U7206 ( .C1(n6197), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6175), 
        .B(n6126), .ZN(n6129) );
  AOI22_X1 U7207 ( .A1(n6229), .A2(n6167), .B1(n6207), .B2(n6127), .ZN(n6128)
         );
  OAI211_X1 U7208 ( .C1(n6193), .C2(n6130), .A(n6129), .B(n6128), .ZN(U2811)
         );
  AOI22_X1 U7209 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6198), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6197), .ZN(n6138) );
  AOI21_X1 U7210 ( .B1(n6215), .B2(n6202), .A(n6175), .ZN(n6137) );
  AOI22_X1 U7211 ( .A1(n6234), .A2(n6167), .B1(n6207), .B2(n6131), .ZN(n6136)
         );
  INV_X1 U7212 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6682) );
  NOR3_X1 U7213 ( .A1(n6139), .A2(n6902), .A3(n6682), .ZN(n6134) );
  OAI211_X1 U7214 ( .C1(REIP_REG_14__SCAN_IN), .C2(n6134), .A(n6133), .B(n6132), .ZN(n6135) );
  NAND4_X1 U7215 ( .A1(n6138), .A2(n6137), .A3(n6136), .A4(n6135), .ZN(U2813)
         );
  NOR2_X1 U7217 ( .A1(n6139), .A2(n6902), .ZN(n6140) );
  NOR2_X1 U7218 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6139), .ZN(n6151) );
  OAI33_X1 U7219 ( .A1(1'b0), .A2(n6140), .A3(REIP_REG_13__SCAN_IN), .B1(n6682), .B2(n6149), .B3(n6151), .ZN(n6147) );
  AOI22_X1 U7220 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6198), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n6197), .ZN(n6142) );
  OAI211_X1 U7221 ( .C1(n6193), .C2(n6143), .A(n6142), .B(n6186), .ZN(n6144)
         );
  AOI21_X1 U7222 ( .B1(n6145), .B2(n6167), .A(n6144), .ZN(n6146) );
  OAI211_X1 U7223 ( .C1(n6148), .C2(n6188), .A(n6147), .B(n6146), .ZN(U2814)
         );
  AOI22_X1 U7224 ( .A1(n6202), .A2(n6150), .B1(REIP_REG_12__SCAN_IN), .B2(
        n6149), .ZN(n6157) );
  AOI211_X1 U7225 ( .C1(n6197), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6175), 
        .B(n6151), .ZN(n6156) );
  INV_X1 U7226 ( .A(n6152), .ZN(n6153) );
  AOI22_X1 U7227 ( .A1(n6238), .A2(n6167), .B1(n6153), .B2(n6207), .ZN(n6155)
         );
  NAND2_X1 U7228 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6198), .ZN(n6154) );
  NAND4_X1 U7229 ( .A1(n6157), .A2(n6156), .A3(n6155), .A4(n6154), .ZN(U2815)
         );
  NAND2_X1 U7230 ( .A1(n6159), .A2(n6158), .ZN(n6160) );
  AND2_X1 U7231 ( .A1(n6161), .A2(n6160), .ZN(n6328) );
  AOI22_X1 U7232 ( .A1(n6202), .A2(n6328), .B1(REIP_REG_9__SCAN_IN), .B2(n6162), .ZN(n6170) );
  OAI22_X1 U7233 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6163), .B1(n4942), .B2(n6171), .ZN(n6164) );
  AOI211_X1 U7234 ( .C1(n6198), .C2(EBX_REG_9__SCAN_IN), .A(n6175), .B(n6164), 
        .ZN(n6169) );
  INV_X1 U7235 ( .A(n6165), .ZN(n6219) );
  AOI22_X1 U7236 ( .A1(n6219), .A2(n6167), .B1(n6207), .B2(n6166), .ZN(n6168)
         );
  NAND3_X1 U7237 ( .A1(n6170), .A2(n6169), .A3(n6168), .ZN(U2818) );
  OAI22_X1 U7238 ( .A1(n6173), .A2(n6172), .B1(n3914), .B2(n6171), .ZN(n6174)
         );
  AOI211_X1 U7239 ( .C1(REIP_REG_6__SCAN_IN), .C2(n6176), .A(n6175), .B(n6174), 
        .ZN(n6182) );
  NOR2_X1 U7240 ( .A1(n6178), .A2(n6177), .ZN(n6180) );
  AOI211_X1 U7241 ( .C1(n6352), .C2(n6202), .A(n6180), .B(n6179), .ZN(n6181)
         );
  OAI211_X1 U7242 ( .C1(n6287), .C2(n6188), .A(n6182), .B(n6181), .ZN(U2821)
         );
  AOI22_X1 U7243 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6198), .B1(n6183), .B2(n6196), 
        .ZN(n6192) );
  OR2_X1 U7244 ( .A1(n6185), .A2(n6184), .ZN(n6211) );
  OAI221_X1 U7245 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6187), .C1(n6669), .C2(
        n6211), .A(n6186), .ZN(n6190) );
  OAI22_X1 U7246 ( .A1(n6293), .A2(n6205), .B1(n6298), .B2(n6188), .ZN(n6189)
         );
  AOI211_X1 U7247 ( .C1(PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n6197), .A(n6190), 
        .B(n6189), .ZN(n6191) );
  OAI211_X1 U7248 ( .C1(n6193), .C2(n6372), .A(n6192), .B(n6191), .ZN(U2823)
         );
  OR2_X1 U7249 ( .A1(n6195), .A2(n6194), .ZN(n6210) );
  INV_X1 U7250 ( .A(n6196), .ZN(n6200) );
  AOI22_X1 U7251 ( .A1(n6198), .A2(EBX_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6197), .ZN(n6199) );
  OAI21_X1 U7252 ( .B1(n6200), .B2(n6407), .A(n6199), .ZN(n6201) );
  AOI21_X1 U7253 ( .B1(n6202), .B2(n6382), .A(n6201), .ZN(n6203) );
  OAI21_X1 U7254 ( .B1(n6205), .B2(n6204), .A(n6203), .ZN(n6206) );
  AOI21_X1 U7255 ( .B1(n6208), .B2(n6207), .A(n6206), .ZN(n6209) );
  OAI221_X1 U7256 ( .B1(n6211), .B2(n6667), .C1(n6211), .C2(n6210), .A(n6209), 
        .ZN(U2824) );
  AOI22_X1 U7257 ( .A1(n6225), .A2(n6218), .B1(n6217), .B2(n6212), .ZN(n6213)
         );
  OAI21_X1 U7258 ( .B1(n6214), .B2(n6221), .A(n6213), .ZN(U2842) );
  INV_X1 U7259 ( .A(EBX_REG_14__SCAN_IN), .ZN(n7030) );
  AOI22_X1 U7260 ( .A1(n6234), .A2(n6218), .B1(n6217), .B2(n6215), .ZN(n6216)
         );
  OAI21_X1 U7261 ( .B1(n7030), .B2(n6221), .A(n6216), .ZN(U2845) );
  AOI22_X1 U7262 ( .A1(n6219), .A2(n6218), .B1(n6217), .B2(n6328), .ZN(n6220)
         );
  OAI21_X1 U7263 ( .B1(n6883), .B2(n6221), .A(n6220), .ZN(U2850) );
  AOI22_X1 U7264 ( .A1(n6222), .A2(n6237), .B1(n6228), .B2(DATAI_18_), .ZN(
        n6224) );
  AOI22_X1 U7265 ( .A1(n6231), .A2(DATAI_2_), .B1(n6230), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7266 ( .A1(n6224), .A2(n6223), .ZN(U2873) );
  AOI22_X1 U7267 ( .A1(n6225), .A2(n6237), .B1(n6228), .B2(DATAI_17_), .ZN(
        n6227) );
  AOI22_X1 U7268 ( .A1(n6231), .A2(DATAI_1_), .B1(n6230), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7269 ( .A1(n6227), .A2(n6226), .ZN(U2874) );
  AOI22_X1 U7270 ( .A1(n6229), .A2(n6237), .B1(n6228), .B2(DATAI_16_), .ZN(
        n6233) );
  AOI22_X1 U7271 ( .A1(n6231), .A2(DATAI_0_), .B1(n6230), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7272 ( .A1(n6233), .A2(n6232), .ZN(U2875) );
  AOI22_X1 U7273 ( .A1(n6234), .A2(n6237), .B1(DATAI_14_), .B2(n6236), .ZN(
        n6235) );
  OAI21_X1 U7274 ( .B1(n7058), .B2(n6240), .A(n6235), .ZN(U2877) );
  AOI22_X1 U7275 ( .A1(n6238), .A2(n6237), .B1(DATAI_12_), .B2(n6236), .ZN(
        n6239) );
  OAI21_X1 U7276 ( .B1(n6841), .B2(n6240), .A(n6239), .ZN(U2879) );
  INV_X1 U7277 ( .A(n6241), .ZN(n6268) );
  AOI22_X1 U7278 ( .A1(n6747), .A2(LWORD_REG_15__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6242) );
  OAI21_X1 U7279 ( .B1(n6243), .B2(n6268), .A(n6242), .ZN(U2908) );
  AOI22_X1 U7280 ( .A1(n6747), .A2(LWORD_REG_14__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6244) );
  OAI21_X1 U7281 ( .B1(n7058), .B2(n6268), .A(n6244), .ZN(U2909) );
  AOI22_X1 U7282 ( .A1(n6747), .A2(LWORD_REG_13__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6245) );
  OAI21_X1 U7283 ( .B1(n6860), .B2(n6268), .A(n6245), .ZN(U2910) );
  AOI22_X1 U7284 ( .A1(n6747), .A2(LWORD_REG_12__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6246) );
  OAI21_X1 U7285 ( .B1(n6841), .B2(n6268), .A(n6246), .ZN(U2911) );
  AOI22_X1 U7286 ( .A1(n6747), .A2(LWORD_REG_11__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6247) );
  OAI21_X1 U7287 ( .B1(n6248), .B2(n6268), .A(n6247), .ZN(U2912) );
  AOI22_X1 U7288 ( .A1(n6747), .A2(LWORD_REG_10__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6249) );
  OAI21_X1 U7289 ( .B1(n6859), .B2(n6268), .A(n6249), .ZN(U2913) );
  AOI22_X1 U7290 ( .A1(n6747), .A2(LWORD_REG_9__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6250) );
  OAI21_X1 U7291 ( .B1(n6251), .B2(n6268), .A(n6250), .ZN(U2914) );
  AOI22_X1 U7292 ( .A1(n6747), .A2(LWORD_REG_8__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6252) );
  OAI21_X1 U7293 ( .B1(n6253), .B2(n6268), .A(n6252), .ZN(U2915) );
  AOI22_X1 U7294 ( .A1(n6747), .A2(LWORD_REG_7__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6254) );
  OAI21_X1 U7295 ( .B1(n3928), .B2(n6268), .A(n6254), .ZN(U2916) );
  AOI22_X1 U7296 ( .A1(n6747), .A2(LWORD_REG_6__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6255) );
  OAI21_X1 U7297 ( .B1(n6256), .B2(n6268), .A(n6255), .ZN(U2917) );
  AOI22_X1 U7298 ( .A1(n6747), .A2(LWORD_REG_5__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6257) );
  OAI21_X1 U7299 ( .B1(n6258), .B2(n6268), .A(n6257), .ZN(U2918) );
  AOI22_X1 U7300 ( .A1(n6747), .A2(LWORD_REG_4__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7301 ( .B1(n6260), .B2(n6268), .A(n6259), .ZN(U2919) );
  AOI22_X1 U7302 ( .A1(n6747), .A2(LWORD_REG_3__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6261) );
  OAI21_X1 U7303 ( .B1(n6827), .B2(n6268), .A(n6261), .ZN(U2920) );
  AOI22_X1 U7304 ( .A1(n6747), .A2(LWORD_REG_2__SCAN_IN), .B1(n6262), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6263) );
  OAI21_X1 U7305 ( .B1(n6973), .B2(n6268), .A(n6263), .ZN(U2921) );
  AOI22_X1 U7306 ( .A1(n6747), .A2(LWORD_REG_1__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6264) );
  OAI21_X1 U7307 ( .B1(n6265), .B2(n6268), .A(n6264), .ZN(U2922) );
  AOI22_X1 U7308 ( .A1(n6747), .A2(LWORD_REG_0__SCAN_IN), .B1(n6266), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6267) );
  OAI21_X1 U7309 ( .B1(n6988), .B2(n6268), .A(n6267), .ZN(U2923) );
  NAND2_X1 U7310 ( .A1(n6270), .A2(n6269), .ZN(n6273) );
  XNOR2_X1 U7311 ( .A(n6271), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6272)
         );
  XNOR2_X1 U7312 ( .A(n6273), .B(n6272), .ZN(n6315) );
  AOI22_X1 U7313 ( .A1(n6353), .A2(REIP_REG_11__SCAN_IN), .B1(n6299), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6279) );
  INV_X1 U7314 ( .A(n6274), .ZN(n6277) );
  AOI22_X1 U7315 ( .A1(n6277), .A2(n4244), .B1(n6276), .B2(n6275), .ZN(n6278)
         );
  OAI211_X1 U7316 ( .C1(n6315), .C2(n6294), .A(n6279), .B(n6278), .ZN(U2975)
         );
  AOI22_X1 U7317 ( .A1(n6353), .A2(REIP_REG_6__SCAN_IN), .B1(n6299), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6286) );
  OAI21_X1 U7318 ( .B1(n6282), .B2(n6281), .A(n6280), .ZN(n6283) );
  INV_X1 U7319 ( .A(n6283), .ZN(n6351) );
  AOI22_X1 U7320 ( .A1(n6351), .A2(n6303), .B1(n4244), .B2(n6284), .ZN(n6285)
         );
  OAI211_X1 U7321 ( .C1(n6308), .C2(n6287), .A(n6286), .B(n6285), .ZN(U2980)
         );
  AOI22_X1 U7322 ( .A1(n6353), .A2(REIP_REG_4__SCAN_IN), .B1(n6299), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6297) );
  OR2_X1 U7323 ( .A1(n6289), .A2(n6288), .ZN(n6290) );
  NAND2_X1 U7324 ( .A1(n6291), .A2(n6290), .ZN(n6371) );
  OAI22_X1 U7325 ( .A1(n6371), .A2(n6294), .B1(n6293), .B2(n6292), .ZN(n6295)
         );
  INV_X1 U7326 ( .A(n6295), .ZN(n6296) );
  OAI211_X1 U7327 ( .C1(n6308), .C2(n6298), .A(n6297), .B(n6296), .ZN(U2982)
         );
  AOI22_X1 U7328 ( .A1(n6353), .A2(REIP_REG_2__SCAN_IN), .B1(n6299), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6306) );
  XNOR2_X1 U7329 ( .A(n6300), .B(n6398), .ZN(n6301) );
  XNOR2_X1 U7330 ( .A(n6302), .B(n6301), .ZN(n6395) );
  AOI22_X1 U7331 ( .A1(n6304), .A2(n4244), .B1(n6303), .B2(n6395), .ZN(n6305)
         );
  OAI211_X1 U7332 ( .C1(n6308), .C2(n6307), .A(n6306), .B(n6305), .ZN(U2984)
         );
  INV_X1 U7333 ( .A(n6309), .ZN(n6310) );
  AOI22_X1 U7334 ( .A1(n6383), .A2(n6310), .B1(n6353), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6314) );
  AOI22_X1 U7335 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6312), .B1(n6311), .B2(n3700), .ZN(n6313) );
  OAI211_X1 U7336 ( .C1(n6315), .C2(n6370), .A(n6314), .B(n6313), .ZN(U3007)
         );
  NAND2_X1 U7337 ( .A1(n6320), .A2(n6338), .ZN(n6333) );
  AOI22_X1 U7338 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n3699), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6316), .ZN(n6325) );
  INV_X1 U7339 ( .A(n6317), .ZN(n6319) );
  AOI21_X1 U7340 ( .B1(n6383), .B2(n6319), .A(n6318), .ZN(n6324) );
  OAI21_X1 U7341 ( .B1(n6321), .B2(n6320), .A(n6343), .ZN(n6329) );
  AOI22_X1 U7342 ( .A1(n6322), .A2(n6396), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6329), .ZN(n6323) );
  OAI211_X1 U7343 ( .C1(n6333), .C2(n6325), .A(n6324), .B(n6323), .ZN(U3008)
         );
  INV_X1 U7344 ( .A(n6326), .ZN(n6327) );
  AOI21_X1 U7345 ( .B1(n6383), .B2(n6328), .A(n6327), .ZN(n6332) );
  AOI22_X1 U7346 ( .A1(n6330), .A2(n6396), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6329), .ZN(n6331) );
  OAI211_X1 U7347 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6333), .A(n6332), 
        .B(n6331), .ZN(U3009) );
  INV_X1 U7348 ( .A(n6334), .ZN(n6335) );
  AOI21_X1 U7349 ( .B1(n6383), .B2(n6336), .A(n6335), .ZN(n6341) );
  INV_X1 U7350 ( .A(n6337), .ZN(n6339) );
  AOI22_X1 U7351 ( .A1(n6339), .A2(n6396), .B1(n6338), .B2(n6342), .ZN(n6340)
         );
  OAI211_X1 U7352 ( .C1(n6343), .C2(n6342), .A(n6341), .B(n6340), .ZN(U3011)
         );
  NAND3_X1 U7353 ( .A1(n6344), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6369), 
        .ZN(n6349) );
  INV_X1 U7354 ( .A(n6349), .ZN(n6346) );
  NAND2_X1 U7355 ( .A1(n6346), .A2(n6345), .ZN(n6356) );
  OAI22_X1 U7356 ( .A1(n6348), .A2(n6393), .B1(n6392), .B2(n6347), .ZN(n6397)
         );
  AOI21_X1 U7357 ( .B1(n6350), .B2(n6349), .A(n6397), .ZN(n6368) );
  AOI222_X1 U7358 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6353), .B1(n6383), .B2(
        n6352), .C1(n6396), .C2(n6351), .ZN(n6354) );
  OAI221_X1 U7359 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6356), .C1(n6355), .C2(n6368), .A(n6354), .ZN(U3012) );
  INV_X1 U7360 ( .A(n6369), .ZN(n6362) );
  NOR2_X1 U7361 ( .A1(n6394), .A2(n6362), .ZN(n6357) );
  AOI21_X1 U7362 ( .B1(n6392), .B2(n6357), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6367) );
  INV_X1 U7363 ( .A(n6358), .ZN(n6360) );
  AOI21_X1 U7364 ( .B1(n6383), .B2(n6360), .A(n6359), .ZN(n6366) );
  NOR3_X1 U7365 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6362), .A3(n6361), 
        .ZN(n6363) );
  AOI21_X1 U7366 ( .B1(n6396), .B2(n6364), .A(n6363), .ZN(n6365) );
  OAI211_X1 U7367 ( .C1(n6368), .C2(n6367), .A(n6366), .B(n6365), .ZN(U3013)
         );
  AOI21_X1 U7368 ( .B1(n6392), .B2(n6394), .A(n6397), .ZN(n6385) );
  AOI211_X1 U7369 ( .C1(n6386), .C2(n6377), .A(n6369), .B(n6387), .ZN(n6375)
         );
  NOR2_X1 U7370 ( .A1(n6371), .A2(n6370), .ZN(n6374) );
  OAI22_X1 U7371 ( .A1(n6390), .A2(n6372), .B1(n6669), .B2(n6388), .ZN(n6373)
         );
  NOR3_X1 U7372 ( .A1(n6375), .A2(n6374), .A3(n6373), .ZN(n6376) );
  OAI21_X1 U7373 ( .B1(n6385), .B2(n6377), .A(n6376), .ZN(U3014) );
  INV_X1 U7374 ( .A(n6378), .ZN(n6381) );
  AND3_X1 U7375 ( .A1(n4466), .A2(n6379), .A3(n6396), .ZN(n6380) );
  AOI211_X1 U7376 ( .C1(n6383), .C2(n6382), .A(n6381), .B(n6380), .ZN(n6384)
         );
  OAI221_X1 U7377 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6387), .C1(n6386), .C2(n6385), .A(n6384), .ZN(U3015) );
  OAI22_X1 U7378 ( .A1(n6390), .A2(n6389), .B1(n6194), .B2(n6388), .ZN(n6391)
         );
  INV_X1 U7379 ( .A(n6391), .ZN(n6403) );
  OAI221_X1 U7380 ( .B1(n6394), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .C1(n6394), .C2(n6393), .A(n6392), .ZN(n6402) );
  AOI22_X1 U7381 ( .A1(n6397), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6396), 
        .B2(n6395), .ZN(n6401) );
  NAND3_X1 U7382 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6399), .A3(n6398), 
        .ZN(n6400) );
  NAND4_X1 U7383 ( .A1(n6403), .A2(n6402), .A3(n6401), .A4(n6400), .ZN(U3016)
         );
  NOR2_X1 U7384 ( .A1(n6611), .A2(n6404), .ZN(U3019) );
  AND2_X1 U7385 ( .A1(n4585), .A2(n6405), .ZN(n6406) );
  NAND3_X1 U7386 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6435), .A3(n6607), .ZN(n6445) );
  NOR2_X1 U7387 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6445), .ZN(n6430)
         );
  NAND2_X1 U7388 ( .A1(n6407), .A2(n3262), .ZN(n6440) );
  OAI22_X1 U7389 ( .A1(n6440), .A2(n6535), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6408), .ZN(n6429) );
  AOI22_X1 U7390 ( .A1(n6526), .A2(n6430), .B1(n6541), .B2(n6429), .ZN(n6414)
         );
  INV_X1 U7391 ( .A(n6474), .ZN(n6456) );
  OAI21_X1 U7392 ( .B1(n6431), .B2(n6456), .A(n6409), .ZN(n6410) );
  AOI21_X1 U7393 ( .B1(n6410), .B2(n6440), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6412) );
  OAI21_X1 U7394 ( .B1(n6430), .B2(n6412), .A(n6411), .ZN(n6432) );
  AOI22_X1 U7395 ( .A1(n6432), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n6527), 
        .B2(n6431), .ZN(n6413) );
  OAI211_X1 U7396 ( .C1(n6544), .C2(n6474), .A(n6414), .B(n6413), .ZN(U3036)
         );
  AOI22_X1 U7397 ( .A1(n6545), .A2(n6430), .B1(n6547), .B2(n6429), .ZN(n6417)
         );
  AOI22_X1 U7398 ( .A1(n6432), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n6415), 
        .B2(n6431), .ZN(n6416) );
  OAI211_X1 U7399 ( .C1(n6474), .C2(n6418), .A(n6417), .B(n6416), .ZN(U3037)
         );
  AOI22_X1 U7400 ( .A1(n6551), .A2(n6430), .B1(n6553), .B2(n6429), .ZN(n6420)
         );
  AOI22_X1 U7401 ( .A1(n6432), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n6552), 
        .B2(n6431), .ZN(n6419) );
  OAI211_X1 U7402 ( .C1(n6474), .C2(n6556), .A(n6420), .B(n6419), .ZN(U3038)
         );
  AOI22_X1 U7403 ( .A1(n6557), .A2(n6430), .B1(n6559), .B2(n6429), .ZN(n6422)
         );
  AOI22_X1 U7404 ( .A1(n6432), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n6558), 
        .B2(n6431), .ZN(n6421) );
  OAI211_X1 U7405 ( .C1(n6474), .C2(n6562), .A(n6422), .B(n6421), .ZN(U3039)
         );
  AOI22_X1 U7406 ( .A1(n6563), .A2(n6430), .B1(n6565), .B2(n6429), .ZN(n6424)
         );
  AOI22_X1 U7407 ( .A1(n6432), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n6564), 
        .B2(n6431), .ZN(n6423) );
  OAI211_X1 U7408 ( .C1(n6474), .C2(n6568), .A(n6424), .B(n6423), .ZN(U3040)
         );
  AOI22_X1 U7409 ( .A1(n6569), .A2(n6430), .B1(n6571), .B2(n6429), .ZN(n6426)
         );
  AOI22_X1 U7410 ( .A1(n6432), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n6570), 
        .B2(n6431), .ZN(n6425) );
  OAI211_X1 U7411 ( .C1(n6474), .C2(n6574), .A(n6426), .B(n6425), .ZN(U3041)
         );
  AOI22_X1 U7412 ( .A1(n6575), .A2(n6430), .B1(n6578), .B2(n6429), .ZN(n6428)
         );
  AOI22_X1 U7413 ( .A1(n6432), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n6510), 
        .B2(n6431), .ZN(n6427) );
  OAI211_X1 U7414 ( .C1(n6474), .C2(n6515), .A(n6428), .B(n6427), .ZN(U3042)
         );
  AOI22_X1 U7415 ( .A1(n6584), .A2(n6430), .B1(n6588), .B2(n6429), .ZN(n6434)
         );
  AOI22_X1 U7416 ( .A1(n6432), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n6585), 
        .B2(n6431), .ZN(n6433) );
  OAI211_X1 U7417 ( .C1(n6474), .C2(n6593), .A(n6434), .B(n6433), .ZN(U3043)
         );
  INV_X1 U7418 ( .A(n6525), .ZN(n6436) );
  NAND2_X1 U7419 ( .A1(n6436), .A2(n6435), .ZN(n6441) );
  INV_X1 U7420 ( .A(n6441), .ZN(n6469) );
  AOI22_X1 U7421 ( .A1(n6526), .A2(n6469), .B1(n6482), .B2(n6468), .ZN(n6449)
         );
  NAND3_X1 U7422 ( .A1(n6437), .A2(n6529), .A3(n4585), .ZN(n6438) );
  NAND2_X1 U7423 ( .A1(n6438), .A2(n6530), .ZN(n6447) );
  INV_X1 U7424 ( .A(n6597), .ZN(n6439) );
  OR2_X1 U7425 ( .A1(n6440), .A2(n6439), .ZN(n6442) );
  NAND2_X1 U7426 ( .A1(n6442), .A2(n6441), .ZN(n6444) );
  AOI21_X1 U7427 ( .B1(n6535), .B2(n6445), .A(n6534), .ZN(n6443) );
  OAI21_X1 U7428 ( .B1(n6447), .B2(n6444), .A(n6443), .ZN(n6471) );
  INV_X1 U7429 ( .A(n6444), .ZN(n6446) );
  OAI22_X1 U7430 ( .A1(n6447), .A2(n6446), .B1(n6445), .B2(n6737), .ZN(n6470)
         );
  AOI22_X1 U7431 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6471), .B1(n6541), 
        .B2(n6470), .ZN(n6448) );
  OAI211_X1 U7432 ( .C1(n6495), .C2(n6474), .A(n6449), .B(n6448), .ZN(U3044)
         );
  AOI22_X1 U7433 ( .A1(n6545), .A2(n6469), .B1(n6546), .B2(n6468), .ZN(n6451)
         );
  AOI22_X1 U7434 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6471), .B1(n6547), 
        .B2(n6470), .ZN(n6450) );
  OAI211_X1 U7435 ( .C1(n6474), .C2(n6550), .A(n6451), .B(n6450), .ZN(U3045)
         );
  AOI22_X1 U7436 ( .A1(n6551), .A2(n6469), .B1(n6452), .B2(n6468), .ZN(n6454)
         );
  AOI22_X1 U7437 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6471), .B1(n6553), 
        .B2(n6470), .ZN(n6453) );
  OAI211_X1 U7438 ( .C1(n6474), .C2(n6455), .A(n6454), .B(n6453), .ZN(U3046)
         );
  AOI22_X1 U7439 ( .A1(n6557), .A2(n6469), .B1(n6558), .B2(n6456), .ZN(n6458)
         );
  AOI22_X1 U7440 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6471), .B1(n6559), 
        .B2(n6470), .ZN(n6457) );
  OAI211_X1 U7441 ( .C1(n6562), .C2(n6459), .A(n6458), .B(n6457), .ZN(U3047)
         );
  AOI22_X1 U7442 ( .A1(n6563), .A2(n6469), .B1(n6460), .B2(n6468), .ZN(n6462)
         );
  AOI22_X1 U7443 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6471), .B1(n6565), 
        .B2(n6470), .ZN(n6461) );
  OAI211_X1 U7444 ( .C1(n6474), .C2(n6463), .A(n6462), .B(n6461), .ZN(U3048)
         );
  AOI22_X1 U7445 ( .A1(n6569), .A2(n6469), .B1(n6506), .B2(n6468), .ZN(n6465)
         );
  AOI22_X1 U7446 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6471), .B1(n6571), 
        .B2(n6470), .ZN(n6464) );
  OAI211_X1 U7447 ( .C1(n6474), .C2(n6509), .A(n6465), .B(n6464), .ZN(U3049)
         );
  AOI22_X1 U7448 ( .A1(n6575), .A2(n6469), .B1(n6576), .B2(n6468), .ZN(n6467)
         );
  AOI22_X1 U7449 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6471), .B1(n6578), 
        .B2(n6470), .ZN(n6466) );
  OAI211_X1 U7450 ( .C1(n6474), .C2(n6582), .A(n6467), .B(n6466), .ZN(U3050)
         );
  AOI22_X1 U7451 ( .A1(n6584), .A2(n6469), .B1(n6516), .B2(n6468), .ZN(n6473)
         );
  AOI22_X1 U7452 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6471), .B1(n6588), 
        .B2(n6470), .ZN(n6472) );
  OAI211_X1 U7453 ( .C1(n6474), .C2(n6524), .A(n6473), .B(n6472), .ZN(U3051)
         );
  AOI22_X1 U7454 ( .A1(n6526), .A2(n6476), .B1(n6541), .B2(n6475), .ZN(n6480)
         );
  AOI22_X1 U7455 ( .A1(n6478), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6527), 
        .B2(n6477), .ZN(n6479) );
  OAI211_X1 U7456 ( .C1(n6544), .C2(n6523), .A(n6480), .B(n6479), .ZN(U3068)
         );
  INV_X1 U7457 ( .A(n6481), .ZN(n6518) );
  AOI22_X1 U7458 ( .A1(n6526), .A2(n6518), .B1(n6517), .B2(n6482), .ZN(n6494)
         );
  INV_X1 U7459 ( .A(n6483), .ZN(n6484) );
  AOI21_X1 U7460 ( .B1(n6485), .B2(n6484), .A(n6518), .ZN(n6492) );
  NAND3_X1 U7461 ( .A1(n6486), .A2(n6492), .A3(n6489), .ZN(n6487) );
  OAI211_X1 U7462 ( .C1(n3578), .C2(n6530), .A(n6488), .B(n6487), .ZN(n6520)
         );
  NAND2_X1 U7463 ( .A1(n6530), .A2(n6489), .ZN(n6491) );
  OAI22_X1 U7464 ( .A1(n6492), .A2(n6491), .B1(n6737), .B2(n6490), .ZN(n6519)
         );
  AOI22_X1 U7465 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6520), .B1(n6541), 
        .B2(n6519), .ZN(n6493) );
  OAI211_X1 U7466 ( .C1(n6495), .C2(n6523), .A(n6494), .B(n6493), .ZN(U3076)
         );
  AOI22_X1 U7467 ( .A1(n6545), .A2(n6518), .B1(n6517), .B2(n6546), .ZN(n6497)
         );
  AOI22_X1 U7468 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6520), .B1(n6547), 
        .B2(n6519), .ZN(n6496) );
  OAI211_X1 U7469 ( .C1(n6550), .C2(n6523), .A(n6497), .B(n6496), .ZN(U3077)
         );
  AOI22_X1 U7470 ( .A1(n6551), .A2(n6518), .B1(n6511), .B2(n6552), .ZN(n6499)
         );
  AOI22_X1 U7471 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6520), .B1(n6553), 
        .B2(n6519), .ZN(n6498) );
  OAI211_X1 U7472 ( .C1(n6556), .C2(n6514), .A(n6499), .B(n6498), .ZN(U3078)
         );
  AOI22_X1 U7473 ( .A1(n6557), .A2(n6518), .B1(n6517), .B2(n6500), .ZN(n6502)
         );
  AOI22_X1 U7474 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6520), .B1(n6559), 
        .B2(n6519), .ZN(n6501) );
  OAI211_X1 U7475 ( .C1(n6503), .C2(n6523), .A(n6502), .B(n6501), .ZN(U3079)
         );
  AOI22_X1 U7476 ( .A1(n6563), .A2(n6518), .B1(n6511), .B2(n6564), .ZN(n6505)
         );
  AOI22_X1 U7477 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6520), .B1(n6565), 
        .B2(n6519), .ZN(n6504) );
  OAI211_X1 U7478 ( .C1(n6568), .C2(n6514), .A(n6505), .B(n6504), .ZN(U3080)
         );
  AOI22_X1 U7479 ( .A1(n6569), .A2(n6518), .B1(n6517), .B2(n6506), .ZN(n6508)
         );
  AOI22_X1 U7480 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6520), .B1(n6571), 
        .B2(n6519), .ZN(n6507) );
  OAI211_X1 U7481 ( .C1(n6509), .C2(n6523), .A(n6508), .B(n6507), .ZN(U3081)
         );
  AOI22_X1 U7482 ( .A1(n6575), .A2(n6518), .B1(n6511), .B2(n6510), .ZN(n6513)
         );
  AOI22_X1 U7483 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6520), .B1(n6578), 
        .B2(n6519), .ZN(n6512) );
  OAI211_X1 U7484 ( .C1(n6515), .C2(n6514), .A(n6513), .B(n6512), .ZN(U3082)
         );
  AOI22_X1 U7485 ( .A1(n6584), .A2(n6518), .B1(n6517), .B2(n6516), .ZN(n6522)
         );
  AOI22_X1 U7486 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6520), .B1(n6588), 
        .B2(n6519), .ZN(n6521) );
  OAI211_X1 U7487 ( .C1(n6524), .C2(n6523), .A(n6522), .B(n6521), .ZN(U3083)
         );
  NOR2_X1 U7488 ( .A1(n6525), .A2(n6435), .ZN(n6583) );
  AOI22_X1 U7489 ( .A1(n6586), .A2(n6527), .B1(n6526), .B2(n6583), .ZN(n6543)
         );
  INV_X1 U7490 ( .A(n6528), .ZN(n6532) );
  INV_X1 U7491 ( .A(n6529), .ZN(n6531) );
  OAI21_X1 U7492 ( .B1(n6532), .B2(n6531), .A(n6530), .ZN(n6540) );
  AOI21_X1 U7493 ( .B1(n6533), .B2(n6597), .A(n6583), .ZN(n6539) );
  INV_X1 U7494 ( .A(n6539), .ZN(n6537) );
  AOI21_X1 U7495 ( .B1(n6535), .B2(n6538), .A(n6534), .ZN(n6536) );
  OAI21_X1 U7496 ( .B1(n6540), .B2(n6537), .A(n6536), .ZN(n6589) );
  OAI22_X1 U7497 ( .A1(n6540), .A2(n6539), .B1(n6538), .B2(n6737), .ZN(n6587)
         );
  AOI22_X1 U7498 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6589), .B1(n6541), 
        .B2(n6587), .ZN(n6542) );
  OAI211_X1 U7499 ( .C1(n6544), .C2(n6592), .A(n6543), .B(n6542), .ZN(U3108)
         );
  INV_X1 U7500 ( .A(n6592), .ZN(n6577) );
  AOI22_X1 U7501 ( .A1(n6577), .A2(n6546), .B1(n6545), .B2(n6583), .ZN(n6549)
         );
  AOI22_X1 U7502 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6589), .B1(n6547), 
        .B2(n6587), .ZN(n6548) );
  OAI211_X1 U7503 ( .C1(n6550), .C2(n6581), .A(n6549), .B(n6548), .ZN(U3109)
         );
  AOI22_X1 U7504 ( .A1(n6586), .A2(n6552), .B1(n6551), .B2(n6583), .ZN(n6555)
         );
  AOI22_X1 U7505 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6589), .B1(n6553), 
        .B2(n6587), .ZN(n6554) );
  OAI211_X1 U7506 ( .C1(n6556), .C2(n6592), .A(n6555), .B(n6554), .ZN(U3110)
         );
  AOI22_X1 U7507 ( .A1(n6586), .A2(n6558), .B1(n6557), .B2(n6583), .ZN(n6561)
         );
  AOI22_X1 U7508 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6589), .B1(n6559), 
        .B2(n6587), .ZN(n6560) );
  OAI211_X1 U7509 ( .C1(n6562), .C2(n6592), .A(n6561), .B(n6560), .ZN(U3111)
         );
  AOI22_X1 U7510 ( .A1(n6586), .A2(n6564), .B1(n6563), .B2(n6583), .ZN(n6567)
         );
  AOI22_X1 U7511 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6589), .B1(n6565), 
        .B2(n6587), .ZN(n6566) );
  OAI211_X1 U7512 ( .C1(n6568), .C2(n6592), .A(n6567), .B(n6566), .ZN(U3112)
         );
  AOI22_X1 U7513 ( .A1(n6586), .A2(n6570), .B1(n6569), .B2(n6583), .ZN(n6573)
         );
  AOI22_X1 U7514 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6589), .B1(n6571), 
        .B2(n6587), .ZN(n6572) );
  OAI211_X1 U7515 ( .C1(n6574), .C2(n6592), .A(n6573), .B(n6572), .ZN(U3113)
         );
  AOI22_X1 U7516 ( .A1(n6577), .A2(n6576), .B1(n6575), .B2(n6583), .ZN(n6580)
         );
  AOI22_X1 U7517 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6589), .B1(n6578), 
        .B2(n6587), .ZN(n6579) );
  OAI211_X1 U7518 ( .C1(n6582), .C2(n6581), .A(n6580), .B(n6579), .ZN(U3114)
         );
  AOI22_X1 U7519 ( .A1(n6586), .A2(n6585), .B1(n6584), .B2(n6583), .ZN(n6591)
         );
  AOI22_X1 U7520 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6589), .B1(n6588), 
        .B2(n6587), .ZN(n6590) );
  OAI211_X1 U7521 ( .C1(n6593), .C2(n6592), .A(n6591), .B(n6590), .ZN(U3115)
         );
  INV_X1 U7522 ( .A(n6594), .ZN(n6595) );
  AOI22_X1 U7523 ( .A1(n6597), .A2(n6596), .B1(n6595), .B2(n3730), .ZN(n6723)
         );
  NAND2_X1 U7524 ( .A1(n6598), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6728) );
  NAND3_X1 U7525 ( .A1(n6723), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6728), .ZN(n6602) );
  OAI211_X1 U7526 ( .C1(n6601), .C2(n6602), .A(n6600), .B(n6599), .ZN(n6604)
         );
  NAND2_X1 U7527 ( .A1(n6602), .A2(n6601), .ZN(n6603) );
  NAND2_X1 U7528 ( .A1(n6604), .A2(n6603), .ZN(n6605) );
  AOI222_X1 U7529 ( .A1(n6607), .A2(n6606), .B1(n6607), .B2(n6605), .C1(n6606), 
        .C2(n6605), .ZN(n6610) );
  OR2_X1 U7530 ( .A1(n6610), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6609)
         );
  NAND2_X1 U7531 ( .A1(n6609), .A2(n6608), .ZN(n6613) );
  NAND2_X1 U7532 ( .A1(n6610), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6612) );
  NAND3_X1 U7533 ( .A1(n6613), .A2(n6612), .A3(n6611), .ZN(n6622) );
  NOR2_X1 U7534 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6617) );
  INV_X1 U7535 ( .A(n6614), .ZN(n6616) );
  OAI211_X1 U7536 ( .C1(n6618), .C2(n6617), .A(n6616), .B(n6615), .ZN(n6619)
         );
  NOR2_X1 U7537 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  NOR2_X1 U7538 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4599), .ZN(n6649) );
  NAND2_X1 U7539 ( .A1(n6639), .A2(n6640), .ZN(n6624) );
  NAND2_X1 U7540 ( .A1(READY_N), .A2(n6747), .ZN(n6623) );
  NAND2_X1 U7541 ( .A1(n6624), .A2(n6623), .ZN(n6628) );
  NAND2_X1 U7542 ( .A1(n6626), .A2(n6625), .ZN(n6627) );
  NOR2_X1 U7543 ( .A1(n6649), .A2(n6719), .ZN(n6635) );
  OAI21_X1 U7544 ( .B1(n6742), .B2(n6629), .A(n6743), .ZN(n6630) );
  OR2_X1 U7545 ( .A1(n6719), .A2(n6630), .ZN(n6634) );
  INV_X1 U7546 ( .A(n6645), .ZN(n6717) );
  AOI21_X1 U7547 ( .B1(n6632), .B2(n6717), .A(n6631), .ZN(n6633) );
  OAI211_X1 U7548 ( .C1(n6635), .C2(n6743), .A(n6634), .B(n6633), .ZN(n6636)
         );
  INV_X1 U7549 ( .A(n6636), .ZN(n6637) );
  OAI21_X1 U7550 ( .B1(n6639), .B2(n6638), .A(n6637), .ZN(U3148) );
  AOI21_X1 U7551 ( .B1(n6641), .B2(n4599), .A(n6640), .ZN(n6644) );
  NAND2_X1 U7552 ( .A1(n6743), .A2(n6737), .ZN(n6646) );
  OAI211_X1 U7553 ( .C1(n6719), .C2(n6649), .A(STATE2_REG_1__SCAN_IN), .B(
        n6646), .ZN(n6642) );
  OAI211_X1 U7554 ( .C1(n6719), .C2(n6644), .A(n6643), .B(n6642), .ZN(U3149)
         );
  NAND3_X1 U7555 ( .A1(n6646), .A2(n6742), .A3(n6645), .ZN(n6648) );
  OAI21_X1 U7556 ( .B1(n6649), .B2(n6648), .A(n6647), .ZN(U3150) );
  INV_X1 U7557 ( .A(n6716), .ZN(n6650) );
  AND2_X1 U7558 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6650), .ZN(U3151) );
  AND2_X1 U7559 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6650), .ZN(U3152) );
  AND2_X1 U7560 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6650), .ZN(U3153) );
  AND2_X1 U7561 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6650), .ZN(U3154) );
  INV_X1 U7562 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6917) );
  NOR2_X1 U7563 ( .A1(n6716), .A2(n6917), .ZN(U3155) );
  AND2_X1 U7564 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6650), .ZN(U3156) );
  INV_X1 U7565 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6854) );
  NOR2_X1 U7566 ( .A1(n6716), .A2(n6854), .ZN(U3157) );
  AND2_X1 U7567 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6650), .ZN(U3158) );
  INV_X1 U7568 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6869) );
  NOR2_X1 U7569 ( .A1(n6716), .A2(n6869), .ZN(U3159) );
  AND2_X1 U7570 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6650), .ZN(U3160) );
  INV_X1 U7571 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6979) );
  NOR2_X1 U7572 ( .A1(n6716), .A2(n6979), .ZN(U3161) );
  AND2_X1 U7573 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6650), .ZN(U3162) );
  AND2_X1 U7574 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6650), .ZN(U3163) );
  AND2_X1 U7575 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6650), .ZN(U3164) );
  AND2_X1 U7576 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6650), .ZN(U3165) );
  AND2_X1 U7577 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6650), .ZN(U3166) );
  AND2_X1 U7578 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6650), .ZN(U3167) );
  AND2_X1 U7579 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6650), .ZN(U3168) );
  AND2_X1 U7580 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6650), .ZN(U3169) );
  AND2_X1 U7581 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6650), .ZN(U3170) );
  AND2_X1 U7582 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6650), .ZN(U3171) );
  AND2_X1 U7583 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6650), .ZN(U3172) );
  AND2_X1 U7584 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6650), .ZN(U3173) );
  AND2_X1 U7585 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6650), .ZN(U3174) );
  INV_X1 U7586 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6970) );
  NOR2_X1 U7587 ( .A1(n6716), .A2(n6970), .ZN(U3175) );
  AND2_X1 U7588 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6650), .ZN(U3176) );
  INV_X1 U7589 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6896) );
  NOR2_X1 U7590 ( .A1(n6716), .A2(n6896), .ZN(U3177) );
  AND2_X1 U7591 ( .A1(n6650), .A2(DATAWIDTH_REG_4__SCAN_IN), .ZN(U3178) );
  INV_X1 U7592 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n7023) );
  NOR2_X1 U7593 ( .A1(n6716), .A2(n7023), .ZN(U3179) );
  AND2_X1 U7594 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6650), .ZN(U3180) );
  INV_X1 U7595 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6654) );
  AOI221_X1 U7596 ( .B1(STATE_REG_1__SCAN_IN), .B2(HOLD), .C1(
        STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n6654), .ZN(n6653) );
  AND2_X1 U7597 ( .A1(n6664), .A2(STATE_REG_1__SCAN_IN), .ZN(n6651) );
  INV_X1 U7598 ( .A(NA_N), .ZN(n6924) );
  AOI221_X1 U7599 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6924), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6663) );
  AOI21_X1 U7600 ( .B1(READY_N), .B2(n6651), .A(n6663), .ZN(n6652) );
  OAI21_X1 U7601 ( .B1(n6712), .B2(n6653), .A(n6652), .ZN(U3181) );
  AND2_X1 U7602 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6657) );
  NOR2_X1 U7603 ( .A1(n4316), .A2(n6654), .ZN(n6659) );
  AOI21_X1 U7604 ( .B1(STATE_REG_1__SCAN_IN), .B2(HOLD), .A(n6659), .ZN(n6656)
         );
  NAND2_X1 U7605 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6660) );
  OAI211_X1 U7606 ( .C1(n6657), .C2(n6656), .A(n6655), .B(n6660), .ZN(U3182)
         );
  AOI221_X1 U7607 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4599), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6658) );
  AOI221_X1 U7608 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6658), .C2(HOLD), .A(n4316), .ZN(n6662) );
  AOI21_X1 U7609 ( .B1(n6659), .B2(n6924), .A(STATE_REG_2__SCAN_IN), .ZN(n6661) );
  OAI22_X1 U7610 ( .A1(n6663), .A2(n6662), .B1(n6661), .B2(n6660), .ZN(U3183)
         );
  NAND2_X1 U7611 ( .A1(n6664), .A2(n6712), .ZN(n6710) );
  NAND2_X1 U7612 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6712), .ZN(n6706) );
  INV_X1 U7613 ( .A(n6706), .ZN(n7147) );
  AOI22_X1 U7614 ( .A1(REIP_REG_1__SCAN_IN), .A2(n7147), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n7148), .ZN(n6665) );
  OAI21_X1 U7615 ( .B1(n6194), .B2(n6710), .A(n6665), .ZN(U3184) );
  AOI22_X1 U7616 ( .A1(REIP_REG_2__SCAN_IN), .A2(n7147), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n7148), .ZN(n6666) );
  OAI21_X1 U7617 ( .B1(n6667), .B2(n6710), .A(n6666), .ZN(U3185) );
  AOI22_X1 U7618 ( .A1(REIP_REG_3__SCAN_IN), .A2(n7147), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n7148), .ZN(n6668) );
  OAI21_X1 U7619 ( .B1(n6669), .B2(n6710), .A(n6668), .ZN(U3186) );
  AOI22_X1 U7620 ( .A1(REIP_REG_4__SCAN_IN), .A2(n7147), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n7148), .ZN(n6670) );
  OAI21_X1 U7621 ( .B1(n6671), .B2(n6710), .A(n6670), .ZN(U3187) );
  AOI22_X1 U7622 ( .A1(REIP_REG_5__SCAN_IN), .A2(n7147), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n7148), .ZN(n6672) );
  OAI21_X1 U7623 ( .B1(n6673), .B2(n6710), .A(n6672), .ZN(U3188) );
  AOI22_X1 U7624 ( .A1(REIP_REG_6__SCAN_IN), .A2(n7147), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n7148), .ZN(n6674) );
  OAI21_X1 U7625 ( .B1(n6993), .B2(n6710), .A(n6674), .ZN(U3189) );
  INV_X1 U7626 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n7007) );
  OAI222_X1 U7627 ( .A1(n6706), .A2(n6993), .B1(n7007), .B2(n6712), .C1(n5303), 
        .C2(n6710), .ZN(U3190) );
  INV_X1 U7628 ( .A(n6710), .ZN(n7146) );
  AOI222_X1 U7629 ( .A1(n7146), .A2(REIP_REG_9__SCAN_IN), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n7148), .C1(REIP_REG_8__SCAN_IN), .C2(
        n7147), .ZN(n6675) );
  INV_X1 U7630 ( .A(n6675), .ZN(U3191) );
  INV_X1 U7631 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6990) );
  AOI22_X1 U7632 ( .A1(REIP_REG_10__SCAN_IN), .A2(n7146), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n7148), .ZN(n6676) );
  OAI21_X1 U7633 ( .B1(n6990), .B2(n6706), .A(n6676), .ZN(U3192) );
  INV_X1 U7634 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6929) );
  AOI22_X1 U7635 ( .A1(REIP_REG_11__SCAN_IN), .A2(n7146), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n7148), .ZN(n6677) );
  OAI21_X1 U7636 ( .B1(n6929), .B2(n6706), .A(n6677), .ZN(U3193) );
  AOI22_X1 U7637 ( .A1(REIP_REG_12__SCAN_IN), .A2(n7146), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n7148), .ZN(n6678) );
  OAI21_X1 U7638 ( .B1(n6679), .B2(n6706), .A(n6678), .ZN(U3194) );
  AOI22_X1 U7639 ( .A1(REIP_REG_13__SCAN_IN), .A2(n7146), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n7148), .ZN(n6680) );
  OAI21_X1 U7640 ( .B1(n6902), .B2(n6706), .A(n6680), .ZN(U3195) );
  AOI22_X1 U7641 ( .A1(REIP_REG_14__SCAN_IN), .A2(n7146), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n7148), .ZN(n6681) );
  OAI21_X1 U7642 ( .B1(n6682), .B2(n6706), .A(n6681), .ZN(U3196) );
  AOI22_X1 U7643 ( .A1(REIP_REG_15__SCAN_IN), .A2(n7146), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n7148), .ZN(n6683) );
  OAI21_X1 U7644 ( .B1(n6684), .B2(n6706), .A(n6683), .ZN(U3197) );
  AOI22_X1 U7645 ( .A1(REIP_REG_16__SCAN_IN), .A2(n7146), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n7148), .ZN(n6685) );
  OAI21_X1 U7646 ( .B1(n6686), .B2(n6706), .A(n6685), .ZN(U3198) );
  INV_X1 U7647 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6688) );
  AOI22_X1 U7648 ( .A1(REIP_REG_17__SCAN_IN), .A2(n7146), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n7148), .ZN(n6687) );
  OAI21_X1 U7649 ( .B1(n6688), .B2(n6706), .A(n6687), .ZN(U3199) );
  AOI22_X1 U7650 ( .A1(REIP_REG_17__SCAN_IN), .A2(n7147), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n7148), .ZN(n6689) );
  OAI21_X1 U7651 ( .B1(n6690), .B2(n6710), .A(n6689), .ZN(U3200) );
  INV_X1 U7652 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6976) );
  OAI222_X1 U7653 ( .A1(n6710), .A2(n6691), .B1(n6976), .B2(n6712), .C1(n6690), 
        .C2(n6706), .ZN(U3201) );
  INV_X1 U7654 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n7053) );
  OAI222_X1 U7655 ( .A1(n6706), .A2(n6691), .B1(n7053), .B2(n6712), .C1(n6693), 
        .C2(n6710), .ZN(U3202) );
  INV_X1 U7656 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n7056) );
  OAI222_X1 U7657 ( .A1(n6706), .A2(n6693), .B1(n7056), .B2(n6712), .C1(n6692), 
        .C2(n6710), .ZN(U3203) );
  AOI22_X1 U7658 ( .A1(REIP_REG_21__SCAN_IN), .A2(n7147), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n7148), .ZN(n6694) );
  OAI21_X1 U7659 ( .B1(n6695), .B2(n6710), .A(n6694), .ZN(U3204) );
  AOI222_X1 U7660 ( .A1(n7147), .A2(REIP_REG_22__SCAN_IN), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n7148), .C1(REIP_REG_23__SCAN_IN), .C2(
        n7146), .ZN(n6696) );
  INV_X1 U7661 ( .A(n6696), .ZN(U3205) );
  AOI22_X1 U7662 ( .A1(REIP_REG_24__SCAN_IN), .A2(n7146), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n7148), .ZN(n6697) );
  OAI21_X1 U7663 ( .B1(n6698), .B2(n6706), .A(n6697), .ZN(U3206) );
  AOI222_X1 U7664 ( .A1(n7146), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n7148), .C1(REIP_REG_24__SCAN_IN), .C2(
        n7147), .ZN(n6699) );
  INV_X1 U7665 ( .A(n6699), .ZN(U3207) );
  AOI22_X1 U7666 ( .A1(REIP_REG_26__SCAN_IN), .A2(n7146), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n7148), .ZN(n6700) );
  OAI21_X1 U7667 ( .B1(n6701), .B2(n6706), .A(n6700), .ZN(U3208) );
  INV_X1 U7668 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6703) );
  AOI22_X1 U7669 ( .A1(REIP_REG_27__SCAN_IN), .A2(n7146), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n7148), .ZN(n6702) );
  OAI21_X1 U7670 ( .B1(n6703), .B2(n6706), .A(n6702), .ZN(U3209) );
  INV_X1 U7671 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n6844) );
  OAI222_X1 U7672 ( .A1(n6706), .A2(n6705), .B1(n6844), .B2(n6712), .C1(n6704), 
        .C2(n6710), .ZN(U3211) );
  AOI22_X1 U7673 ( .A1(REIP_REG_29__SCAN_IN), .A2(n7147), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n7148), .ZN(n6707) );
  OAI21_X1 U7674 ( .B1(n6708), .B2(n6710), .A(n6707), .ZN(U3212) );
  INV_X1 U7675 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6711) );
  AOI22_X1 U7676 ( .A1(REIP_REG_30__SCAN_IN), .A2(n7147), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n7148), .ZN(n6709) );
  OAI21_X1 U7677 ( .B1(n6711), .B2(n6710), .A(n6709), .ZN(U3213) );
  MUX2_X1 U7678 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n7148), .Z(U3445) );
  MUX2_X1 U7679 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n7148), .Z(U3446) );
  MUX2_X1 U7680 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n7148), .Z(U3447) );
  INV_X1 U7681 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6733) );
  INV_X1 U7682 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6898) );
  AOI22_X1 U7683 ( .A1(n6712), .A2(n6733), .B1(n6898), .B2(n7148), .ZN(U3448)
         );
  OAI21_X1 U7684 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6716), .A(n6714), .ZN(
        n6713) );
  INV_X1 U7685 ( .A(n6713), .ZN(U3451) );
  OAI21_X1 U7686 ( .B1(n6716), .B2(n6715), .A(n6714), .ZN(U3452) );
  AOI211_X1 U7687 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6719), .A(n6718), .B(
        n6717), .ZN(n6720) );
  INV_X1 U7688 ( .A(n6720), .ZN(U3453) );
  AOI21_X1 U7689 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n5451), .A(n6721), .ZN(
        n6722) );
  OAI211_X1 U7690 ( .C1(n6723), .C2(n6727), .A(n6725), .B(n6722), .ZN(n6724)
         );
  OAI21_X1 U7691 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6725), .A(n6724), 
        .ZN(n6726) );
  OAI21_X1 U7692 ( .B1(n6728), .B2(n6727), .A(n6726), .ZN(U3461) );
  AOI211_X1 U7693 ( .C1(REIP_REG_0__SCAN_IN), .C2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(REIP_REG_1__SCAN_IN), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6729) );
  AOI21_X1 U7694 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6729), .ZN(n6731) );
  INV_X1 U7695 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6730) );
  AOI22_X1 U7696 ( .A1(n6735), .A2(n6731), .B1(n6730), .B2(n6732), .ZN(U3468)
         );
  NOR2_X1 U7697 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6734) );
  AOI22_X1 U7698 ( .A1(n6735), .A2(n6734), .B1(n6733), .B2(n6732), .ZN(U3469)
         );
  NAND2_X1 U7699 ( .A1(n7148), .A2(W_R_N_REG_SCAN_IN), .ZN(n6736) );
  OAI21_X1 U7700 ( .B1(n7148), .B2(READREQUEST_REG_SCAN_IN), .A(n6736), .ZN(
        U3470) );
  AOI211_X1 U7701 ( .C1(n6739), .C2(n6738), .A(READY_N), .B(n6737), .ZN(n6741)
         );
  AND2_X1 U7702 ( .A1(n6741), .A2(n6740), .ZN(n6744) );
  OAI21_X1 U7703 ( .B1(n6744), .B2(n6743), .A(n6742), .ZN(n6749) );
  AOI211_X1 U7704 ( .C1(n6747), .C2(n4599), .A(n6746), .B(n6745), .ZN(n6748)
         );
  MUX2_X1 U7705 ( .A(n6749), .B(REQUESTPENDING_REG_SCAN_IN), .S(n6748), .Z(
        U3472) );
  MUX2_X1 U7706 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n7148), .Z(U3473) );
  AOI22_X1 U7707 ( .A1(EBX_REG_19__SCAN_IN), .A2(keyinput178), .B1(
        INSTQUEUE_REG_11__4__SCAN_IN), .B2(keyinput166), .ZN(n6750) );
  OAI221_X1 U7708 ( .B1(EBX_REG_19__SCAN_IN), .B2(keyinput178), .C1(
        INSTQUEUE_REG_11__4__SCAN_IN), .C2(keyinput166), .A(n6750), .ZN(n6757)
         );
  AOI22_X1 U7709 ( .A1(EAX_REG_28__SCAN_IN), .A2(keyinput206), .B1(
        INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput238), .ZN(n6751) );
  OAI221_X1 U7710 ( .B1(EAX_REG_28__SCAN_IN), .B2(keyinput206), .C1(
        INSTADDRPOINTER_REG_27__SCAN_IN), .C2(keyinput238), .A(n6751), .ZN(
        n6756) );
  AOI22_X1 U7711 ( .A1(DATAI_2_), .A2(keyinput171), .B1(DATAI_22_), .B2(
        keyinput200), .ZN(n6752) );
  OAI221_X1 U7712 ( .B1(DATAI_2_), .B2(keyinput171), .C1(DATAI_22_), .C2(
        keyinput200), .A(n6752), .ZN(n6755) );
  AOI22_X1 U7713 ( .A1(UWORD_REG_10__SCAN_IN), .A2(keyinput165), .B1(DATAI_12_), .B2(keyinput253), .ZN(n6753) );
  OAI221_X1 U7714 ( .B1(UWORD_REG_10__SCAN_IN), .B2(keyinput165), .C1(
        DATAI_12_), .C2(keyinput253), .A(n6753), .ZN(n6754) );
  NOR4_X1 U7715 ( .A1(n6757), .A2(n6756), .A3(n6755), .A4(n6754), .ZN(n6785)
         );
  AOI22_X1 U7716 ( .A1(LWORD_REG_0__SCAN_IN), .A2(keyinput155), .B1(
        INSTQUEUE_REG_3__6__SCAN_IN), .B2(keyinput164), .ZN(n6758) );
  OAI221_X1 U7717 ( .B1(LWORD_REG_0__SCAN_IN), .B2(keyinput155), .C1(
        INSTQUEUE_REG_3__6__SCAN_IN), .C2(keyinput164), .A(n6758), .ZN(n6765)
         );
  AOI22_X1 U7718 ( .A1(DATAO_REG_18__SCAN_IN), .A2(keyinput252), .B1(
        INSTQUEUE_REG_0__4__SCAN_IN), .B2(keyinput203), .ZN(n6759) );
  OAI221_X1 U7719 ( .B1(DATAO_REG_18__SCAN_IN), .B2(keyinput252), .C1(
        INSTQUEUE_REG_0__4__SCAN_IN), .C2(keyinput203), .A(n6759), .ZN(n6764)
         );
  AOI22_X1 U7720 ( .A1(DATAI_25_), .A2(keyinput215), .B1(
        INSTQUEUE_REG_9__1__SCAN_IN), .B2(keyinput224), .ZN(n6760) );
  OAI221_X1 U7721 ( .B1(DATAI_25_), .B2(keyinput215), .C1(
        INSTQUEUE_REG_9__1__SCAN_IN), .C2(keyinput224), .A(n6760), .ZN(n6763)
         );
  AOI22_X1 U7722 ( .A1(ADDRESS_REG_7__SCAN_IN), .A2(keyinput173), .B1(
        DATAO_REG_21__SCAN_IN), .B2(keyinput157), .ZN(n6761) );
  OAI221_X1 U7723 ( .B1(ADDRESS_REG_7__SCAN_IN), .B2(keyinput173), .C1(
        DATAO_REG_21__SCAN_IN), .C2(keyinput157), .A(n6761), .ZN(n6762) );
  NOR4_X1 U7724 ( .A1(n6765), .A2(n6764), .A3(n6763), .A4(n6762), .ZN(n6784)
         );
  AOI22_X1 U7725 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(keyinput249), .B1(
        INSTQUEUE_REG_4__1__SCAN_IN), .B2(keyinput193), .ZN(n6766) );
  OAI221_X1 U7726 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput249), 
        .C1(INSTQUEUE_REG_4__1__SCAN_IN), .C2(keyinput193), .A(n6766), .ZN(
        n6773) );
  AOI22_X1 U7727 ( .A1(REIP_REG_7__SCAN_IN), .A2(keyinput211), .B1(
        INSTQUEUE_REG_3__1__SCAN_IN), .B2(keyinput158), .ZN(n6767) );
  OAI221_X1 U7728 ( .B1(REIP_REG_7__SCAN_IN), .B2(keyinput211), .C1(
        INSTQUEUE_REG_3__1__SCAN_IN), .C2(keyinput158), .A(n6767), .ZN(n6772)
         );
  AOI22_X1 U7729 ( .A1(BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput219), .B1(
        REIP_REG_9__SCAN_IN), .B2(keyinput223), .ZN(n6768) );
  OAI221_X1 U7730 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput219), .C1(
        REIP_REG_9__SCAN_IN), .C2(keyinput223), .A(n6768), .ZN(n6771) );
  AOI22_X1 U7731 ( .A1(UWORD_REG_3__SCAN_IN), .A2(keyinput179), .B1(
        EBX_REG_25__SCAN_IN), .B2(keyinput180), .ZN(n6769) );
  OAI221_X1 U7732 ( .B1(UWORD_REG_3__SCAN_IN), .B2(keyinput179), .C1(
        EBX_REG_25__SCAN_IN), .C2(keyinput180), .A(n6769), .ZN(n6770) );
  NOR4_X1 U7733 ( .A1(n6773), .A2(n6772), .A3(n6771), .A4(n6770), .ZN(n6783)
         );
  AOI22_X1 U7734 ( .A1(ADS_N_REG_SCAN_IN), .A2(keyinput185), .B1(
        DATAWIDTH_REG_7__SCAN_IN), .B2(keyinput194), .ZN(n6774) );
  OAI221_X1 U7735 ( .B1(ADS_N_REG_SCAN_IN), .B2(keyinput185), .C1(
        DATAWIDTH_REG_7__SCAN_IN), .C2(keyinput194), .A(n6774), .ZN(n6781) );
  AOI22_X1 U7736 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(keyinput136), .B1(
        EBX_REG_14__SCAN_IN), .B2(keyinput246), .ZN(n6775) );
  OAI221_X1 U7737 ( .B1(DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput136), .C1(
        EBX_REG_14__SCAN_IN), .C2(keyinput246), .A(n6775), .ZN(n6780) );
  AOI22_X1 U7738 ( .A1(EAX_REG_19__SCAN_IN), .A2(keyinput210), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(keyinput184), .ZN(n6776) );
  OAI221_X1 U7739 ( .B1(EAX_REG_19__SCAN_IN), .B2(keyinput210), .C1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .C2(keyinput184), .A(n6776), .ZN(
        n6779) );
  AOI22_X1 U7740 ( .A1(LWORD_REG_8__SCAN_IN), .A2(keyinput237), .B1(
        INSTQUEUE_REG_14__6__SCAN_IN), .B2(keyinput192), .ZN(n6777) );
  OAI221_X1 U7741 ( .B1(LWORD_REG_8__SCAN_IN), .B2(keyinput237), .C1(
        INSTQUEUE_REG_14__6__SCAN_IN), .C2(keyinput192), .A(n6777), .ZN(n6778)
         );
  NOR4_X1 U7742 ( .A1(n6781), .A2(n6780), .A3(n6779), .A4(n6778), .ZN(n6782)
         );
  NAND4_X1 U7743 ( .A1(n6785), .A2(n6784), .A3(n6783), .A4(n6782), .ZN(n6942)
         );
  AOI22_X1 U7744 ( .A1(ADDRESS_REG_19__SCAN_IN), .A2(keyinput162), .B1(
        EBX_REG_18__SCAN_IN), .B2(keyinput232), .ZN(n6786) );
  OAI221_X1 U7745 ( .B1(ADDRESS_REG_19__SCAN_IN), .B2(keyinput162), .C1(
        EBX_REG_18__SCAN_IN), .C2(keyinput232), .A(n6786), .ZN(n6793) );
  AOI22_X1 U7746 ( .A1(EAX_REG_22__SCAN_IN), .A2(keyinput245), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput153), .ZN(n6787) );
  OAI221_X1 U7747 ( .B1(EAX_REG_22__SCAN_IN), .B2(keyinput245), .C1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .C2(keyinput153), .A(n6787), .ZN(
        n6792) );
  AOI22_X1 U7748 ( .A1(EAX_REG_24__SCAN_IN), .A2(keyinput214), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(keyinput150), .ZN(n6788) );
  OAI221_X1 U7749 ( .B1(EAX_REG_24__SCAN_IN), .B2(keyinput214), .C1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .C2(keyinput150), .A(n6788), .ZN(
        n6791) );
  AOI22_X1 U7750 ( .A1(ADDRESS_REG_23__SCAN_IN), .A2(keyinput149), .B1(
        REIP_REG_5__SCAN_IN), .B2(keyinput176), .ZN(n6789) );
  OAI221_X1 U7751 ( .B1(ADDRESS_REG_23__SCAN_IN), .B2(keyinput149), .C1(
        REIP_REG_5__SCAN_IN), .C2(keyinput176), .A(n6789), .ZN(n6790) );
  NOR4_X1 U7752 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6824)
         );
  AOI22_X1 U7753 ( .A1(EAX_REG_0__SCAN_IN), .A2(keyinput140), .B1(
        EAX_REG_14__SCAN_IN), .B2(keyinput182), .ZN(n6794) );
  OAI221_X1 U7754 ( .B1(EAX_REG_0__SCAN_IN), .B2(keyinput140), .C1(
        EAX_REG_14__SCAN_IN), .C2(keyinput182), .A(n6794), .ZN(n6801) );
  AOI22_X1 U7755 ( .A1(ADDRESS_REG_18__SCAN_IN), .A2(keyinput145), .B1(
        DATAI_17_), .B2(keyinput240), .ZN(n6795) );
  OAI221_X1 U7756 ( .B1(ADDRESS_REG_18__SCAN_IN), .B2(keyinput145), .C1(
        DATAI_17_), .C2(keyinput240), .A(n6795), .ZN(n6800) );
  AOI22_X1 U7757 ( .A1(EAX_REG_16__SCAN_IN), .A2(keyinput144), .B1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput242), .ZN(n6796) );
  OAI221_X1 U7758 ( .B1(EAX_REG_16__SCAN_IN), .B2(keyinput144), .C1(
        PHYADDRPOINTER_REG_13__SCAN_IN), .C2(keyinput242), .A(n6796), .ZN(
        n6799) );
  AOI22_X1 U7759 ( .A1(LWORD_REG_11__SCAN_IN), .A2(keyinput146), .B1(
        INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput169), .ZN(n6797) );
  OAI221_X1 U7760 ( .B1(LWORD_REG_11__SCAN_IN), .B2(keyinput146), .C1(
        INSTQUEUE_REG_9__4__SCAN_IN), .C2(keyinput169), .A(n6797), .ZN(n6798)
         );
  NOR4_X1 U7761 ( .A1(n6801), .A2(n6800), .A3(n6799), .A4(n6798), .ZN(n6823)
         );
  AOI22_X1 U7762 ( .A1(ADDRESS_REG_21__SCAN_IN), .A2(keyinput213), .B1(
        REIP_REG_18__SCAN_IN), .B2(keyinput235), .ZN(n6802) );
  OAI221_X1 U7763 ( .B1(ADDRESS_REG_21__SCAN_IN), .B2(keyinput213), .C1(
        REIP_REG_18__SCAN_IN), .C2(keyinput235), .A(n6802), .ZN(n6809) );
  AOI22_X1 U7764 ( .A1(DATAO_REG_0__SCAN_IN), .A2(keyinput234), .B1(
        INSTQUEUE_REG_5__6__SCAN_IN), .B2(keyinput205), .ZN(n6803) );
  OAI221_X1 U7765 ( .B1(DATAO_REG_0__SCAN_IN), .B2(keyinput234), .C1(
        INSTQUEUE_REG_5__6__SCAN_IN), .C2(keyinput205), .A(n6803), .ZN(n6808)
         );
  AOI22_X1 U7766 ( .A1(REIP_REG_8__SCAN_IN), .A2(keyinput152), .B1(
        INSTQUEUE_REG_3__0__SCAN_IN), .B2(keyinput129), .ZN(n6804) );
  OAI221_X1 U7767 ( .B1(REIP_REG_8__SCAN_IN), .B2(keyinput152), .C1(
        INSTQUEUE_REG_3__0__SCAN_IN), .C2(keyinput129), .A(n6804), .ZN(n6807)
         );
  AOI22_X1 U7768 ( .A1(EAX_REG_18__SCAN_IN), .A2(keyinput209), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput239), .ZN(n6805) );
  OAI221_X1 U7769 ( .B1(EAX_REG_18__SCAN_IN), .B2(keyinput209), .C1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .C2(keyinput239), .A(n6805), .ZN(n6806) );
  NOR4_X1 U7770 ( .A1(n6809), .A2(n6808), .A3(n6807), .A4(n6806), .ZN(n6822)
         );
  AOI22_X1 U7771 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(keyinput247), 
        .B1(INSTQUEUE_REG_11__6__SCAN_IN), .B2(keyinput147), .ZN(n6810) );
  OAI221_X1 U7772 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput247), 
        .C1(INSTQUEUE_REG_11__6__SCAN_IN), .C2(keyinput147), .A(n6810), .ZN(
        n6820) );
  AOI22_X1 U7773 ( .A1(DATAI_7_), .A2(keyinput131), .B1(
        INSTQUEUE_REG_11__2__SCAN_IN), .B2(keyinput241), .ZN(n6811) );
  OAI221_X1 U7774 ( .B1(DATAI_7_), .B2(keyinput131), .C1(
        INSTQUEUE_REG_11__2__SCAN_IN), .C2(keyinput241), .A(n6811), .ZN(n6819)
         );
  INV_X1 U7775 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6814) );
  AOI22_X1 U7776 ( .A1(n6814), .A2(keyinput148), .B1(keyinput251), .B2(n6813), 
        .ZN(n6812) );
  OAI221_X1 U7777 ( .B1(n6814), .B2(keyinput148), .C1(n6813), .C2(keyinput251), 
        .A(n6812), .ZN(n6818) );
  AOI22_X1 U7778 ( .A1(n7004), .A2(keyinput190), .B1(n6816), .B2(keyinput230), 
        .ZN(n6815) );
  OAI221_X1 U7779 ( .B1(n7004), .B2(keyinput190), .C1(n6816), .C2(keyinput230), 
        .A(n6815), .ZN(n6817) );
  NOR4_X1 U7780 ( .A1(n6820), .A2(n6819), .A3(n6818), .A4(n6817), .ZN(n6821)
         );
  NAND4_X1 U7781 ( .A1(n6824), .A2(n6823), .A3(n6822), .A4(n6821), .ZN(n6941)
         );
  INV_X1 U7782 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6826) );
  AOI22_X1 U7783 ( .A1(n6827), .A2(keyinput244), .B1(n6826), .B2(keyinput170), 
        .ZN(n6825) );
  OAI221_X1 U7784 ( .B1(n6827), .B2(keyinput244), .C1(n6826), .C2(keyinput170), 
        .A(n6825), .ZN(n6838) );
  INV_X1 U7785 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6830) );
  AOI22_X1 U7786 ( .A1(n6830), .A2(keyinput163), .B1(n6829), .B2(keyinput159), 
        .ZN(n6828) );
  OAI221_X1 U7787 ( .B1(n6830), .B2(keyinput163), .C1(n6829), .C2(keyinput159), 
        .A(n6828), .ZN(n6837) );
  INV_X1 U7788 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6833) );
  AOI22_X1 U7789 ( .A1(n6833), .A2(keyinput254), .B1(keyinput135), .B2(n6832), 
        .ZN(n6831) );
  OAI221_X1 U7790 ( .B1(n6833), .B2(keyinput254), .C1(n6832), .C2(keyinput135), 
        .A(n6831), .ZN(n6836) );
  AOI22_X1 U7791 ( .A1(n7023), .A2(keyinput250), .B1(n3914), .B2(keyinput189), 
        .ZN(n6834) );
  OAI221_X1 U7792 ( .B1(n7023), .B2(keyinput250), .C1(n3914), .C2(keyinput189), 
        .A(n6834), .ZN(n6835) );
  NOR4_X1 U7793 ( .A1(n6838), .A2(n6837), .A3(n6836), .A4(n6835), .ZN(n6881)
         );
  INV_X1 U7794 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6986) );
  AOI22_X1 U7795 ( .A1(n6948), .A2(keyinput195), .B1(keyinput128), .B2(n6986), 
        .ZN(n6839) );
  OAI221_X1 U7796 ( .B1(n6948), .B2(keyinput195), .C1(n6986), .C2(keyinput128), 
        .A(n6839), .ZN(n6850) );
  AOI22_X1 U7797 ( .A1(n5062), .A2(keyinput177), .B1(keyinput134), .B2(n6841), 
        .ZN(n6840) );
  OAI221_X1 U7798 ( .B1(n5062), .B2(keyinput177), .C1(n6841), .C2(keyinput134), 
        .A(n6840), .ZN(n6849) );
  AOI22_X1 U7799 ( .A1(n6844), .A2(keyinput225), .B1(n6843), .B2(keyinput168), 
        .ZN(n6842) );
  OAI221_X1 U7800 ( .B1(n6844), .B2(keyinput225), .C1(n6843), .C2(keyinput168), 
        .A(n6842), .ZN(n6848) );
  INV_X1 U7801 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6846) );
  INV_X1 U7802 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6962) );
  AOI22_X1 U7803 ( .A1(n6846), .A2(keyinput248), .B1(keyinput229), .B2(n6962), 
        .ZN(n6845) );
  OAI221_X1 U7804 ( .B1(n6846), .B2(keyinput248), .C1(n6962), .C2(keyinput229), 
        .A(n6845), .ZN(n6847) );
  NOR4_X1 U7805 ( .A1(n6850), .A2(n6849), .A3(n6848), .A4(n6847), .ZN(n6880)
         );
  INV_X1 U7806 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n7012) );
  AOI22_X1 U7807 ( .A1(n6852), .A2(keyinput167), .B1(n7012), .B2(keyinput208), 
        .ZN(n6851) );
  OAI221_X1 U7808 ( .B1(n6852), .B2(keyinput167), .C1(n7012), .C2(keyinput208), 
        .A(n6851), .ZN(n6864) );
  AOI22_X1 U7809 ( .A1(n6854), .A2(keyinput243), .B1(n6975), .B2(keyinput139), 
        .ZN(n6853) );
  OAI221_X1 U7810 ( .B1(n6854), .B2(keyinput243), .C1(n6975), .C2(keyinput139), 
        .A(n6853), .ZN(n6863) );
  INV_X1 U7811 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n6857) );
  INV_X1 U7812 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n6856) );
  AOI22_X1 U7813 ( .A1(n6857), .A2(keyinput220), .B1(n6856), .B2(keyinput188), 
        .ZN(n6855) );
  OAI221_X1 U7814 ( .B1(n6857), .B2(keyinput220), .C1(n6856), .C2(keyinput188), 
        .A(n6855), .ZN(n6862) );
  AOI22_X1 U7815 ( .A1(n6860), .A2(keyinput222), .B1(n6859), .B2(keyinput228), 
        .ZN(n6858) );
  OAI221_X1 U7816 ( .B1(n6860), .B2(keyinput222), .C1(n6859), .C2(keyinput228), 
        .A(n6858), .ZN(n6861) );
  NOR4_X1 U7817 ( .A1(n6864), .A2(n6863), .A3(n6862), .A4(n6861), .ZN(n6879)
         );
  INV_X1 U7818 ( .A(LWORD_REG_1__SCAN_IN), .ZN(n6866) );
  AOI22_X1 U7819 ( .A1(n6866), .A2(keyinput138), .B1(keyinput132), .B2(n6969), 
        .ZN(n6865) );
  OAI221_X1 U7820 ( .B1(n6866), .B2(keyinput138), .C1(n6969), .C2(keyinput132), 
        .A(n6865), .ZN(n6877) );
  AOI22_X1 U7821 ( .A1(n6869), .A2(keyinput172), .B1(n6868), .B2(keyinput207), 
        .ZN(n6867) );
  OAI221_X1 U7822 ( .B1(n6869), .B2(keyinput172), .C1(n6868), .C2(keyinput207), 
        .A(n6867), .ZN(n6876) );
  INV_X1 U7823 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n6871) );
  INV_X1 U7824 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n7021) );
  AOI22_X1 U7825 ( .A1(n6871), .A2(keyinput255), .B1(n7021), .B2(keyinput216), 
        .ZN(n6870) );
  OAI221_X1 U7826 ( .B1(n6871), .B2(keyinput255), .C1(n7021), .C2(keyinput216), 
        .A(n6870), .ZN(n6875) );
  INV_X1 U7827 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6873) );
  AOI22_X1 U7828 ( .A1(n6873), .A2(keyinput217), .B1(n6960), .B2(keyinput218), 
        .ZN(n6872) );
  OAI221_X1 U7829 ( .B1(n6873), .B2(keyinput217), .C1(n6960), .C2(keyinput218), 
        .A(n6872), .ZN(n6874) );
  NOR4_X1 U7830 ( .A1(n6877), .A2(n6876), .A3(n6875), .A4(n6874), .ZN(n6878)
         );
  NAND4_X1 U7831 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n6940)
         );
  AOI22_X1 U7832 ( .A1(n6979), .A2(keyinput212), .B1(n6883), .B2(keyinput197), 
        .ZN(n6882) );
  OAI221_X1 U7833 ( .B1(n6979), .B2(keyinput212), .C1(n6883), .C2(keyinput197), 
        .A(n6882), .ZN(n6894) );
  AOI22_X1 U7834 ( .A1(n6973), .A2(keyinput226), .B1(n6885), .B2(keyinput227), 
        .ZN(n6884) );
  OAI221_X1 U7835 ( .B1(n6973), .B2(keyinput226), .C1(n6885), .C2(keyinput227), 
        .A(n6884), .ZN(n6893) );
  AOI22_X1 U7836 ( .A1(n6888), .A2(keyinput160), .B1(n6887), .B2(keyinput141), 
        .ZN(n6886) );
  OAI221_X1 U7837 ( .B1(n6888), .B2(keyinput160), .C1(n6887), .C2(keyinput141), 
        .A(n6886), .ZN(n6892) );
  XOR2_X1 U7838 ( .A(n7050), .B(keyinput161), .Z(n6890) );
  XNOR2_X1 U7839 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .B(keyinput156), .ZN(n6889) );
  NAND2_X1 U7840 ( .A1(n6890), .A2(n6889), .ZN(n6891) );
  NOR4_X1 U7841 ( .A1(n6894), .A2(n6893), .A3(n6892), .A4(n6891), .ZN(n6938)
         );
  INV_X1 U7842 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n7011) );
  AOI22_X1 U7843 ( .A1(n6896), .A2(keyinput175), .B1(n7011), .B2(keyinput154), 
        .ZN(n6895) );
  OAI221_X1 U7844 ( .B1(n6896), .B2(keyinput175), .C1(n7011), .C2(keyinput154), 
        .A(n6895), .ZN(n6908) );
  AOI22_X1 U7845 ( .A1(n6985), .A2(keyinput137), .B1(keyinput191), .B2(n6898), 
        .ZN(n6897) );
  OAI221_X1 U7846 ( .B1(n6985), .B2(keyinput137), .C1(n6898), .C2(keyinput191), 
        .A(n6897), .ZN(n6907) );
  INV_X1 U7847 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n6901) );
  INV_X1 U7848 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n6900) );
  AOI22_X1 U7849 ( .A1(n6901), .A2(keyinput183), .B1(keyinput196), .B2(n6900), 
        .ZN(n6899) );
  OAI221_X1 U7850 ( .B1(n6901), .B2(keyinput183), .C1(n6900), .C2(keyinput196), 
        .A(n6899), .ZN(n6906) );
  XOR2_X1 U7851 ( .A(n6902), .B(keyinput198), .Z(n6904) );
  XNOR2_X1 U7852 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .B(keyinput236), .ZN(n6903) );
  NAND2_X1 U7853 ( .A1(n6904), .A2(n6903), .ZN(n6905) );
  NOR4_X1 U7854 ( .A1(n6908), .A2(n6907), .A3(n6906), .A4(n6905), .ZN(n6937)
         );
  INV_X1 U7855 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6911) );
  AOI22_X1 U7856 ( .A1(n6911), .A2(keyinput187), .B1(n6910), .B2(keyinput186), 
        .ZN(n6909) );
  OAI221_X1 U7857 ( .B1(n6911), .B2(keyinput187), .C1(n6910), .C2(keyinput186), 
        .A(n6909), .ZN(n6922) );
  INV_X1 U7858 ( .A(DATAI_15_), .ZN(n6913) );
  AOI22_X1 U7859 ( .A1(n7037), .A2(keyinput174), .B1(keyinput130), .B2(n6913), 
        .ZN(n6912) );
  OAI221_X1 U7860 ( .B1(n7037), .B2(keyinput174), .C1(n6913), .C2(keyinput130), 
        .A(n6912), .ZN(n6921) );
  INV_X1 U7861 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6915) );
  AOI22_X1 U7862 ( .A1(n6915), .A2(keyinput221), .B1(keyinput202), .B2(n6976), 
        .ZN(n6914) );
  OAI221_X1 U7863 ( .B1(n6915), .B2(keyinput221), .C1(n6976), .C2(keyinput202), 
        .A(n6914), .ZN(n6920) );
  INV_X1 U7864 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n6918) );
  AOI22_X1 U7865 ( .A1(n6918), .A2(keyinput199), .B1(keyinput181), .B2(n6917), 
        .ZN(n6916) );
  OAI221_X1 U7866 ( .B1(n6918), .B2(keyinput199), .C1(n6917), .C2(keyinput181), 
        .A(n6916), .ZN(n6919) );
  NOR4_X1 U7867 ( .A1(n6922), .A2(n6921), .A3(n6920), .A4(n6919), .ZN(n6936)
         );
  AOI22_X1 U7868 ( .A1(n6925), .A2(keyinput233), .B1(keyinput143), .B2(n6924), 
        .ZN(n6923) );
  OAI221_X1 U7869 ( .B1(n6925), .B2(keyinput233), .C1(n6924), .C2(keyinput143), 
        .A(n6923), .ZN(n6934) );
  INV_X1 U7870 ( .A(LWORD_REG_3__SCAN_IN), .ZN(n6927) );
  AOI22_X1 U7871 ( .A1(n7007), .A2(keyinput201), .B1(n6927), .B2(keyinput142), 
        .ZN(n6926) );
  OAI221_X1 U7872 ( .B1(n7007), .B2(keyinput201), .C1(n6927), .C2(keyinput142), 
        .A(n6926), .ZN(n6933) );
  AOI22_X1 U7873 ( .A1(n6929), .A2(keyinput133), .B1(n6946), .B2(keyinput204), 
        .ZN(n6928) );
  OAI221_X1 U7874 ( .B1(n6929), .B2(keyinput133), .C1(n6946), .C2(keyinput204), 
        .A(n6928), .ZN(n6932) );
  INV_X1 U7875 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n7008) );
  AOI22_X1 U7876 ( .A1(n4599), .A2(keyinput151), .B1(n7008), .B2(keyinput231), 
        .ZN(n6930) );
  OAI221_X1 U7877 ( .B1(n4599), .B2(keyinput151), .C1(n7008), .C2(keyinput231), 
        .A(n6930), .ZN(n6931) );
  NOR4_X1 U7878 ( .A1(n6934), .A2(n6933), .A3(n6932), .A4(n6931), .ZN(n6935)
         );
  NAND4_X1 U7879 ( .A1(n6938), .A2(n6937), .A3(n6936), .A4(n6935), .ZN(n6939)
         );
  NOR4_X1 U7880 ( .A1(n6942), .A2(n6941), .A3(n6940), .A4(n6939), .ZN(n7145)
         );
  AOI22_X1 U7881 ( .A1(DATAI_7_), .A2(keyinput3), .B1(REIP_REG_10__SCAN_IN), 
        .B2(keyinput5), .ZN(n6943) );
  OAI221_X1 U7882 ( .B1(DATAI_7_), .B2(keyinput3), .C1(REIP_REG_10__SCAN_IN), 
        .C2(keyinput5), .A(n6943), .ZN(n6953) );
  AOI22_X1 U7883 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(keyinput8), .B1(
        LWORD_REG_3__SCAN_IN), .B2(keyinput14), .ZN(n6944) );
  OAI221_X1 U7884 ( .B1(DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput8), .C1(
        LWORD_REG_3__SCAN_IN), .C2(keyinput14), .A(n6944), .ZN(n6952) );
  AOI22_X1 U7885 ( .A1(LWORD_REG_8__SCAN_IN), .A2(keyinput109), .B1(n6946), 
        .B2(keyinput76), .ZN(n6945) );
  OAI221_X1 U7886 ( .B1(LWORD_REG_8__SCAN_IN), .B2(keyinput109), .C1(n6946), 
        .C2(keyinput76), .A(n6945), .ZN(n6951) );
  INV_X1 U7887 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6949) );
  AOI22_X1 U7888 ( .A1(n6949), .A2(keyinput38), .B1(keyinput67), .B2(n6948), 
        .ZN(n6947) );
  OAI221_X1 U7889 ( .B1(n6949), .B2(keyinput38), .C1(n6948), .C2(keyinput67), 
        .A(n6947), .ZN(n6950) );
  NOR4_X1 U7890 ( .A1(n6953), .A2(n6952), .A3(n6951), .A4(n6950), .ZN(n7002)
         );
  AOI22_X1 U7891 ( .A1(n6955), .A2(keyinput50), .B1(n5630), .B2(keyinput52), 
        .ZN(n6954) );
  OAI221_X1 U7892 ( .B1(n6955), .B2(keyinput50), .C1(n5630), .C2(keyinput52), 
        .A(n6954), .ZN(n6967) );
  AOI22_X1 U7893 ( .A1(n6958), .A2(keyinput56), .B1(keyinput121), .B2(n6957), 
        .ZN(n6956) );
  OAI221_X1 U7894 ( .B1(n6958), .B2(keyinput56), .C1(n6957), .C2(keyinput121), 
        .A(n6956), .ZN(n6966) );
  AOI22_X1 U7895 ( .A1(n5303), .A2(keyinput24), .B1(n6960), .B2(keyinput90), 
        .ZN(n6959) );
  OAI221_X1 U7896 ( .B1(n5303), .B2(keyinput24), .C1(n6960), .C2(keyinput90), 
        .A(n6959), .ZN(n6965) );
  INV_X1 U7897 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6963) );
  AOI22_X1 U7898 ( .A1(n6963), .A2(keyinput19), .B1(n6962), .B2(keyinput101), 
        .ZN(n6961) );
  OAI221_X1 U7899 ( .B1(n6963), .B2(keyinput19), .C1(n6962), .C2(keyinput101), 
        .A(n6961), .ZN(n6964) );
  NOR4_X1 U7900 ( .A1(n6967), .A2(n6966), .A3(n6965), .A4(n6964), .ZN(n7001)
         );
  AOI22_X1 U7901 ( .A1(n6970), .A2(keyinput66), .B1(n6969), .B2(keyinput4), 
        .ZN(n6968) );
  OAI221_X1 U7902 ( .B1(n6970), .B2(keyinput66), .C1(n6969), .C2(keyinput4), 
        .A(n6968), .ZN(n6983) );
  AOI22_X1 U7903 ( .A1(n6973), .A2(keyinput98), .B1(keyinput86), .B2(n6972), 
        .ZN(n6971) );
  OAI221_X1 U7904 ( .B1(n6973), .B2(keyinput98), .C1(n6972), .C2(keyinput86), 
        .A(n6971), .ZN(n6982) );
  AOI22_X1 U7905 ( .A1(n6976), .A2(keyinput74), .B1(n6975), .B2(keyinput11), 
        .ZN(n6974) );
  OAI221_X1 U7906 ( .B1(n6976), .B2(keyinput74), .C1(n6975), .C2(keyinput11), 
        .A(n6974), .ZN(n6981) );
  AOI22_X1 U7907 ( .A1(n6979), .A2(keyinput84), .B1(n6978), .B2(keyinput75), 
        .ZN(n6977) );
  OAI221_X1 U7908 ( .B1(n6979), .B2(keyinput84), .C1(n6978), .C2(keyinput75), 
        .A(n6977), .ZN(n6980) );
  NOR4_X1 U7909 ( .A1(n6983), .A2(n6982), .A3(n6981), .A4(n6980), .ZN(n7000)
         );
  AOI22_X1 U7910 ( .A1(n6986), .A2(keyinput0), .B1(n6985), .B2(keyinput9), 
        .ZN(n6984) );
  OAI221_X1 U7911 ( .B1(n6986), .B2(keyinput0), .C1(n6985), .C2(keyinput9), 
        .A(n6984), .ZN(n6998) );
  AOI22_X1 U7912 ( .A1(n4599), .A2(keyinput23), .B1(keyinput12), .B2(n6988), 
        .ZN(n6987) );
  OAI221_X1 U7913 ( .B1(n4599), .B2(keyinput23), .C1(n6988), .C2(keyinput12), 
        .A(n6987), .ZN(n6997) );
  INV_X1 U7914 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6991) );
  AOI22_X1 U7915 ( .A1(n6991), .A2(keyinput1), .B1(keyinput95), .B2(n6990), 
        .ZN(n6989) );
  OAI221_X1 U7916 ( .B1(n6991), .B2(keyinput1), .C1(n6990), .C2(keyinput95), 
        .A(n6989), .ZN(n6996) );
  INV_X1 U7917 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n6994) );
  AOI22_X1 U7918 ( .A1(n6994), .A2(keyinput106), .B1(n6993), .B2(keyinput83), 
        .ZN(n6992) );
  OAI221_X1 U7919 ( .B1(n6994), .B2(keyinput106), .C1(n6993), .C2(keyinput83), 
        .A(n6992), .ZN(n6995) );
  NOR4_X1 U7920 ( .A1(n6998), .A2(n6997), .A3(n6996), .A4(n6995), .ZN(n6999)
         );
  NAND4_X1 U7921 ( .A1(n7002), .A2(n7001), .A3(n7000), .A4(n6999), .ZN(n7144)
         );
  INV_X1 U7922 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n7005) );
  AOI22_X1 U7923 ( .A1(n7005), .A2(keyinput64), .B1(keyinput62), .B2(n7004), 
        .ZN(n7003) );
  OAI221_X1 U7924 ( .B1(n7005), .B2(keyinput64), .C1(n7004), .C2(keyinput62), 
        .A(n7003), .ZN(n7018) );
  AOI22_X1 U7925 ( .A1(n7008), .A2(keyinput103), .B1(keyinput73), .B2(n7007), 
        .ZN(n7006) );
  OAI221_X1 U7926 ( .B1(n7008), .B2(keyinput103), .C1(n7007), .C2(keyinput73), 
        .A(n7006), .ZN(n7017) );
  INV_X1 U7927 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n7010) );
  AOI22_X1 U7928 ( .A1(n7011), .A2(keyinput26), .B1(n7010), .B2(keyinput65), 
        .ZN(n7009) );
  OAI221_X1 U7929 ( .B1(n7011), .B2(keyinput26), .C1(n7010), .C2(keyinput65), 
        .A(n7009), .ZN(n7016) );
  XOR2_X1 U7930 ( .A(n7012), .B(keyinput80), .Z(n7014) );
  XNOR2_X1 U7931 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .B(keyinput113), .ZN(
        n7013) );
  NAND2_X1 U7932 ( .A1(n7014), .A2(n7013), .ZN(n7015) );
  NOR4_X1 U7933 ( .A1(n7018), .A2(n7017), .A3(n7016), .A4(n7015), .ZN(n7067)
         );
  INV_X1 U7934 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n7020) );
  AOI22_X1 U7935 ( .A1(n7021), .A2(keyinput88), .B1(keyinput124), .B2(n7020), 
        .ZN(n7019) );
  OAI221_X1 U7936 ( .B1(n7021), .B2(keyinput88), .C1(n7020), .C2(keyinput124), 
        .A(n7019), .ZN(n7034) );
  AOI22_X1 U7937 ( .A1(n7024), .A2(keyinput112), .B1(keyinput122), .B2(n7023), 
        .ZN(n7022) );
  OAI221_X1 U7938 ( .B1(n7024), .B2(keyinput112), .C1(n7023), .C2(keyinput122), 
        .A(n7022), .ZN(n7033) );
  INV_X1 U7939 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n7027) );
  AOI22_X1 U7940 ( .A1(n7027), .A2(keyinput41), .B1(keyinput25), .B2(n7026), 
        .ZN(n7025) );
  OAI221_X1 U7941 ( .B1(n7027), .B2(keyinput41), .C1(n7026), .C2(keyinput25), 
        .A(n7025), .ZN(n7032) );
  AOI22_X1 U7942 ( .A1(n7030), .A2(keyinput118), .B1(keyinput81), .B2(n7029), 
        .ZN(n7028) );
  OAI221_X1 U7943 ( .B1(n7030), .B2(keyinput118), .C1(n7029), .C2(keyinput81), 
        .A(n7028), .ZN(n7031) );
  NOR4_X1 U7944 ( .A1(n7034), .A2(n7033), .A3(n7032), .A4(n7031), .ZN(n7066)
         );
  INV_X1 U7945 ( .A(DATAI_12_), .ZN(n7036) );
  AOI22_X1 U7946 ( .A1(n7037), .A2(keyinput46), .B1(keyinput125), .B2(n7036), 
        .ZN(n7035) );
  OAI221_X1 U7947 ( .B1(n7037), .B2(keyinput46), .C1(n7036), .C2(keyinput125), 
        .A(n7035), .ZN(n7047) );
  INV_X1 U7948 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n7040) );
  AOI22_X1 U7949 ( .A1(n7040), .A2(keyinput30), .B1(keyinput91), .B2(n7039), 
        .ZN(n7038) );
  OAI221_X1 U7950 ( .B1(n7040), .B2(keyinput30), .C1(n7039), .C2(keyinput91), 
        .A(n7038), .ZN(n7046) );
  AOI22_X1 U7951 ( .A1(n4218), .A2(keyinput22), .B1(keyinput87), .B2(n4872), 
        .ZN(n7041) );
  OAI221_X1 U7952 ( .B1(n4218), .B2(keyinput22), .C1(n4872), .C2(keyinput87), 
        .A(n7041), .ZN(n7045) );
  XNOR2_X1 U7953 ( .A(EAX_REG_22__SCAN_IN), .B(keyinput117), .ZN(n7043) );
  XNOR2_X1 U7954 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .B(keyinput28), .ZN(n7042)
         );
  NAND2_X1 U7955 ( .A1(n7043), .A2(n7042), .ZN(n7044) );
  NOR4_X1 U7956 ( .A1(n7047), .A2(n7046), .A3(n7045), .A4(n7044), .ZN(n7065)
         );
  INV_X1 U7957 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n7049) );
  AOI22_X1 U7958 ( .A1(n7050), .A2(keyinput33), .B1(keyinput29), .B2(n7049), 
        .ZN(n7048) );
  OAI221_X1 U7959 ( .B1(n7050), .B2(keyinput33), .C1(n7049), .C2(keyinput29), 
        .A(n7048), .ZN(n7063) );
  INV_X1 U7960 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n7052) );
  AOI22_X1 U7961 ( .A1(n7053), .A2(keyinput17), .B1(n7052), .B2(keyinput37), 
        .ZN(n7051) );
  OAI221_X1 U7962 ( .B1(n7053), .B2(keyinput17), .C1(n7052), .C2(keyinput37), 
        .A(n7051), .ZN(n7062) );
  AOI22_X1 U7963 ( .A1(n7056), .A2(keyinput34), .B1(n7055), .B2(keyinput43), 
        .ZN(n7054) );
  OAI221_X1 U7964 ( .B1(n7056), .B2(keyinput34), .C1(n7055), .C2(keyinput43), 
        .A(n7054), .ZN(n7061) );
  INV_X1 U7965 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n7059) );
  AOI22_X1 U7966 ( .A1(n7059), .A2(keyinput51), .B1(n7058), .B2(keyinput54), 
        .ZN(n7057) );
  OAI221_X1 U7967 ( .B1(n7059), .B2(keyinput51), .C1(n7058), .C2(keyinput54), 
        .A(n7057), .ZN(n7060) );
  NOR4_X1 U7968 ( .A1(n7063), .A2(n7062), .A3(n7061), .A4(n7060), .ZN(n7064)
         );
  NAND4_X1 U7969 ( .A1(n7067), .A2(n7066), .A3(n7065), .A4(n7064), .ZN(n7143)
         );
  OAI22_X1 U7970 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(keyinput36), .B1(
        INSTQUEUE_REG_11__7__SCAN_IN), .B2(keyinput55), .ZN(n7068) );
  AOI221_X1 U7971 ( .B1(INSTQUEUE_REG_3__6__SCAN_IN), .B2(keyinput36), .C1(
        keyinput55), .C2(INSTQUEUE_REG_11__7__SCAN_IN), .A(n7068), .ZN(n7075)
         );
  OAI22_X1 U7972 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(keyinput108), .B1(
        DATAI_6_), .B2(keyinput79), .ZN(n7069) );
  AOI221_X1 U7973 ( .B1(INSTQUEUE_REG_4__0__SCAN_IN), .B2(keyinput108), .C1(
        keyinput79), .C2(DATAI_6_), .A(n7069), .ZN(n7074) );
  OAI22_X1 U7974 ( .A1(DATAI_15_), .A2(keyinput2), .B1(DATAO_REG_25__SCAN_IN), 
        .B2(keyinput71), .ZN(n7070) );
  AOI221_X1 U7975 ( .B1(DATAI_15_), .B2(keyinput2), .C1(keyinput71), .C2(
        DATAO_REG_25__SCAN_IN), .A(n7070), .ZN(n7073) );
  OAI22_X1 U7976 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(keyinput114), .B1(
        keyinput27), .B2(LWORD_REG_0__SCAN_IN), .ZN(n7071) );
  AOI221_X1 U7977 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput114), 
        .C1(LWORD_REG_0__SCAN_IN), .C2(keyinput27), .A(n7071), .ZN(n7072) );
  NAND4_X1 U7978 ( .A1(n7075), .A2(n7074), .A3(n7073), .A4(n7072), .ZN(n7103)
         );
  OAI22_X1 U7979 ( .A1(EAX_REG_17__SCAN_IN), .A2(keyinput31), .B1(keyinput82), 
        .B2(EAX_REG_19__SCAN_IN), .ZN(n7076) );
  AOI221_X1 U7980 ( .B1(EAX_REG_17__SCAN_IN), .B2(keyinput31), .C1(
        EAX_REG_19__SCAN_IN), .C2(keyinput82), .A(n7076), .ZN(n7083) );
  OAI22_X1 U7981 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(keyinput110), 
        .B1(UWORD_REG_7__SCAN_IN), .B2(keyinput60), .ZN(n7077) );
  AOI221_X1 U7982 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput110), 
        .C1(keyinput60), .C2(UWORD_REG_7__SCAN_IN), .A(n7077), .ZN(n7082) );
  OAI22_X1 U7983 ( .A1(EAX_REG_16__SCAN_IN), .A2(keyinput16), .B1(keyinput78), 
        .B2(EAX_REG_28__SCAN_IN), .ZN(n7078) );
  AOI221_X1 U7984 ( .B1(EAX_REG_16__SCAN_IN), .B2(keyinput16), .C1(
        EAX_REG_28__SCAN_IN), .C2(keyinput78), .A(n7078), .ZN(n7081) );
  OAI22_X1 U7985 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(keyinput58), .B1(
        keyinput105), .B2(EAX_REG_27__SCAN_IN), .ZN(n7079) );
  AOI221_X1 U7986 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(keyinput58), 
        .C1(EAX_REG_27__SCAN_IN), .C2(keyinput105), .A(n7079), .ZN(n7080) );
  NAND4_X1 U7987 ( .A1(n7083), .A2(n7082), .A3(n7081), .A4(n7080), .ZN(n7102)
         );
  OAI22_X1 U7988 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(keyinput49), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(keyinput97), .ZN(n7084) );
  AOI221_X1 U7989 ( .B1(INSTQUEUE_REG_14__1__SCAN_IN), .B2(keyinput49), .C1(
        keyinput97), .C2(ADDRESS_REG_27__SCAN_IN), .A(n7084), .ZN(n7091) );
  OAI22_X1 U7990 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(keyinput13), .B1(
        keyinput45), .B2(ADDRESS_REG_7__SCAN_IN), .ZN(n7085) );
  AOI221_X1 U7991 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(keyinput13), 
        .C1(ADDRESS_REG_7__SCAN_IN), .C2(keyinput45), .A(n7085), .ZN(n7090) );
  OAI22_X1 U7992 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(keyinput120), .B1(
        DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput44), .ZN(n7086) );
  AOI221_X1 U7993 ( .B1(INSTQUEUE_REG_1__5__SCAN_IN), .B2(keyinput120), .C1(
        keyinput44), .C2(DATAWIDTH_REG_23__SCAN_IN), .A(n7086), .ZN(n7089) );
  OAI22_X1 U7994 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(keyinput42), .B1(
        keyinput100), .B2(EAX_REG_10__SCAN_IN), .ZN(n7087) );
  AOI221_X1 U7995 ( .B1(INSTQUEUE_REG_3__7__SCAN_IN), .B2(keyinput42), .C1(
        EAX_REG_10__SCAN_IN), .C2(keyinput100), .A(n7087), .ZN(n7088) );
  NAND4_X1 U7996 ( .A1(n7091), .A2(n7090), .A3(n7089), .A4(n7088), .ZN(n7101)
         );
  OAI22_X1 U7997 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(keyinput39), .B1(
        keyinput115), .B2(DATAWIDTH_REG_25__SCAN_IN), .ZN(n7092) );
  AOI221_X1 U7998 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(keyinput39), .C1(
        DATAWIDTH_REG_25__SCAN_IN), .C2(keyinput115), .A(n7092), .ZN(n7099) );
  OAI22_X1 U7999 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(keyinput61), .B1(
        keyinput48), .B2(REIP_REG_5__SCAN_IN), .ZN(n7093) );
  AOI221_X1 U8000 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput61), .C1(
        REIP_REG_5__SCAN_IN), .C2(keyinput48), .A(n7093), .ZN(n7098) );
  OAI22_X1 U8001 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(keyinput126), .B1(
        EAX_REG_12__SCAN_IN), .B2(keyinput6), .ZN(n7094) );
  AOI221_X1 U8002 ( .B1(INSTQUEUE_REG_2__2__SCAN_IN), .B2(keyinput126), .C1(
        keyinput6), .C2(EAX_REG_12__SCAN_IN), .A(n7094), .ZN(n7097) );
  OAI22_X1 U8003 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(keyinput77), .B1(
        keyinput21), .B2(ADDRESS_REG_23__SCAN_IN), .ZN(n7095) );
  AOI221_X1 U8004 ( .B1(INSTQUEUE_REG_5__6__SCAN_IN), .B2(keyinput77), .C1(
        ADDRESS_REG_23__SCAN_IN), .C2(keyinput21), .A(n7095), .ZN(n7096) );
  NAND4_X1 U8005 ( .A1(n7099), .A2(n7098), .A3(n7097), .A4(n7096), .ZN(n7100)
         );
  NOR4_X1 U8006 ( .A1(n7103), .A2(n7102), .A3(n7101), .A4(n7100), .ZN(n7141)
         );
  OAI22_X1 U8007 ( .A1(EBX_REG_18__SCAN_IN), .A2(keyinput104), .B1(keyinput53), 
        .B2(DATAWIDTH_REG_27__SCAN_IN), .ZN(n7104) );
  AOI221_X1 U8008 ( .B1(EBX_REG_18__SCAN_IN), .B2(keyinput104), .C1(
        DATAWIDTH_REG_27__SCAN_IN), .C2(keyinput53), .A(n7104), .ZN(n7111) );
  OAI22_X1 U8009 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(keyinput93), .B1(
        keyinput116), .B2(EAX_REG_3__SCAN_IN), .ZN(n7105) );
  AOI221_X1 U8010 ( .B1(INSTQUEUE_REG_8__0__SCAN_IN), .B2(keyinput93), .C1(
        EAX_REG_3__SCAN_IN), .C2(keyinput116), .A(n7105), .ZN(n7110) );
  OAI22_X1 U8011 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(keyinput20), .B1(
        INSTADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput119), .ZN(n7106) );
  AOI221_X1 U8012 ( .B1(INSTQUEUE_REG_12__6__SCAN_IN), .B2(keyinput20), .C1(
        keyinput119), .C2(INSTADDRPOINTER_REG_14__SCAN_IN), .A(n7106), .ZN(
        n7109) );
  OAI22_X1 U8013 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(keyinput59), .B1(
        keyinput72), .B2(DATAI_22_), .ZN(n7107) );
  AOI221_X1 U8014 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(keyinput59), .C1(
        DATAI_22_), .C2(keyinput72), .A(n7107), .ZN(n7108) );
  NAND4_X1 U8015 ( .A1(n7111), .A2(n7110), .A3(n7109), .A4(n7108), .ZN(n7139)
         );
  OAI22_X1 U8016 ( .A1(DATAO_REG_16__SCAN_IN), .A2(keyinput68), .B1(keyinput10), .B2(LWORD_REG_1__SCAN_IN), .ZN(n7112) );
  AOI221_X1 U8017 ( .B1(DATAO_REG_16__SCAN_IN), .B2(keyinput68), .C1(
        LWORD_REG_1__SCAN_IN), .C2(keyinput10), .A(n7112), .ZN(n7119) );
  OAI22_X1 U8018 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(keyinput99), .B1(
        REIP_REG_12__SCAN_IN), .B2(keyinput70), .ZN(n7113) );
  AOI221_X1 U8019 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput99), 
        .C1(keyinput70), .C2(REIP_REG_12__SCAN_IN), .A(n7113), .ZN(n7118) );
  OAI22_X1 U8020 ( .A1(LWORD_REG_5__SCAN_IN), .A2(keyinput35), .B1(keyinput85), 
        .B2(ADDRESS_REG_21__SCAN_IN), .ZN(n7114) );
  AOI221_X1 U8021 ( .B1(LWORD_REG_5__SCAN_IN), .B2(keyinput35), .C1(
        ADDRESS_REG_21__SCAN_IN), .C2(keyinput85), .A(n7114), .ZN(n7117) );
  OAI22_X1 U8022 ( .A1(EBX_REG_9__SCAN_IN), .A2(keyinput69), .B1(keyinput63), 
        .B2(BE_N_REG_0__SCAN_IN), .ZN(n7115) );
  AOI221_X1 U8023 ( .B1(EBX_REG_9__SCAN_IN), .B2(keyinput69), .C1(
        BE_N_REG_0__SCAN_IN), .C2(keyinput63), .A(n7115), .ZN(n7116) );
  NAND4_X1 U8024 ( .A1(n7119), .A2(n7118), .A3(n7117), .A4(n7116), .ZN(n7138)
         );
  OAI22_X1 U8025 ( .A1(LWORD_REG_11__SCAN_IN), .A2(keyinput18), .B1(
        ADS_N_REG_SCAN_IN), .B2(keyinput57), .ZN(n7120) );
  AOI221_X1 U8026 ( .B1(LWORD_REG_11__SCAN_IN), .B2(keyinput18), .C1(
        keyinput57), .C2(ADS_N_REG_SCAN_IN), .A(n7120), .ZN(n7127) );
  OAI22_X1 U8027 ( .A1(DATAO_REG_27__SCAN_IN), .A2(keyinput127), .B1(
        DATAO_REG_31__SCAN_IN), .B2(keyinput92), .ZN(n7121) );
  AOI221_X1 U8028 ( .B1(DATAO_REG_27__SCAN_IN), .B2(keyinput127), .C1(
        keyinput92), .C2(DATAO_REG_31__SCAN_IN), .A(n7121), .ZN(n7126) );
  OAI22_X1 U8029 ( .A1(EBX_REG_23__SCAN_IN), .A2(keyinput32), .B1(
        DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput47), .ZN(n7122) );
  AOI221_X1 U8030 ( .B1(EBX_REG_23__SCAN_IN), .B2(keyinput32), .C1(keyinput47), 
        .C2(DATAWIDTH_REG_5__SCAN_IN), .A(n7122), .ZN(n7125) );
  OAI22_X1 U8031 ( .A1(EAX_REG_13__SCAN_IN), .A2(keyinput94), .B1(keyinput15), 
        .B2(NA_N), .ZN(n7123) );
  AOI221_X1 U8032 ( .B1(EAX_REG_13__SCAN_IN), .B2(keyinput94), .C1(NA_N), .C2(
        keyinput15), .A(n7123), .ZN(n7124) );
  NAND4_X1 U8033 ( .A1(n7127), .A2(n7126), .A3(n7125), .A4(n7124), .ZN(n7137)
         );
  OAI22_X1 U8034 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput7), .B1(
        keyinput107), .B2(REIP_REG_18__SCAN_IN), .ZN(n7128) );
  AOI221_X1 U8035 ( .B1(PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput7), .C1(
        REIP_REG_18__SCAN_IN), .C2(keyinput107), .A(n7128), .ZN(n7135) );
  OAI22_X1 U8036 ( .A1(EBX_REG_30__SCAN_IN), .A2(keyinput40), .B1(keyinput89), 
        .B2(UWORD_REG_4__SCAN_IN), .ZN(n7129) );
  AOI221_X1 U8037 ( .B1(EBX_REG_30__SCAN_IN), .B2(keyinput40), .C1(
        UWORD_REG_4__SCAN_IN), .C2(keyinput89), .A(n7129), .ZN(n7134) );
  OAI22_X1 U8038 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(keyinput96), .B1(
        keyinput123), .B2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n7130) );
  AOI221_X1 U8039 ( .B1(INSTQUEUE_REG_9__1__SCAN_IN), .B2(keyinput96), .C1(
        INSTADDRPOINTER_REG_5__SCAN_IN), .C2(keyinput123), .A(n7130), .ZN(
        n7133) );
  OAI22_X1 U8040 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(keyinput111), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(keyinput102), .ZN(n7131) );
  AOI221_X1 U8041 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(keyinput111), .C1(
        keyinput102), .C2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n7131), .ZN(n7132) );
  NAND4_X1 U8042 ( .A1(n7135), .A2(n7134), .A3(n7133), .A4(n7132), .ZN(n7136)
         );
  NOR4_X1 U8043 ( .A1(n7139), .A2(n7138), .A3(n7137), .A4(n7136), .ZN(n7140)
         );
  NAND2_X1 U8044 ( .A1(n7141), .A2(n7140), .ZN(n7142) );
  NOR4_X1 U8045 ( .A1(n7145), .A2(n7144), .A3(n7143), .A4(n7142), .ZN(n7150)
         );
  AOI222_X1 U8046 ( .A1(n7148), .A2(ADDRESS_REG_26__SCAN_IN), .B1(
        REIP_REG_27__SCAN_IN), .B2(n7147), .C1(REIP_REG_28__SCAN_IN), .C2(
        n7146), .ZN(n7149) );
  XNOR2_X1 U8047 ( .A(n7150), .B(n7149), .ZN(U3210) );
  CLKBUF_X1 U3643 ( .A(n3536), .Z(n3577) );
  CLKBUF_X3 U3688 ( .A(n3406), .Z(n4603) );
  CLKBUF_X1 U3865 ( .A(n4522), .Z(n3172) );
endmodule

