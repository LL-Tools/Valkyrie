

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8854, n8855, n8856, n8857,
         n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
         n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877,
         n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887,
         n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897,
         n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907,
         n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917,
         n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927,
         n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937,
         n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947,
         n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957,
         n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967,
         n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977,
         n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987,
         n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997,
         n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
         n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
         n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
         n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
         n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
         n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
         n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
         n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
         n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
         n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
         n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
         n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
         n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
         n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
         n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
         n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
         n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
         n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
         n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
         n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
         n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
         n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
         n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
         n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
         n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
         n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
         n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
         n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
         n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
         n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647,
         n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657,
         n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667,
         n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677,
         n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687,
         n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697,
         n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707,
         n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717,
         n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919;

  AND2_X1 U4752 ( .A1(n9580), .A2(n4475), .ZN(n7381) );
  CLKBUF_X2 U4753 ( .A(n5789), .Z(n6043) );
  INV_X1 U4754 ( .A(n5590), .ZN(n5894) );
  CLKBUF_X2 U4755 ( .A(n5060), .Z(n5348) );
  AND4_X1 U4756 ( .A1(n4885), .A2(n4884), .A3(n4883), .A4(n4882), .ZN(n6485)
         );
  INV_X1 U4757 ( .A(n5574), .ZN(n6057) );
  CLKBUF_X2 U4758 ( .A(n4974), .Z(n4253) );
  CLKBUF_X2 U4759 ( .A(n4881), .Z(n4251) );
  CLKBUF_X2 U4760 ( .A(n4881), .Z(n4250) );
  AND2_X1 U4761 ( .A1(n8850), .A2(n4812), .ZN(n4881) );
  XNOR2_X1 U4762 ( .A(n5446), .B(n4834), .ZN(n6366) );
  INV_X1 U4763 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5535) );
  INV_X1 U4764 ( .A(n8274), .ZN(n8267) );
  AND2_X1 U4767 ( .A1(n9579), .A2(n9578), .ZN(n9580) );
  OR2_X2 U4768 ( .A1(n6160), .A2(n6125), .ZN(n6055) );
  INV_X1 U4769 ( .A(n6870), .ZN(n5983) );
  NOR2_X1 U4770 ( .A1(n9206), .A2(n9296), .ZN(n9191) );
  AOI21_X1 U4771 ( .B1(n7274), .B2(n4503), .A(n4502), .ZN(n4501) );
  INV_X1 U4772 ( .A(n4251), .ZN(n5276) );
  BUF_X1 U4773 ( .A(n4265), .Z(n4248) );
  INV_X1 U4774 ( .A(n4864), .ZN(n8567) );
  AND3_X1 U4775 ( .A1(n4954), .A2(n4953), .A3(n4952), .ZN(n6778) );
  INV_X1 U4776 ( .A(n6480), .ZN(n9640) );
  INV_X2 U4777 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8845) );
  INV_X1 U4778 ( .A(n5736), .ZN(n6025) );
  AND4_X1 U4779 ( .A1(n4943), .A2(n4942), .A3(n4941), .A4(n4940), .ZN(n8696)
         );
  NAND2_X1 U4780 ( .A1(n8588), .A2(n8590), .ZN(n8587) );
  NAND2_X1 U4781 ( .A1(n7110), .A2(n8300), .ZN(n8818) );
  OAI211_X1 U4782 ( .C1(n4944), .C2(n6203), .A(n4896), .B(n4895), .ZN(n6450)
         );
  INV_X1 U4783 ( .A(n4822), .ZN(n8850) );
  NOR2_X1 U4784 ( .A1(n4894), .A2(n4797), .ZN(n7310) );
  AND4_X1 U4785 ( .A1(n5602), .A2(n5601), .A3(n5600), .A4(n5599), .ZN(n6832)
         );
  NAND2_X1 U4786 ( .A1(n5551), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5536) );
  INV_X1 U4787 ( .A(n6163), .ZN(n9527) );
  BUF_X1 U4788 ( .A(n6131), .Z(n8976) );
  XNOR2_X1 U4789 ( .A(n5536), .B(n5535), .ZN(n7777) );
  INV_X1 U4790 ( .A(n5641), .ZN(n5744) );
  AOI21_X2 U4791 ( .B1(n6817), .B2(n5659), .A(n4786), .ZN(n6889) );
  AND2_X2 U4792 ( .A1(n5523), .A2(n9367), .ZN(n5598) );
  XNOR2_X2 U4793 ( .A(n5195), .B(n5220), .ZN(n6566) );
  AND2_X4 U4794 ( .A1(n5524), .A2(n8331), .ZN(n5641) );
  NAND2_X2 U4795 ( .A1(n5521), .A2(n9362), .ZN(n8331) );
  AOI21_X2 U4796 ( .B1(n9054), .B2(n9053), .A(n9052), .ZN(n9231) );
  OAI22_X2 U4797 ( .A1(n7502), .A2(n7501), .B1(n7521), .B2(n7548), .ZN(n9054)
         );
  NOR2_X2 U4798 ( .A1(n5515), .A2(n5514), .ZN(n5516) );
  NOR2_X2 U4799 ( .A1(n4338), .A2(n4340), .ZN(n5452) );
  OAI22_X1 U4801 ( .A1(n8577), .A2(n4325), .B1(n4254), .B2(n4328), .ZN(n8528)
         );
  NAND2_X1 U4802 ( .A1(n4346), .A2(n4344), .ZN(n7424) );
  AND2_X1 U4803 ( .A1(n4523), .A2(n4322), .ZN(n7196) );
  NAND2_X1 U4804 ( .A1(n6746), .A2(n6745), .ZN(n6744) );
  NAND2_X2 U4805 ( .A1(n8970), .A2(n9533), .ZN(n7621) );
  NOR2_X1 U4806 ( .A1(n6653), .A2(n4977), .ZN(n4499) );
  AND2_X1 U4807 ( .A1(n4872), .A2(n4880), .ZN(n6453) );
  INV_X1 U4808 ( .A(n9519), .ZN(n6135) );
  AND2_X1 U4809 ( .A1(n8152), .A2(n8132), .ZN(n8146) );
  INV_X1 U4810 ( .A(n7704), .ZN(n7708) );
  OR2_X1 U4811 ( .A1(n5276), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n4901) );
  INV_X1 U4812 ( .A(n6832), .ZN(n8974) );
  CLKBUF_X2 U4813 ( .A(n4886), .Z(n6421) );
  AND2_X2 U4814 ( .A1(n4878), .A2(n7577), .ZN(n4974) );
  INV_X2 U4815 ( .A(n8315), .ZN(n8114) );
  INV_X2 U4816 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NAND2_X1 U4817 ( .A1(n5989), .A2(n5988), .ZN(n8895) );
  CLKBUF_X1 U4818 ( .A(n8380), .Z(n8381) );
  NOR2_X1 U4819 ( .A1(n8528), .A2(n8257), .ZN(n8506) );
  NAND2_X1 U4820 ( .A1(n7272), .A2(n4505), .ZN(n4504) );
  NAND2_X1 U4821 ( .A1(n5991), .A2(n5990), .ZN(n9279) );
  INV_X1 U4822 ( .A(n9166), .ZN(n9285) );
  AND2_X1 U4823 ( .A1(n5974), .A2(n5973), .ZN(n9166) );
  OR2_X1 U4824 ( .A1(n9217), .A2(n9303), .ZN(n9206) );
  NAND2_X1 U4825 ( .A1(n7424), .A2(n4613), .ZN(n4618) );
  NOR2_X1 U4826 ( .A1(n4507), .A2(n4506), .ZN(n4505) );
  OR2_X1 U4827 ( .A1(n7301), .A2(n4345), .ZN(n4344) );
  NAND2_X1 U4828 ( .A1(n5859), .A2(n5858), .ZN(n9323) );
  OR2_X1 U4829 ( .A1(n9421), .A2(n9416), .ZN(n9422) );
  AND2_X1 U4830 ( .A1(n6977), .A2(n4332), .ZN(n9565) );
  NAND2_X1 U4831 ( .A1(n6777), .A2(n8291), .ZN(n6799) );
  NAND2_X1 U4832 ( .A1(n5125), .A2(n5124), .ZN(n8820) );
  AND2_X1 U4833 ( .A1(n7619), .A2(n7621), .ZN(n7803) );
  AOI21_X1 U4834 ( .B1(n8688), .B2(n6785), .A(n4792), .ZN(n8691) );
  AND2_X1 U4835 ( .A1(n8170), .A2(n8169), .ZN(n8294) );
  NAND2_X1 U4836 ( .A1(n5147), .A2(n5146), .ZN(n5161) );
  NAND2_X1 U4837 ( .A1(n5699), .A2(n5698), .ZN(n7075) );
  NOR2_X1 U4838 ( .A1(n8709), .A2(n4777), .ZN(n4776) );
  INV_X1 U4839 ( .A(n8290), .ZN(n8709) );
  NAND2_X1 U4840 ( .A1(n5596), .A2(n5595), .ZN(n6605) );
  NAND2_X1 U4841 ( .A1(n8160), .A2(n8156), .ZN(n8290) );
  INV_X2 U4842 ( .A(n8699), .ZN(n9588) );
  NAND2_X1 U4843 ( .A1(n8700), .A2(n8436), .ZN(n8156) );
  AND2_X1 U4844 ( .A1(n6537), .A2(n9640), .ZN(n6779) );
  NAND2_X1 U4845 ( .A1(n4612), .A2(n4610), .ZN(n9649) );
  NOR2_X1 U4846 ( .A1(n6538), .A2(n8720), .ZN(n6537) );
  NAND2_X1 U4847 ( .A1(n4429), .A2(n7834), .ZN(n7747) );
  OAI211_X1 U4848 ( .C1(n5736), .C2(n9867), .A(n5650), .B(n5649), .ZN(n9519)
         );
  NAND2_X1 U4849 ( .A1(n4973), .A2(n4972), .ZN(n4987) );
  BUF_X1 U4850 ( .A(n6367), .Z(n6457) );
  OAI211_X1 U4851 ( .C1(n4944), .C2(n6210), .A(n4917), .B(n4916), .ZN(n8720)
         );
  AND4_X1 U4852 ( .A1(n4923), .A2(n4922), .A3(n4921), .A4(n4920), .ZN(n6628)
         );
  AND4_X1 U4853 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n6788)
         );
  AND4_X1 U4854 ( .A1(n4984), .A2(n4983), .A3(n4982), .A4(n4981), .ZN(n8694)
         );
  AND4_X1 U4855 ( .A1(n5003), .A2(n5002), .A3(n5001), .A4(n5000), .ZN(n6966)
         );
  NAND2_X1 U4856 ( .A1(n4950), .A2(n4949), .ZN(n4970) );
  NAND2_X1 U4857 ( .A1(n4929), .A2(n4928), .ZN(n4946) );
  AND4_X1 U4858 ( .A1(n5615), .A2(n5614), .A3(n5613), .A4(n5612), .ZN(n6950)
         );
  BUF_X2 U4859 ( .A(n4974), .Z(n4252) );
  NAND2_X2 U4860 ( .A1(n6160), .A2(n6092), .ZN(n5574) );
  AND2_X2 U4861 ( .A1(n4822), .A2(n4812), .ZN(n4265) );
  BUF_X4 U4862 ( .A(n4900), .Z(n5418) );
  NAND2_X1 U4863 ( .A1(n4878), .A2(n6196), .ZN(n4944) );
  AND2_X2 U4864 ( .A1(n8850), .A2(n8854), .ZN(n4900) );
  NAND2_X1 U4865 ( .A1(n4811), .A2(n8846), .ZN(n8854) );
  BUF_X4 U4866 ( .A(n5598), .Z(n4247) );
  NAND2_X1 U4867 ( .A1(n4833), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5446) );
  XNOR2_X1 U4868 ( .A(n4807), .B(n4806), .ZN(n4822) );
  XNOR2_X1 U4869 ( .A(n4830), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8315) );
  XNOR2_X1 U4870 ( .A(n4843), .B(n4842), .ZN(n4864) );
  XNOR2_X1 U4871 ( .A(n5522), .B(P1_IR_REG_30__SCAN_IN), .ZN(n9367) );
  OR2_X1 U4872 ( .A1(n4810), .A2(n8845), .ZN(n4807) );
  MUX2_X1 U4873 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5520), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5521) );
  NAND2_X1 U4874 ( .A1(n9362), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5522) );
  NAND2_X2 U4875 ( .A1(n7577), .A2(P1_U3084), .ZN(n8334) );
  NOR2_X1 U4876 ( .A1(n7577), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9366) );
  OR2_X1 U4877 ( .A1(n5560), .A2(n5519), .ZN(n5520) );
  NOR2_X1 U4878 ( .A1(n5226), .A2(n4828), .ZN(n4835) );
  INV_X4 U4879 ( .A(n6196), .ZN(n7577) );
  NAND2_X1 U4880 ( .A1(n5758), .A2(n4609), .ZN(n5829) );
  AND2_X1 U4881 ( .A1(n4803), .A2(n4797), .ZN(n4342) );
  AND2_X1 U4882 ( .A1(n4753), .A2(n4341), .ZN(n4337) );
  AND2_X1 U4883 ( .A1(n4796), .A2(n4798), .ZN(n4753) );
  INV_X1 U4884 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5095) );
  NOR2_X1 U4885 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5512) );
  INV_X1 U4886 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5094) );
  INV_X1 U4887 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5121) );
  INV_X1 U4888 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5148) );
  INV_X1 U4889 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5166) );
  NOR2_X1 U4890 ( .A1(P1_RD_REG_SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n4855) );
  INV_X1 U4891 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5808) );
  INV_X1 U4892 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5506) );
  INV_X1 U4893 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5670) );
  INV_X4 U4894 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4895 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4667) );
  INV_X1 U4896 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4796) );
  XNOR2_X2 U4897 ( .A(n5318), .B(n5319), .ZN(n8401) );
  NAND2_X2 U4898 ( .A1(n8363), .A2(n5298), .ZN(n5318) );
  OAI21_X2 U4899 ( .B1(n8880), .B2(n8881), .A(n5907), .ZN(n8909) );
  INV_X1 U4900 ( .A(n5574), .ZN(n4249) );
  INV_X2 U4901 ( .A(n4878), .ZN(n4912) );
  NAND2_X2 U4902 ( .A1(n7269), .A2(n5492), .ZN(n4878) );
  INV_X1 U4903 ( .A(n5179), .ZN(n4557) );
  INV_X1 U4904 ( .A(n8854), .ZN(n4812) );
  OR2_X1 U4905 ( .A1(n8741), .A2(n8423), .ZN(n8488) );
  INV_X1 U4906 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4341) );
  INV_X1 U4907 ( .A(n4706), .ZN(n4415) );
  AND2_X1 U4908 ( .A1(n9043), .A2(n9041), .ZN(n7779) );
  OAI21_X1 U4909 ( .B1(n5264), .B2(n5263), .A(n5262), .ZN(n5285) );
  NAND2_X1 U4910 ( .A1(n5113), .A2(n5092), .ZN(n5114) );
  OAI21_X1 U4911 ( .B1(n5044), .B2(n5043), .A(n4293), .ZN(n5069) );
  OR2_X1 U4912 ( .A1(n5042), .A2(n5046), .ZN(n5043) );
  OR2_X1 U4913 ( .A1(n5046), .A2(n5045), .ZN(n5047) );
  NAND2_X1 U4914 ( .A1(n8462), .A2(n8573), .ZN(n8562) );
  INV_X1 U4915 ( .A(n4733), .ZN(n8588) );
  NAND2_X1 U4916 ( .A1(n4737), .A2(n8483), .ZN(n4736) );
  INV_X1 U4917 ( .A(n4735), .ZN(n4734) );
  NAND3_X1 U4918 ( .A1(n4618), .A2(n4614), .A3(n8101), .ZN(n8660) );
  NAND2_X1 U4919 ( .A1(n4638), .A2(n8189), .ZN(n4637) );
  NOR2_X1 U4920 ( .A1(n4642), .A2(n4648), .ZN(n4640) );
  AOI21_X1 U4921 ( .B1(n4776), .B2(n4774), .A(n4291), .ZN(n4773) );
  INV_X1 U4922 ( .A(n4776), .ZN(n4775) );
  BUF_X1 U4923 ( .A(n5721), .Z(n7588) );
  AND2_X1 U4924 ( .A1(n9367), .A2(n8331), .ZN(n5721) );
  OAI21_X1 U4925 ( .B1(n7659), .B2(n7719), .A(n7718), .ZN(n7661) );
  NAND2_X1 U4926 ( .A1(n6488), .A2(n8720), .ZN(n8132) );
  NAND2_X1 U4927 ( .A1(n5031), .A2(n5030), .ZN(n5048) );
  NOR2_X1 U4928 ( .A1(n8741), .A2(n8746), .ZN(n4474) );
  AND2_X1 U4929 ( .A1(n8792), .A2(n8475), .ZN(n8222) );
  AOI21_X1 U4930 ( .B1(n4766), .B2(n4762), .A(n4292), .ZN(n4761) );
  NAND2_X1 U4931 ( .A1(n4636), .A2(n8188), .ZN(n4638) );
  OR2_X1 U4932 ( .A1(n5103), .A2(n4818), .ZN(n5127) );
  INV_X1 U4933 ( .A(n4342), .ZN(n4338) );
  OR2_X1 U4934 ( .A1(n9258), .A2(n9105), .ZN(n7781) );
  OR2_X1 U4935 ( .A1(n9269), .A2(n9135), .ZN(n9079) );
  OR2_X1 U4936 ( .A1(n9275), .A2(n9121), .ZN(n9077) );
  NAND2_X1 U4937 ( .A1(n9195), .A2(n9205), .ZN(n4691) );
  OAI21_X1 U4938 ( .B1(n4436), .B2(n7470), .A(n4434), .ZN(n4433) );
  AND2_X1 U4939 ( .A1(n7411), .A2(n4712), .ZN(n4710) );
  OR2_X1 U4940 ( .A1(n9331), .A2(n8965), .ZN(n7411) );
  XNOR2_X1 U4941 ( .A(n7579), .B(n7578), .ZN(n7585) );
  OAI21_X1 U4942 ( .B1(n5324), .B2(n5323), .A(n5322), .ZN(n5332) );
  NAND2_X1 U4943 ( .A1(n5244), .A2(n5243), .ZN(n5264) );
  NAND2_X1 U4944 ( .A1(n4550), .A2(n4549), .ZN(n5244) );
  AOI21_X1 U4945 ( .B1(n4551), .B2(n4552), .A(n5240), .ZN(n4549) );
  NAND2_X1 U4946 ( .A1(n4553), .A2(n4556), .ZN(n5225) );
  NAND2_X1 U4947 ( .A1(n5161), .A2(n4558), .ZN(n4553) );
  NAND2_X1 U4948 ( .A1(n5179), .A2(n5165), .ZN(n5180) );
  NAND2_X1 U4949 ( .A1(n5085), .A2(SI_11_), .ZN(n5086) );
  NAND2_X1 U4950 ( .A1(n5069), .A2(n4785), .ZN(n5071) );
  NAND2_X1 U4951 ( .A1(n5012), .A2(n5011), .ZN(n5045) );
  NAND2_X1 U4952 ( .A1(n5009), .A2(n5008), .ZN(n5044) );
  NAND2_X1 U4953 ( .A1(n4524), .A2(n7078), .ZN(n4523) );
  INV_X1 U4954 ( .A(n4323), .ZN(n4322) );
  INV_X1 U4955 ( .A(n4527), .ZN(n4524) );
  NAND2_X1 U4956 ( .A1(n8470), .A2(n8115), .ZN(n4655) );
  AOI21_X1 U4957 ( .B1(n4658), .B2(n8510), .A(n4657), .ZN(n4656) );
  INV_X1 U4958 ( .A(n8269), .ZN(n4657) );
  NOR2_X1 U4959 ( .A1(n4661), .A2(n8115), .ZN(n4654) );
  AND4_X1 U4960 ( .A1(n5211), .A2(n5210), .A3(n5209), .A4(n5208), .ZN(n7425)
         );
  OR2_X1 U4961 ( .A1(n8746), .A2(n8549), .ZN(n8487) );
  AND2_X1 U4962 ( .A1(n8510), .A2(n4731), .ZN(n4730) );
  OR2_X1 U4963 ( .A1(n8530), .A2(n4732), .ZN(n4731) );
  OR2_X1 U4964 ( .A1(n4254), .A2(n8556), .ZN(n4325) );
  OR2_X1 U4965 ( .A1(n8752), .A2(n8486), .ZN(n4324) );
  NAND2_X1 U4966 ( .A1(n8239), .A2(n8237), .ZN(n8590) );
  NOR2_X1 U4967 ( .A1(n8788), .A2(n8681), .ZN(n8478) );
  OR2_X1 U4968 ( .A1(n4348), .A2(n7395), .ZN(n4346) );
  OR2_X1 U4969 ( .A1(n7295), .A2(n7302), .ZN(n4782) );
  NAND2_X1 U4970 ( .A1(n5100), .A2(n5099), .ZN(n7107) );
  NAND2_X1 U4971 ( .A1(n8291), .A2(n8164), .ZN(n4336) );
  NAND2_X1 U4972 ( .A1(n6775), .A2(n4269), .ZN(n4778) );
  INV_X1 U4973 ( .A(n4771), .ZN(n4769) );
  AND2_X1 U4974 ( .A1(n5562), .A2(n5561), .ZN(n5571) );
  XNOR2_X1 U4975 ( .A(n6283), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6302) );
  NAND2_X1 U4976 ( .A1(n9081), .A2(n7770), .ZN(n9103) );
  NAND2_X1 U4977 ( .A1(n7783), .A2(n9075), .ZN(n9148) );
  NAND2_X1 U4978 ( .A1(n9058), .A2(n4783), .ZN(n9198) );
  OR2_X1 U4979 ( .A1(n9306), .A2(n9242), .ZN(n9057) );
  AND2_X1 U4980 ( .A1(n9339), .A2(n8966), .ZN(n7409) );
  NAND2_X1 U4981 ( .A1(n7228), .A2(n4781), .ZN(n7410) );
  NAND2_X1 U4982 ( .A1(n7875), .A2(n9033), .ZN(n4607) );
  XNOR2_X1 U4983 ( .A(n5181), .B(n5180), .ZN(n6562) );
  OAI21_X1 U4984 ( .B1(n5161), .B2(n5160), .A(n5159), .ZN(n5181) );
  NAND2_X1 U4985 ( .A1(n5347), .A2(n5346), .ZN(n8761) );
  INV_X1 U4986 ( .A(n4326), .ZN(n8547) );
  AOI22_X1 U4987 ( .A1(n8577), .A2(n4327), .B1(n8556), .B2(n4331), .ZN(n4326)
         );
  NAND2_X1 U4988 ( .A1(n6212), .A2(n8116), .ZN(n4612) );
  NOR2_X1 U4989 ( .A1(n4277), .A2(n4611), .ZN(n4610) );
  NOR2_X1 U4990 ( .A1(n4878), .A2(n7985), .ZN(n4611) );
  AND4_X1 U4991 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), .ZN(n9161)
         );
  OAI211_X1 U4992 ( .C1(n4361), .C2(n4321), .A(n4360), .B(n4356), .ZN(n4355)
         );
  NOR2_X1 U4993 ( .A1(n7872), .A2(n7871), .ZN(n4360) );
  NAND2_X1 U4994 ( .A1(n4361), .A2(n4357), .ZN(n4356) );
  AND2_X1 U4995 ( .A1(n7653), .A2(n7652), .ZN(n4372) );
  NAND2_X1 U4996 ( .A1(n7648), .A2(n7649), .ZN(n4373) );
  NOR2_X1 U4997 ( .A1(n8346), .A2(n8345), .ZN(n4484) );
  NOR2_X1 U4998 ( .A1(n4484), .A2(n4483), .ZN(n4482) );
  INV_X1 U4999 ( .A(n8402), .ZN(n4483) );
  NAND2_X1 U5000 ( .A1(n5321), .A2(n4485), .ZN(n4480) );
  NAND2_X1 U5001 ( .A1(n8346), .A2(n8345), .ZN(n4485) );
  NAND2_X1 U5002 ( .A1(n7692), .A2(n7691), .ZN(n4378) );
  INV_X1 U5003 ( .A(n5407), .ZN(n4571) );
  INV_X1 U5004 ( .A(n4558), .ZN(n4555) );
  NOR2_X1 U5005 ( .A1(n5180), .A2(n4559), .ZN(n4558) );
  INV_X1 U5006 ( .A(n5159), .ZN(n4559) );
  INV_X1 U5007 ( .A(n5144), .ZN(n4540) );
  NAND2_X1 U5008 ( .A1(n4664), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4668) );
  INV_X1 U5009 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4664) );
  NAND2_X1 U5010 ( .A1(n4496), .A2(n4497), .ZN(n4495) );
  INV_X1 U5011 ( .A(n4499), .ZN(n4496) );
  OR2_X1 U5012 ( .A1(n8727), .A2(n8465), .ZN(n8273) );
  NAND2_X1 U5013 ( .A1(n4663), .A2(n8423), .ZN(n4662) );
  OR2_X1 U5014 ( .A1(n8499), .A2(n8110), .ZN(n8268) );
  INV_X1 U5015 ( .A(n8244), .ZN(n4329) );
  NOR2_X1 U5016 ( .A1(n8578), .A2(n4752), .ZN(n4751) );
  INV_X1 U5017 ( .A(n4790), .ZN(n4752) );
  NAND2_X1 U5018 ( .A1(n4632), .A2(n4630), .ZN(n4629) );
  INV_X1 U5019 ( .A(n8590), .ZN(n4630) );
  INV_X1 U5020 ( .A(n8105), .ZN(n4635) );
  NOR2_X1 U5021 ( .A1(n8783), .A2(n8788), .ZN(n4469) );
  NOR2_X1 U5022 ( .A1(n8301), .A2(n4765), .ZN(n4764) );
  INV_X1 U5023 ( .A(n4782), .ZN(n4765) );
  AND2_X1 U5024 ( .A1(n4477), .A2(n7295), .ZN(n4476) );
  NOR2_X1 U5025 ( .A1(n7084), .A2(n7107), .ZN(n4477) );
  NAND2_X1 U5026 ( .A1(n4723), .A2(n6798), .ZN(n4722) );
  INV_X1 U5027 ( .A(n6968), .ZN(n4723) );
  INV_X1 U5028 ( .A(n9567), .ZN(n4725) );
  NAND2_X1 U5029 ( .A1(n6471), .A2(n8146), .ZN(n6532) );
  NOR2_X1 U5030 ( .A1(n4771), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4770) );
  NAND2_X1 U5031 ( .A1(n4804), .A2(n4772), .ZN(n4771) );
  INV_X1 U5032 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4772) );
  NOR2_X1 U5033 ( .A1(n6913), .A2(n4407), .ZN(n7173) );
  AND2_X1 U5034 ( .A1(n6914), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4407) );
  INV_X1 U5035 ( .A(n6092), .ZN(n6125) );
  NAND2_X1 U5036 ( .A1(n9100), .A2(n9116), .ZN(n4427) );
  INV_X1 U5037 ( .A(n9133), .ZN(n4458) );
  INV_X1 U5038 ( .A(n9187), .ZN(n4449) );
  NOR2_X1 U5039 ( .A1(n9201), .A2(n4448), .ZN(n4447) );
  INV_X1 U5040 ( .A(n9069), .ZN(n4448) );
  OR2_X1 U5041 ( .A1(n9303), .A2(n9189), .ZN(n7787) );
  OR2_X1 U5042 ( .A1(n9416), .A2(n7210), .ZN(n7634) );
  NAND2_X1 U5043 ( .A1(n4421), .A2(n9398), .ZN(n4420) );
  NOR2_X1 U5044 ( .A1(n7075), .A2(n6999), .ZN(n4421) );
  AND2_X1 U5045 ( .A1(n7739), .A2(n7836), .ZN(n7795) );
  NAND2_X1 U5046 ( .A1(n9191), .A2(n9182), .ZN(n9176) );
  NAND2_X1 U5047 ( .A1(n5518), .A2(n4707), .ZN(n4706) );
  INV_X1 U5048 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4707) );
  NAND2_X1 U5049 ( .A1(n4561), .A2(n4560), .ZN(n7694) );
  AOI21_X1 U5050 ( .B1(n4563), .B2(n4565), .A(n4318), .ZN(n4560) );
  NAND2_X1 U5051 ( .A1(n5429), .A2(n4563), .ZN(n4561) );
  NOR2_X1 U5052 ( .A1(n5362), .A2(n4579), .ZN(n4578) );
  INV_X1 U5053 ( .A(n5344), .ZN(n4579) );
  NAND2_X1 U5054 ( .A1(n5332), .A2(n5331), .ZN(n5345) );
  NAND2_X1 U5055 ( .A1(n5304), .A2(n5303), .ZN(n5324) );
  NAND2_X1 U5056 ( .A1(n4546), .A2(n5086), .ZN(n4545) );
  INV_X1 U5057 ( .A(n5114), .ZN(n4546) );
  INV_X1 U5058 ( .A(n4544), .ZN(n4543) );
  OAI21_X1 U5059 ( .B1(n4547), .B2(n4545), .A(n5113), .ZN(n4544) );
  INV_X1 U5060 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5511) );
  XNOR2_X1 U5061 ( .A(n5084), .B(SI_11_), .ZN(n5083) );
  NAND2_X1 U5062 ( .A1(n5050), .A2(n5049), .ZN(n5070) );
  NAND2_X1 U5063 ( .A1(n5048), .A2(n5033), .ZN(n5046) );
  NAND2_X1 U5064 ( .A1(n5045), .A2(n5014), .ZN(n5042) );
  NAND2_X1 U5065 ( .A1(n4990), .A2(n4989), .ZN(n5006) );
  AND2_X1 U5066 ( .A1(n4490), .A2(n8339), .ZN(n4489) );
  OR2_X1 U5067 ( .A1(n8412), .A2(n5405), .ZN(n4490) );
  AND2_X1 U5068 ( .A1(n4536), .A2(n4537), .ZN(n4533) );
  NOR2_X1 U5069 ( .A1(n7274), .A2(n4510), .ZN(n4509) );
  NAND2_X1 U5070 ( .A1(n4521), .A2(n4536), .ZN(n4532) );
  NAND2_X1 U5071 ( .A1(n6922), .A2(n4537), .ZN(n4535) );
  OR2_X1 U5072 ( .A1(n5290), .A2(n5289), .ZN(n5312) );
  NAND2_X1 U5073 ( .A1(n5067), .A2(n5068), .ZN(n4537) );
  OR2_X1 U5074 ( .A1(n7436), .A2(n5191), .ZN(n4507) );
  NOR2_X1 U5075 ( .A1(n4654), .A2(n4653), .ZN(n4652) );
  INV_X1 U5076 ( .A(n4658), .ZN(n4653) );
  OR3_X1 U5077 ( .A1(n7064), .A2(n7226), .A3(n7192), .ZN(n6175) );
  AND3_X1 U5078 ( .A1(n5279), .A2(n5278), .A3(n5277), .ZN(n8480) );
  OR2_X1 U5079 ( .A1(n7989), .A2(n7988), .ZN(n4386) );
  AND2_X1 U5080 ( .A1(n4386), .A2(n4385), .ZN(n8076) );
  NAND2_X1 U5081 ( .A1(n7340), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4385) );
  OR2_X1 U5082 ( .A1(n8076), .A2(n8075), .ZN(n4384) );
  AND2_X1 U5083 ( .A1(n8734), .A2(n4474), .ZN(n4473) );
  AND2_X1 U5084 ( .A1(n8541), .A2(n4471), .ZN(n8468) );
  AND2_X1 U5085 ( .A1(n4473), .A2(n4472), .ZN(n4471) );
  NAND2_X1 U5086 ( .A1(n8268), .A2(n8269), .ZN(n8490) );
  INV_X1 U5087 ( .A(n8488), .ZN(n4728) );
  AND2_X1 U5088 ( .A1(n8488), .A2(n8107), .ZN(n8510) );
  OAI21_X1 U5089 ( .B1(n8577), .B2(n8556), .A(n4328), .ZN(n8546) );
  NAND2_X1 U5090 ( .A1(n8587), .A2(n4751), .ZN(n4747) );
  OR2_X1 U5091 ( .A1(n8761), .A2(n8484), .ZN(n8485) );
  INV_X1 U5092 ( .A(n4749), .ZN(n4748) );
  OAI21_X1 U5093 ( .B1(n4751), .B2(n4750), .A(n8556), .ZN(n4749) );
  INV_X1 U5094 ( .A(n8485), .ZN(n4750) );
  INV_X1 U5095 ( .A(n4629), .ZN(n4625) );
  INV_X1 U5096 ( .A(n4633), .ZN(n4632) );
  OAI21_X1 U5097 ( .B1(n8105), .B2(n4634), .A(n8234), .ZN(n4633) );
  INV_X1 U5098 ( .A(n8104), .ZN(n4634) );
  NAND2_X1 U5099 ( .A1(n8642), .A2(n4635), .ZN(n4631) );
  OR2_X1 U5100 ( .A1(n4741), .A2(n4739), .ZN(n4738) );
  INV_X1 U5101 ( .A(n4744), .ZN(n4739) );
  INV_X1 U5102 ( .A(n4742), .ZN(n4741) );
  OAI21_X1 U5103 ( .B1(n8645), .B2(n4743), .A(n8482), .ZN(n4742) );
  NAND2_X1 U5104 ( .A1(n4780), .A2(n4744), .ZN(n4740) );
  NAND2_X1 U5105 ( .A1(n8229), .A2(n8227), .ZN(n8645) );
  NAND2_X1 U5106 ( .A1(n8637), .A2(n8645), .ZN(n8636) );
  NAND2_X1 U5107 ( .A1(n4622), .A2(n8129), .ZN(n4621) );
  INV_X1 U5108 ( .A(n4619), .ZN(n4617) );
  NOR2_X1 U5109 ( .A1(n4620), .A2(n4619), .ZN(n4613) );
  NAND2_X1 U5110 ( .A1(n8676), .A2(n4615), .ZN(n4614) );
  INV_X1 U5111 ( .A(n4621), .ZN(n4615) );
  NOR2_X1 U5112 ( .A1(n7387), .A2(n4352), .ZN(n4351) );
  INV_X1 U5113 ( .A(n8196), .ZN(n4352) );
  NAND2_X1 U5114 ( .A1(n8818), .A2(n4764), .ZN(n4763) );
  INV_X1 U5115 ( .A(n4638), .ZN(n4643) );
  AND4_X1 U5116 ( .A1(n5132), .A2(n5131), .A3(n5130), .A4(n5129), .ZN(n7302)
         );
  NAND2_X1 U5117 ( .A1(n8178), .A2(n8181), .ZN(n4646) );
  AND4_X1 U5118 ( .A1(n5108), .A2(n5107), .A3(n5106), .A4(n5105), .ZN(n7087)
         );
  NOR2_X1 U5119 ( .A1(n8173), .A2(n4333), .ZN(n4332) );
  INV_X1 U5120 ( .A(n8169), .ZN(n4333) );
  OR2_X1 U5121 ( .A1(n5023), .A2(n4816), .ZN(n5061) );
  NAND2_X1 U5122 ( .A1(n8696), .A2(n6778), .ZN(n4779) );
  NOR2_X1 U5123 ( .A1(n8290), .A2(n4624), .ZN(n6785) );
  INV_X1 U5124 ( .A(n8687), .ZN(n4624) );
  NAND2_X1 U5125 ( .A1(n6630), .A2(n6629), .ZN(n6775) );
  NAND2_X1 U5126 ( .A1(n6484), .A2(n6483), .ZN(n4720) );
  INV_X1 U5127 ( .A(n8146), .ZN(n8284) );
  OAI211_X1 U5128 ( .C1(n4944), .C2(n6208), .A(n4863), .B(n4862), .ZN(n6367)
         );
  NAND2_X1 U5129 ( .A1(n4974), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4863) );
  NAND2_X1 U5130 ( .A1(n5392), .A2(n5391), .ZN(n8752) );
  NAND2_X1 U5131 ( .A1(n7221), .A2(n8116), .ZN(n5392) );
  NAND2_X1 U5132 ( .A1(n5188), .A2(n5187), .ZN(n8802) );
  NAND2_X1 U5133 ( .A1(n4838), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U5134 ( .A1(n5845), .A2(n4592), .ZN(n4591) );
  NAND2_X1 U5135 ( .A1(n5849), .A2(n5850), .ZN(n4592) );
  AOI21_X1 U5136 ( .B1(n4584), .B2(n4588), .A(n4307), .ZN(n4582) );
  NAND2_X1 U5137 ( .A1(n7182), .A2(n4283), .ZN(n7284) );
  INV_X1 U5138 ( .A(n7287), .ZN(n4606) );
  NAND2_X1 U5139 ( .A1(n8919), .A2(n5957), .ZN(n8921) );
  OAI21_X1 U5140 ( .B1(n7529), .B2(n5850), .A(n5849), .ZN(n7533) );
  AND2_X1 U5141 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U5142 ( .A1(n7701), .A2(n7708), .ZN(n4567) );
  OR2_X1 U5143 ( .A1(n6302), .A2(n6303), .ZN(n4404) );
  OR2_X1 U5144 ( .A1(n7176), .A2(n9821), .ZN(n4400) );
  AND2_X1 U5145 ( .A1(n9128), .A2(n4423), .ZN(n9046) );
  NOR2_X1 U5146 ( .A1(n4424), .A2(n9049), .ZN(n4423) );
  INV_X1 U5147 ( .A(n4426), .ZN(n4424) );
  AOI21_X1 U5148 ( .B1(n9127), .B2(n9064), .A(n4699), .ZN(n9110) );
  NAND2_X1 U5149 ( .A1(n9079), .A2(n7767), .ZN(n9118) );
  AND4_X1 U5150 ( .A1(n6035), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n9135)
         );
  AOI21_X1 U5151 ( .B1(n7783), .B2(n9074), .A(n4461), .ZN(n4460) );
  INV_X1 U5152 ( .A(n9075), .ZN(n4461) );
  NAND2_X1 U5153 ( .A1(n9157), .A2(n7783), .ZN(n4459) );
  AND2_X1 U5154 ( .A1(n4459), .A2(n4456), .ZN(n9132) );
  NOR2_X1 U5155 ( .A1(n9159), .A2(n9158), .ZN(n9157) );
  NAND2_X1 U5156 ( .A1(n4683), .A2(n4689), .ZN(n4680) );
  AND2_X1 U5157 ( .A1(n9072), .A2(n7762), .ZN(n9172) );
  NAND2_X1 U5158 ( .A1(n9070), .A2(n4447), .ZN(n4446) );
  NAND2_X1 U5159 ( .A1(n7787), .A2(n7786), .ZN(n9201) );
  AND2_X1 U5160 ( .A1(n9069), .A2(n7789), .ZN(n9222) );
  AND2_X1 U5161 ( .A1(n9316), .A2(n9745), .ZN(n9052) );
  NAND2_X1 U5162 ( .A1(n7755), .A2(n7757), .ZN(n4437) );
  NAND2_X1 U5163 ( .A1(n4296), .A2(n7757), .ZN(n4436) );
  NAND2_X1 U5164 ( .A1(n4439), .A2(n7755), .ZN(n4438) );
  INV_X1 U5165 ( .A(n7642), .ZN(n4439) );
  NAND2_X1 U5166 ( .A1(n7463), .A2(n7479), .ZN(n4712) );
  NAND2_X1 U5167 ( .A1(n7412), .A2(n7642), .ZN(n7478) );
  AND2_X1 U5168 ( .A1(n7642), .A2(n7640), .ZN(n7811) );
  INV_X1 U5169 ( .A(n4675), .ZN(n4674) );
  AOI21_X1 U5170 ( .B1(n4675), .B2(n4673), .A(n4285), .ZN(n4672) );
  AND2_X1 U5171 ( .A1(n9418), .A2(n4676), .ZN(n4675) );
  NAND2_X1 U5172 ( .A1(n7628), .A2(n7205), .ZN(n4676) );
  NAND2_X1 U5173 ( .A1(n7019), .A2(n7205), .ZN(n4671) );
  NAND2_X1 U5174 ( .A1(n4677), .A2(n7806), .ZN(n7206) );
  INV_X1 U5175 ( .A(n7019), .ZN(n4677) );
  OR2_X1 U5176 ( .A1(n5719), .A2(n9819), .ZN(n5742) );
  INV_X1 U5177 ( .A(n4714), .ZN(n4713) );
  OAI21_X1 U5178 ( .B1(n7000), .B2(n7803), .A(n7001), .ZN(n4714) );
  NAND2_X1 U5179 ( .A1(n6572), .A2(n6132), .ZN(n7828) );
  INV_X1 U5180 ( .A(n7793), .ZN(n6935) );
  NAND3_X1 U5181 ( .A1(n6568), .A2(n6139), .A3(n6935), .ZN(n6934) );
  NAND2_X1 U5182 ( .A1(n7799), .A2(n6569), .ZN(n6568) );
  INV_X1 U5183 ( .A(n5571), .ZN(n4363) );
  XNOR2_X1 U5184 ( .A(n6131), .B(n7831), .ZN(n6574) );
  NAND2_X1 U5185 ( .A1(n6573), .A2(n6574), .ZN(n6572) );
  INV_X1 U5186 ( .A(n9043), .ZN(n9248) );
  AND2_X1 U5187 ( .A1(n9258), .A2(n9520), .ZN(n9259) );
  INV_X1 U5188 ( .A(n9131), .ZN(n9275) );
  NAND2_X1 U5189 ( .A1(n5896), .A2(n5895), .ZN(n9312) );
  NAND2_X1 U5190 ( .A1(n5793), .A2(n5792), .ZN(n9339) );
  OR2_X1 U5191 ( .A1(n7704), .A2(n7869), .ZN(n9335) );
  XNOR2_X1 U5192 ( .A(n4580), .B(n7582), .ZN(n8844) );
  OAI21_X1 U5193 ( .B1(n7585), .B2(n9881), .A(n7580), .ZN(n4580) );
  XNOR2_X1 U5194 ( .A(n7585), .B(SI_30_), .ZN(n8849) );
  XNOR2_X1 U5195 ( .A(n5408), .B(n5407), .ZN(n7221) );
  OAI21_X1 U5196 ( .B1(n5345), .B2(n4576), .A(n4574), .ZN(n5408) );
  NAND2_X1 U5197 ( .A1(n4569), .A2(n5286), .ZN(n5299) );
  NAND2_X1 U5198 ( .A1(n4542), .A2(n5086), .ZN(n5115) );
  NAND2_X1 U5199 ( .A1(n5071), .A2(n4547), .ZN(n4542) );
  OR2_X1 U5200 ( .A1(n5688), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5693) );
  CLKBUF_X1 U5201 ( .A(n5633), .Z(n5634) );
  XNOR2_X1 U5202 ( .A(n5572), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U5203 ( .A1(n7240), .A2(n8116), .ZN(n5416) );
  INV_X1 U5204 ( .A(n8601), .ZN(n8767) );
  AND4_X1 U5205 ( .A1(n5079), .A2(n5078), .A3(n5077), .A4(n5076), .ZN(n7118)
         );
  AND4_X1 U5206 ( .A1(n4826), .A2(n4825), .A3(n4824), .A4(n4823), .ZN(n7449)
         );
  AND4_X1 U5207 ( .A1(n5066), .A2(n5065), .A3(n5064), .A4(n5063), .ZN(n6980)
         );
  AND4_X1 U5208 ( .A1(n5257), .A2(n5256), .A3(n5255), .A4(n5254), .ZN(n8477)
         );
  INV_X1 U5209 ( .A(n6207), .ZN(n8093) );
  XNOR2_X1 U5210 ( .A(n4389), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U5211 ( .A1(n8445), .A2(n4390), .ZN(n4389) );
  OR2_X1 U5212 ( .A1(n8446), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4390) );
  NAND2_X1 U5213 ( .A1(n5369), .A2(n5368), .ZN(n8758) );
  NAND2_X1 U5214 ( .A1(n7189), .A2(n8116), .ZN(n5369) );
  NAND2_X1 U5215 ( .A1(n8577), .A2(n8244), .ZN(n8559) );
  NAND2_X1 U5216 ( .A1(n8587), .A2(n4790), .ZN(n8572) );
  NAND2_X1 U5217 ( .A1(n4851), .A2(n4850), .ZN(n7269) );
  NAND2_X1 U5218 ( .A1(n4841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4843) );
  AND4_X1 U5219 ( .A1(n6017), .A2(n6016), .A3(n6015), .A4(n6014), .ZN(n9121)
         );
  NAND2_X1 U5220 ( .A1(n6027), .A2(n6026), .ZN(n9269) );
  NAND2_X1 U5221 ( .A1(n7240), .A2(n5894), .ZN(n6027) );
  INV_X1 U5222 ( .A(n9182), .ZN(n9292) );
  AOI21_X1 U5223 ( .B1(n4599), .B2(n4598), .A(n4597), .ZN(n4596) );
  INV_X1 U5224 ( .A(n5715), .ZN(n4597) );
  INV_X1 U5225 ( .A(n4603), .ZN(n4598) );
  AND2_X1 U5226 ( .A1(n8950), .A2(n4593), .ZN(n6090) );
  NOR2_X1 U5227 ( .A1(n8862), .A2(n4594), .ZN(n4593) );
  INV_X1 U5228 ( .A(n6024), .ZN(n4594) );
  INV_X1 U5229 ( .A(n7831), .ZN(n7568) );
  NAND2_X1 U5230 ( .A1(n7182), .A2(n5755), .ZN(n7286) );
  AND4_X1 U5231 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .ZN(n8882)
         );
  NAND2_X1 U5232 ( .A1(n5909), .A2(n5908), .ZN(n9306) );
  NAND2_X1 U5233 ( .A1(n5812), .A2(n5811), .ZN(n9331) );
  NAND2_X1 U5234 ( .A1(n5547), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U5235 ( .A1(n6313), .A2(n4402), .ZN(n9474) );
  OR2_X1 U5236 ( .A1(n6321), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4402) );
  NAND2_X1 U5237 ( .A1(n4298), .A2(n4442), .ZN(n4441) );
  NAND2_X1 U5238 ( .A1(n4694), .A2(n4692), .ZN(n9066) );
  INV_X1 U5239 ( .A(n4693), .ZN(n4692) );
  NAND2_X1 U5240 ( .A1(n5778), .A2(n5777), .ZN(n7376) );
  INV_X1 U5241 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U5242 ( .A1(n4376), .A2(n4375), .ZN(n4374) );
  NOR2_X1 U5243 ( .A1(n7597), .A2(n7704), .ZN(n4375) );
  AOI21_X1 U5244 ( .B1(n4372), .B2(n4373), .A(n4284), .ZN(n4370) );
  INV_X1 U5245 ( .A(n4372), .ZN(n4371) );
  NAND2_X1 U5246 ( .A1(n4366), .A2(n7704), .ZN(n4365) );
  OAI21_X1 U5247 ( .B1(n7665), .B2(n7664), .A(n4368), .ZN(n4367) );
  NOR2_X1 U5248 ( .A1(n4369), .A2(n7704), .ZN(n4368) );
  NOR2_X1 U5249 ( .A1(n8303), .A2(n4760), .ZN(n4759) );
  INV_X1 U5250 ( .A(n4764), .ZN(n4760) );
  INV_X1 U5251 ( .A(n7379), .ZN(n4762) );
  NAND2_X1 U5252 ( .A1(n8972), .A2(n9527), .ZN(n7608) );
  OAI21_X1 U5253 ( .B1(n7694), .B2(n7576), .A(n7575), .ZN(n7579) );
  INV_X1 U5254 ( .A(n4564), .ZN(n4563) );
  OAI21_X1 U5255 ( .B1(n5428), .B2(n4565), .A(n7569), .ZN(n4564) );
  INV_X1 U5256 ( .A(n5430), .ZN(n4565) );
  OAI21_X1 U5257 ( .B1(n4525), .B2(n6923), .A(n4294), .ZN(n4323) );
  NAND2_X1 U5258 ( .A1(n4532), .A2(n4274), .ZN(n4525) );
  NAND2_X1 U5259 ( .A1(n4481), .A2(n4478), .ZN(n5356) );
  NAND2_X1 U5260 ( .A1(n4480), .A2(n4479), .ZN(n4478) );
  INV_X1 U5261 ( .A(n4484), .ZN(n4479) );
  XNOR2_X1 U5262 ( .A(n8758), .B(n5417), .ZN(n5381) );
  NOR2_X1 U5263 ( .A1(n8111), .A2(n4659), .ZN(n4658) );
  INV_X1 U5264 ( .A(n4662), .ZN(n4659) );
  NOR2_X1 U5265 ( .A1(n4330), .A2(n4286), .ZN(n4328) );
  NAND2_X1 U5266 ( .A1(n8548), .A2(n4331), .ZN(n4330) );
  OR2_X1 U5267 ( .A1(n8752), .A2(n8561), .ZN(n8254) );
  OR2_X1 U5268 ( .A1(n8774), .A2(n8593), .ZN(n8234) );
  OAI21_X1 U5269 ( .B1(n4738), .B2(n8607), .A(n4310), .ZN(n4735) );
  INV_X1 U5270 ( .A(n4740), .ZN(n4737) );
  NAND2_X1 U5271 ( .A1(n8103), .A2(n8229), .ZN(n8104) );
  INV_X1 U5272 ( .A(n8625), .ZN(n8103) );
  NOR2_X1 U5273 ( .A1(n8777), .A2(n4468), .ZN(n4467) );
  INV_X1 U5274 ( .A(n4469), .ZN(n4468) );
  OR2_X1 U5275 ( .A1(n5252), .A2(n5251), .ZN(n5274) );
  AND2_X1 U5276 ( .A1(n8788), .A2(n8477), .ZN(n8223) );
  NAND2_X1 U5277 ( .A1(n8129), .A2(n8210), .ZN(n4619) );
  NAND2_X1 U5278 ( .A1(n8206), .A2(n4353), .ZN(n4345) );
  INV_X1 U5279 ( .A(n4349), .ZN(n4348) );
  OAI21_X1 U5280 ( .B1(n4351), .B2(n4350), .A(n8205), .ZN(n4349) );
  OR2_X1 U5281 ( .A1(n5137), .A2(n5136), .ZN(n5139) );
  INV_X1 U5282 ( .A(n8189), .ZN(n4642) );
  NAND2_X1 U5283 ( .A1(n6799), .A2(n6798), .ZN(n6969) );
  INV_X1 U5284 ( .A(n4269), .ZN(n4774) );
  NAND2_X1 U5285 ( .A1(n6427), .A2(n6457), .ZN(n8136) );
  AND2_X1 U5286 ( .A1(n4793), .A2(n4794), .ZN(n4343) );
  OR3_X1 U5287 ( .A1(n5015), .A2(P2_IR_REG_7__SCAN_IN), .A3(
        P2_IR_REG_6__SCAN_IN), .ZN(n5097) );
  INV_X1 U5288 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4795) );
  AOI21_X1 U5289 ( .B1(n4587), .B2(n5957), .A(n4585), .ZN(n4584) );
  AND2_X1 U5290 ( .A1(n5960), .A2(n4586), .ZN(n4585) );
  INV_X1 U5291 ( .A(n5949), .ZN(n4587) );
  INV_X1 U5292 ( .A(n8889), .ZN(n4586) );
  OAI21_X1 U5293 ( .B1(n7706), .B2(n4377), .A(n7773), .ZN(n7702) );
  NAND2_X1 U5294 ( .A1(n7776), .A2(n9258), .ZN(n4377) );
  NOR2_X1 U5295 ( .A1(n9258), .A2(n4427), .ZN(n4426) );
  NAND2_X1 U5296 ( .A1(n9292), .A2(n9060), .ZN(n4689) );
  NAND2_X1 U5297 ( .A1(n4414), .A2(n9238), .ZN(n4413) );
  NOR2_X1 U5298 ( .A1(n9316), .A2(n9323), .ZN(n4414) );
  INV_X1 U5299 ( .A(n7205), .ZN(n4673) );
  OAI22_X1 U5300 ( .A1(n7016), .A2(n7015), .B1(n7075), .B2(n8969), .ZN(n9381)
         );
  NOR2_X1 U5301 ( .A1(n9422), .A2(n7376), .ZN(n7234) );
  AND2_X1 U5302 ( .A1(n7610), .A2(n7608), .ZN(n7801) );
  NAND2_X1 U5303 ( .A1(n5410), .A2(n5409), .ZN(n5429) );
  NAND2_X1 U5304 ( .A1(n4572), .A2(n4570), .ZN(n5410) );
  AOI21_X1 U5305 ( .B1(n4574), .B2(n4576), .A(n4571), .ZN(n4570) );
  NAND2_X1 U5306 ( .A1(n4577), .A2(n5361), .ZN(n4576) );
  INV_X1 U5307 ( .A(n5385), .ZN(n4577) );
  INV_X1 U5308 ( .A(n4575), .ZN(n4574) );
  OAI21_X1 U5309 ( .B1(n4578), .B2(n4576), .A(n5384), .ZN(n4575) );
  AND2_X1 U5310 ( .A1(n4715), .A2(n5517), .ZN(n4416) );
  NAND2_X1 U5311 ( .A1(n5285), .A2(n5284), .ZN(n4569) );
  NAND2_X1 U5312 ( .A1(n4299), .A2(n4255), .ZN(n4551) );
  AND2_X1 U5313 ( .A1(n5218), .A2(n5219), .ZN(n5224) );
  NAND2_X1 U5314 ( .A1(n4556), .A2(n4555), .ZN(n4554) );
  NAND2_X1 U5315 ( .A1(n4556), .A2(n4255), .ZN(n4552) );
  INV_X1 U5316 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4609) );
  XNOR2_X1 U5317 ( .A(n5157), .B(SI_14_), .ZN(n5156) );
  NAND2_X1 U5318 ( .A1(n4541), .A2(n4539), .ZN(n5147) );
  AOI21_X1 U5319 ( .B1(n4543), .B2(n4545), .A(n4540), .ZN(n4539) );
  NOR2_X1 U5320 ( .A1(n5087), .A2(n4548), .ZN(n4547) );
  INV_X1 U5321 ( .A(n5070), .ZN(n4548) );
  XNOR2_X1 U5322 ( .A(n5007), .B(SI_7_), .ZN(n5004) );
  XNOR2_X1 U5323 ( .A(n4988), .B(SI_6_), .ZN(n4985) );
  INV_X1 U5324 ( .A(n4968), .ZN(n4969) );
  XNOR2_X1 U5325 ( .A(n4971), .B(SI_5_), .ZN(n4968) );
  OAI21_X1 U5326 ( .B1(n4855), .B2(P1_ADDR_REG_19__SCAN_IN), .A(n4665), .ZN(
        n4857) );
  INV_X1 U5327 ( .A(n6347), .ZN(n4520) );
  INV_X1 U5328 ( .A(n6434), .ZN(n4514) );
  NAND2_X1 U5329 ( .A1(n4497), .A2(n4500), .ZN(n4493) );
  NAND2_X1 U5330 ( .A1(n5019), .A2(n5020), .ZN(n4500) );
  AND2_X1 U5331 ( .A1(n5261), .A2(n5260), .ZN(n8353) );
  INV_X1 U5332 ( .A(n7114), .ZN(n4531) );
  AOI21_X1 U5333 ( .B1(n4532), .B2(n4529), .A(n4528), .ZN(n4527) );
  NOR2_X1 U5334 ( .A1(n5112), .A2(n5111), .ZN(n4528) );
  NOR2_X1 U5335 ( .A1(n4533), .A2(n7114), .ZN(n4529) );
  XNOR2_X1 U5336 ( .A(n4897), .B(n4898), .ZN(n6428) );
  INV_X1 U5337 ( .A(n7275), .ZN(n4506) );
  OAI22_X1 U5338 ( .A1(n4507), .A2(n7446), .B1(n5215), .B2(n5214), .ZN(n4502)
         );
  INV_X1 U5339 ( .A(n4507), .ZN(n4503) );
  AOI21_X1 U5340 ( .B1(n8279), .B2(n8278), .A(n8277), .ZN(n8317) );
  INV_X1 U5341 ( .A(n6366), .ZN(n5486) );
  AND2_X1 U5342 ( .A1(n5424), .A2(n5423), .ZN(n8415) );
  AND4_X1 U5343 ( .A1(n5028), .A2(n5027), .A3(n5026), .A4(n5025), .ZN(n6965)
         );
  NAND2_X1 U5344 ( .A1(n8080), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4383) );
  NOR2_X1 U5345 ( .A1(n7976), .A2(n4388), .ZN(n7966) );
  NOR2_X1 U5346 ( .A1(n7985), .A2(n7313), .ZN(n4388) );
  NOR2_X1 U5347 ( .A1(n7966), .A2(n7965), .ZN(n7964) );
  NOR2_X1 U5348 ( .A1(n7964), .A2(n4387), .ZN(n7954) );
  AND2_X1 U5349 ( .A1(n7334), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4387) );
  NOR2_X1 U5350 ( .A1(n7954), .A2(n7953), .ZN(n7952) );
  NOR2_X1 U5351 ( .A1(n7940), .A2(n4393), .ZN(n7929) );
  AND2_X1 U5352 ( .A1(n7328), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4393) );
  NOR2_X1 U5353 ( .A1(n7929), .A2(n7930), .ZN(n7928) );
  NOR2_X1 U5354 ( .A1(n7928), .A2(n4392), .ZN(n8061) );
  AND2_X1 U5355 ( .A1(n7325), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4392) );
  NOR2_X1 U5356 ( .A1(n8061), .A2(n8062), .ZN(n8060) );
  NAND2_X1 U5357 ( .A1(n7899), .A2(n4382), .ZN(n8048) );
  OR2_X1 U5358 ( .A1(n7350), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4382) );
  NAND2_X1 U5359 ( .A1(n8048), .A2(n8049), .ZN(n8047) );
  XNOR2_X1 U5360 ( .A(n7321), .B(n8039), .ZN(n8035) );
  NAND2_X1 U5361 ( .A1(n8047), .A2(n4381), .ZN(n7321) );
  OR2_X1 U5362 ( .A1(n8053), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4381) );
  NOR2_X1 U5363 ( .A1(n8019), .A2(n4391), .ZN(n8023) );
  AND2_X1 U5364 ( .A1(n8020), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4391) );
  NAND2_X1 U5365 ( .A1(n8023), .A2(n8022), .ZN(n8445) );
  NAND2_X1 U5366 ( .A1(n4660), .A2(n4662), .ZN(n8491) );
  NAND2_X1 U5367 ( .A1(n8541), .A2(n8526), .ZN(n8521) );
  INV_X1 U5368 ( .A(n8538), .ZN(n8548) );
  NOR2_X1 U5369 ( .A1(n8247), .A2(n4329), .ZN(n4327) );
  NAND2_X1 U5370 ( .A1(n8254), .A2(n8527), .ZN(n8538) );
  AOI21_X1 U5371 ( .B1(n4748), .B2(n4750), .A(n4257), .ZN(n4746) );
  OR2_X1 U5372 ( .A1(n8761), .A2(n8592), .ZN(n8244) );
  NAND2_X1 U5373 ( .A1(n4628), .A2(n4626), .ZN(n8579) );
  NAND2_X1 U5374 ( .A1(n4629), .A2(n8237), .ZN(n4628) );
  AND2_X1 U5375 ( .A1(n4635), .A2(n8237), .ZN(n4627) );
  AND2_X1 U5376 ( .A1(n8244), .A2(n8245), .ZN(n8578) );
  NOR2_X1 U5377 ( .A1(n8642), .A2(n8104), .ZN(n8624) );
  NAND2_X1 U5378 ( .A1(n8670), .A2(n4467), .ZN(n8620) );
  NAND2_X1 U5379 ( .A1(n8670), .A2(n8658), .ZN(n8653) );
  NOR2_X1 U5380 ( .A1(n8224), .A2(n8223), .ZN(n8661) );
  AND2_X1 U5381 ( .A1(n4476), .A2(n4354), .ZN(n4475) );
  NAND2_X1 U5382 ( .A1(n9580), .A2(n4476), .ZN(n7298) );
  NOR2_X1 U5383 ( .A1(n6971), .A2(n4722), .ZN(n4721) );
  AND2_X1 U5384 ( .A1(n6978), .A2(n8181), .ZN(n9567) );
  NAND2_X1 U5385 ( .A1(n4817), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U5386 ( .A1(n6977), .A2(n8169), .ZN(n7043) );
  AOI21_X1 U5387 ( .B1(n8691), .B2(n8160), .A(n8291), .ZN(n6802) );
  INV_X1 U5388 ( .A(n4779), .ZN(n4777) );
  NAND2_X1 U5389 ( .A1(n6632), .A2(n8133), .ZN(n8688) );
  AOI21_X1 U5390 ( .B1(n8284), .B2(n4719), .A(n4288), .ZN(n4718) );
  INV_X1 U5391 ( .A(n6486), .ZN(n4719) );
  INV_X1 U5392 ( .A(n8286), .ZN(n6481) );
  AND2_X1 U5393 ( .A1(n6444), .A2(n8140), .ZN(n6445) );
  NAND2_X1 U5394 ( .A1(n6379), .A2(n9627), .ZN(n6368) );
  NAND2_X1 U5395 ( .A1(n7281), .A2(n8116), .ZN(n5433) );
  NAND2_X1 U5396 ( .A1(n5270), .A2(n5269), .ZN(n8783) );
  INV_X1 U5397 ( .A(n9690), .ZN(n9677) );
  AND2_X1 U5398 ( .A1(n5452), .A2(n4300), .ZN(n4810) );
  INV_X1 U5399 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4768) );
  INV_X1 U5400 ( .A(n5452), .ZN(n5455) );
  OR2_X1 U5401 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4828) );
  AND2_X1 U5402 ( .A1(n4343), .A2(n4753), .ZN(n4755) );
  INV_X1 U5403 ( .A(n4754), .ZN(n4757) );
  INV_X1 U5404 ( .A(n7069), .ZN(n4604) );
  OR2_X1 U5405 ( .A1(n6899), .A2(n6900), .ZN(n4603) );
  OAI22_X1 U5406 ( .A1(n6950), .A2(n6055), .B1(n9511), .B2(n5574), .ZN(n5620)
         );
  NAND2_X1 U5407 ( .A1(n6899), .A2(n6900), .ZN(n4602) );
  NAND2_X1 U5408 ( .A1(n6898), .A2(n4603), .ZN(n4601) );
  AOI21_X1 U5409 ( .B1(n6575), .B2(n5947), .A(n5563), .ZN(n6402) );
  NOR2_X1 U5410 ( .A1(n7779), .A2(n4358), .ZN(n4357) );
  NAND2_X1 U5411 ( .A1(n4359), .A2(n6827), .ZN(n4358) );
  INV_X1 U5412 ( .A(n7714), .ZN(n4359) );
  AND3_X1 U5413 ( .A1(n5569), .A2(n5570), .A3(n5568), .ZN(n4670) );
  NAND2_X1 U5414 ( .A1(n5665), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U5415 ( .A1(n6283), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4403) );
  OR2_X1 U5416 ( .A1(n6334), .A2(n6333), .ZN(n6336) );
  NOR2_X1 U5417 ( .A1(n9464), .A2(n4305), .ZN(n6290) );
  NAND2_X1 U5418 ( .A1(n6290), .A2(n6291), .ZN(n6313) );
  NOR2_X1 U5419 ( .A1(n9491), .A2(n4406), .ZN(n6317) );
  AND2_X1 U5420 ( .A1(n9498), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4406) );
  NOR2_X1 U5421 ( .A1(n6317), .A2(n6316), .ZN(n6588) );
  NOR2_X1 U5422 ( .A1(n6588), .A2(n4405), .ZN(n8978) );
  AND2_X1 U5423 ( .A1(n6589), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U5424 ( .A1(n8978), .A2(n8979), .ZN(n8977) );
  NOR2_X1 U5425 ( .A1(n6673), .A2(n4408), .ZN(n6677) );
  AND2_X1 U5426 ( .A1(n6674), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4408) );
  NOR2_X1 U5427 ( .A1(n6677), .A2(n6676), .ZN(n6913) );
  XNOR2_X1 U5428 ( .A(n7173), .B(n7172), .ZN(n6916) );
  NOR2_X1 U5429 ( .A1(n9012), .A2(n4319), .ZN(n9016) );
  NOR2_X1 U5430 ( .A1(n9016), .A2(n9015), .ZN(n9022) );
  INV_X1 U5431 ( .A(n4443), .ZN(n4442) );
  OAI21_X1 U5432 ( .B1(n9083), .B2(n9081), .A(n9412), .ZN(n4443) );
  NOR2_X1 U5433 ( .A1(n4701), .A2(n4696), .ZN(n4695) );
  INV_X1 U5434 ( .A(n9064), .ZN(n4696) );
  OAI21_X1 U5435 ( .B1(n4701), .B2(n4704), .A(n4697), .ZN(n4693) );
  AOI21_X1 U5436 ( .B1(n4700), .B2(n4698), .A(n4259), .ZN(n4697) );
  INV_X1 U5437 ( .A(n9118), .ZN(n4698) );
  INV_X1 U5438 ( .A(n4427), .ZN(n4425) );
  AND4_X1 U5439 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(n9105)
         );
  INV_X1 U5440 ( .A(n4462), .ZN(n9119) );
  AOI21_X1 U5441 ( .B1(n4456), .B2(n9076), .A(n9078), .ZN(n4455) );
  NOR2_X1 U5442 ( .A1(n9142), .A2(n9275), .ZN(n9128) );
  NOR2_X1 U5443 ( .A1(n9176), .A2(n9285), .ZN(n9162) );
  NAND2_X1 U5444 ( .A1(n9162), .A2(n9147), .ZN(n9142) );
  NAND2_X1 U5445 ( .A1(n9063), .A2(n9062), .ZN(n9141) );
  NAND2_X1 U5446 ( .A1(n9166), .A2(n9175), .ZN(n9062) );
  NAND2_X1 U5447 ( .A1(n4679), .A2(n4678), .ZN(n9063) );
  AOI21_X1 U5448 ( .B1(n4680), .B2(n4681), .A(n4260), .ZN(n4678) );
  NAND2_X1 U5449 ( .A1(n4685), .A2(n4689), .ZN(n4681) );
  AND2_X1 U5450 ( .A1(n5928), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U5451 ( .A1(n4449), .A2(n9071), .ZN(n4445) );
  AOI22_X1 U5452 ( .A1(n9231), .A2(n9056), .B1(n9055), .B2(n9238), .ZN(n9216)
         );
  INV_X1 U5453 ( .A(n4431), .ZN(n7507) );
  OR2_X1 U5454 ( .A1(n4437), .A2(n7470), .ZN(n4435) );
  INV_X1 U5455 ( .A(n4433), .ZN(n4432) );
  NOR2_X1 U5456 ( .A1(n7473), .A2(n9323), .ZN(n7503) );
  NOR2_X1 U5457 ( .A1(n7473), .A2(n4412), .ZN(n9232) );
  INV_X1 U5458 ( .A(n4414), .ZN(n4412) );
  AOI21_X1 U5459 ( .B1(n4710), .B2(n7409), .A(n4287), .ZN(n4709) );
  AND2_X1 U5460 ( .A1(n7234), .A2(n7463), .ZN(n7484) );
  NOR2_X1 U5461 ( .A1(n5795), .A2(n5794), .ZN(n5813) );
  OAI21_X1 U5462 ( .B1(n9406), .B2(n7209), .A(n7752), .ZN(n7230) );
  AND2_X1 U5463 ( .A1(n7632), .A2(n7629), .ZN(n7809) );
  NOR2_X1 U5464 ( .A1(n4420), .A2(n7204), .ZN(n4418) );
  OAI211_X1 U5465 ( .C1(n4454), .C2(n4452), .A(n4315), .B(n7749), .ZN(n7208)
         );
  NOR2_X1 U5466 ( .A1(n6863), .A2(n4420), .ZN(n9390) );
  NOR2_X1 U5467 ( .A1(n6863), .A2(n4419), .ZN(n9392) );
  INV_X1 U5468 ( .A(n4421), .ZN(n4419) );
  AND4_X1 U5469 ( .A1(n5725), .A2(n5724), .A3(n5723), .A4(n5722), .ZN(n7023)
         );
  NAND2_X1 U5470 ( .A1(n6829), .A2(n6142), .ZN(n6998) );
  AND2_X1 U5471 ( .A1(n7741), .A2(n7604), .ZN(n7797) );
  NAND2_X1 U5472 ( .A1(n6934), .A2(n6140), .ZN(n6698) );
  INV_X1 U5473 ( .A(n7795), .ZN(n6699) );
  AND2_X1 U5474 ( .A1(n6938), .A2(n6937), .ZN(n6940) );
  INV_X1 U5475 ( .A(n6941), .ZN(n6937) );
  NAND2_X1 U5476 ( .A1(n5939), .A2(n5938), .ZN(n9296) );
  AND2_X1 U5477 ( .A1(n6062), .A2(n6061), .ZN(n9520) );
  NOR2_X1 U5478 ( .A1(n4258), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4465) );
  XNOR2_X1 U5479 ( .A(n7694), .B(n7696), .ZN(n8330) );
  XNOR2_X1 U5480 ( .A(n7570), .B(n7569), .ZN(n7281) );
  NAND2_X1 U5481 ( .A1(n4562), .A2(n5430), .ZN(n7570) );
  NAND2_X1 U5482 ( .A1(n5429), .A2(n5428), .ZN(n4562) );
  XNOR2_X1 U5483 ( .A(n5429), .B(n5428), .ZN(n7240) );
  XNOR2_X1 U5484 ( .A(n5386), .B(n5385), .ZN(n7189) );
  NAND2_X1 U5485 ( .A1(n4573), .A2(n5361), .ZN(n5386) );
  XNOR2_X1 U5486 ( .A(n5363), .B(n5358), .ZN(n7062) );
  NAND2_X1 U5487 ( .A1(n4538), .A2(n4543), .ZN(n5145) );
  OR2_X1 U5488 ( .A1(n5071), .A2(n4545), .ZN(n4538) );
  NAND2_X1 U5489 ( .A1(n5071), .A2(n5070), .ZN(n5088) );
  XNOR2_X1 U5490 ( .A(n5035), .B(n5034), .ZN(n6226) );
  XNOR2_X1 U5491 ( .A(n4987), .B(n4985), .ZN(n6212) );
  NAND2_X1 U5492 ( .A1(n6620), .A2(n4978), .ZN(n6654) );
  NAND2_X1 U5493 ( .A1(n8411), .A2(n5406), .ZN(n8337) );
  NAND2_X1 U5494 ( .A1(n4488), .A2(n4487), .ZN(n5490) );
  AOI21_X1 U5495 ( .B1(n4489), .B2(n5405), .A(n5427), .ZN(n4487) );
  INV_X1 U5496 ( .A(n4494), .ZN(n6692) );
  AOI21_X1 U5497 ( .B1(n6620), .B2(n4499), .A(n4498), .ZN(n4494) );
  NAND2_X1 U5498 ( .A1(n4526), .A2(n4532), .ZN(n7113) );
  NAND2_X1 U5499 ( .A1(n6923), .A2(n4533), .ZN(n4526) );
  NOR2_X1 U5500 ( .A1(n4508), .A2(n7274), .ZN(n7445) );
  INV_X1 U5501 ( .A(n4511), .ZN(n4508) );
  NAND2_X1 U5502 ( .A1(n7444), .A2(n5192), .ZN(n7437) );
  NAND2_X1 U5503 ( .A1(n4518), .A2(n4520), .ZN(n4517) );
  INV_X1 U5504 ( .A(n6348), .ZN(n4518) );
  NAND2_X1 U5505 ( .A1(n4517), .A2(n4519), .ZN(n6433) );
  NAND2_X1 U5506 ( .A1(n4522), .A2(n4527), .ZN(n7079) );
  OR2_X1 U5507 ( .A1(n6923), .A2(n4530), .ZN(n4522) );
  NAND2_X1 U5508 ( .A1(n4532), .A2(n4531), .ZN(n4530) );
  AND3_X1 U5509 ( .A1(n5294), .A2(n5293), .A3(n5292), .ZN(n8610) );
  NAND2_X1 U5510 ( .A1(n4534), .A2(n4537), .ZN(n7035) );
  OR2_X1 U5511 ( .A1(n6923), .A2(n6922), .ZN(n4534) );
  INV_X1 U5512 ( .A(n6441), .ZN(n6427) );
  NAND2_X1 U5513 ( .A1(n5229), .A2(n5228), .ZN(n8792) );
  OR3_X1 U5514 ( .A1(n5491), .A2(n9677), .A3(n6178), .ZN(n8408) );
  INV_X1 U5515 ( .A(n8422), .ZN(n8406) );
  NAND2_X1 U5516 ( .A1(n5171), .A2(n5170), .ZN(n8807) );
  OR2_X1 U5517 ( .A1(n4654), .A2(n4301), .ZN(n4650) );
  CLKBUF_X1 U5518 ( .A(n5486), .Z(n8326) );
  INV_X1 U5519 ( .A(n4386), .ZN(n7987) );
  INV_X1 U5520 ( .A(n4384), .ZN(n8074) );
  NAND2_X1 U5521 ( .A1(n8118), .A2(n8117), .ZN(n8727) );
  NAND2_X1 U5522 ( .A1(n8541), .A2(n4473), .ZN(n8469) );
  NAND2_X1 U5523 ( .A1(n4729), .A2(n4727), .ZN(n8489) );
  AOI21_X1 U5524 ( .B1(n4730), .B2(n4732), .A(n4728), .ZN(n4727) );
  NAND2_X1 U5525 ( .A1(n8518), .A2(n8487), .ZN(n8511) );
  OAI21_X1 U5526 ( .B1(n8587), .B2(n4750), .A(n4748), .ZN(n8555) );
  NAND2_X1 U5527 ( .A1(n4747), .A2(n8485), .ZN(n8554) );
  AND2_X1 U5528 ( .A1(n5335), .A2(n5334), .ZN(n8601) );
  NAND2_X1 U5529 ( .A1(n4631), .A2(n4632), .ZN(n8589) );
  OAI21_X1 U5530 ( .B1(n8637), .B2(n4740), .A(n4738), .ZN(n8604) );
  NAND2_X1 U5531 ( .A1(n8636), .A2(n4780), .ZN(n8619) );
  NAND2_X1 U5532 ( .A1(n4616), .A2(n4621), .ZN(n8677) );
  NAND2_X1 U5533 ( .A1(n5201), .A2(n5200), .ZN(n8799) );
  NAND2_X1 U5534 ( .A1(n4347), .A2(n4353), .ZN(n7396) );
  NAND2_X1 U5535 ( .A1(n7301), .A2(n4351), .ZN(n4347) );
  INV_X1 U5536 ( .A(n8807), .ZN(n7386) );
  NAND2_X1 U5537 ( .A1(n7301), .A2(n8196), .ZN(n7388) );
  NAND2_X1 U5538 ( .A1(n8818), .A2(n4782), .ZN(n7297) );
  INV_X1 U5539 ( .A(n4763), .ZN(n7380) );
  NAND2_X1 U5540 ( .A1(n4641), .A2(n8189), .ZN(n7101) );
  NAND2_X1 U5541 ( .A1(n4644), .A2(n4643), .ZN(n4641) );
  NAND2_X1 U5542 ( .A1(n4644), .A2(n4636), .ZN(n7100) );
  OAI21_X1 U5543 ( .B1(n9565), .B2(n8178), .A(n8181), .ZN(n7093) );
  NAND2_X1 U5544 ( .A1(n4778), .A2(n4779), .ZN(n8710) );
  NAND2_X1 U5545 ( .A1(n4778), .A2(n4776), .ZN(n9647) );
  NAND2_X1 U5546 ( .A1(n6527), .A2(n8284), .ZN(n6529) );
  NAND2_X1 U5547 ( .A1(n4720), .A2(n6486), .ZN(n6527) );
  OR2_X1 U5548 ( .A1(n9589), .A2(n5480), .ZN(n8705) );
  INV_X1 U5549 ( .A(n8674), .ZN(n9577) );
  NAND2_X1 U5550 ( .A1(n4853), .A2(n4852), .ZN(n4854) );
  NAND2_X1 U5551 ( .A1(n4861), .A2(n4379), .ZN(n6207) );
  AOI22_X1 U5552 ( .A1(n4295), .A2(n8859), .B1(n4380), .B2(n8845), .ZN(n4379)
         );
  INV_X1 U5553 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4380) );
  CLKBUF_X1 U5554 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n8859) );
  AND4_X1 U5555 ( .A1(n5632), .A2(n5631), .A3(n5630), .A4(n5629), .ZN(n6949)
         );
  AND4_X1 U5556 ( .A1(n5748), .A2(n5747), .A3(n5746), .A4(n5745), .ZN(n9377)
         );
  NAND2_X1 U5557 ( .A1(n7529), .A2(n5821), .ZN(n7513) );
  INV_X1 U5558 ( .A(n4590), .ZN(n4589) );
  OAI21_X1 U5559 ( .B1(n4591), .B2(n4289), .A(n7515), .ZN(n4590) );
  NAND2_X1 U5560 ( .A1(n8871), .A2(n5972), .ZN(n8902) );
  AND4_X1 U5561 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .ZN(n7073)
         );
  NAND2_X1 U5562 ( .A1(n4601), .A2(n4602), .ZN(n7068) );
  AND4_X1 U5563 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .ZN(n9189)
         );
  INV_X1 U5564 ( .A(n7123), .ZN(n4605) );
  NAND2_X1 U5565 ( .A1(n5735), .A2(n7123), .ZN(n7181) );
  INV_X1 U5566 ( .A(n6608), .ZN(n5596) );
  AND4_X1 U5567 ( .A1(n5669), .A2(n5668), .A3(n5667), .A4(n5666), .ZN(n6906)
         );
  AND2_X1 U5568 ( .A1(n6816), .A2(n5658), .ZN(n5659) );
  NAND2_X1 U5569 ( .A1(n6008), .A2(n4309), .ZN(n8950) );
  INV_X1 U5570 ( .A(n8948), .ZN(n4595) );
  NAND2_X1 U5571 ( .A1(n6008), .A2(n6007), .ZN(n8949) );
  INV_X1 U5572 ( .A(n7541), .ZN(n8957) );
  AND2_X1 U5573 ( .A1(n6609), .A2(n9520), .ZN(n8914) );
  INV_X1 U5574 ( .A(n7073), .ZN(n8970) );
  INV_X1 U5575 ( .A(n4404), .ZN(n6301) );
  NAND2_X1 U5576 ( .A1(n9474), .A2(n9475), .ZN(n9473) );
  INV_X1 U5577 ( .A(n4400), .ZN(n7244) );
  OAI21_X1 U5578 ( .B1(n7176), .B2(n4398), .A(n4397), .ZN(n8995) );
  NAND2_X1 U5579 ( .A1(n4401), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4398) );
  NAND2_X1 U5580 ( .A1(n7245), .A2(n4401), .ZN(n4397) );
  INV_X1 U5581 ( .A(n7247), .ZN(n4401) );
  INV_X1 U5582 ( .A(n7245), .ZN(n4399) );
  XNOR2_X1 U5583 ( .A(n4395), .B(n4394), .ZN(n9032) );
  INV_X1 U5584 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4394) );
  OR2_X1 U5585 ( .A1(n9022), .A2(n4396), .ZN(n4395) );
  AND2_X1 U5586 ( .A1(n9025), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4396) );
  AND2_X1 U5587 ( .A1(n7584), .A2(n7583), .ZN(n9043) );
  NAND2_X1 U5588 ( .A1(n7587), .A2(n7586), .ZN(n9049) );
  NAND2_X1 U5589 ( .A1(n4702), .A2(n4700), .ZN(n9096) );
  NAND2_X1 U5590 ( .A1(n9110), .A2(n9118), .ZN(n4702) );
  NAND2_X1 U5591 ( .A1(n4459), .A2(n4460), .ZN(n9134) );
  AND2_X1 U5592 ( .A1(n6010), .A2(n6009), .ZN(n9131) );
  NOR2_X1 U5593 ( .A1(n9157), .A2(n9074), .ZN(n9149) );
  INV_X1 U5594 ( .A(n9279), .ZN(n9147) );
  AND2_X1 U5595 ( .A1(n5962), .A2(n5961), .ZN(n9182) );
  NAND2_X1 U5596 ( .A1(n4682), .A2(n4685), .ZN(n9170) );
  NAND2_X1 U5597 ( .A1(n9198), .A2(n4270), .ZN(n4682) );
  AND2_X1 U5598 ( .A1(n4686), .A2(n4690), .ZN(n9185) );
  NAND2_X1 U5599 ( .A1(n9198), .A2(n9201), .ZN(n4686) );
  NAND2_X1 U5600 ( .A1(n5927), .A2(n5926), .ZN(n9303) );
  NAND2_X1 U5601 ( .A1(n9070), .A2(n9069), .ZN(n9200) );
  INV_X1 U5602 ( .A(n4446), .ZN(n9199) );
  INV_X1 U5603 ( .A(n9312), .ZN(n9238) );
  NAND2_X1 U5604 ( .A1(n4430), .A2(n4436), .ZN(n7506) );
  OR2_X1 U5605 ( .A1(n7412), .A2(n4437), .ZN(n4430) );
  NAND2_X1 U5606 ( .A1(n5832), .A2(n5831), .ZN(n9328) );
  NAND2_X1 U5607 ( .A1(n7478), .A2(n7755), .ZN(n7471) );
  INV_X1 U5608 ( .A(n9331), .ZN(n7490) );
  AND2_X1 U5609 ( .A1(n4711), .A2(n4712), .ZN(n7480) );
  OR2_X1 U5610 ( .A1(n7410), .A2(n7409), .ZN(n4711) );
  INV_X1 U5611 ( .A(n9339), .ZN(n7463) );
  NAND2_X1 U5612 ( .A1(n5761), .A2(n5760), .ZN(n9416) );
  NAND2_X1 U5613 ( .A1(n4671), .A2(n4675), .ZN(n9417) );
  NAND2_X1 U5614 ( .A1(n7206), .A2(n7205), .ZN(n9419) );
  AND2_X1 U5615 ( .A1(n6568), .A2(n6139), .ZN(n6936) );
  INV_X1 U5616 ( .A(n9033), .ZN(n9211) );
  AOI22_X1 U5617 ( .A1(n6128), .A2(n6283), .B1(n5674), .B2(n4362), .ZN(n4409)
         );
  INV_X1 U5618 ( .A(n6208), .ZN(n4362) );
  NOR2_X1 U5619 ( .A1(n9260), .A2(n9259), .ZN(n9261) );
  INV_X1 U5620 ( .A(n9255), .ZN(n9263) );
  NAND2_X1 U5621 ( .A1(n5538), .A2(n4463), .ZN(n9362) );
  AND2_X1 U5622 ( .A1(n4465), .A2(n4464), .ZN(n4463) );
  INV_X1 U5623 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4464) );
  INV_X1 U5624 ( .A(n5758), .ZN(n5775) );
  AND2_X1 U5625 ( .A1(n5633), .A2(n5510), .ZN(n5756) );
  XNOR2_X1 U5626 ( .A(n5689), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9484) );
  XNOR2_X1 U5627 ( .A(n5671), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6321) );
  AND2_X1 U5628 ( .A1(n5648), .A2(n5647), .ZN(n9458) );
  NAND2_X1 U5629 ( .A1(n4705), .A2(n5587), .ZN(n5616) );
  INV_X1 U5630 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8461) );
  INV_X1 U5631 ( .A(n4355), .ZN(n7878) );
  NOR2_X1 U5632 ( .A1(n4865), .A2(n5493), .ZN(n4886) );
  NAND2_X1 U5633 ( .A1(n8106), .A2(n8527), .ZN(n4254) );
  INV_X1 U5634 ( .A(n8556), .ZN(n8558) );
  XNOR2_X1 U5635 ( .A(n8758), .B(n8424), .ZN(n8556) );
  OR2_X1 U5636 ( .A1(n5223), .A2(n5222), .ZN(n4255) );
  INV_X1 U5637 ( .A(n4701), .ZN(n4700) );
  NAND2_X1 U5638 ( .A1(n9103), .A2(n4268), .ZN(n4701) );
  AND2_X1 U5639 ( .A1(n8164), .A2(n8165), .ZN(n8159) );
  OR2_X1 U5640 ( .A1(n8807), .A2(n7449), .ZN(n8206) );
  AND4_X1 U5641 ( .A1(n5095), .A2(n5166), .A3(n4965), .A4(n4966), .ZN(n4256)
         );
  INV_X1 U5642 ( .A(n7656), .ZN(n4434) );
  OR2_X1 U5643 ( .A1(n9264), .A2(n9120), .ZN(n9081) );
  INV_X1 U5644 ( .A(n8483), .ZN(n8607) );
  AND2_X1 U5645 ( .A1(n5288), .A2(n5287), .ZN(n8623) );
  INV_X1 U5646 ( .A(n8623), .ZN(n8777) );
  AND4_X1 U5647 ( .A1(n5645), .A2(n5644), .A3(n5643), .A4(n5642), .ZN(n6831)
         );
  AND2_X1 U5648 ( .A1(n8462), .A2(n8424), .ZN(n4257) );
  OR2_X1 U5649 ( .A1(n4278), .A2(n4706), .ZN(n4258) );
  NAND2_X1 U5650 ( .A1(n5081), .A2(n5082), .ZN(n4536) );
  AND2_X1 U5651 ( .A1(n9264), .A2(n4703), .ZN(n4259) );
  AND2_X1 U5652 ( .A1(n9285), .A2(n4688), .ZN(n4260) );
  AND2_X1 U5653 ( .A1(n4467), .A2(n4466), .ZN(n4261) );
  NOR2_X1 U5654 ( .A1(n6801), .A2(n4335), .ZN(n4262) );
  AND2_X1 U5655 ( .A1(n7803), .A2(n7611), .ZN(n4454) );
  NAND2_X1 U5656 ( .A1(n9580), .A2(n4477), .ZN(n4263) );
  NOR2_X1 U5657 ( .A1(n4757), .A2(n4756), .ZN(n4264) );
  INV_X1 U5658 ( .A(n6055), .ZN(n5789) );
  INV_X1 U5659 ( .A(n5673), .ZN(n5736) );
  AND2_X1 U5660 ( .A1(n6455), .A2(n4880), .ZN(n4266) );
  OR2_X1 U5661 ( .A1(n9279), .A2(n9161), .ZN(n7783) );
  NOR2_X1 U5662 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4860) );
  NAND2_X1 U5663 ( .A1(n4936), .A2(n4935), .ZN(n4937) );
  AND4_X1 U5664 ( .A1(n5053), .A2(n5148), .A3(n5121), .A4(n5094), .ZN(n4267)
         );
  OR2_X1 U5665 ( .A1(n9269), .A2(n9065), .ZN(n4268) );
  OR2_X1 U5666 ( .A1(n8696), .A2(n6778), .ZN(n4269) );
  OR2_X1 U5667 ( .A1(n8812), .A2(n8428), .ZN(n7379) );
  INV_X1 U5668 ( .A(n8247), .ZN(n4331) );
  AND2_X1 U5669 ( .A1(n4691), .A2(n9201), .ZN(n4270) );
  INV_X1 U5670 ( .A(n4893), .ZN(n4797) );
  OR2_X1 U5671 ( .A1(n8799), .A2(n7425), .ZN(n8129) );
  NOR2_X1 U5672 ( .A1(n4999), .A2(n4998), .ZN(n4498) );
  AND2_X1 U5673 ( .A1(n7690), .A2(n7689), .ZN(n4271) );
  AND2_X1 U5674 ( .A1(n4956), .A2(n4957), .ZN(n4272) );
  INV_X1 U5675 ( .A(n8125), .ZN(n4661) );
  XNOR2_X1 U5676 ( .A(n8746), .B(n8415), .ZN(n8530) );
  OR2_X1 U5677 ( .A1(n5541), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4273) );
  NAND2_X1 U5678 ( .A1(n8767), .A2(n8611), .ZN(n8237) );
  INV_X1 U5679 ( .A(n8181), .ZN(n4649) );
  NAND2_X1 U5680 ( .A1(n4486), .A2(n5321), .ZN(n8344) );
  NAND4_X1 U5681 ( .A1(n4876), .A2(n4875), .A3(n4874), .A4(n4873), .ZN(n6379)
         );
  NAND2_X1 U5682 ( .A1(n7698), .A2(n7697), .ZN(n9258) );
  NOR2_X1 U5683 ( .A1(n4340), .A2(n4339), .ZN(n4849) );
  AND2_X1 U5684 ( .A1(n4531), .A2(n7078), .ZN(n4274) );
  AND2_X1 U5685 ( .A1(n4384), .A2(n4383), .ZN(n4275) );
  AND2_X1 U5686 ( .A1(n4404), .A2(n4403), .ZN(n4276) );
  OAI21_X1 U5687 ( .B1(n8413), .B2(n5405), .A(n4489), .ZN(n8338) );
  INV_X1 U5688 ( .A(n7446), .ZN(n4510) );
  AND2_X1 U5689 ( .A1(n4253), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n4277) );
  OR2_X1 U5690 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n4278) );
  AND2_X1 U5691 ( .A1(n9296), .A2(n9059), .ZN(n4279) );
  NAND2_X1 U5692 ( .A1(n5878), .A2(n5877), .ZN(n9316) );
  NOR2_X1 U5693 ( .A1(n7180), .A2(n4605), .ZN(n4280) );
  INV_X1 U5694 ( .A(n6196), .ZN(n4930) );
  AND2_X1 U5695 ( .A1(n5250), .A2(n5249), .ZN(n8658) );
  INV_X1 U5696 ( .A(n8658), .ZN(n8788) );
  AND2_X1 U5697 ( .A1(n4446), .A2(n7786), .ZN(n4281) );
  NAND2_X1 U5698 ( .A1(n5416), .A2(n5415), .ZN(n8746) );
  AND2_X1 U5699 ( .A1(n4336), .A2(n8294), .ZN(n4282) );
  AND2_X1 U5700 ( .A1(n4606), .A2(n5755), .ZN(n4283) );
  OR2_X1 U5701 ( .A1(n8783), .A2(n8480), .ZN(n8229) );
  INV_X1 U5702 ( .A(n8303), .ZN(n4766) );
  AND2_X1 U5703 ( .A1(n8206), .A2(n8205), .ZN(n8303) );
  INV_X1 U5704 ( .A(n4353), .ZN(n4350) );
  NAND2_X1 U5705 ( .A1(n4354), .A2(n8428), .ZN(n4353) );
  AND2_X1 U5706 ( .A1(n7759), .A2(n7708), .ZN(n4284) );
  AND2_X1 U5707 ( .A1(n9416), .A2(n8967), .ZN(n4285) );
  AND2_X1 U5708 ( .A1(n8558), .A2(n4329), .ZN(n4286) );
  NOR2_X1 U5709 ( .A1(n7490), .A2(n7462), .ZN(n4287) );
  AND2_X1 U5710 ( .A1(n6488), .A2(n6487), .ZN(n4288) );
  OR2_X1 U5711 ( .A1(n5849), .A2(n5821), .ZN(n4289) );
  AND2_X1 U5712 ( .A1(n4625), .A2(n4631), .ZN(n4290) );
  NAND2_X1 U5713 ( .A1(n6042), .A2(n6041), .ZN(n9264) );
  AND2_X1 U5714 ( .A1(n8436), .A2(n9649), .ZN(n4291) );
  AOI21_X1 U5715 ( .B1(n4558), .B2(n5160), .A(n4557), .ZN(n4556) );
  NOR2_X1 U5716 ( .A1(n8807), .A2(n8427), .ZN(n4292) );
  INV_X1 U5717 ( .A(n4648), .ZN(n4647) );
  OR2_X1 U5718 ( .A1(n7092), .A2(n4649), .ZN(n4648) );
  AND2_X1 U5719 ( .A1(n5047), .A2(n5048), .ZN(n4293) );
  NAND2_X1 U5720 ( .A1(n5134), .A2(n5135), .ZN(n4294) );
  AND2_X1 U5721 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4295) );
  INV_X1 U5722 ( .A(n4780), .ZN(n4743) );
  OAI21_X1 U5723 ( .B1(n4270), .B2(n4684), .A(n9061), .ZN(n4683) );
  INV_X1 U5724 ( .A(n4685), .ZN(n4684) );
  NAND2_X1 U5725 ( .A1(n4297), .A2(n4691), .ZN(n4685) );
  NAND2_X1 U5726 ( .A1(n7736), .A2(n4438), .ZN(n4296) );
  INV_X1 U5727 ( .A(n4498), .ZN(n4497) );
  OR2_X1 U5728 ( .A1(n4687), .A2(n4279), .ZN(n4297) );
  NAND2_X1 U5729 ( .A1(n9083), .A2(n9081), .ZN(n4298) );
  NAND2_X1 U5730 ( .A1(n4554), .A2(n5224), .ZN(n4299) );
  AND2_X1 U5731 ( .A1(n4770), .A2(n4768), .ZN(n4300) );
  AND2_X1 U5732 ( .A1(n4656), .A2(n4655), .ZN(n4301) );
  AND2_X1 U5733 ( .A1(n4449), .A2(n4447), .ZN(n4302) );
  AND2_X1 U5734 ( .A1(n4702), .A2(n4268), .ZN(n4303) );
  NAND2_X1 U5735 ( .A1(n8109), .A2(n8108), .ZN(n8499) );
  AND2_X1 U5736 ( .A1(n4416), .A2(n4415), .ZN(n4304) );
  INV_X1 U5737 ( .A(n4600), .ZN(n4599) );
  NAND2_X1 U5738 ( .A1(n4604), .A2(n4602), .ZN(n4600) );
  INV_X1 U5739 ( .A(n4457), .ZN(n4456) );
  NAND2_X1 U5740 ( .A1(n4460), .A2(n4458), .ZN(n4457) );
  NAND2_X1 U5741 ( .A1(n5433), .A2(n5432), .ZN(n8741) );
  NAND2_X1 U5742 ( .A1(n7272), .A2(n7275), .ZN(n4511) );
  NAND2_X1 U5743 ( .A1(n9565), .A2(n4647), .ZN(n4644) );
  INV_X1 U5744 ( .A(n9175), .ZN(n4688) );
  NAND2_X1 U5745 ( .A1(n8113), .A2(n8112), .ZN(n8470) );
  INV_X1 U5746 ( .A(n8470), .ZN(n4472) );
  AND2_X1 U5747 ( .A1(n5379), .A2(n5378), .ZN(n8424) );
  AND2_X1 U5748 ( .A1(n9470), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4305) );
  NAND2_X1 U5749 ( .A1(n4504), .A2(n4501), .ZN(n7495) );
  AND2_X1 U5750 ( .A1(n4763), .A2(n7379), .ZN(n4306) );
  XOR2_X1 U5751 ( .A(n5970), .B(n6870), .Z(n4307) );
  INV_X1 U5752 ( .A(n9171), .ZN(n4369) );
  INV_X1 U5753 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4965) );
  AND3_X1 U5754 ( .A1(n4754), .A2(n4755), .A3(n4797), .ZN(n5196) );
  INV_X1 U5755 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4966) );
  NAND2_X1 U5756 ( .A1(n7196), .A2(n7197), .ZN(n7195) );
  NAND2_X1 U5757 ( .A1(n4509), .A2(n4511), .ZN(n7444) );
  OAI21_X1 U5758 ( .B1(n7092), .B2(n4646), .A(n8187), .ZN(n4645) );
  INV_X1 U5759 ( .A(n4645), .ZN(n4636) );
  AND4_X1 U5760 ( .A1(n6050), .A2(n6049), .A3(n6048), .A4(n6047), .ZN(n9120)
         );
  INV_X1 U5761 ( .A(n9120), .ZN(n4703) );
  NOR3_X1 U5762 ( .A1(n7473), .A2(n9306), .A3(n4413), .ZN(n4410) );
  NAND2_X1 U5763 ( .A1(n8670), .A2(n4469), .ZN(n4470) );
  AND2_X1 U5764 ( .A1(n4400), .A2(n4399), .ZN(n4308) );
  INV_X1 U5765 ( .A(n4411), .ZN(n9233) );
  NOR2_X1 U5766 ( .A1(n7473), .A2(n4413), .ZN(n4411) );
  AND2_X1 U5767 ( .A1(n4595), .A2(n6007), .ZN(n4309) );
  OR2_X1 U5768 ( .A1(n8774), .A2(n8629), .ZN(n4310) );
  AND2_X1 U5769 ( .A1(n5286), .A2(n5268), .ZN(n5284) );
  INV_X1 U5770 ( .A(n4704), .ZN(n4699) );
  NAND2_X1 U5771 ( .A1(n9275), .A2(n9150), .ZN(n4704) );
  AND3_X1 U5772 ( .A1(n4793), .A2(n4794), .A3(n4796), .ZN(n4311) );
  AND2_X1 U5773 ( .A1(n5300), .A2(n5286), .ZN(n4312) );
  AND2_X1 U5774 ( .A1(n4618), .A2(n4614), .ZN(n4313) );
  INV_X1 U5775 ( .A(n4690), .ZN(n4687) );
  NAND2_X1 U5776 ( .A1(n9303), .A2(n9225), .ZN(n4690) );
  AND2_X1 U5777 ( .A1(n4267), .A2(n4256), .ZN(n4754) );
  AND2_X1 U5778 ( .A1(n6165), .A2(n9209), .ZN(n9386) );
  INV_X1 U5779 ( .A(n9386), .ZN(n7027) );
  NAND2_X1 U5780 ( .A1(n5152), .A2(n5151), .ZN(n8812) );
  INV_X1 U5781 ( .A(n8812), .ZN(n4354) );
  NAND2_X1 U5782 ( .A1(n6817), .A2(n6816), .ZN(n4314) );
  INV_X1 U5783 ( .A(n8160), .ZN(n4335) );
  OAI21_X1 U5784 ( .B1(n6998), .B2(n6997), .A(n4713), .ZN(n7016) );
  NAND2_X1 U5785 ( .A1(n5310), .A2(n5309), .ZN(n8774) );
  INV_X1 U5786 ( .A(n8774), .ZN(n4466) );
  AND2_X1 U5787 ( .A1(n7633), .A2(n7750), .ZN(n7628) );
  NAND2_X1 U5788 ( .A1(n4334), .A2(n4282), .ZN(n6977) );
  OR2_X1 U5789 ( .A1(n6858), .A2(n4452), .ZN(n4315) );
  AND2_X1 U5790 ( .A1(n4601), .A2(n4599), .ZN(n4316) );
  AND2_X1 U5791 ( .A1(n9580), .A2(n9684), .ZN(n4317) );
  AND2_X1 U5792 ( .A1(n7572), .A2(n7571), .ZN(n4318) );
  INV_X1 U5793 ( .A(n4422), .ZN(n7003) );
  NOR2_X1 U5794 ( .A1(n6863), .A2(n6999), .ZN(n4422) );
  XNOR2_X1 U5795 ( .A(n4608), .B(P1_IR_REG_22__SCAN_IN), .ZN(n7875) );
  NAND2_X1 U5796 ( .A1(n4854), .A2(n4808), .ZN(n5492) );
  INV_X1 U5797 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4715) );
  AND2_X1 U5798 ( .A1(n9013), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4319) );
  AND2_X1 U5799 ( .A1(n4517), .A2(n4516), .ZN(n4320) );
  OR2_X1 U5800 ( .A1(n7716), .A2(n7715), .ZN(n4321) );
  INV_X2 U5801 ( .A(n8851), .ZN(n8856) );
  NAND2_X1 U5802 ( .A1(n4910), .A2(n4909), .ZN(n4925) );
  NAND2_X1 U5803 ( .A1(n4364), .A2(n7679), .ZN(n7688) );
  MUX2_X1 U5804 ( .A(n7615), .B(n7614), .S(n7704), .Z(n7622) );
  NAND2_X2 U5805 ( .A1(n8537), .A2(n4324), .ZN(n8519) );
  NAND2_X2 U5806 ( .A1(n8539), .A2(n8538), .ZN(n8537) );
  OAI22_X2 U5807 ( .A1(n8669), .A2(n8476), .B1(n8675), .B2(n8475), .ZN(n8652)
         );
  AND4_X2 U5808 ( .A1(n4716), .A2(n5633), .A3(n5516), .A4(n4715), .ZN(n5538)
         );
  NAND2_X1 U5809 ( .A1(n4726), .A2(n4730), .ZN(n8509) );
  AND2_X4 U5810 ( .A1(n5524), .A2(n5523), .ZN(n5665) );
  INV_X1 U5811 ( .A(n7598), .ZN(n4376) );
  NOR2_X2 U5812 ( .A1(n7423), .A2(n8304), .ZN(n7422) );
  OAI21_X2 U5813 ( .B1(n7650), .B2(n4371), .A(n4370), .ZN(n7659) );
  NAND2_X1 U5814 ( .A1(n7793), .A2(n7828), .ZN(n4429) );
  NAND2_X2 U5815 ( .A1(n5037), .A2(n5036), .ZN(n7056) );
  OAI211_X1 U5816 ( .C1(n7599), .C2(n7708), .A(n7603), .B(n4374), .ZN(n7607)
         );
  AND2_X1 U5817 ( .A1(n7672), .A2(n7717), .ZN(n4366) );
  NAND2_X1 U5818 ( .A1(n4566), .A2(n7713), .ZN(n4361) );
  NAND2_X1 U5819 ( .A1(n6487), .A2(n8439), .ZN(n8152) );
  NAND2_X1 U5820 ( .A1(n8691), .A2(n4262), .ZN(n4334) );
  NAND4_X1 U5821 ( .A1(n4343), .A2(n4267), .A3(n4256), .A4(n4337), .ZN(n4340)
         );
  NAND3_X1 U5822 ( .A1(n4803), .A2(n4797), .A3(n4769), .ZN(n4339) );
  NAND3_X1 U5823 ( .A1(n4342), .A2(n4755), .A3(n4754), .ZN(n5450) );
  NOR2_X2 U5824 ( .A1(n4363), .A2(n6196), .ZN(n5674) );
  NAND4_X1 U5825 ( .A1(n4367), .A2(n4365), .A3(n7673), .A4(n9172), .ZN(n4364)
         );
  NAND2_X1 U5826 ( .A1(n7598), .A2(n7742), .ZN(n7599) );
  NAND2_X1 U5827 ( .A1(n6134), .A2(n7836), .ZN(n7598) );
  OAI21_X2 U5828 ( .B1(n4271), .B2(n4378), .A(n7693), .ZN(n7706) );
  XNOR2_X1 U5829 ( .A(n7243), .B(n7249), .ZN(n7176) );
  NOR2_X4 U5830 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4705) );
  NAND3_X2 U5831 ( .A1(n5587), .A2(n4705), .A3(n5506), .ZN(n4428) );
  NOR2_X4 U5832 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5587) );
  NAND2_X1 U5833 ( .A1(n5573), .A2(n4409), .ZN(n7831) );
  INV_X2 U5834 ( .A(n5571), .ZN(n6128) );
  INV_X1 U5835 ( .A(n4410), .ZN(n9217) );
  NAND4_X1 U5836 ( .A1(n4716), .A2(n5634), .A3(n4304), .A4(n5516), .ZN(n6101)
         );
  NAND4_X1 U5837 ( .A1(n4716), .A2(n5633), .A3(n5516), .A4(n4416), .ZN(n5541)
         );
  INV_X1 U5838 ( .A(n6863), .ZN(n4417) );
  NAND2_X1 U5839 ( .A1(n4418), .A2(n4417), .ZN(n9421) );
  AND2_X1 U5840 ( .A1(n9128), .A2(n4425), .ZN(n9097) );
  NAND2_X1 U5841 ( .A1(n9128), .A2(n4426), .ZN(n9087) );
  NAND2_X1 U5842 ( .A1(n9128), .A2(n9116), .ZN(n9111) );
  NAND2_X1 U5843 ( .A1(n4428), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5646) );
  NOR2_X4 U5844 ( .A1(n4428), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5633) );
  AND2_X1 U5845 ( .A1(n7838), .A2(n7834), .ZN(n7793) );
  OAI21_X1 U5846 ( .B1(n7412), .B2(n4435), .A(n4432), .ZN(n4431) );
  OAI211_X1 U5847 ( .C1(n9102), .C2(n4441), .A(n9086), .B(n4440), .ZN(n9255)
         );
  NAND3_X1 U5848 ( .A1(n9102), .A2(n9083), .A3(n4442), .ZN(n4440) );
  NAND2_X1 U5849 ( .A1(n9070), .A2(n4302), .ZN(n4444) );
  NAND2_X1 U5850 ( .A1(n4444), .A2(n4445), .ZN(n9186) );
  NAND3_X1 U5851 ( .A1(n4451), .A2(n4450), .A3(n7633), .ZN(n9406) );
  NAND3_X1 U5852 ( .A1(n7749), .A2(n4452), .A3(n7750), .ZN(n4450) );
  NAND4_X1 U5853 ( .A1(n7749), .A2(n4454), .A3(n6858), .A4(n7750), .ZN(n4451)
         );
  NAND2_X1 U5854 ( .A1(n9374), .A2(n7621), .ZN(n7022) );
  NAND2_X1 U5855 ( .A1(n6858), .A2(n4454), .ZN(n9374) );
  NAND2_X1 U5856 ( .A1(n4453), .A2(n7621), .ZN(n4452) );
  INV_X1 U5857 ( .A(n7624), .ZN(n4453) );
  OAI21_X1 U5858 ( .B1(n9157), .B2(n4457), .A(n4455), .ZN(n4462) );
  AND2_X1 U5859 ( .A1(n5538), .A2(n4465), .ZN(n5560) );
  NAND2_X1 U5860 ( .A1(n5452), .A2(n4804), .ZN(n5457) );
  AND2_X2 U5861 ( .A1(n8670), .A2(n4261), .ZN(n8612) );
  INV_X1 U5862 ( .A(n4470), .ZN(n8638) );
  AND2_X1 U5863 ( .A1(n8541), .A2(n4474), .ZN(n8512) );
  NAND2_X1 U5864 ( .A1(n8401), .A2(n8402), .ZN(n4486) );
  NAND2_X1 U5865 ( .A1(n8401), .A2(n4482), .ZN(n4481) );
  NAND2_X1 U5866 ( .A1(n8413), .A2(n4489), .ZN(n4488) );
  NAND2_X1 U5867 ( .A1(n8413), .A2(n8412), .ZN(n8411) );
  OAI21_X2 U5868 ( .B1(n6620), .B2(n4493), .A(n4491), .ZN(n6746) );
  NAND2_X1 U5869 ( .A1(n4492), .A2(n4500), .ZN(n4491) );
  NAND2_X1 U5870 ( .A1(n6691), .A2(n4495), .ZN(n4492) );
  OAI21_X2 U5871 ( .B1(n6348), .B2(n4513), .A(n4512), .ZN(n6463) );
  NAND2_X1 U5872 ( .A1(n4515), .A2(n4937), .ZN(n4512) );
  NAND2_X1 U5873 ( .A1(n4514), .A2(n4519), .ZN(n4515) );
  NAND2_X1 U5874 ( .A1(n4520), .A2(n4937), .ZN(n4513) );
  INV_X1 U5875 ( .A(n4515), .ZN(n4516) );
  AOI21_X2 U5876 ( .B1(n6463), .B2(n6462), .A(n4272), .ZN(n6621) );
  OR2_X1 U5877 ( .A1(n4918), .A2(n4919), .ZN(n4519) );
  NAND4_X1 U5878 ( .A1(n4754), .A2(n4755), .A3(n4797), .A4(n4827), .ZN(n5226)
         );
  INV_X1 U5879 ( .A(n5226), .ZN(n5198) );
  NAND2_X1 U5880 ( .A1(n7034), .A2(n4535), .ZN(n4521) );
  NAND2_X1 U5881 ( .A1(n5172), .A2(n5174), .ZN(n7272) );
  NAND2_X2 U5882 ( .A1(n6744), .A2(n5041), .ZN(n6923) );
  NAND2_X1 U5883 ( .A1(n6621), .A2(n6622), .ZN(n6620) );
  AOI21_X1 U5884 ( .B1(n8357), .B2(n8354), .A(n8353), .ZN(n8392) );
  NAND2_X2 U5885 ( .A1(n8371), .A2(n5383), .ZN(n8413) );
  AND2_X2 U5886 ( .A1(n7195), .A2(n4791), .ZN(n7274) );
  NAND2_X1 U5887 ( .A1(n5071), .A2(n4543), .ZN(n4541) );
  NAND2_X1 U5888 ( .A1(n5161), .A2(n4551), .ZN(n4550) );
  OAI21_X1 U5889 ( .B1(n5161), .B2(n4552), .A(n4551), .ZN(n5241) );
  NAND3_X1 U5890 ( .A1(n7702), .A2(n7704), .A3(n7865), .ZN(n4568) );
  NAND2_X1 U5891 ( .A1(n4569), .A2(n4312), .ZN(n5304) );
  NAND2_X1 U5892 ( .A1(n5345), .A2(n4574), .ZN(n4572) );
  NAND2_X1 U5893 ( .A1(n5345), .A2(n4578), .ZN(n4573) );
  NAND2_X1 U5894 ( .A1(n5345), .A2(n5344), .ZN(n5363) );
  NAND2_X1 U5895 ( .A1(n8888), .A2(n4584), .ZN(n4581) );
  NAND2_X1 U5896 ( .A1(n4581), .A2(n4582), .ZN(n8872) );
  NAND2_X2 U5897 ( .A1(n4583), .A2(n5960), .ZN(n8917) );
  NAND2_X1 U5898 ( .A1(n8888), .A2(n8889), .ZN(n4583) );
  NOR2_X1 U5899 ( .A1(n5957), .A2(n5960), .ZN(n4588) );
  NAND2_X1 U5900 ( .A1(n8888), .A2(n5949), .ZN(n8919) );
  OAI21_X2 U5901 ( .B1(n7529), .B2(n4591), .A(n4589), .ZN(n7545) );
  NAND2_X1 U5902 ( .A1(n8950), .A2(n6024), .ZN(n8865) );
  OAI21_X1 U5903 ( .B1(n6898), .B2(n4600), .A(n4596), .ZN(n7126) );
  NAND2_X2 U5904 ( .A1(n5735), .A2(n4280), .ZN(n7182) );
  NAND2_X4 U5905 ( .A1(n6160), .A2(n4607), .ZN(n6870) );
  NOR2_X2 U5906 ( .A1(n5829), .A2(n5532), .ZN(n5548) );
  AND2_X2 U5907 ( .A1(n4716), .A2(n5633), .ZN(n5758) );
  NAND2_X1 U5908 ( .A1(n7424), .A2(n4617), .ZN(n4616) );
  INV_X1 U5909 ( .A(n8676), .ZN(n4620) );
  OAI21_X1 U5910 ( .B1(n7424), .B2(n7397), .A(n8210), .ZN(n8100) );
  NAND2_X1 U5911 ( .A1(n8306), .A2(n4623), .ZN(n4622) );
  NAND2_X1 U5912 ( .A1(n7397), .A2(n8210), .ZN(n4623) );
  NAND2_X1 U5913 ( .A1(n4627), .A2(n8642), .ZN(n4626) );
  NAND2_X1 U5914 ( .A1(n9565), .A2(n4640), .ZN(n4639) );
  NAND3_X1 U5915 ( .A1(n4639), .A2(n4637), .A3(n8194), .ZN(n7301) );
  NAND2_X1 U5916 ( .A1(n4651), .A2(n4650), .ZN(n8119) );
  NAND2_X1 U5917 ( .A1(n8506), .A2(n4652), .ZN(n4651) );
  OR2_X1 U5918 ( .A1(n8506), .A2(n8510), .ZN(n4660) );
  INV_X1 U5919 ( .A(n8741), .ZN(n4663) );
  NAND2_X1 U5920 ( .A1(n4668), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4665) );
  NAND2_X1 U5921 ( .A1(n4855), .A2(n4667), .ZN(n4666) );
  OAI21_X2 U5922 ( .B1(n4668), .B2(n4667), .A(n4666), .ZN(n4911) );
  NAND2_X1 U5923 ( .A1(n4670), .A2(n4669), .ZN(n6131) );
  OAI21_X1 U5924 ( .B1(n7019), .B2(n4674), .A(n4672), .ZN(n7227) );
  NAND2_X1 U5925 ( .A1(n9198), .A2(n4680), .ZN(n4679) );
  OAI21_X1 U5926 ( .B1(n9198), .B2(n4681), .A(n4680), .ZN(n9156) );
  NAND2_X1 U5927 ( .A1(n9127), .A2(n4695), .ZN(n4694) );
  NAND2_X1 U5928 ( .A1(n7410), .A2(n4710), .ZN(n4708) );
  NAND2_X1 U5929 ( .A1(n4708), .A2(n4709), .ZN(n7469) );
  NAND3_X1 U5930 ( .A1(n5633), .A2(n4716), .A3(n5516), .ZN(n6063) );
  AND2_X2 U5931 ( .A1(n5510), .A2(n5511), .ZN(n4716) );
  NAND2_X1 U5932 ( .A1(n4717), .A2(n4718), .ZN(n6490) );
  NAND3_X1 U5933 ( .A1(n6484), .A2(n6483), .A3(n8284), .ZN(n4717) );
  NAND2_X1 U5934 ( .A1(n6799), .A2(n4721), .ZN(n4724) );
  NAND2_X1 U5935 ( .A1(n8297), .A2(n4725), .ZN(n6971) );
  AND2_X2 U5936 ( .A1(n4724), .A2(n6972), .ZN(n7090) );
  OR2_X1 U5937 ( .A1(n8519), .A2(n4732), .ZN(n4726) );
  NAND2_X1 U5938 ( .A1(n8519), .A2(n4730), .ZN(n4729) );
  INV_X1 U5939 ( .A(n8487), .ZN(n4732) );
  NAND2_X1 U5940 ( .A1(n8519), .A2(n8530), .ZN(n8518) );
  OAI21_X1 U5941 ( .B1(n8637), .B2(n4736), .A(n4734), .ZN(n4733) );
  NAND2_X1 U5942 ( .A1(n8777), .A2(n8481), .ZN(n4744) );
  NAND2_X1 U5943 ( .A1(n8587), .A2(n4748), .ZN(n4745) );
  NAND2_X1 U5944 ( .A1(n4745), .A2(n4746), .ZN(n8539) );
  NAND2_X1 U5945 ( .A1(n4797), .A2(n4796), .ZN(n4914) );
  NAND2_X1 U5946 ( .A1(n4797), .A2(n4311), .ZN(n4756) );
  NAND2_X1 U5947 ( .A1(n8818), .A2(n4759), .ZN(n4758) );
  NAND2_X1 U5948 ( .A1(n4758), .A2(n4761), .ZN(n7423) );
  NAND3_X1 U5949 ( .A1(n4845), .A2(n4767), .A3(n4844), .ZN(n6441) );
  AND2_X1 U5950 ( .A1(n4847), .A2(n4846), .ZN(n4767) );
  NAND2_X1 U5951 ( .A1(n5452), .A2(n4770), .ZN(n4808) );
  OAI21_X1 U5952 ( .B1(n6775), .B2(n4775), .A(n4773), .ZN(n6776) );
  AND2_X1 U5953 ( .A1(n6716), .A2(n6712), .ZN(n6713) );
  CLKBUF_X1 U5954 ( .A(n8371), .Z(n8372) );
  OR2_X1 U5955 ( .A1(n6996), .A2(n7803), .ZN(n6997) );
  NAND2_X1 U5956 ( .A1(n6889), .A2(n6882), .ZN(n6730) );
  NAND2_X1 U5957 ( .A1(n6485), .A2(n6450), .ZN(n8142) );
  NAND2_X1 U5958 ( .A1(n9216), .A2(n9057), .ZN(n9058) );
  AOI22_X1 U5959 ( .A1(n7469), .A2(n7814), .B1(n9328), .B2(n8964), .ZN(n7502)
         );
  OR2_X1 U5960 ( .A1(n8641), .A2(n8480), .ZN(n4780) );
  OR2_X1 U5961 ( .A1(n7260), .A2(n7290), .ZN(n4781) );
  OR2_X1 U5962 ( .A1(n9220), .A2(n9204), .ZN(n4783) );
  NOR2_X1 U5963 ( .A1(n7056), .A2(n8433), .ZN(n4784) );
  AND2_X1 U5964 ( .A1(n5070), .A2(n5052), .ZN(n4785) );
  AND4_X1 U5965 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n9175)
         );
  AND2_X1 U5966 ( .A1(n5658), .A2(n5657), .ZN(n4786) );
  AND2_X1 U5967 ( .A1(n5504), .A2(n5503), .ZN(n4787) );
  OR2_X1 U5968 ( .A1(n8658), .A2(n8477), .ZN(n4788) );
  NAND2_X1 U5969 ( .A1(n6372), .A2(n9627), .ZN(n6373) );
  AND2_X1 U5970 ( .A1(n4899), .A2(n4898), .ZN(n4789) );
  OR2_X1 U5971 ( .A1(n8611), .A2(n8601), .ZN(n4790) );
  XNOR2_X1 U5972 ( .A(n8601), .B(n5348), .ZN(n8346) );
  NOR2_X1 U5973 ( .A1(n5174), .A2(n5173), .ZN(n4791) );
  NOR2_X1 U5974 ( .A1(n8290), .A2(n8689), .ZN(n4792) );
  INV_X1 U5975 ( .A(n8643), .ZN(n8492) );
  AND4_X1 U5976 ( .A1(n4802), .A2(n4801), .A3(n4800), .A4(n4799), .ZN(n4803)
         );
  INV_X1 U5977 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5053) );
  NAND2_X1 U5978 ( .A1(n4868), .A2(n4869), .ZN(n4872) );
  NOR2_X1 U5979 ( .A1(n6248), .A2(n8114), .ZN(n8115) );
  AND2_X1 U5980 ( .A1(n5221), .A2(n5220), .ZN(n5222) );
  OR2_X1 U5981 ( .A1(n5139), .A2(n4820), .ZN(n5206) );
  OR2_X1 U5982 ( .A1(n6982), .A2(n6981), .ZN(n7052) );
  INV_X1 U5983 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4804) );
  AND2_X1 U5984 ( .A1(n8922), .A2(n8918), .ZN(n5957) );
  INV_X1 U5985 ( .A(n8331), .ZN(n5523) );
  INV_X1 U5986 ( .A(n7783), .ZN(n9076) );
  INV_X1 U5987 ( .A(n5156), .ZN(n5160) );
  INV_X1 U5988 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5507) );
  INV_X1 U5989 ( .A(n5004), .ZN(n5005) );
  OR2_X1 U5990 ( .A1(n5349), .A2(n8384), .ZN(n5372) );
  OR2_X1 U5991 ( .A1(n5336), .A2(n8348), .ZN(n5349) );
  OAI22_X1 U5992 ( .A1(n8531), .A2(n8695), .B1(n8495), .B2(n8494), .ZN(n8496)
         );
  NAND2_X1 U5993 ( .A1(n8752), .A2(n8561), .ZN(n8527) );
  INV_X1 U5994 ( .A(n5061), .ZN(n4817) );
  OR2_X1 U5995 ( .A1(n8703), .A2(n6782), .ZN(n6982) );
  NAND2_X1 U5996 ( .A1(n4805), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4852) );
  AND2_X1 U5997 ( .A1(n5833), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5860) );
  INV_X1 U5998 ( .A(n6607), .ZN(n5595) );
  AND2_X1 U5999 ( .A1(n5813), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5833) );
  AND3_X1 U6000 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_REG3_REG_20__SCAN_IN), 
        .A3(n5911), .ZN(n5928) );
  OR2_X1 U6001 ( .A1(n5780), .A2(n5779), .ZN(n5795) );
  OR2_X1 U6002 ( .A1(n5701), .A2(n5700), .ZN(n5719) );
  AND2_X1 U6003 ( .A1(n7781), .A2(n7864), .ZN(n9082) );
  OR2_X1 U6004 ( .A1(n6955), .A2(n9519), .ZN(n6956) );
  OR2_X1 U6005 ( .A1(n6837), .A2(n6840), .ZN(n6955) );
  NAND2_X1 U6006 ( .A1(n5163), .A2(n5162), .ZN(n5179) );
  INV_X1 U6007 ( .A(n5083), .ZN(n5087) );
  NOR2_X1 U6008 ( .A1(n5381), .A2(n5380), .ZN(n5382) );
  NOR2_X1 U6009 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  OR2_X1 U6010 ( .A1(n8396), .A2(n8695), .ZN(n8416) );
  OR2_X1 U6011 ( .A1(n8396), .A2(n8693), .ZN(n8414) );
  AND2_X1 U6012 ( .A1(n5438), .A2(n5497), .ZN(n8513) );
  INV_X1 U6013 ( .A(n8496), .ZN(n8497) );
  AND2_X1 U6014 ( .A1(n8210), .A2(n8209), .ZN(n8304) );
  OR2_X1 U6015 ( .A1(n9568), .A2(n9567), .ZN(n9570) );
  INV_X1 U6016 ( .A(n7084), .ZN(n9684) );
  INV_X1 U6017 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4834) );
  AND2_X1 U6018 ( .A1(n6083), .A2(n6084), .ZN(n8862) );
  NAND2_X1 U6019 ( .A1(n8902), .A2(n8903), .ZN(n5989) );
  AND2_X1 U6020 ( .A1(n5860), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5879) );
  NOR2_X1 U6021 ( .A1(n5742), .A2(n5741), .ZN(n5762) );
  NAND2_X1 U6022 ( .A1(n5893), .A2(n5892), .ZN(n8935) );
  INV_X1 U6023 ( .A(n9258), .ZN(n9091) );
  NAND2_X1 U6024 ( .A1(n9269), .A2(n9135), .ZN(n7767) );
  INV_X1 U6025 ( .A(n6768), .ZN(n6875) );
  AND3_X1 U6026 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5639) );
  OR2_X1 U6027 ( .A1(n7716), .A2(n6495), .ZN(n9376) );
  AND2_X1 U6028 ( .A1(n5221), .A2(n5185), .ZN(n5218) );
  AND2_X1 U6029 ( .A1(n5146), .A2(n5120), .ZN(n5144) );
  INV_X1 U6030 ( .A(n8408), .ZN(n8410) );
  AND2_X1 U6031 ( .A1(n5402), .A2(n5401), .ZN(n8561) );
  AND4_X1 U6032 ( .A1(n5178), .A2(n5177), .A3(n5176), .A4(n5175), .ZN(n7438)
         );
  NAND2_X1 U6033 ( .A1(n6410), .A2(n8705), .ZN(n8699) );
  AND2_X1 U6034 ( .A1(n5460), .A2(n5459), .ZN(n9590) );
  AND2_X1 U6035 ( .A1(n5072), .A2(n5057), .ZN(n7325) );
  NAND2_X1 U6036 ( .A1(n8938), .A2(n8935), .ZN(n8880) );
  MUX2_X1 U6037 ( .A(n7827), .B(n7826), .S(n7825), .Z(n7872) );
  AND4_X1 U6038 ( .A1(n5969), .A2(n5968), .A3(n5967), .A4(n5966), .ZN(n9190)
         );
  AND4_X1 U6039 ( .A1(n5838), .A2(n5837), .A3(n5836), .A4(n5835), .ZN(n7537)
         );
  AND4_X1 U6040 ( .A1(n5767), .A2(n5766), .A3(n5765), .A4(n5764), .ZN(n7210)
         );
  INV_X1 U6041 ( .A(n6227), .ZN(n9498) );
  NAND2_X1 U6042 ( .A1(n9077), .A2(n7782), .ZN(n9133) );
  OR2_X1 U6043 ( .A1(n9430), .A2(n6166), .ZN(n9237) );
  OR2_X1 U6044 ( .A1(n9335), .A2(n6159), .ZN(n9209) );
  INV_X1 U6045 ( .A(n9237), .ZN(n9415) );
  OR2_X1 U6046 ( .A1(n6552), .A2(n7869), .ZN(n9542) );
  OR2_X1 U6047 ( .A1(n6096), .A2(n6095), .ZN(n6558) );
  AND2_X1 U6048 ( .A1(n5481), .A2(n8705), .ZN(n8422) );
  INV_X1 U6049 ( .A(n8561), .ZN(n8486) );
  INV_X1 U6050 ( .A(n6485), .ZN(n8440) );
  OR2_X1 U6051 ( .A1(n6385), .A2(n6405), .ZN(n9713) );
  OR2_X1 U6052 ( .A1(n6385), .A2(n6363), .ZN(n9698) );
  CLKBUF_X1 U6053 ( .A(n9604), .Z(n9625) );
  INV_X1 U6054 ( .A(n6705), .ZN(n6991) );
  INV_X1 U6055 ( .A(n8914), .ZN(n8960) );
  OR2_X1 U6056 ( .A1(n9430), .A2(n6872), .ZN(n9247) );
  OR2_X1 U6057 ( .A1(n6558), .A2(n6557), .ZN(n9559) );
  OR2_X1 U6058 ( .A1(n6558), .A2(n6548), .ZN(n9548) );
  INV_X1 U6059 ( .A(n9503), .ZN(n9504) );
  NOR2_X1 U6060 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n4794) );
  NOR2_X1 U6061 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n4793) );
  NAND2_X1 U6062 ( .A1(n4860), .A2(n4795), .ZN(n4893) );
  INV_X1 U6063 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4798) );
  NOR2_X1 U6064 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n4802) );
  NOR2_X1 U6065 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n4801) );
  NOR2_X1 U6066 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4800) );
  NOR2_X1 U6067 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4799) );
  INV_X1 U6068 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4805) );
  INV_X1 U6069 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4806) );
  NAND2_X1 U6070 ( .A1(n4808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4809) );
  MUX2_X1 U6071 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4809), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n4811) );
  INV_X1 U6072 ( .A(n4810), .ZN(n8846) );
  NAND2_X1 U6073 ( .A1(n4900), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4826) );
  NAND2_X1 U6074 ( .A1(n4248), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4825) );
  NAND2_X1 U6075 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n4938) );
  INV_X1 U6076 ( .A(n4938), .ZN(n4813) );
  NAND2_X1 U6077 ( .A1(n4813), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n4959) );
  INV_X1 U6078 ( .A(n4959), .ZN(n4814) );
  NAND2_X1 U6079 ( .A1(n4814), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n4979) );
  INV_X1 U6080 ( .A(n4979), .ZN(n4815) );
  NAND2_X1 U6081 ( .A1(n4815), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5023) );
  NAND2_X1 U6082 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n4816) );
  NAND2_X1 U6083 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n4818) );
  INV_X1 U6084 ( .A(n5127), .ZN(n4819) );
  NAND2_X1 U6085 ( .A1(n4819), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5137) );
  INV_X1 U6086 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5136) );
  INV_X1 U6087 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n4820) );
  NAND2_X1 U6088 ( .A1(n5139), .A2(n4820), .ZN(n4821) );
  AND2_X1 U6089 ( .A1(n5206), .A2(n4821), .ZN(n7384) );
  NAND2_X1 U6090 ( .A1(n4250), .A2(n7384), .ZN(n4824) );
  AND2_X4 U6091 ( .A1(n4822), .A2(n8854), .ZN(n5314) );
  NAND2_X1 U6092 ( .A1(n5314), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n4823) );
  INV_X1 U6093 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4827) );
  INV_X1 U6094 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4829) );
  NAND2_X1 U6095 ( .A1(n4835), .A2(n4829), .ZN(n4838) );
  INV_X1 U6096 ( .A(n4838), .ZN(n4832) );
  INV_X1 U6097 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4831) );
  NAND2_X1 U6098 ( .A1(n4832), .A2(n4831), .ZN(n4833) );
  NAND2_X2 U6099 ( .A1(n8114), .A2(n6366), .ZN(n4865) );
  INV_X1 U6100 ( .A(n4835), .ZN(n4836) );
  NAND2_X1 U6101 ( .A1(n4836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4837) );
  MUX2_X1 U6102 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4837), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n4839) );
  NAND2_X1 U6103 ( .A1(n4839), .A2(n4838), .ZN(n8282) );
  INV_X1 U6104 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U6105 ( .A1(n5198), .A2(n4840), .ZN(n4841) );
  INV_X1 U6106 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4842) );
  NAND2_X1 U6107 ( .A1(n8282), .A2(n4864), .ZN(n5493) );
  NOR2_X1 U6108 ( .A1(n7449), .A2(n6421), .ZN(n7275) );
  NAND2_X1 U6109 ( .A1(n5314), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4845) );
  NAND2_X1 U6110 ( .A1(n4265), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4844) );
  NAND2_X1 U6111 ( .A1(n4881), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U6112 ( .A1(n4900), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4846) );
  NAND2_X1 U6113 ( .A1(n6441), .A2(n8122), .ZN(n4871) );
  INV_X1 U6114 ( .A(n4871), .ZN(n4868) );
  NAND2_X1 U6115 ( .A1(n5457), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4848) );
  MUX2_X1 U6116 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4848), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n4851) );
  INV_X1 U6117 ( .A(n4849), .ZN(n4850) );
  OAI21_X1 U6118 ( .B1(n4849), .B2(n8845), .A(P2_IR_REG_28__SCAN_IN), .ZN(
        n4853) );
  AND2_X1 U6120 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4856) );
  NAND2_X1 U6121 ( .A1(n4911), .A2(n4856), .ZN(n5556) );
  NAND3_X1 U6122 ( .A1(n4857), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n4858) );
  NAND2_X1 U6123 ( .A1(n5556), .A2(n4858), .ZN(n4889) );
  INV_X1 U6124 ( .A(SI_1_), .ZN(n4859) );
  XNOR2_X1 U6125 ( .A(n4889), .B(n4859), .ZN(n4888) );
  MUX2_X1 U6126 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4911), .Z(n4887) );
  XNOR2_X1 U6127 ( .A(n4888), .B(n4887), .ZN(n6208) );
  INV_X1 U6128 ( .A(n4860), .ZN(n4861) );
  NAND2_X1 U6129 ( .A1(n4912), .A2(n8093), .ZN(n4862) );
  NAND2_X1 U6130 ( .A1(n5486), .A2(n8567), .ZN(n6376) );
  NAND2_X1 U6131 ( .A1(n4865), .A2(n6376), .ZN(n8280) );
  INV_X1 U6132 ( .A(n8280), .ZN(n4866) );
  NAND2_X1 U6133 ( .A1(n4866), .A2(n8114), .ZN(n4867) );
  NAND2_X1 U6134 ( .A1(n8315), .A2(n8282), .ZN(n6364) );
  NAND2_X2 U6135 ( .A1(n4867), .A2(n6364), .ZN(n5060) );
  XNOR2_X1 U6136 ( .A(n6367), .B(n5060), .ZN(n4869) );
  INV_X1 U6137 ( .A(n4869), .ZN(n4870) );
  NAND2_X1 U6138 ( .A1(n4871), .A2(n4870), .ZN(n4880) );
  NAND2_X1 U6139 ( .A1(n4265), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4876) );
  NAND2_X1 U6140 ( .A1(n4250), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U6141 ( .A1(n4900), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4874) );
  NAND2_X1 U6142 ( .A1(n5314), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4873) );
  NAND2_X1 U6143 ( .A1(n6196), .A2(SI_0_), .ZN(n4877) );
  XNOR2_X1 U6144 ( .A(n4877), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8860) );
  MUX2_X1 U6145 ( .A(n8859), .B(n8860), .S(n4878), .Z(n9627) );
  INV_X1 U6146 ( .A(n6368), .ZN(n6442) );
  INV_X1 U6147 ( .A(n4886), .ZN(n8122) );
  NOR2_X1 U6148 ( .A1(n5060), .A2(n9627), .ZN(n4879) );
  AOI21_X1 U6149 ( .B1(n6442), .B2(n8122), .A(n4879), .ZN(n6454) );
  NAND2_X1 U6150 ( .A1(n6453), .A2(n6454), .ZN(n6455) );
  NAND2_X1 U6151 ( .A1(n5314), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U6152 ( .A1(n4251), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U6153 ( .A1(n5418), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4883) );
  NAND2_X1 U6154 ( .A1(n4265), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4882) );
  OR2_X1 U6155 ( .A1(n6485), .A2(n6421), .ZN(n4897) );
  NAND2_X1 U6156 ( .A1(n4888), .A2(n4887), .ZN(n4891) );
  NAND2_X1 U6157 ( .A1(n4889), .A2(SI_1_), .ZN(n4890) );
  NAND2_X1 U6158 ( .A1(n4891), .A2(n4890), .ZN(n4906) );
  INV_X1 U6159 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9751) );
  INV_X1 U6160 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6204) );
  MUX2_X1 U6161 ( .A(n9751), .B(n6204), .S(n4911), .Z(n4907) );
  XNOR2_X1 U6162 ( .A(n4907), .B(SI_2_), .ZN(n4905) );
  XNOR2_X1 U6163 ( .A(n4906), .B(n4905), .ZN(n6203) );
  NAND2_X1 U6164 ( .A1(n4252), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n4896) );
  NOR2_X1 U6165 ( .A1(n4860), .A2(n8845), .ZN(n4892) );
  MUX2_X1 U6166 ( .A(n8845), .B(n4892), .S(P2_IR_REG_2__SCAN_IN), .Z(n4894) );
  NAND2_X1 U6167 ( .A1(n4912), .A2(n7310), .ZN(n4895) );
  XNOR2_X1 U6168 ( .A(n6450), .B(n5060), .ZN(n4898) );
  INV_X1 U6169 ( .A(n4897), .ZN(n4899) );
  AOI21_X2 U6170 ( .B1(n4266), .B2(n6428), .A(n4789), .ZN(n6348) );
  NAND2_X1 U6171 ( .A1(n6244), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U6172 ( .A1(n5314), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n4903) );
  NAND2_X1 U6173 ( .A1(n5418), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4902) );
  AND4_X2 U6174 ( .A1(n4904), .A2(n4903), .A3(n4902), .A4(n4901), .ZN(n6488)
         );
  OR2_X1 U6175 ( .A1(n6488), .A2(n6421), .ZN(n4918) );
  INV_X2 U6176 ( .A(n5060), .ZN(n5417) );
  NAND2_X1 U6177 ( .A1(n4906), .A2(n4905), .ZN(n4910) );
  INV_X1 U6178 ( .A(n4907), .ZN(n4908) );
  NAND2_X1 U6179 ( .A1(n4908), .A2(SI_2_), .ZN(n4909) );
  INV_X1 U6180 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6211) );
  INV_X1 U6181 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6202) );
  MUX2_X1 U6182 ( .A(n6211), .B(n6202), .S(n4911), .Z(n4926) );
  XNOR2_X1 U6183 ( .A(n4926), .B(SI_3_), .ZN(n4924) );
  XNOR2_X1 U6184 ( .A(n4925), .B(n4924), .ZN(n6210) );
  NAND2_X1 U6185 ( .A1(n4252), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U6186 ( .A1(n4893), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4913) );
  MUX2_X1 U6187 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4913), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n4915) );
  AND2_X1 U6188 ( .A1(n4915), .A2(n4914), .ZN(n8006) );
  NAND2_X1 U6189 ( .A1(n4912), .A2(n8006), .ZN(n4916) );
  XNOR2_X1 U6190 ( .A(n5417), .B(n8720), .ZN(n4919) );
  XNOR2_X1 U6191 ( .A(n4918), .B(n4919), .ZN(n6347) );
  NAND2_X1 U6192 ( .A1(n4248), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U6193 ( .A1(n5314), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n4922) );
  NAND2_X1 U6194 ( .A1(n5418), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4921) );
  OAI21_X1 U6195 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n4938), .ZN(n6476) );
  INV_X1 U6196 ( .A(n6476), .ZN(n6437) );
  NAND2_X1 U6197 ( .A1(n4251), .A2(n6437), .ZN(n4920) );
  OR2_X1 U6198 ( .A1(n6628), .A2(n6421), .ZN(n4936) );
  NAND2_X1 U6199 ( .A1(n4925), .A2(n4924), .ZN(n4929) );
  INV_X1 U6200 ( .A(n4926), .ZN(n4927) );
  NAND2_X1 U6201 ( .A1(n4927), .A2(SI_3_), .ZN(n4928) );
  INV_X1 U6202 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6198) );
  INV_X1 U6203 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4931) );
  MUX2_X1 U6204 ( .A(n6198), .B(n4931), .S(n4930), .Z(n4947) );
  XNOR2_X1 U6205 ( .A(n4947), .B(SI_4_), .ZN(n4945) );
  XNOR2_X1 U6206 ( .A(n4946), .B(n4945), .ZN(n6197) );
  NAND2_X1 U6207 ( .A1(n4253), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n4934) );
  NAND2_X1 U6208 ( .A1(n4914), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4932) );
  XNOR2_X1 U6209 ( .A(n4932), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U6210 ( .A1(n4912), .A2(n7340), .ZN(n4933) );
  OAI211_X1 U6211 ( .C1(n4944), .C2(n6197), .A(n4934), .B(n4933), .ZN(n6480)
         );
  XNOR2_X1 U6212 ( .A(n5417), .B(n6480), .ZN(n4935) );
  OAI21_X1 U6213 ( .B1(n4936), .B2(n4935), .A(n4937), .ZN(n6434) );
  NAND2_X1 U6214 ( .A1(n4248), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4943) );
  NAND2_X1 U6215 ( .A1(n5418), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4942) );
  INV_X1 U6216 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U6217 ( .A1(n4938), .A2(n8073), .ZN(n4939) );
  AND2_X1 U6218 ( .A1(n4959), .A2(n4939), .ZN(n6644) );
  NAND2_X1 U6219 ( .A1(n4250), .A2(n6644), .ZN(n4941) );
  NAND2_X1 U6220 ( .A1(n5314), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n4940) );
  NOR2_X1 U6221 ( .A1(n8696), .A2(n6421), .ZN(n4957) );
  INV_X4 U6222 ( .A(n4944), .ZN(n8116) );
  NAND2_X1 U6223 ( .A1(n4946), .A2(n4945), .ZN(n4950) );
  INV_X1 U6224 ( .A(n4947), .ZN(n4948) );
  NAND2_X1 U6225 ( .A1(n4948), .A2(SI_4_), .ZN(n4949) );
  MUX2_X1 U6226 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n4930), .Z(n4971) );
  XNOR2_X1 U6227 ( .A(n4970), .B(n4968), .ZN(n6199) );
  NAND2_X1 U6228 ( .A1(n8116), .A2(n6199), .ZN(n4954) );
  NAND2_X1 U6229 ( .A1(n4253), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n4953) );
  NOR2_X1 U6230 ( .A1(n4914), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n4967) );
  OR2_X1 U6231 ( .A1(n4967), .A2(n8845), .ZN(n4951) );
  XNOR2_X1 U6232 ( .A(n4951), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8080) );
  NAND2_X1 U6233 ( .A1(n4912), .A2(n8080), .ZN(n4952) );
  XNOR2_X1 U6234 ( .A(n6778), .B(n5060), .ZN(n4955) );
  XNOR2_X1 U6235 ( .A(n4957), .B(n4955), .ZN(n6462) );
  INV_X1 U6236 ( .A(n4955), .ZN(n4956) );
  NAND2_X1 U6237 ( .A1(n4248), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4964) );
  NAND2_X1 U6238 ( .A1(n5418), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4963) );
  INV_X1 U6239 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4958) );
  NAND2_X1 U6240 ( .A1(n4959), .A2(n4958), .ZN(n4960) );
  AND2_X1 U6241 ( .A1(n4979), .A2(n4960), .ZN(n8704) );
  NAND2_X1 U6242 ( .A1(n4250), .A2(n8704), .ZN(n4962) );
  NAND2_X1 U6243 ( .A1(n5314), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n4961) );
  NOR2_X1 U6244 ( .A1(n6788), .A2(n6421), .ZN(n4976) );
  NAND2_X1 U6245 ( .A1(n4967), .A2(n4966), .ZN(n5015) );
  NAND2_X1 U6246 ( .A1(n5015), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4991) );
  XNOR2_X1 U6247 ( .A(n4965), .B(n4991), .ZN(n7985) );
  NAND2_X1 U6248 ( .A1(n4970), .A2(n4969), .ZN(n4973) );
  NAND2_X1 U6249 ( .A1(n4971), .A2(SI_5_), .ZN(n4972) );
  MUX2_X1 U6250 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7577), .Z(n4988) );
  XNOR2_X1 U6251 ( .A(n9649), .B(n5348), .ZN(n4975) );
  NOR2_X1 U6252 ( .A1(n4976), .A2(n4975), .ZN(n4977) );
  AOI21_X1 U6253 ( .B1(n4976), .B2(n4975), .A(n4977), .ZN(n6622) );
  INV_X1 U6254 ( .A(n4977), .ZN(n4978) );
  NAND2_X1 U6255 ( .A1(n5418), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6256 ( .A1(n4248), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4983) );
  INV_X1 U6257 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7963) );
  NAND2_X1 U6258 ( .A1(n4979), .A2(n7963), .ZN(n4980) );
  AND2_X1 U6259 ( .A1(n5023), .A2(n4980), .ZN(n6781) );
  NAND2_X1 U6260 ( .A1(n4250), .A2(n6781), .ZN(n4982) );
  NAND2_X1 U6261 ( .A1(n5314), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n4981) );
  NOR2_X1 U6262 ( .A1(n8694), .A2(n6421), .ZN(n4997) );
  INV_X1 U6263 ( .A(n4985), .ZN(n4986) );
  NAND2_X1 U6264 ( .A1(n4987), .A2(n4986), .ZN(n4990) );
  NAND2_X1 U6265 ( .A1(n4988), .A2(SI_6_), .ZN(n4989) );
  MUX2_X1 U6266 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n7577), .Z(n5007) );
  XNOR2_X1 U6267 ( .A(n5006), .B(n5004), .ZN(n6216) );
  NAND2_X1 U6268 ( .A1(n6216), .A2(n8116), .ZN(n4995) );
  NAND2_X1 U6269 ( .A1(n4991), .A2(n4965), .ZN(n4992) );
  NAND2_X1 U6270 ( .A1(n4992), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4993) );
  XNOR2_X1 U6271 ( .A(n4993), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7334) );
  AOI22_X1 U6272 ( .A1(n4252), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n4912), .B2(
        n7334), .ZN(n4994) );
  NAND2_X1 U6273 ( .A1(n4995), .A2(n4994), .ZN(n6782) );
  XNOR2_X1 U6274 ( .A(n6782), .B(n5348), .ZN(n4996) );
  XNOR2_X1 U6275 ( .A(n4997), .B(n4996), .ZN(n6653) );
  INV_X1 U6276 ( .A(n4996), .ZN(n4999) );
  INV_X1 U6277 ( .A(n4997), .ZN(n4998) );
  NAND2_X1 U6278 ( .A1(n6244), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5003) );
  NAND2_X1 U6279 ( .A1(n5314), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5002) );
  XNOR2_X1 U6280 ( .A(n5023), .B(P2_REG3_REG_8__SCAN_IN), .ZN(n6810) );
  NAND2_X1 U6281 ( .A1(n4250), .A2(n6810), .ZN(n5001) );
  NAND2_X1 U6282 ( .A1(n5418), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5000) );
  NOR2_X1 U6283 ( .A1(n6966), .A2(n6421), .ZN(n5020) );
  NAND2_X1 U6284 ( .A1(n5006), .A2(n5005), .ZN(n5009) );
  NAND2_X1 U6285 ( .A1(n5007), .A2(SI_7_), .ZN(n5008) );
  INV_X1 U6286 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9805) );
  INV_X1 U6287 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5010) );
  MUX2_X1 U6288 ( .A(n9805), .B(n5010), .S(n7577), .Z(n5012) );
  INV_X1 U6289 ( .A(SI_8_), .ZN(n5011) );
  INV_X1 U6290 ( .A(n5012), .ZN(n5013) );
  NAND2_X1 U6291 ( .A1(n5013), .A2(SI_8_), .ZN(n5014) );
  XNOR2_X1 U6292 ( .A(n5044), .B(n5042), .ZN(n6220) );
  NAND2_X1 U6293 ( .A1(n6220), .A2(n8116), .ZN(n5018) );
  NAND2_X1 U6294 ( .A1(n5097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5016) );
  XNOR2_X1 U6295 ( .A(n5016), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7331) );
  AOI22_X1 U6296 ( .A1(n4253), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4912), .B2(
        n7331), .ZN(n5017) );
  NAND2_X1 U6297 ( .A1(n5018), .A2(n5017), .ZN(n6981) );
  XNOR2_X1 U6298 ( .A(n6981), .B(n5060), .ZN(n5019) );
  XOR2_X1 U6299 ( .A(n5020), .B(n5019), .Z(n6691) );
  NAND2_X1 U6300 ( .A1(n6244), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5028) );
  NAND2_X1 U6301 ( .A1(n5314), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5027) );
  INV_X1 U6302 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5022) );
  INV_X1 U6303 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5021) );
  OAI21_X1 U6304 ( .B1(n5023), .B2(n5022), .A(n5021), .ZN(n5024) );
  AND2_X1 U6305 ( .A1(n5024), .A2(n5061), .ZN(n7055) );
  NAND2_X1 U6306 ( .A1(n4251), .A2(n7055), .ZN(n5026) );
  NAND2_X1 U6307 ( .A1(n5418), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5025) );
  NOR2_X1 U6308 ( .A1(n6965), .A2(n6421), .ZN(n5039) );
  OR2_X1 U6309 ( .A1(n5044), .A2(n5042), .ZN(n5029) );
  NAND2_X1 U6310 ( .A1(n5029), .A2(n5045), .ZN(n5035) );
  INV_X1 U6311 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6230) );
  INV_X1 U6312 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6228) );
  MUX2_X1 U6313 ( .A(n6230), .B(n6228), .S(n7577), .Z(n5031) );
  INV_X1 U6314 ( .A(SI_9_), .ZN(n5030) );
  INV_X1 U6315 ( .A(n5031), .ZN(n5032) );
  NAND2_X1 U6316 ( .A1(n5032), .A2(SI_9_), .ZN(n5033) );
  INV_X1 U6317 ( .A(n5046), .ZN(n5034) );
  NAND2_X1 U6318 ( .A1(n6226), .A2(n8116), .ZN(n5037) );
  OAI21_X1 U6319 ( .B1(n5097), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5054) );
  XNOR2_X1 U6320 ( .A(n5054), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7328) );
  AOI22_X1 U6321 ( .A1(n4252), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4912), .B2(
        n7328), .ZN(n5036) );
  XNOR2_X1 U6322 ( .A(n7056), .B(n5348), .ZN(n5038) );
  NOR2_X1 U6323 ( .A1(n5038), .A2(n5039), .ZN(n5040) );
  AOI21_X1 U6324 ( .B1(n5039), .B2(n5038), .A(n5040), .ZN(n6745) );
  INV_X1 U6325 ( .A(n5040), .ZN(n5041) );
  INV_X1 U6326 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6238) );
  INV_X1 U6327 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6236) );
  MUX2_X1 U6328 ( .A(n6238), .B(n6236), .S(n7577), .Z(n5050) );
  INV_X1 U6329 ( .A(SI_10_), .ZN(n5049) );
  INV_X1 U6330 ( .A(n5050), .ZN(n5051) );
  NAND2_X1 U6331 ( .A1(n5051), .A2(SI_10_), .ZN(n5052) );
  XNOR2_X1 U6332 ( .A(n5069), .B(n4785), .ZN(n6235) );
  NAND2_X1 U6333 ( .A1(n6235), .A2(n8116), .ZN(n5059) );
  NAND2_X1 U6334 ( .A1(n5054), .A2(n5053), .ZN(n5055) );
  NAND2_X1 U6335 ( .A1(n5055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5056) );
  NAND2_X1 U6336 ( .A1(n5056), .A2(n5095), .ZN(n5072) );
  OR2_X1 U6337 ( .A1(n5056), .A2(n5095), .ZN(n5057) );
  AOI22_X1 U6338 ( .A1(n4253), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4912), .B2(
        n7325), .ZN(n5058) );
  NAND2_X1 U6339 ( .A1(n5059), .A2(n5058), .ZN(n9676) );
  XNOR2_X1 U6340 ( .A(n9676), .B(n5348), .ZN(n5067) );
  INV_X1 U6341 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7931) );
  NAND2_X1 U6342 ( .A1(n5061), .A2(n7931), .ZN(n5062) );
  AND2_X1 U6343 ( .A1(n5103), .A2(n5062), .ZN(n9575) );
  NAND2_X1 U6344 ( .A1(n4250), .A2(n9575), .ZN(n5066) );
  NAND2_X1 U6345 ( .A1(n6244), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5065) );
  NAND2_X1 U6346 ( .A1(n5314), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U6347 ( .A1(n5418), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5063) );
  NOR2_X1 U6348 ( .A1(n6980), .A2(n6421), .ZN(n5068) );
  XNOR2_X1 U6349 ( .A(n5067), .B(n5068), .ZN(n6922) );
  INV_X1 U6350 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6242) );
  INV_X1 U6351 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6240) );
  MUX2_X1 U6352 ( .A(n6242), .B(n6240), .S(n7577), .Z(n5084) );
  XNOR2_X1 U6353 ( .A(n5088), .B(n5083), .ZN(n6239) );
  NAND2_X1 U6354 ( .A1(n6239), .A2(n8116), .ZN(n5075) );
  NAND2_X1 U6355 ( .A1(n5072), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5073) );
  XNOR2_X1 U6356 ( .A(n5073), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7347) );
  AOI22_X1 U6357 ( .A1(n4253), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n4912), .B2(
        n7347), .ZN(n5074) );
  NAND2_X1 U6358 ( .A1(n5075), .A2(n5074), .ZN(n7084) );
  XNOR2_X1 U6359 ( .A(n9684), .B(n5348), .ZN(n5080) );
  NAND2_X1 U6360 ( .A1(n5418), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5079) );
  NAND2_X1 U6361 ( .A1(n4248), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5078) );
  XNOR2_X1 U6362 ( .A(n5103), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n7036) );
  NAND2_X1 U6363 ( .A1(n4251), .A2(n7036), .ZN(n5077) );
  NAND2_X1 U6364 ( .A1(n5314), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5076) );
  NOR2_X1 U6365 ( .A1(n7118), .A2(n6421), .ZN(n5082) );
  XNOR2_X1 U6366 ( .A(n5080), .B(n5082), .ZN(n7034) );
  INV_X1 U6367 ( .A(n5080), .ZN(n5081) );
  INV_X1 U6368 ( .A(n5084), .ZN(n5085) );
  INV_X1 U6369 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6254) );
  INV_X1 U6370 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6252) );
  MUX2_X1 U6371 ( .A(n6254), .B(n6252), .S(n7577), .Z(n5090) );
  INV_X1 U6372 ( .A(SI_12_), .ZN(n5089) );
  NAND2_X1 U6373 ( .A1(n5090), .A2(n5089), .ZN(n5113) );
  INV_X1 U6374 ( .A(n5090), .ZN(n5091) );
  NAND2_X1 U6375 ( .A1(n5091), .A2(SI_12_), .ZN(n5092) );
  XNOR2_X1 U6376 ( .A(n5115), .B(n5114), .ZN(n6251) );
  NAND2_X1 U6377 ( .A1(n6251), .A2(n8116), .ZN(n5100) );
  INV_X1 U6378 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5093) );
  NAND4_X1 U6379 ( .A1(n5095), .A2(n5053), .A3(n5094), .A4(n5093), .ZN(n5096)
         );
  NOR2_X1 U6380 ( .A1(n5097), .A2(n5096), .ZN(n5122) );
  OR2_X1 U6381 ( .A1(n5122), .A2(n8845), .ZN(n5098) );
  XNOR2_X1 U6382 ( .A(n5098), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7917) );
  AOI22_X1 U6383 ( .A1(n4252), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n4912), .B2(
        n7917), .ZN(n5099) );
  XNOR2_X1 U6384 ( .A(n7107), .B(n5348), .ZN(n5109) );
  NAND2_X1 U6385 ( .A1(n5418), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6386 ( .A1(n6244), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5107) );
  INV_X1 U6387 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5102) );
  INV_X1 U6388 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5101) );
  OAI21_X1 U6389 ( .B1(n5103), .B2(n5102), .A(n5101), .ZN(n5104) );
  AND2_X1 U6390 ( .A1(n5104), .A2(n5127), .ZN(n7116) );
  NAND2_X1 U6391 ( .A1(n4250), .A2(n7116), .ZN(n5106) );
  NAND2_X1 U6392 ( .A1(n5314), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5105) );
  NOR2_X1 U6393 ( .A1(n7087), .A2(n6421), .ZN(n5110) );
  XNOR2_X1 U6394 ( .A(n5109), .B(n5110), .ZN(n7114) );
  INV_X1 U6395 ( .A(n5109), .ZN(n5112) );
  INV_X1 U6396 ( .A(n5110), .ZN(n5111) );
  INV_X1 U6397 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6343) );
  INV_X1 U6398 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5116) );
  MUX2_X1 U6399 ( .A(n6343), .B(n5116), .S(n7577), .Z(n5118) );
  INV_X1 U6400 ( .A(SI_13_), .ZN(n5117) );
  NAND2_X1 U6401 ( .A1(n5118), .A2(n5117), .ZN(n5146) );
  INV_X1 U6402 ( .A(n5118), .ZN(n5119) );
  NAND2_X1 U6403 ( .A1(n5119), .A2(SI_13_), .ZN(n5120) );
  XNOR2_X1 U6404 ( .A(n5145), .B(n5144), .ZN(n6310) );
  NAND2_X1 U6405 ( .A1(n6310), .A2(n8116), .ZN(n5125) );
  NAND2_X1 U6406 ( .A1(n5122), .A2(n5121), .ZN(n5123) );
  NAND2_X1 U6407 ( .A1(n5123), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5149) );
  XNOR2_X1 U6408 ( .A(n5149), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7350) );
  AOI22_X1 U6409 ( .A1(n4253), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n4912), .B2(
        n7350), .ZN(n5124) );
  XNOR2_X1 U6410 ( .A(n8820), .B(n5417), .ZN(n5133) );
  NAND2_X1 U6411 ( .A1(n4248), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U6412 ( .A1(n5418), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5131) );
  INV_X1 U6413 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5126) );
  NAND2_X1 U6414 ( .A1(n5127), .A2(n5126), .ZN(n5128) );
  AND2_X1 U6415 ( .A1(n5137), .A2(n5128), .ZN(n7104) );
  NAND2_X1 U6416 ( .A1(n4251), .A2(n7104), .ZN(n5130) );
  NAND2_X1 U6417 ( .A1(n5314), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5129) );
  NOR2_X1 U6418 ( .A1(n7302), .A2(n6421), .ZN(n5135) );
  XNOR2_X1 U6419 ( .A(n5133), .B(n5135), .ZN(n7078) );
  INV_X1 U6420 ( .A(n5133), .ZN(n5134) );
  NAND2_X1 U6421 ( .A1(n5418), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5143) );
  NAND2_X1 U6422 ( .A1(n4265), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6423 ( .A1(n5137), .A2(n5136), .ZN(n5138) );
  AND2_X1 U6424 ( .A1(n5139), .A2(n5138), .ZN(n7299) );
  NAND2_X1 U6425 ( .A1(n4251), .A2(n7299), .ZN(n5141) );
  NAND2_X1 U6426 ( .A1(n5314), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5140) );
  NAND4_X1 U6427 ( .A1(n5143), .A2(n5142), .A3(n5141), .A4(n5140), .ZN(n8428)
         );
  AND2_X1 U6428 ( .A1(n8428), .A2(n8122), .ZN(n5154) );
  INV_X1 U6429 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6345) );
  INV_X1 U6430 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9759) );
  MUX2_X1 U6431 ( .A(n6345), .B(n9759), .S(n7577), .Z(n5157) );
  XNOR2_X1 U6432 ( .A(n5161), .B(n5156), .ZN(n6344) );
  NAND2_X1 U6433 ( .A1(n6344), .A2(n8116), .ZN(n5152) );
  NAND2_X1 U6434 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  NAND2_X1 U6435 ( .A1(n5150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5167) );
  XNOR2_X1 U6436 ( .A(n5167), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8053) );
  AOI22_X1 U6437 ( .A1(n4252), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n4912), .B2(
        n8053), .ZN(n5151) );
  XNOR2_X1 U6438 ( .A(n8812), .B(n5348), .ZN(n5153) );
  NOR2_X1 U6439 ( .A1(n5153), .A2(n5154), .ZN(n5173) );
  AOI21_X1 U6440 ( .B1(n5154), .B2(n5153), .A(n5173), .ZN(n7197) );
  INV_X1 U6441 ( .A(n5173), .ZN(n5155) );
  NAND2_X1 U6442 ( .A1(n7195), .A2(n5155), .ZN(n5172) );
  INV_X1 U6443 ( .A(n5157), .ZN(n5158) );
  NAND2_X1 U6444 ( .A1(n5158), .A2(SI_14_), .ZN(n5159) );
  INV_X1 U6445 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6565) );
  INV_X1 U6446 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6563) );
  MUX2_X1 U6447 ( .A(n6565), .B(n6563), .S(n7577), .Z(n5163) );
  INV_X1 U6448 ( .A(SI_15_), .ZN(n5162) );
  INV_X1 U6449 ( .A(n5163), .ZN(n5164) );
  NAND2_X1 U6450 ( .A1(n5164), .A2(SI_15_), .ZN(n5165) );
  NAND2_X1 U6451 ( .A1(n6562), .A2(n8116), .ZN(n5171) );
  NAND2_X1 U6452 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  NAND2_X1 U6453 ( .A1(n5168), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5169) );
  XNOR2_X1 U6454 ( .A(n5169), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7354) );
  AOI22_X1 U6455 ( .A1(n4252), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n4912), .B2(
        n7354), .ZN(n5170) );
  XNOR2_X1 U6456 ( .A(n7386), .B(n5060), .ZN(n5174) );
  NAND2_X1 U6457 ( .A1(n4900), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6458 ( .A1(n6244), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5177) );
  XNOR2_X1 U6459 ( .A(n5206), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n7448) );
  NAND2_X1 U6460 ( .A1(n4251), .A2(n7448), .ZN(n5176) );
  NAND2_X1 U6461 ( .A1(n5314), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5175) );
  NOR2_X1 U6462 ( .A1(n7438), .A2(n6421), .ZN(n5190) );
  INV_X1 U6463 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9838) );
  INV_X1 U6464 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6599) );
  MUX2_X1 U6465 ( .A(n9838), .B(n6599), .S(n7577), .Z(n5183) );
  INV_X1 U6466 ( .A(SI_16_), .ZN(n5182) );
  NAND2_X1 U6467 ( .A1(n5183), .A2(n5182), .ZN(n5221) );
  INV_X1 U6468 ( .A(n5183), .ZN(n5184) );
  NAND2_X1 U6469 ( .A1(n5184), .A2(SI_16_), .ZN(n5185) );
  XNOR2_X1 U6470 ( .A(n5225), .B(n5218), .ZN(n6598) );
  NAND2_X1 U6471 ( .A1(n6598), .A2(n8116), .ZN(n5188) );
  OR2_X1 U6472 ( .A1(n4264), .A2(n8845), .ZN(n5186) );
  XNOR2_X1 U6473 ( .A(n5186), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7884) );
  AOI22_X1 U6474 ( .A1(n4253), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n4912), .B2(
        n7884), .ZN(n5187) );
  XNOR2_X1 U6475 ( .A(n8802), .B(n5348), .ZN(n5189) );
  NOR2_X1 U6476 ( .A1(n5189), .A2(n5190), .ZN(n5191) );
  AOI21_X1 U6477 ( .B1(n5190), .B2(n5189), .A(n5191), .ZN(n7446) );
  INV_X1 U6478 ( .A(n5191), .ZN(n5192) );
  NAND2_X1 U6479 ( .A1(n5225), .A2(n5218), .ZN(n5193) );
  NAND2_X1 U6480 ( .A1(n5193), .A2(n5221), .ZN(n5195) );
  INV_X1 U6481 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6604) );
  INV_X1 U6482 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5194) );
  MUX2_X1 U6483 ( .A(n6604), .B(n5194), .S(n7577), .Z(n5216) );
  XNOR2_X1 U6484 ( .A(n5216), .B(SI_17_), .ZN(n5220) );
  NAND2_X1 U6485 ( .A1(n6566), .A2(n8116), .ZN(n5201) );
  NOR2_X1 U6486 ( .A1(n5196), .A2(n8845), .ZN(n5197) );
  MUX2_X1 U6487 ( .A(n8845), .B(n5197), .S(P2_IR_REG_17__SCAN_IN), .Z(n5199)
         );
  OR2_X1 U6488 ( .A1(n5199), .A2(n5198), .ZN(n8016) );
  INV_X1 U6489 ( .A(n8016), .ZN(n8020) );
  AOI22_X1 U6490 ( .A1(n4252), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n4912), .B2(
        n8020), .ZN(n5200) );
  XNOR2_X1 U6491 ( .A(n8799), .B(n5348), .ZN(n5212) );
  NAND2_X1 U6492 ( .A1(n4265), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6493 ( .A1(n5314), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5210) );
  INV_X1 U6494 ( .A(n5206), .ZN(n5203) );
  AND2_X1 U6495 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n5202) );
  NAND2_X1 U6496 ( .A1(n5203), .A2(n5202), .ZN(n5231) );
  INV_X1 U6497 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5205) );
  INV_X1 U6498 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5204) );
  OAI21_X1 U6499 ( .B1(n5206), .B2(n5205), .A(n5204), .ZN(n5207) );
  AND2_X1 U6500 ( .A1(n5231), .A2(n5207), .ZN(n7404) );
  NAND2_X1 U6501 ( .A1(n4250), .A2(n7404), .ZN(n5209) );
  NAND2_X1 U6502 ( .A1(n4900), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5208) );
  NOR2_X1 U6503 ( .A1(n7425), .A2(n6421), .ZN(n5213) );
  XNOR2_X1 U6504 ( .A(n5212), .B(n5213), .ZN(n7436) );
  INV_X1 U6505 ( .A(n5212), .ZN(n5215) );
  INV_X1 U6506 ( .A(n5213), .ZN(n5214) );
  INV_X1 U6507 ( .A(n5216), .ZN(n5217) );
  NAND2_X1 U6508 ( .A1(n5217), .A2(SI_17_), .ZN(n5219) );
  INV_X1 U6509 ( .A(n5219), .ZN(n5223) );
  MUX2_X1 U6510 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7577), .Z(n5242) );
  XNOR2_X1 U6511 ( .A(n5242), .B(SI_18_), .ZN(n5240) );
  XNOR2_X1 U6512 ( .A(n5241), .B(n5240), .ZN(n6601) );
  NAND2_X1 U6513 ( .A1(n6601), .A2(n8116), .ZN(n5229) );
  NAND2_X1 U6514 ( .A1(n5226), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5227) );
  XNOR2_X1 U6515 ( .A(n5227), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8446) );
  AOI22_X1 U6516 ( .A1(n4253), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4912), .B2(
        n8446), .ZN(n5228) );
  XNOR2_X1 U6517 ( .A(n8792), .B(n5348), .ZN(n5238) );
  NAND2_X1 U6518 ( .A1(n4248), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6519 ( .A1(n4900), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5235) );
  INV_X1 U6520 ( .A(n5231), .ZN(n5230) );
  NAND2_X1 U6521 ( .A1(n5230), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5252) );
  INV_X1 U6522 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9777) );
  NAND2_X1 U6523 ( .A1(n5231), .A2(n9777), .ZN(n5232) );
  AND2_X1 U6524 ( .A1(n5252), .A2(n5232), .ZN(n8672) );
  NAND2_X1 U6525 ( .A1(n4251), .A2(n8672), .ZN(n5234) );
  NAND2_X1 U6526 ( .A1(n5314), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5233) );
  NAND4_X1 U6527 ( .A1(n5236), .A2(n5235), .A3(n5234), .A4(n5233), .ZN(n8662)
         );
  NAND2_X1 U6528 ( .A1(n8662), .A2(n8122), .ZN(n5237) );
  XNOR2_X1 U6529 ( .A(n5238), .B(n5237), .ZN(n7496) );
  INV_X1 U6530 ( .A(n5237), .ZN(n5239) );
  AOI22_X2 U6531 ( .A1(n7495), .A2(n7496), .B1(n5239), .B2(n5238), .ZN(n8357)
         );
  NAND2_X1 U6532 ( .A1(n5242), .A2(SI_18_), .ZN(n5243) );
  INV_X1 U6533 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6665) );
  INV_X1 U6534 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6667) );
  MUX2_X1 U6535 ( .A(n6665), .B(n6667), .S(n7577), .Z(n5246) );
  INV_X1 U6536 ( .A(SI_19_), .ZN(n5245) );
  NAND2_X1 U6537 ( .A1(n5246), .A2(n5245), .ZN(n5262) );
  INV_X1 U6538 ( .A(n5246), .ZN(n5247) );
  NAND2_X1 U6539 ( .A1(n5247), .A2(SI_19_), .ZN(n5248) );
  NAND2_X1 U6540 ( .A1(n5262), .A2(n5248), .ZN(n5263) );
  XNOR2_X1 U6541 ( .A(n5264), .B(n5263), .ZN(n6664) );
  NAND2_X1 U6542 ( .A1(n6664), .A2(n8116), .ZN(n5250) );
  AOI22_X1 U6543 ( .A1(n4252), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n4912), .B2(
        n8567), .ZN(n5249) );
  XNOR2_X1 U6544 ( .A(n8658), .B(n5348), .ZN(n5261) );
  INV_X1 U6545 ( .A(n5261), .ZN(n5259) );
  NAND2_X1 U6546 ( .A1(n5418), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U6547 ( .A1(n4248), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5256) );
  INV_X1 U6548 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5251) );
  NAND2_X1 U6549 ( .A1(n5252), .A2(n5251), .ZN(n5253) );
  AND2_X1 U6550 ( .A1(n5274), .A2(n5253), .ZN(n8656) );
  NAND2_X1 U6551 ( .A1(n4251), .A2(n8656), .ZN(n5255) );
  NAND2_X1 U6552 ( .A1(n5314), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5254) );
  OR2_X1 U6553 ( .A1(n8477), .A2(n6421), .ZN(n5260) );
  INV_X1 U6554 ( .A(n5260), .ZN(n5258) );
  NAND2_X1 U6555 ( .A1(n5259), .A2(n5258), .ZN(n8354) );
  INV_X1 U6556 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6726) );
  INV_X1 U6557 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6724) );
  MUX2_X1 U6558 ( .A(n6726), .B(n6724), .S(n7577), .Z(n5266) );
  INV_X1 U6559 ( .A(SI_20_), .ZN(n5265) );
  NAND2_X1 U6560 ( .A1(n5266), .A2(n5265), .ZN(n5286) );
  INV_X1 U6561 ( .A(n5266), .ZN(n5267) );
  NAND2_X1 U6562 ( .A1(n5267), .A2(SI_20_), .ZN(n5268) );
  XNOR2_X1 U6563 ( .A(n5285), .B(n5284), .ZN(n6723) );
  NAND2_X1 U6564 ( .A1(n6723), .A2(n8116), .ZN(n5270) );
  NAND2_X1 U6565 ( .A1(n4253), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5269) );
  XNOR2_X1 U6566 ( .A(n8783), .B(n5417), .ZN(n5281) );
  NAND2_X1 U6567 ( .A1(n4900), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5272) );
  NAND2_X1 U6568 ( .A1(n6244), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5271) );
  AND2_X1 U6569 ( .A1(n5272), .A2(n5271), .ZN(n5279) );
  INV_X1 U6570 ( .A(n5274), .ZN(n5273) );
  NAND2_X1 U6571 ( .A1(n5273), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5290) );
  INV_X1 U6572 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U6573 ( .A1(n5274), .A2(n8394), .ZN(n5275) );
  NAND2_X1 U6574 ( .A1(n5290), .A2(n5275), .ZN(n8393) );
  OR2_X1 U6575 ( .A1(n8393), .A2(n5276), .ZN(n5278) );
  NAND2_X1 U6576 ( .A1(n5314), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5277) );
  INV_X1 U6577 ( .A(n8480), .ZN(n8663) );
  NAND2_X1 U6578 ( .A1(n8663), .A2(n8122), .ZN(n5280) );
  AOI21_X1 U6579 ( .B1(n5281), .B2(n5280), .A(n5282), .ZN(n8391) );
  NAND2_X1 U6580 ( .A1(n8392), .A2(n8391), .ZN(n8390) );
  INV_X1 U6581 ( .A(n5282), .ZN(n5283) );
  NAND2_X1 U6582 ( .A1(n8390), .A2(n5283), .ZN(n8365) );
  INV_X1 U6583 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6755) );
  INV_X1 U6584 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6753) );
  MUX2_X1 U6585 ( .A(n6755), .B(n6753), .S(n7577), .Z(n5301) );
  XNOR2_X1 U6586 ( .A(n5301), .B(SI_21_), .ZN(n5300) );
  XNOR2_X1 U6587 ( .A(n5299), .B(n5300), .ZN(n6752) );
  NAND2_X1 U6588 ( .A1(n6752), .A2(n8116), .ZN(n5288) );
  NAND2_X1 U6589 ( .A1(n4253), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5287) );
  XNOR2_X1 U6590 ( .A(n8623), .B(n5348), .ZN(n5295) );
  INV_X1 U6591 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6592 ( .A1(n5290), .A2(n5289), .ZN(n5291) );
  AND2_X1 U6593 ( .A1(n5312), .A2(n5291), .ZN(n8631) );
  NAND2_X1 U6594 ( .A1(n8631), .A2(n4250), .ZN(n5294) );
  AOI22_X1 U6595 ( .A1(n6244), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5418), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6596 ( .A1(n5314), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5292) );
  NOR2_X1 U6597 ( .A1(n8610), .A2(n6421), .ZN(n5296) );
  XNOR2_X1 U6598 ( .A(n5295), .B(n5296), .ZN(n8364) );
  NAND2_X1 U6599 ( .A1(n8365), .A2(n8364), .ZN(n8363) );
  INV_X1 U6600 ( .A(n5295), .ZN(n5297) );
  NAND2_X1 U6601 ( .A1(n5297), .A2(n5296), .ZN(n5298) );
  INV_X1 U6602 ( .A(n5301), .ZN(n5302) );
  NAND2_X1 U6603 ( .A1(n5302), .A2(SI_21_), .ZN(n5303) );
  INV_X1 U6604 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8099) );
  INV_X1 U6605 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n6828) );
  MUX2_X1 U6606 ( .A(n8099), .B(n6828), .S(n7577), .Z(n5306) );
  INV_X1 U6607 ( .A(SI_22_), .ZN(n5305) );
  NAND2_X1 U6608 ( .A1(n5306), .A2(n5305), .ZN(n5322) );
  INV_X1 U6609 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U6610 ( .A1(n5307), .A2(SI_22_), .ZN(n5308) );
  NAND2_X1 U6611 ( .A1(n5322), .A2(n5308), .ZN(n5323) );
  XNOR2_X1 U6612 ( .A(n5324), .B(n5323), .ZN(n6826) );
  NAND2_X1 U6613 ( .A1(n6826), .A2(n8116), .ZN(n5310) );
  NAND2_X1 U6614 ( .A1(n4252), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5309) );
  XNOR2_X1 U6615 ( .A(n8774), .B(n5417), .ZN(n5319) );
  INV_X1 U6616 ( .A(n5312), .ZN(n5311) );
  NAND2_X1 U6617 ( .A1(n5311), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5336) );
  INV_X1 U6618 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U6619 ( .A1(n5312), .A2(n8403), .ZN(n5313) );
  NAND2_X1 U6620 ( .A1(n5336), .A2(n5313), .ZN(n8613) );
  OR2_X1 U6621 ( .A1(n8613), .A2(n5276), .ZN(n5317) );
  AOI22_X1 U6622 ( .A1(n4265), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n4900), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6623 ( .A1(n5314), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5315) );
  AND3_X1 U6624 ( .A1(n5317), .A2(n5316), .A3(n5315), .ZN(n8593) );
  INV_X1 U6625 ( .A(n8593), .ZN(n8629) );
  NAND2_X1 U6626 ( .A1(n8629), .A2(n8122), .ZN(n8402) );
  INV_X1 U6627 ( .A(n5318), .ZN(n5320) );
  NAND2_X1 U6628 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  INV_X1 U6629 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5326) );
  INV_X1 U6630 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5325) );
  MUX2_X1 U6631 ( .A(n5326), .B(n5325), .S(n7577), .Z(n5328) );
  INV_X1 U6632 ( .A(SI_23_), .ZN(n5327) );
  NAND2_X1 U6633 ( .A1(n5328), .A2(n5327), .ZN(n5344) );
  INV_X1 U6634 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U6635 ( .A1(n5329), .A2(SI_23_), .ZN(n5330) );
  AND2_X1 U6636 ( .A1(n5344), .A2(n5330), .ZN(n5331) );
  OR2_X1 U6637 ( .A1(n5332), .A2(n5331), .ZN(n5333) );
  NAND2_X1 U6638 ( .A1(n5345), .A2(n5333), .ZN(n7010) );
  NAND2_X1 U6639 ( .A1(n7010), .A2(n8116), .ZN(n5335) );
  NAND2_X1 U6640 ( .A1(n4252), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5334) );
  INV_X1 U6641 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U6642 ( .A1(n5336), .A2(n8348), .ZN(n5337) );
  NAND2_X1 U6643 ( .A1(n5349), .A2(n5337), .ZN(n8597) );
  OR2_X1 U6644 ( .A1(n8597), .A2(n5276), .ZN(n5343) );
  INV_X1 U6645 ( .A(n5314), .ZN(n5501) );
  INV_X1 U6646 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U6647 ( .A1(n4265), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6648 ( .A1(n5418), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5338) );
  OAI211_X1 U6649 ( .C1(n5501), .C2(n5340), .A(n5339), .B(n5338), .ZN(n5341)
         );
  INV_X1 U6650 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U6651 ( .A1(n5343), .A2(n5342), .ZN(n8580) );
  NAND2_X1 U6652 ( .A1(n8580), .A2(n8122), .ZN(n8345) );
  INV_X1 U6653 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7063) );
  INV_X1 U6654 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7065) );
  MUX2_X1 U6655 ( .A(n7063), .B(n7065), .S(n7577), .Z(n5359) );
  XNOR2_X1 U6656 ( .A(n5359), .B(SI_24_), .ZN(n5358) );
  NAND2_X1 U6657 ( .A1(n7062), .A2(n8116), .ZN(n5347) );
  NAND2_X1 U6658 ( .A1(n4253), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5346) );
  XNOR2_X1 U6659 ( .A(n8761), .B(n5348), .ZN(n5354) );
  XNOR2_X1 U6660 ( .A(n5356), .B(n5354), .ZN(n8380) );
  INV_X1 U6661 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8384) );
  NAND2_X1 U6662 ( .A1(n5349), .A2(n8384), .ZN(n5350) );
  NAND2_X1 U6663 ( .A1(n5372), .A2(n5350), .ZN(n8385) );
  INV_X1 U6664 ( .A(n8385), .ZN(n8574) );
  INV_X1 U6665 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9775) );
  NAND2_X1 U6666 ( .A1(n4900), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U6667 ( .A1(n4248), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5351) );
  OAI211_X1 U6668 ( .C1(n9775), .C2(n5501), .A(n5352), .B(n5351), .ZN(n5353)
         );
  AOI21_X1 U6669 ( .B1(n8574), .B2(n4250), .A(n5353), .ZN(n8592) );
  NOR2_X1 U6670 ( .A1(n8592), .A2(n6421), .ZN(n8383) );
  NAND2_X1 U6671 ( .A1(n8380), .A2(n8383), .ZN(n8382) );
  INV_X1 U6672 ( .A(n5354), .ZN(n5355) );
  OR2_X1 U6673 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U6674 ( .A1(n8382), .A2(n5357), .ZN(n8370) );
  INV_X1 U6675 ( .A(n5358), .ZN(n5362) );
  INV_X1 U6676 ( .A(n5359), .ZN(n5360) );
  NAND2_X1 U6677 ( .A1(n5360), .A2(SI_24_), .ZN(n5361) );
  INV_X1 U6678 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7194) );
  INV_X1 U6679 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7191) );
  MUX2_X1 U6680 ( .A(n7194), .B(n7191), .S(n7577), .Z(n5365) );
  INV_X1 U6681 ( .A(SI_25_), .ZN(n5364) );
  NAND2_X1 U6682 ( .A1(n5365), .A2(n5364), .ZN(n5384) );
  INV_X1 U6683 ( .A(n5365), .ZN(n5366) );
  NAND2_X1 U6684 ( .A1(n5366), .A2(SI_25_), .ZN(n5367) );
  NAND2_X1 U6685 ( .A1(n5384), .A2(n5367), .ZN(n5385) );
  NAND2_X1 U6686 ( .A1(n4253), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5368) );
  INV_X1 U6687 ( .A(n5372), .ZN(n5370) );
  NAND2_X1 U6688 ( .A1(n5370), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5395) );
  INV_X1 U6689 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5371) );
  NAND2_X1 U6690 ( .A1(n5372), .A2(n5371), .ZN(n5373) );
  AND2_X1 U6691 ( .A1(n5395), .A2(n5373), .ZN(n8565) );
  NAND2_X1 U6692 ( .A1(n8565), .A2(n4251), .ZN(n5379) );
  INV_X1 U6693 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6694 ( .A1(n4900), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6695 ( .A1(n4248), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5374) );
  OAI211_X1 U6696 ( .C1(n5376), .C2(n5501), .A(n5375), .B(n5374), .ZN(n5377)
         );
  INV_X1 U6697 ( .A(n5377), .ZN(n5378) );
  OR2_X1 U6698 ( .A1(n8424), .A2(n6421), .ZN(n5380) );
  AOI21_X1 U6699 ( .B1(n5381), .B2(n5380), .A(n5382), .ZN(n8373) );
  NAND2_X1 U6700 ( .A1(n8370), .A2(n8373), .ZN(n8371) );
  INV_X1 U6701 ( .A(n5382), .ZN(n5383) );
  INV_X1 U6702 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7224) );
  INV_X1 U6703 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7222) );
  MUX2_X1 U6704 ( .A(n7224), .B(n7222), .S(n7577), .Z(n5388) );
  INV_X1 U6705 ( .A(SI_26_), .ZN(n5387) );
  NAND2_X1 U6706 ( .A1(n5388), .A2(n5387), .ZN(n5409) );
  INV_X1 U6707 ( .A(n5388), .ZN(n5389) );
  NAND2_X1 U6708 ( .A1(n5389), .A2(SI_26_), .ZN(n5390) );
  AND2_X1 U6709 ( .A1(n5409), .A2(n5390), .ZN(n5407) );
  NAND2_X1 U6710 ( .A1(n4252), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5391) );
  XNOR2_X1 U6711 ( .A(n8752), .B(n5417), .ZN(n5404) );
  INV_X1 U6712 ( .A(n5395), .ZN(n5393) );
  NAND2_X1 U6713 ( .A1(n5393), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5437) );
  INV_X1 U6714 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U6715 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  NAND2_X1 U6716 ( .A1(n5437), .A2(n5396), .ZN(n8542) );
  OR2_X1 U6717 ( .A1(n8542), .A2(n5276), .ZN(n5402) );
  INV_X1 U6718 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6719 ( .A1(n5418), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U6720 ( .A1(n4265), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5397) );
  OAI211_X1 U6721 ( .C1(n5399), .C2(n5501), .A(n5398), .B(n5397), .ZN(n5400)
         );
  INV_X1 U6722 ( .A(n5400), .ZN(n5401) );
  NAND2_X1 U6723 ( .A1(n8486), .A2(n8122), .ZN(n5403) );
  NOR2_X1 U6724 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  AOI21_X1 U6725 ( .B1(n5404), .B2(n5403), .A(n5405), .ZN(n8412) );
  INV_X1 U6726 ( .A(n5405), .ZN(n5406) );
  INV_X1 U6727 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7271) );
  INV_X1 U6728 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5411) );
  MUX2_X1 U6729 ( .A(n7271), .B(n5411), .S(n7577), .Z(n5412) );
  INV_X1 U6730 ( .A(SI_27_), .ZN(n9804) );
  NAND2_X1 U6731 ( .A1(n5412), .A2(n9804), .ZN(n5430) );
  INV_X1 U6732 ( .A(n5412), .ZN(n5413) );
  NAND2_X1 U6733 ( .A1(n5413), .A2(SI_27_), .ZN(n5414) );
  AND2_X1 U6734 ( .A1(n5430), .A2(n5414), .ZN(n5428) );
  NAND2_X1 U6735 ( .A1(n4252), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5415) );
  XNOR2_X1 U6736 ( .A(n8746), .B(n5417), .ZN(n5426) );
  XNOR2_X1 U6737 ( .A(n5437), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8524) );
  NAND2_X1 U6738 ( .A1(n8524), .A2(n4250), .ZN(n5424) );
  INV_X1 U6739 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6740 ( .A1(n6244), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6741 ( .A1(n5418), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5419) );
  OAI211_X1 U6742 ( .C1(n5421), .C2(n5501), .A(n5420), .B(n5419), .ZN(n5422)
         );
  INV_X1 U6743 ( .A(n5422), .ZN(n5423) );
  OR2_X1 U6744 ( .A1(n8415), .A2(n6421), .ZN(n5425) );
  NOR2_X1 U6745 ( .A1(n5426), .A2(n5425), .ZN(n5427) );
  AOI21_X1 U6746 ( .B1(n5426), .B2(n5425), .A(n5427), .ZN(n8339) );
  INV_X1 U6747 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8336) );
  INV_X1 U6748 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5431) );
  MUX2_X1 U6749 ( .A(n8336), .B(n5431), .S(n7577), .Z(n7572) );
  XNOR2_X1 U6750 ( .A(n7572), .B(SI_28_), .ZN(n7569) );
  NAND2_X1 U6751 ( .A1(n4253), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5432) );
  INV_X1 U6752 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5435) );
  INV_X1 U6753 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5434) );
  OAI21_X1 U6754 ( .B1(n5437), .B2(n5435), .A(n5434), .ZN(n5438) );
  NAND2_X1 U6755 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n5436) );
  OR2_X1 U6756 ( .A1(n5437), .A2(n5436), .ZN(n5497) );
  NAND2_X1 U6757 ( .A1(n8513), .A2(n4251), .ZN(n5444) );
  INV_X1 U6758 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6759 ( .A1(n6244), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U6760 ( .A1(n4900), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5439) );
  OAI211_X1 U6761 ( .C1(n5441), .C2(n5501), .A(n5440), .B(n5439), .ZN(n5442)
         );
  INV_X1 U6762 ( .A(n5442), .ZN(n5443) );
  NAND2_X1 U6763 ( .A1(n5444), .A2(n5443), .ZN(n8423) );
  NAND2_X1 U6764 ( .A1(n8423), .A2(n8122), .ZN(n5445) );
  XNOR2_X1 U6765 ( .A(n5445), .B(n5348), .ZN(n5484) );
  NAND2_X1 U6766 ( .A1(n5446), .A2(n4834), .ZN(n5447) );
  NAND2_X1 U6767 ( .A1(n5447), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5475) );
  INV_X1 U6768 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U6769 ( .A1(n5475), .A2(n9789), .ZN(n5477) );
  NAND2_X1 U6770 ( .A1(n5477), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5449) );
  INV_X1 U6771 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5448) );
  XNOR2_X1 U6772 ( .A(n5449), .B(n5448), .ZN(n7064) );
  XNOR2_X1 U6773 ( .A(n7064), .B(P2_B_REG_SCAN_IN), .ZN(n5454) );
  NAND2_X1 U6774 ( .A1(n5450), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5451) );
  MUX2_X1 U6775 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5451), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5453) );
  NAND2_X1 U6776 ( .A1(n5453), .A2(n5455), .ZN(n7192) );
  NAND2_X1 U6777 ( .A1(n5454), .A2(n7192), .ZN(n5460) );
  NAND2_X1 U6778 ( .A1(n5455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5456) );
  MUX2_X1 U6779 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5456), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5458) );
  NAND2_X1 U6780 ( .A1(n5458), .A2(n5457), .ZN(n7226) );
  INV_X1 U6781 ( .A(n7226), .ZN(n5459) );
  INV_X1 U6782 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6783 ( .A1(n9590), .A2(n5461), .ZN(n5462) );
  NAND2_X1 U6784 ( .A1(n7064), .A2(n7226), .ZN(n9621) );
  NAND2_X1 U6785 ( .A1(n5462), .A2(n9621), .ZN(n6405) );
  INV_X1 U6786 ( .A(n6405), .ZN(n6363) );
  INV_X1 U6787 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6788 ( .A1(n7226), .A2(n7192), .ZN(n9623) );
  INV_X1 U6789 ( .A(n9623), .ZN(n5463) );
  AOI21_X1 U6790 ( .B1(n9590), .B2(n5464), .A(n5463), .ZN(n6406) );
  NOR4_X1 U6791 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5473) );
  INV_X1 U6792 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n9839) );
  INV_X1 U6793 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9620) );
  INV_X1 U6794 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9619) );
  INV_X1 U6795 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n9618) );
  NAND4_X1 U6796 ( .A1(n9839), .A2(n9620), .A3(n9619), .A4(n9618), .ZN(n5470)
         );
  NOR4_X1 U6797 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n5468) );
  NOR4_X1 U6798 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5467) );
  NOR4_X1 U6799 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5466) );
  NOR4_X1 U6800 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n5465) );
  NAND4_X1 U6801 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n5465), .ZN(n5469)
         );
  NOR4_X1 U6802 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n5470), .A4(n5469), .ZN(n5472) );
  NOR4_X1 U6803 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n5471) );
  NAND3_X1 U6804 ( .A1(n5473), .A2(n5472), .A3(n5471), .ZN(n5474) );
  NAND2_X1 U6805 ( .A1(n9590), .A2(n5474), .ZN(n6361) );
  NAND3_X1 U6806 ( .A1(n6363), .A2(n6406), .A3(n6361), .ZN(n5496) );
  OR2_X1 U6807 ( .A1(n5475), .A2(n9789), .ZN(n5476) );
  NAND2_X1 U6808 ( .A1(n5477), .A2(n5476), .ZN(n6174) );
  NAND2_X1 U6809 ( .A1(n6174), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9624) );
  INV_X1 U6810 ( .A(n9624), .ZN(n5478) );
  NAND2_X1 U6811 ( .A1(n6175), .A2(n5478), .ZN(n9589) );
  OR2_X1 U6812 ( .A1(n5496), .A2(n9589), .ZN(n5491) );
  NOR2_X1 U6813 ( .A1(n4865), .A2(n8282), .ZN(n6417) );
  INV_X1 U6814 ( .A(n6417), .ZN(n5479) );
  OR2_X1 U6815 ( .A1(n5491), .A2(n5479), .ZN(n5481) );
  NAND2_X1 U6816 ( .A1(n8282), .A2(n8567), .ZN(n8319) );
  NOR2_X1 U6817 ( .A1(n4865), .A2(n8319), .ZN(n6362) );
  INV_X1 U6818 ( .A(n6362), .ZN(n5480) );
  NOR3_X1 U6819 ( .A1(n4663), .A2(n5484), .A3(n8406), .ZN(n5482) );
  AOI21_X1 U6820 ( .B1(n4663), .B2(n5484), .A(n5482), .ZN(n5489) );
  NAND3_X1 U6821 ( .A1(n8741), .A2(n8422), .A3(n5484), .ZN(n5483) );
  OAI21_X1 U6822 ( .B1(n8741), .B2(n5484), .A(n5483), .ZN(n5485) );
  NAND2_X1 U6823 ( .A1(n5490), .A2(n5485), .ZN(n5488) );
  INV_X1 U6824 ( .A(n4865), .ZN(n9628) );
  NAND2_X1 U6825 ( .A1(n9628), .A2(n5493), .ZN(n9690) );
  AND2_X1 U6826 ( .A1(n8326), .A2(n8315), .ZN(n6178) );
  OAI21_X1 U6827 ( .B1(n4663), .B2(n8422), .A(n8408), .ZN(n5487) );
  OAI211_X1 U6828 ( .C1(n5490), .C2(n5489), .A(n5488), .B(n5487), .ZN(n5505)
         );
  INV_X1 U6829 ( .A(n8415), .ZN(n8549) );
  OR2_X1 U6830 ( .A1(n5491), .A2(n5493), .ZN(n8396) );
  INV_X1 U6831 ( .A(n6178), .ZN(n6187) );
  OR2_X1 U6832 ( .A1(n6187), .A2(n5492), .ZN(n8695) );
  INV_X1 U6833 ( .A(n8416), .ZN(n8375) );
  AOI22_X1 U6834 ( .A1(n8549), .A2(n8375), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5504) );
  AND2_X1 U6835 ( .A1(n6178), .A2(n5493), .ZN(n6360) );
  INV_X1 U6836 ( .A(n6360), .ZN(n5494) );
  NAND3_X1 U6837 ( .A1(n6175), .A2(n6174), .A3(n5494), .ZN(n5495) );
  AOI21_X1 U6838 ( .B1(n5496), .B2(n9690), .A(n5495), .ZN(n6349) );
  NAND2_X1 U6839 ( .A1(n5496), .A2(n6417), .ZN(n6350) );
  AOI21_X1 U6840 ( .B1(n6349), .B2(n6350), .A(P2_U3152), .ZN(n8398) );
  AND2_X1 U6841 ( .A1(n5492), .A2(n6178), .ZN(n8680) );
  INV_X1 U6842 ( .A(n8680), .ZN(n8693) );
  INV_X1 U6843 ( .A(n8414), .ZN(n8374) );
  INV_X1 U6844 ( .A(n5497), .ZN(n8500) );
  INV_X1 U6845 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U6846 ( .A1(n4248), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5499) );
  NAND2_X1 U6847 ( .A1(n5418), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5498) );
  OAI211_X1 U6848 ( .C1(n5501), .C2(n5500), .A(n5499), .B(n5498), .ZN(n5502)
         );
  AOI21_X1 U6849 ( .B1(n8500), .B2(n4250), .A(n5502), .ZN(n8110) );
  INV_X1 U6850 ( .A(n8110), .ZN(n8507) );
  AOI22_X1 U6851 ( .A1(n8513), .A2(n8398), .B1(n8374), .B2(n8507), .ZN(n5503)
         );
  NAND2_X1 U6852 ( .A1(n5505), .A2(n4787), .ZN(P2_U3222) );
  NOR2_X1 U6853 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5509) );
  NOR2_X1 U6854 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5508) );
  AND4_X2 U6855 ( .A1(n5509), .A2(n5508), .A3(n5670), .A4(n5507), .ZN(n5510)
         );
  NOR2_X1 U6856 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5513) );
  INV_X1 U6857 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5545) );
  INV_X2 U6858 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9864) );
  NAND4_X1 U6859 ( .A1(n5513), .A2(n5512), .A3(n5545), .A4(n9864), .ZN(n5515)
         );
  INV_X1 U6860 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5529) );
  INV_X1 U6861 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5530) );
  NAND4_X1 U6862 ( .A1(n5529), .A2(n5808), .A3(n5530), .A4(n5535), .ZN(n5514)
         );
  INV_X1 U6863 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5517) );
  INV_X1 U6864 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U6865 ( .A1(n4247), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5528) );
  INV_X1 U6866 ( .A(n9367), .ZN(n5524) );
  NAND2_X1 U6867 ( .A1(n5665), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U6868 ( .A1(n5721), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U6869 ( .A1(n5641), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5525) );
  NAND4_X2 U6870 ( .A1(n5528), .A2(n5527), .A3(n5526), .A4(n5525), .ZN(n6575)
         );
  INV_X1 U6871 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U6872 ( .A1(n5805), .A2(n5808), .ZN(n5828) );
  NAND3_X1 U6873 ( .A1(n9864), .A2(n5530), .A3(n5529), .ZN(n5531) );
  OR2_X1 U6874 ( .A1(n5828), .A2(n5531), .ZN(n5532) );
  INV_X1 U6875 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U6876 ( .A1(n5548), .A2(n5533), .ZN(n5551) );
  NAND2_X1 U6877 ( .A1(n5536), .A2(n5535), .ZN(n5534) );
  NAND2_X2 U6878 ( .A1(n5534), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5546) );
  XNOR2_X2 U6879 ( .A(n5546), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6060) );
  NAND2_X2 U6880 ( .A1(n6060), .A2(n7777), .ZN(n6160) );
  NAND2_X1 U6881 ( .A1(n4273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5537) );
  XNOR2_X1 U6882 ( .A(n5537), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6080) );
  INV_X1 U6883 ( .A(n5538), .ZN(n5539) );
  NAND2_X1 U6884 ( .A1(n5539), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5540) );
  MUX2_X1 U6885 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5540), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5542) );
  NAND2_X1 U6886 ( .A1(n5542), .A2(n5541), .ZN(n7067) );
  INV_X1 U6887 ( .A(n7067), .ZN(n6067) );
  NAND2_X1 U6888 ( .A1(n5541), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5543) );
  MUX2_X1 U6889 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5543), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5544) );
  AND2_X1 U6890 ( .A1(n5544), .A2(n4273), .ZN(n6070) );
  NAND3_X1 U6891 ( .A1(n6080), .A2(n6067), .A3(n6070), .ZN(n6092) );
  NAND2_X1 U6892 ( .A1(n5546), .A2(n5545), .ZN(n5547) );
  INV_X1 U6893 ( .A(n5548), .ZN(n5549) );
  NAND2_X1 U6894 ( .A1(n5549), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5550) );
  MUX2_X1 U6895 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5550), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n5552) );
  NAND2_X1 U6896 ( .A1(n5552), .A2(n5551), .ZN(n9033) );
  AND2_X1 U6897 ( .A1(n7777), .A2(n9033), .ZN(n6091) );
  INV_X1 U6898 ( .A(n6091), .ZN(n6061) );
  OR2_X1 U6899 ( .A1(n7875), .A2(n6061), .ZN(n5553) );
  NAND2_X4 U6900 ( .A1(n4249), .A2(n5553), .ZN(n6051) );
  NAND2_X1 U6902 ( .A1(n7577), .A2(SI_0_), .ZN(n5555) );
  INV_X1 U6903 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U6904 ( .A1(n5555), .A2(n5554), .ZN(n5557) );
  AND2_X1 U6905 ( .A1(n5557), .A2(n5556), .ZN(n9370) );
  NAND2_X1 U6906 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n6102) );
  INV_X1 U6907 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n6103) );
  NOR2_X1 U6908 ( .A1(n6102), .A2(n6103), .ZN(n5559) );
  NOR2_X1 U6909 ( .A1(n4278), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5558) );
  AOI21_X1 U6910 ( .B1(n6101), .B2(n5559), .A(n5558), .ZN(n5562) );
  INV_X1 U6911 ( .A(n5560), .ZN(n5561) );
  MUX2_X1 U6912 ( .A(n9370), .B(P1_IR_REG_0__SCAN_IN), .S(n6128), .Z(n6795) );
  INV_X1 U6913 ( .A(n6795), .ZN(n6570) );
  INV_X1 U6914 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6282) );
  OAI22_X1 U6915 ( .A1(n6570), .A2(n6055), .B1(n6282), .B2(n6092), .ZN(n5563)
         );
  NAND2_X1 U6916 ( .A1(n6575), .A2(n5789), .ZN(n5565) );
  AOI22_X1 U6917 ( .A1(n6057), .A2(n6795), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n6125), .ZN(n5564) );
  NAND2_X1 U6918 ( .A1(n5565), .A2(n5564), .ZN(n6401) );
  NAND2_X1 U6919 ( .A1(n6402), .A2(n6401), .ZN(n6400) );
  INV_X1 U6920 ( .A(n6401), .ZN(n5566) );
  NAND2_X1 U6921 ( .A1(n5566), .A2(n6870), .ZN(n5567) );
  NAND2_X1 U6922 ( .A1(n6400), .A2(n5567), .ZN(n7554) );
  NAND2_X1 U6923 ( .A1(n5598), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U6924 ( .A1(n5721), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5569) );
  NAND2_X1 U6925 ( .A1(n5641), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U6926 ( .A1(n8976), .A2(n5789), .ZN(n5576) );
  AND2_X1 U6927 ( .A1(n5571), .A2(n6196), .ZN(n5673) );
  NAND2_X1 U6928 ( .A1(n5673), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U6929 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5572) );
  OR2_X1 U6930 ( .A1(n7568), .A2(n5574), .ZN(n5575) );
  NAND2_X1 U6931 ( .A1(n5576), .A2(n5575), .ZN(n5577) );
  XNOR2_X1 U6932 ( .A(n5577), .B(n5983), .ZN(n5581) );
  NAND2_X1 U6933 ( .A1(n7554), .A2(n5581), .ZN(n5580) );
  NAND2_X1 U6934 ( .A1(n8976), .A2(n5947), .ZN(n5579) );
  OR2_X1 U6935 ( .A1(n7568), .A2(n6055), .ZN(n5578) );
  NAND2_X1 U6936 ( .A1(n5579), .A2(n5578), .ZN(n7557) );
  NAND2_X1 U6937 ( .A1(n5580), .A2(n7557), .ZN(n7556) );
  INV_X1 U6938 ( .A(n7554), .ZN(n5582) );
  INV_X1 U6939 ( .A(n5581), .ZN(n7555) );
  NAND2_X1 U6940 ( .A1(n5582), .A2(n7555), .ZN(n7560) );
  NAND2_X1 U6941 ( .A1(n7556), .A2(n7560), .ZN(n6608) );
  NAND2_X1 U6942 ( .A1(n5665), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5586) );
  NAND2_X1 U6943 ( .A1(n5598), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U6944 ( .A1(n5721), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U6945 ( .A1(n5641), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5583) );
  AND4_X2 U6946 ( .A1(n5586), .A2(n5585), .A3(n5584), .A4(n5583), .ZN(n6133)
         );
  INV_X1 U6947 ( .A(n5674), .ZN(n5590) );
  NAND2_X1 U6948 ( .A1(n5673), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5589) );
  OR2_X1 U6949 ( .A1(n5587), .A2(n5519), .ZN(n5604) );
  XNOR2_X1 U6950 ( .A(n5604), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6284) );
  NAND2_X1 U6951 ( .A1(n6128), .A2(n6284), .ZN(n5588) );
  OAI211_X1 U6952 ( .C1(n5590), .C2(n6203), .A(n5589), .B(n5588), .ZN(n6941)
         );
  OAI22_X1 U6953 ( .A1(n6133), .A2(n6055), .B1(n6937), .B2(n5574), .ZN(n5591)
         );
  XNOR2_X1 U6954 ( .A(n5591), .B(n6870), .ZN(n5593) );
  OAI22_X1 U6955 ( .A1(n6133), .A2(n6051), .B1(n6937), .B2(n6055), .ZN(n5592)
         );
  OR2_X1 U6956 ( .A1(n5593), .A2(n5592), .ZN(n5597) );
  NAND2_X1 U6957 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  NAND2_X1 U6958 ( .A1(n5597), .A2(n5594), .ZN(n6607) );
  NAND2_X1 U6959 ( .A1(n6605), .A2(n5597), .ZN(n6683) );
  NAND2_X1 U6960 ( .A1(n5665), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5602) );
  INV_X1 U6961 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6988) );
  NAND2_X1 U6962 ( .A1(n4247), .A2(n6988), .ZN(n5601) );
  NAND2_X1 U6963 ( .A1(n5721), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U6964 ( .A1(n5641), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U6965 ( .A1(n5673), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5608) );
  INV_X1 U6966 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5603) );
  NAND2_X1 U6967 ( .A1(n5604), .A2(n5603), .ZN(n5605) );
  NAND2_X1 U6968 ( .A1(n5605), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5606) );
  XNOR2_X1 U6969 ( .A(n5606), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U6970 ( .A1(n6128), .A2(n6340), .ZN(n5607) );
  OAI211_X1 U6971 ( .C1(n5590), .C2(n6210), .A(n5608), .B(n5607), .ZN(n6705)
         );
  OAI22_X1 U6972 ( .A1(n6832), .A2(n6055), .B1(n6991), .B2(n5574), .ZN(n5609)
         );
  XNOR2_X1 U6973 ( .A(n5609), .B(n6870), .ZN(n5627) );
  INV_X1 U6974 ( .A(n5627), .ZN(n5610) );
  OAI22_X1 U6975 ( .A1(n6832), .A2(n6051), .B1(n6991), .B2(n6055), .ZN(n5626)
         );
  XNOR2_X1 U6976 ( .A(n5610), .B(n5626), .ZN(n6684) );
  INV_X1 U6977 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5611) );
  XNOR2_X1 U6978 ( .A(n5611), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6839) );
  NAND2_X1 U6979 ( .A1(n4247), .A2(n6839), .ZN(n5615) );
  NAND2_X1 U6980 ( .A1(n5665), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U6981 ( .A1(n5641), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U6982 ( .A1(n5721), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U6983 ( .A1(n5673), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U6984 ( .A1(n5616), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5617) );
  XNOR2_X1 U6985 ( .A(n5617), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U6986 ( .A1(n6128), .A2(n6509), .ZN(n5618) );
  OAI211_X1 U6987 ( .C1(n5590), .C2(n6197), .A(n5619), .B(n5618), .ZN(n6840)
         );
  INV_X1 U6988 ( .A(n6840), .ZN(n9511) );
  XNOR2_X1 U6989 ( .A(n5620), .B(n5983), .ZN(n5625) );
  INV_X1 U6990 ( .A(n5625), .ZN(n5621) );
  OAI22_X1 U6991 ( .A1(n6950), .A2(n6051), .B1(n9511), .B2(n6055), .ZN(n5624)
         );
  NAND2_X1 U6992 ( .A1(n5621), .A2(n5624), .ZN(n5623) );
  AND2_X1 U6993 ( .A1(n6684), .A2(n5623), .ZN(n5622) );
  NAND2_X1 U6994 ( .A1(n6683), .A2(n5622), .ZN(n6817) );
  INV_X1 U6995 ( .A(n5623), .ZN(n5628) );
  XNOR2_X1 U6996 ( .A(n5625), .B(n5624), .ZN(n6716) );
  OR2_X1 U6997 ( .A1(n5627), .A2(n5626), .ZN(n6712) );
  OR2_X1 U6998 ( .A1(n5628), .A2(n6713), .ZN(n6816) );
  NAND2_X1 U6999 ( .A1(n5639), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5663) );
  OAI21_X1 U7000 ( .B1(n5639), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5663), .ZN(
        n6167) );
  INV_X1 U7001 ( .A(n6167), .ZN(n6895) );
  NAND2_X1 U7002 ( .A1(n4247), .A2(n6895), .ZN(n5632) );
  NAND2_X1 U7003 ( .A1(n5665), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7004 ( .A1(n5641), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7005 ( .A1(n5721), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5629) );
  INV_X1 U7006 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7007 ( .A1(n5674), .A2(n6212), .ZN(n5637) );
  OR2_X1 U7008 ( .A1(n5634), .A2(n5519), .ZN(n5635) );
  XNOR2_X1 U7009 ( .A(n5635), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U7010 ( .A1(n6128), .A2(n9470), .ZN(n5636) );
  OAI22_X1 U7011 ( .A1(n6949), .A2(n6055), .B1(n9527), .B2(n6018), .ZN(n5638)
         );
  XNOR2_X1 U7012 ( .A(n5638), .B(n6870), .ZN(n5661) );
  OAI22_X1 U7013 ( .A1(n6949), .A2(n6051), .B1(n9527), .B2(n6055), .ZN(n5660)
         );
  OR2_X1 U7014 ( .A1(n5661), .A2(n5660), .ZN(n6884) );
  NAND2_X1 U7015 ( .A1(n5665), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5645) );
  AOI21_X1 U7016 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5640) );
  NOR2_X1 U7017 ( .A1(n5640), .A2(n5639), .ZN(n6958) );
  NAND2_X1 U7018 ( .A1(n4247), .A2(n6958), .ZN(n5644) );
  NAND2_X1 U7019 ( .A1(n5721), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U7020 ( .A1(n5641), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5642) );
  INV_X1 U7021 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9867) );
  NAND2_X1 U7022 ( .A1(n5674), .A2(n6199), .ZN(n5650) );
  MUX2_X1 U7023 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5646), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5648) );
  INV_X1 U7024 ( .A(n5634), .ZN(n5647) );
  NAND2_X1 U7025 ( .A1(n6128), .A2(n9458), .ZN(n5649) );
  OAI22_X1 U7026 ( .A1(n6831), .A2(n6055), .B1(n6135), .B2(n6018), .ZN(n5651)
         );
  XNOR2_X1 U7027 ( .A(n5651), .B(n6870), .ZN(n5656) );
  INV_X1 U7028 ( .A(n5656), .ZN(n6818) );
  OR2_X1 U7029 ( .A1(n6831), .A2(n6051), .ZN(n5653) );
  NAND2_X1 U7030 ( .A1(n9519), .A2(n6043), .ZN(n5652) );
  NAND2_X1 U7031 ( .A1(n5653), .A2(n5652), .ZN(n6820) );
  INV_X1 U7032 ( .A(n6820), .ZN(n5654) );
  NAND2_X1 U7033 ( .A1(n6818), .A2(n5654), .ZN(n5655) );
  AND2_X1 U7034 ( .A1(n6884), .A2(n5655), .ZN(n5658) );
  AND2_X1 U7035 ( .A1(n5656), .A2(n6820), .ZN(n5657) );
  NAND2_X1 U7036 ( .A1(n5661), .A2(n5660), .ZN(n6882) );
  INV_X1 U7037 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5662) );
  NOR2_X1 U7038 ( .A1(n5663), .A2(n5662), .ZN(n5682) );
  AND2_X1 U7039 ( .A1(n5663), .A2(n5662), .ZN(n5664) );
  NOR2_X1 U7040 ( .A1(n5682), .A2(n5664), .ZN(n6873) );
  NAND2_X1 U7041 ( .A1(n4247), .A2(n6873), .ZN(n5669) );
  NAND2_X1 U7042 ( .A1(n5665), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5668) );
  NAND2_X1 U7043 ( .A1(n5641), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U7044 ( .A1(n5721), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5666) );
  OR2_X1 U7045 ( .A1(n6906), .A2(n6051), .ZN(n5678) );
  NAND2_X1 U7046 ( .A1(n5634), .A2(n5670), .ZN(n5688) );
  NAND2_X1 U7047 ( .A1(n5688), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5671) );
  AND2_X1 U7048 ( .A1(n6128), .A2(n6321), .ZN(n5672) );
  AOI21_X1 U7049 ( .B1(n5673), .B2(P2_DATAO_REG_7__SCAN_IN), .A(n5672), .ZN(
        n5676) );
  NAND2_X1 U7050 ( .A1(n6216), .A2(n5674), .ZN(n5675) );
  NAND2_X1 U7051 ( .A1(n5676), .A2(n5675), .ZN(n6768) );
  NAND2_X1 U7052 ( .A1(n6768), .A2(n6043), .ZN(n5677) );
  NAND2_X1 U7053 ( .A1(n5678), .A2(n5677), .ZN(n6728) );
  OAI22_X1 U7054 ( .A1(n6906), .A2(n6055), .B1(n6875), .B2(n6018), .ZN(n5679)
         );
  XNOR2_X1 U7055 ( .A(n5679), .B(n6870), .ZN(n6727) );
  OAI21_X1 U7056 ( .B1(n6730), .B2(n6728), .A(n6727), .ZN(n5681) );
  NAND2_X1 U7057 ( .A1(n6730), .A2(n6728), .ZN(n5680) );
  NAND2_X1 U7058 ( .A1(n5681), .A2(n5680), .ZN(n6898) );
  NAND2_X1 U7059 ( .A1(n5682), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5701) );
  OR2_X1 U7060 ( .A1(n5682), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5683) );
  AND2_X1 U7061 ( .A1(n5701), .A2(n5683), .ZN(n6902) );
  NAND2_X1 U7062 ( .A1(n4247), .A2(n6902), .ZN(n5687) );
  NAND2_X1 U7063 ( .A1(n5665), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U7064 ( .A1(n7588), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7065 ( .A1(n5641), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7066 ( .A1(n6220), .A2(n5894), .ZN(n5691) );
  NAND2_X1 U7067 ( .A1(n5693), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5689) );
  AOI22_X1 U7068 ( .A1(n6025), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n9484), .B2(
        n6128), .ZN(n5690) );
  NAND2_X1 U7069 ( .A1(n5691), .A2(n5690), .ZN(n6999) );
  INV_X1 U7070 ( .A(n6999), .ZN(n9533) );
  OAI22_X1 U7071 ( .A1(n7073), .A2(n6055), .B1(n9533), .B2(n6018), .ZN(n5692)
         );
  XNOR2_X1 U7072 ( .A(n5692), .B(n6870), .ZN(n6899) );
  OAI22_X1 U7073 ( .A1(n7073), .A2(n6051), .B1(n9533), .B2(n6055), .ZN(n6900)
         );
  NAND2_X1 U7074 ( .A1(n6226), .A2(n5894), .ZN(n5699) );
  NOR2_X1 U7075 ( .A1(n5693), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5696) );
  OR2_X1 U7076 ( .A1(n5696), .A2(n5519), .ZN(n5694) );
  INV_X1 U7077 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5695) );
  MUX2_X1 U7078 ( .A(n5694), .B(P1_IR_REG_31__SCAN_IN), .S(n5695), .Z(n5697)
         );
  NAND2_X1 U7079 ( .A1(n5696), .A2(n5695), .ZN(n5737) );
  NAND2_X1 U7080 ( .A1(n5697), .A2(n5737), .ZN(n6227) );
  AOI22_X1 U7081 ( .A1(n6025), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n9498), .B2(
        n6128), .ZN(n5698) );
  NAND2_X1 U7082 ( .A1(n7075), .A2(n6057), .ZN(n5708) );
  INV_X1 U7083 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7084 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  AND2_X1 U7085 ( .A1(n5719), .A2(n5702), .ZN(n7070) );
  NAND2_X1 U7086 ( .A1(n4247), .A2(n7070), .ZN(n5706) );
  NAND2_X1 U7087 ( .A1(n5665), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7088 ( .A1(n7588), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U7089 ( .A1(n5641), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5703) );
  NAND4_X1 U7090 ( .A1(n5706), .A2(n5705), .A3(n5704), .A4(n5703), .ZN(n8969)
         );
  NAND2_X1 U7091 ( .A1(n8969), .A2(n6043), .ZN(n5707) );
  NAND2_X1 U7092 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  XNOR2_X1 U7093 ( .A(n5709), .B(n5983), .ZN(n5710) );
  AOI22_X1 U7094 ( .A1(n7075), .A2(n6043), .B1(n8969), .B2(n5947), .ZN(n5711)
         );
  NAND2_X1 U7095 ( .A1(n5710), .A2(n5711), .ZN(n5715) );
  INV_X1 U7096 ( .A(n5710), .ZN(n5713) );
  INV_X1 U7097 ( .A(n5711), .ZN(n5712) );
  NAND2_X1 U7098 ( .A1(n5713), .A2(n5712), .ZN(n5714) );
  NAND2_X1 U7099 ( .A1(n5715), .A2(n5714), .ZN(n7069) );
  NAND2_X1 U7100 ( .A1(n6235), .A2(n5894), .ZN(n5718) );
  NAND2_X1 U7101 ( .A1(n5737), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5716) );
  XNOR2_X1 U7102 ( .A(n5716), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6589) );
  AOI22_X1 U7103 ( .A1(n6025), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6589), .B2(
        n6128), .ZN(n5717) );
  NAND2_X1 U7104 ( .A1(n5718), .A2(n5717), .ZN(n9388) );
  NAND2_X1 U7105 ( .A1(n9388), .A2(n6057), .ZN(n5727) );
  INV_X1 U7106 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9819) );
  NAND2_X1 U7107 ( .A1(n5719), .A2(n9819), .ZN(n5720) );
  AND2_X1 U7108 ( .A1(n5742), .A2(n5720), .ZN(n9387) );
  NAND2_X1 U7109 ( .A1(n4247), .A2(n9387), .ZN(n5725) );
  NAND2_X1 U7110 ( .A1(n5665), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U7111 ( .A1(n5641), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U7112 ( .A1(n7588), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5722) );
  OR2_X1 U7113 ( .A1(n7023), .A2(n6055), .ZN(n5726) );
  NAND2_X1 U7114 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  XNOR2_X1 U7115 ( .A(n5728), .B(n6870), .ZN(n5731) );
  NAND2_X1 U7116 ( .A1(n9388), .A2(n6043), .ZN(n5730) );
  OR2_X1 U7117 ( .A1(n7023), .A2(n6051), .ZN(n5729) );
  NAND2_X1 U7118 ( .A1(n5730), .A2(n5729), .ZN(n5732) );
  NAND2_X1 U7119 ( .A1(n5731), .A2(n5732), .ZN(n7124) );
  NAND2_X1 U7120 ( .A1(n7126), .A2(n7124), .ZN(n5735) );
  INV_X1 U7121 ( .A(n5731), .ZN(n5734) );
  INV_X1 U7122 ( .A(n5732), .ZN(n5733) );
  NAND2_X1 U7123 ( .A1(n5734), .A2(n5733), .ZN(n7123) );
  NAND2_X1 U7124 ( .A1(n6239), .A2(n5894), .ZN(n5740) );
  OAI21_X1 U7125 ( .B1(n5737), .B2(P1_IR_REG_10__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5738) );
  XNOR2_X1 U7126 ( .A(n5738), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6590) );
  AOI22_X1 U7127 ( .A1(n6025), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6590), .B2(
        n6128), .ZN(n5739) );
  NAND2_X1 U7128 ( .A1(n5740), .A2(n5739), .ZN(n7204) );
  NAND2_X1 U7129 ( .A1(n7204), .A2(n6057), .ZN(n5750) );
  INV_X1 U7130 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5741) );
  AND2_X1 U7131 ( .A1(n5742), .A2(n5741), .ZN(n5743) );
  NOR2_X1 U7132 ( .A1(n5762), .A2(n5743), .ZN(n7186) );
  NAND2_X1 U7133 ( .A1(n4247), .A2(n7186), .ZN(n5748) );
  NAND2_X1 U7134 ( .A1(n5665), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5747) );
  NAND2_X1 U7135 ( .A1(n5641), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U7136 ( .A1(n7588), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5745) );
  OR2_X1 U7137 ( .A1(n9377), .A2(n6055), .ZN(n5749) );
  NAND2_X1 U7138 ( .A1(n5750), .A2(n5749), .ZN(n5751) );
  XNOR2_X1 U7139 ( .A(n5751), .B(n5983), .ZN(n5754) );
  NOR2_X1 U7140 ( .A1(n9377), .A2(n6051), .ZN(n5752) );
  AOI21_X1 U7141 ( .B1(n7204), .B2(n6043), .A(n5752), .ZN(n5753) );
  XNOR2_X1 U7142 ( .A(n5754), .B(n5753), .ZN(n7180) );
  OR2_X1 U7143 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  NAND2_X1 U7144 ( .A1(n6251), .A2(n5894), .ZN(n5761) );
  NOR2_X1 U7145 ( .A1(n5756), .A2(n5519), .ZN(n5757) );
  MUX2_X1 U7146 ( .A(n5519), .B(n5757), .S(P1_IR_REG_12__SCAN_IN), .Z(n5759)
         );
  OR2_X1 U7147 ( .A1(n5759), .A2(n5758), .ZN(n6586) );
  INV_X1 U7148 ( .A(n6586), .ZN(n6674) );
  AOI22_X1 U7149 ( .A1(n6025), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6674), .B2(
        n6128), .ZN(n5760) );
  NAND2_X1 U7150 ( .A1(n9416), .A2(n6057), .ZN(n5769) );
  NAND2_X1 U7151 ( .A1(n5665), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5767) );
  OR2_X1 U7152 ( .A1(n5762), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7153 ( .A1(n5762), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5780) );
  AND2_X1 U7154 ( .A1(n5763), .A2(n5780), .ZN(n9413) );
  NAND2_X1 U7155 ( .A1(n4247), .A2(n9413), .ZN(n5766) );
  NAND2_X1 U7156 ( .A1(n7588), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7157 ( .A1(n5641), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5764) );
  OR2_X1 U7158 ( .A1(n7210), .A2(n6055), .ZN(n5768) );
  NAND2_X1 U7159 ( .A1(n5769), .A2(n5768), .ZN(n5770) );
  XNOR2_X1 U7160 ( .A(n5770), .B(n5983), .ZN(n5773) );
  NOR2_X1 U7161 ( .A1(n7210), .A2(n6051), .ZN(n5771) );
  AOI21_X1 U7162 ( .B1(n9416), .B2(n6043), .A(n5771), .ZN(n5772) );
  XNOR2_X1 U7163 ( .A(n5773), .B(n5772), .ZN(n7287) );
  NAND2_X1 U7164 ( .A1(n5773), .A2(n5772), .ZN(n5774) );
  NAND2_X2 U7165 ( .A1(n7284), .A2(n5774), .ZN(n7370) );
  NAND2_X1 U7166 ( .A1(n6310), .A2(n5894), .ZN(n5778) );
  NAND2_X1 U7167 ( .A1(n5775), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5776) );
  XNOR2_X1 U7168 ( .A(n5776), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6914) );
  AOI22_X1 U7169 ( .A1(n6025), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6914), .B2(
        n6128), .ZN(n5777) );
  NAND2_X1 U7170 ( .A1(n7376), .A2(n6057), .ZN(n5787) );
  NAND2_X1 U7171 ( .A1(n5665), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5785) );
  INV_X1 U7172 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7173 ( .A1(n5780), .A2(n5779), .ZN(n5781) );
  AND2_X1 U7174 ( .A1(n5795), .A2(n5781), .ZN(n7214) );
  NAND2_X1 U7175 ( .A1(n4247), .A2(n7214), .ZN(n5784) );
  NAND2_X1 U7176 ( .A1(n7588), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U7177 ( .A1(n5641), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5782) );
  NAND4_X1 U7178 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n9408)
         );
  NAND2_X1 U7179 ( .A1(n9408), .A2(n6043), .ZN(n5786) );
  NAND2_X1 U7180 ( .A1(n5787), .A2(n5786), .ZN(n5788) );
  XNOR2_X1 U7181 ( .A(n5788), .B(n5983), .ZN(n7368) );
  AND2_X1 U7182 ( .A1(n9408), .A2(n5947), .ZN(n5790) );
  AOI21_X1 U7183 ( .B1(n7376), .B2(n6043), .A(n5790), .ZN(n7367) );
  AND2_X1 U7184 ( .A1(n7368), .A2(n7367), .ZN(n5791) );
  OAI22_X2 U7185 ( .A1(n7370), .A2(n5791), .B1(n7368), .B2(n7367), .ZN(n7529)
         );
  NAND2_X1 U7186 ( .A1(n6344), .A2(n5894), .ZN(n5793) );
  NAND2_X1 U7187 ( .A1(n5829), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5806) );
  XNOR2_X1 U7188 ( .A(n5806), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7166) );
  AOI22_X1 U7189 ( .A1(n6025), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7166), .B2(
        n6128), .ZN(n5792) );
  NAND2_X1 U7190 ( .A1(n9339), .A2(n6057), .ZN(n5802) );
  INV_X1 U7191 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5794) );
  AND2_X1 U7192 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  NOR2_X1 U7193 ( .A1(n5813), .A2(n5796), .ZN(n7466) );
  NAND2_X1 U7194 ( .A1(n4247), .A2(n7466), .ZN(n5800) );
  NAND2_X1 U7195 ( .A1(n5665), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7196 ( .A1(n5641), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7197 ( .A1(n7588), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5797) );
  NAND4_X1 U7198 ( .A1(n5800), .A2(n5799), .A3(n5798), .A4(n5797), .ZN(n8966)
         );
  NAND2_X1 U7199 ( .A1(n8966), .A2(n6043), .ZN(n5801) );
  NAND2_X1 U7200 ( .A1(n5802), .A2(n5801), .ZN(n5803) );
  XNOR2_X1 U7201 ( .A(n5803), .B(n5983), .ZN(n7458) );
  AND2_X1 U7202 ( .A1(n8966), .A2(n5947), .ZN(n5804) );
  AOI21_X1 U7203 ( .B1(n9339), .B2(n6043), .A(n5804), .ZN(n5825) );
  NAND2_X1 U7204 ( .A1(n7458), .A2(n5825), .ZN(n7528) );
  NAND2_X1 U7205 ( .A1(n6562), .A2(n5894), .ZN(n5812) );
  NAND2_X1 U7206 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  NAND2_X1 U7207 ( .A1(n5807), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5809) );
  XNOR2_X1 U7208 ( .A(n5809), .B(n5808), .ZN(n7249) );
  INV_X1 U7209 ( .A(n7249), .ZN(n5810) );
  AOI22_X1 U7210 ( .A1(n6025), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5810), .B2(
        n6128), .ZN(n5811) );
  NAND2_X1 U7211 ( .A1(n9331), .A2(n6043), .ZN(n5820) );
  NOR2_X1 U7212 ( .A1(n5813), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5814) );
  OR2_X1 U7213 ( .A1(n5833), .A2(n5814), .ZN(n7540) );
  INV_X1 U7214 ( .A(n7540), .ZN(n7488) );
  NAND2_X1 U7215 ( .A1(n4247), .A2(n7488), .ZN(n5818) );
  NAND2_X1 U7216 ( .A1(n5665), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5817) );
  NAND2_X1 U7217 ( .A1(n7588), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U7218 ( .A1(n5641), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5815) );
  NAND4_X1 U7219 ( .A1(n5818), .A2(n5817), .A3(n5816), .A4(n5815), .ZN(n8965)
         );
  NAND2_X1 U7220 ( .A1(n8965), .A2(n5947), .ZN(n5819) );
  NAND2_X1 U7221 ( .A1(n5820), .A2(n5819), .ZN(n7535) );
  AND2_X1 U7222 ( .A1(n7528), .A2(n7535), .ZN(n5821) );
  INV_X1 U7223 ( .A(n7535), .ZN(n5827) );
  NAND2_X1 U7224 ( .A1(n9331), .A2(n6057), .ZN(n5823) );
  NAND2_X1 U7225 ( .A1(n8965), .A2(n6043), .ZN(n5822) );
  NAND2_X1 U7226 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  XNOR2_X1 U7227 ( .A(n5824), .B(n5983), .ZN(n5847) );
  INV_X1 U7228 ( .A(n7458), .ZN(n5826) );
  INV_X1 U7229 ( .A(n5825), .ZN(n7457) );
  NAND2_X1 U7230 ( .A1(n5826), .A2(n7457), .ZN(n5846) );
  AND2_X1 U7231 ( .A1(n5847), .A2(n5846), .ZN(n7530) );
  OR2_X1 U7232 ( .A1(n5827), .A2(n7530), .ZN(n7512) );
  NAND2_X1 U7233 ( .A1(n6598), .A2(n5894), .ZN(n5832) );
  OR2_X1 U7234 ( .A1(n5829), .A2(n5828), .ZN(n5855) );
  NAND2_X1 U7235 ( .A1(n5855), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5830) );
  XNOR2_X1 U7236 ( .A(n5830), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8996) );
  AOI22_X1 U7237 ( .A1(n6025), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8996), .B2(
        n6128), .ZN(n5831) );
  NAND2_X1 U7238 ( .A1(n9328), .A2(n6057), .ZN(n5840) );
  NAND2_X1 U7239 ( .A1(n5665), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5838) );
  NOR2_X1 U7240 ( .A1(n5833), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5834) );
  OR2_X1 U7241 ( .A1(n5860), .A2(n5834), .ZN(n7524) );
  INV_X1 U7242 ( .A(n7524), .ZN(n7416) );
  NAND2_X1 U7243 ( .A1(n4247), .A2(n7416), .ZN(n5837) );
  NAND2_X1 U7244 ( .A1(n7588), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U7245 ( .A1(n5641), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5835) );
  OR2_X1 U7246 ( .A1(n7537), .A2(n6055), .ZN(n5839) );
  NAND2_X1 U7247 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  XNOR2_X1 U7248 ( .A(n5841), .B(n6870), .ZN(n5851) );
  NAND2_X1 U7249 ( .A1(n9328), .A2(n6043), .ZN(n5843) );
  OR2_X1 U7250 ( .A1(n7537), .A2(n6051), .ZN(n5842) );
  NAND2_X1 U7251 ( .A1(n5843), .A2(n5842), .ZN(n5852) );
  AND2_X1 U7252 ( .A1(n5851), .A2(n5852), .ZN(n7516) );
  INV_X1 U7253 ( .A(n7516), .ZN(n5844) );
  AND2_X1 U7254 ( .A1(n7512), .A2(n5844), .ZN(n5845) );
  INV_X1 U7255 ( .A(n5846), .ZN(n5850) );
  INV_X1 U7256 ( .A(n5847), .ZN(n5848) );
  AND2_X1 U7257 ( .A1(n5848), .A2(n7528), .ZN(n5849) );
  INV_X1 U7258 ( .A(n5851), .ZN(n5854) );
  INV_X1 U7259 ( .A(n5852), .ZN(n5853) );
  NAND2_X1 U7260 ( .A1(n5854), .A2(n5853), .ZN(n7515) );
  NAND2_X1 U7261 ( .A1(n6566), .A2(n5894), .ZN(n5859) );
  OAI21_X1 U7262 ( .B1(n5855), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5856) );
  OR2_X1 U7263 ( .A1(n5856), .A2(n9864), .ZN(n5857) );
  NAND2_X1 U7264 ( .A1(n5856), .A2(n9864), .ZN(n5875) );
  AND2_X1 U7265 ( .A1(n5857), .A2(n5875), .ZN(n9013) );
  AOI22_X1 U7266 ( .A1(n6025), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9013), .B2(
        n6128), .ZN(n5858) );
  NAND2_X1 U7267 ( .A1(n9323), .A2(n6057), .ZN(n5867) );
  NAND2_X1 U7268 ( .A1(n5665), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5865) );
  NOR2_X1 U7269 ( .A1(n5860), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5861) );
  NOR2_X1 U7270 ( .A1(n5879), .A2(n5861), .ZN(n7551) );
  NAND2_X1 U7271 ( .A1(n4247), .A2(n7551), .ZN(n5864) );
  NAND2_X1 U7272 ( .A1(n7588), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7273 ( .A1(n5641), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5862) );
  NAND4_X1 U7274 ( .A1(n5865), .A2(n5864), .A3(n5863), .A4(n5862), .ZN(n8963)
         );
  NAND2_X1 U7275 ( .A1(n8963), .A2(n6043), .ZN(n5866) );
  NAND2_X1 U7276 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  XNOR2_X1 U7277 ( .A(n5868), .B(n6870), .ZN(n5870) );
  AND2_X1 U7278 ( .A1(n8963), .A2(n5947), .ZN(n5869) );
  AOI21_X1 U7279 ( .B1(n9323), .B2(n6043), .A(n5869), .ZN(n5871) );
  XNOR2_X1 U7280 ( .A(n5870), .B(n5871), .ZN(n7546) );
  NAND2_X1 U7281 ( .A1(n7545), .A2(n7546), .ZN(n5874) );
  INV_X1 U7282 ( .A(n5870), .ZN(n5872) );
  NAND2_X1 U7283 ( .A1(n5872), .A2(n5871), .ZN(n5873) );
  NAND2_X1 U7284 ( .A1(n5874), .A2(n5873), .ZN(n5890) );
  NAND2_X1 U7285 ( .A1(n6601), .A2(n5894), .ZN(n5878) );
  NAND2_X1 U7286 ( .A1(n5875), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5876) );
  XNOR2_X1 U7287 ( .A(n5876), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9025) );
  AOI22_X1 U7288 ( .A1(n6025), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9025), .B2(
        n6128), .ZN(n5877) );
  NAND2_X1 U7289 ( .A1(n9316), .A2(n6057), .ZN(n5886) );
  OR2_X1 U7290 ( .A1(n5879), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5880) );
  NAND2_X1 U7291 ( .A1(n5879), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5910) );
  AND2_X1 U7292 ( .A1(n5880), .A2(n5910), .ZN(n8943) );
  NAND2_X1 U7293 ( .A1(n4247), .A2(n8943), .ZN(n5884) );
  NAND2_X1 U7294 ( .A1(n5665), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U7295 ( .A1(n5641), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5882) );
  NAND2_X1 U7296 ( .A1(n7588), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5881) );
  OR2_X1 U7297 ( .A1(n8882), .A2(n6055), .ZN(n5885) );
  NAND2_X1 U7298 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  XNOR2_X1 U7299 ( .A(n5887), .B(n5983), .ZN(n5891) );
  NAND2_X1 U7300 ( .A1(n5890), .A2(n5891), .ZN(n8934) );
  NAND2_X1 U7301 ( .A1(n9316), .A2(n6043), .ZN(n5889) );
  OR2_X1 U7302 ( .A1(n8882), .A2(n6051), .ZN(n5888) );
  NAND2_X1 U7303 ( .A1(n5889), .A2(n5888), .ZN(n8933) );
  NAND2_X1 U7304 ( .A1(n8934), .A2(n8933), .ZN(n8938) );
  INV_X1 U7305 ( .A(n5890), .ZN(n5893) );
  INV_X1 U7306 ( .A(n5891), .ZN(n5892) );
  NAND2_X1 U7307 ( .A1(n6664), .A2(n5894), .ZN(n5896) );
  AOI22_X1 U7308 ( .A1(n6025), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9211), .B2(
        n6128), .ZN(n5895) );
  NAND2_X1 U7309 ( .A1(n9312), .A2(n6057), .ZN(n5902) );
  NAND2_X1 U7310 ( .A1(n5665), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U7311 ( .A(P1_REG3_REG_19__SCAN_IN), .B(n5910), .ZN(n9235) );
  NAND2_X1 U7312 ( .A1(n4247), .A2(n9235), .ZN(n5899) );
  NAND2_X1 U7313 ( .A1(n7588), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7314 ( .A1(n5641), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5897) );
  NAND4_X1 U7315 ( .A1(n5900), .A2(n5899), .A3(n5898), .A4(n5897), .ZN(n9224)
         );
  NAND2_X1 U7316 ( .A1(n9224), .A2(n6043), .ZN(n5901) );
  NAND2_X1 U7317 ( .A1(n5902), .A2(n5901), .ZN(n5903) );
  XNOR2_X1 U7318 ( .A(n5903), .B(n5983), .ZN(n5906) );
  AND2_X1 U7319 ( .A1(n9224), .A2(n5947), .ZN(n5904) );
  AOI21_X1 U7320 ( .B1(n9312), .B2(n6043), .A(n5904), .ZN(n5905) );
  XNOR2_X1 U7321 ( .A(n5906), .B(n5905), .ZN(n8881) );
  NAND2_X1 U7322 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  NAND2_X1 U7323 ( .A1(n6723), .A2(n5894), .ZN(n5909) );
  NAND2_X1 U7324 ( .A1(n6025), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5908) );
  NAND2_X1 U7325 ( .A1(n9306), .A2(n6057), .ZN(n5918) );
  NAND2_X1 U7326 ( .A1(n5665), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5916) );
  INV_X1 U7327 ( .A(n5910), .ZN(n5911) );
  AOI21_X1 U7328 ( .B1(P1_REG3_REG_19__SCAN_IN), .B2(n5911), .A(
        P1_REG3_REG_20__SCAN_IN), .ZN(n5912) );
  NOR2_X1 U7329 ( .A1(n5912), .A2(n5928), .ZN(n9218) );
  NAND2_X1 U7330 ( .A1(n4247), .A2(n9218), .ZN(n5915) );
  NAND2_X1 U7331 ( .A1(n7588), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5914) );
  NAND2_X1 U7332 ( .A1(n5641), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5913) );
  NAND4_X1 U7333 ( .A1(n5916), .A2(n5915), .A3(n5914), .A4(n5913), .ZN(n9242)
         );
  NAND2_X1 U7334 ( .A1(n9242), .A2(n6043), .ZN(n5917) );
  NAND2_X1 U7335 ( .A1(n5918), .A2(n5917), .ZN(n5919) );
  XNOR2_X1 U7336 ( .A(n5919), .B(n6870), .ZN(n5921) );
  AND2_X1 U7337 ( .A1(n9242), .A2(n5947), .ZN(n5920) );
  AOI21_X1 U7338 ( .B1(n9306), .B2(n6043), .A(n5920), .ZN(n5922) );
  XNOR2_X1 U7339 ( .A(n5921), .B(n5922), .ZN(n8910) );
  NAND2_X1 U7340 ( .A1(n8909), .A2(n8910), .ZN(n5925) );
  INV_X1 U7341 ( .A(n5921), .ZN(n5923) );
  NAND2_X1 U7342 ( .A1(n5923), .A2(n5922), .ZN(n5924) );
  NAND2_X2 U7343 ( .A1(n5925), .A2(n5924), .ZN(n8888) );
  NAND2_X1 U7344 ( .A1(n6752), .A2(n5894), .ZN(n5927) );
  NAND2_X1 U7345 ( .A1(n6025), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7346 ( .A1(n9303), .A2(n6057), .ZN(n5935) );
  NAND2_X1 U7347 ( .A1(n5665), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5933) );
  NOR2_X1 U7348 ( .A1(n5928), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5929) );
  NOR2_X1 U7349 ( .A1(n5940), .A2(n5929), .ZN(n9208) );
  NAND2_X1 U7350 ( .A1(n4247), .A2(n9208), .ZN(n5932) );
  NAND2_X1 U7351 ( .A1(n7588), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7352 ( .A1(n5641), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5930) );
  OR2_X1 U7353 ( .A1(n9189), .A2(n6055), .ZN(n5934) );
  NAND2_X1 U7354 ( .A1(n5935), .A2(n5934), .ZN(n5936) );
  XNOR2_X1 U7355 ( .A(n5936), .B(n6870), .ZN(n5954) );
  NOR2_X1 U7356 ( .A1(n9189), .A2(n6051), .ZN(n5937) );
  AOI21_X1 U7357 ( .B1(n9303), .B2(n6043), .A(n5937), .ZN(n5955) );
  XNOR2_X1 U7358 ( .A(n5954), .B(n5955), .ZN(n8889) );
  NAND2_X1 U7359 ( .A1(n6826), .A2(n5894), .ZN(n5939) );
  NAND2_X1 U7360 ( .A1(n6025), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5938) );
  INV_X1 U7361 ( .A(n5940), .ZN(n5942) );
  INV_X1 U7362 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7363 ( .A1(n5940), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5964) );
  INV_X1 U7364 ( .A(n5964), .ZN(n5963) );
  AOI21_X1 U7365 ( .B1(n5942), .B2(n5941), .A(n5963), .ZN(n9192) );
  NAND2_X1 U7366 ( .A1(n4247), .A2(n9192), .ZN(n5946) );
  NAND2_X1 U7367 ( .A1(n5665), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5945) );
  NAND2_X1 U7368 ( .A1(n5641), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7369 ( .A1(n7588), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5943) );
  NAND4_X1 U7370 ( .A1(n5946), .A2(n5945), .A3(n5944), .A4(n5943), .ZN(n9059)
         );
  AND2_X1 U7371 ( .A1(n9059), .A2(n5947), .ZN(n5948) );
  AOI21_X1 U7372 ( .B1(n9296), .B2(n6043), .A(n5948), .ZN(n5953) );
  AND2_X1 U7373 ( .A1(n8889), .A2(n5953), .ZN(n5949) );
  NAND2_X1 U7374 ( .A1(n9296), .A2(n6057), .ZN(n5951) );
  NAND2_X1 U7375 ( .A1(n9059), .A2(n6043), .ZN(n5950) );
  NAND2_X1 U7376 ( .A1(n5951), .A2(n5950), .ZN(n5952) );
  XNOR2_X1 U7377 ( .A(n5952), .B(n6870), .ZN(n8922) );
  INV_X1 U7378 ( .A(n5953), .ZN(n5959) );
  INV_X1 U7379 ( .A(n5954), .ZN(n5956) );
  NAND2_X1 U7380 ( .A1(n5956), .A2(n5955), .ZN(n5958) );
  OR2_X1 U7381 ( .A1(n5959), .A2(n5958), .ZN(n8918) );
  AND2_X1 U7382 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  NAND2_X1 U7383 ( .A1(n7010), .A2(n5894), .ZN(n5962) );
  NAND2_X1 U7384 ( .A1(n6025), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5961) );
  INV_X1 U7385 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7386 ( .A1(n5963), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5975) );
  INV_X1 U7387 ( .A(n5975), .ZN(n5977) );
  AOI21_X1 U7388 ( .B1(n5965), .B2(n5964), .A(n5977), .ZN(n9179) );
  NAND2_X1 U7389 ( .A1(n4247), .A2(n9179), .ZN(n5969) );
  NAND2_X1 U7390 ( .A1(n5665), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7391 ( .A1(n7588), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7392 ( .A1(n5641), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5966) );
  OAI22_X1 U7393 ( .A1(n9182), .A2(n6018), .B1(n9190), .B2(n6055), .ZN(n5970)
         );
  NOR2_X1 U7394 ( .A1(n9190), .A2(n6051), .ZN(n5971) );
  AOI21_X1 U7395 ( .B1(n9292), .B2(n6043), .A(n5971), .ZN(n8873) );
  NAND2_X1 U7396 ( .A1(n8872), .A2(n8873), .ZN(n5972) );
  NAND3_X1 U7397 ( .A1(n8921), .A2(n4307), .A3(n8917), .ZN(n8871) );
  NAND2_X1 U7398 ( .A1(n7062), .A2(n5894), .ZN(n5974) );
  NAND2_X1 U7399 ( .A1(n6025), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5973) );
  INV_X1 U7400 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5976) );
  NAND2_X1 U7401 ( .A1(n5976), .A2(n5975), .ZN(n5978) );
  NAND2_X1 U7402 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n5977), .ZN(n5994) );
  AND2_X1 U7403 ( .A1(n5978), .A2(n5994), .ZN(n9163) );
  NAND2_X1 U7404 ( .A1(n4247), .A2(n9163), .ZN(n5982) );
  NAND2_X1 U7405 ( .A1(n5665), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7406 ( .A1(n5641), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7407 ( .A1(n7588), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5979) );
  OAI22_X1 U7408 ( .A1(n9166), .A2(n6018), .B1(n9175), .B2(n6055), .ZN(n5984)
         );
  XNOR2_X1 U7409 ( .A(n5984), .B(n5983), .ZN(n5985) );
  OAI22_X1 U7410 ( .A1(n9166), .A2(n6055), .B1(n9175), .B2(n6051), .ZN(n5986)
         );
  XNOR2_X1 U7411 ( .A(n5985), .B(n5986), .ZN(n8903) );
  INV_X1 U7412 ( .A(n5985), .ZN(n5987) );
  OR2_X1 U7413 ( .A1(n5987), .A2(n5986), .ZN(n5988) );
  NAND2_X1 U7414 ( .A1(n7189), .A2(n5894), .ZN(n5991) );
  NAND2_X1 U7415 ( .A1(n6025), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7416 ( .A1(n9279), .A2(n6057), .ZN(n6001) );
  INV_X1 U7417 ( .A(n5994), .ZN(n5992) );
  NAND2_X1 U7418 ( .A1(n5992), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6012) );
  INV_X1 U7419 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7420 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  AND2_X1 U7421 ( .A1(n6012), .A2(n5995), .ZN(n9145) );
  NAND2_X1 U7422 ( .A1(n4247), .A2(n9145), .ZN(n5999) );
  NAND2_X1 U7423 ( .A1(n5665), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7424 ( .A1(n5641), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7425 ( .A1(n7588), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5996) );
  OR2_X1 U7426 ( .A1(n9161), .A2(n6055), .ZN(n6000) );
  NAND2_X1 U7427 ( .A1(n6001), .A2(n6000), .ZN(n6002) );
  XNOR2_X1 U7428 ( .A(n6002), .B(n6870), .ZN(n6004) );
  NOR2_X1 U7429 ( .A1(n9161), .A2(n6051), .ZN(n6003) );
  AOI21_X1 U7430 ( .B1(n9279), .B2(n6043), .A(n6003), .ZN(n6005) );
  XNOR2_X1 U7431 ( .A(n6004), .B(n6005), .ZN(n8896) );
  NAND2_X1 U7432 ( .A1(n8895), .A2(n8896), .ZN(n6008) );
  INV_X1 U7433 ( .A(n6004), .ZN(n6006) );
  NAND2_X1 U7434 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  NAND2_X1 U7435 ( .A1(n7221), .A2(n5894), .ZN(n6010) );
  NAND2_X1 U7436 ( .A1(n6025), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6009) );
  INV_X1 U7437 ( .A(n6012), .ZN(n6011) );
  NAND2_X1 U7438 ( .A1(n6011), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6030) );
  INV_X1 U7439 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8953) );
  NAND2_X1 U7440 ( .A1(n6012), .A2(n8953), .ZN(n6013) );
  AND2_X1 U7441 ( .A1(n6030), .A2(n6013), .ZN(n9129) );
  NAND2_X1 U7442 ( .A1(n4247), .A2(n9129), .ZN(n6017) );
  NAND2_X1 U7443 ( .A1(n5665), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7444 ( .A1(n5641), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7445 ( .A1(n7588), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6014) );
  OAI22_X1 U7446 ( .A1(n9131), .A2(n6018), .B1(n9121), .B2(n6055), .ZN(n6019)
         );
  XNOR2_X1 U7447 ( .A(n6019), .B(n6870), .ZN(n6023) );
  OR2_X1 U7448 ( .A1(n9131), .A2(n6055), .ZN(n6021) );
  OR2_X1 U7449 ( .A1(n9121), .A2(n6051), .ZN(n6020) );
  NAND2_X1 U7450 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  XNOR2_X1 U7451 ( .A(n6023), .B(n6022), .ZN(n8948) );
  NAND2_X1 U7452 ( .A1(n6023), .A2(n6022), .ZN(n6024) );
  NAND2_X1 U7453 ( .A1(n6025), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7454 ( .A1(n9269), .A2(n6057), .ZN(n6037) );
  INV_X1 U7455 ( .A(n6030), .ZN(n6028) );
  NAND2_X1 U7456 ( .A1(n6028), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6045) );
  INV_X1 U7457 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U7458 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  AND2_X1 U7459 ( .A1(n6045), .A2(n6031), .ZN(n9114) );
  NAND2_X1 U7460 ( .A1(n4247), .A2(n9114), .ZN(n6035) );
  NAND2_X1 U7461 ( .A1(n5665), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7462 ( .A1(n7588), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6033) );
  NAND2_X1 U7463 ( .A1(n5641), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6032) );
  OR2_X1 U7464 ( .A1(n9135), .A2(n6055), .ZN(n6036) );
  NAND2_X1 U7465 ( .A1(n6037), .A2(n6036), .ZN(n6038) );
  XNOR2_X1 U7466 ( .A(n6038), .B(n6870), .ZN(n6083) );
  NAND2_X1 U7467 ( .A1(n9269), .A2(n6043), .ZN(n6040) );
  OR2_X1 U7468 ( .A1(n9135), .A2(n6051), .ZN(n6039) );
  NAND2_X1 U7469 ( .A1(n6040), .A2(n6039), .ZN(n6084) );
  NAND2_X1 U7470 ( .A1(n7281), .A2(n5894), .ZN(n6042) );
  NAND2_X1 U7471 ( .A1(n6025), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7472 ( .A1(n9264), .A2(n6043), .ZN(n6053) );
  NAND2_X1 U7473 ( .A1(n5665), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6050) );
  INV_X1 U7474 ( .A(n6045), .ZN(n6044) );
  NAND2_X1 U7475 ( .A1(n6044), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6107) );
  INV_X1 U7476 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7477 ( .A1(n6045), .A2(n6115), .ZN(n6046) );
  AND2_X1 U7478 ( .A1(n6107), .A2(n6046), .ZN(n9098) );
  NAND2_X1 U7479 ( .A1(n4247), .A2(n9098), .ZN(n6049) );
  NAND2_X1 U7480 ( .A1(n7588), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7481 ( .A1(n5641), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6047) );
  OR2_X1 U7482 ( .A1(n9120), .A2(n6051), .ZN(n6052) );
  NAND2_X1 U7483 ( .A1(n6053), .A2(n6052), .ZN(n6054) );
  XNOR2_X1 U7484 ( .A(n6054), .B(n6870), .ZN(n6059) );
  NOR2_X1 U7485 ( .A1(n9120), .A2(n6055), .ZN(n6056) );
  AOI21_X1 U7486 ( .B1(n9264), .B2(n6057), .A(n6056), .ZN(n6058) );
  XNOR2_X1 U7487 ( .A(n6059), .B(n6058), .ZN(n6088) );
  INV_X1 U7488 ( .A(n6088), .ZN(n6119) );
  INV_X1 U7489 ( .A(n7875), .ZN(n6827) );
  INV_X1 U7490 ( .A(n6060), .ZN(n7823) );
  NAND2_X1 U7491 ( .A1(n6827), .A2(n7823), .ZN(n6552) );
  INV_X1 U7492 ( .A(n6552), .ZN(n6062) );
  NAND2_X1 U7493 ( .A1(n7875), .A2(n6060), .ZN(n7716) );
  NAND2_X1 U7494 ( .A1(n6063), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6064) );
  XNOR2_X1 U7495 ( .A(n6064), .B(n4715), .ZN(n6126) );
  AND2_X1 U7496 ( .A1(n6126), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6065) );
  AND2_X1 U7497 ( .A1(n6092), .A2(n6065), .ZN(n9360) );
  NAND2_X1 U7498 ( .A1(n7716), .A2(n9360), .ZN(n6082) );
  INV_X1 U7499 ( .A(n6070), .ZN(n7190) );
  NAND3_X1 U7500 ( .A1(n7190), .A2(P1_B_REG_SCAN_IN), .A3(n7067), .ZN(n6069)
         );
  INV_X1 U7501 ( .A(P1_B_REG_SCAN_IN), .ZN(n6066) );
  NAND2_X1 U7502 ( .A1(n6067), .A2(n6066), .ZN(n6068) );
  AND3_X1 U7503 ( .A1(n6080), .A2(n6069), .A3(n6068), .ZN(n6155) );
  INV_X1 U7504 ( .A(n6155), .ZN(n6222) );
  OAI22_X1 U7505 ( .A1(n6222), .A2(P1_D_REG_1__SCAN_IN), .B1(n6080), .B2(n6070), .ZN(n6555) );
  INV_X1 U7506 ( .A(n6555), .ZN(n9361) );
  NOR4_X1 U7507 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6074) );
  NOR4_X1 U7508 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6073) );
  NOR4_X1 U7509 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6072) );
  NOR4_X1 U7510 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6071) );
  NAND4_X1 U7511 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n6079)
         );
  NOR2_X1 U7512 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n9758) );
  NOR4_X1 U7513 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6077) );
  NOR4_X1 U7514 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6076) );
  NOR4_X1 U7515 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6075) );
  NAND4_X1 U7516 ( .A1(n9758), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n6078)
         );
  NOR2_X1 U7517 ( .A1(n6079), .A2(n6078), .ZN(n6153) );
  NAND2_X1 U7518 ( .A1(n6153), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6081) );
  INV_X1 U7519 ( .A(n6080), .ZN(n7223) );
  AND2_X1 U7520 ( .A1(n7223), .A2(n7067), .ZN(n6152) );
  AOI21_X1 U7521 ( .B1(n6155), .B2(n6081), .A(n6152), .ZN(n6556) );
  NAND2_X1 U7522 ( .A1(n9361), .A2(n6556), .ZN(n6112) );
  OR3_X1 U7523 ( .A1(n9520), .A2(n6082), .A3(n6112), .ZN(n8947) );
  INV_X1 U7524 ( .A(n8947), .ZN(n8926) );
  INV_X1 U7525 ( .A(n6083), .ZN(n6086) );
  INV_X1 U7526 ( .A(n6084), .ZN(n6085) );
  NAND2_X1 U7527 ( .A1(n6086), .A2(n6085), .ZN(n8861) );
  NAND3_X1 U7528 ( .A1(n6119), .A2(n8926), .A3(n8861), .ZN(n6087) );
  OR2_X1 U7529 ( .A1(n6090), .A2(n6087), .ZN(n6124) );
  AND2_X1 U7530 ( .A1(n6088), .A2(n8926), .ZN(n6089) );
  NAND2_X1 U7531 ( .A1(n6090), .A2(n6089), .ZN(n6123) );
  OR2_X1 U7532 ( .A1(n7716), .A2(n6091), .ZN(n6094) );
  AND2_X1 U7533 ( .A1(n6092), .A2(n6126), .ZN(n6093) );
  NAND2_X1 U7534 ( .A1(n6094), .A2(n6093), .ZN(n6158) );
  OR2_X1 U7535 ( .A1(n6158), .A2(P1_U3084), .ZN(n6096) );
  NAND2_X2 U7536 ( .A1(n6827), .A2(n9211), .ZN(n7704) );
  INV_X1 U7537 ( .A(n7777), .ZN(n7869) );
  NOR2_X1 U7538 ( .A1(n9335), .A2(n6060), .ZN(n6095) );
  INV_X1 U7539 ( .A(n6112), .ZN(n6106) );
  NOR2_X1 U7540 ( .A1(n6558), .A2(n6106), .ZN(n6099) );
  INV_X1 U7541 ( .A(n6099), .ZN(n6098) );
  INV_X1 U7542 ( .A(n6096), .ZN(n6097) );
  AND2_X1 U7543 ( .A1(n6098), .A2(n6097), .ZN(n6609) );
  AOI21_X1 U7544 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6158), .A(n6099), .ZN(n7541) );
  INV_X1 U7545 ( .A(n9098), .ZN(n6118) );
  OR3_X1 U7546 ( .A1(n6827), .A2(n9211), .A3(n6160), .ZN(n6871) );
  INV_X1 U7547 ( .A(n9360), .ZN(n6100) );
  NOR2_X1 U7548 ( .A1(n6871), .A2(n6100), .ZN(n6114) );
  INV_X1 U7549 ( .A(n6114), .ZN(n6105) );
  NAND2_X1 U7550 ( .A1(n6101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7551 ( .A1(n6257), .A2(n6102), .ZN(n6104) );
  XNOR2_X1 U7552 ( .A(n6104), .B(n6103), .ZN(n6495) );
  INV_X1 U7553 ( .A(n6495), .ZN(n6258) );
  NOR2_X1 U7554 ( .A1(n6105), .A2(n6258), .ZN(n7873) );
  AND2_X1 U7555 ( .A1(n7873), .A2(n6106), .ZN(n8940) );
  INV_X1 U7556 ( .A(n9135), .ZN(n9065) );
  INV_X1 U7557 ( .A(n6107), .ZN(n9089) );
  NAND2_X1 U7558 ( .A1(n4247), .A2(n9089), .ZN(n6111) );
  NAND2_X1 U7559 ( .A1(n5665), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6110) );
  NAND2_X1 U7560 ( .A1(n5641), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7561 ( .A1(n7588), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6108) );
  NOR2_X1 U7562 ( .A1(n6112), .A2(n6495), .ZN(n6113) );
  NAND2_X1 U7563 ( .A1(n6114), .A2(n6113), .ZN(n8954) );
  OAI22_X1 U7564 ( .A1(n9105), .A2(n8954), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6115), .ZN(n6116) );
  AOI21_X1 U7565 ( .B1(n8940), .B2(n9065), .A(n6116), .ZN(n6117) );
  OAI21_X1 U7566 ( .B1(n7541), .B2(n6118), .A(n6117), .ZN(n6121) );
  NOR3_X1 U7567 ( .A1(n6119), .A2(n8947), .A3(n8861), .ZN(n6120) );
  AOI211_X1 U7568 ( .C1(n8914), .C2(n9264), .A(n6121), .B(n6120), .ZN(n6122)
         );
  NAND3_X1 U7569 ( .A1(n6124), .A2(n6123), .A3(n6122), .ZN(P1_U3218) );
  NAND2_X1 U7570 ( .A1(n6125), .A2(n6126), .ZN(n6255) );
  OR2_X1 U7571 ( .A1(n6255), .A2(P1_U3084), .ZN(n8961) );
  INV_X1 U7572 ( .A(n8961), .ZN(P1_U4006) );
  INV_X1 U7573 ( .A(n6126), .ZN(n7011) );
  OR2_X1 U7574 ( .A1(n7716), .A2(n7011), .ZN(n6127) );
  NAND2_X1 U7575 ( .A1(n6127), .A2(n6255), .ZN(n6265) );
  OR2_X1 U7576 ( .A1(n6265), .A2(n6128), .ZN(n6129) );
  NAND2_X1 U7577 ( .A1(n6129), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  OR2_X1 U7578 ( .A1(n6175), .A2(n9624), .ZN(n8425) );
  INV_X2 U7579 ( .A(n8425), .ZN(P2_U3966) );
  NAND2_X1 U7580 ( .A1(n7875), .A2(n9211), .ZN(n6130) );
  NAND2_X1 U7581 ( .A1(n6060), .A2(n7869), .ZN(n7714) );
  AND2_X1 U7582 ( .A1(n6130), .A2(n7714), .ZN(n9203) );
  NOR2_X1 U7583 ( .A1(n6575), .A2(n6570), .ZN(n6573) );
  INV_X1 U7584 ( .A(n8976), .ZN(n7832) );
  NAND2_X1 U7585 ( .A1(n7832), .A2(n7831), .ZN(n6132) );
  NAND2_X1 U7586 ( .A1(n6133), .A2(n6941), .ZN(n7834) );
  INV_X1 U7587 ( .A(n6133), .ZN(n8975) );
  NAND2_X1 U7588 ( .A1(n8975), .A2(n6937), .ZN(n7838) );
  NAND2_X1 U7589 ( .A1(n8974), .A2(n6991), .ZN(n7739) );
  NAND2_X1 U7590 ( .A1(n6832), .A2(n6705), .ZN(n7836) );
  NAND2_X1 U7591 ( .A1(n7747), .A2(n7795), .ZN(n6134) );
  INV_X1 U7592 ( .A(n6950), .ZN(n8973) );
  NAND2_X1 U7593 ( .A1(n8973), .A2(n9511), .ZN(n7742) );
  NAND2_X1 U7594 ( .A1(n6950), .A2(n6840), .ZN(n7596) );
  NAND2_X1 U7595 ( .A1(n7599), .A2(n7596), .ZN(n6948) );
  NAND2_X1 U7596 ( .A1(n6831), .A2(n9519), .ZN(n7741) );
  INV_X1 U7597 ( .A(n6831), .ZN(n6136) );
  NAND2_X1 U7598 ( .A1(n6136), .A2(n6135), .ZN(n7604) );
  NAND2_X1 U7599 ( .A1(n6948), .A2(n7797), .ZN(n6947) );
  NAND2_X1 U7600 ( .A1(n6947), .A2(n7741), .ZN(n6138) );
  NAND2_X1 U7601 ( .A1(n6949), .A2(n6163), .ZN(n7610) );
  INV_X1 U7602 ( .A(n6949), .ZN(n8972) );
  INV_X1 U7603 ( .A(n7801), .ZN(n6137) );
  XNOR2_X1 U7604 ( .A(n6138), .B(n6137), .ZN(n6151) );
  INV_X1 U7605 ( .A(n6574), .ZN(n7799) );
  AND2_X1 U7606 ( .A1(n6575), .A2(n6795), .ZN(n6569) );
  NAND2_X1 U7607 ( .A1(n8976), .A2(n7831), .ZN(n6139) );
  NAND2_X1 U7608 ( .A1(n6133), .A2(n6937), .ZN(n6140) );
  NAND2_X1 U7609 ( .A1(n6698), .A2(n6699), .ZN(n6697) );
  NAND2_X1 U7610 ( .A1(n6832), .A2(n6991), .ZN(n6141) );
  NAND2_X1 U7611 ( .A1(n6697), .A2(n6141), .ZN(n6830) );
  NAND2_X1 U7612 ( .A1(n7596), .A2(n7742), .ZN(n7792) );
  NAND2_X1 U7613 ( .A1(n6830), .A2(n7792), .ZN(n6829) );
  NAND2_X1 U7614 ( .A1(n6950), .A2(n9511), .ZN(n6142) );
  OR2_X1 U7615 ( .A1(n6998), .A2(n7797), .ZN(n6954) );
  NAND2_X1 U7616 ( .A1(n6136), .A2(n9519), .ZN(n6756) );
  NAND2_X1 U7617 ( .A1(n6954), .A2(n6756), .ZN(n6143) );
  OR2_X1 U7618 ( .A1(n6143), .A2(n7801), .ZN(n6145) );
  NAND2_X1 U7619 ( .A1(n6143), .A2(n7801), .ZN(n6144) );
  NAND2_X1 U7620 ( .A1(n6145), .A2(n6144), .ZN(n9531) );
  XNOR2_X1 U7621 ( .A(n7875), .B(n6160), .ZN(n6146) );
  NAND2_X1 U7622 ( .A1(n6146), .A2(n9033), .ZN(n9382) );
  INV_X1 U7623 ( .A(n9382), .ZN(n6834) );
  NAND2_X1 U7624 ( .A1(n9531), .A2(n6834), .ZN(n6150) );
  INV_X1 U7625 ( .A(n7716), .ZN(n6147) );
  AND2_X1 U7626 ( .A1(n6147), .A2(n6495), .ZN(n9409) );
  INV_X1 U7627 ( .A(n9409), .ZN(n9378) );
  OAI22_X1 U7628 ( .A1(n6831), .A2(n9378), .B1(n6906), .B2(n9376), .ZN(n6148)
         );
  INV_X1 U7629 ( .A(n6148), .ZN(n6149) );
  OAI211_X1 U7630 ( .C1(n9203), .C2(n6151), .A(n6150), .B(n6149), .ZN(n9529)
         );
  INV_X1 U7631 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9787) );
  NAND2_X1 U7632 ( .A1(n6155), .A2(n9787), .ZN(n6156) );
  INV_X1 U7633 ( .A(n6152), .ZN(n6223) );
  INV_X1 U7634 ( .A(n6153), .ZN(n6154) );
  AOI22_X1 U7635 ( .A1(n6156), .A2(n6223), .B1(n6155), .B2(n6154), .ZN(n6547)
         );
  NAND3_X1 U7636 ( .A1(n6547), .A2(n9361), .A3(P1_STATE_REG_SCAN_IN), .ZN(
        n6157) );
  OR2_X1 U7637 ( .A1(n6158), .A2(n6157), .ZN(n6165) );
  NAND2_X1 U7638 ( .A1(n7823), .A2(n9360), .ZN(n6159) );
  INV_X2 U7639 ( .A(n7027), .ZN(n9430) );
  MUX2_X1 U7640 ( .A(n9529), .B(P1_REG2_REG_6__SCAN_IN), .S(n9430), .Z(n6171)
         );
  INV_X1 U7641 ( .A(n9531), .ZN(n6162) );
  OR2_X1 U7642 ( .A1(n6160), .A2(n9033), .ZN(n6161) );
  OR2_X1 U7643 ( .A1(n9430), .A2(n6161), .ZN(n7491) );
  NOR2_X1 U7644 ( .A1(n6162), .A2(n7491), .ZN(n6170) );
  NOR2_X1 U7645 ( .A1(n7831), .A2(n6795), .ZN(n6938) );
  NAND2_X1 U7646 ( .A1(n6940), .A2(n6991), .ZN(n6837) );
  NOR2_X1 U7647 ( .A1(n6956), .A2(n6163), .ZN(n6766) );
  INV_X1 U7648 ( .A(n6766), .ZN(n6767) );
  NAND2_X1 U7649 ( .A1(n6956), .A2(n6163), .ZN(n6164) );
  NAND2_X1 U7650 ( .A1(n6767), .A2(n6164), .ZN(n9528) );
  NOR2_X1 U7651 ( .A1(n6165), .A2(n9211), .ZN(n9426) );
  INV_X1 U7652 ( .A(n9426), .ZN(n6961) );
  INV_X1 U7653 ( .A(n9542), .ZN(n9423) );
  NAND2_X1 U7654 ( .A1(n9426), .A2(n9423), .ZN(n9088) );
  NOR2_X1 U7655 ( .A1(n9528), .A2(n9088), .ZN(n6169) );
  OR2_X1 U7656 ( .A1(n6552), .A2(n7777), .ZN(n6166) );
  OAI22_X1 U7657 ( .A1(n9237), .A2(n9527), .B1(n6167), .B2(n9209), .ZN(n6168)
         );
  OR4_X1 U7658 ( .A1(n6171), .A2(n6170), .A3(n6169), .A4(n6168), .ZN(P1_U3285)
         );
  INV_X1 U7659 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6409) );
  XNOR2_X1 U7660 ( .A(n6207), .B(n6409), .ZN(n8085) );
  NAND2_X1 U7661 ( .A1(n8859), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8084) );
  NOR2_X1 U7662 ( .A1(n8085), .A2(n8084), .ZN(n6172) );
  AOI21_X1 U7663 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n8093), .A(n6172), .ZN(
        n6182) );
  INV_X1 U7664 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6173) );
  MUX2_X1 U7665 ( .A(n6173), .B(P2_REG2_REG_2__SCAN_IN), .S(n7310), .Z(n6181)
         );
  NOR2_X1 U7666 ( .A1(n6182), .A2(n6181), .ZN(n8011) );
  OR2_X1 U7667 ( .A1(n6174), .A2(P2_U3152), .ZN(n8328) );
  INV_X1 U7668 ( .A(n6175), .ZN(n6176) );
  NAND2_X1 U7669 ( .A1(n6176), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6177) );
  OAI211_X1 U7670 ( .C1(n9589), .C2(n6178), .A(n8328), .B(n6177), .ZN(n6179)
         );
  AND2_X1 U7671 ( .A1(n6179), .A2(n4878), .ZN(n6183) );
  INV_X1 U7672 ( .A(n6183), .ZN(n6180) );
  NAND2_X1 U7673 ( .A1(n6180), .A2(n8425), .ZN(n6186) );
  INV_X1 U7674 ( .A(n7269), .ZN(n8463) );
  NAND2_X1 U7675 ( .A1(n6186), .A2(n8463), .ZN(n6391) );
  OR2_X1 U7676 ( .A1(n6391), .A2(n5492), .ZN(n8450) );
  AOI211_X1 U7677 ( .C1(n6182), .C2(n6181), .A(n8011), .B(n8450), .ZN(n6194)
         );
  XNOR2_X1 U7678 ( .A(n8093), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n8089) );
  NAND2_X1 U7679 ( .A1(n8859), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8090) );
  NOR2_X1 U7680 ( .A1(n8089), .A2(n8090), .ZN(n8088) );
  AOI21_X1 U7681 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n8093), .A(n8088), .ZN(
        n6185) );
  XNOR2_X1 U7682 ( .A(n7310), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6184) );
  NOR2_X1 U7683 ( .A1(n6185), .A2(n6184), .ZN(n7309) );
  AND2_X1 U7684 ( .A1(n6183), .A2(n7269), .ZN(n8453) );
  INV_X1 U7685 ( .A(n8453), .ZN(n8087) );
  AOI211_X1 U7686 ( .C1(n6185), .C2(n6184), .A(n7309), .B(n8087), .ZN(n6193)
         );
  NAND2_X1 U7687 ( .A1(n6186), .A2(n5492), .ZN(n8448) );
  INV_X1 U7688 ( .A(n7310), .ZN(n7337) );
  NOR2_X1 U7689 ( .A1(n8448), .A2(n7337), .ZN(n6192) );
  OAI21_X1 U7690 ( .B1(n9589), .B2(n6187), .A(n4878), .ZN(n6189) );
  NAND2_X1 U7691 ( .A1(n9589), .A2(n8328), .ZN(n6188) );
  NAND2_X1 U7692 ( .A1(n6189), .A2(n6188), .ZN(n8460) );
  INV_X1 U7693 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6190) );
  INV_X1 U7694 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6448) );
  OAI22_X1 U7695 ( .A1(n8460), .A2(n6190), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6448), .ZN(n6191) );
  OR4_X1 U7696 ( .A1(n6194), .A2(n6193), .A3(n6192), .A4(n6191), .ZN(P2_U3247)
         );
  AOI22_X1 U7697 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n9366), .B1(n6509), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6195) );
  OAI21_X1 U7698 ( .B1(n6197), .B2(n8334), .A(n6195), .ZN(P1_U3349) );
  NOR2_X1 U7699 ( .A1(n6196), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8851) );
  NAND2_X1 U7700 ( .A1(n6196), .A2(P2_U3152), .ZN(n8858) );
  INV_X1 U7701 ( .A(n7340), .ZN(n7999) );
  OAI222_X1 U7702 ( .A1(n8856), .A2(n6198), .B1(n8858), .B2(n6197), .C1(
        P2_U3152), .C2(n7999), .ZN(P2_U3354) );
  OAI222_X1 U7703 ( .A1(n8856), .A2(n9751), .B1(n8858), .B2(n6203), .C1(
        P2_U3152), .C2(n7337), .ZN(P2_U3356) );
  INV_X1 U7704 ( .A(n6199), .ZN(n6206) );
  AOI22_X1 U7705 ( .A1(n8080), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n8851), .ZN(n6200) );
  OAI21_X1 U7706 ( .B1(n6206), .B2(n8858), .A(n6200), .ZN(P2_U3353) );
  INV_X1 U7707 ( .A(n9366), .ZN(n8333) );
  INV_X1 U7708 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6201) );
  INV_X1 U7709 ( .A(n6283), .ZN(n6304) );
  OAI222_X1 U7710 ( .A1(n8333), .A2(n6201), .B1(n8334), .B2(n6208), .C1(
        P1_U3084), .C2(n6304), .ZN(P1_U3352) );
  INV_X1 U7711 ( .A(n6340), .ZN(n6285) );
  OAI222_X1 U7712 ( .A1(n8333), .A2(n6202), .B1(n8334), .B2(n6210), .C1(
        P1_U3084), .C2(n6285), .ZN(P1_U3350) );
  INV_X1 U7713 ( .A(n6284), .ZN(n6520) );
  OAI222_X1 U7714 ( .A1(n8333), .A2(n6204), .B1(n8334), .B2(n6203), .C1(
        P1_U3084), .C2(n6520), .ZN(P1_U3351) );
  INV_X1 U7715 ( .A(n9458), .ZN(n6205) );
  OAI222_X1 U7716 ( .A1(n8333), .A2(n9867), .B1(n8334), .B2(n6206), .C1(
        P1_U3084), .C2(n6205), .ZN(P1_U3348) );
  INV_X1 U7717 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6209) );
  CLKBUF_X1 U7718 ( .A(n8858), .Z(n8098) );
  OAI222_X1 U7719 ( .A1(n8856), .A2(n6209), .B1(n8098), .B2(n6208), .C1(
        P2_U3152), .C2(n6207), .ZN(P2_U3357) );
  INV_X1 U7720 ( .A(n8006), .ZN(n8014) );
  OAI222_X1 U7721 ( .A1(n8856), .A2(n6211), .B1(n8098), .B2(n6210), .C1(
        P2_U3152), .C2(n8014), .ZN(P2_U3355) );
  INV_X1 U7722 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6213) );
  INV_X1 U7723 ( .A(n6212), .ZN(n6214) );
  OAI222_X1 U7724 ( .A1(n8856), .A2(n6213), .B1(n8858), .B2(n6214), .C1(
        P2_U3152), .C2(n7985), .ZN(P2_U3352) );
  INV_X1 U7725 ( .A(n9470), .ZN(n6276) );
  OAI222_X1 U7726 ( .A1(n8333), .A2(n6215), .B1(n8334), .B2(n6214), .C1(
        P1_U3084), .C2(n6276), .ZN(P1_U3347) );
  INV_X1 U7727 ( .A(n6216), .ZN(n6218) );
  AOI22_X1 U7728 ( .A1(n6321), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9366), .ZN(n6217) );
  OAI21_X1 U7729 ( .B1(n6218), .B2(n8334), .A(n6217), .ZN(P1_U3346) );
  INV_X1 U7730 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6219) );
  INV_X1 U7731 ( .A(n7334), .ZN(n7974) );
  OAI222_X1 U7732 ( .A1(n8856), .A2(n6219), .B1(n8098), .B2(n6218), .C1(
        P2_U3152), .C2(n7974), .ZN(P2_U3351) );
  INV_X1 U7733 ( .A(n6220), .ZN(n6225) );
  AOI22_X1 U7734 ( .A1(n9484), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9366), .ZN(n6221) );
  OAI21_X1 U7735 ( .B1(n6225), .B2(n8334), .A(n6221), .ZN(P1_U3345) );
  AND2_X1 U7736 ( .A1(n6222), .A2(n9360), .ZN(n9503) );
  NAND2_X1 U7737 ( .A1(n9503), .A2(n6223), .ZN(n6224) );
  OAI21_X1 U7738 ( .B1(n9503), .B2(n9787), .A(n6224), .ZN(P1_U3440) );
  INV_X1 U7739 ( .A(n7331), .ZN(n7962) );
  OAI222_X1 U7740 ( .A1(n8856), .A2(n9805), .B1(n8098), .B2(n6225), .C1(
        P2_U3152), .C2(n7962), .ZN(P2_U3350) );
  INV_X1 U7741 ( .A(n6226), .ZN(n6229) );
  OAI222_X1 U7742 ( .A1(n8333), .A2(n6228), .B1(n8334), .B2(n6229), .C1(n6227), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U7743 ( .A(n7328), .ZN(n7950) );
  OAI222_X1 U7744 ( .A1(n8856), .A2(n6230), .B1(n8858), .B2(n6229), .C1(n7950), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  NAND2_X1 U7745 ( .A1(n4900), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U7746 ( .A1(n4265), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7747 ( .A1(n5314), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6231) );
  AND3_X1 U7748 ( .A1(n6233), .A2(n6232), .A3(n6231), .ZN(n8494) );
  NAND2_X1 U7749 ( .A1(n8425), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6234) );
  OAI21_X1 U7750 ( .B1(n8425), .B2(n8494), .A(n6234), .ZN(P2_U3582) );
  INV_X1 U7751 ( .A(n6235), .ZN(n6237) );
  INV_X1 U7752 ( .A(n6589), .ZN(n6323) );
  OAI222_X1 U7753 ( .A1(n8333), .A2(n6236), .B1(n8334), .B2(n6237), .C1(n6323), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U7754 ( .A(n7325), .ZN(n7938) );
  OAI222_X1 U7755 ( .A1(n8856), .A2(n6238), .B1(n8098), .B2(n6237), .C1(n7938), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U7756 ( .A(n6239), .ZN(n6241) );
  INV_X1 U7757 ( .A(n6590), .ZN(n8982) );
  OAI222_X1 U7758 ( .A1(n8333), .A2(n6240), .B1(n8334), .B2(n6241), .C1(n8982), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  INV_X1 U7759 ( .A(n7347), .ZN(n8067) );
  OAI222_X1 U7760 ( .A1(n8856), .A2(n6242), .B1(n8098), .B2(n6241), .C1(n8067), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U7761 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9834) );
  NAND2_X1 U7762 ( .A1(n6575), .A2(P1_U4006), .ZN(n6243) );
  OAI21_X1 U7763 ( .B1(P1_U4006), .B2(n9834), .A(n6243), .ZN(P1_U3555) );
  INV_X1 U7764 ( .A(n8460), .ZN(n8079) );
  NOR2_X1 U7765 ( .A1(n8079), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7766 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7767 ( .A1(n6244), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7768 ( .A1(n4900), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7769 ( .A1(n5314), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6245) );
  AND3_X1 U7770 ( .A1(n6247), .A2(n6246), .A3(n6245), .ZN(n8465) );
  INV_X1 U7771 ( .A(n8465), .ZN(n6248) );
  NAND2_X1 U7772 ( .A1(n6248), .A2(P2_U3966), .ZN(n6249) );
  OAI21_X1 U7773 ( .B1(P2_U3966), .B2(n6250), .A(n6249), .ZN(P2_U3583) );
  INV_X1 U7774 ( .A(n6251), .ZN(n6253) );
  OAI222_X1 U7775 ( .A1(n8333), .A2(n6252), .B1(n8334), .B2(n6253), .C1(
        P1_U3084), .C2(n6586), .ZN(P1_U3341) );
  INV_X1 U7776 ( .A(n7917), .ZN(n7924) );
  OAI222_X1 U7777 ( .A1(n8856), .A2(n6254), .B1(n8098), .B2(n6253), .C1(
        P2_U3152), .C2(n7924), .ZN(P2_U3346) );
  INV_X1 U7778 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6264) );
  INV_X1 U7779 ( .A(n6255), .ZN(n6256) );
  OR2_X1 U7780 ( .A1(P1_U3083), .A2(n6256), .ZN(n9038) );
  INV_X1 U7781 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6561) );
  XNOR2_X1 U7782 ( .A(n6257), .B(P1_IR_REG_27__SCAN_IN), .ZN(n9039) );
  INV_X1 U7783 ( .A(n9039), .ZN(n6497) );
  INV_X1 U7784 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6259) );
  AOI21_X1 U7785 ( .B1(n9039), .B2(n6259), .A(n6258), .ZN(n6500) );
  XNOR2_X1 U7786 ( .A(n6500), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6260) );
  AOI211_X1 U7787 ( .C1(n6561), .C2(n6497), .A(P1_U3084), .B(n6260), .ZN(n6261) );
  AOI22_X1 U7788 ( .A1(n6261), .A2(P1_U3083), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3084), .ZN(n6263) );
  NAND2_X1 U7789 ( .A1(n6495), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7283) );
  OR2_X1 U7790 ( .A1(n6265), .A2(n7283), .ZN(n6280) );
  OR2_X1 U7791 ( .A1(n6280), .A2(n9039), .ZN(n9476) );
  INV_X1 U7792 ( .A(n9476), .ZN(n9497) );
  NAND3_X1 U7793 ( .A1(n9497), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6561), .ZN(
        n6262) );
  OAI211_X1 U7794 ( .C1(n6264), .C2(n9038), .A(n6263), .B(n6262), .ZN(P1_U3241) );
  INV_X1 U7795 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U7796 ( .A1(n9039), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7242) );
  OR2_X1 U7797 ( .A1(n6265), .A2(n7242), .ZN(n9023) );
  OR2_X1 U7798 ( .A1(n9023), .A2(n6495), .ZN(n9027) );
  INV_X1 U7799 ( .A(n9027), .ZN(n9499) );
  NOR2_X1 U7800 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6321), .ZN(n6266) );
  AOI21_X1 U7801 ( .B1(n6321), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6266), .ZN(
        n6278) );
  INV_X1 U7802 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6267) );
  XNOR2_X1 U7803 ( .A(n6284), .B(n6267), .ZN(n6515) );
  INV_X1 U7804 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9750) );
  XNOR2_X1 U7805 ( .A(n6283), .B(n9750), .ZN(n6296) );
  NAND2_X1 U7806 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6300) );
  INV_X1 U7807 ( .A(n6300), .ZN(n6268) );
  NAND2_X1 U7808 ( .A1(n6296), .A2(n6268), .ZN(n6297) );
  NAND2_X1 U7809 ( .A1(n6283), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7810 ( .A1(n6297), .A2(n6269), .ZN(n6514) );
  AND2_X1 U7811 ( .A1(n6515), .A2(n6514), .ZN(n6516) );
  INV_X1 U7812 ( .A(n6516), .ZN(n6271) );
  NAND2_X1 U7813 ( .A1(n6284), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7814 ( .A1(n6271), .A2(n6270), .ZN(n6331) );
  INV_X1 U7815 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6272) );
  XNOR2_X1 U7816 ( .A(n6340), .B(n6272), .ZN(n6332) );
  NAND2_X1 U7817 ( .A1(n6331), .A2(n6332), .ZN(n6330) );
  NAND2_X1 U7818 ( .A1(n6340), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7819 ( .A1(n6330), .A2(n6273), .ZN(n6504) );
  XNOR2_X1 U7820 ( .A(n6509), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n6505) );
  NOR2_X1 U7821 ( .A1(n6504), .A2(n6505), .ZN(n6503) );
  NOR2_X1 U7822 ( .A1(n6509), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6274) );
  OR2_X1 U7823 ( .A1(n6503), .A2(n6274), .ZN(n9449) );
  NAND2_X1 U7824 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9458), .ZN(n6275) );
  OAI21_X1 U7825 ( .B1(n9458), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6275), .ZN(
        n9448) );
  NOR2_X1 U7826 ( .A1(n9449), .A2(n9448), .ZN(n9447) );
  AOI21_X1 U7827 ( .B1(n9458), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9447), .ZN(
        n9463) );
  INV_X1 U7828 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9862) );
  AOI22_X1 U7829 ( .A1(n9470), .A2(P1_REG1_REG_6__SCAN_IN), .B1(n9862), .B2(
        n6276), .ZN(n9462) );
  NAND2_X1 U7830 ( .A1(n9463), .A2(n9462), .ZN(n9461) );
  OAI21_X1 U7831 ( .B1(n9470), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9461), .ZN(
        n6277) );
  NAND2_X1 U7832 ( .A1(n6278), .A2(n6277), .ZN(n6320) );
  OAI21_X1 U7833 ( .B1(n6278), .B2(n6277), .A(n6320), .ZN(n6279) );
  AOI22_X1 U7834 ( .A1(n6321), .A2(n9499), .B1(n9497), .B2(n6279), .ZN(n6294)
         );
  OR2_X1 U7835 ( .A1(n6280), .A2(n6497), .ZN(n9490) );
  INV_X1 U7836 ( .A(n9490), .ZN(n9483) );
  NOR2_X1 U7837 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6321), .ZN(n6281) );
  AOI21_X1 U7838 ( .B1(n6321), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6281), .ZN(
        n6291) );
  INV_X1 U7839 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6286) );
  NOR2_X1 U7840 ( .A1(n6282), .A2(n6259), .ZN(n6498) );
  INV_X1 U7841 ( .A(n6498), .ZN(n6303) );
  XNOR2_X1 U7842 ( .A(n6284), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6513) );
  NOR2_X1 U7843 ( .A1(n4276), .A2(n6513), .ZN(n6512) );
  AOI21_X1 U7844 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6284), .A(n6512), .ZN(
        n6334) );
  XNOR2_X1 U7845 ( .A(n6340), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n6333) );
  OAI21_X1 U7846 ( .B1(n6286), .B2(n6285), .A(n6336), .ZN(n6501) );
  XNOR2_X1 U7847 ( .A(n6509), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n6502) );
  NOR2_X1 U7848 ( .A1(n6501), .A2(n6502), .ZN(n9452) );
  NOR2_X1 U7849 ( .A1(n6509), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9451) );
  NOR2_X1 U7850 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9458), .ZN(n6287) );
  AOI21_X1 U7851 ( .B1(n9458), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6287), .ZN(
        n9450) );
  OAI21_X1 U7852 ( .B1(n9452), .B2(n9451), .A(n9450), .ZN(n9454) );
  OAI21_X1 U7853 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n9458), .A(n9454), .ZN(
        n9466) );
  INV_X1 U7854 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6288) );
  MUX2_X1 U7855 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6288), .S(n9470), .Z(n6289)
         );
  INV_X1 U7856 ( .A(n6289), .ZN(n9465) );
  NOR2_X1 U7857 ( .A1(n9466), .A2(n9465), .ZN(n9464) );
  OAI21_X1 U7858 ( .B1(n6291), .B2(n6290), .A(n6313), .ZN(n6292) );
  AND2_X1 U7859 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6731) );
  AOI21_X1 U7860 ( .B1(n9483), .B2(n6292), .A(n6731), .ZN(n6293) );
  OAI211_X1 U7861 ( .C1(n9038), .C2(n6295), .A(n6294), .B(n6293), .ZN(P1_U3248) );
  INV_X1 U7862 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6309) );
  INV_X1 U7863 ( .A(n6296), .ZN(n6299) );
  INV_X1 U7864 ( .A(n6297), .ZN(n6298) );
  AOI211_X1 U7865 ( .C1(n6300), .C2(n6299), .A(n6298), .B(n9476), .ZN(n6307)
         );
  AOI211_X1 U7866 ( .C1(n6303), .C2(n6302), .A(n6301), .B(n9490), .ZN(n6306)
         );
  INV_X1 U7867 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6737) );
  OAI22_X1 U7868 ( .A1(n9027), .A2(n6304), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6737), .ZN(n6305) );
  NOR3_X1 U7869 ( .A1(n6307), .A2(n6306), .A3(n6305), .ZN(n6308) );
  OAI21_X1 U7870 ( .B1(n9038), .B2(n6309), .A(n6308), .ZN(P1_U3242) );
  INV_X1 U7871 ( .A(n6310), .ZN(n6342) );
  AOI22_X1 U7872 ( .A1(n6914), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9366), .ZN(n6311) );
  OAI21_X1 U7873 ( .B1(n6342), .B2(n8334), .A(n6311), .ZN(P1_U3340) );
  INV_X1 U7874 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6329) );
  NOR2_X1 U7875 ( .A1(n9819), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7127) );
  NOR2_X1 U7876 ( .A1(n9484), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6312) );
  AOI21_X1 U7877 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9484), .A(n6312), .ZN(
        n9475) );
  OAI21_X1 U7878 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9484), .A(n9473), .ZN(
        n9493) );
  NAND2_X1 U7879 ( .A1(n9498), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6314) );
  OAI21_X1 U7880 ( .B1(n9498), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6314), .ZN(
        n9492) );
  NOR2_X1 U7881 ( .A1(n9493), .A2(n9492), .ZN(n9491) );
  NAND2_X1 U7882 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6589), .ZN(n6315) );
  OAI21_X1 U7883 ( .B1(n6589), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6315), .ZN(
        n6316) );
  AOI211_X1 U7884 ( .C1(n6317), .C2(n6316), .A(n6588), .B(n9490), .ZN(n6318)
         );
  AOI211_X1 U7885 ( .C1(n9499), .C2(n6589), .A(n7127), .B(n6318), .ZN(n6328)
         );
  NAND2_X1 U7886 ( .A1(n9484), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6319) );
  OAI21_X1 U7887 ( .B1(n9484), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6319), .ZN(
        n9478) );
  OAI21_X1 U7888 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6321), .A(n6320), .ZN(
        n9479) );
  NOR2_X1 U7889 ( .A1(n9478), .A2(n9479), .ZN(n9477) );
  AOI21_X1 U7890 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9484), .A(n9477), .ZN(
        n9489) );
  NOR2_X1 U7891 ( .A1(n9498), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6322) );
  AOI21_X1 U7892 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9498), .A(n6322), .ZN(
        n9488) );
  NAND2_X1 U7893 ( .A1(n9489), .A2(n9488), .ZN(n9487) );
  OAI21_X1 U7894 ( .B1(n9498), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9487), .ZN(
        n6325) );
  INV_X1 U7895 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9404) );
  AOI22_X1 U7896 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6589), .B1(n6323), .B2(
        n9404), .ZN(n6324) );
  NAND2_X1 U7897 ( .A1(n6324), .A2(n6325), .ZN(n6582) );
  OAI21_X1 U7898 ( .B1(n6325), .B2(n6324), .A(n6582), .ZN(n6326) );
  NAND2_X1 U7899 ( .A1(n6326), .A2(n9497), .ZN(n6327) );
  OAI211_X1 U7900 ( .C1(n9038), .C2(n6329), .A(n6328), .B(n6327), .ZN(P1_U3251) );
  INV_X1 U7901 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n7139) );
  AND2_X1 U7902 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6686) );
  OAI211_X1 U7903 ( .C1(n6332), .C2(n6331), .A(n9497), .B(n6330), .ZN(n6338)
         );
  NAND2_X1 U7904 ( .A1(n6334), .A2(n6333), .ZN(n6335) );
  NAND3_X1 U7905 ( .A1(n9483), .A2(n6336), .A3(n6335), .ZN(n6337) );
  NAND2_X1 U7906 ( .A1(n6338), .A2(n6337), .ZN(n6339) );
  AOI211_X1 U7907 ( .C1(n9499), .C2(n6340), .A(n6686), .B(n6339), .ZN(n6341)
         );
  OAI21_X1 U7908 ( .B1(n7139), .B2(n9038), .A(n6341), .ZN(P1_U3244) );
  INV_X1 U7909 ( .A(n7350), .ZN(n7908) );
  OAI222_X1 U7910 ( .A1(n8856), .A2(n6343), .B1(n8098), .B2(n6342), .C1(n7908), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U7911 ( .A(n6344), .ZN(n6346) );
  INV_X1 U7912 ( .A(n8053), .ZN(n7353) );
  OAI222_X1 U7913 ( .A1(n8856), .A2(n6345), .B1(n8098), .B2(n6346), .C1(n7353), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U7914 ( .A(n7166), .ZN(n7172) );
  OAI222_X1 U7915 ( .A1(n8333), .A2(n9759), .B1(n8334), .B2(n6346), .C1(n7172), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  XNOR2_X1 U7916 ( .A(n6348), .B(n6347), .ZN(n6359) );
  INV_X1 U7917 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8717) );
  OR2_X1 U7918 ( .A1(n6349), .A2(P2_U3152), .ZN(n6352) );
  OR2_X1 U7919 ( .A1(n6350), .A2(n9589), .ZN(n6351) );
  NAND2_X1 U7920 ( .A1(n6352), .A2(n6351), .ZN(n8358) );
  INV_X1 U7921 ( .A(n8720), .ZN(n6487) );
  INV_X1 U7922 ( .A(n8396), .ZN(n6355) );
  OR2_X1 U7923 ( .A1(n6628), .A2(n8693), .ZN(n6354) );
  OR2_X1 U7924 ( .A1(n6485), .A2(n8695), .ZN(n6353) );
  NAND2_X1 U7925 ( .A1(n6354), .A2(n6353), .ZN(n6533) );
  AOI22_X1 U7926 ( .A1(n6355), .A2(n6533), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3152), .ZN(n6356) );
  OAI21_X1 U7927 ( .B1(n6487), .B2(n8422), .A(n6356), .ZN(n6357) );
  AOI21_X1 U7928 ( .B1(n8717), .B2(n8358), .A(n6357), .ZN(n6358) );
  OAI21_X1 U7929 ( .B1(n8408), .B2(n6359), .A(n6358), .ZN(P2_U3220) );
  NOR2_X1 U7930 ( .A1(n9589), .A2(n6360), .ZN(n8324) );
  NAND2_X1 U7931 ( .A1(n6361), .A2(n8324), .ZN(n6407) );
  OR3_X1 U7932 ( .A1(n6406), .A2(n6362), .A3(n6407), .ZN(n6385) );
  INV_X2 U7933 ( .A(n9698), .ZN(n9700) );
  INV_X1 U7934 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6384) );
  XNOR2_X1 U7935 ( .A(n8326), .B(n6364), .ZN(n6365) );
  NAND2_X1 U7936 ( .A1(n6365), .A2(n4864), .ZN(n9571) );
  INV_X1 U7937 ( .A(n8319), .ZN(n6415) );
  NAND2_X1 U7938 ( .A1(n6366), .A2(n6415), .ZN(n9681) );
  NAND2_X1 U7939 ( .A1(n9571), .A2(n9681), .ZN(n9697) );
  INV_X1 U7940 ( .A(n6367), .ZN(n6371) );
  NAND2_X1 U7941 ( .A1(n6441), .A2(n6371), .ZN(n8140) );
  NAND2_X1 U7942 ( .A1(n8136), .A2(n8140), .ZN(n6375) );
  NAND2_X1 U7943 ( .A1(n6375), .A2(n6368), .ZN(n6440) );
  OAI21_X1 U7944 ( .B1(n6375), .B2(n6368), .A(n6440), .ZN(n6418) );
  NAND2_X1 U7945 ( .A1(n6457), .A2(n9627), .ZN(n6369) );
  INV_X1 U7946 ( .A(n8282), .ZN(n8318) );
  OR2_X1 U7947 ( .A1(n4865), .A2(n8318), .ZN(n9692) );
  INV_X1 U7948 ( .A(n9692), .ZN(n9650) );
  NAND2_X1 U7949 ( .A1(n6369), .A2(n9650), .ZN(n6370) );
  NOR2_X1 U7950 ( .A1(n6457), .A2(n9627), .ZN(n6447) );
  OR2_X1 U7951 ( .A1(n6370), .A2(n6447), .ZN(n6411) );
  OAI21_X1 U7952 ( .B1(n6371), .B2(n9690), .A(n6411), .ZN(n6382) );
  INV_X1 U7953 ( .A(n6379), .ZN(n6372) );
  NAND2_X1 U7954 ( .A1(n6373), .A2(n8136), .ZN(n6444) );
  INV_X1 U7955 ( .A(n8140), .ZN(n6378) );
  INV_X1 U7956 ( .A(n6373), .ZN(n6374) );
  NAND2_X1 U7957 ( .A1(n6375), .A2(n6374), .ZN(n6377) );
  NAND2_X1 U7958 ( .A1(n8318), .A2(n8315), .ZN(n8121) );
  AND2_X1 U7959 ( .A1(n6376), .A2(n8121), .ZN(n8643) );
  OAI211_X1 U7960 ( .C1(n6444), .C2(n6378), .A(n6377), .B(n8492), .ZN(n6381)
         );
  INV_X1 U7961 ( .A(n8695), .ZN(n8678) );
  AOI22_X1 U7962 ( .A1(n8440), .A2(n8680), .B1(n8678), .B2(n6379), .ZN(n6380)
         );
  NAND2_X1 U7963 ( .A1(n6381), .A2(n6380), .ZN(n6414) );
  AOI211_X1 U7964 ( .C1(n9697), .C2(n6418), .A(n6382), .B(n6414), .ZN(n6386)
         );
  OR2_X1 U7965 ( .A1(n6386), .A2(n9698), .ZN(n6383) );
  OAI21_X1 U7966 ( .B1(n9700), .B2(n6384), .A(n6383), .ZN(P2_U3454) );
  INV_X2 U7967 ( .A(n9713), .ZN(n9715) );
  INV_X1 U7968 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6388) );
  OR2_X1 U7969 ( .A1(n6386), .A2(n9713), .ZN(n6387) );
  OAI21_X1 U7970 ( .B1(n9715), .B2(n6388), .A(n6387), .ZN(P2_U3521) );
  INV_X1 U7971 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6389) );
  NAND2_X1 U7972 ( .A1(n8453), .A2(n6389), .ZN(n6390) );
  OAI211_X1 U7973 ( .C1(n6391), .C2(P2_REG2_REG_0__SCAN_IN), .A(n6390), .B(
        n8448), .ZN(n6396) );
  INV_X1 U7974 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U7975 ( .A1(n8453), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6392) );
  OAI21_X1 U7976 ( .B1(n8450), .B2(n6393), .A(n6392), .ZN(n6395) );
  INV_X1 U7977 ( .A(n8859), .ZN(n6394) );
  MUX2_X1 U7978 ( .A(n6396), .B(n6395), .S(n6394), .Z(n6399) );
  INV_X1 U7979 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6397) );
  INV_X1 U7980 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6659) );
  OAI22_X1 U7981 ( .A1(n8460), .A2(n6397), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6659), .ZN(n6398) );
  OR2_X1 U7982 ( .A1(n6399), .A2(n6398), .ZN(P2_U3245) );
  OAI21_X1 U7983 ( .B1(n6402), .B2(n6401), .A(n6400), .ZN(n6494) );
  INV_X1 U7984 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6793) );
  OAI22_X1 U7985 ( .A1(n6609), .A2(n6793), .B1(n7832), .B2(n8954), .ZN(n6403)
         );
  AOI21_X1 U7986 ( .B1(n8926), .B2(n6494), .A(n6403), .ZN(n6404) );
  OAI21_X1 U7987 ( .B1(n6570), .B2(n8960), .A(n6404), .ZN(P1_U3230) );
  NAND2_X1 U7988 ( .A1(n6406), .A2(n6405), .ZN(n6408) );
  OR2_X1 U7989 ( .A1(n6408), .A2(n6407), .ZN(n6410) );
  NOR2_X1 U7990 ( .A1(n8699), .A2(n6409), .ZN(n6413) );
  OR2_X1 U7991 ( .A1(n6410), .A2(n8567), .ZN(n9583) );
  INV_X1 U7992 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n8086) );
  OAI22_X1 U7993 ( .A1(n9583), .A2(n6411), .B1(n8086), .B2(n8705), .ZN(n6412)
         );
  AOI211_X1 U7994 ( .C1(n8699), .C2(n6414), .A(n6413), .B(n6412), .ZN(n6420)
         );
  NAND2_X1 U7995 ( .A1(n6415), .A2(n8315), .ZN(n6808) );
  NAND2_X1 U7996 ( .A1(n9571), .A2(n6808), .ZN(n6416) );
  NAND2_X1 U7997 ( .A1(n8699), .A2(n6416), .ZN(n8686) );
  INV_X1 U7998 ( .A(n8686), .ZN(n8711) );
  NAND2_X1 U7999 ( .A1(n8699), .A2(n6417), .ZN(n8674) );
  AOI22_X1 U8000 ( .A1(n8711), .A2(n6418), .B1(n9577), .B2(n6457), .ZN(n6419)
         );
  NAND2_X1 U8001 ( .A1(n6420), .A2(n6419), .ZN(P2_U3295) );
  NOR2_X1 U8002 ( .A1(n8358), .A2(P2_U3152), .ZN(n6460) );
  INV_X1 U8003 ( .A(n9627), .ZN(n6422) );
  NAND2_X1 U8004 ( .A1(n6379), .A2(n6422), .ZN(n8139) );
  MUX2_X1 U8005 ( .A(n8139), .B(n6422), .S(n6421), .Z(n6423) );
  AOI21_X1 U8006 ( .B1(n6373), .B2(n6423), .A(n8408), .ZN(n6425) );
  NOR2_X1 U8007 ( .A1(n8414), .A2(n6427), .ZN(n6424) );
  AOI211_X1 U8008 ( .C1(n9627), .C2(n8406), .A(n6425), .B(n6424), .ZN(n6426)
         );
  OAI21_X1 U8009 ( .B1(n6460), .B2(n6659), .A(n6426), .ZN(P2_U3234) );
  OAI22_X1 U8010 ( .A1(n6427), .A2(n8416), .B1(n8414), .B2(n6488), .ZN(n6431)
         );
  INV_X1 U8011 ( .A(n6450), .ZN(n9636) );
  XNOR2_X1 U8012 ( .A(n6428), .B(n4266), .ZN(n6429) );
  OAI22_X1 U8013 ( .A1(n8422), .A2(n9636), .B1(n6429), .B2(n8408), .ZN(n6430)
         );
  NOR2_X1 U8014 ( .A1(n6431), .A2(n6430), .ZN(n6432) );
  OAI21_X1 U8015 ( .B1(n6460), .B2(n6448), .A(n6432), .ZN(P2_U3239) );
  AOI21_X1 U8016 ( .B1(n6434), .B2(n6433), .A(n4320), .ZN(n6439) );
  NAND2_X1 U8017 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7986) );
  OAI21_X1 U8018 ( .B1(n8422), .B2(n9640), .A(n7986), .ZN(n6436) );
  OAI22_X1 U8019 ( .A1(n6488), .A2(n8416), .B1(n8414), .B2(n8696), .ZN(n6435)
         );
  AOI211_X1 U8020 ( .C1(n6437), .C2(n8358), .A(n6436), .B(n6435), .ZN(n6438)
         );
  OAI21_X1 U8021 ( .B1(n6439), .B2(n8408), .A(n6438), .ZN(P2_U3232) );
  NAND2_X1 U8022 ( .A1(n6440), .A2(n6457), .ZN(n6484) );
  NAND2_X1 U8023 ( .A1(n6442), .A2(n6441), .ZN(n6482) );
  NAND2_X1 U8024 ( .A1(n6484), .A2(n6482), .ZN(n6443) );
  NAND2_X1 U8025 ( .A1(n8440), .A2(n9636), .ZN(n8137) );
  AND2_X1 U8026 ( .A1(n8137), .A2(n8142), .ZN(n8286) );
  XNOR2_X1 U8027 ( .A(n6443), .B(n6481), .ZN(n9633) );
  NAND2_X1 U8028 ( .A1(n6445), .A2(n8286), .ZN(n6530) );
  OAI21_X1 U8029 ( .B1(n6445), .B2(n8286), .A(n6530), .ZN(n6446) );
  INV_X1 U8030 ( .A(n6488), .ZN(n8439) );
  AOI222_X1 U8031 ( .A1(n8492), .A2(n6446), .B1(n8439), .B2(n8680), .C1(n6441), 
        .C2(n8678), .ZN(n9635) );
  MUX2_X1 U8032 ( .A(n6173), .B(n9635), .S(n8699), .Z(n6452) );
  NAND2_X1 U8033 ( .A1(n6447), .A2(n9636), .ZN(n6538) );
  OAI211_X1 U8034 ( .C1(n6447), .C2(n9636), .A(n6538), .B(n9650), .ZN(n9634)
         );
  OAI22_X1 U8035 ( .A1(n9583), .A2(n9634), .B1(n6448), .B2(n8705), .ZN(n6449)
         );
  AOI21_X1 U8036 ( .B1(n9577), .B2(n6450), .A(n6449), .ZN(n6451) );
  OAI211_X1 U8037 ( .C1(n8686), .C2(n9633), .A(n6452), .B(n6451), .ZN(P2_U3294) );
  AOI22_X1 U8038 ( .A1(n8375), .A2(n6379), .B1(n8374), .B2(n8440), .ZN(n6459)
         );
  OAI21_X1 U8039 ( .B1(n6453), .B2(n6454), .A(n6455), .ZN(n6456) );
  AOI22_X1 U8040 ( .A1(n8406), .A2(n6457), .B1(n8410), .B2(n6456), .ZN(n6458)
         );
  OAI211_X1 U8041 ( .C1(n6460), .C2(n8086), .A(n6459), .B(n6458), .ZN(P2_U3224) );
  INV_X1 U8042 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U8043 ( .A1(n8507), .A2(P2_U3966), .ZN(n6461) );
  OAI21_X1 U8044 ( .B1(n8332), .B2(P2_U3966), .A(n6461), .ZN(P2_U3581) );
  XNOR2_X1 U8045 ( .A(n6463), .B(n6462), .ZN(n6470) );
  INV_X1 U8046 ( .A(n6778), .ZN(n6637) );
  OR2_X1 U8047 ( .A1(n6628), .A2(n8695), .ZN(n6465) );
  OR2_X1 U8048 ( .A1(n6788), .A2(n8693), .ZN(n6464) );
  NAND2_X1 U8049 ( .A1(n6465), .A2(n6464), .ZN(n6634) );
  INV_X1 U8050 ( .A(n6634), .ZN(n6466) );
  OAI22_X1 U8051 ( .A1(n8396), .A2(n6466), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8073), .ZN(n6467) );
  AOI21_X1 U8052 ( .B1(n8406), .B2(n6637), .A(n6467), .ZN(n6469) );
  NAND2_X1 U8053 ( .A1(n8358), .A2(n6644), .ZN(n6468) );
  OAI211_X1 U8054 ( .C1(n6470), .C2(n8408), .A(n6469), .B(n6468), .ZN(P2_U3229) );
  NAND2_X1 U8055 ( .A1(n6530), .A2(n8142), .ZN(n6471) );
  NAND2_X1 U8056 ( .A1(n6532), .A2(n8132), .ZN(n6631) );
  NAND2_X1 U8057 ( .A1(n6628), .A2(n6480), .ZN(n8133) );
  INV_X1 U8058 ( .A(n6628), .ZN(n8438) );
  NAND2_X1 U8059 ( .A1(n8438), .A2(n9640), .ZN(n6784) );
  NAND2_X1 U8060 ( .A1(n8133), .A2(n6784), .ZN(n6489) );
  INV_X1 U8061 ( .A(n6489), .ZN(n8287) );
  XNOR2_X1 U8062 ( .A(n6631), .B(n8287), .ZN(n6472) );
  NAND2_X1 U8063 ( .A1(n6472), .A2(n8492), .ZN(n6475) );
  OAI22_X1 U8064 ( .A1(n6488), .A2(n8695), .B1(n8696), .B2(n8693), .ZN(n6473)
         );
  INV_X1 U8065 ( .A(n6473), .ZN(n6474) );
  NAND2_X1 U8066 ( .A1(n6475), .A2(n6474), .ZN(n9642) );
  INV_X1 U8067 ( .A(n9642), .ZN(n6493) );
  INV_X1 U8068 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n9847) );
  OAI22_X1 U8069 ( .A1(n8705), .A2(n6476), .B1(n9847), .B2(n8699), .ZN(n6479)
         );
  OR2_X1 U8070 ( .A1(n9583), .A2(n9692), .ZN(n8707) );
  INV_X1 U8071 ( .A(n6779), .ZN(n6477) );
  OAI21_X1 U8072 ( .B1(n9640), .B2(n6537), .A(n6477), .ZN(n9641) );
  NOR2_X1 U8073 ( .A1(n8707), .A2(n9641), .ZN(n6478) );
  AOI211_X1 U8074 ( .C1(n9577), .C2(n6480), .A(n6479), .B(n6478), .ZN(n6492)
         );
  AND2_X1 U8075 ( .A1(n6482), .A2(n6481), .ZN(n6483) );
  NAND2_X1 U8076 ( .A1(n6485), .A2(n9636), .ZN(n6486) );
  NAND2_X1 U8077 ( .A1(n6490), .A2(n6489), .ZN(n6630) );
  OAI21_X1 U8078 ( .B1(n6490), .B2(n6489), .A(n6630), .ZN(n9644) );
  NAND2_X1 U8079 ( .A1(n9644), .A2(n8711), .ZN(n6491) );
  OAI211_X1 U8080 ( .C1(n9588), .C2(n6493), .A(n6492), .B(n6491), .ZN(P2_U3292) );
  INV_X1 U8081 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U8082 ( .A1(n6494), .A2(n6497), .ZN(n6496) );
  OAI211_X1 U8083 ( .C1(n6498), .C2(n6497), .A(n6496), .B(n6495), .ZN(n6499)
         );
  OAI211_X1 U8084 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6500), .A(n6499), .B(
        P1_U4006), .ZN(n6525) );
  AND2_X1 U8085 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6718) );
  AOI21_X1 U8086 ( .B1(n6502), .B2(n6501), .A(n9452), .ZN(n6507) );
  AOI21_X1 U8087 ( .B1(n6505), .B2(n6504), .A(n6503), .ZN(n6506) );
  OAI22_X1 U8088 ( .A1(n6507), .A2(n9490), .B1(n9476), .B2(n6506), .ZN(n6508)
         );
  AOI211_X1 U8089 ( .C1(n9499), .C2(n6509), .A(n6718), .B(n6508), .ZN(n6510)
         );
  OAI211_X1 U8090 ( .C1(n9038), .C2(n6511), .A(n6525), .B(n6510), .ZN(P1_U3245) );
  INV_X1 U8091 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6526) );
  AOI211_X1 U8092 ( .C1(n4276), .C2(n6513), .A(n6512), .B(n9490), .ZN(n6523)
         );
  INV_X1 U8093 ( .A(n6514), .ZN(n6518) );
  INV_X1 U8094 ( .A(n6515), .ZN(n6517) );
  AOI211_X1 U8095 ( .C1(n6518), .C2(n6517), .A(n6516), .B(n9476), .ZN(n6522)
         );
  INV_X1 U8096 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6519) );
  OAI22_X1 U8097 ( .A1(n9027), .A2(n6520), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6519), .ZN(n6521) );
  NOR3_X1 U8098 ( .A1(n6523), .A2(n6522), .A3(n6521), .ZN(n6524) );
  OAI211_X1 U8099 ( .C1(n9038), .C2(n6526), .A(n6525), .B(n6524), .ZN(P1_U3243) );
  INV_X1 U8100 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6543) );
  OR2_X1 U8101 ( .A1(n6527), .A2(n8284), .ZN(n6528) );
  NAND2_X1 U8102 ( .A1(n6529), .A2(n6528), .ZN(n8721) );
  INV_X1 U8103 ( .A(n8721), .ZN(n6541) );
  INV_X1 U8104 ( .A(n9571), .ZN(n7429) );
  NAND2_X1 U8105 ( .A1(n8721), .A2(n7429), .ZN(n6536) );
  NAND3_X1 U8106 ( .A1(n6530), .A2(n8284), .A3(n8142), .ZN(n6531) );
  NAND2_X1 U8107 ( .A1(n6532), .A2(n6531), .ZN(n6534) );
  AOI21_X1 U8108 ( .B1(n6534), .B2(n8492), .A(n6533), .ZN(n6535) );
  NAND2_X1 U8109 ( .A1(n6536), .A2(n6535), .ZN(n8715) );
  INV_X1 U8110 ( .A(n8715), .ZN(n6540) );
  AOI21_X1 U8111 ( .B1(n8720), .B2(n6538), .A(n6537), .ZN(n8718) );
  AOI22_X1 U8112 ( .A1(n8718), .A2(n9650), .B1(n9677), .B2(n8720), .ZN(n6539)
         );
  OAI211_X1 U8113 ( .C1(n6541), .C2(n9681), .A(n6540), .B(n6539), .ZN(n6544)
         );
  NAND2_X1 U8114 ( .A1(n6544), .A2(n9700), .ZN(n6542) );
  OAI21_X1 U8115 ( .B1(n9700), .B2(n6543), .A(n6542), .ZN(P2_U3460) );
  INV_X1 U8116 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8117 ( .A1(n6544), .A2(n9715), .ZN(n6545) );
  OAI21_X1 U8118 ( .B1(n9715), .B2(n6546), .A(n6545), .ZN(P2_U3523) );
  NAND2_X1 U8119 ( .A1(n6547), .A2(n6555), .ZN(n6548) );
  INV_X2 U8120 ( .A(n9548), .ZN(n9550) );
  INV_X1 U8121 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6554) );
  AND2_X1 U8122 ( .A1(n6575), .A2(n6570), .ZN(n7829) );
  NOR2_X1 U8123 ( .A1(n6573), .A2(n7829), .ZN(n7794) );
  NAND2_X1 U8124 ( .A1(n6871), .A2(n6552), .ZN(n6549) );
  OR2_X1 U8125 ( .A1(n7794), .A2(n6549), .ZN(n6551) );
  INV_X1 U8126 ( .A(n9376), .ZN(n9407) );
  NAND2_X1 U8127 ( .A1(n8976), .A2(n9407), .ZN(n6550) );
  AND2_X1 U8128 ( .A1(n6551), .A2(n6550), .ZN(n6792) );
  OAI21_X1 U8129 ( .B1(n6570), .B2(n6552), .A(n6792), .ZN(n6559) );
  NAND2_X1 U8130 ( .A1(n6559), .A2(n9550), .ZN(n6553) );
  OAI21_X1 U8131 ( .B1(n9550), .B2(n6554), .A(n6553), .ZN(P1_U3454) );
  NAND2_X1 U8132 ( .A1(n6556), .A2(n6555), .ZN(n6557) );
  INV_X2 U8133 ( .A(n9559), .ZN(n9562) );
  NAND2_X1 U8134 ( .A1(n6559), .A2(n9562), .ZN(n6560) );
  OAI21_X1 U8135 ( .B1(n9562), .B2(n6561), .A(n6560), .ZN(P1_U3523) );
  INV_X1 U8136 ( .A(n6562), .ZN(n6564) );
  OAI222_X1 U8137 ( .A1(n8333), .A2(n6563), .B1(n8334), .B2(n6564), .C1(
        P1_U3084), .C2(n7249), .ZN(P1_U3338) );
  INV_X1 U8138 ( .A(n7354), .ZN(n8039) );
  OAI222_X1 U8139 ( .A1(n8856), .A2(n6565), .B1(n8098), .B2(n6564), .C1(
        P2_U3152), .C2(n8039), .ZN(P2_U3343) );
  INV_X1 U8140 ( .A(n6566), .ZN(n6603) );
  AOI22_X1 U8141 ( .A1(n9013), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9366), .ZN(n6567) );
  OAI21_X1 U8142 ( .B1(n6603), .B2(n8334), .A(n6567), .ZN(P1_U3336) );
  INV_X1 U8143 ( .A(n9335), .ZN(n9538) );
  OAI21_X1 U8144 ( .B1(n7799), .B2(n6569), .A(n6568), .ZN(n6743) );
  INV_X1 U8145 ( .A(n6743), .ZN(n6580) );
  INV_X1 U8146 ( .A(n9520), .ZN(n9540) );
  NOR2_X1 U8147 ( .A1(n7568), .A2(n6570), .ZN(n6571) );
  OR3_X1 U8148 ( .A1(n6571), .A2(n6938), .A3(n9542), .ZN(n6738) );
  OAI21_X1 U8149 ( .B1(n7568), .B2(n9540), .A(n6738), .ZN(n6579) );
  OAI21_X1 U8150 ( .B1(n6574), .B2(n6573), .A(n6572), .ZN(n6577) );
  INV_X1 U8151 ( .A(n9203), .ZN(n9412) );
  INV_X1 U8152 ( .A(n6575), .ZN(n7563) );
  OAI22_X1 U8153 ( .A1(n7563), .A2(n9378), .B1(n6133), .B2(n9376), .ZN(n6576)
         );
  AOI21_X1 U8154 ( .B1(n6577), .B2(n9412), .A(n6576), .ZN(n6578) );
  OAI21_X1 U8155 ( .B1(n9382), .B2(n6743), .A(n6578), .ZN(n6740) );
  AOI211_X1 U8156 ( .C1(n9538), .C2(n6580), .A(n6579), .B(n6740), .ZN(n6617)
         );
  NAND2_X1 U8157 ( .A1(n9559), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6581) );
  OAI21_X1 U8158 ( .B1(n6617), .B2(n9559), .A(n6581), .ZN(P1_U3524) );
  INV_X1 U8159 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9443) );
  AOI22_X1 U8160 ( .A1(n6590), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n9443), .B2(
        n8982), .ZN(n8987) );
  OAI21_X1 U8161 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6589), .A(n6582), .ZN(
        n8986) );
  NAND2_X1 U8162 ( .A1(n8987), .A2(n8986), .ZN(n8985) );
  OAI21_X1 U8163 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6590), .A(n8985), .ZN(
        n6584) );
  MUX2_X1 U8164 ( .A(n9436), .B(P1_REG1_REG_12__SCAN_IN), .S(n6586), .Z(n6583)
         );
  NAND2_X1 U8165 ( .A1(n6583), .A2(n6584), .ZN(n6669) );
  OAI21_X1 U8166 ( .B1(n6584), .B2(n6583), .A(n6669), .ZN(n6596) );
  INV_X1 U8167 ( .A(n9038), .ZN(n9500) );
  NAND2_X1 U8168 ( .A1(n9500), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6585) );
  NAND2_X1 U8169 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3084), .ZN(n7288) );
  OAI211_X1 U8170 ( .C1(n9027), .C2(n6586), .A(n6585), .B(n7288), .ZN(n6595)
         );
  INV_X1 U8171 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6587) );
  AOI22_X1 U8172 ( .A1(n6590), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n6587), .B2(
        n8982), .ZN(n8979) );
  OAI21_X1 U8173 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6590), .A(n8977), .ZN(
        n6593) );
  NAND2_X1 U8174 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6674), .ZN(n6591) );
  OAI21_X1 U8175 ( .B1(n6674), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6591), .ZN(
        n6592) );
  NOR2_X1 U8176 ( .A1(n6592), .A2(n6593), .ZN(n6673) );
  AOI211_X1 U8177 ( .C1(n6593), .C2(n6592), .A(n6673), .B(n9490), .ZN(n6594)
         );
  AOI211_X1 U8178 ( .C1(n9497), .C2(n6596), .A(n6595), .B(n6594), .ZN(n6597)
         );
  INV_X1 U8179 ( .A(n6597), .ZN(P1_U3253) );
  INV_X1 U8180 ( .A(n8996), .ZN(n7255) );
  INV_X1 U8181 ( .A(n6598), .ZN(n6600) );
  OAI222_X1 U8182 ( .A1(P1_U3084), .A2(n7255), .B1(n8334), .B2(n6600), .C1(
        n6599), .C2(n8333), .ZN(P1_U3337) );
  INV_X1 U8183 ( .A(n7884), .ZN(n7363) );
  OAI222_X1 U8184 ( .A1(n8856), .A2(n9838), .B1(n8098), .B2(n6600), .C1(n7363), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8185 ( .A(n6601), .ZN(n6615) );
  AOI22_X1 U8186 ( .A1(n9025), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9366), .ZN(n6602) );
  OAI21_X1 U8187 ( .B1(n6615), .B2(n8334), .A(n6602), .ZN(P1_U3335) );
  OAI222_X1 U8188 ( .A1(n8856), .A2(n6604), .B1(n8098), .B2(n6603), .C1(n8016), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8189 ( .A(n6605), .ZN(n6606) );
  AOI21_X1 U8190 ( .B1(n6608), .B2(n6607), .A(n6606), .ZN(n6613) );
  INV_X1 U8191 ( .A(n6609), .ZN(n7565) );
  NAND2_X1 U8192 ( .A1(n9520), .A2(n6941), .ZN(n9505) );
  INV_X1 U8193 ( .A(n8954), .ZN(n8928) );
  AOI22_X1 U8194 ( .A1(n8974), .A2(n8928), .B1(n8940), .B2(n8976), .ZN(n6610)
         );
  OAI21_X1 U8195 ( .B1(n7565), .B2(n9505), .A(n6610), .ZN(n6611) );
  AOI21_X1 U8196 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7565), .A(n6611), .ZN(
        n6612) );
  OAI21_X1 U8197 ( .B1(n6613), .B2(n8947), .A(n6612), .ZN(P1_U3235) );
  INV_X1 U8198 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8855) );
  INV_X1 U8199 ( .A(n9105), .ZN(n7707) );
  NAND2_X1 U8200 ( .A1(n7707), .A2(P1_U4006), .ZN(n6614) );
  OAI21_X1 U8201 ( .B1(n8855), .B2(P1_U4006), .A(n6614), .ZN(P1_U3584) );
  INV_X1 U8202 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6616) );
  INV_X1 U8203 ( .A(n8446), .ZN(n8026) );
  OAI222_X1 U8204 ( .A1(n8856), .A2(n6616), .B1(n8098), .B2(n6615), .C1(
        P2_U3152), .C2(n8026), .ZN(P2_U3340) );
  INV_X1 U8205 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6619) );
  OR2_X1 U8206 ( .A1(n6617), .A2(n9548), .ZN(n6618) );
  OAI21_X1 U8207 ( .B1(n9550), .B2(n6619), .A(n6618), .ZN(P1_U3457) );
  OAI21_X1 U8208 ( .B1(n6622), .B2(n6621), .A(n6620), .ZN(n6626) );
  OAI22_X1 U8209 ( .A1(n8696), .A2(n8416), .B1(n8414), .B2(n8694), .ZN(n6625)
         );
  INV_X1 U8210 ( .A(n9649), .ZN(n8700) );
  NAND2_X1 U8211 ( .A1(n8358), .A2(n8704), .ZN(n6623) );
  NAND2_X1 U8212 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7975) );
  OAI211_X1 U8213 ( .C1(n8700), .C2(n8422), .A(n6623), .B(n7975), .ZN(n6624)
         );
  AOI211_X1 U8214 ( .C1(n6626), .C2(n8410), .A(n6625), .B(n6624), .ZN(n6627)
         );
  INV_X1 U8215 ( .A(n6627), .ZN(P2_U3241) );
  INV_X1 U8216 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6640) );
  NAND2_X1 U8217 ( .A1(n8696), .A2(n6637), .ZN(n8689) );
  INV_X1 U8218 ( .A(n8696), .ZN(n8437) );
  NAND2_X1 U8219 ( .A1(n8437), .A2(n6778), .ZN(n8151) );
  NAND2_X1 U8220 ( .A1(n8689), .A2(n8151), .ZN(n8289) );
  NAND2_X1 U8221 ( .A1(n6628), .A2(n9640), .ZN(n6629) );
  XOR2_X1 U8222 ( .A(n8289), .B(n6775), .Z(n6652) );
  INV_X1 U8223 ( .A(n9697), .ZN(n8816) );
  INV_X1 U8224 ( .A(n6631), .ZN(n6632) );
  NAND2_X1 U8225 ( .A1(n8688), .A2(n6784), .ZN(n6633) );
  XNOR2_X1 U8226 ( .A(n6633), .B(n8289), .ZN(n6635) );
  AOI21_X1 U8227 ( .B1(n6635), .B2(n8492), .A(n6634), .ZN(n6648) );
  XNOR2_X1 U8228 ( .A(n6779), .B(n6778), .ZN(n6636) );
  NOR2_X1 U8229 ( .A1(n6636), .A2(n9692), .ZN(n6645) );
  AOI21_X1 U8230 ( .B1(n9677), .B2(n6637), .A(n6645), .ZN(n6638) );
  OAI211_X1 U8231 ( .C1(n6652), .C2(n8816), .A(n6648), .B(n6638), .ZN(n6641)
         );
  NAND2_X1 U8232 ( .A1(n6641), .A2(n9700), .ZN(n6639) );
  OAI21_X1 U8233 ( .B1(n9700), .B2(n6640), .A(n6639), .ZN(P2_U3466) );
  INV_X1 U8234 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U8235 ( .A1(n6641), .A2(n9715), .ZN(n6642) );
  OAI21_X1 U8236 ( .B1(n9715), .B2(n6643), .A(n6642), .ZN(P2_U3525) );
  NOR2_X1 U8237 ( .A1(n9588), .A2(n8567), .ZN(n8667) );
  INV_X1 U8238 ( .A(n8705), .ZN(n9576) );
  AOI22_X1 U8239 ( .A1(n8667), .A2(n6645), .B1(n6644), .B2(n9576), .ZN(n6646)
         );
  OAI21_X1 U8240 ( .B1(n6778), .B2(n8674), .A(n6646), .ZN(n6647) );
  INV_X1 U8241 ( .A(n6647), .ZN(n6651) );
  INV_X1 U8242 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6649) );
  MUX2_X1 U8243 ( .A(n6649), .B(n6648), .S(n8699), .Z(n6650) );
  OAI211_X1 U8244 ( .C1(n6652), .C2(n8686), .A(n6651), .B(n6650), .ZN(P2_U3291) );
  XNOR2_X1 U8245 ( .A(n6654), .B(n6653), .ZN(n6658) );
  INV_X1 U8246 ( .A(n6782), .ZN(n9657) );
  OAI22_X1 U8247 ( .A1(n8422), .A2(n9657), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7963), .ZN(n6656) );
  OAI22_X1 U8248 ( .A1(n6788), .A2(n8416), .B1(n8414), .B2(n6966), .ZN(n6655)
         );
  AOI211_X1 U8249 ( .C1(n6781), .C2(n8358), .A(n6656), .B(n6655), .ZN(n6657)
         );
  OAI21_X1 U8250 ( .B1(n6658), .B2(n8408), .A(n6657), .ZN(P2_U3215) );
  NAND2_X1 U8251 ( .A1(n6373), .A2(n8139), .ZN(n9629) );
  INV_X1 U8252 ( .A(n9629), .ZN(n6663) );
  AOI22_X1 U8253 ( .A1(n9629), .A2(n8492), .B1(n8680), .B2(n6441), .ZN(n9631)
         );
  OAI22_X1 U8254 ( .A1(n9588), .A2(n9631), .B1(n6659), .B2(n8705), .ZN(n6660)
         );
  AOI21_X1 U8255 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n9588), .A(n6660), .ZN(
        n6662) );
  INV_X1 U8256 ( .A(n8707), .ZN(n8719) );
  OAI21_X1 U8257 ( .B1(n8719), .B2(n9577), .A(n9627), .ZN(n6661) );
  OAI211_X1 U8258 ( .C1(n6663), .C2(n8686), .A(n6662), .B(n6661), .ZN(P2_U3296) );
  INV_X1 U8259 ( .A(n6664), .ZN(n6666) );
  OAI222_X1 U8260 ( .A1(n8856), .A2(n6665), .B1(n8098), .B2(n6666), .C1(n4864), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8261 ( .A1(n8333), .A2(n6667), .B1(n8334), .B2(n6666), .C1(
        P1_U3084), .C2(n9033), .ZN(P1_U3334) );
  INV_X1 U8262 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6682) );
  INV_X1 U8263 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6668) );
  MUX2_X1 U8264 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6668), .S(n6914), .Z(n6671)
         );
  OAI21_X1 U8265 ( .B1(n6674), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6669), .ZN(
        n6670) );
  NAND2_X1 U8266 ( .A1(n6671), .A2(n6670), .ZN(n6910) );
  OAI21_X1 U8267 ( .B1(n6671), .B2(n6670), .A(n6910), .ZN(n6680) );
  INV_X1 U8268 ( .A(n6914), .ZN(n6672) );
  NAND2_X1 U8269 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3084), .ZN(n7371) );
  OAI21_X1 U8270 ( .B1(n9027), .B2(n6672), .A(n7371), .ZN(n6679) );
  NAND2_X1 U8271 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n6914), .ZN(n6675) );
  OAI21_X1 U8272 ( .B1(n6914), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6675), .ZN(
        n6676) );
  AOI211_X1 U8273 ( .C1(n6677), .C2(n6676), .A(n6913), .B(n9490), .ZN(n6678)
         );
  AOI211_X1 U8274 ( .C1(n9497), .C2(n6680), .A(n6679), .B(n6678), .ZN(n6681)
         );
  OAI21_X1 U8275 ( .B1(n9038), .B2(n6682), .A(n6681), .ZN(P1_U3254) );
  NAND2_X1 U8276 ( .A1(n6683), .A2(n6684), .ZN(n6714) );
  OAI21_X1 U8277 ( .B1(n6684), .B2(n6683), .A(n6714), .ZN(n6685) );
  NAND2_X1 U8278 ( .A1(n6685), .A2(n8926), .ZN(n6690) );
  INV_X1 U8279 ( .A(n8940), .ZN(n8952) );
  AOI21_X1 U8280 ( .B1(n8973), .B2(n8928), .A(n6686), .ZN(n6687) );
  OAI21_X1 U8281 ( .B1(n6133), .B2(n8952), .A(n6687), .ZN(n6688) );
  AOI21_X1 U8282 ( .B1(n8957), .B2(n6988), .A(n6688), .ZN(n6689) );
  OAI211_X1 U8283 ( .C1(n6991), .C2(n8960), .A(n6690), .B(n6689), .ZN(P1_U3216) );
  XNOR2_X1 U8284 ( .A(n6692), .B(n6691), .ZN(n6696) );
  INV_X1 U8285 ( .A(n6981), .ZN(n9662) );
  NAND2_X1 U8286 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n7951) );
  OAI21_X1 U8287 ( .B1(n8422), .B2(n9662), .A(n7951), .ZN(n6694) );
  OAI22_X1 U8288 ( .A1(n8694), .A2(n8416), .B1(n8414), .B2(n6965), .ZN(n6693)
         );
  AOI211_X1 U8289 ( .C1(n6810), .C2(n8358), .A(n6694), .B(n6693), .ZN(n6695)
         );
  OAI21_X1 U8290 ( .B1(n6696), .B2(n8408), .A(n6695), .ZN(P2_U3223) );
  INV_X1 U8291 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6709) );
  OAI21_X1 U8292 ( .B1(n6698), .B2(n6699), .A(n6697), .ZN(n6993) );
  INV_X1 U8293 ( .A(n6993), .ZN(n6707) );
  OAI22_X1 U8294 ( .A1(n6133), .A2(n9378), .B1(n6950), .B2(n9376), .ZN(n6702)
         );
  XNOR2_X1 U8295 ( .A(n7747), .B(n6699), .ZN(n6700) );
  NOR2_X1 U8296 ( .A1(n6700), .A2(n9203), .ZN(n6701) );
  AOI211_X1 U8297 ( .C1(n6834), .C2(n6993), .A(n6702), .B(n6701), .ZN(n6995)
         );
  INV_X1 U8298 ( .A(n6940), .ZN(n6704) );
  INV_X1 U8299 ( .A(n6837), .ZN(n6703) );
  AOI21_X1 U8300 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(n6987) );
  AOI22_X1 U8301 ( .A1(n6987), .A2(n9423), .B1(n9520), .B2(n6705), .ZN(n6706)
         );
  OAI211_X1 U8302 ( .C1(n6707), .C2(n9335), .A(n6995), .B(n6706), .ZN(n6710)
         );
  NAND2_X1 U8303 ( .A1(n6710), .A2(n9550), .ZN(n6708) );
  OAI21_X1 U8304 ( .B1(n9550), .B2(n6709), .A(n6708), .ZN(P1_U3463) );
  NAND2_X1 U8305 ( .A1(n6710), .A2(n9562), .ZN(n6711) );
  OAI21_X1 U8306 ( .B1(n9562), .B2(n6272), .A(n6711), .ZN(P1_U3526) );
  AND2_X1 U8307 ( .A1(n6714), .A2(n6712), .ZN(n6717) );
  NAND2_X1 U8308 ( .A1(n6714), .A2(n6713), .ZN(n6715) );
  OAI211_X1 U8309 ( .C1(n6717), .C2(n6716), .A(n8926), .B(n6715), .ZN(n6722)
         );
  AOI21_X1 U8310 ( .B1(n6136), .B2(n8928), .A(n6718), .ZN(n6719) );
  OAI21_X1 U8311 ( .B1(n6832), .B2(n8952), .A(n6719), .ZN(n6720) );
  AOI21_X1 U8312 ( .B1(n8957), .B2(n6839), .A(n6720), .ZN(n6721) );
  OAI211_X1 U8313 ( .C1(n9511), .C2(n8960), .A(n6722), .B(n6721), .ZN(P1_U3228) );
  INV_X1 U8314 ( .A(n6723), .ZN(n6725) );
  OAI222_X1 U8315 ( .A1(P1_U3084), .A2(n7777), .B1(n8334), .B2(n6725), .C1(
        n6724), .C2(n8333), .ZN(P1_U3333) );
  OAI222_X1 U8316 ( .A1(n8856), .A2(n6726), .B1(P2_U3152), .B2(n8282), .C1(
        n8098), .C2(n6725), .ZN(P2_U3338) );
  XOR2_X1 U8317 ( .A(n6728), .B(n6727), .Z(n6729) );
  XNOR2_X1 U8318 ( .A(n6730), .B(n6729), .ZN(n6736) );
  NAND2_X1 U8319 ( .A1(n8957), .A2(n6873), .ZN(n6733) );
  AOI21_X1 U8320 ( .B1(n8970), .B2(n8928), .A(n6731), .ZN(n6732) );
  OAI211_X1 U8321 ( .C1(n6949), .C2(n8952), .A(n6733), .B(n6732), .ZN(n6734)
         );
  AOI21_X1 U8322 ( .B1(n8914), .B2(n6768), .A(n6734), .ZN(n6735) );
  OAI21_X1 U8323 ( .B1(n6736), .B2(n8947), .A(n6735), .ZN(P1_U3211) );
  OAI22_X1 U8324 ( .A1(n6738), .A2(n9211), .B1(n9209), .B2(n6737), .ZN(n6739)
         );
  OAI21_X1 U8325 ( .B1(n6740), .B2(n6739), .A(n7027), .ZN(n6742) );
  AOI22_X1 U8326 ( .A1(n9415), .A2(n7831), .B1(n9430), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6741) );
  OAI211_X1 U8327 ( .C1(n6743), .C2(n7491), .A(n6742), .B(n6741), .ZN(P1_U3290) );
  OAI21_X1 U8328 ( .B1(n6746), .B2(n6745), .A(n6744), .ZN(n6750) );
  INV_X1 U8329 ( .A(n7056), .ZN(n9668) );
  OAI22_X1 U8330 ( .A1(n9668), .A2(n8422), .B1(n8416), .B2(n6966), .ZN(n6749)
         );
  NAND2_X1 U8331 ( .A1(n8358), .A2(n7055), .ZN(n6747) );
  NAND2_X1 U8332 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7939) );
  OAI211_X1 U8333 ( .C1(n6980), .C2(n8414), .A(n6747), .B(n7939), .ZN(n6748)
         );
  AOI211_X1 U8334 ( .C1(n6750), .C2(n8410), .A(n6749), .B(n6748), .ZN(n6751)
         );
  INV_X1 U8335 ( .A(n6751), .ZN(P2_U3233) );
  INV_X1 U8336 ( .A(n6752), .ZN(n6754) );
  OAI222_X1 U8337 ( .A1(P1_U3084), .A2(n7823), .B1(n8334), .B2(n6754), .C1(
        n6753), .C2(n8333), .ZN(P1_U3332) );
  OAI222_X1 U8338 ( .A1(n8856), .A2(n6755), .B1(P2_U3152), .B2(n8114), .C1(
        n8098), .C2(n6754), .ZN(P2_U3337) );
  INV_X1 U8339 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6771) );
  AND2_X1 U8340 ( .A1(n6949), .A2(n9527), .ZN(n6847) );
  OR2_X1 U8341 ( .A1(n7797), .A2(n6847), .ZN(n6846) );
  OR2_X1 U8342 ( .A1(n6998), .A2(n6846), .ZN(n6759) );
  AND2_X1 U8343 ( .A1(n6137), .A2(n6756), .ZN(n6849) );
  OR2_X1 U8344 ( .A1(n6847), .A2(n6849), .ZN(n6757) );
  AND2_X1 U8345 ( .A1(n6759), .A2(n6757), .ZN(n6761) );
  NAND2_X1 U8346 ( .A1(n6906), .A2(n6768), .ZN(n7611) );
  INV_X1 U8347 ( .A(n6906), .ZN(n8971) );
  NAND2_X1 U8348 ( .A1(n8971), .A2(n6875), .ZN(n7845) );
  NAND2_X1 U8349 ( .A1(n7611), .A2(n7845), .ZN(n6850) );
  AND2_X1 U8350 ( .A1(n6850), .A2(n6757), .ZN(n6758) );
  NAND2_X1 U8351 ( .A1(n6759), .A2(n6758), .ZN(n6760) );
  OAI21_X1 U8352 ( .B1(n6761), .B2(n6850), .A(n6760), .ZN(n6762) );
  INV_X1 U8353 ( .A(n6762), .ZN(n6881) );
  NAND2_X1 U8354 ( .A1(n9382), .A2(n9335), .ZN(n9546) );
  INV_X1 U8355 ( .A(n9546), .ZN(n9517) );
  INV_X1 U8356 ( .A(n6850), .ZN(n7802) );
  NAND2_X1 U8357 ( .A1(n7741), .A2(n7596), .ZN(n7600) );
  INV_X1 U8358 ( .A(n7610), .ZN(n7744) );
  NOR2_X1 U8359 ( .A1(n7600), .A2(n7744), .ZN(n7842) );
  NAND2_X1 U8360 ( .A1(n7604), .A2(n7608), .ZN(n6763) );
  AND2_X1 U8361 ( .A1(n7610), .A2(n6763), .ZN(n7841) );
  AOI21_X1 U8362 ( .B1(n7599), .B2(n7842), .A(n7841), .ZN(n6764) );
  NAND2_X1 U8363 ( .A1(n6764), .A2(n7802), .ZN(n6858) );
  OAI21_X1 U8364 ( .B1(n7802), .B2(n6764), .A(n6858), .ZN(n6765) );
  AOI222_X1 U8365 ( .A1(n9412), .A2(n6765), .B1(n8970), .B2(n9407), .C1(n8972), 
        .C2(n9409), .ZN(n6876) );
  NAND2_X1 U8366 ( .A1(n6766), .A2(n6875), .ZN(n6863) );
  AOI211_X1 U8367 ( .C1(n6768), .C2(n6767), .A(n9542), .B(n4417), .ZN(n6879)
         );
  AOI21_X1 U8368 ( .B1(n9520), .B2(n6768), .A(n6879), .ZN(n6769) );
  OAI211_X1 U8369 ( .C1(n6881), .C2(n9517), .A(n6876), .B(n6769), .ZN(n6772)
         );
  NAND2_X1 U8370 ( .A1(n6772), .A2(n9562), .ZN(n6770) );
  OAI21_X1 U8371 ( .B1(n9562), .B2(n6771), .A(n6770), .ZN(P1_U3530) );
  INV_X1 U8372 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U8373 ( .A1(n6772), .A2(n9550), .ZN(n6773) );
  OAI21_X1 U8374 ( .B1(n9550), .B2(n6774), .A(n6773), .ZN(P1_U3475) );
  INV_X1 U8375 ( .A(n6788), .ZN(n8436) );
  NAND2_X1 U8376 ( .A1(n6788), .A2(n9649), .ZN(n8160) );
  INV_X1 U8377 ( .A(n6776), .ZN(n6777) );
  NAND2_X1 U8378 ( .A1(n8694), .A2(n6782), .ZN(n8164) );
  INV_X1 U8379 ( .A(n8694), .ZN(n8435) );
  NAND2_X1 U8380 ( .A1(n9657), .A2(n8435), .ZN(n8165) );
  INV_X1 U8381 ( .A(n8159), .ZN(n8291) );
  OAI21_X1 U8382 ( .B1(n6777), .B2(n8291), .A(n6799), .ZN(n9660) );
  AND2_X1 U8383 ( .A1(n6779), .A2(n6778), .ZN(n8701) );
  NAND2_X1 U8384 ( .A1(n8701), .A2(n8700), .ZN(n8703) );
  INV_X1 U8385 ( .A(n8703), .ZN(n6780) );
  OAI211_X1 U8386 ( .C1(n6780), .C2(n9657), .A(n9650), .B(n6982), .ZN(n9656)
         );
  AOI22_X1 U8387 ( .A1(n9577), .A2(n6782), .B1(n9576), .B2(n6781), .ZN(n6783)
         );
  OAI21_X1 U8388 ( .B1(n9656), .B2(n9583), .A(n6783), .ZN(n6790) );
  NOR2_X1 U8389 ( .A1(n8159), .A2(n4335), .ZN(n6786) );
  AND2_X1 U8390 ( .A1(n6784), .A2(n8151), .ZN(n8687) );
  AOI21_X1 U8391 ( .B1(n6786), .B2(n8691), .A(n6802), .ZN(n6787) );
  OAI222_X1 U8392 ( .A1(n8693), .A2(n6966), .B1(n8695), .B2(n6788), .C1(n8643), 
        .C2(n6787), .ZN(n9658) );
  MUX2_X1 U8393 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9658), .S(n8699), .Z(n6789)
         );
  AOI211_X1 U8394 ( .C1(n8711), .C2(n9660), .A(n6790), .B(n6789), .ZN(n6791)
         );
  INV_X1 U8395 ( .A(n6791), .ZN(P2_U3289) );
  OAI21_X1 U8396 ( .B1(n6793), .B2(n9209), .A(n6792), .ZN(n6794) );
  NAND2_X1 U8397 ( .A1(n6794), .A2(n7027), .ZN(n6797) );
  INV_X1 U8398 ( .A(n9088), .ZN(n9229) );
  OAI21_X1 U8399 ( .B1(n9229), .B2(n9415), .A(n6795), .ZN(n6796) );
  OAI211_X1 U8400 ( .C1(n6259), .C2(n7027), .A(n6797), .B(n6796), .ZN(P1_U3291) );
  NAND2_X1 U8401 ( .A1(n8694), .A2(n9657), .ZN(n6798) );
  OR2_X1 U8402 ( .A1(n6981), .A2(n6966), .ZN(n8170) );
  NAND2_X1 U8403 ( .A1(n6981), .A2(n6966), .ZN(n8169) );
  OR2_X1 U8404 ( .A1(n6969), .A2(n8294), .ZN(n7046) );
  NAND2_X1 U8405 ( .A1(n6969), .A2(n8294), .ZN(n6800) );
  NAND2_X1 U8406 ( .A1(n7046), .A2(n6800), .ZN(n6807) );
  INV_X1 U8407 ( .A(n6965), .ZN(n8433) );
  AOI22_X1 U8408 ( .A1(n8678), .A2(n8435), .B1(n8433), .B2(n8680), .ZN(n6806)
         );
  INV_X1 U8409 ( .A(n8164), .ZN(n6801) );
  INV_X1 U8410 ( .A(n6977), .ZN(n6804) );
  NOR3_X1 U8411 ( .A1(n6802), .A2(n8294), .A3(n6801), .ZN(n6803) );
  OAI21_X1 U8412 ( .B1(n6804), .B2(n6803), .A(n8492), .ZN(n6805) );
  OAI211_X1 U8413 ( .C1(n6807), .C2(n9571), .A(n6806), .B(n6805), .ZN(n9664)
         );
  INV_X1 U8414 ( .A(n9664), .ZN(n6815) );
  INV_X1 U8415 ( .A(n6807), .ZN(n9666) );
  INV_X1 U8416 ( .A(n6808), .ZN(n6809) );
  NAND2_X1 U8417 ( .A1(n8699), .A2(n6809), .ZN(n9584) );
  INV_X1 U8418 ( .A(n9584), .ZN(n8722) );
  XNOR2_X1 U8419 ( .A(n6982), .B(n6981), .ZN(n9663) );
  AOI22_X1 U8420 ( .A1(n9588), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n6810), .B2(
        n9576), .ZN(n6812) );
  NAND2_X1 U8421 ( .A1(n9577), .A2(n6981), .ZN(n6811) );
  OAI211_X1 U8422 ( .C1(n9663), .C2(n8707), .A(n6812), .B(n6811), .ZN(n6813)
         );
  AOI21_X1 U8423 ( .B1(n9666), .B2(n8722), .A(n6813), .ZN(n6814) );
  OAI21_X1 U8424 ( .B1(n6815), .B2(n9588), .A(n6814), .ZN(P2_U3288) );
  NAND2_X1 U8425 ( .A1(n4314), .A2(n6818), .ZN(n6883) );
  OAI21_X1 U8426 ( .B1(n4314), .B2(n6818), .A(n6883), .ZN(n6819) );
  NOR2_X1 U8427 ( .A1(n6819), .A2(n6820), .ZN(n6887) );
  AOI21_X1 U8428 ( .B1(n6820), .B2(n6819), .A(n6887), .ZN(n6825) );
  NAND2_X1 U8429 ( .A1(n8957), .A2(n6958), .ZN(n6822) );
  INV_X1 U8430 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9801) );
  NOR2_X1 U8431 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9801), .ZN(n9456) );
  AOI21_X1 U8432 ( .B1(n8972), .B2(n8928), .A(n9456), .ZN(n6821) );
  OAI211_X1 U8433 ( .C1(n6950), .C2(n8952), .A(n6822), .B(n6821), .ZN(n6823)
         );
  AOI21_X1 U8434 ( .B1(n8914), .B2(n9519), .A(n6823), .ZN(n6824) );
  OAI21_X1 U8435 ( .B1(n6825), .B2(n8947), .A(n6824), .ZN(P1_U3225) );
  INV_X1 U8436 ( .A(n6826), .ZN(n8097) );
  OAI222_X1 U8437 ( .A1(n8333), .A2(n6828), .B1(n8334), .B2(n8097), .C1(
        P1_U3084), .C2(n6827), .ZN(P1_U3331) );
  XNOR2_X1 U8438 ( .A(n7598), .B(n7792), .ZN(n6836) );
  OAI21_X1 U8439 ( .B1(n6830), .B2(n7792), .A(n6829), .ZN(n9515) );
  OAI22_X1 U8440 ( .A1(n6832), .A2(n9378), .B1(n6831), .B2(n9376), .ZN(n6833)
         );
  AOI21_X1 U8441 ( .B1(n9515), .B2(n6834), .A(n6833), .ZN(n6835) );
  OAI21_X1 U8442 ( .B1(n9203), .B2(n6836), .A(n6835), .ZN(n9513) );
  INV_X1 U8443 ( .A(n9513), .ZN(n6845) );
  INV_X1 U8444 ( .A(n7491), .ZN(n9394) );
  NAND2_X1 U8445 ( .A1(n6837), .A2(n6840), .ZN(n6838) );
  NAND2_X1 U8446 ( .A1(n6955), .A2(n6838), .ZN(n9512) );
  INV_X1 U8447 ( .A(n9209), .ZN(n9414) );
  AOI22_X1 U8448 ( .A1(n9386), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n6839), .B2(
        n9414), .ZN(n6842) );
  NAND2_X1 U8449 ( .A1(n9415), .A2(n6840), .ZN(n6841) );
  OAI211_X1 U8450 ( .C1(n9088), .C2(n9512), .A(n6842), .B(n6841), .ZN(n6843)
         );
  AOI21_X1 U8451 ( .B1(n9515), .B2(n9394), .A(n6843), .ZN(n6844) );
  OAI21_X1 U8452 ( .B1(n6845), .B2(n9386), .A(n6844), .ZN(P1_U3287) );
  AND2_X1 U8453 ( .A1(n6906), .A2(n6875), .ZN(n6851) );
  OR2_X1 U8454 ( .A1(n6846), .A2(n6851), .ZN(n6996) );
  OR2_X1 U8455 ( .A1(n6998), .A2(n6996), .ZN(n6854) );
  OR2_X1 U8456 ( .A1(n6847), .A2(n6851), .ZN(n6848) );
  OR2_X1 U8457 ( .A1(n6849), .A2(n6848), .ZN(n6853) );
  OR2_X1 U8458 ( .A1(n6851), .A2(n6850), .ZN(n6852) );
  AND2_X1 U8459 ( .A1(n6853), .A2(n6852), .ZN(n7000) );
  AND2_X1 U8460 ( .A1(n6854), .A2(n7000), .ZN(n6855) );
  NAND2_X1 U8461 ( .A1(n7073), .A2(n6999), .ZN(n7619) );
  OR2_X1 U8462 ( .A1(n6855), .A2(n7803), .ZN(n6857) );
  NAND2_X1 U8463 ( .A1(n6855), .A2(n7803), .ZN(n6856) );
  NAND2_X1 U8464 ( .A1(n6857), .A2(n6856), .ZN(n6862) );
  AOI22_X1 U8465 ( .A1(n8971), .A2(n9409), .B1(n9407), .B2(n8969), .ZN(n6861)
         );
  AND2_X1 U8466 ( .A1(n6858), .A2(n7611), .ZN(n6859) );
  OAI211_X1 U8467 ( .C1(n6859), .C2(n7803), .A(n9374), .B(n9412), .ZN(n6860)
         );
  OAI211_X1 U8468 ( .C1(n6862), .C2(n9382), .A(n6861), .B(n6860), .ZN(n9535)
         );
  INV_X1 U8469 ( .A(n9535), .ZN(n6869) );
  INV_X1 U8470 ( .A(n6862), .ZN(n9537) );
  NAND2_X1 U8471 ( .A1(n6863), .A2(n6999), .ZN(n6864) );
  NAND2_X1 U8472 ( .A1(n7003), .A2(n6864), .ZN(n9534) );
  AOI22_X1 U8473 ( .A1(n9386), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n6902), .B2(
        n9414), .ZN(n6866) );
  NAND2_X1 U8474 ( .A1(n9415), .A2(n6999), .ZN(n6865) );
  OAI211_X1 U8475 ( .C1(n9534), .C2(n9088), .A(n6866), .B(n6865), .ZN(n6867)
         );
  AOI21_X1 U8476 ( .B1(n9537), .B2(n9394), .A(n6867), .ZN(n6868) );
  OAI21_X1 U8477 ( .B1(n6869), .B2(n9386), .A(n6868), .ZN(P1_U3283) );
  NAND2_X1 U8478 ( .A1(n6871), .A2(n6870), .ZN(n6872) );
  AOI22_X1 U8479 ( .A1(n9386), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6873), .B2(
        n9414), .ZN(n6874) );
  OAI21_X1 U8480 ( .B1(n9237), .B2(n6875), .A(n6874), .ZN(n6878) );
  NOR2_X1 U8481 ( .A1(n6876), .A2(n9386), .ZN(n6877) );
  AOI211_X1 U8482 ( .C1(n6879), .C2(n9426), .A(n6878), .B(n6877), .ZN(n6880)
         );
  OAI21_X1 U8483 ( .B1(n6881), .B2(n9247), .A(n6880), .ZN(P1_U3284) );
  INV_X1 U8484 ( .A(n6882), .ZN(n6890) );
  INV_X1 U8485 ( .A(n6883), .ZN(n6886) );
  INV_X1 U8486 ( .A(n6884), .ZN(n6885) );
  OAI22_X1 U8487 ( .A1(n6887), .A2(n6886), .B1(n6890), .B2(n6885), .ZN(n6888)
         );
  OAI211_X1 U8488 ( .C1(n6890), .C2(n6889), .A(n6888), .B(n8926), .ZN(n6897)
         );
  NAND2_X1 U8489 ( .A1(n6136), .A2(n8940), .ZN(n6893) );
  INV_X1 U8490 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6891) );
  NOR2_X1 U8491 ( .A1(n6891), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9468) );
  INV_X1 U8492 ( .A(n9468), .ZN(n6892) );
  OAI211_X1 U8493 ( .C1(n6906), .C2(n8954), .A(n6893), .B(n6892), .ZN(n6894)
         );
  AOI21_X1 U8494 ( .B1(n8957), .B2(n6895), .A(n6894), .ZN(n6896) );
  OAI211_X1 U8495 ( .C1(n9527), .C2(n8960), .A(n6897), .B(n6896), .ZN(P1_U3237) );
  XOR2_X1 U8496 ( .A(n6900), .B(n6899), .Z(n6901) );
  XNOR2_X1 U8497 ( .A(n6898), .B(n6901), .ZN(n6909) );
  NAND2_X1 U8498 ( .A1(n8957), .A2(n6902), .ZN(n6905) );
  INV_X1 U8499 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6903) );
  NOR2_X1 U8500 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6903), .ZN(n9481) );
  AOI21_X1 U8501 ( .B1(n8928), .B2(n8969), .A(n9481), .ZN(n6904) );
  OAI211_X1 U8502 ( .C1(n6906), .C2(n8952), .A(n6905), .B(n6904), .ZN(n6907)
         );
  AOI21_X1 U8503 ( .B1(n8914), .B2(n6999), .A(n6907), .ZN(n6908) );
  OAI21_X1 U8504 ( .B1(n6909), .B2(n8947), .A(n6908), .ZN(P1_U3219) );
  INV_X1 U8505 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n6921) );
  XNOR2_X1 U8506 ( .A(n7172), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n6912) );
  OAI21_X1 U8507 ( .B1(n6914), .B2(P1_REG1_REG_13__SCAN_IN), .A(n6910), .ZN(
        n6911) );
  NAND2_X1 U8508 ( .A1(n6912), .A2(n6911), .ZN(n7165) );
  OAI21_X1 U8509 ( .B1(n6912), .B2(n6911), .A(n7165), .ZN(n6919) );
  NAND2_X1 U8510 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7460) );
  OAI21_X1 U8511 ( .B1(n9027), .B2(n7172), .A(n7460), .ZN(n6918) );
  INV_X1 U8512 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6915) );
  NOR2_X1 U8513 ( .A1(n6915), .A2(n6916), .ZN(n7174) );
  AOI211_X1 U8514 ( .C1(n6916), .C2(n6915), .A(n7174), .B(n9490), .ZN(n6917)
         );
  AOI211_X1 U8515 ( .C1(n9497), .C2(n6919), .A(n6918), .B(n6917), .ZN(n6920)
         );
  OAI21_X1 U8516 ( .B1(n9038), .B2(n6921), .A(n6920), .ZN(P1_U3255) );
  INV_X1 U8517 ( .A(n9676), .ZN(n9578) );
  XOR2_X1 U8518 ( .A(n6923), .B(n6922), .Z(n6924) );
  NAND2_X1 U8519 ( .A1(n6924), .A2(n8410), .ZN(n6930) );
  OR2_X1 U8520 ( .A1(n7118), .A2(n8693), .ZN(n6926) );
  OR2_X1 U8521 ( .A1(n6965), .A2(n8695), .ZN(n6925) );
  NAND2_X1 U8522 ( .A1(n6926), .A2(n6925), .ZN(n9573) );
  INV_X1 U8523 ( .A(n9573), .ZN(n6927) );
  OAI22_X1 U8524 ( .A1(n8396), .A2(n6927), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7931), .ZN(n6928) );
  AOI21_X1 U8525 ( .B1(n9575), .B2(n8358), .A(n6928), .ZN(n6929) );
  OAI211_X1 U8526 ( .C1(n9578), .C2(n8422), .A(n6930), .B(n6929), .ZN(P2_U3219) );
  XNOR2_X1 U8527 ( .A(n7828), .B(n7793), .ZN(n6931) );
  NAND2_X1 U8528 ( .A1(n6931), .A2(n9412), .ZN(n6933) );
  AOI22_X1 U8529 ( .A1(n8974), .A2(n9407), .B1(n9409), .B2(n8976), .ZN(n6932)
         );
  NAND2_X1 U8530 ( .A1(n6933), .A2(n6932), .ZN(n9507) );
  INV_X1 U8531 ( .A(n9507), .ZN(n6946) );
  OAI21_X1 U8532 ( .B1(n6936), .B2(n6935), .A(n6934), .ZN(n9509) );
  INV_X1 U8533 ( .A(n9247), .ZN(n9427) );
  NOR2_X1 U8534 ( .A1(n6938), .A2(n6937), .ZN(n6939) );
  OR2_X1 U8535 ( .A1(n6940), .A2(n6939), .ZN(n9506) );
  AOI22_X1 U8536 ( .A1(n9430), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9414), .ZN(n6943) );
  NAND2_X1 U8537 ( .A1(n9415), .A2(n6941), .ZN(n6942) );
  OAI211_X1 U8538 ( .C1(n9088), .C2(n9506), .A(n6943), .B(n6942), .ZN(n6944)
         );
  AOI21_X1 U8539 ( .B1(n9509), .B2(n9427), .A(n6944), .ZN(n6945) );
  OAI21_X1 U8540 ( .B1(n6946), .B2(n9386), .A(n6945), .ZN(P1_U3289) );
  OAI21_X1 U8541 ( .B1(n7797), .B2(n6948), .A(n6947), .ZN(n6952) );
  OAI22_X1 U8542 ( .A1(n6950), .A2(n9378), .B1(n6949), .B2(n9376), .ZN(n6951)
         );
  AOI21_X1 U8543 ( .B1(n6952), .B2(n9412), .A(n6951), .ZN(n9525) );
  NAND2_X1 U8544 ( .A1(n6998), .A2(n7797), .ZN(n6953) );
  NAND2_X1 U8545 ( .A1(n6954), .A2(n6953), .ZN(n9518) );
  INV_X1 U8546 ( .A(n9518), .ZN(n6963) );
  AOI21_X1 U8547 ( .B1(n6955), .B2(n9519), .A(n9542), .ZN(n6957) );
  NAND2_X1 U8548 ( .A1(n6957), .A2(n6956), .ZN(n9522) );
  AOI22_X1 U8549 ( .A1(n9430), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6958), .B2(
        n9414), .ZN(n6960) );
  NAND2_X1 U8550 ( .A1(n9415), .A2(n9519), .ZN(n6959) );
  OAI211_X1 U8551 ( .C1(n9522), .C2(n6961), .A(n6960), .B(n6959), .ZN(n6962)
         );
  AOI21_X1 U8552 ( .B1(n6963), .B2(n9427), .A(n6962), .ZN(n6964) );
  OAI21_X1 U8553 ( .B1(n9430), .B2(n9525), .A(n6964), .ZN(P1_U3286) );
  OR2_X1 U8554 ( .A1(n8294), .A2(n4784), .ZN(n6968) );
  OR2_X1 U8555 ( .A1(n6969), .A2(n6968), .ZN(n6967) );
  OR2_X1 U8556 ( .A1(n7056), .A2(n6965), .ZN(n9563) );
  NAND2_X1 U8557 ( .A1(n7056), .A2(n6965), .ZN(n8179) );
  NAND2_X1 U8558 ( .A1(n9563), .A2(n8179), .ZN(n8293) );
  INV_X1 U8559 ( .A(n6966), .ZN(n8434) );
  NAND2_X1 U8560 ( .A1(n6981), .A2(n8434), .ZN(n7044) );
  AND2_X1 U8561 ( .A1(n8293), .A2(n7044), .ZN(n7045) );
  OR2_X1 U8562 ( .A1(n4784), .A2(n7045), .ZN(n6970) );
  AND2_X1 U8563 ( .A1(n6967), .A2(n6970), .ZN(n9568) );
  OR2_X1 U8564 ( .A1(n9676), .A2(n6980), .ZN(n6978) );
  NAND2_X1 U8565 ( .A1(n9676), .A2(n6980), .ZN(n8181) );
  INV_X1 U8566 ( .A(n6980), .ZN(n8432) );
  NAND2_X1 U8567 ( .A1(n9676), .A2(n8432), .ZN(n6973) );
  NAND2_X1 U8568 ( .A1(n9570), .A2(n6973), .ZN(n6976) );
  OR2_X1 U8569 ( .A1(n7084), .A2(n7118), .ZN(n8187) );
  NAND2_X1 U8570 ( .A1(n7084), .A2(n7118), .ZN(n8185) );
  NAND2_X1 U8571 ( .A1(n8187), .A2(n8185), .ZN(n8297) );
  INV_X1 U8572 ( .A(n8297), .ZN(n6974) );
  OR2_X1 U8573 ( .A1(n6971), .A2(n6970), .ZN(n6972) );
  OR2_X1 U8574 ( .A1(n6974), .A2(n6973), .ZN(n7086) );
  AND2_X1 U8575 ( .A1(n7090), .A2(n7086), .ZN(n6975) );
  OAI21_X1 U8576 ( .B1(n6976), .B2(n8297), .A(n6975), .ZN(n9683) );
  INV_X1 U8577 ( .A(n8179), .ZN(n8173) );
  NAND2_X1 U8578 ( .A1(n6978), .A2(n9563), .ZN(n8178) );
  XNOR2_X1 U8579 ( .A(n7093), .B(n8297), .ZN(n6979) );
  OAI222_X1 U8580 ( .A1(n8693), .A2(n7087), .B1(n8695), .B2(n6980), .C1(n6979), 
        .C2(n8643), .ZN(n9686) );
  NOR2_X2 U8581 ( .A1(n7052), .A2(n7056), .ZN(n9579) );
  XNOR2_X1 U8582 ( .A(n9580), .B(n9684), .ZN(n9685) );
  AOI22_X1 U8583 ( .A1(n9588), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7036), .B2(
        n9576), .ZN(n6984) );
  NAND2_X1 U8584 ( .A1(n9577), .A2(n7084), .ZN(n6983) );
  OAI211_X1 U8585 ( .C1(n9685), .C2(n8707), .A(n6984), .B(n6983), .ZN(n6985)
         );
  AOI21_X1 U8586 ( .B1(n9686), .B2(n8699), .A(n6985), .ZN(n6986) );
  OAI21_X1 U8587 ( .B1(n8686), .B2(n9683), .A(n6986), .ZN(P2_U3285) );
  NAND2_X1 U8588 ( .A1(n6987), .A2(n9229), .ZN(n6990) );
  AOI22_X1 U8589 ( .A1(n9430), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9414), .B2(
        n6988), .ZN(n6989) );
  OAI211_X1 U8590 ( .C1(n6991), .C2(n9237), .A(n6990), .B(n6989), .ZN(n6992)
         );
  AOI21_X1 U8591 ( .B1(n6993), .B2(n9394), .A(n6992), .ZN(n6994) );
  OAI21_X1 U8592 ( .B1(n6995), .B2(n9386), .A(n6994), .ZN(P1_U3288) );
  INV_X1 U8593 ( .A(n7075), .ZN(n9541) );
  NAND2_X1 U8594 ( .A1(n9541), .A2(n8969), .ZN(n7616) );
  INV_X1 U8595 ( .A(n8969), .ZN(n9379) );
  NAND2_X1 U8596 ( .A1(n9379), .A2(n7075), .ZN(n9371) );
  NAND2_X1 U8597 ( .A1(n7616), .A2(n9371), .ZN(n7805) );
  NAND2_X1 U8598 ( .A1(n8970), .A2(n6999), .ZN(n7001) );
  XOR2_X1 U8599 ( .A(n7805), .B(n7016), .Z(n9547) );
  INV_X1 U8600 ( .A(n9547), .ZN(n7009) );
  XOR2_X1 U8601 ( .A(n7805), .B(n7022), .Z(n7002) );
  OAI222_X1 U8602 ( .A1(n9378), .A2(n7073), .B1(n9376), .B2(n7023), .C1(n9203), 
        .C2(n7002), .ZN(n9544) );
  INV_X1 U8603 ( .A(n9392), .ZN(n7004) );
  OAI21_X1 U8604 ( .B1(n9541), .B2(n4422), .A(n7004), .ZN(n9543) );
  AOI22_X1 U8605 ( .A1(n9430), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7070), .B2(
        n9414), .ZN(n7006) );
  NAND2_X1 U8606 ( .A1(n9415), .A2(n7075), .ZN(n7005) );
  OAI211_X1 U8607 ( .C1(n9543), .C2(n9088), .A(n7006), .B(n7005), .ZN(n7007)
         );
  AOI21_X1 U8608 ( .B1(n9544), .B2(n7027), .A(n7007), .ZN(n7008) );
  OAI21_X1 U8609 ( .B1(n7009), .B2(n9247), .A(n7008), .ZN(P1_U3282) );
  INV_X1 U8610 ( .A(n7010), .ZN(n7014) );
  NAND2_X1 U8611 ( .A1(n9366), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7012) );
  NAND2_X1 U8612 ( .A1(n7011), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7877) );
  OAI211_X1 U8613 ( .C1(n7014), .C2(n8334), .A(n7012), .B(n7877), .ZN(P1_U3330) );
  NAND2_X1 U8614 ( .A1(n8851), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7013) );
  OAI211_X1 U8615 ( .C1(n7014), .C2(n8858), .A(n7013), .B(n8328), .ZN(P2_U3335) );
  AND2_X1 U8616 ( .A1(n7075), .A2(n8969), .ZN(n7015) );
  OR2_X1 U8617 ( .A1(n9388), .A2(n7023), .ZN(n7617) );
  NAND2_X1 U8618 ( .A1(n9388), .A2(n7023), .ZN(n7623) );
  NAND2_X1 U8619 ( .A1(n7617), .A2(n7623), .ZN(n9380) );
  NAND2_X1 U8620 ( .A1(n9381), .A2(n9380), .ZN(n7018) );
  INV_X1 U8621 ( .A(n7023), .ZN(n8968) );
  OR2_X1 U8622 ( .A1(n9388), .A2(n8968), .ZN(n7017) );
  NAND2_X1 U8623 ( .A1(n7018), .A2(n7017), .ZN(n7019) );
  OR2_X1 U8624 ( .A1(n7204), .A2(n9377), .ZN(n7633) );
  NAND2_X1 U8625 ( .A1(n7204), .A2(n9377), .ZN(n7750) );
  NAND2_X1 U8626 ( .A1(n7019), .A2(n7628), .ZN(n7020) );
  NAND2_X1 U8627 ( .A1(n7206), .A2(n7020), .ZN(n9437) );
  NAND2_X1 U8628 ( .A1(n7617), .A2(n7616), .ZN(n7624) );
  NAND2_X1 U8629 ( .A1(n7623), .A2(n9371), .ZN(n7021) );
  NAND2_X1 U8630 ( .A1(n7021), .A2(n7617), .ZN(n7749) );
  XNOR2_X1 U8631 ( .A(n7208), .B(n7628), .ZN(n7025) );
  OAI22_X1 U8632 ( .A1(n7023), .A2(n9378), .B1(n7210), .B2(n9376), .ZN(n7024)
         );
  AOI21_X1 U8633 ( .B1(n7025), .B2(n9412), .A(n7024), .ZN(n7026) );
  OAI21_X1 U8634 ( .B1(n9437), .B2(n9382), .A(n7026), .ZN(n9440) );
  NAND2_X1 U8635 ( .A1(n9440), .A2(n7027), .ZN(n7033) );
  INV_X1 U8636 ( .A(n9388), .ZN(n9398) );
  INV_X1 U8637 ( .A(n7204), .ZN(n9438) );
  OR2_X1 U8638 ( .A1(n9390), .A2(n9438), .ZN(n7028) );
  NAND2_X1 U8639 ( .A1(n9421), .A2(n7028), .ZN(n9439) );
  INV_X1 U8640 ( .A(n9439), .ZN(n7031) );
  AOI22_X1 U8641 ( .A1(n9386), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7186), .B2(
        n9414), .ZN(n7029) );
  OAI21_X1 U8642 ( .B1(n9438), .B2(n9237), .A(n7029), .ZN(n7030) );
  AOI21_X1 U8643 ( .B1(n7031), .B2(n9229), .A(n7030), .ZN(n7032) );
  OAI211_X1 U8644 ( .C1(n9437), .C2(n7491), .A(n7033), .B(n7032), .ZN(P1_U3280) );
  XOR2_X1 U8645 ( .A(n7035), .B(n7034), .Z(n7041) );
  AOI22_X1 U8646 ( .A1(n8375), .A2(n8432), .B1(n8358), .B2(n7036), .ZN(n7039)
         );
  OAI22_X1 U8647 ( .A1(n8414), .A2(n7087), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5102), .ZN(n7037) );
  INV_X1 U8648 ( .A(n7037), .ZN(n7038) );
  OAI211_X1 U8649 ( .C1(n9684), .C2(n8422), .A(n7039), .B(n7038), .ZN(n7040)
         );
  AOI21_X1 U8650 ( .B1(n7041), .B2(n8410), .A(n7040), .ZN(n7042) );
  INV_X1 U8651 ( .A(n7042), .ZN(P2_U3238) );
  XNOR2_X1 U8652 ( .A(n8293), .B(n7043), .ZN(n7051) );
  AND2_X1 U8653 ( .A1(n7046), .A2(n7044), .ZN(n7048) );
  NAND2_X1 U8654 ( .A1(n7046), .A2(n7045), .ZN(n7047) );
  OAI21_X1 U8655 ( .B1(n7048), .B2(n8293), .A(n7047), .ZN(n9672) );
  NAND2_X1 U8656 ( .A1(n9672), .A2(n7429), .ZN(n7050) );
  AOI22_X1 U8657 ( .A1(n8678), .A2(n8434), .B1(n8432), .B2(n8680), .ZN(n7049)
         );
  OAI211_X1 U8658 ( .C1(n8643), .C2(n7051), .A(n7050), .B(n7049), .ZN(n9670)
         );
  INV_X1 U8659 ( .A(n9670), .ZN(n7061) );
  INV_X1 U8660 ( .A(n9579), .ZN(n7054) );
  NAND2_X1 U8661 ( .A1(n7052), .A2(n7056), .ZN(n7053) );
  NAND2_X1 U8662 ( .A1(n7054), .A2(n7053), .ZN(n9669) );
  AOI22_X1 U8663 ( .A1(n9588), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7055), .B2(
        n9576), .ZN(n7058) );
  NAND2_X1 U8664 ( .A1(n9577), .A2(n7056), .ZN(n7057) );
  OAI211_X1 U8665 ( .C1(n9669), .C2(n8707), .A(n7058), .B(n7057), .ZN(n7059)
         );
  AOI21_X1 U8666 ( .B1(n9672), .B2(n8722), .A(n7059), .ZN(n7060) );
  OAI21_X1 U8667 ( .B1(n7061), .B2(n9588), .A(n7060), .ZN(P2_U3287) );
  INV_X1 U8668 ( .A(n7062), .ZN(n7066) );
  OAI222_X1 U8669 ( .A1(n7064), .A2(P2_U3152), .B1(n8098), .B2(n7066), .C1(
        n7063), .C2(n8856), .ZN(P2_U3334) );
  OAI222_X1 U8670 ( .A1(n7067), .A2(P1_U3084), .B1(n8334), .B2(n7066), .C1(
        n7065), .C2(n8333), .ZN(P1_U3329) );
  AOI21_X1 U8671 ( .B1(n7069), .B2(n7068), .A(n4316), .ZN(n7077) );
  NAND2_X1 U8672 ( .A1(n8957), .A2(n7070), .ZN(n7072) );
  AND2_X1 U8673 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9495) );
  AOI21_X1 U8674 ( .B1(n8968), .B2(n8928), .A(n9495), .ZN(n7071) );
  OAI211_X1 U8675 ( .C1(n7073), .C2(n8952), .A(n7072), .B(n7071), .ZN(n7074)
         );
  AOI21_X1 U8676 ( .B1(n8914), .B2(n7075), .A(n7074), .ZN(n7076) );
  OAI21_X1 U8677 ( .B1(n7077), .B2(n8947), .A(n7076), .ZN(P1_U3229) );
  XNOR2_X1 U8678 ( .A(n7079), .B(n7078), .ZN(n7083) );
  INV_X1 U8679 ( .A(n8428), .ZN(n8200) );
  INV_X1 U8680 ( .A(n7087), .ZN(n8430) );
  AOI22_X1 U8681 ( .A1(n8375), .A2(n8430), .B1(n8358), .B2(n7104), .ZN(n7080)
         );
  NAND2_X1 U8682 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7902) );
  OAI211_X1 U8683 ( .C1(n8200), .C2(n8414), .A(n7080), .B(n7902), .ZN(n7081)
         );
  AOI21_X1 U8684 ( .B1(n8820), .B2(n8406), .A(n7081), .ZN(n7082) );
  OAI21_X1 U8685 ( .B1(n7083), .B2(n8408), .A(n7082), .ZN(P2_U3236) );
  INV_X1 U8686 ( .A(n7118), .ZN(n8431) );
  NAND2_X1 U8687 ( .A1(n7084), .A2(n8431), .ZN(n7085) );
  AND2_X1 U8688 ( .A1(n7086), .A2(n7085), .ZN(n7088) );
  AND2_X1 U8689 ( .A1(n7090), .A2(n7088), .ZN(n7091) );
  OR2_X1 U8690 ( .A1(n7107), .A2(n7087), .ZN(n8188) );
  NAND2_X1 U8691 ( .A1(n7107), .A2(n7087), .ZN(n8189) );
  NAND2_X1 U8692 ( .A1(n8188), .A2(n8189), .ZN(n8299) );
  AND2_X1 U8693 ( .A1(n8299), .A2(n7088), .ZN(n7089) );
  NAND2_X1 U8694 ( .A1(n7090), .A2(n7089), .ZN(n7109) );
  OAI21_X1 U8695 ( .B1(n7091), .B2(n8299), .A(n7109), .ZN(n9696) );
  INV_X1 U8696 ( .A(n9696), .ZN(n7099) );
  INV_X1 U8697 ( .A(n8185), .ZN(n7092) );
  XOR2_X1 U8698 ( .A(n8299), .B(n7100), .Z(n7094) );
  OAI222_X1 U8699 ( .A1(n8693), .A2(n7302), .B1(n8695), .B2(n7118), .C1(n8643), 
        .C2(n7094), .ZN(n9694) );
  INV_X1 U8700 ( .A(n7107), .ZN(n9691) );
  OAI21_X1 U8701 ( .B1(n9691), .B2(n4317), .A(n4263), .ZN(n9693) );
  AOI22_X1 U8702 ( .A1(n9588), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7116), .B2(
        n9576), .ZN(n7096) );
  NAND2_X1 U8703 ( .A1(n9577), .A2(n7107), .ZN(n7095) );
  OAI211_X1 U8704 ( .C1(n9693), .C2(n8707), .A(n7096), .B(n7095), .ZN(n7097)
         );
  AOI21_X1 U8705 ( .B1(n9694), .B2(n8699), .A(n7097), .ZN(n7098) );
  OAI21_X1 U8706 ( .B1(n7099), .B2(n8686), .A(n7098), .ZN(P2_U3284) );
  OR2_X1 U8707 ( .A1(n8820), .A2(n7302), .ZN(n8197) );
  NAND2_X1 U8708 ( .A1(n8820), .A2(n7302), .ZN(n8196) );
  NAND2_X1 U8709 ( .A1(n8197), .A2(n8196), .ZN(n8300) );
  INV_X1 U8710 ( .A(n8300), .ZN(n8194) );
  OAI21_X1 U8711 ( .B1(n8194), .B2(n7101), .A(n7301), .ZN(n7102) );
  AOI222_X1 U8712 ( .A1(n8492), .A2(n7102), .B1(n8428), .B2(n8680), .C1(n8430), 
        .C2(n8678), .ZN(n8823) );
  INV_X1 U8713 ( .A(n8820), .ZN(n7295) );
  INV_X1 U8714 ( .A(n7298), .ZN(n7103) );
  AOI21_X1 U8715 ( .B1(n8820), .B2(n4263), .A(n7103), .ZN(n8821) );
  AOI22_X1 U8716 ( .A1(n9588), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7104), .B2(
        n9576), .ZN(n7105) );
  OAI21_X1 U8717 ( .B1(n7295), .B2(n8674), .A(n7105), .ZN(n7106) );
  AOI21_X1 U8718 ( .B1(n8821), .B2(n8719), .A(n7106), .ZN(n7112) );
  OR2_X1 U8719 ( .A1(n7107), .A2(n8430), .ZN(n7108) );
  AND2_X2 U8720 ( .A1(n7109), .A2(n7108), .ZN(n7110) );
  OR2_X1 U8721 ( .A1(n7110), .A2(n8300), .ZN(n8819) );
  NAND3_X1 U8722 ( .A1(n8819), .A2(n8711), .A3(n8818), .ZN(n7111) );
  OAI211_X1 U8723 ( .C1(n8823), .C2(n9588), .A(n7112), .B(n7111), .ZN(P2_U3283) );
  XOR2_X1 U8724 ( .A(n7114), .B(n7113), .Z(n7115) );
  NAND2_X1 U8725 ( .A1(n7115), .A2(n8410), .ZN(n7122) );
  NAND2_X1 U8726 ( .A1(n8358), .A2(n7116), .ZN(n7117) );
  OAI21_X1 U8727 ( .B1(n7118), .B2(n8416), .A(n7117), .ZN(n7120) );
  NAND2_X1 U8728 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7912) );
  OAI21_X1 U8729 ( .B1(n8414), .B2(n7302), .A(n7912), .ZN(n7119) );
  NOR2_X1 U8730 ( .A1(n7120), .A2(n7119), .ZN(n7121) );
  OAI211_X1 U8731 ( .C1(n9691), .C2(n8422), .A(n7122), .B(n7121), .ZN(P2_U3226) );
  NAND2_X1 U8732 ( .A1(n7124), .A2(n7123), .ZN(n7125) );
  XNOR2_X1 U8733 ( .A(n7126), .B(n7125), .ZN(n7133) );
  NAND2_X1 U8734 ( .A1(n8940), .A2(n8969), .ZN(n7129) );
  INV_X1 U8735 ( .A(n7127), .ZN(n7128) );
  OAI211_X1 U8736 ( .C1(n9377), .C2(n8954), .A(n7129), .B(n7128), .ZN(n7131)
         );
  NOR2_X1 U8737 ( .A1(n8960), .A2(n9398), .ZN(n7130) );
  AOI211_X1 U8738 ( .C1(n9387), .C2(n8957), .A(n7131), .B(n7130), .ZN(n7132)
         );
  OAI21_X1 U8739 ( .B1(n7133), .B2(n8947), .A(n7132), .ZN(P1_U3215) );
  INV_X1 U8740 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9908) );
  NOR2_X1 U8741 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7134) );
  AOI21_X1 U8742 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7134), .ZN(n9723) );
  NOR2_X1 U8743 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7135) );
  AOI21_X1 U8744 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7135), .ZN(n9726) );
  NOR2_X1 U8745 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7136) );
  AOI21_X1 U8746 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7136), .ZN(n9729) );
  NOR2_X1 U8747 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7137) );
  AOI21_X1 U8748 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7137), .ZN(n9732) );
  NOR2_X1 U8749 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7138) );
  AOI21_X1 U8750 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7138), .ZN(n9735) );
  NOR2_X1 U8751 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7145) );
  XNOR2_X1 U8752 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9919) );
  NAND2_X1 U8753 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7143) );
  XNOR2_X1 U8754 ( .A(n7139), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U8755 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7141) );
  XOR2_X1 U8756 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n9915) );
  AOI21_X1 U8757 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9716) );
  INV_X1 U8758 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9720) );
  NAND3_X1 U8759 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9718) );
  OAI21_X1 U8760 ( .B1(n9716), .B2(n9720), .A(n9718), .ZN(n9914) );
  NAND2_X1 U8761 ( .A1(n9915), .A2(n9914), .ZN(n7140) );
  NAND2_X1 U8762 ( .A1(n7141), .A2(n7140), .ZN(n9916) );
  NAND2_X1 U8763 ( .A1(n9917), .A2(n9916), .ZN(n7142) );
  NAND2_X1 U8764 ( .A1(n7143), .A2(n7142), .ZN(n9918) );
  NOR2_X1 U8765 ( .A1(n9919), .A2(n9918), .ZN(n7144) );
  NOR2_X1 U8766 ( .A1(n7145), .A2(n7144), .ZN(n7146) );
  NOR2_X1 U8767 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7146), .ZN(n9903) );
  AND2_X1 U8768 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7146), .ZN(n9904) );
  NOR2_X1 U8769 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9904), .ZN(n7147) );
  NOR2_X1 U8770 ( .A1(n9903), .A2(n7147), .ZN(n7148) );
  NAND2_X1 U8771 ( .A1(n7148), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7150) );
  XOR2_X1 U8772 ( .A(n7148), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n9902) );
  NAND2_X1 U8773 ( .A1(n9902), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7149) );
  NAND2_X1 U8774 ( .A1(n7150), .A2(n7149), .ZN(n7151) );
  NAND2_X1 U8775 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7151), .ZN(n7153) );
  XOR2_X1 U8776 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7151), .Z(n9901) );
  NAND2_X1 U8777 ( .A1(n9901), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7152) );
  NAND2_X1 U8778 ( .A1(n7153), .A2(n7152), .ZN(n7154) );
  NAND2_X1 U8779 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7154), .ZN(n7156) );
  XOR2_X1 U8780 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7154), .Z(n9913) );
  NAND2_X1 U8781 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9913), .ZN(n7155) );
  NAND2_X1 U8782 ( .A1(n7156), .A2(n7155), .ZN(n7157) );
  AND2_X1 U8783 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7157), .ZN(n7158) );
  INV_X1 U8784 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9912) );
  XNOR2_X1 U8785 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7157), .ZN(n9911) );
  NOR2_X1 U8786 ( .A1(n9912), .A2(n9911), .ZN(n9910) );
  NOR2_X1 U8787 ( .A1(n7158), .A2(n9910), .ZN(n9744) );
  NAND2_X1 U8788 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7159) );
  OAI21_X1 U8789 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7159), .ZN(n9743) );
  NOR2_X1 U8790 ( .A1(n9744), .A2(n9743), .ZN(n9742) );
  AOI21_X1 U8791 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9742), .ZN(n9741) );
  NAND2_X1 U8792 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7160) );
  OAI21_X1 U8793 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7160), .ZN(n9740) );
  NOR2_X1 U8794 ( .A1(n9741), .A2(n9740), .ZN(n9739) );
  AOI21_X1 U8795 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9739), .ZN(n9738) );
  NOR2_X1 U8796 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7161) );
  AOI21_X1 U8797 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7161), .ZN(n9737) );
  NAND2_X1 U8798 ( .A1(n9738), .A2(n9737), .ZN(n9736) );
  OAI21_X1 U8799 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9736), .ZN(n9734) );
  NAND2_X1 U8800 ( .A1(n9735), .A2(n9734), .ZN(n9733) );
  OAI21_X1 U8801 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9733), .ZN(n9731) );
  NAND2_X1 U8802 ( .A1(n9732), .A2(n9731), .ZN(n9730) );
  OAI21_X1 U8803 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9730), .ZN(n9728) );
  NAND2_X1 U8804 ( .A1(n9729), .A2(n9728), .ZN(n9727) );
  OAI21_X1 U8805 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9727), .ZN(n9725) );
  NAND2_X1 U8806 ( .A1(n9726), .A2(n9725), .ZN(n9724) );
  OAI21_X1 U8807 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9724), .ZN(n9722) );
  NAND2_X1 U8808 ( .A1(n9723), .A2(n9722), .ZN(n9721) );
  OAI21_X1 U8809 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9721), .ZN(n9907) );
  NOR2_X1 U8810 ( .A1(n9908), .A2(n9907), .ZN(n7162) );
  NAND2_X1 U8811 ( .A1(n9908), .A2(n9907), .ZN(n9906) );
  OAI21_X1 U8812 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7162), .A(n9906), .ZN(
        n7164) );
  XNOR2_X1 U8813 ( .A(n4667), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7163) );
  XNOR2_X1 U8814 ( .A(n7164), .B(n7163), .ZN(ADD_1071_U4) );
  OAI21_X1 U8815 ( .B1(n7166), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7165), .ZN(
        n7248) );
  XNOR2_X1 U8816 ( .A(n7249), .B(n7248), .ZN(n7167) );
  INV_X1 U8817 ( .A(n7167), .ZN(n7170) );
  INV_X1 U8818 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7168) );
  NOR2_X1 U8819 ( .A1(n7168), .A2(n7167), .ZN(n7250) );
  INV_X1 U8820 ( .A(n7250), .ZN(n7169) );
  OAI211_X1 U8821 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7170), .A(n9497), .B(
        n7169), .ZN(n7171) );
  NAND2_X1 U8822 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7536) );
  OAI211_X1 U8823 ( .C1(n9027), .C2(n7249), .A(n7171), .B(n7536), .ZN(n7178)
         );
  NOR2_X1 U8824 ( .A1(n7173), .A2(n7172), .ZN(n7175) );
  NOR2_X1 U8825 ( .A1(n7175), .A2(n7174), .ZN(n7243) );
  INV_X1 U8826 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9821) );
  AOI211_X1 U8827 ( .C1(n7176), .C2(n9821), .A(n7244), .B(n9490), .ZN(n7177)
         );
  AOI211_X1 U8828 ( .C1(n9500), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7178), .B(
        n7177), .ZN(n7179) );
  INV_X1 U8829 ( .A(n7179), .ZN(P1_U3256) );
  AOI21_X1 U8830 ( .B1(n7181), .B2(n7180), .A(n8947), .ZN(n7183) );
  NAND2_X1 U8831 ( .A1(n7183), .A2(n7182), .ZN(n7188) );
  NAND2_X1 U8832 ( .A1(n8968), .A2(n8940), .ZN(n7184) );
  NAND2_X1 U8833 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3084), .ZN(n8981) );
  OAI211_X1 U8834 ( .C1(n7210), .C2(n8954), .A(n7184), .B(n8981), .ZN(n7185)
         );
  AOI21_X1 U8835 ( .B1(n8957), .B2(n7186), .A(n7185), .ZN(n7187) );
  OAI211_X1 U8836 ( .C1(n9438), .C2(n8960), .A(n7188), .B(n7187), .ZN(P1_U3234) );
  INV_X1 U8837 ( .A(n7189), .ZN(n7193) );
  OAI222_X1 U8838 ( .A1(n8333), .A2(n7191), .B1(n8334), .B2(n7193), .C1(n7190), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U8839 ( .A1(n8856), .A2(n7194), .B1(n8098), .B2(n7193), .C1(n7192), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI21_X1 U8840 ( .B1(n7197), .B2(n7196), .A(n7195), .ZN(n7198) );
  NAND2_X1 U8841 ( .A1(n7198), .A2(n8410), .ZN(n7203) );
  INV_X1 U8842 ( .A(n7449), .ZN(n8427) );
  NAND2_X1 U8843 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n8051) );
  INV_X1 U8844 ( .A(n8051), .ZN(n7201) );
  INV_X1 U8845 ( .A(n8358), .ZN(n7451) );
  INV_X1 U8846 ( .A(n7299), .ZN(n7199) );
  OAI22_X1 U8847 ( .A1(n7451), .A2(n7199), .B1(n7302), .B2(n8416), .ZN(n7200)
         );
  AOI211_X1 U8848 ( .C1(n8374), .C2(n8427), .A(n7201), .B(n7200), .ZN(n7202)
         );
  OAI211_X1 U8849 ( .C1(n4354), .C2(n8422), .A(n7203), .B(n7202), .ZN(P2_U3217) );
  INV_X1 U8850 ( .A(n9377), .ZN(n9410) );
  NAND2_X1 U8851 ( .A1(n7204), .A2(n9410), .ZN(n7205) );
  NAND2_X1 U8852 ( .A1(n9416), .A2(n7210), .ZN(n7752) );
  NAND2_X1 U8853 ( .A1(n7634), .A2(n7752), .ZN(n9418) );
  INV_X1 U8854 ( .A(n7210), .ZN(n8967) );
  INV_X1 U8855 ( .A(n9408), .ZN(n7290) );
  OR2_X1 U8856 ( .A1(n7376), .A2(n7290), .ZN(n7632) );
  NAND2_X1 U8857 ( .A1(n7376), .A2(n7290), .ZN(n7629) );
  INV_X1 U8858 ( .A(n7809), .ZN(n7207) );
  XNOR2_X1 U8859 ( .A(n7227), .B(n7207), .ZN(n7259) );
  INV_X1 U8860 ( .A(n7634), .ZN(n7209) );
  XNOR2_X1 U8861 ( .A(n7230), .B(n7809), .ZN(n7212) );
  INV_X1 U8862 ( .A(n8966), .ZN(n7479) );
  OAI22_X1 U8863 ( .A1(n7479), .A2(n9376), .B1(n7210), .B2(n9378), .ZN(n7211)
         );
  AOI21_X1 U8864 ( .B1(n7212), .B2(n9412), .A(n7211), .ZN(n7213) );
  OAI21_X1 U8865 ( .B1(n7259), .B2(n9382), .A(n7213), .ZN(n7262) );
  NAND2_X1 U8866 ( .A1(n7262), .A2(n7027), .ZN(n7220) );
  INV_X1 U8867 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7215) );
  INV_X1 U8868 ( .A(n7214), .ZN(n7374) );
  OAI22_X1 U8869 ( .A1(n7027), .A2(n7215), .B1(n7374), .B2(n9209), .ZN(n7218)
         );
  AND2_X1 U8870 ( .A1(n9422), .A2(n7376), .ZN(n7216) );
  OR2_X1 U8871 ( .A1(n7216), .A2(n7234), .ZN(n7261) );
  NOR2_X1 U8872 ( .A1(n7261), .A2(n9088), .ZN(n7217) );
  AOI211_X1 U8873 ( .C1(n9415), .C2(n7376), .A(n7218), .B(n7217), .ZN(n7219)
         );
  OAI211_X1 U8874 ( .C1(n7259), .C2(n7491), .A(n7220), .B(n7219), .ZN(P1_U3278) );
  INV_X1 U8875 ( .A(n7221), .ZN(n7225) );
  OAI222_X1 U8876 ( .A1(n7223), .A2(P1_U3084), .B1(n8334), .B2(n7225), .C1(
        n7222), .C2(n8333), .ZN(P1_U3327) );
  OAI222_X1 U8877 ( .A1(n7226), .A2(P2_U3152), .B1(n8858), .B2(n7225), .C1(
        n7224), .C2(n8856), .ZN(P2_U3332) );
  OR2_X1 U8878 ( .A1(n9339), .A2(n7479), .ZN(n7642) );
  NAND2_X1 U8879 ( .A1(n9339), .A2(n7479), .ZN(n7640) );
  OAI21_X1 U8880 ( .B1(n7376), .B2(n9408), .A(n7227), .ZN(n7228) );
  INV_X1 U8881 ( .A(n7376), .ZN(n7260) );
  XOR2_X1 U8882 ( .A(n7811), .B(n7410), .Z(n9341) );
  INV_X1 U8883 ( .A(n7629), .ZN(n7229) );
  AOI21_X1 U8884 ( .B1(n7230), .B2(n7809), .A(n7229), .ZN(n7231) );
  NAND2_X1 U8885 ( .A1(n7231), .A2(n7811), .ZN(n7412) );
  OAI211_X1 U8886 ( .C1(n7231), .C2(n7811), .A(n7412), .B(n9412), .ZN(n7233)
         );
  AOI22_X1 U8887 ( .A1(n9409), .A2(n9408), .B1(n8965), .B2(n9407), .ZN(n7232)
         );
  NAND2_X1 U8888 ( .A1(n7233), .A2(n7232), .ZN(n9337) );
  INV_X1 U8889 ( .A(n7234), .ZN(n7235) );
  AOI211_X1 U8890 ( .C1(n9339), .C2(n7235), .A(n9542), .B(n7484), .ZN(n9338)
         );
  NAND2_X1 U8891 ( .A1(n9338), .A2(n9426), .ZN(n7237) );
  AOI22_X1 U8892 ( .A1(n9386), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7466), .B2(
        n9414), .ZN(n7236) );
  OAI211_X1 U8893 ( .C1(n7463), .C2(n9237), .A(n7237), .B(n7236), .ZN(n7238)
         );
  AOI21_X1 U8894 ( .B1(n9337), .B2(n7027), .A(n7238), .ZN(n7239) );
  OAI21_X1 U8895 ( .B1(n9341), .B2(n9247), .A(n7239), .ZN(P1_U3277) );
  INV_X1 U8896 ( .A(n7240), .ZN(n7270) );
  NAND2_X1 U8897 ( .A1(n9366), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n7241) );
  OAI211_X1 U8898 ( .C1(n7270), .C2(n8334), .A(n7242), .B(n7241), .ZN(P1_U3326) );
  NOR2_X1 U8899 ( .A1(n7243), .A2(n7249), .ZN(n7245) );
  NAND2_X1 U8900 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8996), .ZN(n7246) );
  OAI21_X1 U8901 ( .B1(n8996), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7246), .ZN(
        n7247) );
  AOI211_X1 U8902 ( .C1(n4308), .C2(n7247), .A(n8995), .B(n9490), .ZN(n7258)
         );
  NOR2_X1 U8903 ( .A1(n7249), .A2(n7248), .ZN(n7251) );
  NOR2_X1 U8904 ( .A1(n7251), .A2(n7250), .ZN(n7253) );
  XNOR2_X1 U8905 ( .A(n8996), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7252) );
  NOR2_X1 U8906 ( .A1(n7253), .A2(n7252), .ZN(n8992) );
  AOI211_X1 U8907 ( .C1(n7253), .C2(n7252), .A(n8992), .B(n9476), .ZN(n7257)
         );
  NAND2_X1 U8908 ( .A1(n9500), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7254) );
  NAND2_X1 U8909 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n7520) );
  OAI211_X1 U8910 ( .C1(n9027), .C2(n7255), .A(n7254), .B(n7520), .ZN(n7256)
         );
  OR3_X1 U8911 ( .A1(n7258), .A2(n7257), .A3(n7256), .ZN(P1_U3257) );
  INV_X1 U8912 ( .A(n7259), .ZN(n7264) );
  OAI22_X1 U8913 ( .A1(n7261), .A2(n9542), .B1(n7260), .B2(n9540), .ZN(n7263)
         );
  AOI211_X1 U8914 ( .C1(n9538), .C2(n7264), .A(n7263), .B(n7262), .ZN(n7266)
         );
  MUX2_X1 U8915 ( .A(n6668), .B(n7266), .S(n9562), .Z(n7265) );
  INV_X1 U8916 ( .A(n7265), .ZN(P1_U3536) );
  INV_X1 U8917 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7267) );
  MUX2_X1 U8918 ( .A(n7267), .B(n7266), .S(n9550), .Z(n7268) );
  INV_X1 U8919 ( .A(n7268), .ZN(P1_U3493) );
  OAI222_X1 U8920 ( .A1(n8856), .A2(n7271), .B1(n8858), .B2(n7270), .C1(n7269), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U8921 ( .A(n7272), .ZN(n7273) );
  NOR2_X1 U8922 ( .A1(n7274), .A2(n7273), .ZN(n7276) );
  XNOR2_X1 U8923 ( .A(n7276), .B(n7275), .ZN(n7280) );
  AOI22_X1 U8924 ( .A1(n8375), .A2(n8428), .B1(n8358), .B2(n7384), .ZN(n7277)
         );
  NAND2_X1 U8925 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8036) );
  OAI211_X1 U8926 ( .C1(n7438), .C2(n8414), .A(n7277), .B(n8036), .ZN(n7278)
         );
  AOI21_X1 U8927 ( .B1(n8807), .B2(n8406), .A(n7278), .ZN(n7279) );
  OAI21_X1 U8928 ( .B1(n7280), .B2(n8408), .A(n7279), .ZN(P2_U3243) );
  INV_X1 U8929 ( .A(n7281), .ZN(n8335) );
  NAND2_X1 U8930 ( .A1(n9366), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n7282) );
  OAI211_X1 U8931 ( .C1(n8335), .C2(n8334), .A(n7283), .B(n7282), .ZN(P1_U3325) );
  INV_X1 U8932 ( .A(n7284), .ZN(n7285) );
  AOI21_X1 U8933 ( .B1(n7287), .B2(n7286), .A(n7285), .ZN(n7294) );
  NAND2_X1 U8934 ( .A1(n9410), .A2(n8940), .ZN(n7289) );
  OAI211_X1 U8935 ( .C1(n7290), .C2(n8954), .A(n7289), .B(n7288), .ZN(n7292)
         );
  INV_X1 U8936 ( .A(n9416), .ZN(n9433) );
  NOR2_X1 U8937 ( .A1(n9433), .A2(n8960), .ZN(n7291) );
  AOI211_X1 U8938 ( .C1(n9413), .C2(n8957), .A(n7292), .B(n7291), .ZN(n7293)
         );
  OAI21_X1 U8939 ( .B1(n7294), .B2(n8947), .A(n7293), .ZN(P1_U3222) );
  NAND2_X1 U8940 ( .A1(n8812), .A2(n8428), .ZN(n7296) );
  NAND2_X1 U8941 ( .A1(n7379), .A2(n7296), .ZN(n8301) );
  AOI21_X1 U8942 ( .B1(n7297), .B2(n8301), .A(n7380), .ZN(n8817) );
  AOI21_X1 U8943 ( .B1(n8812), .B2(n7298), .A(n7381), .ZN(n8813) );
  AOI22_X1 U8944 ( .A1(n9588), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7299), .B2(
        n9576), .ZN(n7300) );
  OAI21_X1 U8945 ( .B1(n4354), .B2(n8674), .A(n7300), .ZN(n7305) );
  XNOR2_X1 U8946 ( .A(n7388), .B(n8301), .ZN(n7303) );
  INV_X1 U8947 ( .A(n7302), .ZN(n8429) );
  AOI222_X1 U8948 ( .A1(n8492), .A2(n7303), .B1(n8429), .B2(n8678), .C1(n8427), 
        .C2(n8680), .ZN(n8815) );
  NOR2_X1 U8949 ( .A1(n8815), .A2(n9588), .ZN(n7304) );
  AOI211_X1 U8950 ( .C1(n8813), .C2(n8719), .A(n7305), .B(n7304), .ZN(n7306)
         );
  OAI21_X1 U8951 ( .B1(n8817), .B2(n8686), .A(n7306), .ZN(P2_U3282) );
  INV_X1 U8952 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7307) );
  AOI22_X1 U8953 ( .A1(n8053), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n7307), .B2(
        n7353), .ZN(n8049) );
  INV_X1 U8954 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7308) );
  AOI22_X1 U8955 ( .A1(n7350), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n7308), .B2(
        n7908), .ZN(n7900) );
  AOI21_X1 U8956 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n7310), .A(n7309), .ZN(
        n8002) );
  XNOR2_X1 U8957 ( .A(n8006), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n8001) );
  NOR2_X1 U8958 ( .A1(n8002), .A2(n8001), .ZN(n8000) );
  AOI21_X1 U8959 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n8006), .A(n8000), .ZN(
        n7989) );
  XNOR2_X1 U8960 ( .A(n7340), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n7988) );
  OR2_X1 U8961 ( .A1(n8080), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7312) );
  NAND2_X1 U8962 ( .A1(n8080), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7311) );
  NAND2_X1 U8963 ( .A1(n7312), .A2(n7311), .ZN(n8075) );
  INV_X1 U8964 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7313) );
  MUX2_X1 U8965 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7313), .S(n7985), .Z(n7977)
         );
  NOR2_X1 U8966 ( .A1(n4275), .A2(n7977), .ZN(n7976) );
  NAND2_X1 U8967 ( .A1(n7334), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7314) );
  OAI21_X1 U8968 ( .B1(n7334), .B2(P2_REG1_REG_7__SCAN_IN), .A(n7314), .ZN(
        n7965) );
  INV_X1 U8969 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7315) );
  MUX2_X1 U8970 ( .A(n7315), .B(P2_REG1_REG_8__SCAN_IN), .S(n7331), .Z(n7953)
         );
  AOI21_X1 U8971 ( .B1(n7331), .B2(P2_REG1_REG_8__SCAN_IN), .A(n7952), .ZN(
        n7942) );
  INV_X1 U8972 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7316) );
  MUX2_X1 U8973 ( .A(n7316), .B(P2_REG1_REG_9__SCAN_IN), .S(n7328), .Z(n7941)
         );
  NOR2_X1 U8974 ( .A1(n7942), .A2(n7941), .ZN(n7940) );
  INV_X1 U8975 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7317) );
  MUX2_X1 U8976 ( .A(n7317), .B(P2_REG1_REG_10__SCAN_IN), .S(n7325), .Z(n7930)
         );
  INV_X1 U8977 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7318) );
  MUX2_X1 U8978 ( .A(n7318), .B(P2_REG1_REG_11__SCAN_IN), .S(n7347), .Z(n8062)
         );
  AOI21_X1 U8979 ( .B1(n7347), .B2(P2_REG1_REG_11__SCAN_IN), .A(n8060), .ZN(
        n7911) );
  INV_X1 U8980 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7319) );
  MUX2_X1 U8981 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7319), .S(n7917), .Z(n7910)
         );
  NAND2_X1 U8982 ( .A1(n7911), .A2(n7910), .ZN(n7909) );
  NAND2_X1 U8983 ( .A1(n7924), .A2(n7319), .ZN(n7320) );
  NAND2_X1 U8984 ( .A1(n7909), .A2(n7320), .ZN(n7901) );
  NAND2_X1 U8985 ( .A1(n7900), .A2(n7901), .ZN(n7899) );
  NOR2_X1 U8986 ( .A1(n8039), .A2(n7321), .ZN(n7322) );
  INV_X1 U8987 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8034) );
  NOR2_X1 U8988 ( .A1(n8034), .A2(n8035), .ZN(n8033) );
  NOR2_X1 U8989 ( .A1(n7322), .A2(n8033), .ZN(n7324) );
  XOR2_X1 U8990 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n7884), .Z(n7323) );
  NAND2_X1 U8991 ( .A1(n7323), .A2(n7324), .ZN(n7885) );
  OAI21_X1 U8992 ( .B1(n7324), .B2(n7323), .A(n7885), .ZN(n7365) );
  INV_X1 U8993 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7352) );
  INV_X1 U8994 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7351) );
  NAND2_X1 U8995 ( .A1(n7917), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7349) );
  INV_X1 U8996 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7918) );
  INV_X1 U8997 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7348) );
  NAND2_X1 U8998 ( .A1(n7325), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7346) );
  INV_X1 U8999 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7326) );
  MUX2_X1 U9000 ( .A(n7326), .B(P2_REG2_REG_10__SCAN_IN), .S(n7325), .Z(n7327)
         );
  INV_X1 U9001 ( .A(n7327), .ZN(n7926) );
  NAND2_X1 U9002 ( .A1(n7328), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7345) );
  INV_X1 U9003 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7329) );
  MUX2_X1 U9004 ( .A(n7329), .B(P2_REG2_REG_9__SCAN_IN), .S(n7328), .Z(n7330)
         );
  INV_X1 U9005 ( .A(n7330), .ZN(n7946) );
  NAND2_X1 U9006 ( .A1(n7331), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7344) );
  INV_X1 U9007 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7332) );
  MUX2_X1 U9008 ( .A(n7332), .B(P2_REG2_REG_8__SCAN_IN), .S(n7331), .Z(n7333)
         );
  INV_X1 U9009 ( .A(n7333), .ZN(n7958) );
  NAND2_X1 U9010 ( .A1(n7334), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7343) );
  INV_X1 U9011 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7335) );
  MUX2_X1 U9012 ( .A(n7335), .B(P2_REG2_REG_7__SCAN_IN), .S(n7334), .Z(n7336)
         );
  INV_X1 U9013 ( .A(n7336), .ZN(n7971) );
  INV_X1 U9014 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9817) );
  MUX2_X1 U9015 ( .A(n9817), .B(P2_REG2_REG_6__SCAN_IN), .S(n7985), .Z(n7981)
         );
  NAND2_X1 U9016 ( .A1(n8080), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7342) );
  NOR2_X1 U9017 ( .A1(n7337), .A2(n6173), .ZN(n8005) );
  INV_X1 U9018 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7338) );
  MUX2_X1 U9019 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n7338), .S(n8006), .Z(n7339)
         );
  OAI21_X1 U9020 ( .B1(n8011), .B2(n8005), .A(n7339), .ZN(n8009) );
  NAND2_X1 U9021 ( .A1(n8006), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7994) );
  MUX2_X1 U9022 ( .A(n9847), .B(P2_REG2_REG_4__SCAN_IN), .S(n7340), .Z(n7993)
         );
  AOI21_X1 U9023 ( .B1(n8009), .B2(n7994), .A(n7993), .ZN(n7992) );
  AOI21_X1 U9024 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n7340), .A(n7992), .ZN(
        n8072) );
  MUX2_X1 U9025 ( .A(n6649), .B(P2_REG2_REG_5__SCAN_IN), .S(n8080), .Z(n8071)
         );
  OR2_X1 U9026 ( .A1(n8072), .A2(n8071), .ZN(n7341) );
  NAND2_X1 U9027 ( .A1(n7342), .A2(n7341), .ZN(n7982) );
  NAND2_X1 U9028 ( .A1(n7981), .A2(n7982), .ZN(n7980) );
  OAI21_X1 U9029 ( .B1(n7985), .B2(n9817), .A(n7980), .ZN(n7970) );
  NAND2_X1 U9030 ( .A1(n7971), .A2(n7970), .ZN(n7969) );
  NAND2_X1 U9031 ( .A1(n7343), .A2(n7969), .ZN(n7959) );
  NAND2_X1 U9032 ( .A1(n7958), .A2(n7959), .ZN(n7957) );
  NAND2_X1 U9033 ( .A1(n7344), .A2(n7957), .ZN(n7947) );
  NAND2_X1 U9034 ( .A1(n7946), .A2(n7947), .ZN(n7945) );
  NAND2_X1 U9035 ( .A1(n7345), .A2(n7945), .ZN(n7927) );
  NAND2_X1 U9036 ( .A1(n7926), .A2(n7927), .ZN(n7925) );
  NAND2_X1 U9037 ( .A1(n7346), .A2(n7925), .ZN(n8059) );
  MUX2_X1 U9038 ( .A(n7348), .B(P2_REG2_REG_11__SCAN_IN), .S(n7347), .Z(n8058)
         );
  NOR2_X1 U9039 ( .A1(n8059), .A2(n8058), .ZN(n8057) );
  AOI21_X1 U9040 ( .B1(n8067), .B2(n7348), .A(n8057), .ZN(n7921) );
  OAI211_X1 U9041 ( .C1(n7917), .C2(P2_REG2_REG_12__SCAN_IN), .A(n7921), .B(
        n7349), .ZN(n7919) );
  NAND2_X1 U9042 ( .A1(n7349), .A2(n7919), .ZN(n7897) );
  AOI22_X1 U9043 ( .A1(n7350), .A2(n7351), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7908), .ZN(n7896) );
  NOR2_X1 U9044 ( .A1(n7897), .A2(n7896), .ZN(n7895) );
  AOI21_X1 U9045 ( .B1(n7908), .B2(n7351), .A(n7895), .ZN(n8046) );
  AOI22_X1 U9046 ( .A1(n8053), .A2(n7352), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7353), .ZN(n8045) );
  NOR2_X1 U9047 ( .A1(n8046), .A2(n8045), .ZN(n8044) );
  AOI21_X1 U9048 ( .B1(n7353), .B2(n7352), .A(n8044), .ZN(n7355) );
  NOR2_X1 U9049 ( .A1(n7354), .A2(n7355), .ZN(n7356) );
  XNOR2_X1 U9050 ( .A(n7355), .B(n7354), .ZN(n8032) );
  NOR2_X1 U9051 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8032), .ZN(n8031) );
  NOR2_X1 U9052 ( .A1(n7356), .A2(n8031), .ZN(n7360) );
  INV_X1 U9053 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7358) );
  NAND2_X1 U9054 ( .A1(n7884), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7880) );
  INV_X1 U9055 ( .A(n7880), .ZN(n7357) );
  AOI21_X1 U9056 ( .B1(n7358), .B2(n7363), .A(n7357), .ZN(n7359) );
  INV_X1 U9057 ( .A(n8450), .ZN(n8454) );
  NAND2_X1 U9058 ( .A1(n7359), .A2(n7360), .ZN(n7879) );
  OAI211_X1 U9059 ( .C1(n7360), .C2(n7359), .A(n8454), .B(n7879), .ZN(n7362)
         );
  AND2_X1 U9060 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n7453) );
  AOI21_X1 U9061 ( .B1(n8079), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7453), .ZN(
        n7361) );
  OAI211_X1 U9062 ( .C1(n8448), .C2(n7363), .A(n7362), .B(n7361), .ZN(n7364)
         );
  AOI21_X1 U9063 ( .B1(n8453), .B2(n7365), .A(n7364), .ZN(n7366) );
  INV_X1 U9064 ( .A(n7366), .ZN(P2_U3261) );
  XNOR2_X1 U9065 ( .A(n7368), .B(n7367), .ZN(n7369) );
  XNOR2_X1 U9066 ( .A(n7370), .B(n7369), .ZN(n7378) );
  OAI21_X1 U9067 ( .B1(n7479), .B2(n8954), .A(n7371), .ZN(n7372) );
  AOI21_X1 U9068 ( .B1(n8940), .B2(n8967), .A(n7372), .ZN(n7373) );
  OAI21_X1 U9069 ( .B1(n7541), .B2(n7374), .A(n7373), .ZN(n7375) );
  AOI21_X1 U9070 ( .B1(n7376), .B2(n8914), .A(n7375), .ZN(n7377) );
  OAI21_X1 U9071 ( .B1(n7378), .B2(n8947), .A(n7377), .ZN(P1_U3232) );
  NAND2_X1 U9072 ( .A1(n8807), .A2(n7449), .ZN(n8205) );
  XOR2_X1 U9073 ( .A(n8303), .B(n4306), .Z(n8811) );
  INV_X1 U9074 ( .A(n7381), .ZN(n7383) );
  NAND2_X1 U9075 ( .A1(n7381), .A2(n7386), .ZN(n7430) );
  INV_X1 U9076 ( .A(n7430), .ZN(n7382) );
  AOI21_X1 U9077 ( .B1(n8807), .B2(n7383), .A(n7382), .ZN(n8808) );
  AOI22_X1 U9078 ( .A1(n9588), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7384), .B2(
        n9576), .ZN(n7385) );
  OAI21_X1 U9079 ( .B1(n7386), .B2(n8674), .A(n7385), .ZN(n7391) );
  INV_X1 U9080 ( .A(n8301), .ZN(n7387) );
  XOR2_X1 U9081 ( .A(n8303), .B(n7396), .Z(n7389) );
  INV_X1 U9082 ( .A(n7438), .ZN(n8426) );
  AOI222_X1 U9083 ( .A1(n8492), .A2(n7389), .B1(n8426), .B2(n8680), .C1(n8428), 
        .C2(n8678), .ZN(n8810) );
  NOR2_X1 U9084 ( .A1(n8810), .A2(n9588), .ZN(n7390) );
  AOI211_X1 U9085 ( .C1(n8808), .C2(n8719), .A(n7391), .B(n7390), .ZN(n7392)
         );
  OAI21_X1 U9086 ( .B1(n8811), .B2(n8686), .A(n7392), .ZN(P2_U3281) );
  OR2_X1 U9087 ( .A1(n8802), .A2(n7438), .ZN(n8210) );
  NAND2_X1 U9088 ( .A1(n8802), .A2(n7438), .ZN(n8209) );
  AOI21_X1 U9089 ( .B1(n8802), .B2(n8426), .A(n7422), .ZN(n7393) );
  NAND2_X1 U9090 ( .A1(n8799), .A2(n7425), .ZN(n8126) );
  NAND2_X1 U9091 ( .A1(n8129), .A2(n8126), .ZN(n7398) );
  NAND2_X1 U9092 ( .A1(n7393), .A2(n7398), .ZN(n8474) );
  OAI21_X1 U9093 ( .B1(n7393), .B2(n7398), .A(n8474), .ZN(n7394) );
  INV_X1 U9094 ( .A(n7394), .ZN(n8801) );
  AOI22_X1 U9095 ( .A1(n8799), .A2(n9577), .B1(n9588), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n7408) );
  INV_X1 U9096 ( .A(n8662), .ZN(n8475) );
  INV_X1 U9097 ( .A(n8206), .ZN(n7395) );
  INV_X1 U9098 ( .A(n8209), .ZN(n7397) );
  INV_X1 U9099 ( .A(n7398), .ZN(n8306) );
  XNOR2_X1 U9100 ( .A(n8100), .B(n8306), .ZN(n7399) );
  OAI222_X1 U9101 ( .A1(n8693), .A2(n8475), .B1(n8695), .B2(n7438), .C1(n8643), 
        .C2(n7399), .ZN(n8797) );
  NOR2_X1 U9102 ( .A1(n7430), .A2(n8802), .ZN(n7401) );
  INV_X1 U9103 ( .A(n7401), .ZN(n7403) );
  INV_X1 U9104 ( .A(n8799), .ZN(n7400) );
  NAND2_X1 U9105 ( .A1(n7401), .A2(n7400), .ZN(n8671) );
  INV_X1 U9106 ( .A(n8671), .ZN(n7402) );
  AOI211_X1 U9107 ( .C1(n8799), .C2(n7403), .A(n9692), .B(n7402), .ZN(n8798)
         );
  INV_X1 U9108 ( .A(n8798), .ZN(n7405) );
  INV_X1 U9109 ( .A(n7404), .ZN(n7439) );
  OAI22_X1 U9110 ( .A1(n7405), .A2(n8567), .B1(n8705), .B2(n7439), .ZN(n7406)
         );
  OAI21_X1 U9111 ( .B1(n8797), .B2(n7406), .A(n8699), .ZN(n7407) );
  OAI211_X1 U9112 ( .C1(n8801), .C2(n8686), .A(n7408), .B(n7407), .ZN(P2_U3279) );
  INV_X1 U9113 ( .A(n8965), .ZN(n7462) );
  OR2_X1 U9114 ( .A1(n9328), .A2(n7537), .ZN(n7651) );
  NAND2_X1 U9115 ( .A1(n9328), .A2(n7537), .ZN(n7757) );
  NAND2_X1 U9116 ( .A1(n7651), .A2(n7757), .ZN(n7814) );
  XNOR2_X1 U9117 ( .A(n7469), .B(n7814), .ZN(n9330) );
  INV_X1 U9118 ( .A(n8963), .ZN(n7521) );
  NAND2_X1 U9119 ( .A1(n9331), .A2(n7462), .ZN(n7755) );
  OR2_X1 U9120 ( .A1(n9331), .A2(n7462), .ZN(n7647) );
  NAND2_X1 U9121 ( .A1(n7471), .A2(n7647), .ZN(n7413) );
  INV_X1 U9122 ( .A(n7814), .ZN(n7649) );
  XNOR2_X1 U9123 ( .A(n7413), .B(n7649), .ZN(n7414) );
  OAI222_X1 U9124 ( .A1(n9378), .A2(n7462), .B1(n9376), .B2(n7521), .C1(n9203), 
        .C2(n7414), .ZN(n9326) );
  INV_X1 U9125 ( .A(n9328), .ZN(n7419) );
  NAND2_X1 U9126 ( .A1(n7484), .A2(n7490), .ZN(n7485) );
  OR2_X2 U9127 ( .A1(n7485), .A2(n9328), .ZN(n7473) );
  INV_X1 U9128 ( .A(n7473), .ZN(n7415) );
  AOI211_X1 U9129 ( .C1(n9328), .C2(n7485), .A(n9542), .B(n7415), .ZN(n9327)
         );
  NAND2_X1 U9130 ( .A1(n9327), .A2(n9426), .ZN(n7418) );
  AOI22_X1 U9131 ( .A1(n9386), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7416), .B2(
        n9414), .ZN(n7417) );
  OAI211_X1 U9132 ( .C1(n7419), .C2(n9237), .A(n7418), .B(n7417), .ZN(n7420)
         );
  AOI21_X1 U9133 ( .B1(n9326), .B2(n7027), .A(n7420), .ZN(n7421) );
  OAI21_X1 U9134 ( .B1(n9330), .B2(n9247), .A(n7421), .ZN(P1_U3275) );
  AOI21_X1 U9135 ( .B1(n8304), .B2(n7423), .A(n7422), .ZN(n7432) );
  XOR2_X1 U9136 ( .A(n8304), .B(n7424), .Z(n7427) );
  INV_X1 U9137 ( .A(n7425), .ZN(n8679) );
  AOI22_X1 U9138 ( .A1(n8678), .A2(n8427), .B1(n8679), .B2(n8680), .ZN(n7426)
         );
  OAI21_X1 U9139 ( .B1(n7427), .B2(n8643), .A(n7426), .ZN(n7428) );
  AOI21_X1 U9140 ( .B1(n7432), .B2(n7429), .A(n7428), .ZN(n8805) );
  XOR2_X1 U9141 ( .A(n8802), .B(n7430), .Z(n8803) );
  INV_X1 U9142 ( .A(n8802), .ZN(n7456) );
  AOI22_X1 U9143 ( .A1(n9588), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n7448), .B2(
        n9576), .ZN(n7431) );
  OAI21_X1 U9144 ( .B1(n7456), .B2(n8674), .A(n7431), .ZN(n7434) );
  INV_X1 U9145 ( .A(n7432), .ZN(n8806) );
  NOR2_X1 U9146 ( .A1(n8806), .A2(n9584), .ZN(n7433) );
  AOI211_X1 U9147 ( .C1(n8803), .C2(n8719), .A(n7434), .B(n7433), .ZN(n7435)
         );
  OAI21_X1 U9148 ( .B1(n9588), .B2(n8805), .A(n7435), .ZN(P2_U3280) );
  XNOR2_X1 U9149 ( .A(n7437), .B(n7436), .ZN(n7443) );
  OAI22_X1 U9150 ( .A1(n8414), .A2(n8475), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5204), .ZN(n7441) );
  OAI22_X1 U9151 ( .A1(n7451), .A2(n7439), .B1(n7438), .B2(n8416), .ZN(n7440)
         );
  AOI211_X1 U9152 ( .C1(n8799), .C2(n8406), .A(n7441), .B(n7440), .ZN(n7442)
         );
  OAI21_X1 U9153 ( .B1(n7443), .B2(n8408), .A(n7442), .ZN(P2_U3230) );
  OAI21_X1 U9154 ( .B1(n7446), .B2(n7445), .A(n7444), .ZN(n7447) );
  NAND2_X1 U9155 ( .A1(n7447), .A2(n8410), .ZN(n7455) );
  INV_X1 U9156 ( .A(n7448), .ZN(n7450) );
  OAI22_X1 U9157 ( .A1(n7451), .A2(n7450), .B1(n7449), .B2(n8416), .ZN(n7452)
         );
  AOI211_X1 U9158 ( .C1(n8374), .C2(n8679), .A(n7453), .B(n7452), .ZN(n7454)
         );
  OAI211_X1 U9159 ( .C1(n7456), .C2(n8422), .A(n7455), .B(n7454), .ZN(P2_U3228) );
  XNOR2_X1 U9160 ( .A(n7458), .B(n7457), .ZN(n7459) );
  XNOR2_X1 U9161 ( .A(n7529), .B(n7459), .ZN(n7468) );
  NAND2_X1 U9162 ( .A1(n8940), .A2(n9408), .ZN(n7461) );
  OAI211_X1 U9163 ( .C1(n7462), .C2(n8954), .A(n7461), .B(n7460), .ZN(n7465)
         );
  NOR2_X1 U9164 ( .A1(n7463), .A2(n8960), .ZN(n7464) );
  AOI211_X1 U9165 ( .C1(n7466), .C2(n8957), .A(n7465), .B(n7464), .ZN(n7467)
         );
  OAI21_X1 U9166 ( .B1(n7468), .B2(n8947), .A(n7467), .ZN(P1_U3213) );
  INV_X1 U9167 ( .A(n7537), .ZN(n8964) );
  NOR2_X1 U9168 ( .A1(n9323), .A2(n7521), .ZN(n7656) );
  NAND2_X1 U9169 ( .A1(n9323), .A2(n7521), .ZN(n7654) );
  INV_X1 U9170 ( .A(n7654), .ZN(n7470) );
  OR2_X1 U9171 ( .A1(n7656), .A2(n7470), .ZN(n7815) );
  INV_X1 U9172 ( .A(n7815), .ZN(n7653) );
  XNOR2_X1 U9173 ( .A(n7502), .B(n7653), .ZN(n9325) );
  AND2_X1 U9174 ( .A1(n7651), .A2(n7647), .ZN(n7736) );
  XNOR2_X1 U9175 ( .A(n7506), .B(n7653), .ZN(n7472) );
  OAI222_X1 U9176 ( .A1(n9376), .A2(n8882), .B1(n9378), .B2(n7537), .C1(n7472), 
        .C2(n9203), .ZN(n9321) );
  INV_X1 U9177 ( .A(n9323), .ZN(n7548) );
  AOI211_X1 U9178 ( .C1(n9323), .C2(n7473), .A(n9542), .B(n7503), .ZN(n9322)
         );
  NAND2_X1 U9179 ( .A1(n9322), .A2(n9426), .ZN(n7475) );
  AOI22_X1 U9180 ( .A1(n9386), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n7551), .B2(
        n9414), .ZN(n7474) );
  OAI211_X1 U9181 ( .C1(n7548), .C2(n9237), .A(n7475), .B(n7474), .ZN(n7476)
         );
  AOI21_X1 U9182 ( .B1(n9321), .B2(n7027), .A(n7476), .ZN(n7477) );
  OAI21_X1 U9183 ( .B1(n9325), .B2(n9247), .A(n7477), .ZN(P1_U3274) );
  AND2_X1 U9184 ( .A1(n7647), .A2(n7755), .ZN(n7645) );
  INV_X1 U9185 ( .A(n7645), .ZN(n7813) );
  XNOR2_X1 U9186 ( .A(n7478), .B(n7813), .ZN(n7483) );
  OAI22_X1 U9187 ( .A1(n7479), .A2(n9378), .B1(n7537), .B2(n9376), .ZN(n7482)
         );
  XNOR2_X1 U9188 ( .A(n7480), .B(n7813), .ZN(n9336) );
  NOR2_X1 U9189 ( .A1(n9336), .A2(n9382), .ZN(n7481) );
  AOI211_X1 U9190 ( .C1(n9412), .C2(n7483), .A(n7482), .B(n7481), .ZN(n9334)
         );
  INV_X1 U9191 ( .A(n7484), .ZN(n7487) );
  INV_X1 U9192 ( .A(n7485), .ZN(n7486) );
  AOI21_X1 U9193 ( .B1(n9331), .B2(n7487), .A(n7486), .ZN(n9332) );
  AOI22_X1 U9194 ( .A1(n9430), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7488), .B2(
        n9414), .ZN(n7489) );
  OAI21_X1 U9195 ( .B1(n7490), .B2(n9237), .A(n7489), .ZN(n7493) );
  NOR2_X1 U9196 ( .A1(n9336), .A2(n7491), .ZN(n7492) );
  AOI211_X1 U9197 ( .C1(n9332), .C2(n9229), .A(n7493), .B(n7492), .ZN(n7494)
         );
  OAI21_X1 U9198 ( .B1(n9334), .B2(n9386), .A(n7494), .ZN(P1_U3276) );
  XNOR2_X1 U9199 ( .A(n7495), .B(n7496), .ZN(n7500) );
  AOI22_X1 U9200 ( .A1(n8375), .A2(n8679), .B1(n8358), .B2(n8672), .ZN(n7497)
         );
  NAND2_X1 U9201 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8025) );
  OAI211_X1 U9202 ( .C1(n8477), .C2(n8414), .A(n7497), .B(n8025), .ZN(n7498)
         );
  AOI21_X1 U9203 ( .B1(n8792), .B2(n8406), .A(n7498), .ZN(n7499) );
  OAI21_X1 U9204 ( .B1(n7500), .B2(n8408), .A(n7499), .ZN(P2_U3240) );
  NOR2_X1 U9205 ( .A1(n9323), .A2(n8963), .ZN(n7501) );
  OR2_X1 U9206 ( .A1(n9316), .A2(n8882), .ZN(n7657) );
  NAND2_X1 U9207 ( .A1(n9316), .A2(n8882), .ZN(n9067) );
  NAND2_X1 U9208 ( .A1(n7657), .A2(n9067), .ZN(n9053) );
  XNOR2_X1 U9209 ( .A(n9054), .B(n9053), .ZN(n9320) );
  INV_X1 U9210 ( .A(n7503), .ZN(n7504) );
  INV_X1 U9211 ( .A(n9316), .ZN(n8946) );
  AOI21_X1 U9212 ( .B1(n9316), .B2(n7504), .A(n9232), .ZN(n9317) );
  AOI22_X1 U9213 ( .A1(n9430), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n8943), .B2(
        n9414), .ZN(n7505) );
  OAI21_X1 U9214 ( .B1(n8946), .B2(n9237), .A(n7505), .ZN(n7510) );
  INV_X1 U9215 ( .A(n9053), .ZN(n7817) );
  NAND2_X1 U9216 ( .A1(n7507), .A2(n7817), .ZN(n9068) );
  OAI21_X1 U9217 ( .B1(n7817), .B2(n7507), .A(n9068), .ZN(n7508) );
  AOI222_X1 U9218 ( .A1(n9412), .A2(n7508), .B1(n9224), .B2(n9407), .C1(n8963), 
        .C2(n9409), .ZN(n9319) );
  NOR2_X1 U9219 ( .A1(n9319), .A2(n9430), .ZN(n7509) );
  AOI211_X1 U9220 ( .C1(n9317), .C2(n9229), .A(n7510), .B(n7509), .ZN(n7511)
         );
  OAI21_X1 U9221 ( .B1(n9320), .B2(n9247), .A(n7511), .ZN(P1_U3273) );
  AND2_X1 U9222 ( .A1(n7513), .A2(n7512), .ZN(n7514) );
  NAND2_X1 U9223 ( .A1(n7514), .A2(n7533), .ZN(n7519) );
  INV_X1 U9224 ( .A(n7515), .ZN(n7517) );
  NOR2_X1 U9225 ( .A1(n7517), .A2(n7516), .ZN(n7518) );
  XNOR2_X1 U9226 ( .A(n7519), .B(n7518), .ZN(n7527) );
  OAI21_X1 U9227 ( .B1(n7521), .B2(n8954), .A(n7520), .ZN(n7522) );
  AOI21_X1 U9228 ( .B1(n8940), .B2(n8965), .A(n7522), .ZN(n7523) );
  OAI21_X1 U9229 ( .B1(n7541), .B2(n7524), .A(n7523), .ZN(n7525) );
  AOI21_X1 U9230 ( .B1(n9328), .B2(n8914), .A(n7525), .ZN(n7526) );
  OAI21_X1 U9231 ( .B1(n7527), .B2(n8947), .A(n7526), .ZN(P1_U3224) );
  NAND2_X1 U9232 ( .A1(n7529), .A2(n7528), .ZN(n7531) );
  NAND2_X1 U9233 ( .A1(n7531), .A2(n7530), .ZN(n7532) );
  NAND2_X1 U9234 ( .A1(n7533), .A2(n7532), .ZN(n7534) );
  XOR2_X1 U9235 ( .A(n7535), .B(n7534), .Z(n7544) );
  OAI21_X1 U9236 ( .B1(n7537), .B2(n8954), .A(n7536), .ZN(n7538) );
  AOI21_X1 U9237 ( .B1(n8940), .B2(n8966), .A(n7538), .ZN(n7539) );
  OAI21_X1 U9238 ( .B1(n7541), .B2(n7540), .A(n7539), .ZN(n7542) );
  AOI21_X1 U9239 ( .B1(n9331), .B2(n8914), .A(n7542), .ZN(n7543) );
  OAI21_X1 U9240 ( .B1(n7544), .B2(n8947), .A(n7543), .ZN(P1_U3239) );
  XOR2_X1 U9241 ( .A(n7546), .B(n7545), .Z(n7553) );
  NAND2_X1 U9242 ( .A1(n8964), .A2(n8940), .ZN(n7547) );
  NAND2_X1 U9243 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9000) );
  OAI211_X1 U9244 ( .C1(n8882), .C2(n8954), .A(n7547), .B(n9000), .ZN(n7550)
         );
  NOR2_X1 U9245 ( .A1(n7548), .A2(n8960), .ZN(n7549) );
  AOI211_X1 U9246 ( .C1(n7551), .C2(n8957), .A(n7550), .B(n7549), .ZN(n7552)
         );
  OAI21_X1 U9247 ( .B1(n7553), .B2(n8947), .A(n7552), .ZN(P1_U3226) );
  INV_X1 U9248 ( .A(n7557), .ZN(n7561) );
  XNOR2_X1 U9249 ( .A(n7555), .B(n7554), .ZN(n7558) );
  OAI21_X1 U9250 ( .B1(n7558), .B2(n7557), .A(n7556), .ZN(n7559) );
  OAI21_X1 U9251 ( .B1(n7561), .B2(n7560), .A(n7559), .ZN(n7562) );
  NAND2_X1 U9252 ( .A1(n7562), .A2(n8926), .ZN(n7567) );
  OAI22_X1 U9253 ( .A1(n8952), .A2(n7563), .B1(n6133), .B2(n8954), .ZN(n7564)
         );
  AOI21_X1 U9254 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n7565), .A(n7564), .ZN(
        n7566) );
  OAI211_X1 U9255 ( .C1(n7568), .C2(n8960), .A(n7567), .B(n7566), .ZN(P1_U3220) );
  INV_X1 U9256 ( .A(SI_28_), .ZN(n7571) );
  MUX2_X1 U9257 ( .A(n8855), .B(n8332), .S(n7577), .Z(n7695) );
  INV_X1 U9258 ( .A(SI_29_), .ZN(n7573) );
  AND2_X1 U9259 ( .A1(n7695), .A2(n7573), .ZN(n7576) );
  INV_X1 U9260 ( .A(n7695), .ZN(n7574) );
  NAND2_X1 U9261 ( .A1(n7574), .A2(SI_29_), .ZN(n7575) );
  MUX2_X1 U9262 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7577), .Z(n7578) );
  NAND2_X1 U9263 ( .A1(n7579), .A2(n7578), .ZN(n7580) );
  MUX2_X1 U9264 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7577), .Z(n7581) );
  XNOR2_X1 U9265 ( .A(n7581), .B(SI_31_), .ZN(n7582) );
  NAND2_X1 U9266 ( .A1(n8844), .A2(n5894), .ZN(n7584) );
  NAND2_X1 U9267 ( .A1(n6025), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7583) );
  NAND2_X1 U9268 ( .A1(n8849), .A2(n5894), .ZN(n7587) );
  NAND2_X1 U9269 ( .A1(n6025), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7586) );
  INV_X1 U9270 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9786) );
  NAND2_X1 U9271 ( .A1(n5665), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7590) );
  NAND2_X1 U9272 ( .A1(n7588), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n7589) );
  OAI211_X1 U9273 ( .C1(n5744), .C2(n9786), .A(n7590), .B(n7589), .ZN(n9085)
         );
  INV_X1 U9274 ( .A(n9085), .ZN(n7591) );
  OR2_X1 U9275 ( .A1(n9049), .A2(n7591), .ZN(n7861) );
  OR2_X1 U9276 ( .A1(n9043), .A2(n7861), .ZN(n7595) );
  NAND2_X1 U9277 ( .A1(n5665), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7594) );
  NAND2_X1 U9278 ( .A1(n7588), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U9279 ( .A1(n5641), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7592) );
  AND3_X1 U9280 ( .A1(n7594), .A2(n7593), .A3(n7592), .ZN(n7699) );
  NAND2_X1 U9281 ( .A1(n9248), .A2(n7699), .ZN(n7865) );
  NAND2_X1 U9282 ( .A1(n7595), .A2(n7865), .ZN(n7701) );
  INV_X1 U9283 ( .A(n7701), .ZN(n7776) );
  INV_X1 U9284 ( .A(n7596), .ZN(n7597) );
  NAND2_X1 U9285 ( .A1(n7604), .A2(n7742), .ZN(n7601) );
  MUX2_X1 U9286 ( .A(n7601), .B(n7600), .S(n7704), .Z(n7602) );
  INV_X1 U9287 ( .A(n7602), .ZN(n7603) );
  MUX2_X1 U9288 ( .A(n7604), .B(n7741), .S(n7708), .Z(n7605) );
  AND2_X1 U9289 ( .A1(n7605), .A2(n7801), .ZN(n7606) );
  NAND2_X1 U9290 ( .A1(n7607), .A2(n7606), .ZN(n7613) );
  AND2_X1 U9291 ( .A1(n7845), .A2(n7608), .ZN(n7609) );
  NAND2_X1 U9292 ( .A1(n7611), .A2(n7619), .ZN(n7748) );
  AOI21_X1 U9293 ( .B1(n7613), .B2(n7609), .A(n7748), .ZN(n7615) );
  AND2_X1 U9294 ( .A1(n7611), .A2(n7610), .ZN(n7612) );
  INV_X1 U9295 ( .A(n7845), .ZN(n7761) );
  AOI21_X1 U9296 ( .B1(n7613), .B2(n7612), .A(n7761), .ZN(n7614) );
  AND2_X1 U9297 ( .A1(n7616), .A2(n7621), .ZN(n9373) );
  NAND2_X1 U9298 ( .A1(n9373), .A2(n7617), .ZN(n7731) );
  OAI21_X1 U9299 ( .B1(n7622), .B2(n7731), .A(n7749), .ZN(n7618) );
  NAND2_X1 U9300 ( .A1(n7618), .A2(n7634), .ZN(n7627) );
  NAND2_X1 U9301 ( .A1(n9371), .A2(n7619), .ZN(n7620) );
  AOI21_X1 U9302 ( .B1(n7622), .B2(n7621), .A(n7620), .ZN(n7625) );
  OAI211_X1 U9303 ( .C1(n7625), .C2(n7624), .A(n7752), .B(n7623), .ZN(n7626)
         );
  MUX2_X1 U9304 ( .A(n7627), .B(n7626), .S(n7704), .Z(n7639) );
  INV_X1 U9305 ( .A(n7628), .ZN(n7806) );
  NAND2_X1 U9306 ( .A1(n7640), .A2(n7629), .ZN(n7754) );
  NAND2_X1 U9307 ( .A1(n7752), .A2(n7750), .ZN(n7630) );
  AND2_X1 U9308 ( .A1(n7630), .A2(n7634), .ZN(n7631) );
  NOR2_X1 U9309 ( .A1(n7754), .A2(n7631), .ZN(n7637) );
  NAND2_X1 U9310 ( .A1(n7642), .A2(n7632), .ZN(n7641) );
  NAND2_X1 U9311 ( .A1(n7634), .A2(n7633), .ZN(n7635) );
  AND2_X1 U9312 ( .A1(n7635), .A2(n7752), .ZN(n7636) );
  NOR2_X1 U9313 ( .A1(n7641), .A2(n7636), .ZN(n7730) );
  MUX2_X1 U9314 ( .A(n7637), .B(n7730), .S(n7704), .Z(n7638) );
  OAI21_X1 U9315 ( .B1(n7639), .B2(n7806), .A(n7638), .ZN(n7646) );
  NAND2_X1 U9316 ( .A1(n7641), .A2(n7640), .ZN(n7643) );
  NAND2_X1 U9317 ( .A1(n7754), .A2(n7642), .ZN(n7732) );
  MUX2_X1 U9318 ( .A(n7643), .B(n7732), .S(n7704), .Z(n7644) );
  NAND3_X1 U9319 ( .A1(n7646), .A2(n7645), .A3(n7644), .ZN(n7650) );
  MUX2_X1 U9320 ( .A(n7755), .B(n7647), .S(n7704), .Z(n7648) );
  MUX2_X1 U9321 ( .A(n7651), .B(n7757), .S(n7704), .Z(n7652) );
  NAND2_X1 U9322 ( .A1(n9067), .A2(n7654), .ZN(n7759) );
  INV_X1 U9323 ( .A(n9224), .ZN(n9055) );
  NOR2_X1 U9324 ( .A1(n9312), .A2(n9055), .ZN(n7791) );
  INV_X1 U9325 ( .A(n7791), .ZN(n7660) );
  NAND3_X1 U9326 ( .A1(n7659), .A2(n7657), .A3(n7660), .ZN(n7655) );
  AND2_X1 U9327 ( .A1(n9312), .A2(n9055), .ZN(n7790) );
  INV_X1 U9328 ( .A(n7790), .ZN(n9221) );
  INV_X1 U9329 ( .A(n9242), .ZN(n9204) );
  NAND2_X1 U9330 ( .A1(n9306), .A2(n9204), .ZN(n7789) );
  NAND3_X1 U9331 ( .A1(n7655), .A2(n9221), .A3(n7789), .ZN(n7663) );
  NAND2_X1 U9332 ( .A1(n7657), .A2(n4434), .ZN(n7719) );
  INV_X1 U9333 ( .A(n9067), .ZN(n7658) );
  NOR2_X1 U9334 ( .A1(n7790), .A2(n7658), .ZN(n7718) );
  OR2_X1 U9335 ( .A1(n9306), .A2(n9204), .ZN(n9069) );
  AND2_X1 U9336 ( .A1(n9069), .A2(n7660), .ZN(n7722) );
  NAND2_X1 U9337 ( .A1(n7661), .A2(n7722), .ZN(n7662) );
  MUX2_X1 U9338 ( .A(n7663), .B(n7662), .S(n7704), .Z(n7669) );
  NAND2_X1 U9339 ( .A1(n9303), .A2(n9189), .ZN(n7786) );
  INV_X1 U9340 ( .A(n7786), .ZN(n9071) );
  AOI21_X1 U9341 ( .B1(n7669), .B2(n9069), .A(n9071), .ZN(n7665) );
  INV_X1 U9342 ( .A(n9059), .ZN(n9205) );
  OR2_X1 U9343 ( .A1(n9296), .A2(n9205), .ZN(n7788) );
  NAND2_X1 U9344 ( .A1(n7788), .A2(n7787), .ZN(n7664) );
  NAND2_X1 U9345 ( .A1(n9296), .A2(n9205), .ZN(n9171) );
  INV_X1 U9346 ( .A(n7789), .ZN(n7666) );
  NAND2_X1 U9347 ( .A1(n7787), .A2(n7666), .ZN(n7667) );
  AND2_X1 U9348 ( .A1(n7667), .A2(n7786), .ZN(n7668) );
  AND2_X1 U9349 ( .A1(n9171), .A2(n7668), .ZN(n7763) );
  NAND2_X1 U9350 ( .A1(n7669), .A2(n7763), .ZN(n7672) );
  INV_X1 U9351 ( .A(n7787), .ZN(n7670) );
  NAND2_X1 U9352 ( .A1(n7763), .A2(n7670), .ZN(n7671) );
  AND2_X1 U9353 ( .A1(n7671), .A2(n7788), .ZN(n7717) );
  INV_X1 U9354 ( .A(n9190), .ZN(n9060) );
  NAND2_X1 U9355 ( .A1(n9182), .A2(n9060), .ZN(n9072) );
  NAND2_X1 U9356 ( .A1(n9292), .A2(n9190), .ZN(n7762) );
  OR2_X1 U9357 ( .A1(n9285), .A2(n9175), .ZN(n7785) );
  NAND2_X1 U9358 ( .A1(n9285), .A2(n9175), .ZN(n7784) );
  MUX2_X1 U9359 ( .A(n7785), .B(n7784), .S(n7704), .Z(n7673) );
  NAND2_X1 U9360 ( .A1(n9279), .A2(n9161), .ZN(n9075) );
  NAND2_X1 U9361 ( .A1(n9075), .A2(n7784), .ZN(n7765) );
  INV_X1 U9362 ( .A(n7762), .ZN(n7674) );
  AND2_X1 U9363 ( .A1(n7785), .A2(n7674), .ZN(n7675) );
  NOR2_X1 U9364 ( .A1(n7765), .A2(n7675), .ZN(n7678) );
  INV_X1 U9365 ( .A(n7784), .ZN(n9074) );
  OAI211_X1 U9366 ( .C1(n9074), .C2(n9072), .A(n7783), .B(n7785), .ZN(n7676)
         );
  INV_X1 U9367 ( .A(n7676), .ZN(n7677) );
  MUX2_X1 U9368 ( .A(n7678), .B(n7677), .S(n7704), .Z(n7679) );
  OAI22_X1 U9369 ( .A1(n7688), .A2(n9275), .B1(n7708), .B2(n9075), .ZN(n7680)
         );
  NAND2_X1 U9370 ( .A1(n7680), .A2(n9121), .ZN(n7683) );
  INV_X1 U9371 ( .A(n9121), .ZN(n9150) );
  AOI21_X1 U9372 ( .B1(n9131), .B2(n9076), .A(n9150), .ZN(n7681) );
  MUX2_X1 U9373 ( .A(n9131), .B(n7681), .S(n7708), .Z(n7682) );
  NAND2_X1 U9374 ( .A1(n7683), .A2(n7682), .ZN(n7690) );
  OAI21_X1 U9375 ( .B1(n9131), .B2(n9076), .A(n7767), .ZN(n7686) );
  NAND2_X1 U9376 ( .A1(n9075), .A2(n9150), .ZN(n7684) );
  NAND2_X1 U9377 ( .A1(n9079), .A2(n7684), .ZN(n7685) );
  MUX2_X1 U9378 ( .A(n7686), .B(n7685), .S(n7704), .Z(n7687) );
  OAI21_X1 U9379 ( .B1(n7688), .B2(n9118), .A(n7687), .ZN(n7689) );
  NAND2_X1 U9380 ( .A1(n9264), .A2(n9120), .ZN(n7770) );
  INV_X1 U9381 ( .A(n9103), .ZN(n7692) );
  MUX2_X1 U9382 ( .A(n7767), .B(n9079), .S(n7708), .Z(n7691) );
  MUX2_X1 U9383 ( .A(n7770), .B(n9081), .S(n7704), .Z(n7693) );
  XNOR2_X1 U9384 ( .A(n7695), .B(SI_29_), .ZN(n7696) );
  NAND2_X1 U9385 ( .A1(n8330), .A2(n5894), .ZN(n7698) );
  NAND2_X1 U9386 ( .A1(n6025), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7697) );
  INV_X1 U9387 ( .A(n7699), .ZN(n9041) );
  NAND2_X1 U9388 ( .A1(n9041), .A2(n9085), .ZN(n7700) );
  NAND2_X1 U9389 ( .A1(n9049), .A2(n7700), .ZN(n7773) );
  NAND2_X1 U9390 ( .A1(n7706), .A2(n9105), .ZN(n7703) );
  MUX2_X1 U9391 ( .A(n7704), .B(n7703), .S(n9091), .Z(n7705) );
  OAI211_X1 U9392 ( .C1(n9105), .C2(n7708), .A(n7776), .B(n7705), .ZN(n7711)
         );
  INV_X1 U9393 ( .A(n7706), .ZN(n7709) );
  NAND3_X1 U9394 ( .A1(n7709), .A2(n7708), .A3(n7707), .ZN(n7710) );
  NAND2_X1 U9395 ( .A1(n7711), .A2(n7710), .ZN(n7712) );
  AOI21_X1 U9396 ( .B1(n7712), .B2(n7773), .A(n7779), .ZN(n7713) );
  NOR2_X1 U9397 ( .A1(n7777), .A2(n9033), .ZN(n7827) );
  INV_X1 U9398 ( .A(n7827), .ZN(n7715) );
  INV_X1 U9399 ( .A(n7717), .ZN(n7728) );
  INV_X1 U9400 ( .A(n7763), .ZN(n7726) );
  INV_X1 U9401 ( .A(n7718), .ZN(n7721) );
  INV_X1 U9402 ( .A(n7719), .ZN(n7720) );
  NOR2_X1 U9403 ( .A1(n7721), .A2(n7720), .ZN(n7724) );
  INV_X1 U9404 ( .A(n7722), .ZN(n7723) );
  NOR2_X1 U9405 ( .A1(n7724), .A2(n7723), .ZN(n7725) );
  NOR2_X1 U9406 ( .A1(n7726), .A2(n7725), .ZN(n7727) );
  OAI21_X1 U9407 ( .B1(n7728), .B2(n7727), .A(n7762), .ZN(n7729) );
  NAND3_X1 U9408 ( .A1(n7729), .A2(n9072), .A3(n7785), .ZN(n7851) );
  INV_X1 U9409 ( .A(n7730), .ZN(n7734) );
  AND4_X1 U9410 ( .A1(n7752), .A2(n7750), .A3(n7749), .A4(n7731), .ZN(n7733)
         );
  OAI211_X1 U9411 ( .C1(n7734), .C2(n7733), .A(n7755), .B(n7732), .ZN(n7735)
         );
  NAND2_X1 U9412 ( .A1(n7736), .A2(n7735), .ZN(n7737) );
  NAND2_X1 U9413 ( .A1(n7737), .A2(n7757), .ZN(n7738) );
  OR2_X1 U9414 ( .A1(n7759), .A2(n7738), .ZN(n7847) );
  NAND2_X1 U9415 ( .A1(n7742), .A2(n7739), .ZN(n7740) );
  NOR2_X1 U9416 ( .A1(n7841), .A2(n7740), .ZN(n7840) );
  INV_X1 U9417 ( .A(n7741), .ZN(n7743) );
  NOR3_X1 U9418 ( .A1(n7744), .A2(n7743), .A3(n7742), .ZN(n7745) );
  AOI211_X1 U9419 ( .C1(n7842), .C2(n7836), .A(n7841), .B(n7745), .ZN(n7746)
         );
  AOI21_X1 U9420 ( .B1(n7840), .B2(n7747), .A(n7746), .ZN(n7760) );
  INV_X1 U9421 ( .A(n7748), .ZN(n7751) );
  NAND4_X1 U9422 ( .A1(n7752), .A2(n7751), .A3(n7750), .A4(n7749), .ZN(n7753)
         );
  NOR2_X1 U9423 ( .A1(n7754), .A2(n7753), .ZN(n7756) );
  NAND3_X1 U9424 ( .A1(n7757), .A2(n7756), .A3(n7755), .ZN(n7758) );
  NOR2_X1 U9425 ( .A1(n7759), .A2(n7758), .ZN(n7850) );
  OAI21_X1 U9426 ( .B1(n7761), .B2(n7760), .A(n7850), .ZN(n7764) );
  NAND3_X1 U9427 ( .A1(n7763), .A2(n9221), .A3(n7762), .ZN(n7853) );
  AOI21_X1 U9428 ( .B1(n7847), .B2(n7764), .A(n7853), .ZN(n7766) );
  INV_X1 U9429 ( .A(n7765), .ZN(n7856) );
  OAI21_X1 U9430 ( .B1(n7851), .B2(n7766), .A(n7856), .ZN(n7771) );
  NAND2_X1 U9431 ( .A1(n9275), .A2(n9121), .ZN(n7782) );
  NAND2_X1 U9432 ( .A1(n7767), .A2(n7782), .ZN(n7768) );
  NAND2_X1 U9433 ( .A1(n7768), .A2(n9079), .ZN(n7769) );
  NAND2_X1 U9434 ( .A1(n7770), .A2(n7769), .ZN(n7859) );
  AOI21_X1 U9435 ( .B1(n9079), .B2(n7771), .A(n7859), .ZN(n7774) );
  AND2_X1 U9436 ( .A1(n9077), .A2(n7783), .ZN(n7772) );
  OAI211_X1 U9437 ( .C1(n7859), .C2(n7772), .A(n7781), .B(n9081), .ZN(n7857)
         );
  NAND2_X1 U9438 ( .A1(n9258), .A2(n9105), .ZN(n7864) );
  OAI211_X1 U9439 ( .C1(n7774), .C2(n7857), .A(n7773), .B(n7864), .ZN(n7775)
         );
  AOI211_X1 U9440 ( .C1(n7776), .C2(n7775), .A(n7823), .B(n7779), .ZN(n7778)
         );
  NOR3_X1 U9441 ( .A1(n7778), .A2(n9211), .A3(n7777), .ZN(n7826) );
  INV_X1 U9442 ( .A(n9049), .ZN(n9254) );
  INV_X1 U9443 ( .A(n7779), .ZN(n7780) );
  OAI21_X1 U9444 ( .B1(n9254), .B2(n9085), .A(n7780), .ZN(n7866) );
  INV_X1 U9445 ( .A(n9148), .ZN(n7820) );
  NAND2_X1 U9446 ( .A1(n7785), .A2(n7784), .ZN(n9158) );
  INV_X1 U9447 ( .A(n9158), .ZN(n9155) );
  INV_X1 U9448 ( .A(n9172), .ZN(n9169) );
  NAND2_X1 U9449 ( .A1(n7788), .A2(n9171), .ZN(n9187) );
  NOR2_X1 U9450 ( .A1(n7791), .A2(n7790), .ZN(n9241) );
  INV_X1 U9451 ( .A(n9418), .ZN(n7810) );
  INV_X1 U9452 ( .A(n7792), .ZN(n7796) );
  NAND4_X1 U9453 ( .A1(n7796), .A2(n7795), .A3(n7794), .A4(n7793), .ZN(n7800)
         );
  INV_X1 U9454 ( .A(n7797), .ZN(n7798) );
  NOR3_X1 U9455 ( .A1(n7800), .A2(n7799), .A3(n7798), .ZN(n7804) );
  NAND4_X1 U9456 ( .A1(n7804), .A2(n7803), .A3(n7802), .A4(n7801), .ZN(n7807)
         );
  NOR4_X1 U9457 ( .A1(n7807), .A2(n7806), .A3(n9380), .A4(n7805), .ZN(n7808)
         );
  NAND4_X1 U9458 ( .A1(n7811), .A2(n7810), .A3(n7809), .A4(n7808), .ZN(n7812)
         );
  NOR4_X1 U9459 ( .A1(n7815), .A2(n7814), .A3(n7813), .A4(n7812), .ZN(n7816)
         );
  NAND4_X1 U9460 ( .A1(n9222), .A2(n7817), .A3(n9241), .A4(n7816), .ZN(n7818)
         );
  NOR4_X1 U9461 ( .A1(n9169), .A2(n9201), .A3(n9187), .A4(n7818), .ZN(n7819)
         );
  NAND3_X1 U9462 ( .A1(n7820), .A2(n9155), .A3(n7819), .ZN(n7821) );
  NOR4_X1 U9463 ( .A1(n9103), .A2(n9118), .A3(n9133), .A4(n7821), .ZN(n7822)
         );
  NAND4_X1 U9464 ( .A1(n7861), .A2(n9082), .A3(n7822), .A4(n7865), .ZN(n7824)
         );
  OAI21_X1 U9465 ( .B1(n7866), .B2(n7824), .A(n7823), .ZN(n7825) );
  INV_X1 U9466 ( .A(n7828), .ZN(n7835) );
  INV_X1 U9467 ( .A(n7829), .ZN(n7830) );
  OAI211_X1 U9468 ( .C1(n7832), .C2(n7831), .A(n6060), .B(n7830), .ZN(n7833)
         );
  NAND3_X1 U9469 ( .A1(n7835), .A2(n7834), .A3(n7833), .ZN(n7839) );
  INV_X1 U9470 ( .A(n7836), .ZN(n7837) );
  AOI21_X1 U9471 ( .B1(n7839), .B2(n7838), .A(n7837), .ZN(n7844) );
  INV_X1 U9472 ( .A(n7840), .ZN(n7843) );
  OAI22_X1 U9473 ( .A1(n7844), .A2(n7843), .B1(n7842), .B2(n7841), .ZN(n7846)
         );
  NAND2_X1 U9474 ( .A1(n7846), .A2(n7845), .ZN(n7849) );
  INV_X1 U9475 ( .A(n7847), .ZN(n7848) );
  AOI21_X1 U9476 ( .B1(n7850), .B2(n7849), .A(n7848), .ZN(n7854) );
  INV_X1 U9477 ( .A(n7851), .ZN(n7852) );
  OAI21_X1 U9478 ( .B1(n7854), .B2(n7853), .A(n7852), .ZN(n7855) );
  AOI21_X1 U9479 ( .B1(n7856), .B2(n7855), .A(n9118), .ZN(n7860) );
  INV_X1 U9480 ( .A(n7857), .ZN(n7858) );
  OAI21_X1 U9481 ( .B1(n7860), .B2(n7859), .A(n7858), .ZN(n7863) );
  INV_X1 U9482 ( .A(n7861), .ZN(n7862) );
  AOI21_X1 U9483 ( .B1(n7864), .B2(n7863), .A(n7862), .ZN(n7867) );
  OAI21_X1 U9484 ( .B1(n7867), .B2(n7866), .A(n7865), .ZN(n7868) );
  XNOR2_X1 U9485 ( .A(n7868), .B(n9033), .ZN(n7870) );
  NOR2_X1 U9486 ( .A1(n7870), .A2(n7869), .ZN(n7871) );
  NAND2_X1 U9487 ( .A1(n7873), .A2(n9039), .ZN(n7874) );
  OAI211_X1 U9488 ( .C1(n7875), .C2(n7877), .A(n7874), .B(P1_B_REG_SCAN_IN), 
        .ZN(n7876) );
  OAI21_X1 U9489 ( .B1(n7878), .B2(n7877), .A(n7876), .ZN(P1_U3240) );
  NAND2_X1 U9490 ( .A1(n7880), .A2(n7879), .ZN(n7882) );
  XNOR2_X1 U9491 ( .A(n8016), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n7881) );
  NAND2_X1 U9492 ( .A1(n7881), .A2(n7882), .ZN(n8015) );
  OAI211_X1 U9493 ( .C1(n7882), .C2(n7881), .A(n8454), .B(n8015), .ZN(n7894)
         );
  INV_X1 U9494 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7883) );
  XNOR2_X1 U9495 ( .A(n8016), .B(n7883), .ZN(n7888) );
  OR2_X1 U9496 ( .A1(n7884), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U9497 ( .A1(n7886), .A2(n7885), .ZN(n7887) );
  NOR2_X1 U9498 ( .A1(n7888), .A2(n7887), .ZN(n8019) );
  AOI21_X1 U9499 ( .B1(n7888), .B2(n7887), .A(n8019), .ZN(n7892) );
  INV_X1 U9500 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7890) );
  OR2_X1 U9501 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5204), .ZN(n7889) );
  OAI21_X1 U9502 ( .B1(n8460), .B2(n7890), .A(n7889), .ZN(n7891) );
  AOI21_X1 U9503 ( .B1(n8453), .B2(n7892), .A(n7891), .ZN(n7893) );
  OAI211_X1 U9504 ( .C1(n8448), .C2(n8016), .A(n7894), .B(n7893), .ZN(P2_U3262) );
  AOI21_X1 U9505 ( .B1(n7897), .B2(n7896), .A(n7895), .ZN(n7898) );
  OR2_X1 U9506 ( .A1(n7898), .A2(n8450), .ZN(n7907) );
  OAI21_X1 U9507 ( .B1(n7901), .B2(n7900), .A(n7899), .ZN(n7905) );
  INV_X1 U9508 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7903) );
  OAI21_X1 U9509 ( .B1(n8460), .B2(n7903), .A(n7902), .ZN(n7904) );
  AOI21_X1 U9510 ( .B1(n8453), .B2(n7905), .A(n7904), .ZN(n7906) );
  OAI211_X1 U9511 ( .C1(n8448), .C2(n7908), .A(n7907), .B(n7906), .ZN(P2_U3258) );
  OAI21_X1 U9512 ( .B1(n7911), .B2(n7910), .A(n7909), .ZN(n7916) );
  INV_X1 U9513 ( .A(n7912), .ZN(n7915) );
  INV_X1 U9514 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7913) );
  NOR2_X1 U9515 ( .A1(n8460), .A2(n7913), .ZN(n7914) );
  AOI211_X1 U9516 ( .C1(n8453), .C2(n7916), .A(n7915), .B(n7914), .ZN(n7923)
         );
  MUX2_X1 U9517 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7918), .S(n7917), .Z(n7920)
         );
  OAI211_X1 U9518 ( .C1(n7921), .C2(n7920), .A(n8454), .B(n7919), .ZN(n7922)
         );
  OAI211_X1 U9519 ( .C1(n8448), .C2(n7924), .A(n7923), .B(n7922), .ZN(P2_U3257) );
  OAI211_X1 U9520 ( .C1(n7927), .C2(n7926), .A(n8454), .B(n7925), .ZN(n7937)
         );
  AOI21_X1 U9521 ( .B1(n7930), .B2(n7929), .A(n7928), .ZN(n7935) );
  INV_X1 U9522 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7933) );
  OR2_X1 U9523 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7931), .ZN(n7932) );
  OAI21_X1 U9524 ( .B1(n8460), .B2(n7933), .A(n7932), .ZN(n7934) );
  AOI21_X1 U9525 ( .B1(n8453), .B2(n7935), .A(n7934), .ZN(n7936) );
  OAI211_X1 U9526 ( .C1(n8448), .C2(n7938), .A(n7937), .B(n7936), .ZN(P2_U3255) );
  INV_X1 U9527 ( .A(n7939), .ZN(n7944) );
  AOI211_X1 U9528 ( .C1(n7942), .C2(n7941), .A(n7940), .B(n8087), .ZN(n7943)
         );
  AOI211_X1 U9529 ( .C1(n8079), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7944), .B(
        n7943), .ZN(n7949) );
  OAI211_X1 U9530 ( .C1(n7947), .C2(n7946), .A(n8454), .B(n7945), .ZN(n7948)
         );
  OAI211_X1 U9531 ( .C1(n8448), .C2(n7950), .A(n7949), .B(n7948), .ZN(P2_U3254) );
  INV_X1 U9532 ( .A(n7951), .ZN(n7956) );
  AOI211_X1 U9533 ( .C1(n7954), .C2(n7953), .A(n7952), .B(n8087), .ZN(n7955)
         );
  AOI211_X1 U9534 ( .C1(n8079), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7956), .B(
        n7955), .ZN(n7961) );
  OAI211_X1 U9535 ( .C1(n7959), .C2(n7958), .A(n8454), .B(n7957), .ZN(n7960)
         );
  OAI211_X1 U9536 ( .C1(n8448), .C2(n7962), .A(n7961), .B(n7960), .ZN(P2_U3253) );
  NOR2_X1 U9537 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7963), .ZN(n7968) );
  AOI211_X1 U9538 ( .C1(n7966), .C2(n7965), .A(n7964), .B(n8087), .ZN(n7967)
         );
  AOI211_X1 U9539 ( .C1(n8079), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n7968), .B(
        n7967), .ZN(n7973) );
  OAI211_X1 U9540 ( .C1(n7971), .C2(n7970), .A(n8454), .B(n7969), .ZN(n7972)
         );
  OAI211_X1 U9541 ( .C1(n8448), .C2(n7974), .A(n7973), .B(n7972), .ZN(P2_U3252) );
  INV_X1 U9542 ( .A(n7975), .ZN(n7979) );
  AOI211_X1 U9543 ( .C1(n4275), .C2(n7977), .A(n7976), .B(n8087), .ZN(n7978)
         );
  AOI211_X1 U9544 ( .C1(n8079), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n7979), .B(
        n7978), .ZN(n7984) );
  OAI211_X1 U9545 ( .C1(n7982), .C2(n7981), .A(n8454), .B(n7980), .ZN(n7983)
         );
  OAI211_X1 U9546 ( .C1(n8448), .C2(n7985), .A(n7984), .B(n7983), .ZN(P2_U3251) );
  INV_X1 U9547 ( .A(n7986), .ZN(n7991) );
  AOI211_X1 U9548 ( .C1(n7989), .C2(n7988), .A(n7987), .B(n8087), .ZN(n7990)
         );
  AOI211_X1 U9549 ( .C1(n8079), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7991), .B(
        n7990), .ZN(n7998) );
  INV_X1 U9550 ( .A(n7992), .ZN(n7996) );
  NAND3_X1 U9551 ( .A1(n8009), .A2(n7994), .A3(n7993), .ZN(n7995) );
  NAND3_X1 U9552 ( .A1(n8454), .A2(n7996), .A3(n7995), .ZN(n7997) );
  OAI211_X1 U9553 ( .C1(n8448), .C2(n7999), .A(n7998), .B(n7997), .ZN(P2_U3249) );
  NOR2_X1 U9554 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8717), .ZN(n8004) );
  AOI211_X1 U9555 ( .C1(n8002), .C2(n8001), .A(n8000), .B(n8087), .ZN(n8003)
         );
  AOI211_X1 U9556 ( .C1(n8079), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n8004), .B(
        n8003), .ZN(n8013) );
  INV_X1 U9557 ( .A(n8005), .ZN(n8008) );
  MUX2_X1 U9558 ( .A(n7338), .B(P2_REG2_REG_3__SCAN_IN), .S(n8006), .Z(n8007)
         );
  NAND2_X1 U9559 ( .A1(n8008), .A2(n8007), .ZN(n8010) );
  OAI211_X1 U9560 ( .C1(n8011), .C2(n8010), .A(n8454), .B(n8009), .ZN(n8012)
         );
  OAI211_X1 U9561 ( .C1(n8448), .C2(n8014), .A(n8013), .B(n8012), .ZN(P2_U3248) );
  INV_X1 U9562 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8017) );
  OAI21_X1 U9563 ( .B1(n8017), .B2(n8016), .A(n8015), .ZN(n8441) );
  XNOR2_X1 U9564 ( .A(n8446), .B(n8441), .ZN(n8018) );
  NOR2_X1 U9565 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8018), .ZN(n8443) );
  AOI21_X1 U9566 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8018), .A(n8443), .ZN(
        n8030) );
  INV_X1 U9567 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8021) );
  AOI22_X1 U9568 ( .A1(n8446), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8021), .B2(
        n8026), .ZN(n8022) );
  OAI21_X1 U9569 ( .B1(n8023), .B2(n8022), .A(n8445), .ZN(n8028) );
  NAND2_X1 U9570 ( .A1(n8079), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8024) );
  OAI211_X1 U9571 ( .C1(n8448), .C2(n8026), .A(n8025), .B(n8024), .ZN(n8027)
         );
  AOI21_X1 U9572 ( .B1(n8028), .B2(n8453), .A(n8027), .ZN(n8029) );
  OAI21_X1 U9573 ( .B1(n8030), .B2(n8450), .A(n8029), .ZN(P2_U3263) );
  AOI21_X1 U9574 ( .B1(n8032), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8031), .ZN(
        n8043) );
  AOI211_X1 U9575 ( .C1(n8035), .C2(n8034), .A(n8033), .B(n8087), .ZN(n8041)
         );
  INV_X1 U9576 ( .A(n8036), .ZN(n8037) );
  AOI21_X1 U9577 ( .B1(n8079), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8037), .ZN(
        n8038) );
  OAI21_X1 U9578 ( .B1(n8448), .B2(n8039), .A(n8038), .ZN(n8040) );
  NOR2_X1 U9579 ( .A1(n8041), .A2(n8040), .ZN(n8042) );
  OAI21_X1 U9580 ( .B1(n8043), .B2(n8450), .A(n8042), .ZN(P2_U3260) );
  AOI21_X1 U9581 ( .B1(n8046), .B2(n8045), .A(n8044), .ZN(n8056) );
  OAI21_X1 U9582 ( .B1(n8049), .B2(n8048), .A(n8047), .ZN(n8050) );
  NAND2_X1 U9583 ( .A1(n8050), .A2(n8453), .ZN(n8055) );
  INV_X1 U9584 ( .A(n8448), .ZN(n8094) );
  INV_X1 U9585 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n9861) );
  OAI21_X1 U9586 ( .B1(n8460), .B2(n9861), .A(n8051), .ZN(n8052) );
  AOI21_X1 U9587 ( .B1(n8094), .B2(n8053), .A(n8052), .ZN(n8054) );
  OAI211_X1 U9588 ( .C1(n8056), .C2(n8450), .A(n8055), .B(n8054), .ZN(P2_U3259) );
  AOI21_X1 U9589 ( .B1(n8059), .B2(n8058), .A(n8057), .ZN(n8070) );
  AOI21_X1 U9590 ( .B1(n8062), .B2(n8061), .A(n8060), .ZN(n8063) );
  NAND2_X1 U9591 ( .A1(n8453), .A2(n8063), .ZN(n8066) );
  NOR2_X1 U9592 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5102), .ZN(n8064) );
  AOI21_X1 U9593 ( .B1(n8079), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8064), .ZN(
        n8065) );
  OAI211_X1 U9594 ( .C1(n8448), .C2(n8067), .A(n8066), .B(n8065), .ZN(n8068)
         );
  INV_X1 U9595 ( .A(n8068), .ZN(n8069) );
  OAI21_X1 U9596 ( .B1(n8070), .B2(n8450), .A(n8069), .ZN(P2_U3256) );
  XNOR2_X1 U9597 ( .A(n8072), .B(n8071), .ZN(n8083) );
  NOR2_X1 U9598 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8073), .ZN(n8078) );
  AOI211_X1 U9599 ( .C1(n8076), .C2(n8075), .A(n8087), .B(n8074), .ZN(n8077)
         );
  AOI211_X1 U9600 ( .C1(n8079), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n8078), .B(
        n8077), .ZN(n8082) );
  NAND2_X1 U9601 ( .A1(n8094), .A2(n8080), .ZN(n8081) );
  OAI211_X1 U9602 ( .C1(n8083), .C2(n8450), .A(n8082), .B(n8081), .ZN(P2_U3250) );
  XNOR2_X1 U9603 ( .A(n8085), .B(n8084), .ZN(n8096) );
  OAI22_X1 U9604 ( .A1(n8460), .A2(n9720), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8086), .ZN(n8092) );
  AOI211_X1 U9605 ( .C1(n8090), .C2(n8089), .A(n8088), .B(n8087), .ZN(n8091)
         );
  AOI211_X1 U9606 ( .C1(n8094), .C2(n8093), .A(n8092), .B(n8091), .ZN(n8095)
         );
  OAI21_X1 U9607 ( .B1(n8450), .B2(n8096), .A(n8095), .ZN(P2_U3246) );
  OAI222_X1 U9608 ( .A1(n8856), .A2(n8099), .B1(n8098), .B2(n8097), .C1(n6366), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  NOR2_X1 U9609 ( .A1(n8792), .A2(n8475), .ZN(n8130) );
  NOR2_X1 U9610 ( .A1(n8130), .A2(n8222), .ZN(n8676) );
  INV_X1 U9611 ( .A(n8222), .ZN(n8101) );
  NOR2_X1 U9612 ( .A1(n8788), .A2(n8477), .ZN(n8224) );
  NAND2_X1 U9613 ( .A1(n8660), .A2(n8661), .ZN(n8659) );
  INV_X1 U9614 ( .A(n8223), .ZN(n8102) );
  NAND2_X1 U9615 ( .A1(n8659), .A2(n8102), .ZN(n8644) );
  NAND2_X1 U9616 ( .A1(n8783), .A2(n8480), .ZN(n8227) );
  NOR2_X2 U9617 ( .A1(n8644), .A2(n8645), .ZN(n8642) );
  OR2_X1 U9618 ( .A1(n8777), .A2(n8610), .ZN(n8228) );
  NAND2_X1 U9619 ( .A1(n8777), .A2(n8610), .ZN(n8605) );
  NAND2_X1 U9620 ( .A1(n8228), .A2(n8605), .ZN(n8625) );
  INV_X1 U9621 ( .A(n8229), .ZN(n8626) );
  NAND2_X1 U9622 ( .A1(n8774), .A2(n8593), .ZN(n8221) );
  NAND2_X1 U9623 ( .A1(n8234), .A2(n8221), .ZN(n8483) );
  NAND2_X1 U9624 ( .A1(n8607), .A2(n8605), .ZN(n8105) );
  NAND2_X1 U9625 ( .A1(n8601), .A2(n8580), .ZN(n8239) );
  INV_X1 U9626 ( .A(n8580), .ZN(n8611) );
  NAND2_X1 U9627 ( .A1(n8761), .A2(n8592), .ZN(n8245) );
  NAND2_X1 U9628 ( .A1(n8579), .A2(n8578), .ZN(n8577) );
  NOR2_X1 U9629 ( .A1(n8758), .A2(n8424), .ZN(n8247) );
  INV_X1 U9630 ( .A(n8530), .ZN(n8106) );
  NOR2_X1 U9631 ( .A1(n8746), .A2(n8415), .ZN(n8257) );
  NAND2_X1 U9632 ( .A1(n8741), .A2(n8423), .ZN(n8107) );
  INV_X1 U9633 ( .A(n8423), .ZN(n8531) );
  NAND2_X1 U9634 ( .A1(n8330), .A2(n8116), .ZN(n8109) );
  NAND2_X1 U9635 ( .A1(n4252), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8108) );
  INV_X1 U9636 ( .A(n8268), .ZN(n8111) );
  NAND2_X1 U9637 ( .A1(n8499), .A2(n8110), .ZN(n8269) );
  NAND2_X1 U9638 ( .A1(n8849), .A2(n8116), .ZN(n8113) );
  NAND2_X1 U9639 ( .A1(n4252), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8112) );
  NOR2_X1 U9640 ( .A1(n8470), .A2(n8494), .ZN(n8125) );
  NAND2_X1 U9641 ( .A1(n8844), .A2(n8116), .ZN(n8118) );
  NAND2_X1 U9642 ( .A1(n4253), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U9643 ( .A1(n8470), .A2(n8494), .ZN(n8272) );
  NAND2_X1 U9644 ( .A1(n8273), .A2(n8272), .ZN(n8123) );
  NAND2_X1 U9645 ( .A1(n8727), .A2(n8465), .ZN(n8124) );
  OAI21_X1 U9646 ( .B1(n8119), .B2(n8123), .A(n8124), .ZN(n8120) );
  XNOR2_X1 U9647 ( .A(n8120), .B(n8567), .ZN(n8323) );
  NAND2_X1 U9648 ( .A1(n8122), .A2(n8121), .ZN(n8322) );
  INV_X1 U9649 ( .A(n8123), .ZN(n8311) );
  INV_X1 U9650 ( .A(n8124), .ZN(n8276) );
  NOR2_X1 U9651 ( .A1(n8276), .A2(n8125), .ZN(n8313) );
  OR2_X1 U9652 ( .A1(n8280), .A2(n4864), .ZN(n8274) );
  MUX2_X1 U9653 ( .A(n8311), .B(n8313), .S(n8274), .Z(n8279) );
  INV_X1 U9654 ( .A(n8490), .ZN(n8312) );
  INV_X1 U9655 ( .A(n8510), .ZN(n8262) );
  INV_X1 U9656 ( .A(n8126), .ZN(n8127) );
  NOR2_X1 U9657 ( .A1(n8222), .A2(n8127), .ZN(n8128) );
  MUX2_X1 U9658 ( .A(n8129), .B(n8128), .S(n8267), .Z(n8215) );
  INV_X1 U9659 ( .A(n8130), .ZN(n8216) );
  AND2_X1 U9660 ( .A1(n8133), .A2(n8689), .ZN(n8131) );
  MUX2_X1 U9661 ( .A(n8687), .B(n8131), .S(n8267), .Z(n8155) );
  NAND2_X1 U9662 ( .A1(n8133), .A2(n8132), .ZN(n8135) );
  NAND2_X1 U9663 ( .A1(n8160), .A2(n8689), .ZN(n8134) );
  AOI21_X1 U9664 ( .B1(n8155), .B2(n8135), .A(n8134), .ZN(n8149) );
  NAND2_X1 U9665 ( .A1(n8140), .A2(n8139), .ZN(n8283) );
  NAND3_X1 U9666 ( .A1(n8283), .A2(n8142), .A3(n8136), .ZN(n8138) );
  NAND2_X1 U9667 ( .A1(n8138), .A2(n8137), .ZN(n8145) );
  AND2_X1 U9668 ( .A1(n8139), .A2(n8315), .ZN(n8141) );
  OAI211_X1 U9669 ( .C1(n6444), .C2(n8141), .A(n8137), .B(n8140), .ZN(n8143)
         );
  NAND2_X1 U9670 ( .A1(n8143), .A2(n8142), .ZN(n8144) );
  MUX2_X1 U9671 ( .A(n8145), .B(n8144), .S(n8274), .Z(n8147) );
  NAND3_X1 U9672 ( .A1(n8147), .A2(n8155), .A3(n8146), .ZN(n8148) );
  OAI21_X1 U9673 ( .B1(n8267), .B2(n8149), .A(n8148), .ZN(n8150) );
  NAND2_X1 U9674 ( .A1(n8150), .A2(n8156), .ZN(n8163) );
  INV_X1 U9675 ( .A(n8151), .ZN(n8154) );
  NAND2_X1 U9676 ( .A1(n8687), .A2(n8152), .ZN(n8153) );
  OAI21_X1 U9677 ( .B1(n8155), .B2(n8154), .A(n8153), .ZN(n8157) );
  NAND2_X1 U9678 ( .A1(n8157), .A2(n8156), .ZN(n8158) );
  NAND2_X1 U9679 ( .A1(n8158), .A2(n8267), .ZN(n8162) );
  OAI21_X1 U9680 ( .B1(n8160), .B2(n8274), .A(n8159), .ZN(n8161) );
  AOI21_X1 U9681 ( .B1(n8163), .B2(n8162), .A(n8161), .ZN(n8168) );
  MUX2_X1 U9682 ( .A(n8165), .B(n8164), .S(n8274), .Z(n8166) );
  NAND2_X1 U9683 ( .A1(n8294), .A2(n8166), .ZN(n8167) );
  OR2_X1 U9684 ( .A1(n8168), .A2(n8167), .ZN(n8175) );
  MUX2_X1 U9685 ( .A(n8170), .B(n8169), .S(n8267), .Z(n8171) );
  INV_X1 U9686 ( .A(n8171), .ZN(n8172) );
  NOR2_X1 U9687 ( .A1(n8173), .A2(n8172), .ZN(n8174) );
  NAND2_X1 U9688 ( .A1(n8175), .A2(n8174), .ZN(n8180) );
  INV_X1 U9689 ( .A(n8178), .ZN(n8176) );
  NAND2_X1 U9690 ( .A1(n8180), .A2(n8176), .ZN(n8177) );
  NAND3_X1 U9691 ( .A1(n8177), .A2(n8185), .A3(n8181), .ZN(n8184) );
  AOI21_X1 U9692 ( .B1(n8180), .B2(n8179), .A(n8178), .ZN(n8182) );
  OAI21_X1 U9693 ( .B1(n8182), .B2(n4649), .A(n8187), .ZN(n8183) );
  MUX2_X1 U9694 ( .A(n8184), .B(n8183), .S(n8274), .Z(n8195) );
  NAND2_X1 U9695 ( .A1(n8189), .A2(n8185), .ZN(n8186) );
  NAND2_X1 U9696 ( .A1(n8186), .A2(n8188), .ZN(n8192) );
  NAND2_X1 U9697 ( .A1(n8188), .A2(n8187), .ZN(n8190) );
  NAND2_X1 U9698 ( .A1(n8190), .A2(n8189), .ZN(n8191) );
  MUX2_X1 U9699 ( .A(n8192), .B(n8191), .S(n8267), .Z(n8193) );
  OAI211_X1 U9700 ( .C1(n8195), .C2(n8299), .A(n8194), .B(n8193), .ZN(n8199)
         );
  MUX2_X1 U9701 ( .A(n8197), .B(n8196), .S(n8267), .Z(n8198) );
  NAND3_X1 U9702 ( .A1(n8199), .A2(n8301), .A3(n8198), .ZN(n8204) );
  OR2_X1 U9703 ( .A1(n8812), .A2(n8274), .ZN(n8202) );
  NAND2_X1 U9704 ( .A1(n8812), .A2(n8274), .ZN(n8201) );
  MUX2_X1 U9705 ( .A(n8202), .B(n8201), .S(n8200), .Z(n8203) );
  NAND3_X1 U9706 ( .A1(n8204), .A2(n8303), .A3(n8203), .ZN(n8208) );
  MUX2_X1 U9707 ( .A(n8206), .B(n8205), .S(n8267), .Z(n8207) );
  NAND3_X1 U9708 ( .A1(n8208), .A2(n8304), .A3(n8207), .ZN(n8212) );
  MUX2_X1 U9709 ( .A(n8210), .B(n8209), .S(n8274), .Z(n8211) );
  NAND3_X1 U9710 ( .A1(n8212), .A2(n8306), .A3(n8211), .ZN(n8213) );
  AND2_X1 U9711 ( .A1(n8216), .A2(n8213), .ZN(n8214) );
  NAND2_X1 U9712 ( .A1(n8215), .A2(n8214), .ZN(n8226) );
  AOI21_X1 U9713 ( .B1(n8226), .B2(n8216), .A(n8223), .ZN(n8219) );
  INV_X1 U9714 ( .A(n8224), .ZN(n8217) );
  NAND2_X1 U9715 ( .A1(n8229), .A2(n8217), .ZN(n8218) );
  OAI211_X1 U9716 ( .C1(n8219), .C2(n8218), .A(n8227), .B(n8605), .ZN(n8220)
         );
  NAND4_X1 U9717 ( .A1(n8220), .A2(n8234), .A3(n8267), .A4(n8228), .ZN(n8243)
         );
  INV_X1 U9718 ( .A(n8221), .ZN(n8236) );
  NOR2_X1 U9719 ( .A1(n8223), .A2(n8222), .ZN(n8225) );
  AOI21_X1 U9720 ( .B1(n8226), .B2(n8225), .A(n8224), .ZN(n8231) );
  INV_X1 U9721 ( .A(n8227), .ZN(n8230) );
  OAI211_X1 U9722 ( .C1(n8231), .C2(n8230), .A(n8229), .B(n8228), .ZN(n8232)
         );
  NAND2_X1 U9723 ( .A1(n8232), .A2(n8605), .ZN(n8233) );
  AOI21_X1 U9724 ( .B1(n8234), .B2(n8233), .A(n8236), .ZN(n8235) );
  MUX2_X1 U9725 ( .A(n8236), .B(n8235), .S(n8274), .Z(n8238) );
  OAI22_X1 U9726 ( .A1(n8238), .A2(n8590), .B1(n8267), .B2(n8237), .ZN(n8242)
         );
  NAND2_X1 U9727 ( .A1(n8578), .A2(n8239), .ZN(n8241) );
  NAND2_X1 U9728 ( .A1(n8245), .A2(n8274), .ZN(n8240) );
  AOI22_X1 U9729 ( .A1(n8243), .A2(n8242), .B1(n8241), .B2(n8240), .ZN(n8253)
         );
  MUX2_X1 U9730 ( .A(n8245), .B(n8244), .S(n8274), .Z(n8246) );
  NAND2_X1 U9731 ( .A1(n8558), .A2(n8246), .ZN(n8252) );
  AND2_X1 U9732 ( .A1(n8254), .A2(n4331), .ZN(n8250) );
  AND2_X1 U9733 ( .A1(n8758), .A2(n8424), .ZN(n8248) );
  NOR2_X1 U9734 ( .A1(n8538), .A2(n8248), .ZN(n8249) );
  MUX2_X1 U9735 ( .A(n8250), .B(n8249), .S(n8274), .Z(n8251) );
  OAI21_X1 U9736 ( .B1(n8253), .B2(n8252), .A(n8251), .ZN(n8256) );
  MUX2_X1 U9737 ( .A(n8527), .B(n8254), .S(n8274), .Z(n8255) );
  NAND3_X1 U9738 ( .A1(n8256), .A2(n8106), .A3(n8255), .ZN(n8261) );
  AND2_X1 U9739 ( .A1(n8746), .A2(n8415), .ZN(n8258) );
  MUX2_X1 U9740 ( .A(n8258), .B(n8257), .S(n8267), .Z(n8259) );
  INV_X1 U9741 ( .A(n8259), .ZN(n8260) );
  NAND3_X1 U9742 ( .A1(n8262), .A2(n8261), .A3(n8260), .ZN(n8266) );
  NAND2_X1 U9743 ( .A1(n8423), .A2(n8274), .ZN(n8264) );
  NAND2_X1 U9744 ( .A1(n8531), .A2(n8267), .ZN(n8263) );
  MUX2_X1 U9745 ( .A(n8264), .B(n8263), .S(n8741), .Z(n8265) );
  NAND3_X1 U9746 ( .A1(n8312), .A2(n8266), .A3(n8265), .ZN(n8271) );
  MUX2_X1 U9747 ( .A(n8269), .B(n8268), .S(n8267), .Z(n8270) );
  NAND4_X1 U9748 ( .A1(n4661), .A2(n8272), .A3(n8271), .A4(n8270), .ZN(n8278)
         );
  INV_X1 U9749 ( .A(n8273), .ZN(n8275) );
  MUX2_X1 U9750 ( .A(n8276), .B(n8275), .S(n8274), .Z(n8277) );
  INV_X1 U9751 ( .A(n8317), .ZN(n8281) );
  NAND3_X1 U9752 ( .A1(n8281), .A2(n8282), .A3(n8280), .ZN(n8321) );
  NOR3_X1 U9753 ( .A1(n8284), .A2(n8283), .A3(n8282), .ZN(n8288) );
  INV_X1 U9754 ( .A(n6444), .ZN(n8285) );
  NAND4_X1 U9755 ( .A1(n8288), .A2(n8287), .A3(n8286), .A4(n8285), .ZN(n8292)
         );
  NOR4_X1 U9756 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), .ZN(n8296)
         );
  INV_X1 U9757 ( .A(n8293), .ZN(n8295) );
  NAND4_X1 U9758 ( .A1(n8296), .A2(n9567), .A3(n8295), .A4(n8294), .ZN(n8298)
         );
  NOR4_X1 U9759 ( .A1(n8300), .A2(n8299), .A3(n8298), .A4(n8297), .ZN(n8302)
         );
  AND4_X1 U9760 ( .A1(n8304), .A2(n8303), .A3(n8302), .A4(n8301), .ZN(n8305)
         );
  NAND4_X1 U9761 ( .A1(n8661), .A2(n8306), .A3(n8676), .A4(n8305), .ZN(n8307)
         );
  NOR4_X1 U9762 ( .A1(n8590), .A2(n8645), .A3(n8625), .A4(n8307), .ZN(n8308)
         );
  NAND4_X1 U9763 ( .A1(n8548), .A2(n8578), .A3(n8607), .A4(n8308), .ZN(n8309)
         );
  NOR4_X1 U9764 ( .A1(n8510), .A2(n8309), .A3(n8530), .A4(n8556), .ZN(n8310)
         );
  NAND4_X1 U9765 ( .A1(n8313), .A2(n8312), .A3(n8311), .A4(n8310), .ZN(n8314)
         );
  XNOR2_X1 U9766 ( .A(n8314), .B(n4864), .ZN(n8316) );
  OAI222_X1 U9767 ( .A1(n6366), .A2(n8319), .B1(n8318), .B2(n8317), .C1(n8316), 
        .C2(n8315), .ZN(n8320) );
  AOI22_X1 U9768 ( .A1(n8323), .A2(n8322), .B1(n8321), .B2(n8320), .ZN(n8329)
         );
  NAND3_X1 U9769 ( .A1(n8324), .A2(n8463), .A3(n8678), .ZN(n8325) );
  OAI211_X1 U9770 ( .C1(n8326), .C2(n8328), .A(n8325), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8327) );
  OAI21_X1 U9771 ( .B1(n8329), .B2(n8328), .A(n8327), .ZN(P2_U3244) );
  INV_X1 U9772 ( .A(n8330), .ZN(n8857) );
  OAI222_X1 U9773 ( .A1(n8334), .A2(n8857), .B1(n8333), .B2(n8332), .C1(n8331), 
        .C2(P1_U3084), .ZN(P1_U3324) );
  OAI222_X1 U9774 ( .A1(n8856), .A2(n8336), .B1(P2_U3152), .B2(n5492), .C1(
        n8858), .C2(n8335), .ZN(P2_U3330) );
  OAI211_X1 U9775 ( .C1(n8337), .C2(n8339), .A(n8338), .B(n8410), .ZN(n8343)
         );
  AOI22_X1 U9776 ( .A1(n8374), .A2(n8423), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8342) );
  AOI22_X1 U9777 ( .A1(n8524), .A2(n8398), .B1(n8375), .B2(n8486), .ZN(n8341)
         );
  NAND2_X1 U9778 ( .A1(n8746), .A2(n8406), .ZN(n8340) );
  NAND4_X1 U9779 ( .A1(n8343), .A2(n8342), .A3(n8341), .A4(n8340), .ZN(
        P2_U3216) );
  XNOR2_X1 U9780 ( .A(n8346), .B(n8345), .ZN(n8347) );
  XNOR2_X1 U9781 ( .A(n8344), .B(n8347), .ZN(n8352) );
  OAI22_X1 U9782 ( .A1(n8416), .A2(n8593), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8348), .ZN(n8350) );
  INV_X1 U9783 ( .A(n8398), .ZN(n8417) );
  OAI22_X1 U9784 ( .A1(n8417), .A2(n8597), .B1(n8592), .B2(n8414), .ZN(n8349)
         );
  AOI211_X1 U9785 ( .C1(n8767), .C2(n8406), .A(n8350), .B(n8349), .ZN(n8351)
         );
  OAI21_X1 U9786 ( .B1(n8352), .B2(n8408), .A(n8351), .ZN(P2_U3218) );
  INV_X1 U9787 ( .A(n8353), .ZN(n8355) );
  NAND2_X1 U9788 ( .A1(n8355), .A2(n8354), .ZN(n8356) );
  XNOR2_X1 U9789 ( .A(n8357), .B(n8356), .ZN(n8362) );
  AOI22_X1 U9790 ( .A1(n8374), .A2(n8663), .B1(n8358), .B2(n8656), .ZN(n8359)
         );
  NAND2_X1 U9791 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8458) );
  OAI211_X1 U9792 ( .C1(n8475), .C2(n8416), .A(n8359), .B(n8458), .ZN(n8360)
         );
  AOI21_X1 U9793 ( .B1(n8788), .B2(n8406), .A(n8360), .ZN(n8361) );
  OAI21_X1 U9794 ( .B1(n8362), .B2(n8408), .A(n8361), .ZN(P2_U3221) );
  OAI211_X1 U9795 ( .C1(n8365), .C2(n8364), .A(n8363), .B(n8410), .ZN(n8369)
         );
  AOI22_X1 U9796 ( .A1(n8374), .A2(n8629), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8368) );
  AOI22_X1 U9797 ( .A1(n8398), .A2(n8631), .B1(n8375), .B2(n8663), .ZN(n8367)
         );
  NAND2_X1 U9798 ( .A1(n8777), .A2(n8406), .ZN(n8366) );
  NAND4_X1 U9799 ( .A1(n8369), .A2(n8368), .A3(n8367), .A4(n8366), .ZN(
        P2_U3225) );
  OAI211_X1 U9800 ( .C1(n8370), .C2(n8373), .A(n8372), .B(n8410), .ZN(n8379)
         );
  AOI22_X1 U9801 ( .A1(n8374), .A2(n8486), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8378) );
  INV_X1 U9802 ( .A(n8592), .ZN(n8484) );
  AOI22_X1 U9803 ( .A1(n8565), .A2(n8398), .B1(n8375), .B2(n8484), .ZN(n8377)
         );
  NAND2_X1 U9804 ( .A1(n8758), .A2(n8406), .ZN(n8376) );
  NAND4_X1 U9805 ( .A1(n8379), .A2(n8378), .A3(n8377), .A4(n8376), .ZN(
        P2_U3227) );
  OAI211_X1 U9806 ( .C1(n8381), .C2(n8383), .A(n8382), .B(n8410), .ZN(n8389)
         );
  OAI22_X1 U9807 ( .A1(n8414), .A2(n8424), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8384), .ZN(n8387) );
  OAI22_X1 U9808 ( .A1(n8417), .A2(n8385), .B1(n8611), .B2(n8416), .ZN(n8386)
         );
  AOI211_X1 U9809 ( .C1(n8761), .C2(n8406), .A(n8387), .B(n8386), .ZN(n8388)
         );
  NAND2_X1 U9810 ( .A1(n8389), .A2(n8388), .ZN(P2_U3231) );
  INV_X1 U9811 ( .A(n8783), .ZN(n8641) );
  OAI211_X1 U9812 ( .C1(n8392), .C2(n8391), .A(n8390), .B(n8410), .ZN(n8400)
         );
  INV_X1 U9813 ( .A(n8393), .ZN(n8639) );
  OAI22_X1 U9814 ( .A1(n8610), .A2(n8693), .B1(n8477), .B2(n8695), .ZN(n8646)
         );
  INV_X1 U9815 ( .A(n8646), .ZN(n8395) );
  OAI22_X1 U9816 ( .A1(n8396), .A2(n8395), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8394), .ZN(n8397) );
  AOI21_X1 U9817 ( .B1(n8398), .B2(n8639), .A(n8397), .ZN(n8399) );
  OAI211_X1 U9818 ( .C1(n8641), .C2(n8422), .A(n8400), .B(n8399), .ZN(P2_U3235) );
  XOR2_X1 U9819 ( .A(n8402), .B(n8401), .Z(n8409) );
  OAI22_X1 U9820 ( .A1(n8414), .A2(n8611), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8403), .ZN(n8405) );
  OAI22_X1 U9821 ( .A1(n8417), .A2(n8613), .B1(n8610), .B2(n8416), .ZN(n8404)
         );
  AOI211_X1 U9822 ( .C1(n8774), .C2(n8406), .A(n8405), .B(n8404), .ZN(n8407)
         );
  OAI21_X1 U9823 ( .B1(n8409), .B2(n8408), .A(n8407), .ZN(P2_U3237) );
  INV_X1 U9824 ( .A(n8752), .ZN(n8545) );
  OAI211_X1 U9825 ( .C1(n8413), .C2(n8412), .A(n8411), .B(n8410), .ZN(n8421)
         );
  NOR2_X1 U9826 ( .A1(n8415), .A2(n8414), .ZN(n8419) );
  OAI22_X1 U9827 ( .A1(n8417), .A2(n8542), .B1(n8424), .B2(n8416), .ZN(n8418)
         );
  AOI211_X1 U9828 ( .C1(P2_REG3_REG_26__SCAN_IN), .C2(P2_U3152), .A(n8419), 
        .B(n8418), .ZN(n8420) );
  OAI211_X1 U9829 ( .C1(n8545), .C2(n8422), .A(n8421), .B(n8420), .ZN(P2_U3242) );
  MUX2_X1 U9830 ( .A(n8423), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8425), .Z(
        P2_U3580) );
  MUX2_X1 U9831 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8549), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9832 ( .A(n8486), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8425), .Z(
        P2_U3578) );
  INV_X1 U9833 ( .A(n8424), .ZN(n8581) );
  MUX2_X1 U9834 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8581), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9835 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8484), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U9836 ( .A(n8580), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8425), .Z(
        P2_U3575) );
  MUX2_X1 U9837 ( .A(n8629), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8425), .Z(
        P2_U3574) );
  INV_X1 U9838 ( .A(n8610), .ZN(n8481) );
  MUX2_X1 U9839 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8481), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9840 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8663), .S(P2_U3966), .Z(
        P2_U3572) );
  INV_X1 U9841 ( .A(n8477), .ZN(n8681) );
  MUX2_X1 U9842 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8681), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9843 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8662), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9844 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8679), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9845 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8426), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9846 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8427), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9847 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8428), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9848 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8429), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9849 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8430), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9850 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8431), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9851 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8432), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9852 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8433), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9853 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8434), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9854 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8435), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9855 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8436), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9856 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8437), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9857 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8438), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9858 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8439), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9859 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8440), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9860 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6441), .S(P2_U3966), .Z(
        P2_U3553) );
  MUX2_X1 U9861 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n6379), .S(P2_U3966), .Z(
        P2_U3552) );
  NOR2_X1 U9862 ( .A1(n8446), .A2(n8441), .ZN(n8442) );
  NOR2_X1 U9863 ( .A1(n8443), .A2(n8442), .ZN(n8444) );
  XOR2_X1 U9864 ( .A(n8444), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8455) );
  INV_X1 U9865 ( .A(n8452), .ZN(n8447) );
  NAND2_X1 U9866 ( .A1(n8447), .A2(n8453), .ZN(n8449) );
  OAI211_X1 U9867 ( .C1(n8455), .C2(n8450), .A(n8449), .B(n8448), .ZN(n8451)
         );
  INV_X1 U9868 ( .A(n8451), .ZN(n8457) );
  AOI22_X1 U9869 ( .A1(n8455), .A2(n8454), .B1(n8453), .B2(n8452), .ZN(n8456)
         );
  MUX2_X1 U9870 ( .A(n8457), .B(n8456), .S(n4864), .Z(n8459) );
  OAI211_X1 U9871 ( .C1(n8461), .C2(n8460), .A(n8459), .B(n8458), .ZN(P2_U3264) );
  INV_X1 U9872 ( .A(n8746), .ZN(n8526) );
  INV_X1 U9873 ( .A(n8758), .ZN(n8462) );
  NOR2_X2 U9874 ( .A1(n8671), .A2(n8792), .ZN(n8670) );
  NAND2_X1 U9875 ( .A1(n8601), .A2(n8612), .ZN(n8594) );
  NOR2_X2 U9876 ( .A1(n8594), .A2(n8761), .ZN(n8573) );
  NOR2_X2 U9877 ( .A1(n8562), .A2(n8752), .ZN(n8541) );
  INV_X1 U9878 ( .A(n8499), .ZN(n8734) );
  XOR2_X1 U9879 ( .A(n8727), .B(n8468), .Z(n8729) );
  NAND2_X1 U9880 ( .A1(n8463), .A2(P2_B_REG_SCAN_IN), .ZN(n8464) );
  NAND2_X1 U9881 ( .A1(n8680), .A2(n8464), .ZN(n8495) );
  NOR2_X1 U9882 ( .A1(n8465), .A2(n8495), .ZN(n8726) );
  INV_X1 U9883 ( .A(n8726), .ZN(n8731) );
  NOR2_X1 U9884 ( .A1(n9588), .A2(n8731), .ZN(n8471) );
  AOI21_X1 U9885 ( .B1(n9588), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8471), .ZN(
        n8467) );
  NAND2_X1 U9886 ( .A1(n8727), .A2(n9577), .ZN(n8466) );
  OAI211_X1 U9887 ( .C1(n8729), .C2(n8707), .A(n8467), .B(n8466), .ZN(P2_U3265) );
  AOI21_X1 U9888 ( .B1(n8470), .B2(n8469), .A(n8468), .ZN(n8730) );
  NAND2_X1 U9889 ( .A1(n8730), .A2(n8719), .ZN(n8473) );
  AOI21_X1 U9890 ( .B1(n9588), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8471), .ZN(
        n8472) );
  OAI211_X1 U9891 ( .C1(n4472), .C2(n8674), .A(n8473), .B(n8472), .ZN(P2_U3266) );
  OAI21_X1 U9892 ( .B1(n8679), .B2(n8799), .A(n8474), .ZN(n8669) );
  NOR2_X1 U9893 ( .A1(n8792), .A2(n8662), .ZN(n8476) );
  INV_X1 U9894 ( .A(n8792), .ZN(n8675) );
  INV_X1 U9895 ( .A(n8652), .ZN(n8479) );
  AOI21_X2 U9896 ( .B1(n8479), .B2(n4788), .A(n8478), .ZN(n8637) );
  NAND2_X1 U9897 ( .A1(n8623), .A2(n8610), .ZN(n8482) );
  XNOR2_X1 U9898 ( .A(n8489), .B(n8490), .ZN(n8733) );
  INV_X1 U9899 ( .A(n8733), .ZN(n8505) );
  XNOR2_X1 U9900 ( .A(n8491), .B(n8490), .ZN(n8493) );
  NAND2_X1 U9901 ( .A1(n8493), .A2(n8492), .ZN(n8498) );
  NAND2_X1 U9902 ( .A1(n8498), .A2(n8497), .ZN(n8737) );
  XOR2_X1 U9903 ( .A(n8499), .B(n8512), .Z(n8735) );
  NOR2_X1 U9904 ( .A1(n8735), .A2(n8707), .ZN(n8503) );
  AOI22_X1 U9905 ( .A1(n9588), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8500), .B2(
        n9576), .ZN(n8501) );
  OAI21_X1 U9906 ( .B1(n8734), .B2(n8674), .A(n8501), .ZN(n8502) );
  AOI211_X1 U9907 ( .C1(n8737), .C2(n8699), .A(n8503), .B(n8502), .ZN(n8504)
         );
  OAI21_X1 U9908 ( .B1(n8505), .B2(n8686), .A(n8504), .ZN(P2_U3267) );
  XOR2_X1 U9909 ( .A(n8510), .B(n8506), .Z(n8508) );
  AOI222_X1 U9910 ( .A1(n8492), .A2(n8508), .B1(n8549), .B2(n8678), .C1(n8507), 
        .C2(n8680), .ZN(n8744) );
  OAI21_X1 U9911 ( .B1(n8511), .B2(n8510), .A(n8509), .ZN(n8740) );
  NAND2_X1 U9912 ( .A1(n8740), .A2(n8711), .ZN(n8517) );
  AOI21_X1 U9913 ( .B1(n8741), .B2(n8521), .A(n8512), .ZN(n8742) );
  AOI22_X1 U9914 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(n9588), .B1(n8513), .B2(
        n9576), .ZN(n8514) );
  OAI21_X1 U9915 ( .B1(n4663), .B2(n8674), .A(n8514), .ZN(n8515) );
  AOI21_X1 U9916 ( .B1(n8742), .B2(n8719), .A(n8515), .ZN(n8516) );
  OAI211_X1 U9917 ( .C1(n9588), .C2(n8744), .A(n8517), .B(n8516), .ZN(P2_U3268) );
  OAI21_X1 U9918 ( .B1(n8519), .B2(n8530), .A(n8518), .ZN(n8520) );
  INV_X1 U9919 ( .A(n8520), .ZN(n8750) );
  INV_X1 U9920 ( .A(n8541), .ZN(n8523) );
  INV_X1 U9921 ( .A(n8521), .ZN(n8522) );
  AOI21_X1 U9922 ( .B1(n8746), .B2(n8523), .A(n8522), .ZN(n8747) );
  AOI22_X1 U9923 ( .A1(n9588), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8524), .B2(
        n9576), .ZN(n8525) );
  OAI21_X1 U9924 ( .B1(n8526), .B2(n8674), .A(n8525), .ZN(n8535) );
  NAND2_X1 U9925 ( .A1(n8546), .A2(n8527), .ZN(n8529) );
  AOI211_X1 U9926 ( .C1(n8530), .C2(n8529), .A(n8643), .B(n8528), .ZN(n8533)
         );
  OAI22_X1 U9927 ( .A1(n8531), .A2(n8693), .B1(n8561), .B2(n8695), .ZN(n8532)
         );
  NOR2_X1 U9928 ( .A1(n8533), .A2(n8532), .ZN(n8749) );
  NOR2_X1 U9929 ( .A1(n8749), .A2(n9588), .ZN(n8534) );
  AOI211_X1 U9930 ( .C1(n8747), .C2(n8719), .A(n8535), .B(n8534), .ZN(n8536)
         );
  OAI21_X1 U9931 ( .B1(n8750), .B2(n8686), .A(n8536), .ZN(P2_U3269) );
  OAI21_X1 U9932 ( .B1(n8539), .B2(n8538), .A(n8537), .ZN(n8540) );
  INV_X1 U9933 ( .A(n8540), .ZN(n8755) );
  AOI211_X1 U9934 ( .C1(n8752), .C2(n8562), .A(n9692), .B(n8541), .ZN(n8751)
         );
  INV_X1 U9935 ( .A(n8542), .ZN(n8543) );
  AOI22_X1 U9936 ( .A1(n9588), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8543), .B2(
        n9576), .ZN(n8544) );
  OAI21_X1 U9937 ( .B1(n8545), .B2(n8674), .A(n8544), .ZN(n8552) );
  OAI21_X1 U9938 ( .B1(n8548), .B2(n8547), .A(n8546), .ZN(n8550) );
  AOI222_X1 U9939 ( .A1(n8492), .A2(n8550), .B1(n8549), .B2(n8680), .C1(n8581), 
        .C2(n8678), .ZN(n8754) );
  NOR2_X1 U9940 ( .A1(n8754), .A2(n9588), .ZN(n8551) );
  AOI211_X1 U9941 ( .C1(n8751), .C2(n8667), .A(n8552), .B(n8551), .ZN(n8553)
         );
  OAI21_X1 U9942 ( .B1(n8755), .B2(n8686), .A(n8553), .ZN(P2_U3270) );
  OAI21_X1 U9943 ( .B1(n8554), .B2(n8556), .A(n8555), .ZN(n8557) );
  INV_X1 U9944 ( .A(n8557), .ZN(n8760) );
  AOI22_X1 U9945 ( .A1(n8758), .A2(n9577), .B1(n9588), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8571) );
  XNOR2_X1 U9946 ( .A(n8559), .B(n8558), .ZN(n8560) );
  OAI222_X1 U9947 ( .A1(n8693), .A2(n8561), .B1(n8695), .B2(n8592), .C1(n8560), 
        .C2(n8643), .ZN(n8756) );
  INV_X1 U9948 ( .A(n8573), .ZN(n8564) );
  INV_X1 U9949 ( .A(n8562), .ZN(n8563) );
  AOI211_X1 U9950 ( .C1(n8758), .C2(n8564), .A(n9692), .B(n8563), .ZN(n8757)
         );
  INV_X1 U9951 ( .A(n8757), .ZN(n8568) );
  INV_X1 U9952 ( .A(n8565), .ZN(n8566) );
  OAI22_X1 U9953 ( .A1(n8568), .A2(n8567), .B1(n8705), .B2(n8566), .ZN(n8569)
         );
  OAI21_X1 U9954 ( .B1(n8756), .B2(n8569), .A(n8699), .ZN(n8570) );
  OAI211_X1 U9955 ( .C1(n8760), .C2(n8686), .A(n8571), .B(n8570), .ZN(P2_U3271) );
  XOR2_X1 U9956 ( .A(n8578), .B(n8572), .Z(n8765) );
  AOI21_X1 U9957 ( .B1(n8761), .B2(n8594), .A(n8573), .ZN(n8762) );
  INV_X1 U9958 ( .A(n8761), .ZN(n8576) );
  AOI22_X1 U9959 ( .A1(n9588), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8574), .B2(
        n9576), .ZN(n8575) );
  OAI21_X1 U9960 ( .B1(n8576), .B2(n8674), .A(n8575), .ZN(n8585) );
  OAI211_X1 U9961 ( .C1(n8579), .C2(n8578), .A(n8577), .B(n8492), .ZN(n8583)
         );
  AOI22_X1 U9962 ( .A1(n8581), .A2(n8680), .B1(n8678), .B2(n8580), .ZN(n8582)
         );
  AND2_X1 U9963 ( .A1(n8583), .A2(n8582), .ZN(n8764) );
  NOR2_X1 U9964 ( .A1(n8764), .A2(n9588), .ZN(n8584) );
  AOI211_X1 U9965 ( .C1(n8762), .C2(n8719), .A(n8585), .B(n8584), .ZN(n8586)
         );
  OAI21_X1 U9966 ( .B1(n8765), .B2(n8686), .A(n8586), .ZN(P2_U3272) );
  OAI21_X1 U9967 ( .B1(n8588), .B2(n8590), .A(n8587), .ZN(n8771) );
  AOI21_X1 U9968 ( .B1(n8590), .B2(n8589), .A(n4290), .ZN(n8591) );
  OAI222_X1 U9969 ( .A1(n8695), .A2(n8593), .B1(n8693), .B2(n8592), .C1(n8643), 
        .C2(n8591), .ZN(n8766) );
  INV_X1 U9970 ( .A(n8612), .ZN(n8596) );
  INV_X1 U9971 ( .A(n8594), .ZN(n8595) );
  AOI21_X1 U9972 ( .B1(n8767), .B2(n8596), .A(n8595), .ZN(n8768) );
  NAND2_X1 U9973 ( .A1(n8768), .A2(n8719), .ZN(n8600) );
  INV_X1 U9974 ( .A(n8597), .ZN(n8598) );
  AOI22_X1 U9975 ( .A1(n9588), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8598), .B2(
        n9576), .ZN(n8599) );
  OAI211_X1 U9976 ( .C1(n8601), .C2(n8674), .A(n8600), .B(n8599), .ZN(n8602)
         );
  AOI21_X1 U9977 ( .B1(n8766), .B2(n8699), .A(n8602), .ZN(n8603) );
  OAI21_X1 U9978 ( .B1(n8771), .B2(n8686), .A(n8603), .ZN(P2_U3273) );
  XNOR2_X1 U9979 ( .A(n8604), .B(n8607), .ZN(n8776) );
  INV_X1 U9980 ( .A(n8605), .ZN(n8606) );
  NOR2_X1 U9981 ( .A1(n8624), .A2(n8606), .ZN(n8608) );
  XNOR2_X1 U9982 ( .A(n8608), .B(n8607), .ZN(n8609) );
  OAI222_X1 U9983 ( .A1(n8693), .A2(n8611), .B1(n8695), .B2(n8610), .C1(n8609), 
        .C2(n8643), .ZN(n8772) );
  AOI211_X1 U9984 ( .C1(n8774), .C2(n8620), .A(n9692), .B(n8612), .ZN(n8773)
         );
  INV_X1 U9985 ( .A(n9583), .ZN(n8650) );
  NAND2_X1 U9986 ( .A1(n8773), .A2(n8650), .ZN(n8616) );
  INV_X1 U9987 ( .A(n8613), .ZN(n8614) );
  AOI22_X1 U9988 ( .A1(n9588), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8614), .B2(
        n9576), .ZN(n8615) );
  OAI211_X1 U9989 ( .C1(n4466), .C2(n8674), .A(n8616), .B(n8615), .ZN(n8617)
         );
  AOI21_X1 U9990 ( .B1(n8772), .B2(n8699), .A(n8617), .ZN(n8618) );
  OAI21_X1 U9991 ( .B1(n8776), .B2(n8686), .A(n8618), .ZN(P2_U3274) );
  XNOR2_X1 U9992 ( .A(n8619), .B(n8625), .ZN(n8781) );
  INV_X1 U9993 ( .A(n8620), .ZN(n8621) );
  AOI21_X1 U9994 ( .B1(n8777), .B2(n4470), .A(n8621), .ZN(n8778) );
  INV_X1 U9995 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8622) );
  OAI22_X1 U9996 ( .A1(n8623), .A2(n8674), .B1(n8622), .B2(n8699), .ZN(n8634)
         );
  INV_X1 U9997 ( .A(n8624), .ZN(n8628) );
  OAI21_X1 U9998 ( .B1(n8642), .B2(n8626), .A(n8625), .ZN(n8627) );
  NAND2_X1 U9999 ( .A1(n8628), .A2(n8627), .ZN(n8630) );
  AOI222_X1 U10000 ( .A1(n8492), .A2(n8630), .B1(n8629), .B2(n8680), .C1(n8663), .C2(n8678), .ZN(n8780) );
  NAND2_X1 U10001 ( .A1(n9576), .A2(n8631), .ZN(n8632) );
  AOI21_X1 U10002 ( .B1(n8780), .B2(n8632), .A(n9588), .ZN(n8633) );
  AOI211_X1 U10003 ( .C1(n8778), .C2(n8719), .A(n8634), .B(n8633), .ZN(n8635)
         );
  OAI21_X1 U10004 ( .B1(n8686), .B2(n8781), .A(n8635), .ZN(P2_U3275) );
  OAI21_X1 U10005 ( .B1(n8637), .B2(n8645), .A(n8636), .ZN(n8786) );
  AOI211_X1 U10006 ( .C1(n8783), .C2(n8653), .A(n9692), .B(n8638), .ZN(n8782)
         );
  AOI22_X1 U10007 ( .A1(n9588), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8639), .B2(
        n9576), .ZN(n8640) );
  OAI21_X1 U10008 ( .B1(n8641), .B2(n8674), .A(n8640), .ZN(n8649) );
  AOI211_X1 U10009 ( .C1(n8645), .C2(n8644), .A(n8643), .B(n8642), .ZN(n8647)
         );
  NOR2_X1 U10010 ( .A1(n8647), .A2(n8646), .ZN(n8785) );
  NOR2_X1 U10011 ( .A1(n8785), .A2(n9588), .ZN(n8648) );
  AOI211_X1 U10012 ( .C1(n8782), .C2(n8650), .A(n8649), .B(n8648), .ZN(n8651)
         );
  OAI21_X1 U10013 ( .B1(n8686), .B2(n8786), .A(n8651), .ZN(P2_U3276) );
  XOR2_X1 U10014 ( .A(n8661), .B(n8652), .Z(n8791) );
  INV_X1 U10015 ( .A(n8670), .ZN(n8655) );
  INV_X1 U10016 ( .A(n8653), .ZN(n8654) );
  AOI211_X1 U10017 ( .C1(n8788), .C2(n8655), .A(n9692), .B(n8654), .ZN(n8787)
         );
  AOI22_X1 U10018 ( .A1(n9588), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8656), .B2(
        n9576), .ZN(n8657) );
  OAI21_X1 U10019 ( .B1(n8658), .B2(n8674), .A(n8657), .ZN(n8666) );
  OAI21_X1 U10020 ( .B1(n8661), .B2(n8660), .A(n8659), .ZN(n8664) );
  AOI222_X1 U10021 ( .A1(n8492), .A2(n8664), .B1(n8663), .B2(n8680), .C1(n8662), .C2(n8678), .ZN(n8790) );
  NOR2_X1 U10022 ( .A1(n8790), .A2(n9588), .ZN(n8665) );
  AOI211_X1 U10023 ( .C1(n8787), .C2(n8667), .A(n8666), .B(n8665), .ZN(n8668)
         );
  OAI21_X1 U10024 ( .B1(n8791), .B2(n8686), .A(n8668), .ZN(P2_U3277) );
  XNOR2_X1 U10025 ( .A(n8669), .B(n8676), .ZN(n8796) );
  AOI21_X1 U10026 ( .B1(n8792), .B2(n8671), .A(n8670), .ZN(n8793) );
  AOI22_X1 U10027 ( .A1(n9588), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8672), .B2(
        n9576), .ZN(n8673) );
  OAI21_X1 U10028 ( .B1(n8675), .B2(n8674), .A(n8673), .ZN(n8684) );
  OAI21_X1 U10029 ( .B1(n8677), .B2(n8676), .A(n4313), .ZN(n8682) );
  AOI222_X1 U10030 ( .A1(n8492), .A2(n8682), .B1(n8681), .B2(n8680), .C1(n8679), .C2(n8678), .ZN(n8795) );
  NOR2_X1 U10031 ( .A1(n8795), .A2(n9588), .ZN(n8683) );
  AOI211_X1 U10032 ( .C1(n8793), .C2(n8719), .A(n8684), .B(n8683), .ZN(n8685)
         );
  OAI21_X1 U10033 ( .B1(n8796), .B2(n8686), .A(n8685), .ZN(P2_U3278) );
  NAND2_X1 U10034 ( .A1(n8688), .A2(n8687), .ZN(n8690) );
  NAND2_X1 U10035 ( .A1(n8690), .A2(n8689), .ZN(n8692) );
  OAI21_X1 U10036 ( .B1(n8709), .B2(n8692), .A(n8691), .ZN(n8698) );
  OAI22_X1 U10037 ( .A1(n8696), .A2(n8695), .B1(n8694), .B2(n8693), .ZN(n8697)
         );
  AOI21_X1 U10038 ( .B1(n8698), .B2(n8492), .A(n8697), .ZN(n9653) );
  MUX2_X1 U10039 ( .A(n9817), .B(n9653), .S(n8699), .Z(n8714) );
  OR2_X1 U10040 ( .A1(n8701), .A2(n8700), .ZN(n8702) );
  NAND2_X1 U10041 ( .A1(n8703), .A2(n8702), .ZN(n9648) );
  INV_X1 U10042 ( .A(n8704), .ZN(n8706) );
  OAI22_X1 U10043 ( .A1(n8707), .A2(n9648), .B1(n8706), .B2(n8705), .ZN(n8708)
         );
  AOI21_X1 U10044 ( .B1(n9577), .B2(n9649), .A(n8708), .ZN(n8713) );
  NAND2_X1 U10045 ( .A1(n8710), .A2(n8709), .ZN(n9646) );
  NAND3_X1 U10046 ( .A1(n9647), .A2(n9646), .A3(n8711), .ZN(n8712) );
  NAND3_X1 U10047 ( .A1(n8714), .A2(n8713), .A3(n8712), .ZN(P2_U3290) );
  MUX2_X1 U10048 ( .A(n8715), .B(P2_REG2_REG_3__SCAN_IN), .S(n9588), .Z(n8716)
         );
  INV_X1 U10049 ( .A(n8716), .ZN(n8725) );
  AOI22_X1 U10050 ( .A1(n8719), .A2(n8718), .B1(n9576), .B2(n8717), .ZN(n8724)
         );
  AOI22_X1 U10051 ( .A1(n8722), .A2(n8721), .B1(n9577), .B2(n8720), .ZN(n8723)
         );
  NAND3_X1 U10052 ( .A1(n8725), .A2(n8724), .A3(n8723), .ZN(P2_U3293) );
  AOI21_X1 U10053 ( .B1(n8727), .B2(n9677), .A(n8726), .ZN(n8728) );
  OAI21_X1 U10054 ( .B1(n8729), .B2(n9692), .A(n8728), .ZN(n8825) );
  MUX2_X1 U10055 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8825), .S(n9715), .Z(
        P2_U3551) );
  NAND2_X1 U10056 ( .A1(n8730), .A2(n9650), .ZN(n8732) );
  OAI211_X1 U10057 ( .C1(n4472), .C2(n9690), .A(n8732), .B(n8731), .ZN(n8826)
         );
  MUX2_X1 U10058 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8826), .S(n9715), .Z(
        P2_U3550) );
  NAND2_X1 U10059 ( .A1(n8733), .A2(n9697), .ZN(n8739) );
  OAI22_X1 U10060 ( .A1(n8735), .A2(n9692), .B1(n8734), .B2(n9690), .ZN(n8736)
         );
  NOR2_X1 U10061 ( .A1(n8737), .A2(n8736), .ZN(n8738) );
  NAND2_X1 U10062 ( .A1(n8739), .A2(n8738), .ZN(n8827) );
  MUX2_X1 U10063 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8827), .S(n9715), .Z(
        P2_U3549) );
  INV_X1 U10064 ( .A(n8740), .ZN(n8745) );
  AOI22_X1 U10065 ( .A1(n8742), .A2(n9650), .B1(n9677), .B2(n8741), .ZN(n8743)
         );
  OAI211_X1 U10066 ( .C1(n8745), .C2(n8816), .A(n8744), .B(n8743), .ZN(n8828)
         );
  MUX2_X1 U10067 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8828), .S(n9715), .Z(
        P2_U3548) );
  AOI22_X1 U10068 ( .A1(n8747), .A2(n9650), .B1(n9677), .B2(n8746), .ZN(n8748)
         );
  OAI211_X1 U10069 ( .C1(n8750), .C2(n8816), .A(n8749), .B(n8748), .ZN(n8829)
         );
  MUX2_X1 U10070 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8829), .S(n9715), .Z(
        P2_U3547) );
  AOI21_X1 U10071 ( .B1(n9677), .B2(n8752), .A(n8751), .ZN(n8753) );
  OAI211_X1 U10072 ( .C1(n8755), .C2(n8816), .A(n8754), .B(n8753), .ZN(n8830)
         );
  MUX2_X1 U10073 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8830), .S(n9715), .Z(
        P2_U3546) );
  AOI211_X1 U10074 ( .C1(n9677), .C2(n8758), .A(n8757), .B(n8756), .ZN(n8759)
         );
  OAI21_X1 U10075 ( .B1(n8760), .B2(n8816), .A(n8759), .ZN(n8831) );
  MUX2_X1 U10076 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8831), .S(n9715), .Z(
        P2_U3545) );
  AOI22_X1 U10077 ( .A1(n8762), .A2(n9650), .B1(n9677), .B2(n8761), .ZN(n8763)
         );
  OAI211_X1 U10078 ( .C1(n8765), .C2(n8816), .A(n8764), .B(n8763), .ZN(n8832)
         );
  MUX2_X1 U10079 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8832), .S(n9715), .Z(
        P2_U3544) );
  INV_X1 U10080 ( .A(n8766), .ZN(n8770) );
  AOI22_X1 U10081 ( .A1(n8768), .A2(n9650), .B1(n9677), .B2(n8767), .ZN(n8769)
         );
  OAI211_X1 U10082 ( .C1(n8771), .C2(n8816), .A(n8770), .B(n8769), .ZN(n8833)
         );
  MUX2_X1 U10083 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8833), .S(n9715), .Z(
        P2_U3543) );
  AOI211_X1 U10084 ( .C1(n9677), .C2(n8774), .A(n8773), .B(n8772), .ZN(n8775)
         );
  OAI21_X1 U10085 ( .B1(n8776), .B2(n8816), .A(n8775), .ZN(n8834) );
  MUX2_X1 U10086 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8834), .S(n9715), .Z(
        P2_U3542) );
  AOI22_X1 U10087 ( .A1(n8778), .A2(n9650), .B1(n9677), .B2(n8777), .ZN(n8779)
         );
  OAI211_X1 U10088 ( .C1(n8781), .C2(n8816), .A(n8780), .B(n8779), .ZN(n8835)
         );
  MUX2_X1 U10089 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8835), .S(n9715), .Z(
        P2_U3541) );
  AOI21_X1 U10090 ( .B1(n9677), .B2(n8783), .A(n8782), .ZN(n8784) );
  OAI211_X1 U10091 ( .C1(n8786), .C2(n8816), .A(n8785), .B(n8784), .ZN(n8836)
         );
  MUX2_X1 U10092 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8836), .S(n9715), .Z(
        P2_U3540) );
  AOI21_X1 U10093 ( .B1(n9677), .B2(n8788), .A(n8787), .ZN(n8789) );
  OAI211_X1 U10094 ( .C1(n8791), .C2(n8816), .A(n8790), .B(n8789), .ZN(n8837)
         );
  MUX2_X1 U10095 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8837), .S(n9715), .Z(
        P2_U3539) );
  AOI22_X1 U10096 ( .A1(n8793), .A2(n9650), .B1(n9677), .B2(n8792), .ZN(n8794)
         );
  OAI211_X1 U10097 ( .C1(n8796), .C2(n8816), .A(n8795), .B(n8794), .ZN(n8838)
         );
  MUX2_X1 U10098 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8838), .S(n9715), .Z(
        P2_U3538) );
  AOI211_X1 U10099 ( .C1(n9677), .C2(n8799), .A(n8798), .B(n8797), .ZN(n8800)
         );
  OAI21_X1 U10100 ( .B1(n8801), .B2(n8816), .A(n8800), .ZN(n8839) );
  MUX2_X1 U10101 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8839), .S(n9715), .Z(
        P2_U3537) );
  AOI22_X1 U10102 ( .A1(n8803), .A2(n9650), .B1(n9677), .B2(n8802), .ZN(n8804)
         );
  OAI211_X1 U10103 ( .C1(n8806), .C2(n9681), .A(n8805), .B(n8804), .ZN(n8840)
         );
  MUX2_X1 U10104 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8840), .S(n9715), .Z(
        P2_U3536) );
  AOI22_X1 U10105 ( .A1(n8808), .A2(n9650), .B1(n9677), .B2(n8807), .ZN(n8809)
         );
  OAI211_X1 U10106 ( .C1(n8811), .C2(n8816), .A(n8810), .B(n8809), .ZN(n8841)
         );
  MUX2_X1 U10107 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8841), .S(n9715), .Z(
        P2_U3535) );
  AOI22_X1 U10108 ( .A1(n8813), .A2(n9650), .B1(n9677), .B2(n8812), .ZN(n8814)
         );
  OAI211_X1 U10109 ( .C1(n8817), .C2(n8816), .A(n8815), .B(n8814), .ZN(n8842)
         );
  MUX2_X1 U10110 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8842), .S(n9715), .Z(
        P2_U3534) );
  NAND3_X1 U10111 ( .A1(n8819), .A2(n9697), .A3(n8818), .ZN(n8824) );
  AOI22_X1 U10112 ( .A1(n8821), .A2(n9650), .B1(n9677), .B2(n8820), .ZN(n8822)
         );
  NAND3_X1 U10113 ( .A1(n8824), .A2(n8823), .A3(n8822), .ZN(n8843) );
  MUX2_X1 U10114 ( .A(n8843), .B(P2_REG1_REG_13__SCAN_IN), .S(n9713), .Z(
        P2_U3533) );
  MUX2_X1 U10115 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8825), .S(n9700), .Z(
        P2_U3519) );
  MUX2_X1 U10116 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8826), .S(n9700), .Z(
        P2_U3518) );
  MUX2_X1 U10117 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8827), .S(n9700), .Z(
        P2_U3517) );
  MUX2_X1 U10118 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8828), .S(n9700), .Z(
        P2_U3516) );
  MUX2_X1 U10119 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8829), .S(n9700), .Z(
        P2_U3515) );
  MUX2_X1 U10120 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8830), .S(n9700), .Z(
        P2_U3514) );
  MUX2_X1 U10121 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8831), .S(n9700), .Z(
        P2_U3513) );
  MUX2_X1 U10122 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8832), .S(n9700), .Z(
        P2_U3512) );
  MUX2_X1 U10123 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8833), .S(n9700), .Z(
        P2_U3511) );
  MUX2_X1 U10124 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8834), .S(n9700), .Z(
        P2_U3510) );
  MUX2_X1 U10125 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8835), .S(n9700), .Z(
        P2_U3509) );
  MUX2_X1 U10126 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8836), .S(n9700), .Z(
        P2_U3508) );
  MUX2_X1 U10127 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8837), .S(n9700), .Z(
        P2_U3507) );
  MUX2_X1 U10128 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8838), .S(n9700), .Z(
        P2_U3505) );
  MUX2_X1 U10129 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8839), .S(n9700), .Z(
        P2_U3502) );
  MUX2_X1 U10130 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8840), .S(n9700), .Z(
        P2_U3499) );
  MUX2_X1 U10131 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8841), .S(n9700), .Z(
        P2_U3496) );
  MUX2_X1 U10132 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8842), .S(n9700), .Z(
        P2_U3493) );
  MUX2_X1 U10133 ( .A(n8843), .B(P2_REG0_REG_13__SCAN_IN), .S(n9698), .Z(
        P2_U3490) );
  INV_X1 U10134 ( .A(n8844), .ZN(n9365) );
  NOR4_X1 U10135 ( .A1(n8846), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8845), .A4(
        P2_U3152), .ZN(n8847) );
  AOI21_X1 U10136 ( .B1(n8851), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8847), .ZN(
        n8848) );
  OAI21_X1 U10137 ( .B1(n9365), .B2(n8858), .A(n8848), .ZN(P2_U3327) );
  INV_X1 U10138 ( .A(n8849), .ZN(n9369) );
  AOI22_X1 U10139 ( .A1(n8850), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8851), .ZN(n8852) );
  OAI21_X1 U10140 ( .B1(n9369), .B2(n8858), .A(n8852), .ZN(P2_U3328) );
  OAI222_X1 U10141 ( .A1(n8858), .A2(n8857), .B1(n8856), .B2(n8855), .C1(n8854), .C2(P2_U3152), .ZN(P2_U3329) );
  MUX2_X1 U10142 ( .A(n8860), .B(n8859), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10143 ( .A(n8861), .ZN(n8863) );
  NOR2_X1 U10144 ( .A1(n8863), .A2(n8862), .ZN(n8864) );
  XNOR2_X1 U10145 ( .A(n8865), .B(n8864), .ZN(n8870) );
  NAND2_X1 U10146 ( .A1(n8957), .A2(n9114), .ZN(n8867) );
  AOI22_X1 U10147 ( .A1(n4703), .A2(n8928), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8866) );
  OAI211_X1 U10148 ( .C1(n9121), .C2(n8952), .A(n8867), .B(n8866), .ZN(n8868)
         );
  AOI21_X1 U10149 ( .B1(n9269), .B2(n8914), .A(n8868), .ZN(n8869) );
  OAI21_X1 U10150 ( .B1(n8870), .B2(n8947), .A(n8869), .ZN(P1_U3212) );
  NAND2_X1 U10151 ( .A1(n8872), .A2(n8871), .ZN(n8874) );
  XNOR2_X1 U10152 ( .A(n8874), .B(n8873), .ZN(n8879) );
  NAND2_X1 U10153 ( .A1(n8957), .A2(n9179), .ZN(n8876) );
  AOI22_X1 U10154 ( .A1(n4688), .A2(n8928), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8875) );
  OAI211_X1 U10155 ( .C1(n9205), .C2(n8952), .A(n8876), .B(n8875), .ZN(n8877)
         );
  AOI21_X1 U10156 ( .B1(n9292), .B2(n8914), .A(n8877), .ZN(n8878) );
  OAI21_X1 U10157 ( .B1(n8879), .B2(n8947), .A(n8878), .ZN(P1_U3214) );
  XOR2_X1 U10158 ( .A(n8881), .B(n8880), .Z(n8887) );
  INV_X1 U10159 ( .A(n8882), .ZN(n9745) );
  NAND2_X1 U10160 ( .A1(n9745), .A2(n8940), .ZN(n8883) );
  NAND2_X1 U10161 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9036) );
  OAI211_X1 U10162 ( .C1(n9204), .C2(n8954), .A(n8883), .B(n9036), .ZN(n8885)
         );
  NOR2_X1 U10163 ( .A1(n9238), .A2(n8960), .ZN(n8884) );
  AOI211_X1 U10164 ( .C1(n9235), .C2(n8957), .A(n8885), .B(n8884), .ZN(n8886)
         );
  OAI21_X1 U10165 ( .B1(n8887), .B2(n8947), .A(n8886), .ZN(P1_U3217) );
  XOR2_X1 U10166 ( .A(n8889), .B(n8888), .Z(n8894) );
  NAND2_X1 U10167 ( .A1(n8957), .A2(n9208), .ZN(n8891) );
  AOI22_X1 U10168 ( .A1(n8928), .A2(n9059), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8890) );
  OAI211_X1 U10169 ( .C1(n9204), .C2(n8952), .A(n8891), .B(n8890), .ZN(n8892)
         );
  AOI21_X1 U10170 ( .B1(n9303), .B2(n8914), .A(n8892), .ZN(n8893) );
  OAI21_X1 U10171 ( .B1(n8894), .B2(n8947), .A(n8893), .ZN(P1_U3221) );
  XOR2_X1 U10172 ( .A(n8896), .B(n8895), .Z(n8901) );
  NAND2_X1 U10173 ( .A1(n8957), .A2(n9145), .ZN(n8898) );
  AOI22_X1 U10174 ( .A1(n9150), .A2(n8928), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8897) );
  OAI211_X1 U10175 ( .C1(n9175), .C2(n8952), .A(n8898), .B(n8897), .ZN(n8899)
         );
  AOI21_X1 U10176 ( .B1(n9279), .B2(n8914), .A(n8899), .ZN(n8900) );
  OAI21_X1 U10177 ( .B1(n8901), .B2(n8947), .A(n8900), .ZN(P1_U3223) );
  XOR2_X1 U10178 ( .A(n8903), .B(n8902), .Z(n8908) );
  NAND2_X1 U10179 ( .A1(n8957), .A2(n9163), .ZN(n8905) );
  INV_X1 U10180 ( .A(n9161), .ZN(n8962) );
  AOI22_X1 U10181 ( .A1(n8962), .A2(n8928), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8904) );
  OAI211_X1 U10182 ( .C1(n9190), .C2(n8952), .A(n8905), .B(n8904), .ZN(n8906)
         );
  AOI21_X1 U10183 ( .B1(n9285), .B2(n8914), .A(n8906), .ZN(n8907) );
  OAI21_X1 U10184 ( .B1(n8908), .B2(n8947), .A(n8907), .ZN(P1_U3227) );
  XOR2_X1 U10185 ( .A(n8910), .B(n8909), .Z(n8916) );
  NAND2_X1 U10186 ( .A1(n8957), .A2(n9218), .ZN(n8912) );
  INV_X1 U10187 ( .A(n9189), .ZN(n9225) );
  AOI22_X1 U10188 ( .A1(n9225), .A2(n8928), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8911) );
  OAI211_X1 U10189 ( .C1(n9055), .C2(n8952), .A(n8912), .B(n8911), .ZN(n8913)
         );
  AOI21_X1 U10190 ( .B1(n9306), .B2(n8914), .A(n8913), .ZN(n8915) );
  OAI21_X1 U10191 ( .B1(n8916), .B2(n8947), .A(n8915), .ZN(P1_U3231) );
  INV_X1 U10192 ( .A(n9296), .ZN(n9195) );
  AND2_X1 U10193 ( .A1(n8919), .A2(n8918), .ZN(n8920) );
  AOI21_X1 U10194 ( .B1(n8917), .B2(n8920), .A(n8922), .ZN(n8925) );
  INV_X1 U10195 ( .A(n8921), .ZN(n8924) );
  INV_X1 U10196 ( .A(n8922), .ZN(n8923) );
  OAI22_X1 U10197 ( .A1(n8925), .A2(n8924), .B1(n8923), .B2(n8917), .ZN(n8927)
         );
  NAND2_X1 U10198 ( .A1(n8927), .A2(n8926), .ZN(n8932) );
  AOI22_X1 U10199 ( .A1(n9060), .A2(n8928), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n8929) );
  OAI21_X1 U10200 ( .B1(n9189), .B2(n8952), .A(n8929), .ZN(n8930) );
  AOI21_X1 U10201 ( .B1(n8957), .B2(n9192), .A(n8930), .ZN(n8931) );
  OAI211_X1 U10202 ( .C1(n9195), .C2(n8960), .A(n8932), .B(n8931), .ZN(
        P1_U3233) );
  INV_X1 U10203 ( .A(n8935), .ZN(n8939) );
  AOI21_X1 U10204 ( .B1(n8935), .B2(n8934), .A(n8933), .ZN(n8936) );
  NOR2_X1 U10205 ( .A1(n8936), .A2(n8947), .ZN(n8937) );
  OAI21_X1 U10206 ( .B1(n8939), .B2(n8938), .A(n8937), .ZN(n8945) );
  NAND2_X1 U10207 ( .A1(n8940), .A2(n8963), .ZN(n8941) );
  NAND2_X1 U10208 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9010) );
  OAI211_X1 U10209 ( .C1(n9055), .C2(n8954), .A(n8941), .B(n9010), .ZN(n8942)
         );
  AOI21_X1 U10210 ( .B1(n8957), .B2(n8943), .A(n8942), .ZN(n8944) );
  OAI211_X1 U10211 ( .C1(n8946), .C2(n8960), .A(n8945), .B(n8944), .ZN(
        P1_U3236) );
  AOI21_X1 U10212 ( .B1(n8949), .B2(n8948), .A(n8947), .ZN(n8951) );
  NAND2_X1 U10213 ( .A1(n8951), .A2(n8950), .ZN(n8959) );
  NOR2_X1 U10214 ( .A1(n8952), .A2(n9161), .ZN(n8956) );
  OAI22_X1 U10215 ( .A1(n9135), .A2(n8954), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8953), .ZN(n8955) );
  AOI211_X1 U10216 ( .C1(n8957), .C2(n9129), .A(n8956), .B(n8955), .ZN(n8958)
         );
  OAI211_X1 U10217 ( .C1(n9131), .C2(n8960), .A(n8959), .B(n8958), .ZN(
        P1_U3238) );
  MUX2_X1 U10218 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9041), .S(P1_U4006), .Z(
        P1_U3586) );
  MUX2_X1 U10219 ( .A(n9085), .B(P1_DATAO_REG_30__SCAN_IN), .S(n8961), .Z(
        P1_U3585) );
  MUX2_X1 U10220 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n4703), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10221 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9065), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10222 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9150), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10223 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n8962), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10224 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n4688), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10225 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9060), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10226 ( .A(n9059), .B(P1_DATAO_REG_22__SCAN_IN), .S(n8961), .Z(
        P1_U3577) );
  MUX2_X1 U10227 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9225), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10228 ( .A(n9242), .B(P1_DATAO_REG_20__SCAN_IN), .S(n8961), .Z(
        P1_U3575) );
  MUX2_X1 U10229 ( .A(n9224), .B(P1_DATAO_REG_19__SCAN_IN), .S(n8961), .Z(
        P1_U3574) );
  MUX2_X1 U10230 ( .A(n8963), .B(P1_DATAO_REG_17__SCAN_IN), .S(n8961), .Z(
        P1_U3572) );
  MUX2_X1 U10231 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8964), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10232 ( .A(n8965), .B(P1_DATAO_REG_15__SCAN_IN), .S(n8961), .Z(
        P1_U3570) );
  MUX2_X1 U10233 ( .A(n8966), .B(P1_DATAO_REG_14__SCAN_IN), .S(n8961), .Z(
        P1_U3569) );
  MUX2_X1 U10234 ( .A(n9408), .B(P1_DATAO_REG_13__SCAN_IN), .S(n8961), .Z(
        P1_U3568) );
  MUX2_X1 U10235 ( .A(n8967), .B(P1_DATAO_REG_12__SCAN_IN), .S(n8961), .Z(
        P1_U3567) );
  MUX2_X1 U10236 ( .A(n9410), .B(P1_DATAO_REG_11__SCAN_IN), .S(n8961), .Z(
        P1_U3566) );
  MUX2_X1 U10237 ( .A(n8968), .B(P1_DATAO_REG_10__SCAN_IN), .S(n8961), .Z(
        P1_U3565) );
  MUX2_X1 U10238 ( .A(n8969), .B(P1_DATAO_REG_9__SCAN_IN), .S(n8961), .Z(
        P1_U3564) );
  MUX2_X1 U10239 ( .A(n8970), .B(P1_DATAO_REG_8__SCAN_IN), .S(n8961), .Z(
        P1_U3563) );
  MUX2_X1 U10240 ( .A(n8971), .B(P1_DATAO_REG_7__SCAN_IN), .S(n8961), .Z(
        P1_U3562) );
  MUX2_X1 U10241 ( .A(n8972), .B(P1_DATAO_REG_6__SCAN_IN), .S(n8961), .Z(
        P1_U3561) );
  MUX2_X1 U10242 ( .A(n6136), .B(P1_DATAO_REG_5__SCAN_IN), .S(n8961), .Z(
        P1_U3560) );
  MUX2_X1 U10243 ( .A(n8973), .B(P1_DATAO_REG_4__SCAN_IN), .S(n8961), .Z(
        P1_U3559) );
  MUX2_X1 U10244 ( .A(n8974), .B(P1_DATAO_REG_3__SCAN_IN), .S(n8961), .Z(
        P1_U3558) );
  MUX2_X1 U10245 ( .A(n8975), .B(P1_DATAO_REG_2__SCAN_IN), .S(n8961), .Z(
        P1_U3557) );
  MUX2_X1 U10246 ( .A(n8976), .B(P1_DATAO_REG_1__SCAN_IN), .S(n8961), .Z(
        P1_U3556) );
  OAI21_X1 U10247 ( .B1(n8979), .B2(n8978), .A(n8977), .ZN(n8980) );
  NAND2_X1 U10248 ( .A1(n8980), .A2(n9483), .ZN(n8991) );
  INV_X1 U10249 ( .A(n8981), .ZN(n8984) );
  NOR2_X1 U10250 ( .A1(n9027), .A2(n8982), .ZN(n8983) );
  AOI211_X1 U10251 ( .C1(P1_ADDR_REG_11__SCAN_IN), .C2(n9500), .A(n8984), .B(
        n8983), .ZN(n8990) );
  OAI21_X1 U10252 ( .B1(n8987), .B2(n8986), .A(n8985), .ZN(n8988) );
  NAND2_X1 U10253 ( .A1(n8988), .A2(n9497), .ZN(n8989) );
  NAND3_X1 U10254 ( .A1(n8991), .A2(n8990), .A3(n8989), .ZN(P1_U3252) );
  INV_X1 U10255 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9006) );
  AOI21_X1 U10256 ( .B1(n8996), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8992), .ZN(
        n8994) );
  XNOR2_X1 U10257 ( .A(n9013), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8993) );
  NOR2_X1 U10258 ( .A1(n8994), .A2(n8993), .ZN(n9007) );
  AOI211_X1 U10259 ( .C1(n8994), .C2(n8993), .A(n9007), .B(n9476), .ZN(n9004)
         );
  AOI21_X1 U10260 ( .B1(n8996), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8995), .ZN(
        n8999) );
  NAND2_X1 U10261 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9013), .ZN(n8997) );
  OAI21_X1 U10262 ( .B1(n9013), .B2(P1_REG2_REG_17__SCAN_IN), .A(n8997), .ZN(
        n8998) );
  NOR2_X1 U10263 ( .A1(n8999), .A2(n8998), .ZN(n9012) );
  AOI211_X1 U10264 ( .C1(n8999), .C2(n8998), .A(n9012), .B(n9490), .ZN(n9003)
         );
  INV_X1 U10265 ( .A(n9013), .ZN(n9001) );
  OAI21_X1 U10266 ( .B1(n9027), .B2(n9001), .A(n9000), .ZN(n9002) );
  NOR3_X1 U10267 ( .A1(n9004), .A2(n9003), .A3(n9002), .ZN(n9005) );
  OAI21_X1 U10268 ( .B1(n9038), .B2(n9006), .A(n9005), .ZN(P1_U3258) );
  INV_X1 U10269 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9021) );
  XOR2_X1 U10270 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9025), .Z(n9009) );
  AOI21_X1 U10271 ( .B1(n9013), .B2(P1_REG1_REG_17__SCAN_IN), .A(n9007), .ZN(
        n9008) );
  NAND2_X1 U10272 ( .A1(n9009), .A2(n9008), .ZN(n9024) );
  OAI21_X1 U10273 ( .B1(n9009), .B2(n9008), .A(n9024), .ZN(n9019) );
  INV_X1 U10274 ( .A(n9025), .ZN(n9011) );
  OAI21_X1 U10275 ( .B1(n9027), .B2(n9011), .A(n9010), .ZN(n9018) );
  NAND2_X1 U10276 ( .A1(n9025), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9014) );
  OAI21_X1 U10277 ( .B1(n9025), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9014), .ZN(
        n9015) );
  AOI211_X1 U10278 ( .C1(n9016), .C2(n9015), .A(n9022), .B(n9490), .ZN(n9017)
         );
  AOI211_X1 U10279 ( .C1(n9497), .C2(n9019), .A(n9018), .B(n9017), .ZN(n9020)
         );
  OAI21_X1 U10280 ( .B1(n9038), .B2(n9021), .A(n9020), .ZN(P1_U3259) );
  INV_X1 U10281 ( .A(n9032), .ZN(n9030) );
  INV_X1 U10282 ( .A(n9023), .ZN(n9029) );
  OAI21_X1 U10283 ( .B1(n9025), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9024), .ZN(
        n9026) );
  INV_X1 U10284 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9778) );
  XOR2_X1 U10285 ( .A(n9026), .B(n9778), .Z(n9031) );
  OAI21_X1 U10286 ( .B1(n9031), .B2(n9476), .A(n9027), .ZN(n9028) );
  AOI21_X1 U10287 ( .B1(n9030), .B2(n9029), .A(n9028), .ZN(n9035) );
  AOI22_X1 U10288 ( .A1(n9032), .A2(n9483), .B1(n9497), .B2(n9031), .ZN(n9034)
         );
  MUX2_X1 U10289 ( .A(n9035), .B(n9034), .S(n9033), .Z(n9037) );
  OAI211_X1 U10290 ( .C1(n4667), .C2(n9038), .A(n9037), .B(n9036), .ZN(
        P1_U3260) );
  INV_X1 U10291 ( .A(n9269), .ZN(n9116) );
  XNOR2_X1 U10292 ( .A(n9046), .B(n9043), .ZN(n9250) );
  NAND2_X1 U10293 ( .A1(n9430), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9042) );
  AND2_X1 U10294 ( .A1(n9039), .A2(P1_B_REG_SCAN_IN), .ZN(n9040) );
  NOR2_X1 U10295 ( .A1(n9376), .A2(n9040), .ZN(n9084) );
  NAND2_X1 U10296 ( .A1(n9041), .A2(n9084), .ZN(n9252) );
  OR2_X1 U10297 ( .A1(n9252), .A2(n9430), .ZN(n9047) );
  OAI211_X1 U10298 ( .C1(n9043), .C2(n9237), .A(n9042), .B(n9047), .ZN(n9044)
         );
  INV_X1 U10299 ( .A(n9044), .ZN(n9045) );
  OAI21_X1 U10300 ( .B1(n9250), .B2(n9088), .A(n9045), .ZN(P1_U3261) );
  AOI21_X1 U10301 ( .B1(n9087), .B2(n9049), .A(n9046), .ZN(n9251) );
  INV_X1 U10302 ( .A(n9251), .ZN(n9051) );
  INV_X1 U10303 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9802) );
  OAI21_X1 U10304 ( .B1(n7027), .B2(n9802), .A(n9047), .ZN(n9048) );
  AOI21_X1 U10305 ( .B1(n9049), .B2(n9415), .A(n9048), .ZN(n9050) );
  OAI21_X1 U10306 ( .B1(n9051), .B2(n9088), .A(n9050), .ZN(P1_U3262) );
  INV_X1 U10307 ( .A(n9264), .ZN(n9100) );
  NAND2_X1 U10308 ( .A1(n9312), .A2(n9224), .ZN(n9056) );
  INV_X1 U10309 ( .A(n9306), .ZN(n9220) );
  NAND2_X1 U10310 ( .A1(n9182), .A2(n9190), .ZN(n9061) );
  AOI22_X2 U10311 ( .A1(n9141), .A2(n9148), .B1(n9161), .B2(n9147), .ZN(n9127)
         );
  NAND2_X1 U10312 ( .A1(n9131), .A2(n9121), .ZN(n9064) );
  XNOR2_X1 U10313 ( .A(n9066), .B(n9082), .ZN(n9256) );
  INV_X1 U10314 ( .A(n9256), .ZN(n9095) );
  NAND2_X1 U10315 ( .A1(n9068), .A2(n9067), .ZN(n9240) );
  NAND2_X1 U10316 ( .A1(n9240), .A2(n9241), .ZN(n9239) );
  NAND3_X1 U10317 ( .A1(n9239), .A2(n9222), .A3(n9221), .ZN(n9070) );
  NAND2_X1 U10318 ( .A1(n9172), .A2(n9171), .ZN(n9073) );
  OAI21_X1 U10319 ( .B1(n9186), .B2(n9073), .A(n9072), .ZN(n9159) );
  INV_X1 U10320 ( .A(n9077), .ZN(n9078) );
  NOR2_X1 U10321 ( .A1(n9119), .A2(n9118), .ZN(n9117) );
  INV_X1 U10322 ( .A(n9079), .ZN(n9080) );
  NOR2_X1 U10323 ( .A1(n9117), .A2(n9080), .ZN(n9104) );
  NOR2_X1 U10324 ( .A1(n9104), .A2(n9103), .ZN(n9102) );
  INV_X1 U10325 ( .A(n9082), .ZN(n9083) );
  AOI22_X1 U10326 ( .A1(n4703), .A2(n9409), .B1(n9085), .B2(n9084), .ZN(n9086)
         );
  OAI21_X1 U10327 ( .B1(n9097), .B2(n9091), .A(n9087), .ZN(n9257) );
  NOR2_X1 U10328 ( .A1(n9257), .A2(n9088), .ZN(n9093) );
  AOI22_X1 U10329 ( .A1(n9386), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9089), .B2(
        n9414), .ZN(n9090) );
  OAI21_X1 U10330 ( .B1(n9091), .B2(n9237), .A(n9090), .ZN(n9092) );
  AOI211_X1 U10331 ( .C1(n9255), .C2(n7027), .A(n9093), .B(n9092), .ZN(n9094)
         );
  OAI21_X1 U10332 ( .B1(n9095), .B2(n9247), .A(n9094), .ZN(P1_U3355) );
  OAI21_X1 U10333 ( .B1(n4303), .B2(n9103), .A(n9096), .ZN(n9268) );
  AOI21_X1 U10334 ( .B1(n9264), .B2(n9111), .A(n9097), .ZN(n9265) );
  AOI22_X1 U10335 ( .A1(n9430), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9098), .B2(
        n9414), .ZN(n9099) );
  OAI21_X1 U10336 ( .B1(n9100), .B2(n9237), .A(n9099), .ZN(n9101) );
  AOI21_X1 U10337 ( .B1(n9265), .B2(n9229), .A(n9101), .ZN(n9109) );
  AOI211_X1 U10338 ( .C1(n9104), .C2(n9103), .A(n9203), .B(n9102), .ZN(n9107)
         );
  OAI22_X1 U10339 ( .A1(n9135), .A2(n9378), .B1(n9105), .B2(n9376), .ZN(n9106)
         );
  NOR2_X1 U10340 ( .A1(n9107), .A2(n9106), .ZN(n9267) );
  OR2_X1 U10341 ( .A1(n9267), .A2(n9430), .ZN(n9108) );
  OAI211_X1 U10342 ( .C1(n9268), .C2(n9247), .A(n9109), .B(n9108), .ZN(
        P1_U3263) );
  XOR2_X1 U10343 ( .A(n9118), .B(n9110), .Z(n9273) );
  INV_X1 U10344 ( .A(n9128), .ZN(n9113) );
  INV_X1 U10345 ( .A(n9111), .ZN(n9112) );
  AOI21_X1 U10346 ( .B1(n9269), .B2(n9113), .A(n9112), .ZN(n9270) );
  AOI22_X1 U10347 ( .A1(n9386), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9114), .B2(
        n9414), .ZN(n9115) );
  OAI21_X1 U10348 ( .B1(n9116), .B2(n9237), .A(n9115), .ZN(n9125) );
  AOI211_X1 U10349 ( .C1(n9119), .C2(n9118), .A(n9203), .B(n9117), .ZN(n9123)
         );
  OAI22_X1 U10350 ( .A1(n9121), .A2(n9378), .B1(n9120), .B2(n9376), .ZN(n9122)
         );
  NOR2_X1 U10351 ( .A1(n9123), .A2(n9122), .ZN(n9272) );
  NOR2_X1 U10352 ( .A1(n9272), .A2(n9430), .ZN(n9124) );
  AOI211_X1 U10353 ( .C1(n9229), .C2(n9270), .A(n9125), .B(n9124), .ZN(n9126)
         );
  OAI21_X1 U10354 ( .B1(n9273), .B2(n9247), .A(n9126), .ZN(P1_U3264) );
  XNOR2_X1 U10355 ( .A(n9127), .B(n9133), .ZN(n9278) );
  AOI211_X1 U10356 ( .C1(n9275), .C2(n9142), .A(n9542), .B(n9128), .ZN(n9274)
         );
  AOI22_X1 U10357 ( .A1(n9386), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9129), .B2(
        n9414), .ZN(n9130) );
  OAI21_X1 U10358 ( .B1(n9131), .B2(n9237), .A(n9130), .ZN(n9139) );
  AOI211_X1 U10359 ( .C1(n9134), .C2(n9133), .A(n9203), .B(n9132), .ZN(n9137)
         );
  OAI22_X1 U10360 ( .A1(n9161), .A2(n9378), .B1(n9135), .B2(n9376), .ZN(n9136)
         );
  NOR2_X1 U10361 ( .A1(n9137), .A2(n9136), .ZN(n9277) );
  NOR2_X1 U10362 ( .A1(n9277), .A2(n9386), .ZN(n9138) );
  AOI211_X1 U10363 ( .C1(n9274), .C2(n9426), .A(n9139), .B(n9138), .ZN(n9140)
         );
  OAI21_X1 U10364 ( .B1(n9278), .B2(n9247), .A(n9140), .ZN(P1_U3265) );
  XOR2_X1 U10365 ( .A(n9148), .B(n9141), .Z(n9283) );
  INV_X1 U10366 ( .A(n9162), .ZN(n9144) );
  INV_X1 U10367 ( .A(n9142), .ZN(n9143) );
  AOI21_X1 U10368 ( .B1(n9279), .B2(n9144), .A(n9143), .ZN(n9280) );
  AOI22_X1 U10369 ( .A1(n9386), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9145), .B2(
        n9414), .ZN(n9146) );
  OAI21_X1 U10370 ( .B1(n9147), .B2(n9237), .A(n9146), .ZN(n9153) );
  XNOR2_X1 U10371 ( .A(n9149), .B(n9148), .ZN(n9151) );
  AOI222_X1 U10372 ( .A1(n9412), .A2(n9151), .B1(n9150), .B2(n9407), .C1(n4688), .C2(n9409), .ZN(n9282) );
  NOR2_X1 U10373 ( .A1(n9282), .A2(n9386), .ZN(n9152) );
  AOI211_X1 U10374 ( .C1(n9280), .C2(n9229), .A(n9153), .B(n9152), .ZN(n9154)
         );
  OAI21_X1 U10375 ( .B1(n9283), .B2(n9247), .A(n9154), .ZN(P1_U3266) );
  XNOR2_X1 U10376 ( .A(n9156), .B(n9155), .ZN(n9289) );
  AOI21_X1 U10377 ( .B1(n9159), .B2(n9158), .A(n9157), .ZN(n9160) );
  OAI222_X1 U10378 ( .A1(n9376), .A2(n9161), .B1(n9378), .B2(n9190), .C1(n9203), .C2(n9160), .ZN(n9284) );
  AOI21_X1 U10379 ( .B1(n9285), .B2(n9176), .A(n9162), .ZN(n9286) );
  NAND2_X1 U10380 ( .A1(n9286), .A2(n9229), .ZN(n9165) );
  AOI22_X1 U10381 ( .A1(n9430), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9163), .B2(
        n9414), .ZN(n9164) );
  OAI211_X1 U10382 ( .C1(n9166), .C2(n9237), .A(n9165), .B(n9164), .ZN(n9167)
         );
  AOI21_X1 U10383 ( .B1(n9284), .B2(n7027), .A(n9167), .ZN(n9168) );
  OAI21_X1 U10384 ( .B1(n9289), .B2(n9247), .A(n9168), .ZN(P1_U3267) );
  XNOR2_X1 U10385 ( .A(n9170), .B(n9169), .ZN(n9294) );
  NOR2_X1 U10386 ( .A1(n9186), .A2(n4369), .ZN(n9173) );
  XNOR2_X1 U10387 ( .A(n9173), .B(n9172), .ZN(n9174) );
  OAI222_X1 U10388 ( .A1(n9376), .A2(n9175), .B1(n9378), .B2(n9205), .C1(n9174), .C2(n9203), .ZN(n9290) );
  INV_X1 U10389 ( .A(n9191), .ZN(n9178) );
  INV_X1 U10390 ( .A(n9176), .ZN(n9177) );
  AOI211_X1 U10391 ( .C1(n9292), .C2(n9178), .A(n9542), .B(n9177), .ZN(n9291)
         );
  NAND2_X1 U10392 ( .A1(n9291), .A2(n9426), .ZN(n9181) );
  AOI22_X1 U10393 ( .A1(n9430), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9179), .B2(
        n9414), .ZN(n9180) );
  OAI211_X1 U10394 ( .C1(n9182), .C2(n9237), .A(n9181), .B(n9180), .ZN(n9183)
         );
  AOI21_X1 U10395 ( .B1(n9290), .B2(n7027), .A(n9183), .ZN(n9184) );
  OAI21_X1 U10396 ( .B1(n9294), .B2(n9247), .A(n9184), .ZN(P1_U3268) );
  XOR2_X1 U10397 ( .A(n9187), .B(n9185), .Z(n9300) );
  AOI21_X1 U10398 ( .B1(n4281), .B2(n9187), .A(n9186), .ZN(n9188) );
  OAI222_X1 U10399 ( .A1(n9376), .A2(n9190), .B1(n9378), .B2(n9189), .C1(n9203), .C2(n9188), .ZN(n9295) );
  AOI21_X1 U10400 ( .B1(n9296), .B2(n9206), .A(n9191), .ZN(n9297) );
  NAND2_X1 U10401 ( .A1(n9297), .A2(n9229), .ZN(n9194) );
  AOI22_X1 U10402 ( .A1(n9430), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9192), .B2(
        n9414), .ZN(n9193) );
  OAI211_X1 U10403 ( .C1(n9195), .C2(n9237), .A(n9194), .B(n9193), .ZN(n9196)
         );
  AOI21_X1 U10404 ( .B1(n9295), .B2(n7027), .A(n9196), .ZN(n9197) );
  OAI21_X1 U10405 ( .B1(n9300), .B2(n9247), .A(n9197), .ZN(P1_U3269) );
  XNOR2_X1 U10406 ( .A(n9198), .B(n9201), .ZN(n9305) );
  AOI22_X1 U10407 ( .A1(n9303), .A2(n9415), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9386), .ZN(n9215) );
  AOI21_X1 U10408 ( .B1(n9201), .B2(n9200), .A(n9199), .ZN(n9202) );
  OAI222_X1 U10409 ( .A1(n9376), .A2(n9205), .B1(n9378), .B2(n9204), .C1(n9203), .C2(n9202), .ZN(n9301) );
  INV_X1 U10410 ( .A(n9206), .ZN(n9207) );
  AOI211_X1 U10411 ( .C1(n9303), .C2(n9217), .A(n9542), .B(n9207), .ZN(n9302)
         );
  INV_X1 U10412 ( .A(n9302), .ZN(n9212) );
  INV_X1 U10413 ( .A(n9208), .ZN(n9210) );
  OAI22_X1 U10414 ( .A1(n9212), .A2(n9211), .B1(n9210), .B2(n9209), .ZN(n9213)
         );
  OAI21_X1 U10415 ( .B1(n9301), .B2(n9213), .A(n7027), .ZN(n9214) );
  OAI211_X1 U10416 ( .C1(n9305), .C2(n9247), .A(n9215), .B(n9214), .ZN(
        P1_U3270) );
  XOR2_X1 U10417 ( .A(n9222), .B(n9216), .Z(n9310) );
  AOI21_X1 U10418 ( .B1(n9306), .B2(n9233), .A(n4410), .ZN(n9307) );
  AOI22_X1 U10419 ( .A1(n9386), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9218), .B2(
        n9414), .ZN(n9219) );
  OAI21_X1 U10420 ( .B1(n9220), .B2(n9237), .A(n9219), .ZN(n9228) );
  NAND2_X1 U10421 ( .A1(n9239), .A2(n9221), .ZN(n9223) );
  XNOR2_X1 U10422 ( .A(n9223), .B(n9222), .ZN(n9226) );
  AOI222_X1 U10423 ( .A1(n9412), .A2(n9226), .B1(n9225), .B2(n9407), .C1(n9224), .C2(n9409), .ZN(n9309) );
  NOR2_X1 U10424 ( .A1(n9309), .A2(n9430), .ZN(n9227) );
  AOI211_X1 U10425 ( .C1(n9307), .C2(n9229), .A(n9228), .B(n9227), .ZN(n9230)
         );
  OAI21_X1 U10426 ( .B1(n9310), .B2(n9247), .A(n9230), .ZN(P1_U3271) );
  XNOR2_X1 U10427 ( .A(n9231), .B(n9241), .ZN(n9315) );
  INV_X1 U10428 ( .A(n9232), .ZN(n9234) );
  AOI211_X1 U10429 ( .C1(n9312), .C2(n9234), .A(n9542), .B(n4411), .ZN(n9311)
         );
  AOI22_X1 U10430 ( .A1(n9386), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9414), .B2(
        n9235), .ZN(n9236) );
  OAI21_X1 U10431 ( .B1(n9238), .B2(n9237), .A(n9236), .ZN(n9245) );
  OAI21_X1 U10432 ( .B1(n9241), .B2(n9240), .A(n9239), .ZN(n9243) );
  AOI222_X1 U10433 ( .A1(n9412), .A2(n9243), .B1(n9242), .B2(n9407), .C1(n9745), .C2(n9409), .ZN(n9314) );
  NOR2_X1 U10434 ( .A1(n9314), .A2(n9430), .ZN(n9244) );
  AOI211_X1 U10435 ( .C1(n9311), .C2(n9426), .A(n9245), .B(n9244), .ZN(n9246)
         );
  OAI21_X1 U10436 ( .B1(n9315), .B2(n9247), .A(n9246), .ZN(P1_U3272) );
  NAND2_X1 U10437 ( .A1(n9248), .A2(n9520), .ZN(n9249) );
  OAI211_X1 U10438 ( .C1(n9250), .C2(n9542), .A(n9252), .B(n9249), .ZN(n9342)
         );
  MUX2_X1 U10439 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9342), .S(n9562), .Z(
        P1_U3554) );
  NAND2_X1 U10440 ( .A1(n9251), .A2(n9423), .ZN(n9253) );
  OAI211_X1 U10441 ( .C1(n9254), .C2(n9540), .A(n9253), .B(n9252), .ZN(n9343)
         );
  MUX2_X1 U10442 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9343), .S(n9562), .Z(
        P1_U3553) );
  NAND2_X1 U10443 ( .A1(n9256), .A2(n9546), .ZN(n9262) );
  NOR2_X1 U10444 ( .A1(n9257), .A2(n9542), .ZN(n9260) );
  NAND3_X1 U10445 ( .A1(n9263), .A2(n9262), .A3(n9261), .ZN(n9344) );
  MUX2_X1 U10446 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9344), .S(n9562), .Z(
        P1_U3552) );
  AOI22_X1 U10447 ( .A1(n9265), .A2(n9423), .B1(n9520), .B2(n9264), .ZN(n9266)
         );
  OAI211_X1 U10448 ( .C1(n9268), .C2(n9517), .A(n9267), .B(n9266), .ZN(n9345)
         );
  MUX2_X1 U10449 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9345), .S(n9562), .Z(
        P1_U3551) );
  AOI22_X1 U10450 ( .A1(n9270), .A2(n9423), .B1(n9520), .B2(n9269), .ZN(n9271)
         );
  OAI211_X1 U10451 ( .C1(n9273), .C2(n9517), .A(n9272), .B(n9271), .ZN(n9346)
         );
  MUX2_X1 U10452 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9346), .S(n9562), .Z(
        P1_U3550) );
  AOI21_X1 U10453 ( .B1(n9520), .B2(n9275), .A(n9274), .ZN(n9276) );
  OAI211_X1 U10454 ( .C1(n9278), .C2(n9517), .A(n9277), .B(n9276), .ZN(n9347)
         );
  MUX2_X1 U10455 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9347), .S(n9562), .Z(
        P1_U3549) );
  AOI22_X1 U10456 ( .A1(n9280), .A2(n9423), .B1(n9520), .B2(n9279), .ZN(n9281)
         );
  OAI211_X1 U10457 ( .C1(n9283), .C2(n9517), .A(n9282), .B(n9281), .ZN(n9348)
         );
  MUX2_X1 U10458 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9348), .S(n9562), .Z(
        P1_U3548) );
  INV_X1 U10459 ( .A(n9284), .ZN(n9288) );
  AOI22_X1 U10460 ( .A1(n9286), .A2(n9423), .B1(n9520), .B2(n9285), .ZN(n9287)
         );
  OAI211_X1 U10461 ( .C1(n9289), .C2(n9517), .A(n9288), .B(n9287), .ZN(n9349)
         );
  MUX2_X1 U10462 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9349), .S(n9562), .Z(
        P1_U3547) );
  AOI211_X1 U10463 ( .C1(n9520), .C2(n9292), .A(n9291), .B(n9290), .ZN(n9293)
         );
  OAI21_X1 U10464 ( .B1(n9294), .B2(n9517), .A(n9293), .ZN(n9350) );
  MUX2_X1 U10465 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9350), .S(n9562), .Z(
        P1_U3546) );
  INV_X1 U10466 ( .A(n9295), .ZN(n9299) );
  AOI22_X1 U10467 ( .A1(n9297), .A2(n9423), .B1(n9520), .B2(n9296), .ZN(n9298)
         );
  OAI211_X1 U10468 ( .C1(n9300), .C2(n9517), .A(n9299), .B(n9298), .ZN(n9351)
         );
  MUX2_X1 U10469 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9351), .S(n9562), .Z(
        P1_U3545) );
  AOI211_X1 U10470 ( .C1(n9520), .C2(n9303), .A(n9302), .B(n9301), .ZN(n9304)
         );
  OAI21_X1 U10471 ( .B1(n9305), .B2(n9517), .A(n9304), .ZN(n9352) );
  MUX2_X1 U10472 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9352), .S(n9562), .Z(
        P1_U3544) );
  AOI22_X1 U10473 ( .A1(n9307), .A2(n9423), .B1(n9520), .B2(n9306), .ZN(n9308)
         );
  OAI211_X1 U10474 ( .C1(n9310), .C2(n9517), .A(n9309), .B(n9308), .ZN(n9353)
         );
  MUX2_X1 U10475 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9353), .S(n9562), .Z(
        P1_U3543) );
  AOI21_X1 U10476 ( .B1(n9520), .B2(n9312), .A(n9311), .ZN(n9313) );
  OAI211_X1 U10477 ( .C1(n9315), .C2(n9517), .A(n9314), .B(n9313), .ZN(n9354)
         );
  MUX2_X1 U10478 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9354), .S(n9562), .Z(
        P1_U3542) );
  AOI22_X1 U10479 ( .A1(n9317), .A2(n9423), .B1(n9520), .B2(n9316), .ZN(n9318)
         );
  OAI211_X1 U10480 ( .C1(n9320), .C2(n9517), .A(n9319), .B(n9318), .ZN(n9355)
         );
  MUX2_X1 U10481 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9355), .S(n9562), .Z(
        P1_U3541) );
  AOI211_X1 U10482 ( .C1(n9520), .C2(n9323), .A(n9322), .B(n9321), .ZN(n9324)
         );
  OAI21_X1 U10483 ( .B1(n9325), .B2(n9517), .A(n9324), .ZN(n9356) );
  MUX2_X1 U10484 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9356), .S(n9562), .Z(
        P1_U3540) );
  AOI211_X1 U10485 ( .C1(n9520), .C2(n9328), .A(n9327), .B(n9326), .ZN(n9329)
         );
  OAI21_X1 U10486 ( .B1(n9330), .B2(n9517), .A(n9329), .ZN(n9357) );
  MUX2_X1 U10487 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9357), .S(n9562), .Z(
        P1_U3539) );
  AOI22_X1 U10488 ( .A1(n9332), .A2(n9423), .B1(n9520), .B2(n9331), .ZN(n9333)
         );
  OAI211_X1 U10489 ( .C1(n9336), .C2(n9335), .A(n9334), .B(n9333), .ZN(n9358)
         );
  MUX2_X1 U10490 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9358), .S(n9562), .Z(
        P1_U3538) );
  AOI211_X1 U10491 ( .C1(n9520), .C2(n9339), .A(n9338), .B(n9337), .ZN(n9340)
         );
  OAI21_X1 U10492 ( .B1(n9341), .B2(n9517), .A(n9340), .ZN(n9359) );
  MUX2_X1 U10493 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9359), .S(n9562), .Z(
        P1_U3537) );
  MUX2_X1 U10494 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9342), .S(n9550), .Z(
        P1_U3522) );
  MUX2_X1 U10495 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9343), .S(n9550), .Z(
        P1_U3521) );
  MUX2_X1 U10496 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9344), .S(n9550), .Z(
        P1_U3520) );
  MUX2_X1 U10497 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9345), .S(n9550), .Z(
        P1_U3519) );
  MUX2_X1 U10498 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9346), .S(n9550), .Z(
        P1_U3518) );
  MUX2_X1 U10499 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9347), .S(n9550), .Z(
        P1_U3517) );
  MUX2_X1 U10500 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9348), .S(n9550), .Z(
        P1_U3516) );
  MUX2_X1 U10501 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9349), .S(n9550), .Z(
        P1_U3515) );
  MUX2_X1 U10502 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9350), .S(n9550), .Z(
        P1_U3514) );
  MUX2_X1 U10503 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9351), .S(n9550), .Z(
        P1_U3513) );
  MUX2_X1 U10504 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9352), .S(n9550), .Z(
        P1_U3512) );
  MUX2_X1 U10505 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9353), .S(n9550), .Z(
        P1_U3511) );
  MUX2_X1 U10506 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9354), .S(n9550), .Z(
        P1_U3510) );
  MUX2_X1 U10507 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9355), .S(n9550), .Z(
        P1_U3508) );
  MUX2_X1 U10508 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9356), .S(n9550), .Z(
        P1_U3505) );
  MUX2_X1 U10509 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9357), .S(n9550), .Z(
        P1_U3502) );
  MUX2_X1 U10510 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9358), .S(n9550), .Z(
        P1_U3499) );
  MUX2_X1 U10511 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9359), .S(n9550), .Z(
        P1_U3496) );
  MUX2_X1 U10512 ( .A(P1_D_REG_1__SCAN_IN), .B(n9361), .S(n9360), .Z(P1_U3441)
         );
  NOR4_X1 U10513 ( .A1(n9362), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5519), .A4(
        P1_U3084), .ZN(n9363) );
  AOI21_X1 U10514 ( .B1(n9366), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9363), .ZN(
        n9364) );
  OAI21_X1 U10515 ( .B1(n9365), .B2(n8334), .A(n9364), .ZN(P1_U3322) );
  AOI22_X1 U10516 ( .A1(n9367), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9366), .ZN(n9368) );
  OAI21_X1 U10517 ( .B1(n9369), .B2(n8334), .A(n9368), .ZN(P1_U3323) );
  MUX2_X1 U10518 ( .A(n9370), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10519 ( .A(n9371), .ZN(n9372) );
  AOI21_X1 U10520 ( .B1(n9374), .B2(n9373), .A(n9372), .ZN(n9375) );
  XNOR2_X1 U10521 ( .A(n9375), .B(n9380), .ZN(n9385) );
  OAI22_X1 U10522 ( .A1(n9379), .A2(n9378), .B1(n9377), .B2(n9376), .ZN(n9384)
         );
  XOR2_X1 U10523 ( .A(n9381), .B(n9380), .Z(n9389) );
  NOR2_X1 U10524 ( .A1(n9389), .A2(n9382), .ZN(n9383) );
  AOI211_X1 U10525 ( .C1(n9385), .C2(n9412), .A(n9384), .B(n9383), .ZN(n9399)
         );
  AOI222_X1 U10526 ( .A1(n9388), .A2(n9415), .B1(n9387), .B2(n9414), .C1(
        P1_REG2_REG_10__SCAN_IN), .C2(n9386), .ZN(n9396) );
  INV_X1 U10527 ( .A(n9389), .ZN(n9402) );
  INV_X1 U10528 ( .A(n9390), .ZN(n9391) );
  OAI211_X1 U10529 ( .C1(n9398), .C2(n9392), .A(n9391), .B(n9423), .ZN(n9397)
         );
  INV_X1 U10530 ( .A(n9397), .ZN(n9393) );
  AOI22_X1 U10531 ( .A1(n9402), .A2(n9394), .B1(n9426), .B2(n9393), .ZN(n9395)
         );
  OAI211_X1 U10532 ( .C1(n9430), .C2(n9399), .A(n9396), .B(n9395), .ZN(
        P1_U3281) );
  OAI21_X1 U10533 ( .B1(n9398), .B2(n9540), .A(n9397), .ZN(n9401) );
  INV_X1 U10534 ( .A(n9399), .ZN(n9400) );
  AOI211_X1 U10535 ( .C1(n9538), .C2(n9402), .A(n9401), .B(n9400), .ZN(n9405)
         );
  INV_X1 U10536 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9403) );
  AOI22_X1 U10537 ( .A1(n9550), .A2(n9405), .B1(n9403), .B2(n9548), .ZN(
        P1_U3484) );
  AOI22_X1 U10538 ( .A1(n9562), .A2(n9405), .B1(n9404), .B2(n9559), .ZN(
        P1_U3533) );
  XNOR2_X1 U10539 ( .A(n9406), .B(n9418), .ZN(n9411) );
  AOI222_X1 U10540 ( .A1(n9412), .A2(n9411), .B1(n9410), .B2(n9409), .C1(n9408), .C2(n9407), .ZN(n9432) );
  AOI222_X1 U10541 ( .A1(n9416), .A2(n9415), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9430), .C1(n9414), .C2(n9413), .ZN(n9429) );
  OAI21_X1 U10542 ( .B1(n9419), .B2(n9418), .A(n9417), .ZN(n9420) );
  INV_X1 U10543 ( .A(n9420), .ZN(n9435) );
  INV_X1 U10544 ( .A(n9421), .ZN(n9424) );
  OAI211_X1 U10545 ( .C1(n9424), .C2(n9433), .A(n9423), .B(n9422), .ZN(n9431)
         );
  INV_X1 U10546 ( .A(n9431), .ZN(n9425) );
  AOI22_X1 U10547 ( .A1(n9435), .A2(n9427), .B1(n9426), .B2(n9425), .ZN(n9428)
         );
  OAI211_X1 U10548 ( .C1(n9430), .C2(n9432), .A(n9429), .B(n9428), .ZN(
        P1_U3279) );
  OAI211_X1 U10549 ( .C1(n9433), .C2(n9540), .A(n9432), .B(n9431), .ZN(n9434)
         );
  AOI21_X1 U10550 ( .B1(n9435), .B2(n9546), .A(n9434), .ZN(n9445) );
  INV_X1 U10551 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9436) );
  AOI22_X1 U10552 ( .A1(n9562), .A2(n9445), .B1(n9436), .B2(n9559), .ZN(
        P1_U3535) );
  INV_X1 U10553 ( .A(n9437), .ZN(n9442) );
  OAI22_X1 U10554 ( .A1(n9439), .A2(n9542), .B1(n9438), .B2(n9540), .ZN(n9441)
         );
  AOI211_X1 U10555 ( .C1(n9538), .C2(n9442), .A(n9441), .B(n9440), .ZN(n9446)
         );
  AOI22_X1 U10556 ( .A1(n9562), .A2(n9446), .B1(n9443), .B2(n9559), .ZN(
        P1_U3534) );
  INV_X1 U10557 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9444) );
  AOI22_X1 U10558 ( .A1(n9550), .A2(n9445), .B1(n9444), .B2(n9548), .ZN(
        P1_U3490) );
  INV_X1 U10559 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9880) );
  AOI22_X1 U10560 ( .A1(n9550), .A2(n9446), .B1(n9880), .B2(n9548), .ZN(
        P1_U3487) );
  XNOR2_X1 U10561 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10562 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  AOI211_X1 U10563 ( .C1(n9449), .C2(n9448), .A(n9447), .B(n9476), .ZN(n9457)
         );
  OR3_X1 U10564 ( .A1(n9452), .A2(n9451), .A3(n9450), .ZN(n9453) );
  AOI21_X1 U10565 ( .B1(n9454), .B2(n9453), .A(n9490), .ZN(n9455) );
  NOR3_X1 U10566 ( .A1(n9457), .A2(n9456), .A3(n9455), .ZN(n9460) );
  AOI22_X1 U10567 ( .A1(n9500), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9499), .B2(
        n9458), .ZN(n9459) );
  NAND2_X1 U10568 ( .A1(n9460), .A2(n9459), .ZN(P1_U3246) );
  OAI21_X1 U10569 ( .B1(n9463), .B2(n9462), .A(n9461), .ZN(n9469) );
  AOI211_X1 U10570 ( .C1(n9466), .C2(n9465), .A(n9464), .B(n9490), .ZN(n9467)
         );
  AOI211_X1 U10571 ( .C1(n9469), .C2(n9497), .A(n9468), .B(n9467), .ZN(n9472)
         );
  AOI22_X1 U10572 ( .A1(n9500), .A2(P1_ADDR_REG_6__SCAN_IN), .B1(n9499), .B2(
        n9470), .ZN(n9471) );
  NAND2_X1 U10573 ( .A1(n9472), .A2(n9471), .ZN(P1_U3247) );
  OAI21_X1 U10574 ( .B1(n9475), .B2(n9474), .A(n9473), .ZN(n9482) );
  AOI211_X1 U10575 ( .C1(n9479), .C2(n9478), .A(n9477), .B(n9476), .ZN(n9480)
         );
  AOI211_X1 U10576 ( .C1(n9483), .C2(n9482), .A(n9481), .B(n9480), .ZN(n9486)
         );
  AOI22_X1 U10577 ( .A1(n9500), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n9499), .B2(
        n9484), .ZN(n9485) );
  NAND2_X1 U10578 ( .A1(n9486), .A2(n9485), .ZN(P1_U3249) );
  OAI21_X1 U10579 ( .B1(n9489), .B2(n9488), .A(n9487), .ZN(n9496) );
  AOI211_X1 U10580 ( .C1(n9493), .C2(n9492), .A(n9491), .B(n9490), .ZN(n9494)
         );
  AOI211_X1 U10581 ( .C1(n9497), .C2(n9496), .A(n9495), .B(n9494), .ZN(n9502)
         );
  AOI22_X1 U10582 ( .A1(n9500), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(n9499), .B2(
        n9498), .ZN(n9501) );
  NAND2_X1 U10583 ( .A1(n9502), .A2(n9501), .ZN(P1_U3250) );
  INV_X1 U10584 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9870) );
  NOR2_X1 U10585 ( .A1(n9503), .A2(n9870), .ZN(P1_U3292) );
  AND2_X1 U10586 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9504), .ZN(P1_U3293) );
  AND2_X1 U10587 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9504), .ZN(P1_U3294) );
  AND2_X1 U10588 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9504), .ZN(P1_U3295) );
  AND2_X1 U10589 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9504), .ZN(P1_U3296) );
  AND2_X1 U10590 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9504), .ZN(P1_U3297) );
  AND2_X1 U10591 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9504), .ZN(P1_U3298) );
  AND2_X1 U10592 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9504), .ZN(P1_U3299) );
  AND2_X1 U10593 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9504), .ZN(P1_U3300) );
  AND2_X1 U10594 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9504), .ZN(P1_U3301) );
  AND2_X1 U10595 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9504), .ZN(P1_U3302) );
  AND2_X1 U10596 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9504), .ZN(P1_U3303) );
  AND2_X1 U10597 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9504), .ZN(P1_U3304) );
  INV_X1 U10598 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n9836) );
  NOR2_X1 U10599 ( .A1(n9503), .A2(n9836), .ZN(P1_U3305) );
  AND2_X1 U10600 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9504), .ZN(P1_U3306) );
  INV_X1 U10601 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9878) );
  NOR2_X1 U10602 ( .A1(n9503), .A2(n9878), .ZN(P1_U3307) );
  AND2_X1 U10603 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9504), .ZN(P1_U3308) );
  AND2_X1 U10604 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9504), .ZN(P1_U3309) );
  AND2_X1 U10605 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9504), .ZN(P1_U3310) );
  AND2_X1 U10606 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9504), .ZN(P1_U3311) );
  AND2_X1 U10607 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9504), .ZN(P1_U3312) );
  AND2_X1 U10608 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9504), .ZN(P1_U3313) );
  INV_X1 U10609 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9855) );
  NOR2_X1 U10610 ( .A1(n9503), .A2(n9855), .ZN(P1_U3314) );
  AND2_X1 U10611 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9504), .ZN(P1_U3315) );
  AND2_X1 U10612 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9504), .ZN(P1_U3316) );
  AND2_X1 U10613 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9504), .ZN(P1_U3317) );
  AND2_X1 U10614 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9504), .ZN(P1_U3318) );
  AND2_X1 U10615 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9504), .ZN(P1_U3319) );
  AND2_X1 U10616 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9504), .ZN(P1_U3320) );
  AND2_X1 U10617 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9504), .ZN(P1_U3321) );
  OAI21_X1 U10618 ( .B1(n9506), .B2(n9542), .A(n9505), .ZN(n9508) );
  AOI211_X1 U10619 ( .C1(n9546), .C2(n9509), .A(n9508), .B(n9507), .ZN(n9551)
         );
  INV_X1 U10620 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9510) );
  AOI22_X1 U10621 ( .A1(n9550), .A2(n9551), .B1(n9510), .B2(n9548), .ZN(
        P1_U3460) );
  OAI22_X1 U10622 ( .A1(n9512), .A2(n9542), .B1(n9511), .B2(n9540), .ZN(n9514)
         );
  AOI211_X1 U10623 ( .C1(n9538), .C2(n9515), .A(n9514), .B(n9513), .ZN(n9553)
         );
  INV_X1 U10624 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9516) );
  AOI22_X1 U10625 ( .A1(n9550), .A2(n9553), .B1(n9516), .B2(n9548), .ZN(
        P1_U3466) );
  OR2_X1 U10626 ( .A1(n9518), .A2(n9517), .ZN(n9524) );
  NAND2_X1 U10627 ( .A1(n9520), .A2(n9519), .ZN(n9521) );
  AND2_X1 U10628 ( .A1(n9522), .A2(n9521), .ZN(n9523) );
  AND3_X1 U10629 ( .A1(n9525), .A2(n9524), .A3(n9523), .ZN(n9555) );
  INV_X1 U10630 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9526) );
  AOI22_X1 U10631 ( .A1(n9550), .A2(n9555), .B1(n9526), .B2(n9548), .ZN(
        P1_U3469) );
  OAI22_X1 U10632 ( .A1(n9528), .A2(n9542), .B1(n9527), .B2(n9540), .ZN(n9530)
         );
  AOI211_X1 U10633 ( .C1(n9538), .C2(n9531), .A(n9530), .B(n9529), .ZN(n9556)
         );
  INV_X1 U10634 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9532) );
  AOI22_X1 U10635 ( .A1(n9550), .A2(n9556), .B1(n9532), .B2(n9548), .ZN(
        P1_U3472) );
  OAI22_X1 U10636 ( .A1(n9534), .A2(n9542), .B1(n9533), .B2(n9540), .ZN(n9536)
         );
  AOI211_X1 U10637 ( .C1(n9538), .C2(n9537), .A(n9536), .B(n9535), .ZN(n9558)
         );
  INV_X1 U10638 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9539) );
  AOI22_X1 U10639 ( .A1(n9550), .A2(n9558), .B1(n9539), .B2(n9548), .ZN(
        P1_U3478) );
  OAI22_X1 U10640 ( .A1(n9543), .A2(n9542), .B1(n9541), .B2(n9540), .ZN(n9545)
         );
  AOI211_X1 U10641 ( .C1(n9547), .C2(n9546), .A(n9545), .B(n9544), .ZN(n9561)
         );
  INV_X1 U10642 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9549) );
  AOI22_X1 U10643 ( .A1(n9550), .A2(n9561), .B1(n9549), .B2(n9548), .ZN(
        P1_U3481) );
  AOI22_X1 U10644 ( .A1(n9562), .A2(n9551), .B1(n6267), .B2(n9559), .ZN(
        P1_U3525) );
  INV_X1 U10645 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9552) );
  AOI22_X1 U10646 ( .A1(n9562), .A2(n9553), .B1(n9552), .B2(n9559), .ZN(
        P1_U3527) );
  INV_X1 U10647 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9554) );
  AOI22_X1 U10648 ( .A1(n9562), .A2(n9555), .B1(n9554), .B2(n9559), .ZN(
        P1_U3528) );
  AOI22_X1 U10649 ( .A1(n9562), .A2(n9556), .B1(n9862), .B2(n9559), .ZN(
        P1_U3529) );
  INV_X1 U10650 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9557) );
  AOI22_X1 U10651 ( .A1(n9562), .A2(n9558), .B1(n9557), .B2(n9559), .ZN(
        P1_U3531) );
  INV_X1 U10652 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9560) );
  AOI22_X1 U10653 ( .A1(n9562), .A2(n9561), .B1(n9560), .B2(n9559), .ZN(
        P1_U3532) );
  INV_X1 U10654 ( .A(n9563), .ZN(n9564) );
  NOR2_X1 U10655 ( .A1(n9565), .A2(n9564), .ZN(n9566) );
  XNOR2_X1 U10656 ( .A(n9566), .B(n9567), .ZN(n9574) );
  NAND2_X1 U10657 ( .A1(n9568), .A2(n9567), .ZN(n9569) );
  NAND2_X1 U10658 ( .A1(n9570), .A2(n9569), .ZN(n9680) );
  NOR2_X1 U10659 ( .A1(n9680), .A2(n9571), .ZN(n9572) );
  AOI211_X1 U10660 ( .C1(n8492), .C2(n9574), .A(n9573), .B(n9572), .ZN(n9679)
         );
  AOI222_X1 U10661 ( .A1(n9676), .A2(n9577), .B1(P2_REG2_REG_10__SCAN_IN), 
        .B2(n9588), .C1(n9576), .C2(n9575), .ZN(n9587) );
  OAI21_X1 U10662 ( .B1(n9579), .B2(n9578), .A(n9650), .ZN(n9581) );
  NOR2_X1 U10663 ( .A1(n9581), .A2(n9580), .ZN(n9675) );
  INV_X1 U10664 ( .A(n9675), .ZN(n9582) );
  OAI22_X1 U10665 ( .A1(n9680), .A2(n9584), .B1(n9583), .B2(n9582), .ZN(n9585)
         );
  INV_X1 U10666 ( .A(n9585), .ZN(n9586) );
  OAI211_X1 U10667 ( .C1(n9588), .C2(n9679), .A(n9587), .B(n9586), .ZN(
        P2_U3286) );
  NOR2_X1 U10668 ( .A1(n9590), .A2(n9589), .ZN(n9604) );
  INV_X1 U10669 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9591) );
  NOR2_X1 U10670 ( .A1(n9625), .A2(n9591), .ZN(P2_U3297) );
  INV_X1 U10671 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9592) );
  NOR2_X1 U10672 ( .A1(n9625), .A2(n9592), .ZN(P2_U3298) );
  INV_X1 U10673 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9593) );
  NOR2_X1 U10674 ( .A1(n9625), .A2(n9593), .ZN(P2_U3299) );
  INV_X1 U10675 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n9594) );
  NOR2_X1 U10676 ( .A1(n9625), .A2(n9594), .ZN(P2_U3300) );
  INV_X1 U10677 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n9595) );
  NOR2_X1 U10678 ( .A1(n9604), .A2(n9595), .ZN(P2_U3301) );
  INV_X1 U10679 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9596) );
  NOR2_X1 U10680 ( .A1(n9604), .A2(n9596), .ZN(P2_U3302) );
  INV_X1 U10681 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9597) );
  NOR2_X1 U10682 ( .A1(n9604), .A2(n9597), .ZN(P2_U3303) );
  INV_X1 U10683 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n9598) );
  NOR2_X1 U10684 ( .A1(n9604), .A2(n9598), .ZN(P2_U3304) );
  NOR2_X1 U10685 ( .A1(n9604), .A2(n9839), .ZN(P2_U3305) );
  INV_X1 U10686 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n9599) );
  NOR2_X1 U10687 ( .A1(n9604), .A2(n9599), .ZN(P2_U3306) );
  INV_X1 U10688 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n9600) );
  NOR2_X1 U10689 ( .A1(n9604), .A2(n9600), .ZN(P2_U3307) );
  INV_X1 U10690 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n9601) );
  NOR2_X1 U10691 ( .A1(n9604), .A2(n9601), .ZN(P2_U3308) );
  INV_X1 U10692 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9602) );
  NOR2_X1 U10693 ( .A1(n9604), .A2(n9602), .ZN(P2_U3309) );
  INV_X1 U10694 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n9603) );
  NOR2_X1 U10695 ( .A1(n9604), .A2(n9603), .ZN(P2_U3310) );
  INV_X1 U10696 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9605) );
  NOR2_X1 U10697 ( .A1(n9625), .A2(n9605), .ZN(P2_U3311) );
  INV_X1 U10698 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9606) );
  NOR2_X1 U10699 ( .A1(n9625), .A2(n9606), .ZN(P2_U3312) );
  INV_X1 U10700 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n9607) );
  NOR2_X1 U10701 ( .A1(n9625), .A2(n9607), .ZN(P2_U3313) );
  INV_X1 U10702 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n9608) );
  NOR2_X1 U10703 ( .A1(n9625), .A2(n9608), .ZN(P2_U3314) );
  INV_X1 U10704 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9609) );
  NOR2_X1 U10705 ( .A1(n9625), .A2(n9609), .ZN(P2_U3315) );
  INV_X1 U10706 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n9610) );
  NOR2_X1 U10707 ( .A1(n9625), .A2(n9610), .ZN(P2_U3316) );
  INV_X1 U10708 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n9611) );
  NOR2_X1 U10709 ( .A1(n9625), .A2(n9611), .ZN(P2_U3317) );
  INV_X1 U10710 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9612) );
  NOR2_X1 U10711 ( .A1(n9625), .A2(n9612), .ZN(P2_U3318) );
  INV_X1 U10712 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9613) );
  NOR2_X1 U10713 ( .A1(n9625), .A2(n9613), .ZN(P2_U3319) );
  INV_X1 U10714 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9614) );
  NOR2_X1 U10715 ( .A1(n9625), .A2(n9614), .ZN(P2_U3320) );
  INV_X1 U10716 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n9615) );
  NOR2_X1 U10717 ( .A1(n9625), .A2(n9615), .ZN(P2_U3321) );
  INV_X1 U10718 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n9616) );
  NOR2_X1 U10719 ( .A1(n9625), .A2(n9616), .ZN(P2_U3322) );
  INV_X1 U10720 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n9617) );
  NOR2_X1 U10721 ( .A1(n9625), .A2(n9617), .ZN(P2_U3323) );
  NOR2_X1 U10722 ( .A1(n9625), .A2(n9618), .ZN(P2_U3324) );
  NOR2_X1 U10723 ( .A1(n9625), .A2(n9619), .ZN(P2_U3325) );
  NOR2_X1 U10724 ( .A1(n9625), .A2(n9620), .ZN(P2_U3326) );
  OAI22_X1 U10725 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9625), .B1(n9624), .B2(
        n9621), .ZN(n9622) );
  INV_X1 U10726 ( .A(n9622), .ZN(P2_U3437) );
  OAI22_X1 U10727 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n9625), .B1(n9624), .B2(
        n9623), .ZN(n9626) );
  INV_X1 U10728 ( .A(n9626), .ZN(P2_U3438) );
  AOI22_X1 U10729 ( .A1(n9629), .A2(n9697), .B1(n9628), .B2(n9627), .ZN(n9630)
         );
  AND2_X1 U10730 ( .A1(n9631), .A2(n9630), .ZN(n9701) );
  INV_X1 U10731 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9632) );
  AOI22_X1 U10732 ( .A1(n9700), .A2(n9701), .B1(n9632), .B2(n9698), .ZN(
        P2_U3451) );
  INV_X1 U10733 ( .A(n9633), .ZN(n9638) );
  OAI211_X1 U10734 ( .C1(n9636), .C2(n9690), .A(n9635), .B(n9634), .ZN(n9637)
         );
  AOI21_X1 U10735 ( .B1(n9638), .B2(n9697), .A(n9637), .ZN(n9703) );
  INV_X1 U10736 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9639) );
  AOI22_X1 U10737 ( .A1(n9700), .A2(n9703), .B1(n9639), .B2(n9698), .ZN(
        P2_U3457) );
  OAI22_X1 U10738 ( .A1(n9641), .A2(n9692), .B1(n9640), .B2(n9690), .ZN(n9643)
         );
  AOI211_X1 U10739 ( .C1(n9697), .C2(n9644), .A(n9643), .B(n9642), .ZN(n9705)
         );
  INV_X1 U10740 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9645) );
  AOI22_X1 U10741 ( .A1(n9700), .A2(n9705), .B1(n9645), .B2(n9698), .ZN(
        P2_U3463) );
  NAND3_X1 U10742 ( .A1(n9647), .A2(n9646), .A3(n9697), .ZN(n9654) );
  INV_X1 U10743 ( .A(n9648), .ZN(n9651) );
  AOI22_X1 U10744 ( .A1(n9651), .A2(n9650), .B1(n9677), .B2(n9649), .ZN(n9652)
         );
  AND3_X1 U10745 ( .A1(n9654), .A2(n9653), .A3(n9652), .ZN(n9706) );
  INV_X1 U10746 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9655) );
  AOI22_X1 U10747 ( .A1(n9700), .A2(n9706), .B1(n9655), .B2(n9698), .ZN(
        P2_U3469) );
  OAI21_X1 U10748 ( .B1(n9657), .B2(n9690), .A(n9656), .ZN(n9659) );
  AOI211_X1 U10749 ( .C1(n9697), .C2(n9660), .A(n9659), .B(n9658), .ZN(n9708)
         );
  INV_X1 U10750 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9661) );
  AOI22_X1 U10751 ( .A1(n9700), .A2(n9708), .B1(n9661), .B2(n9698), .ZN(
        P2_U3472) );
  INV_X1 U10752 ( .A(n9681), .ZN(n9673) );
  OAI22_X1 U10753 ( .A1(n9663), .A2(n9692), .B1(n9662), .B2(n9690), .ZN(n9665)
         );
  AOI211_X1 U10754 ( .C1(n9673), .C2(n9666), .A(n9665), .B(n9664), .ZN(n9709)
         );
  INV_X1 U10755 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9667) );
  AOI22_X1 U10756 ( .A1(n9700), .A2(n9709), .B1(n9667), .B2(n9698), .ZN(
        P2_U3475) );
  OAI22_X1 U10757 ( .A1(n9669), .A2(n9692), .B1(n9668), .B2(n9690), .ZN(n9671)
         );
  AOI211_X1 U10758 ( .C1(n9673), .C2(n9672), .A(n9671), .B(n9670), .ZN(n9710)
         );
  INV_X1 U10759 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9674) );
  AOI22_X1 U10760 ( .A1(n9700), .A2(n9710), .B1(n9674), .B2(n9698), .ZN(
        P2_U3478) );
  AOI21_X1 U10761 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9678) );
  OAI211_X1 U10762 ( .C1(n9681), .C2(n9680), .A(n9679), .B(n9678), .ZN(n9682)
         );
  INV_X1 U10763 ( .A(n9682), .ZN(n9711) );
  INV_X1 U10764 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9813) );
  AOI22_X1 U10765 ( .A1(n9700), .A2(n9711), .B1(n9813), .B2(n9698), .ZN(
        P2_U3481) );
  INV_X1 U10766 ( .A(n9683), .ZN(n9688) );
  OAI22_X1 U10767 ( .A1(n9685), .A2(n9692), .B1(n9684), .B2(n9690), .ZN(n9687)
         );
  AOI211_X1 U10768 ( .C1(n9688), .C2(n9697), .A(n9687), .B(n9686), .ZN(n9712)
         );
  INV_X1 U10769 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9689) );
  AOI22_X1 U10770 ( .A1(n9700), .A2(n9712), .B1(n9689), .B2(n9698), .ZN(
        P2_U3484) );
  OAI22_X1 U10771 ( .A1(n9693), .A2(n9692), .B1(n9691), .B2(n9690), .ZN(n9695)
         );
  AOI211_X1 U10772 ( .C1(n9697), .C2(n9696), .A(n9695), .B(n9694), .ZN(n9714)
         );
  INV_X1 U10773 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9699) );
  AOI22_X1 U10774 ( .A1(n9700), .A2(n9714), .B1(n9699), .B2(n9698), .ZN(
        P2_U3487) );
  AOI22_X1 U10775 ( .A1(n9715), .A2(n9701), .B1(n6389), .B2(n9713), .ZN(
        P2_U3520) );
  INV_X1 U10776 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9702) );
  AOI22_X1 U10777 ( .A1(n9715), .A2(n9703), .B1(n9702), .B2(n9713), .ZN(
        P2_U3522) );
  INV_X1 U10778 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9704) );
  AOI22_X1 U10779 ( .A1(n9715), .A2(n9705), .B1(n9704), .B2(n9713), .ZN(
        P2_U3524) );
  AOI22_X1 U10780 ( .A1(n9715), .A2(n9706), .B1(n7313), .B2(n9713), .ZN(
        P2_U3526) );
  INV_X1 U10781 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9707) );
  AOI22_X1 U10782 ( .A1(n9715), .A2(n9708), .B1(n9707), .B2(n9713), .ZN(
        P2_U3527) );
  AOI22_X1 U10783 ( .A1(n9715), .A2(n9709), .B1(n7315), .B2(n9713), .ZN(
        P2_U3528) );
  AOI22_X1 U10784 ( .A1(n9715), .A2(n9710), .B1(n7316), .B2(n9713), .ZN(
        P2_U3529) );
  AOI22_X1 U10785 ( .A1(n9715), .A2(n9711), .B1(n7317), .B2(n9713), .ZN(
        P2_U3530) );
  AOI22_X1 U10786 ( .A1(n9715), .A2(n9712), .B1(n7318), .B2(n9713), .ZN(
        P2_U3531) );
  AOI22_X1 U10787 ( .A1(n9715), .A2(n9714), .B1(n7319), .B2(n9713), .ZN(
        P2_U3532) );
  INV_X1 U10788 ( .A(n9716), .ZN(n9717) );
  NAND2_X1 U10789 ( .A1(n9718), .A2(n9717), .ZN(n9719) );
  XOR2_X1 U10790 ( .A(n9720), .B(n9719), .Z(ADD_1071_U5) );
  XOR2_X1 U10791 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10792 ( .B1(n9723), .B2(n9722), .A(n9721), .ZN(ADD_1071_U56) );
  OAI21_X1 U10793 ( .B1(n9726), .B2(n9725), .A(n9724), .ZN(ADD_1071_U57) );
  OAI21_X1 U10794 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(ADD_1071_U58) );
  OAI21_X1 U10795 ( .B1(n9732), .B2(n9731), .A(n9730), .ZN(ADD_1071_U59) );
  OAI21_X1 U10796 ( .B1(n9735), .B2(n9734), .A(n9733), .ZN(ADD_1071_U60) );
  OAI21_X1 U10797 ( .B1(n9738), .B2(n9737), .A(n9736), .ZN(ADD_1071_U61) );
  AOI21_X1 U10798 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(ADD_1071_U62) );
  AOI21_X1 U10799 ( .B1(n9744), .B2(n9743), .A(n9742), .ZN(ADD_1071_U63) );
  MUX2_X1 U10800 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9745), .S(P1_U4006), .Z(
        n9900) );
  INV_X1 U10801 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9746) );
  NOR4_X1 U10802 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), 
        .A3(P2_D_REG_0__SCAN_IN), .A4(n9746), .ZN(n9771) );
  NAND4_X1 U10803 ( .A1(P1_REG1_REG_24__SCAN_IN), .A2(P2_REG2_REG_1__SCAN_IN), 
        .A3(P2_REG0_REG_31__SCAN_IN), .A4(n9834), .ZN(n9749) );
  NAND3_X1 U10804 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_REG0_REG_11__SCAN_IN), 
        .A3(P1_REG0_REG_28__SCAN_IN), .ZN(n9748) );
  INV_X1 U10805 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9884) );
  INV_X1 U10806 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9883) );
  NAND4_X1 U10807 ( .A1(P1_REG1_REG_20__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9884), .A4(n9883), .ZN(n9747) );
  NOR4_X1 U10808 ( .A1(SI_30_), .A2(n9749), .A3(n9748), .A4(n9747), .ZN(n9770)
         );
  NAND4_X1 U10809 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(n9813), .A3(n9821), .A4(
        n9817), .ZN(n9756) );
  NAND4_X1 U10810 ( .A1(n9751), .A2(n9750), .A3(SI_27_), .A4(
        P1_REG1_REG_19__SCAN_IN), .ZN(n9755) );
  NAND4_X1 U10811 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(P2_REG0_REG_15__SCAN_IN), 
        .A3(n9805), .A4(n9802), .ZN(n9752) );
  NOR2_X1 U10812 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n9752), .ZN(n9753) );
  NAND4_X1 U10813 ( .A1(n9753), .A2(P2_REG0_REG_20__SCAN_IN), .A3(
        P2_REG2_REG_5__SCAN_IN), .A4(n9777), .ZN(n9754) );
  NOR3_X1 U10814 ( .A1(n9756), .A2(n9755), .A3(n9754), .ZN(n9769) );
  NAND4_X1 U10815 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG1_REG_27__SCAN_IN), 
        .A3(P2_REG2_REG_4__SCAN_IN), .A4(n9819), .ZN(n9767) );
  NAND4_X1 U10816 ( .A1(P1_REG2_REG_28__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .A3(P2_REG0_REG_16__SCAN_IN), .A4(n9855), .ZN(n9766) );
  NOR4_X1 U10817 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .A3(P1_IR_REG_29__SCAN_IN), .A4(P1_REG3_REG_5__SCAN_IN), .ZN(n9757) );
  INV_X1 U10818 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9799) );
  NAND4_X1 U10819 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n9758), .A3(n9757), .A4(
        n9799), .ZN(n9765) );
  INV_X1 U10820 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9773) );
  NOR4_X1 U10821 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), 
        .A3(n9773), .A4(n9775), .ZN(n9763) );
  NOR4_X1 U10822 ( .A1(P1_D_REG_0__SCAN_IN), .A2(P1_DATAO_REG_1__SCAN_IN), 
        .A3(n9759), .A4(n9786), .ZN(n9762) );
  INV_X1 U10823 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9790) );
  AND4_X1 U10824 ( .A1(n9789), .A2(n9790), .A3(P2_IR_REG_12__SCAN_IN), .A4(
        P2_DATAO_REG_22__SCAN_IN), .ZN(n9761) );
  INV_X1 U10825 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9871) );
  NOR4_X1 U10826 ( .A1(P2_REG2_REG_30__SCAN_IN), .A2(n9862), .A3(n9867), .A4(
        n9871), .ZN(n9760) );
  NAND4_X1 U10827 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(n9764)
         );
  NOR4_X1 U10828 ( .A1(n9767), .A2(n9766), .A3(n9765), .A4(n9764), .ZN(n9768)
         );
  NAND4_X1 U10829 ( .A1(n9771), .A2(n9770), .A3(n9769), .A4(n9768), .ZN(n9898)
         );
  AOI22_X1 U10830 ( .A1(n9773), .A2(keyinput22), .B1(keyinput3), .B2(n5053), 
        .ZN(n9772) );
  OAI221_X1 U10831 ( .B1(n9773), .B2(keyinput22), .C1(n5053), .C2(keyinput3), 
        .A(n9772), .ZN(n9784) );
  AOI22_X1 U10832 ( .A1(n7215), .A2(keyinput37), .B1(keyinput2), .B2(n9775), 
        .ZN(n9774) );
  OAI221_X1 U10833 ( .B1(n7215), .B2(keyinput37), .C1(n9775), .C2(keyinput2), 
        .A(n9774), .ZN(n9783) );
  AOI22_X1 U10834 ( .A1(n9778), .A2(keyinput61), .B1(keyinput55), .B2(n9777), 
        .ZN(n9776) );
  OAI221_X1 U10835 ( .B1(n9778), .B2(keyinput61), .C1(n9777), .C2(keyinput55), 
        .A(n9776), .ZN(n9782) );
  XNOR2_X1 U10836 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput8), .ZN(n9780) );
  XNOR2_X1 U10837 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput36), .ZN(n9779) );
  NAND2_X1 U10838 ( .A1(n9780), .A2(n9779), .ZN(n9781) );
  NOR4_X1 U10839 ( .A1(n9784), .A2(n9783), .A3(n9782), .A4(n9781), .ZN(n9831)
         );
  AOI22_X1 U10840 ( .A1(n9787), .A2(keyinput50), .B1(keyinput49), .B2(n9786), 
        .ZN(n9785) );
  OAI221_X1 U10841 ( .B1(n9787), .B2(keyinput50), .C1(n9786), .C2(keyinput49), 
        .A(n9785), .ZN(n9797) );
  AOI22_X1 U10842 ( .A1(n9790), .A2(keyinput41), .B1(keyinput23), .B2(n9789), 
        .ZN(n9788) );
  OAI221_X1 U10843 ( .B1(n9790), .B2(keyinput41), .C1(n9789), .C2(keyinput23), 
        .A(n9788), .ZN(n9796) );
  XNOR2_X1 U10844 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput32), .ZN(n9794)
         );
  XNOR2_X1 U10845 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput43), .ZN(n9793) );
  XNOR2_X1 U10846 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput42), .ZN(n9792) );
  XNOR2_X1 U10847 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(keyinput26), .ZN(n9791)
         );
  NAND4_X1 U10848 ( .A1(n9794), .A2(n9793), .A3(n9792), .A4(n9791), .ZN(n9795)
         );
  NOR3_X1 U10849 ( .A1(n9797), .A2(n9796), .A3(n9795), .ZN(n9830) );
  AOI22_X1 U10850 ( .A1(n9799), .A2(keyinput11), .B1(n6649), .B2(keyinput29), 
        .ZN(n9798) );
  OAI221_X1 U10851 ( .B1(n9799), .B2(keyinput11), .C1(n6649), .C2(keyinput29), 
        .A(n9798), .ZN(n9811) );
  AOI22_X1 U10852 ( .A1(n9802), .A2(keyinput1), .B1(n9801), .B2(keyinput52), 
        .ZN(n9800) );
  OAI221_X1 U10853 ( .B1(n9802), .B2(keyinput1), .C1(n9801), .C2(keyinput52), 
        .A(n9800), .ZN(n9810) );
  AOI22_X1 U10854 ( .A1(n9805), .A2(keyinput25), .B1(n9804), .B2(keyinput5), 
        .ZN(n9803) );
  OAI221_X1 U10855 ( .B1(n9805), .B2(keyinput25), .C1(n9804), .C2(keyinput5), 
        .A(n9803), .ZN(n9809) );
  XNOR2_X1 U10856 ( .A(P2_REG0_REG_20__SCAN_IN), .B(keyinput62), .ZN(n9807) );
  XNOR2_X1 U10857 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput48), .ZN(n9806) );
  NAND2_X1 U10858 ( .A1(n9807), .A2(n9806), .ZN(n9808) );
  NOR4_X1 U10859 ( .A1(n9811), .A2(n9810), .A3(n9809), .A4(n9808), .ZN(n9829)
         );
  INV_X1 U10860 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9814) );
  AOI22_X1 U10861 ( .A1(n9814), .A2(keyinput44), .B1(keyinput34), .B2(n9813), 
        .ZN(n9812) );
  OAI221_X1 U10862 ( .B1(n9814), .B2(keyinput44), .C1(n9813), .C2(keyinput34), 
        .A(n9812), .ZN(n9827) );
  INV_X1 U10863 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9816) );
  AOI22_X1 U10864 ( .A1(n9817), .A2(keyinput0), .B1(n9816), .B2(keyinput59), 
        .ZN(n9815) );
  OAI221_X1 U10865 ( .B1(n9817), .B2(keyinput0), .C1(n9816), .C2(keyinput59), 
        .A(n9815), .ZN(n9826) );
  INV_X1 U10866 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9820) );
  AOI22_X1 U10867 ( .A1(n9820), .A2(keyinput4), .B1(n9819), .B2(keyinput9), 
        .ZN(n9818) );
  OAI221_X1 U10868 ( .B1(n9820), .B2(keyinput4), .C1(n9819), .C2(keyinput9), 
        .A(n9818), .ZN(n9825) );
  XOR2_X1 U10869 ( .A(n9821), .B(keyinput10), .Z(n9823) );
  XNOR2_X1 U10870 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput24), .ZN(n9822) );
  NAND2_X1 U10871 ( .A1(n9823), .A2(n9822), .ZN(n9824) );
  NOR4_X1 U10872 ( .A1(n9827), .A2(n9826), .A3(n9825), .A4(n9824), .ZN(n9828)
         );
  NAND4_X1 U10873 ( .A1(n9831), .A2(n9830), .A3(n9829), .A4(n9828), .ZN(n9896)
         );
  INV_X1 U10874 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9833) );
  AOI22_X1 U10875 ( .A1(n9834), .A2(keyinput58), .B1(keyinput30), .B2(n9833), 
        .ZN(n9832) );
  OAI221_X1 U10876 ( .B1(n9834), .B2(keyinput58), .C1(n9833), .C2(keyinput30), 
        .A(n9832), .ZN(n9845) );
  AOI22_X1 U10877 ( .A1(n9836), .A2(keyinput7), .B1(keyinput28), .B2(n5461), 
        .ZN(n9835) );
  OAI221_X1 U10878 ( .B1(n9836), .B2(keyinput7), .C1(n5461), .C2(keyinput28), 
        .A(n9835), .ZN(n9844) );
  AOI22_X1 U10879 ( .A1(n9839), .A2(keyinput13), .B1(n9838), .B2(keyinput6), 
        .ZN(n9837) );
  OAI221_X1 U10880 ( .B1(n9839), .B2(keyinput13), .C1(n9838), .C2(keyinput6), 
        .A(n9837), .ZN(n9843) );
  XNOR2_X1 U10881 ( .A(P2_REG2_REG_1__SCAN_IN), .B(keyinput20), .ZN(n9841) );
  XNOR2_X1 U10882 ( .A(P1_REG1_REG_24__SCAN_IN), .B(keyinput16), .ZN(n9840) );
  NAND2_X1 U10883 ( .A1(n9841), .A2(n9840), .ZN(n9842) );
  NOR4_X1 U10884 ( .A1(n9845), .A2(n9844), .A3(n9843), .A4(n9842), .ZN(n9894)
         );
  INV_X1 U10885 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9848) );
  AOI22_X1 U10886 ( .A1(n9848), .A2(keyinput53), .B1(keyinput12), .B2(n9847), 
        .ZN(n9846) );
  OAI221_X1 U10887 ( .B1(n9848), .B2(keyinput53), .C1(n9847), .C2(keyinput12), 
        .A(n9846), .ZN(n9859) );
  INV_X1 U10888 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9851) );
  INV_X1 U10889 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9850) );
  AOI22_X1 U10890 ( .A1(n9851), .A2(keyinput46), .B1(n9850), .B2(keyinput38), 
        .ZN(n9849) );
  OAI221_X1 U10891 ( .B1(n9851), .B2(keyinput46), .C1(n9850), .C2(keyinput38), 
        .A(n9849), .ZN(n9858) );
  XNOR2_X1 U10892 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput51), .ZN(n9854) );
  XNOR2_X1 U10893 ( .A(P1_REG0_REG_14__SCAN_IN), .B(keyinput18), .ZN(n9853) );
  XNOR2_X1 U10894 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput54), .ZN(n9852) );
  NAND3_X1 U10895 ( .A1(n9854), .A2(n9853), .A3(n9852), .ZN(n9857) );
  XNOR2_X1 U10896 ( .A(n9855), .B(keyinput17), .ZN(n9856) );
  NOR4_X1 U10897 ( .A1(n9859), .A2(n9858), .A3(n9857), .A4(n9856), .ZN(n9893)
         );
  AOI22_X1 U10898 ( .A1(n9862), .A2(keyinput14), .B1(keyinput40), .B2(n9861), 
        .ZN(n9860) );
  OAI221_X1 U10899 ( .B1(n9862), .B2(keyinput14), .C1(n9861), .C2(keyinput40), 
        .A(n9860), .ZN(n9875) );
  INV_X1 U10900 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9865) );
  AOI22_X1 U10901 ( .A1(n9865), .A2(keyinput21), .B1(n9864), .B2(keyinput39), 
        .ZN(n9863) );
  OAI221_X1 U10902 ( .B1(n9865), .B2(keyinput21), .C1(n9864), .C2(keyinput39), 
        .A(n9863), .ZN(n9874) );
  INV_X1 U10903 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9868) );
  AOI22_X1 U10904 ( .A1(n9868), .A2(keyinput31), .B1(n9867), .B2(keyinput60), 
        .ZN(n9866) );
  OAI221_X1 U10905 ( .B1(n9868), .B2(keyinput31), .C1(n9867), .C2(keyinput60), 
        .A(n9866), .ZN(n9873) );
  AOI22_X1 U10906 ( .A1(n9871), .A2(keyinput27), .B1(n9870), .B2(keyinput19), 
        .ZN(n9869) );
  OAI221_X1 U10907 ( .B1(n9871), .B2(keyinput27), .C1(n9870), .C2(keyinput19), 
        .A(n9869), .ZN(n9872) );
  NOR4_X1 U10908 ( .A1(n9875), .A2(n9874), .A3(n9873), .A4(n9872), .ZN(n9892)
         );
  INV_X1 U10909 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9877) );
  AOI22_X1 U10910 ( .A1(n9878), .A2(keyinput15), .B1(keyinput35), .B2(n9877), 
        .ZN(n9876) );
  OAI221_X1 U10911 ( .B1(n9878), .B2(keyinput15), .C1(n9877), .C2(keyinput35), 
        .A(n9876), .ZN(n9890) );
  INV_X1 U10912 ( .A(SI_30_), .ZN(n9881) );
  AOI22_X1 U10913 ( .A1(n9881), .A2(keyinput33), .B1(n9880), .B2(keyinput57), 
        .ZN(n9879) );
  OAI221_X1 U10914 ( .B1(n9881), .B2(keyinput33), .C1(n9880), .C2(keyinput57), 
        .A(n9879), .ZN(n9889) );
  AOI22_X1 U10915 ( .A1(n9884), .A2(keyinput45), .B1(keyinput56), .B2(n9883), 
        .ZN(n9882) );
  OAI221_X1 U10916 ( .B1(n9884), .B2(keyinput45), .C1(n9883), .C2(keyinput56), 
        .A(n9882), .ZN(n9888) );
  XNOR2_X1 U10917 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput47), .ZN(n9886) );
  XNOR2_X1 U10918 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput63), .ZN(n9885) );
  NAND2_X1 U10919 ( .A1(n9886), .A2(n9885), .ZN(n9887) );
  NOR4_X1 U10920 ( .A1(n9890), .A2(n9889), .A3(n9888), .A4(n9887), .ZN(n9891)
         );
  NAND4_X1 U10921 ( .A1(n9894), .A2(n9893), .A3(n9892), .A4(n9891), .ZN(n9895)
         );
  NOR2_X1 U10922 ( .A1(n9896), .A2(n9895), .ZN(n9897) );
  XOR2_X1 U10923 ( .A(n9898), .B(n9897), .Z(n9899) );
  XNOR2_X1 U10924 ( .A(n9900), .B(n9899), .ZN(P1_U3573) );
  XOR2_X1 U10925 ( .A(n9901), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U10926 ( .A(n9902), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U10927 ( .A1(n9904), .A2(n9903), .ZN(n9905) );
  XOR2_X1 U10928 ( .A(n9905), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  OAI21_X1 U10929 ( .B1(n9908), .B2(n9907), .A(n9906), .ZN(n9909) );
  XNOR2_X1 U10930 ( .A(n9909), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U10931 ( .B1(n9912), .B2(n9911), .A(n9910), .ZN(ADD_1071_U47) );
  XOR2_X1 U10932 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9913), .Z(ADD_1071_U48) );
  XOR2_X1 U10933 ( .A(n9915), .B(n9914), .Z(ADD_1071_U54) );
  XOR2_X1 U10934 ( .A(n9917), .B(n9916), .Z(ADD_1071_U53) );
  XNOR2_X1 U10935 ( .A(n9919), .B(n9918), .ZN(ADD_1071_U52) );
  OAI211_X1 U4800 ( .C1(n5736), .C2(n6215), .A(n5637), .B(n5636), .ZN(n6163)
         );
  CLKBUF_X1 U4765 ( .A(n5574), .Z(n6018) );
  CLKBUF_X1 U4766 ( .A(n4265), .Z(n6244) );
  INV_X1 U6119 ( .A(n6051), .ZN(n5947) );
  INV_X1 U6901 ( .A(n4911), .ZN(n6196) );
endmodule

