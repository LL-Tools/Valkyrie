

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348;

  CLKBUF_X2 U2541 ( .A(n2931), .Z(n3044) );
  CLKBUF_X2 U2542 ( .A(n2917), .Z(n3704) );
  NAND2_X1 U2543 ( .A1(n2870), .A2(n2869), .ZN(n2800) );
  OR2_X1 U2544 ( .A1(n4630), .A2(n4370), .ZN(n2609) );
  NAND2_X1 U2545 ( .A1(n3553), .A2(n4348), .ZN(n3593) );
  NAND2_X1 U2546 ( .A1(n2601), .A2(n4350), .ZN(n3518) );
  CLKBUF_X2 U2547 ( .A(n2800), .Z(n3300) );
  AOI21_X2 U2548 ( .B1(n4431), .B2(n4810), .A(n3661), .ZN(n4791) );
  OAI21_X2 U2549 ( .B1(n3518), .B2(n3517), .A(n4328), .ZN(n3553) );
  INV_X4 U2550 ( .A(n3004), .ZN(n3726) );
  AND2_X4 U2551 ( .A1(n3288), .A2(n2909), .ZN(n3004) );
  OR2_X1 U2552 ( .A1(n4309), .A2(n4306), .ZN(n3240) );
  NOR2_X1 U2554 ( .A1(n2521), .A2(n4410), .ZN(n3702) );
  OR2_X1 U2555 ( .A1(n4737), .A2(n4366), .ZN(n2610) );
  NAND2_X1 U2556 ( .A1(n3789), .A2(n3788), .ZN(n3787) );
  AND2_X1 U2557 ( .A1(n3395), .A2(n2944), .ZN(n3470) );
  OAI21_X1 U2558 ( .B1(n3269), .B2(n5327), .A(n5300), .ZN(n5267) );
  INV_X1 U2559 ( .A(n3523), .ZN(n3524) );
  AND2_X2 U2560 ( .A1(n3434), .A2(n5300), .ZN(n5348) );
  AND2_X1 U2561 ( .A1(n2936), .A2(n2525), .ZN(n3488) );
  AND4_X1 U2562 ( .A1(n2949), .A2(n2948), .A3(n2947), .A4(n2946), .ZN(n3482)
         );
  NAND3_X1 U2563 ( .A1(n4913), .A2(n4911), .A3(n4912), .ZN(n3288) );
  NAND2_X1 U2564 ( .A1(n2913), .A2(n2912), .ZN(n3727) );
  AND2_X1 U2565 ( .A1(n4909), .A2(n4910), .ZN(n2945) );
  BUF_X2 U2566 ( .A(n2932), .Z(n3040) );
  NAND2_X1 U2567 ( .A1(n2722), .A2(n2784), .ZN(n2869) );
  XNOR2_X1 U2568 ( .A(n2718), .B(n4174), .ZN(n2865) );
  NAND2_X1 U2569 ( .A1(n2876), .A2(n4179), .ZN(n2878) );
  NAND2_X1 U2570 ( .A1(n2863), .A2(IR_REG_31__SCAN_IN), .ZN(n2718) );
  XNOR2_X1 U2571 ( .A(n2853), .B(IR_REG_22__SCAN_IN), .ZN(n4914) );
  OR2_X1 U2572 ( .A1(n2785), .A2(n2841), .ZN(n2876) );
  AND3_X1 U2573 ( .A1(n2685), .A2(n2684), .A3(n2626), .ZN(n2785) );
  AND2_X1 U2574 ( .A1(n2760), .A2(n2627), .ZN(n2626) );
  AND2_X1 U2575 ( .A1(n2686), .A2(n4160), .ZN(n2624) );
  AND2_X1 U2576 ( .A1(n2526), .A2(n2778), .ZN(n2627) );
  AND3_X1 U2577 ( .A1(n2789), .A2(n2771), .A3(n2770), .ZN(n2772) );
  INV_X1 U2578 ( .A(IR_REG_8__SCAN_IN), .ZN(n4141) );
  OAI21_X2 U2579 ( .B1(n4399), .B2(n3419), .A(n4343), .ZN(n3479) );
  NOR2_X2 U2580 ( .A1(n4773), .A2(n4364), .ZN(n4741) );
  AOI21_X2 U2581 ( .B1(n5278), .B2(n4439), .A(n4438), .ZN(n4648) );
  NOR2_X1 U2582 ( .A1(n4599), .A2(n2669), .ZN(n2668) );
  INV_X1 U2583 ( .A(n2673), .ZN(n2669) );
  INV_X1 U2584 ( .A(n2642), .ZN(n2639) );
  AND2_X1 U2585 ( .A1(n3288), .A2(n2913), .ZN(n2959) );
  NAND2_X1 U2586 ( .A1(n2559), .A2(n3306), .ZN(n3307) );
  OAI21_X1 U2587 ( .B1(n3344), .B2(n2691), .A(n2690), .ZN(n2689) );
  NAND2_X1 U2588 ( .A1(n2583), .A2(n4929), .ZN(n2690) );
  AND2_X1 U2589 ( .A1(n2605), .A2(n4383), .ZN(n2603) );
  NAND2_X1 U2590 ( .A1(n2932), .A2(REG1_REG_1__SCAN_IN), .ZN(n2907) );
  AND2_X1 U2591 ( .A1(n2885), .A2(n4911), .ZN(n2900) );
  INV_X1 U2592 ( .A(IR_REG_23__SCAN_IN), .ZN(n3965) );
  OR2_X1 U2593 ( .A1(n3042), .A2(n3041), .ZN(n3055) );
  AOI21_X1 U2594 ( .B1(n2748), .B2(n2753), .A(n2546), .ZN(n2747) );
  NAND2_X1 U2595 ( .A1(n2697), .A2(n2506), .ZN(n4967) );
  AND2_X1 U2596 ( .A1(n4967), .A2(n3304), .ZN(n4987) );
  NAND2_X1 U2597 ( .A1(n2586), .A2(REG2_REG_1__SCAN_IN), .ZN(n3304) );
  XNOR2_X1 U2598 ( .A(n2583), .B(n4929), .ZN(n3344) );
  OR2_X1 U2599 ( .A1(n4556), .A2(n2713), .ZN(n2711) );
  NAND2_X1 U2600 ( .A1(n2715), .A2(n2714), .ZN(n2713) );
  INV_X1 U2601 ( .A(n4557), .ZN(n2714) );
  NAND2_X1 U2602 ( .A1(n2674), .A2(n2527), .ZN(n2673) );
  NAND2_X1 U2603 ( .A1(n2646), .A2(n2644), .ZN(n3611) );
  INV_X1 U2604 ( .A(n2645), .ZN(n2644) );
  OAI21_X1 U2605 ( .B1(n2650), .B2(n2649), .A(n3602), .ZN(n2645) );
  NOR2_X1 U2606 ( .A1(n3564), .A2(n2655), .ZN(n2652) );
  CLKBUF_X1 U2607 ( .A(IR_REG_0__SCAN_IN), .Z(n4958) );
  INV_X1 U2608 ( .A(n4826), .ZN(n2637) );
  INV_X1 U2609 ( .A(IR_REG_17__SCAN_IN), .ZN(n4159) );
  INV_X1 U2610 ( .A(IR_REG_16__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U2611 ( .A1(n2995), .A2(n2996), .ZN(n2745) );
  AOI21_X1 U2612 ( .B1(n2522), .B2(n2982), .A(n2744), .ZN(n2743) );
  INV_X1 U2613 ( .A(n3727), .ZN(n3250) );
  INV_X1 U2614 ( .A(n2668), .ZN(n2667) );
  NAND2_X1 U2615 ( .A1(n2671), .A2(n2540), .ZN(n2660) );
  NOR2_X1 U2616 ( .A1(n2667), .A2(n2663), .ZN(n2662) );
  INV_X1 U2617 ( .A(n2671), .ZN(n2663) );
  INV_X1 U2618 ( .A(n2665), .ZN(n2658) );
  AOI21_X1 U2619 ( .B1(n2668), .B2(n2666), .A(n2532), .ZN(n2665) );
  INV_X1 U2620 ( .A(n2520), .ZN(n2666) );
  INV_X1 U2621 ( .A(n4446), .ZN(n2608) );
  NAND2_X1 U2622 ( .A1(n4604), .A2(n4621), .ZN(n2674) );
  NOR2_X1 U2623 ( .A1(n4408), .A2(n2672), .ZN(n2671) );
  NOR2_X1 U2624 ( .A1(n2540), .A2(n3655), .ZN(n2672) );
  NOR2_X1 U2625 ( .A1(n2617), .A2(n2615), .ZN(n2614) );
  AND2_X1 U2626 ( .A1(n2616), .A2(n4321), .ZN(n2615) );
  INV_X1 U2627 ( .A(n4339), .ZN(n2617) );
  INV_X1 U2628 ( .A(n4332), .ZN(n2616) );
  INV_X1 U2629 ( .A(n4324), .ZN(n2613) );
  AND2_X1 U2630 ( .A1(n5160), .A2(n4832), .ZN(n2631) );
  AOI21_X1 U2631 ( .B1(n4826), .B2(n2643), .A(n2544), .ZN(n2642) );
  INV_X1 U2632 ( .A(n3628), .ZN(n2643) );
  OAI22_X1 U2633 ( .A1(n4393), .A2(n2678), .B1(n3626), .B2(n5108), .ZN(n2677)
         );
  NAND2_X1 U2634 ( .A1(n2679), .A2(n4419), .ZN(n2678) );
  INV_X1 U2635 ( .A(n4418), .ZN(n2679) );
  NAND2_X1 U2636 ( .A1(n2900), .A2(n2896), .ZN(n3260) );
  AND2_X1 U2637 ( .A1(n4345), .A2(n5050), .ZN(n3478) );
  NAND2_X1 U2638 ( .A1(n5018), .A2(n3804), .ZN(n4343) );
  NOR2_X1 U2639 ( .A1(n4914), .A2(n4915), .ZN(n5014) );
  NAND2_X1 U2640 ( .A1(n4172), .A2(IR_REG_31__SCAN_IN), .ZN(n2860) );
  INV_X1 U2641 ( .A(IR_REG_22__SCAN_IN), .ZN(n4164) );
  NAND2_X1 U2642 ( .A1(n2848), .A2(n2777), .ZN(n2857) );
  INV_X1 U2643 ( .A(IR_REG_11__SCAN_IN), .ZN(n4146) );
  INV_X1 U2644 ( .A(IR_REG_7__SCAN_IN), .ZN(n4140) );
  AOI21_X1 U2645 ( .B1(n3418), .B2(n3004), .A(n2767), .ZN(n2926) );
  NAND2_X1 U2646 ( .A1(n3212), .A2(n2731), .ZN(n2730) );
  INV_X1 U2647 ( .A(n3210), .ZN(n2731) );
  INV_X1 U2648 ( .A(n4255), .ZN(n2732) );
  NOR2_X1 U2649 ( .A1(n2733), .A2(n2726), .ZN(n2725) );
  NOR2_X1 U2650 ( .A1(n3212), .A2(n4255), .ZN(n2733) );
  INV_X1 U2651 ( .A(n3198), .ZN(n2726) );
  NAND2_X1 U2652 ( .A1(n3764), .A2(n3198), .ZN(n3767) );
  XNOR2_X1 U2653 ( .A(n2962), .B(n3727), .ZN(n2963) );
  NAND2_X1 U2654 ( .A1(n2961), .A2(n2960), .ZN(n2962) );
  OR2_X1 U2655 ( .A1(n3493), .A2(n3725), .ZN(n2960) );
  NAND2_X1 U2656 ( .A1(n2923), .A2(n2766), .ZN(n3371) );
  NAND2_X1 U2657 ( .A1(n3418), .A2(n3253), .ZN(n2923) );
  NOR2_X1 U2658 ( .A1(n3055), .A2(n3586), .ZN(n3070) );
  NAND2_X1 U2659 ( .A1(n3775), .A2(n3035), .ZN(n3777) );
  NAND2_X1 U2660 ( .A1(n5222), .A2(n5221), .ZN(n5223) );
  AND2_X1 U2661 ( .A1(n3100), .A2(n3099), .ZN(n5190) );
  AND4_X1 U2662 ( .A1(n3048), .A2(n3047), .A3(n3046), .A4(n3045), .ZN(n3809)
         );
  NAND2_X1 U2663 ( .A1(n2557), .A2(n2558), .ZN(n2559) );
  INV_X1 U2664 ( .A(n4987), .ZN(n2558) );
  NAND2_X1 U2665 ( .A1(n2696), .A2(REG2_REG_3__SCAN_IN), .ZN(n2695) );
  NAND2_X1 U2666 ( .A1(n2707), .A2(REG2_REG_4__SCAN_IN), .ZN(n2706) );
  NAND2_X1 U2667 ( .A1(n3311), .A2(n2707), .ZN(n2705) );
  INV_X1 U2668 ( .A(n3365), .ZN(n2707) );
  XNOR2_X1 U2669 ( .A(n2689), .B(n3308), .ZN(n5008) );
  NAND2_X1 U2670 ( .A1(n2592), .A2(n2589), .ZN(n3359) );
  NAND2_X1 U2671 ( .A1(n2591), .A2(n2590), .ZN(n2589) );
  NAND2_X1 U2672 ( .A1(n5008), .A2(n2593), .ZN(n2592) );
  INV_X1 U2673 ( .A(n3360), .ZN(n2590) );
  NOR2_X1 U2674 ( .A1(n3359), .A2(n2595), .ZN(n3322) );
  AND2_X1 U2675 ( .A1(n4928), .A2(REG1_REG_5__SCAN_IN), .ZN(n2595) );
  NAND2_X1 U2676 ( .A1(n2563), .A2(REG2_REG_6__SCAN_IN), .ZN(n2709) );
  AND2_X1 U2677 ( .A1(n4926), .A2(REG2_REG_7__SCAN_IN), .ZN(n3316) );
  INV_X1 U2678 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3586) );
  NOR2_X1 U2679 ( .A1(n3581), .A2(n2708), .ZN(n4495) );
  XNOR2_X1 U2680 ( .A(n4487), .B(n4494), .ZN(n3585) );
  NAND2_X1 U2681 ( .A1(n3583), .A2(n3584), .ZN(n4487) );
  NAND2_X1 U2682 ( .A1(n3585), .A2(REG1_REG_12__SCAN_IN), .ZN(n4488) );
  OR2_X1 U2683 ( .A1(n4509), .A2(n2702), .ZN(n2701) );
  NAND2_X1 U2684 ( .A1(n2704), .A2(REG2_REG_14__SCAN_IN), .ZN(n2702) );
  NAND2_X1 U2685 ( .A1(n4524), .A2(n2704), .ZN(n2703) );
  NAND2_X1 U2686 ( .A1(n4532), .A2(n4531), .ZN(n4539) );
  XNOR2_X1 U2687 ( .A(n4553), .B(n4918), .ZN(n4544) );
  AND3_X1 U2688 ( .A1(n2701), .A2(n4525), .A3(n2703), .ZN(n4553) );
  NAND2_X1 U2689 ( .A1(n4544), .A2(n4543), .ZN(n4555) );
  OR2_X1 U2690 ( .A1(n3712), .A2(n4378), .ZN(n5331) );
  NAND2_X1 U2691 ( .A1(n2521), .A2(n4410), .ZN(n3682) );
  INV_X1 U2692 ( .A(n3702), .ZN(n3683) );
  INV_X1 U2693 ( .A(n3734), .ZN(n3724) );
  OR2_X1 U2694 ( .A1(n4630), .A2(n2606), .ZN(n2604) );
  NAND2_X1 U2695 ( .A1(n2608), .A2(n2607), .ZN(n2606) );
  INV_X1 U2696 ( .A(n4370), .ZN(n2607) );
  NAND2_X1 U2697 ( .A1(n2608), .A2(n4444), .ZN(n2605) );
  AND2_X1 U2698 ( .A1(n4383), .A2(n4375), .ZN(n4599) );
  NAND2_X1 U2699 ( .A1(n2656), .A2(n2671), .ZN(n2664) );
  OR2_X1 U2700 ( .A1(n2540), .A2(n4645), .ZN(n2656) );
  OAI21_X1 U2701 ( .B1(n4648), .B2(n4442), .A(n4414), .ZN(n4630) );
  AND4_X1 U2702 ( .A1(n3232), .A2(n3231), .A3(n3230), .A4(n3229), .ZN(n4634)
         );
  NAND2_X1 U2703 ( .A1(n5279), .A2(n5280), .ZN(n5278) );
  INV_X1 U2704 ( .A(n4323), .ZN(n3661) );
  INV_X1 U2705 ( .A(n4846), .ZN(n4858) );
  INV_X1 U2706 ( .A(n2682), .ZN(n4855) );
  OAI21_X1 U2707 ( .B1(n5102), .B2(n2680), .A(n2676), .ZN(n2682) );
  NAND2_X1 U2708 ( .A1(n2681), .A2(n4419), .ZN(n2680) );
  INV_X1 U2709 ( .A(n2677), .ZN(n2676) );
  OAI21_X1 U2710 ( .B1(n3611), .B2(n3610), .A(n3609), .ZN(n5102) );
  AOI21_X1 U2711 ( .B1(n2652), .B2(n3514), .A(n2524), .ZN(n2650) );
  NAND2_X1 U2712 ( .A1(n4462), .A2(n3260), .ZN(n3430) );
  INV_X1 U2713 ( .A(n5327), .ZN(n5282) );
  INV_X1 U2714 ( .A(n5283), .ZN(n5107) );
  AND2_X1 U2715 ( .A1(n2898), .A2(n3295), .ZN(n2899) );
  INV_X1 U2716 ( .A(n5293), .ZN(n5233) );
  NAND2_X1 U2717 ( .A1(n2862), .A2(n2863), .ZN(n2864) );
  MUX2_X1 U2718 ( .A(IR_REG_31__SCAN_IN), .B(n2782), .S(IR_REG_28__SCAN_IN), 
        .Z(n2784) );
  INV_X1 U2719 ( .A(IR_REG_27__SCAN_IN), .ZN(n3978) );
  INV_X1 U2720 ( .A(IR_REG_26__SCAN_IN), .ZN(n4179) );
  NAND2_X1 U2721 ( .A1(n2779), .A2(n3965), .ZN(n2780) );
  NAND2_X1 U2722 ( .A1(n2880), .A2(n3965), .ZN(n2882) );
  NAND2_X1 U2723 ( .A1(n2857), .A2(n2849), .ZN(n4592) );
  OR2_X1 U2724 ( .A1(n2848), .A2(n2777), .ZN(n2849) );
  INV_X1 U2725 ( .A(IR_REG_15__SCAN_IN), .ZN(n2834) );
  AND3_X1 U2726 ( .A1(n2773), .A2(n2772), .A3(n2717), .ZN(n2824) );
  OR2_X1 U2727 ( .A1(n2819), .A2(IR_REG_6__SCAN_IN), .ZN(n2810) );
  NAND2_X1 U2728 ( .A1(n2734), .A2(n2737), .ZN(n5259) );
  AOI21_X1 U2729 ( .B1(n5245), .B2(n2738), .A(n2514), .ZN(n2737) );
  INV_X1 U2730 ( .A(n4607), .ZN(n4469) );
  INV_X1 U2731 ( .A(n4651), .ZN(n4616) );
  NAND2_X1 U2732 ( .A1(n2697), .A2(n2568), .ZN(n4970) );
  NAND2_X1 U2733 ( .A1(n4973), .A2(n2529), .ZN(n4972) );
  NOR2_X1 U2734 ( .A1(n3582), .A2(n4836), .ZN(n4497) );
  XNOR2_X1 U2735 ( .A(n4495), .B(n4494), .ZN(n3582) );
  OR2_X1 U2736 ( .A1(n4966), .A2(n4979), .ZN(n4550) );
  AND2_X1 U2737 ( .A1(n3303), .A2(n3318), .ZN(n4998) );
  NAND2_X1 U2738 ( .A1(n4589), .A2(n5010), .ZN(n2692) );
  XNOR2_X1 U2739 ( .A(n2599), .B(n2598), .ZN(n4589) );
  INV_X1 U2740 ( .A(n4588), .ZN(n2598) );
  NAND2_X1 U2741 ( .A1(n4587), .A2(n2600), .ZN(n2599) );
  NAND2_X1 U2742 ( .A1(n2711), .A2(n2710), .ZN(n2578) );
  AND2_X1 U2743 ( .A1(n2712), .A2(n2556), .ZN(n2710) );
  NAND2_X1 U2744 ( .A1(n2619), .A2(n5289), .ZN(n2623) );
  AND2_X1 U2745 ( .A1(n2796), .A2(n2797), .ZN(n4929) );
  INV_X1 U2746 ( .A(IR_REG_18__SCAN_IN), .ZN(n4160) );
  INV_X1 U2747 ( .A(IR_REG_2__SCAN_IN), .ZN(n2792) );
  AND2_X1 U2748 ( .A1(n2751), .A2(n2749), .ZN(n2748) );
  INV_X1 U2749 ( .A(n3112), .ZN(n2749) );
  AND2_X1 U2750 ( .A1(n3082), .A2(n2755), .ZN(n2754) );
  INV_X1 U2751 ( .A(n3752), .ZN(n2755) );
  NAND2_X1 U2752 ( .A1(n4992), .A2(n2584), .ZN(n2583) );
  NAND2_X1 U2753 ( .A1(n4989), .A2(REG1_REG_2__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U2754 ( .A1(n2695), .A2(n2530), .ZN(n3309) );
  NAND2_X1 U2755 ( .A1(n3309), .A2(n5002), .ZN(n3310) );
  NOR2_X1 U2756 ( .A1(n3360), .A2(n2594), .ZN(n2593) );
  INV_X1 U2757 ( .A(n2596), .ZN(n2591) );
  NAND2_X1 U2758 ( .A1(n3407), .A2(n3406), .ZN(n3408) );
  NAND2_X1 U2759 ( .A1(n3408), .A2(n4923), .ZN(n3453) );
  INV_X1 U2760 ( .A(n4500), .ZN(n2572) );
  INV_X1 U2761 ( .A(n4526), .ZN(n2704) );
  NAND2_X1 U2762 ( .A1(n4511), .A2(n4512), .ZN(n4527) );
  INV_X1 U2763 ( .A(n4572), .ZN(n2715) );
  NOR2_X1 U2764 ( .A1(n3227), .A2(n4310), .ZN(n3241) );
  NOR2_X1 U2765 ( .A1(n4632), .A2(n4257), .ZN(n2633) );
  NOR2_X1 U2766 ( .A1(n2630), .A2(n5281), .ZN(n2629) );
  INV_X1 U2767 ( .A(n4394), .ZN(n2649) );
  NOR2_X1 U2768 ( .A1(n2649), .A2(n2648), .ZN(n2647) );
  INV_X1 U2769 ( .A(n2652), .ZN(n2648) );
  INV_X1 U2770 ( .A(n3424), .ZN(n3298) );
  NAND2_X1 U2771 ( .A1(n3417), .A2(n3448), .ZN(n4341) );
  AOI21_X1 U2772 ( .B1(n2638), .B2(n2637), .A(n2545), .ZN(n2636) );
  OR2_X1 U2773 ( .A1(n4754), .A2(n4436), .ZN(n4782) );
  NOR2_X1 U2774 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2781)
         );
  INV_X1 U2775 ( .A(IR_REG_30__SCAN_IN), .ZN(n4174) );
  AND2_X1 U2776 ( .A1(n2775), .A2(n4159), .ZN(n2625) );
  AND2_X1 U2777 ( .A1(n2774), .A2(n2717), .ZN(n2686) );
  NOR2_X1 U2778 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2774)
         );
  INV_X1 U2779 ( .A(IR_REG_14__SCAN_IN), .ZN(n4147) );
  INV_X1 U2780 ( .A(IR_REG_10__SCAN_IN), .ZN(n2717) );
  NOR2_X1 U2781 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2771)
         );
  NOR2_X1 U2782 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2770)
         );
  AND3_X1 U2783 ( .A1(n2817), .A2(n4141), .A3(n2792), .ZN(n2773) );
  NAND2_X1 U2784 ( .A1(n3824), .A2(n2756), .ZN(n3723) );
  NOR2_X1 U2785 ( .A1(n3256), .A2(n2757), .ZN(n2756) );
  INV_X1 U2786 ( .A(n3226), .ZN(n2757) );
  NAND2_X1 U2787 ( .A1(n2742), .A2(n2740), .ZN(n3789) );
  NAND2_X1 U2788 ( .A1(n2741), .A2(n2745), .ZN(n2740) );
  OR2_X1 U2789 ( .A1(n3213), .A2(n3918), .ZN(n3227) );
  AND2_X1 U2790 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2967) );
  NOR2_X1 U2791 ( .A1(n2739), .A2(n2736), .ZN(n2735) );
  INV_X1 U2792 ( .A(n5221), .ZN(n2736) );
  INV_X1 U2793 ( .A(n5245), .ZN(n2739) );
  NAND2_X1 U2794 ( .A1(n4275), .A2(n4276), .ZN(n4274) );
  INV_X1 U2795 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3041) );
  OR2_X1 U2796 ( .A1(n3281), .A2(n3302), .ZN(n3269) );
  AOI21_X1 U2797 ( .B1(n2752), .B2(n2754), .A(n2553), .ZN(n2751) );
  INV_X1 U2798 ( .A(n4276), .ZN(n2752) );
  INV_X1 U2799 ( .A(n2754), .ZN(n2753) );
  AND4_X1 U2800 ( .A1(n3087), .A2(n3086), .A3(n3085), .A4(n3084), .ZN(n4792)
         );
  AND4_X1 U2801 ( .A1(n2991), .A2(n2990), .A3(n2989), .A4(n2988), .ZN(n3596)
         );
  XNOR2_X1 U2802 ( .A(n3307), .B(n4929), .ZN(n3347) );
  NOR2_X1 U2803 ( .A1(n5001), .A2(n5000), .ZN(n4999) );
  OR2_X1 U2804 ( .A1(n3389), .A2(n3388), .ZN(n3407) );
  OAI21_X1 U2805 ( .B1(n4923), .B2(n3408), .A(n3453), .ZN(n3409) );
  NOR2_X1 U2806 ( .A1(n3409), .A2(n3622), .ZN(n3455) );
  OAI21_X1 U2807 ( .B1(n3459), .B2(n3458), .A(n2688), .ZN(n3463) );
  NAND2_X1 U2808 ( .A1(n2597), .A2(n4923), .ZN(n2688) );
  NAND2_X1 U2809 ( .A1(n2571), .A2(n2569), .ZN(n4520) );
  AOI21_X1 U2810 ( .B1(n4496), .B2(n2572), .A(n2570), .ZN(n2569) );
  NAND2_X1 U2811 ( .A1(n4497), .A2(n2572), .ZN(n2571) );
  INV_X1 U2812 ( .A(n4508), .ZN(n2570) );
  XNOR2_X1 U2813 ( .A(n4527), .B(n4521), .ZN(n4513) );
  NOR2_X1 U2814 ( .A1(n4559), .A2(n4560), .ZN(n4563) );
  INV_X1 U2815 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4577) );
  AND2_X1 U2816 ( .A1(n4570), .A2(REG2_REG_17__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U2817 ( .A1(n4575), .A2(n4576), .ZN(n4587) );
  NAND2_X1 U2818 ( .A1(n4917), .A2(REG1_REG_18__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U2819 ( .A1(n2715), .A2(n2716), .ZN(n2712) );
  AND2_X1 U2820 ( .A1(n3300), .A2(DATAI_28_), .ZN(n3734) );
  NAND2_X1 U2821 ( .A1(n2661), .A2(n2657), .ZN(n3699) );
  NOR2_X1 U2822 ( .A1(n2659), .A2(n2658), .ZN(n2657) );
  NOR2_X1 U2823 ( .A1(n2667), .A2(n2660), .ZN(n2659) );
  AND2_X1 U2824 ( .A1(n4669), .A2(n2632), .ZN(n4594) );
  AND2_X1 U2825 ( .A1(n2516), .A2(n3657), .ZN(n2632) );
  NAND2_X1 U2826 ( .A1(n4669), .A2(n2516), .ZN(n4622) );
  AND2_X1 U2827 ( .A1(n3300), .A2(DATAI_25_), .ZN(n4632) );
  NAND2_X1 U2828 ( .A1(n4669), .A2(n2633), .ZN(n4637) );
  AND4_X1 U2829 ( .A1(n3218), .A2(n3217), .A3(n3216), .A4(n3215), .ZN(n4651)
         );
  NAND2_X1 U2830 ( .A1(n4669), .A2(n4656), .ZN(n4655) );
  AND2_X1 U2831 ( .A1(n4693), .A2(n4671), .ZN(n4669) );
  INV_X1 U2832 ( .A(n3769), .ZN(n4671) );
  AND2_X1 U2833 ( .A1(n4663), .A2(n3678), .ZN(n4686) );
  AND2_X1 U2834 ( .A1(n4748), .A2(n2628), .ZN(n4693) );
  AND2_X1 U2835 ( .A1(n2515), .A2(n4290), .ZN(n2628) );
  OAI21_X1 U2836 ( .B1(n4700), .B2(n3652), .A(n3653), .ZN(n4681) );
  OR2_X1 U2837 ( .A1(n4681), .A2(n4686), .ZN(n4682) );
  NAND2_X1 U2838 ( .A1(n4748), .A2(n2515), .ZN(n4712) );
  OR2_X1 U2839 ( .A1(n4416), .A2(n4415), .ZN(n4701) );
  NAND2_X1 U2840 ( .A1(REG3_REG_20__SCAN_IN), .A2(n3151), .ZN(n3178) );
  NAND2_X1 U2841 ( .A1(n2610), .A2(n3669), .ZN(n5279) );
  AND2_X1 U2842 ( .A1(n3671), .A2(n3670), .ZN(n5280) );
  NAND2_X1 U2843 ( .A1(n4748), .A2(n2629), .ZN(n5275) );
  AND2_X1 U2844 ( .A1(n4748), .A2(n4729), .ZN(n5277) );
  NOR2_X1 U2845 ( .A1(n4741), .A2(n3674), .ZN(n4737) );
  NOR2_X1 U2846 ( .A1(n2769), .A2(n5227), .ZN(n4748) );
  OR2_X1 U2847 ( .A1(n4781), .A2(n4761), .ZN(n2769) );
  NOR2_X1 U2848 ( .A1(n3101), .A2(n3840), .ZN(n3113) );
  AND4_X1 U2849 ( .A1(n3097), .A2(n3096), .A3(n3095), .A4(n3094), .ZN(n4774)
         );
  AND2_X1 U2850 ( .A1(n4771), .A2(n4770), .ZN(n4773) );
  AND2_X1 U2851 ( .A1(n4856), .A2(n2549), .ZN(n4804) );
  INV_X1 U2852 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4514) );
  NOR2_X1 U2853 ( .A1(n3083), .A2(n4514), .ZN(n3092) );
  AOI21_X1 U2854 ( .B1(n2614), .B2(n2618), .A(n2613), .ZN(n2612) );
  INV_X1 U2855 ( .A(n4321), .ZN(n2618) );
  AND2_X1 U2856 ( .A1(n4323), .A2(n4318), .ZN(n4810) );
  NAND2_X1 U2857 ( .A1(n4856), .A2(n2512), .ZN(n4817) );
  INV_X1 U2858 ( .A(n4810), .ZN(n4815) );
  NAND2_X1 U2859 ( .A1(n4827), .A2(n4321), .ZN(n5156) );
  NAND2_X1 U2860 ( .A1(n4856), .A2(n2631), .ZN(n5166) );
  NAND2_X1 U2861 ( .A1(n2640), .A2(n2642), .ZN(n5154) );
  NAND2_X1 U2862 ( .A1(n2641), .A2(n4826), .ZN(n2640) );
  NAND2_X1 U2863 ( .A1(n4843), .A2(n4332), .ZN(n4827) );
  NAND2_X1 U2864 ( .A1(n4856), .A2(n4832), .ZN(n5164) );
  AND2_X1 U2865 ( .A1(n4859), .A2(n4858), .ZN(n4856) );
  AND4_X1 U2866 ( .A1(n3059), .A2(n3058), .A3(n3057), .A4(n3056), .ZN(n4849)
         );
  AND2_X1 U2867 ( .A1(n4320), .A2(n4332), .ZN(n4844) );
  OAI21_X1 U2868 ( .B1(n5112), .B2(n5111), .A(n4358), .ZN(n3615) );
  NAND2_X1 U2869 ( .A1(n3615), .A2(n4393), .ZN(n3658) );
  AND2_X1 U2870 ( .A1(n2634), .A2(n3560), .ZN(n4859) );
  AND2_X1 U2871 ( .A1(n2511), .A2(n3626), .ZN(n2634) );
  NAND2_X1 U2872 ( .A1(n3560), .A2(n2511), .ZN(n5104) );
  AND2_X1 U2873 ( .A1(n2997), .A2(REG3_REG_8__SCAN_IN), .ZN(n3012) );
  AND2_X1 U2874 ( .A1(n3012), .A2(REG3_REG_9__SCAN_IN), .ZN(n3022) );
  AND4_X1 U2875 ( .A1(n3027), .A2(n3026), .A3(n3025), .A4(n3024), .ZN(n5108)
         );
  OAI21_X1 U2876 ( .B1(n3614), .B2(n4325), .A(n4355), .ZN(n5112) );
  NAND2_X1 U2877 ( .A1(n3560), .A2(n2510), .ZN(n5103) );
  AND2_X1 U2878 ( .A1(n3595), .A2(n3609), .ZN(n4421) );
  AND2_X1 U2879 ( .A1(n3560), .A2(n3554), .ZN(n3603) );
  NOR2_X1 U2880 ( .A1(n3523), .A2(n3573), .ZN(n3560) );
  AND4_X1 U2881 ( .A1(n2972), .A2(n2971), .A3(n2970), .A4(n2969), .ZN(n3504)
         );
  OR2_X1 U2882 ( .A1(n3525), .A2(n3545), .ZN(n3523) );
  NAND2_X1 U2883 ( .A1(n2602), .A2(n4397), .ZN(n3498) );
  NOR2_X1 U2884 ( .A1(n5047), .A2(n5048), .ZN(n5046) );
  NAND2_X1 U2885 ( .A1(n2917), .A2(REG2_REG_1__SCAN_IN), .ZN(n2906) );
  NAND2_X1 U2886 ( .A1(n4869), .A2(n4868), .ZN(n5293) );
  INV_X1 U2887 ( .A(n5291), .ZN(n5335) );
  NOR2_X1 U2888 ( .A1(n3430), .A2(n2897), .ZN(n2902) );
  INV_X1 U2889 ( .A(n2900), .ZN(n3292) );
  NOR2_X1 U2890 ( .A1(n2761), .A2(n2780), .ZN(n2760) );
  NAND2_X1 U2891 ( .A1(n2762), .A2(n4164), .ZN(n2761) );
  INV_X1 U2892 ( .A(IR_REG_25__SCAN_IN), .ZN(n2762) );
  NAND2_X1 U2893 ( .A1(n2882), .A2(n2881), .ZN(n3301) );
  XNOR2_X1 U2894 ( .A(n2858), .B(n2776), .ZN(n4866) );
  NAND2_X1 U2895 ( .A1(n2523), .A2(n2775), .ZN(n2759) );
  NAND2_X1 U2896 ( .A1(n2772), .A2(n2773), .ZN(n2821) );
  NAND2_X1 U2897 ( .A1(n2534), .A2(IR_REG_1__SCAN_IN), .ZN(n2564) );
  OAI21_X1 U2898 ( .B1(n2566), .B2(n2841), .A(n2700), .ZN(n2565) );
  OAI21_X1 U2899 ( .B1(n3572), .B2(n2522), .A(n2982), .ZN(n3742) );
  NAND2_X1 U2900 ( .A1(n4274), .A2(n3082), .ZN(n3754) );
  NAND2_X1 U2901 ( .A1(n2943), .A2(n2942), .ZN(n2944) );
  NAND2_X1 U2902 ( .A1(n5223), .A2(n5225), .ZN(n5244) );
  XOR2_X1 U2903 ( .A(n3730), .B(n3729), .Z(n3731) );
  AND4_X1 U2904 ( .A1(n3183), .A2(n3182), .A3(n3181), .A4(n3180), .ZN(n5316)
         );
  NAND2_X1 U2905 ( .A1(n3068), .A2(n3815), .ZN(n3819) );
  INV_X1 U2906 ( .A(n4829), .ZN(n4832) );
  INV_X1 U2907 ( .A(n5267), .ZN(n5319) );
  INV_X1 U2908 ( .A(n2729), .ZN(n2728) );
  OAI21_X1 U2909 ( .B1(n2539), .B2(n2732), .A(n2730), .ZN(n2729) );
  NAND2_X1 U2910 ( .A1(n3767), .A2(n2539), .ZN(n4254) );
  NAND2_X1 U2911 ( .A1(n2727), .A2(n3212), .ZN(n4253) );
  NAND2_X1 U2912 ( .A1(n3767), .A2(n3210), .ZN(n2727) );
  OAI211_X1 U2913 ( .C1(n2869), .C2(n2721), .A(n2720), .B(n2719), .ZN(n5015)
         );
  NAND2_X1 U2914 ( .A1(n3777), .A2(n2538), .ZN(n4298) );
  INV_X1 U2915 ( .A(n5326), .ZN(n4301) );
  NAND2_X1 U2916 ( .A1(n2800), .A2(DATAI_2_), .ZN(n2791) );
  NAND2_X1 U2917 ( .A1(n3123), .A2(n3125), .ZN(n3126) );
  NAND2_X1 U2918 ( .A1(n2750), .A2(n2751), .ZN(n3833) );
  OR2_X1 U2919 ( .A1(n4275), .A2(n2753), .ZN(n2750) );
  INV_X1 U2920 ( .A(n5319), .ZN(n5246) );
  INV_X1 U2921 ( .A(n5226), .ZN(n5322) );
  AND2_X1 U2922 ( .A1(n3291), .A2(n3277), .ZN(n4462) );
  AND3_X1 U2923 ( .A1(n2868), .A2(n2867), .A3(n2866), .ZN(n4453) );
  INV_X1 U2924 ( .A(n5316), .ZN(n4710) );
  INV_X1 U2925 ( .A(n3596), .ZN(n4482) );
  NAND4_X1 U2926 ( .A1(n2958), .A2(n2957), .A3(n2956), .A4(n2955), .ZN(n5053)
         );
  INV_X1 U2927 ( .A(n3482), .ZN(n4486) );
  INV_X1 U2928 ( .A(n2559), .ZN(n4986) );
  NAND2_X1 U2929 ( .A1(n4972), .A2(n2585), .ZN(n4994) );
  NAND2_X1 U2930 ( .A1(n2586), .A2(REG1_REG_1__SCAN_IN), .ZN(n2585) );
  AND2_X1 U2931 ( .A1(n2588), .A2(n2596), .ZN(n3361) );
  NAND2_X1 U2932 ( .A1(n5008), .A2(REG1_REG_4__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U2933 ( .A1(n2563), .A2(n2562), .ZN(n3354) );
  NOR2_X1 U2934 ( .A1(n2709), .A2(n3314), .ZN(n3353) );
  NOR2_X1 U2935 ( .A1(n3333), .A2(n3332), .ZN(n3331) );
  AND2_X1 U2936 ( .A1(n2709), .A2(n2562), .ZN(n3333) );
  INV_X1 U2937 ( .A(n4925), .ZN(n3383) );
  NOR2_X1 U2938 ( .A1(n3381), .A2(n3380), .ZN(n3400) );
  XNOR2_X1 U2939 ( .A(n2597), .B(n4923), .ZN(n3459) );
  OAI21_X1 U2940 ( .B1(n3409), .B2(n2574), .A(n2573), .ZN(n3581) );
  NAND2_X1 U2941 ( .A1(n2575), .A2(REG2_REG_10__SCAN_IN), .ZN(n2574) );
  NAND2_X1 U2942 ( .A1(n3454), .A2(n2575), .ZN(n2573) );
  INV_X1 U2943 ( .A(n3457), .ZN(n2575) );
  NOR2_X1 U2944 ( .A1(n4497), .A2(n4496), .ZN(n4501) );
  NAND2_X1 U2945 ( .A1(n4488), .A2(n4489), .ZN(n4493) );
  NAND2_X1 U2946 ( .A1(n4493), .A2(n2687), .ZN(n4511) );
  AND2_X1 U2947 ( .A1(n4512), .A2(n4491), .ZN(n2687) );
  XNOR2_X1 U2948 ( .A(n4520), .B(n4920), .ZN(n4509) );
  NOR2_X1 U2949 ( .A1(n4509), .A2(n4510), .ZN(n4523) );
  NAND2_X1 U2950 ( .A1(n2701), .A2(n2703), .ZN(n4542) );
  OAI211_X1 U2951 ( .C1(n4532), .C2(n2519), .A(n2580), .B(n2579), .ZN(n4541)
         );
  INV_X1 U2952 ( .A(n2581), .ZN(n2580) );
  NAND2_X1 U2953 ( .A1(n4532), .A2(n2517), .ZN(n2579) );
  OAI21_X1 U2954 ( .B1(n4531), .B2(n2519), .A(n2582), .ZN(n2581) );
  NOR2_X1 U2955 ( .A1(n4541), .A2(REG1_REG_16__SCAN_IN), .ZN(n4559) );
  NAND2_X1 U2956 ( .A1(n4555), .A2(n4554), .ZN(n4556) );
  NAND2_X1 U2957 ( .A1(n2711), .A2(n2712), .ZN(n4584) );
  NOR2_X1 U2958 ( .A1(n5331), .A2(n4452), .ZN(n2851) );
  AOI21_X1 U2959 ( .B1(n3694), .B2(n5289), .A(n3693), .ZN(n4873) );
  NAND2_X1 U2960 ( .A1(n3683), .A2(n3682), .ZN(n3694) );
  NAND2_X1 U2961 ( .A1(n2604), .A2(n2605), .ZN(n4601) );
  NAND2_X1 U2962 ( .A1(n2670), .A2(n2673), .ZN(n4593) );
  NAND2_X1 U2963 ( .A1(n2664), .A2(n2520), .ZN(n2670) );
  NAND2_X1 U2964 ( .A1(n2664), .A2(n4407), .ZN(n4610) );
  AOI21_X1 U2965 ( .B1(n4645), .B2(n3655), .A(n2540), .ZN(n4629) );
  NAND2_X1 U2966 ( .A1(n4853), .A2(n3628), .ZN(n4825) );
  NAND2_X1 U2967 ( .A1(n2675), .A2(n4419), .ZN(n3627) );
  NAND2_X1 U2968 ( .A1(n5102), .A2(n4418), .ZN(n2675) );
  NAND2_X1 U2969 ( .A1(n5305), .A2(n5177), .ZN(n4841) );
  NAND2_X1 U2970 ( .A1(n3527), .A2(n2652), .ZN(n2651) );
  NAND2_X1 U2971 ( .A1(n3291), .A2(n3268), .ZN(n5300) );
  INV_X1 U2972 ( .A(n3267), .ZN(n3268) );
  NAND2_X1 U2973 ( .A1(n2653), .A2(n2654), .ZN(n3565) );
  OR2_X1 U2974 ( .A1(n3527), .A2(n3514), .ZN(n2653) );
  NAND2_X1 U2975 ( .A1(n5305), .A2(n4592), .ZN(n4733) );
  INV_X1 U2976 ( .A(n4841), .ZN(n4863) );
  INV_X1 U2977 ( .A(n5302), .ZN(n5344) );
  INV_X1 U2978 ( .A(n5300), .ZN(n5178) );
  AND2_X1 U2979 ( .A1(n2621), .A2(n3710), .ZN(n2620) );
  INV_X1 U2980 ( .A(n2622), .ZN(n2621) );
  OAI21_X1 U2981 ( .B1(n4871), .B2(n5233), .A(n4870), .ZN(n2622) );
  INV_X1 U2982 ( .A(n4913), .ZN(n3295) );
  NAND2_X1 U2983 ( .A1(n3292), .A2(n3291), .ZN(n4954) );
  INV_X1 U2984 ( .A(n2864), .ZN(n4910) );
  AND2_X1 U2985 ( .A1(n2878), .A2(n2877), .ZN(n4911) );
  XNOR2_X1 U2986 ( .A(n2879), .B(IR_REG_25__SCAN_IN), .ZN(n4912) );
  XNOR2_X1 U2987 ( .A(n2875), .B(IR_REG_24__SCAN_IN), .ZN(n4913) );
  NAND2_X1 U2988 ( .A1(n2882), .A2(IR_REG_31__SCAN_IN), .ZN(n2875) );
  AND2_X1 U2989 ( .A1(n3301), .A2(STATE_REG_SCAN_IN), .ZN(n4930) );
  INV_X1 U2990 ( .A(n2855), .ZN(n2856) );
  INV_X1 U2991 ( .A(n4866), .ZN(n4916) );
  INV_X1 U2992 ( .A(n4592), .ZN(n5173) );
  AND2_X1 U2993 ( .A1(n2836), .A2(n2838), .ZN(n4919) );
  AND2_X1 U2994 ( .A1(n2827), .A2(n2828), .ZN(n5139) );
  AND2_X1 U2995 ( .A1(n2813), .A2(n2814), .ZN(n4926) );
  NOR2_X1 U2996 ( .A1(n2807), .A2(n2806), .ZN(n4928) );
  NOR2_X1 U2997 ( .A1(n4971), .A2(n2699), .ZN(n4976) );
  NOR2_X1 U2998 ( .A1(n4968), .A2(n2693), .ZN(n3348) );
  OAI21_X1 U2999 ( .B1(n2576), .B2(n4968), .A(n2507), .ZN(U3259) );
  XNOR2_X1 U3000 ( .A(n2578), .B(n2577), .ZN(n2576) );
  INV_X1 U3001 ( .A(n4586), .ZN(n2577) );
  AND2_X1 U3002 ( .A1(n2852), .A2(n2536), .ZN(n2859) );
  OR2_X1 U3003 ( .A1(n3400), .A2(n2548), .ZN(n2597) );
  NAND2_X1 U3004 ( .A1(n2564), .A2(n2565), .ZN(n5031) );
  XNOR2_X1 U3005 ( .A(n2790), .B(IR_REG_2__SCAN_IN), .ZN(n4989) );
  AND2_X1 U3006 ( .A1(n2568), .A2(n2567), .ZN(n2506) );
  AND2_X1 U3007 ( .A1(n2692), .A2(n2554), .ZN(n2507) );
  AND2_X1 U3008 ( .A1(n2781), .A2(n2683), .ZN(n2508) );
  AND3_X1 U3009 ( .A1(n2760), .A2(n2508), .A3(n4172), .ZN(n2509) );
  INV_X1 U3010 ( .A(n4958), .ZN(n2566) );
  AND2_X1 U3011 ( .A1(n3554), .A2(n3613), .ZN(n2510) );
  AND2_X1 U3012 ( .A1(n2510), .A2(n5105), .ZN(n2511) );
  AND2_X1 U3013 ( .A1(n2631), .A2(n4818), .ZN(n2512) );
  OR2_X1 U3014 ( .A1(n2830), .A2(IR_REG_13__SCAN_IN), .ZN(n2513) );
  NOR2_X1 U3015 ( .A1(n3149), .A2(n3148), .ZN(n2514) );
  AND2_X1 U3016 ( .A1(n4928), .A2(REG2_REG_5__SCAN_IN), .ZN(n3313) );
  AND2_X1 U3017 ( .A1(n2629), .A2(n5318), .ZN(n2515) );
  AND2_X1 U3018 ( .A1(n2633), .A2(n3656), .ZN(n2516) );
  AND2_X1 U3019 ( .A1(n4531), .A2(n4918), .ZN(n2517) );
  INV_X1 U3020 ( .A(n3418), .ZN(n3439) );
  NAND4_X1 U3021 ( .A1(n2921), .A2(n2920), .A3(n2919), .A4(n2918), .ZN(n3418)
         );
  AND2_X1 U3022 ( .A1(n3448), .A2(n4340), .ZN(n2518) );
  OR2_X1 U3023 ( .A1(n4530), .A2(n4918), .ZN(n2519) );
  INV_X1 U3024 ( .A(n2562), .ZN(n3314) );
  OAI21_X1 U3025 ( .B1(n3364), .B2(n3313), .A(n2561), .ZN(n2562) );
  AND3_X1 U3026 ( .A1(n2684), .A2(n2685), .A3(n2627), .ZN(n2852) );
  NAND2_X2 U3027 ( .A1(n2959), .A2(n5291), .ZN(n2951) );
  AND2_X1 U3028 ( .A1(n2674), .A2(n4407), .ZN(n2520) );
  AND2_X1 U3029 ( .A1(n2604), .A2(n2603), .ZN(n2521) );
  NOR2_X1 U3030 ( .A1(n3569), .A2(n3570), .ZN(n2522) );
  AND2_X1 U3031 ( .A1(n4909), .A2(n2864), .ZN(n2917) );
  AOI21_X1 U3032 ( .B1(n5259), .B2(n5260), .A(n5261), .ZN(n5308) );
  NOR2_X1 U3033 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2789)
         );
  AND3_X1 U3034 ( .A1(n4147), .A2(n4155), .A3(n2834), .ZN(n2523) );
  AND4_X1 U3035 ( .A1(n2908), .A2(n2906), .A3(n2905), .A4(n2907), .ZN(n5018)
         );
  INV_X1 U3036 ( .A(n5018), .ZN(n3417) );
  INV_X1 U3037 ( .A(n3308), .ZN(n5002) );
  AND2_X1 U3038 ( .A1(n4483), .A2(n3573), .ZN(n2524) );
  AND3_X1 U3039 ( .A1(n2935), .A2(n2934), .A3(n2933), .ZN(n2525) );
  AND2_X1 U3040 ( .A1(n2777), .A2(n2776), .ZN(n2526) );
  AND2_X1 U3041 ( .A1(n4634), .A2(n3656), .ZN(n2527) );
  NAND2_X1 U3042 ( .A1(n2685), .A2(n2684), .ZN(n2847) );
  NOR2_X1 U3043 ( .A1(n4569), .A2(n2716), .ZN(n2528) );
  AND2_X1 U3044 ( .A1(n4958), .A2(REG1_REG_0__SCAN_IN), .ZN(n2529) );
  NAND2_X1 U3045 ( .A1(n4929), .A2(n3307), .ZN(n2530) );
  INV_X1 U3046 ( .A(n2655), .ZN(n2654) );
  NAND2_X1 U3047 ( .A1(n2609), .A2(n4448), .ZN(n2531) );
  NAND2_X1 U3048 ( .A1(n2724), .A2(n2728), .ZN(n3823) );
  NOR2_X1 U3049 ( .A1(n4618), .A2(n3657), .ZN(n2532) );
  OR2_X1 U3050 ( .A1(n2874), .A2(n2780), .ZN(n2533) );
  AND2_X1 U3051 ( .A1(n4958), .A2(IR_REG_31__SCAN_IN), .ZN(n2534) );
  AND2_X1 U3052 ( .A1(n2982), .A2(n2745), .ZN(n2535) );
  AND2_X1 U3053 ( .A1(n2760), .A2(n2508), .ZN(n2536) );
  NOR2_X1 U3054 ( .A1(n2639), .A2(n4797), .ZN(n2638) );
  NAND3_X1 U3055 ( .A1(n2685), .A2(n2684), .A3(n2526), .ZN(n2537) );
  INV_X1 U3056 ( .A(IR_REG_29__SCAN_IN), .ZN(n4172) );
  OR2_X1 U3057 ( .A1(n3039), .A2(n3038), .ZN(n2538) );
  AND2_X1 U3058 ( .A1(n3211), .A2(n3210), .ZN(n2539) );
  AND2_X1 U3059 ( .A1(n4668), .A2(n4257), .ZN(n2540) );
  INV_X1 U3060 ( .A(IR_REG_19__SCAN_IN), .ZN(n2777) );
  AOI21_X1 U3061 ( .B1(n4719), .B2(n3651), .A(n2763), .ZN(n4700) );
  INV_X1 U3062 ( .A(IR_REG_20__SCAN_IN), .ZN(n2776) );
  OAI21_X1 U3063 ( .B1(n2800), .B2(n5039), .A(n2791), .ZN(n3416) );
  INV_X1 U3064 ( .A(n3416), .ZN(n3487) );
  OR2_X1 U3065 ( .A1(n4692), .A2(n4671), .ZN(n2541) );
  INV_X1 U3066 ( .A(n4818), .ZN(n3757) );
  NOR2_X1 U3067 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2817)
         );
  INV_X1 U3068 ( .A(n4796), .ZN(n5193) );
  NOR2_X1 U3069 ( .A1(n3313), .A2(n2561), .ZN(n2542) );
  NOR2_X1 U3070 ( .A1(n4501), .A2(n4500), .ZN(n2543) );
  AND2_X1 U3071 ( .A1(n4849), .A2(n4832), .ZN(n2544) );
  NAND2_X1 U3072 ( .A1(n4815), .A2(n4391), .ZN(n2545) );
  NAND2_X1 U3073 ( .A1(n3111), .A2(n3849), .ZN(n2546) );
  INV_X1 U3074 ( .A(n5160), .ZN(n5163) );
  NOR2_X1 U3075 ( .A1(n4523), .A2(n4524), .ZN(n2547) );
  AND2_X1 U3076 ( .A1(n4924), .A2(REG1_REG_9__SCAN_IN), .ZN(n2548) );
  AND2_X1 U3077 ( .A1(n2512), .A2(n4796), .ZN(n2549) );
  AND2_X1 U3078 ( .A1(n3054), .A2(n2538), .ZN(n2550) );
  INV_X1 U3079 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2698) );
  INV_X1 U3080 ( .A(DATAI_0_), .ZN(n2721) );
  NAND2_X1 U3081 ( .A1(n2651), .A2(n2650), .ZN(n3601) );
  INV_X1 U3082 ( .A(IR_REG_13__SCAN_IN), .ZN(n2775) );
  NOR2_X1 U3083 ( .A1(n2758), .A2(n2830), .ZN(n2843) );
  INV_X1 U3084 ( .A(n5225), .ZN(n2738) );
  NAND2_X1 U3085 ( .A1(n4825), .A2(n4826), .ZN(n4824) );
  NOR2_X1 U3086 ( .A1(n2830), .A2(n2759), .ZN(n2840) );
  AND2_X1 U3087 ( .A1(n4334), .A2(n4331), .ZN(n4393) );
  INV_X1 U3088 ( .A(n4393), .ZN(n2681) );
  NOR2_X1 U3089 ( .A1(n3455), .A2(n3454), .ZN(n2551) );
  AND2_X1 U3090 ( .A1(n3300), .A2(DATAI_22_), .ZN(n4694) );
  XNOR2_X1 U3091 ( .A(n2723), .B(n3978), .ZN(n2870) );
  INV_X1 U3092 ( .A(IR_REG_28__SCAN_IN), .ZN(n2683) );
  INV_X1 U3093 ( .A(n4920), .ZN(n4521) );
  INV_X1 U3094 ( .A(n4729), .ZN(n2630) );
  NAND2_X1 U3095 ( .A1(n2560), .A2(n2542), .ZN(n2563) );
  OR2_X1 U3096 ( .A1(n4591), .A2(n4592), .ZN(n2552) );
  NOR2_X1 U3097 ( .A1(n3091), .A2(n3090), .ZN(n2553) );
  INV_X1 U3098 ( .A(n3804), .ZN(n3448) );
  AND2_X1 U3099 ( .A1(n4590), .A2(n2552), .ZN(n2554) );
  NOR2_X1 U3100 ( .A1(n4999), .A2(n3311), .ZN(n2555) );
  NAND2_X1 U3101 ( .A1(n4917), .A2(REG2_REG_18__SCAN_IN), .ZN(n2556) );
  INV_X1 U3102 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2691) );
  INV_X1 U3103 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2594) );
  INV_X1 U3104 ( .A(n4978), .ZN(n2567) );
  INV_X1 U3105 ( .A(n4988), .ZN(n2557) );
  INV_X1 U3106 ( .A(n3364), .ZN(n2560) );
  INV_X1 U3107 ( .A(n4927), .ZN(n2561) );
  NAND3_X1 U3108 ( .A1(n2564), .A2(n2565), .A3(REG2_REG_1__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U3109 ( .A1(n4539), .A2(n4540), .ZN(n4558) );
  NAND2_X1 U3110 ( .A1(n4530), .A2(n4918), .ZN(n2582) );
  INV_X1 U3111 ( .A(n5031), .ZN(n2586) );
  OAI21_X1 U3112 ( .B1(n5031), .B2(REG1_REG_1__SCAN_IN), .A(n2587), .ZN(n4973)
         );
  NAND2_X1 U3113 ( .A1(n5031), .A2(REG1_REG_1__SCAN_IN), .ZN(n2587) );
  NAND2_X1 U3114 ( .A1(n2689), .A2(n5002), .ZN(n2596) );
  NAND2_X1 U3115 ( .A1(n3498), .A2(n2768), .ZN(n2601) );
  NAND2_X1 U3116 ( .A1(n5049), .A2(n3480), .ZN(n2602) );
  INV_X1 U3117 ( .A(n2609), .ZN(n4613) );
  NAND2_X1 U3118 ( .A1(n4843), .A2(n2614), .ZN(n2611) );
  NAND2_X1 U3119 ( .A1(n2611), .A2(n2612), .ZN(n4431) );
  AND3_X2 U3120 ( .A1(n2862), .A2(n2863), .A3(n2865), .ZN(n2932) );
  XNOR2_X1 U3121 ( .A(n3703), .B(n4427), .ZN(n2619) );
  NAND2_X1 U3122 ( .A1(n2623), .A2(n2620), .ZN(n4899) );
  NAND2_X1 U3123 ( .A1(n2623), .A2(n3710), .ZN(n3711) );
  AND3_X2 U3124 ( .A1(n2624), .A2(n2773), .A3(n2772), .ZN(n2684) );
  NAND2_X1 U3125 ( .A1(n2523), .A2(n2625), .ZN(n2758) );
  NAND3_X1 U3126 ( .A1(n3448), .A2(n3487), .A3(n4340), .ZN(n5047) );
  NAND2_X1 U3127 ( .A1(n2786), .A2(n2586), .ZN(n2788) );
  NAND2_X2 U3128 ( .A1(n4341), .A2(n4343), .ZN(n3419) );
  NOR2_X1 U3129 ( .A1(n3702), .A2(n3701), .ZN(n3703) );
  NAND2_X1 U3130 ( .A1(n3479), .A2(n3478), .ZN(n5049) );
  NAND2_X1 U3131 ( .A1(n2878), .A2(IR_REG_31__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U3132 ( .A1(n3658), .A2(n4331), .ZN(n4845) );
  NAND2_X1 U3133 ( .A1(n2785), .A2(n2781), .ZN(n2783) );
  INV_X1 U3134 ( .A(n4853), .ZN(n2641) );
  NAND2_X1 U3135 ( .A1(n2635), .A2(n2636), .ZN(n3629) );
  NAND2_X1 U3136 ( .A1(n4853), .A2(n2638), .ZN(n2635) );
  NAND2_X1 U3137 ( .A1(n3527), .A2(n2647), .ZN(n2646) );
  NOR2_X1 U3138 ( .A1(n4484), .A2(n3545), .ZN(n2655) );
  NAND2_X1 U3139 ( .A1(n4645), .A2(n2662), .ZN(n2661) );
  NAND2_X1 U3140 ( .A1(n2852), .A2(n2509), .ZN(n2863) );
  INV_X1 U3141 ( .A(n2758), .ZN(n2685) );
  NAND3_X1 U3142 ( .A1(n2773), .A2(n2772), .A3(n2686), .ZN(n2830) );
  NAND2_X1 U3143 ( .A1(n3463), .A2(n3462), .ZN(n3583) );
  NAND2_X1 U3144 ( .A1(n2695), .A2(n2694), .ZN(n2693) );
  NAND2_X1 U3145 ( .A1(n3347), .A2(n5069), .ZN(n2694) );
  INV_X1 U3146 ( .A(n3347), .ZN(n2696) );
  NAND2_X1 U3147 ( .A1(n5031), .A2(n2698), .ZN(n2697) );
  NOR2_X1 U31480 ( .A1(n4591), .A2(n5031), .ZN(n2699) );
  INV_X1 U31490 ( .A(IR_REG_1__SCAN_IN), .ZN(n2700) );
  OAI21_X1 U3150 ( .B1(n5001), .B2(n2706), .A(n2705), .ZN(n3364) );
  AND2_X1 U3151 ( .A1(n5139), .A2(REG2_REG_11__SCAN_IN), .ZN(n2708) );
  NOR2_X1 U3152 ( .A1(n4556), .A2(n4557), .ZN(n4569) );
  NAND3_X1 U3153 ( .A1(n2870), .A2(n2869), .A3(n4958), .ZN(n2719) );
  OR2_X1 U3154 ( .A1(n2870), .A2(n2721), .ZN(n2720) );
  INV_X1 U3155 ( .A(n2859), .ZN(n2722) );
  NAND2_X1 U3156 ( .A1(n3764), .A2(n2725), .ZN(n2724) );
  NAND2_X1 U3157 ( .A1(n3777), .A2(n2550), .ZN(n3814) );
  NAND2_X1 U3158 ( .A1(n5222), .A2(n2735), .ZN(n2734) );
  INV_X1 U3159 ( .A(n2743), .ZN(n2741) );
  NAND2_X1 U3160 ( .A1(n3572), .A2(n2535), .ZN(n2742) );
  INV_X1 U3161 ( .A(n3743), .ZN(n2744) );
  NAND2_X1 U3162 ( .A1(n2746), .A2(n2747), .ZN(n3122) );
  NAND2_X1 U3163 ( .A1(n4275), .A2(n2748), .ZN(n2746) );
  NAND2_X1 U3164 ( .A1(n3225), .A2(n3224), .ZN(n3824) );
  NAND2_X1 U3165 ( .A1(n3824), .A2(n3226), .ZN(n4309) );
  INV_X1 U3166 ( .A(n3723), .ZN(n3718) );
  NAND2_X1 U3167 ( .A1(n2852), .A2(n4164), .ZN(n2874) );
  OAI21_X1 U3168 ( .B1(n5018), .B2(n2951), .A(n2915), .ZN(n2916) );
  NAND2_X1 U3169 ( .A1(n3471), .A2(n3487), .ZN(n4345) );
  OR2_X1 U3170 ( .A1(n2876), .A2(n4179), .ZN(n2877) );
  NOR2_X1 U3171 ( .A1(n3718), .A2(n3258), .ZN(n3264) );
  NAND2_X1 U3172 ( .A1(n2928), .A2(n2916), .ZN(n2930) );
  INV_X2 U3173 ( .A(n5348), .ZN(n5305) );
  AND2_X2 U3174 ( .A1(n2902), .A2(n3431), .ZN(n5343) );
  AND2_X2 U3175 ( .A1(n2902), .A2(n3261), .ZN(n5339) );
  INV_X2 U3176 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  AND2_X1 U3177 ( .A1(n3415), .A2(n3414), .ZN(n5115) );
  NAND2_X1 U3178 ( .A1(n3424), .A2(n3727), .ZN(n4869) );
  INV_X1 U3179 ( .A(U4043), .ZN(n4485) );
  AND2_X1 U3180 ( .A1(n3663), .A2(n3662), .ZN(n4803) );
  INV_X1 U3181 ( .A(n4803), .ZN(n3664) );
  NOR2_X1 U3182 ( .A1(n3650), .A2(n3649), .ZN(n2763) );
  OR2_X1 U3183 ( .A1(n3288), .A2(n2566), .ZN(n2764) );
  NOR2_X1 U3184 ( .A1(n4799), .A2(n4797), .ZN(n2765) );
  AND2_X1 U3185 ( .A1(n2922), .A2(n2764), .ZN(n2766) );
  AND2_X1 U3186 ( .A1(n5015), .A2(n2959), .ZN(n2767) );
  OR2_X1 U3187 ( .A1(n5053), .A2(n3493), .ZN(n2768) );
  INV_X1 U3188 ( .A(n2916), .ZN(n2929) );
  XNOR2_X1 U3189 ( .A(n2914), .B(n3727), .ZN(n2928) );
  AND2_X1 U3190 ( .A1(n4738), .A2(n3665), .ZN(n4752) );
  INV_X1 U3191 ( .A(IR_REG_24__SCAN_IN), .ZN(n2779) );
  INV_X1 U3192 ( .A(n3124), .ZN(n3125) );
  INV_X1 U3193 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4258) );
  INV_X1 U3194 ( .A(IR_REG_21__SCAN_IN), .ZN(n2778) );
  INV_X1 U3195 ( .A(n4287), .ZN(n3185) );
  OR2_X1 U3196 ( .A1(n3199), .A2(n4258), .ZN(n3213) );
  AND2_X1 U3197 ( .A1(n3684), .A2(n3271), .ZN(n3733) );
  NOR2_X1 U3198 ( .A1(n3178), .A2(n3177), .ZN(n3187) );
  INV_X1 U3199 ( .A(n3501), .ZN(n3573) );
  AOI21_X1 U3200 ( .B1(n4469), .B2(n5054), .A(n3709), .ZN(n3710) );
  INV_X1 U3201 ( .A(n5105), .ZN(n5119) );
  AND2_X1 U3202 ( .A1(n4398), .A2(n4397), .ZN(n5058) );
  INV_X1 U3203 ( .A(n5015), .ZN(n4340) );
  INV_X1 U3204 ( .A(n3721), .ZN(n3258) );
  AND2_X1 U3205 ( .A1(n3778), .A2(n3776), .ZN(n3035) );
  NAND2_X1 U3206 ( .A1(n2800), .A2(DATAI_1_), .ZN(n2787) );
  OAI22_X1 U3207 ( .A1(n3827), .A2(n2951), .B1(n3726), .B2(n4656), .ZN(n4255)
         );
  OR2_X1 U3208 ( .A1(n3281), .A2(n3279), .ZN(n3793) );
  AND2_X1 U3209 ( .A1(n3270), .A2(n3243), .ZN(n4595) );
  INV_X1 U32100 ( .A(n3291), .ZN(n3302) );
  NOR2_X1 U32110 ( .A1(n3331), .A2(n3316), .ZN(n3384) );
  INV_X1 U32120 ( .A(n3453), .ZN(n3454) );
  INV_X1 U32130 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3840) );
  INV_X1 U32140 ( .A(n5213), .ZN(n4570) );
  AND2_X1 U32150 ( .A1(n3300), .A2(DATAI_26_), .ZN(n4621) );
  OR2_X1 U32160 ( .A1(n5291), .A2(n4592), .ZN(n3267) );
  INV_X1 U32170 ( .A(n5054), .ZN(n5286) );
  OR2_X1 U32180 ( .A1(n4733), .A2(n5291), .ZN(n5302) );
  OR2_X1 U32190 ( .A1(n3692), .A2(n3691), .ZN(n3693) );
  AND2_X1 U32200 ( .A1(n5174), .A2(n5167), .ZN(n5172) );
  NAND2_X1 U32210 ( .A1(n5014), .A2(n4916), .ZN(n5327) );
  INV_X1 U32220 ( .A(n3657), .ZN(n4603) );
  AND2_X1 U32230 ( .A1(n3300), .A2(DATAI_23_), .ZN(n3769) );
  NOR2_X1 U32240 ( .A1(n3127), .A2(n4577), .ZN(n3140) );
  INV_X1 U32250 ( .A(n3150), .ZN(n3151) );
  INV_X1 U32260 ( .A(n4747), .ZN(n5227) );
  INV_X1 U32270 ( .A(n3793), .ZN(n5243) );
  AND4_X1 U32280 ( .A1(n3275), .A2(n3274), .A3(n3273), .A4(n3272), .ZN(n4607)
         );
  AND4_X1 U32290 ( .A1(n3192), .A2(n3191), .A3(n3190), .A4(n3189), .ZN(n4692)
         );
  AND4_X1 U32300 ( .A1(n3118), .A2(n3117), .A3(n3116), .A4(n3115), .ZN(n4775)
         );
  INV_X1 U32310 ( .A(n4550), .ZN(n5010) );
  INV_X1 U32320 ( .A(n4919), .ZN(n4536) );
  OR2_X1 U32330 ( .A1(n4966), .A2(n3319), .ZN(n4968) );
  AND2_X1 U32340 ( .A1(n2869), .A2(n3298), .ZN(n5283) );
  INV_X1 U32350 ( .A(n4733), .ZN(n4838) );
  INV_X1 U32360 ( .A(n5115), .ZN(n5289) );
  AOI21_X1 U32370 ( .B1(n2900), .B2(n4173), .A(n2899), .ZN(n3261) );
  NAND2_X2 U32380 ( .A1(n5014), .A2(n4866), .ZN(n5291) );
  INV_X1 U32390 ( .A(n3261), .ZN(n3431) );
  AND2_X1 U32400 ( .A1(n3288), .A2(n4930), .ZN(n3291) );
  INV_X1 U32410 ( .A(n4930), .ZN(n3293) );
  NAND2_X1 U32420 ( .A1(n3263), .A2(n3276), .ZN(n5226) );
  AND2_X1 U32430 ( .A1(n3282), .A2(n3374), .ZN(n5326) );
  INV_X1 U32440 ( .A(n4634), .ZN(n4604) );
  INV_X1 U32450 ( .A(n4485), .ZN(n4481) );
  INV_X1 U32460 ( .A(n3504), .ZN(n4484) );
  OR2_X1 U32470 ( .A1(n4966), .A2(n4981), .ZN(n4591) );
  INV_X1 U32480 ( .A(n5339), .ZN(n5337) );
  AND3_X1 U32490 ( .A1(n5087), .A2(n5086), .A3(n5085), .ZN(n5089) );
  INV_X1 U32500 ( .A(n5343), .ZN(n5340) );
  INV_X1 U32510 ( .A(n4954), .ZN(n4956) );
  NOR2_X1 U32520 ( .A1(n3288), .A2(n3293), .ZN(U4043) );
  NAND2_X1 U32530 ( .A1(n2783), .A2(IR_REG_31__SCAN_IN), .ZN(n2782) );
  INV_X1 U32540 ( .A(n2800), .ZN(n2786) );
  NAND2_X2 U32550 ( .A1(n2788), .A2(n2787), .ZN(n3804) );
  OR2_X1 U32560 ( .A1(n2789), .A2(n2841), .ZN(n2790) );
  INV_X1 U32570 ( .A(n4989), .ZN(n5039) );
  AND2_X1 U32580 ( .A1(n2789), .A2(n2792), .ZN(n2802) );
  INV_X1 U32590 ( .A(IR_REG_31__SCAN_IN), .ZN(n2841) );
  NOR2_X1 U32600 ( .A1(n2802), .A2(n2841), .ZN(n2793) );
  NAND2_X1 U32610 ( .A1(n2793), .A2(IR_REG_3__SCAN_IN), .ZN(n2796) );
  INV_X1 U32620 ( .A(n2793), .ZN(n2795) );
  INV_X1 U32630 ( .A(IR_REG_3__SCAN_IN), .ZN(n2794) );
  NAND2_X1 U32640 ( .A1(n2795), .A2(n2794), .ZN(n2797) );
  MUX2_X1 U32650 ( .A(n4929), .B(DATAI_3_), .S(n2800), .Z(n5048) );
  NAND2_X1 U32660 ( .A1(n2797), .A2(IR_REG_31__SCAN_IN), .ZN(n2799) );
  INV_X1 U32670 ( .A(IR_REG_4__SCAN_IN), .ZN(n2798) );
  XNOR2_X1 U32680 ( .A(n2799), .B(n2798), .ZN(n3308) );
  INV_X1 U32690 ( .A(DATAI_4_), .ZN(n4085) );
  MUX2_X1 U32700 ( .A(n3308), .B(n4085), .S(n3300), .Z(n3493) );
  NAND2_X1 U32710 ( .A1(n5046), .A2(n3493), .ZN(n3525) );
  NOR2_X1 U32720 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2801)
         );
  AND2_X1 U32730 ( .A1(n2802), .A2(n2801), .ZN(n2805) );
  NOR2_X1 U32740 ( .A1(n2805), .A2(n2841), .ZN(n2803) );
  MUX2_X1 U32750 ( .A(n2841), .B(n2803), .S(IR_REG_5__SCAN_IN), .Z(n2807) );
  INV_X1 U32760 ( .A(IR_REG_5__SCAN_IN), .ZN(n2804) );
  NAND2_X1 U32770 ( .A1(n2805), .A2(n2804), .ZN(n2819) );
  INV_X1 U32780 ( .A(n2819), .ZN(n2806) );
  MUX2_X1 U32790 ( .A(n4928), .B(DATAI_5_), .S(n3300), .Z(n3545) );
  NAND2_X1 U32800 ( .A1(n2819), .A2(IR_REG_31__SCAN_IN), .ZN(n2809) );
  INV_X1 U32810 ( .A(IR_REG_6__SCAN_IN), .ZN(n2808) );
  XNOR2_X1 U32820 ( .A(n2809), .B(n2808), .ZN(n4927) );
  INV_X1 U32830 ( .A(DATAI_6_), .ZN(n4081) );
  MUX2_X1 U32840 ( .A(n4927), .B(n4081), .S(n3300), .Z(n3501) );
  NAND2_X1 U32850 ( .A1(n2810), .A2(IR_REG_31__SCAN_IN), .ZN(n2812) );
  INV_X1 U32860 ( .A(n2812), .ZN(n2811) );
  NAND2_X1 U32870 ( .A1(n2811), .A2(IR_REG_7__SCAN_IN), .ZN(n2813) );
  NAND2_X1 U32880 ( .A1(n2812), .A2(n4140), .ZN(n2814) );
  MUX2_X1 U32890 ( .A(n4926), .B(DATAI_7_), .S(n3300), .Z(n3745) );
  INV_X1 U32900 ( .A(n3745), .ZN(n3554) );
  NAND2_X1 U32910 ( .A1(n2814), .A2(IR_REG_31__SCAN_IN), .ZN(n2815) );
  XNOR2_X1 U32920 ( .A(n2815), .B(IR_REG_8__SCAN_IN), .ZN(n4925) );
  INV_X1 U32930 ( .A(DATAI_8_), .ZN(n2816) );
  MUX2_X1 U32940 ( .A(n3383), .B(n2816), .S(n3300), .Z(n3613) );
  NAND2_X1 U32950 ( .A1(n2817), .A2(n4141), .ZN(n2818) );
  OAI21_X1 U32960 ( .B1(n2819), .B2(n2818), .A(IR_REG_31__SCAN_IN), .ZN(n2820)
         );
  MUX2_X1 U32970 ( .A(IR_REG_31__SCAN_IN), .B(n2820), .S(IR_REG_9__SCAN_IN), 
        .Z(n2822) );
  NAND2_X1 U32980 ( .A1(n2822), .A2(n2821), .ZN(n3405) );
  INV_X1 U32990 ( .A(DATAI_9_), .ZN(n4071) );
  MUX2_X1 U33000 ( .A(n3405), .B(n4071), .S(n3300), .Z(n5105) );
  NAND2_X1 U33010 ( .A1(n2821), .A2(IR_REG_31__SCAN_IN), .ZN(n2823) );
  XNOR2_X1 U33020 ( .A(n2823), .B(IR_REG_10__SCAN_IN), .ZN(n4923) );
  MUX2_X1 U33030 ( .A(n4923), .B(DATAI_10_), .S(n3300), .Z(n3782) );
  OR2_X1 U33040 ( .A1(n2824), .A2(n2841), .ZN(n2826) );
  INV_X1 U33050 ( .A(n2826), .ZN(n2825) );
  NAND2_X1 U33060 ( .A1(n2825), .A2(IR_REG_11__SCAN_IN), .ZN(n2827) );
  NAND2_X1 U33070 ( .A1(n2826), .A2(n4146), .ZN(n2828) );
  MUX2_X1 U33080 ( .A(n5139), .B(DATAI_11_), .S(n3300), .Z(n4846) );
  NAND2_X1 U33090 ( .A1(n2828), .A2(IR_REG_31__SCAN_IN), .ZN(n2829) );
  XNOR2_X1 U33100 ( .A(n2829), .B(IR_REG_12__SCAN_IN), .ZN(n4922) );
  MUX2_X1 U33110 ( .A(n4922), .B(DATAI_12_), .S(n3300), .Z(n4829) );
  NAND2_X1 U33120 ( .A1(n2830), .A2(IR_REG_31__SCAN_IN), .ZN(n2831) );
  XNOR2_X1 U33130 ( .A(n2831), .B(n2775), .ZN(n4507) );
  INV_X1 U33140 ( .A(DATAI_13_), .ZN(n4070) );
  MUX2_X1 U33150 ( .A(n4507), .B(n4070), .S(n3300), .Z(n5160) );
  NAND2_X1 U33160 ( .A1(n2513), .A2(IR_REG_31__SCAN_IN), .ZN(n2832) );
  XNOR2_X1 U33170 ( .A(n2832), .B(IR_REG_14__SCAN_IN), .ZN(n4920) );
  INV_X1 U33180 ( .A(DATAI_14_), .ZN(n4062) );
  MUX2_X1 U33190 ( .A(n4521), .B(n4062), .S(n3300), .Z(n4818) );
  NAND2_X1 U33200 ( .A1(n2832), .A2(n4147), .ZN(n2833) );
  NAND2_X1 U33210 ( .A1(n2833), .A2(IR_REG_31__SCAN_IN), .ZN(n2835) );
  OR2_X1 U33220 ( .A1(n2835), .A2(n2834), .ZN(n2836) );
  NAND2_X1 U33230 ( .A1(n2835), .A2(n2834), .ZN(n2838) );
  INV_X1 U33240 ( .A(DATAI_15_), .ZN(n2837) );
  MUX2_X1 U33250 ( .A(n4536), .B(n2837), .S(n3300), .Z(n4796) );
  NAND2_X1 U33260 ( .A1(n2838), .A2(IR_REG_31__SCAN_IN), .ZN(n2839) );
  XNOR2_X1 U33270 ( .A(n2839), .B(IR_REG_16__SCAN_IN), .ZN(n4918) );
  INV_X1 U33280 ( .A(n4918), .ZN(n4552) );
  INV_X1 U33290 ( .A(DATAI_16_), .ZN(n3872) );
  MUX2_X1 U33300 ( .A(n4552), .B(n3872), .S(n3300), .Z(n4779) );
  NAND2_X1 U33310 ( .A1(n4804), .A2(n4779), .ZN(n4781) );
  NOR2_X1 U33320 ( .A1(n2840), .A2(n2841), .ZN(n2842) );
  MUX2_X1 U33330 ( .A(n2841), .B(n2842), .S(IR_REG_17__SCAN_IN), .Z(n2844) );
  OR2_X1 U33340 ( .A1(n2844), .A2(n2843), .ZN(n5213) );
  MUX2_X1 U33350 ( .A(n4570), .B(DATAI_17_), .S(n3300), .Z(n4761) );
  OR2_X1 U33360 ( .A1(n2843), .A2(n2841), .ZN(n2845) );
  XNOR2_X1 U33370 ( .A(n2845), .B(IR_REG_18__SCAN_IN), .ZN(n4917) );
  INV_X1 U33380 ( .A(n4917), .ZN(n4581) );
  INV_X1 U33390 ( .A(DATAI_18_), .ZN(n2846) );
  MUX2_X1 U33400 ( .A(n4581), .B(n2846), .S(n3300), .Z(n4747) );
  NAND2_X1 U33410 ( .A1(n2847), .A2(IR_REG_31__SCAN_IN), .ZN(n2848) );
  INV_X1 U33420 ( .A(DATAI_19_), .ZN(n2850) );
  MUX2_X1 U33430 ( .A(n4592), .B(n2850), .S(n3300), .Z(n4729) );
  NAND2_X1 U33440 ( .A1(n3300), .A2(DATAI_20_), .ZN(n5276) );
  NAND2_X1 U33450 ( .A1(n3300), .A2(DATAI_21_), .ZN(n5318) );
  INV_X1 U33460 ( .A(n5318), .ZN(n4711) );
  NAND2_X1 U33470 ( .A1(n3300), .A2(DATAI_24_), .ZN(n4656) );
  NAND2_X1 U33480 ( .A1(n3300), .A2(DATAI_27_), .ZN(n3657) );
  NAND2_X1 U33490 ( .A1(n4594), .A2(n3724), .ZN(n3712) );
  NAND2_X1 U33500 ( .A1(n3300), .A2(DATAI_29_), .ZN(n4372) );
  INV_X1 U33510 ( .A(n4372), .ZN(n4378) );
  NAND2_X1 U33520 ( .A1(n3300), .A2(DATAI_30_), .ZN(n5330) );
  INV_X1 U3353 ( .A(n5330), .ZN(n4452) );
  AND2_X1 U33540 ( .A1(n3300), .A2(DATAI_31_), .ZN(n4456) );
  XNOR2_X1 U3355 ( .A(n2851), .B(n4456), .ZN(n5345) );
  OR2_X1 U3356 ( .A1(n2852), .A2(n2841), .ZN(n2853) );
  NAND2_X1 U3357 ( .A1(n2537), .A2(IR_REG_31__SCAN_IN), .ZN(n2854) );
  MUX2_X1 U3358 ( .A(IR_REG_31__SCAN_IN), .B(n2854), .S(IR_REG_21__SCAN_IN), 
        .Z(n2855) );
  NOR2_X2 U3359 ( .A1(n2856), .A2(n2852), .ZN(n4915) );
  NAND2_X1 U3360 ( .A1(n2857), .A2(IR_REG_31__SCAN_IN), .ZN(n2858) );
  OAI21_X1 U3361 ( .B1(n2859), .B2(n2841), .A(IR_REG_29__SCAN_IN), .ZN(n2861)
         );
  NAND2_X1 U3362 ( .A1(n2861), .A2(n2860), .ZN(n2862) );
  NAND2_X1 U3363 ( .A1(n2932), .A2(REG1_REG_31__SCAN_IN), .ZN(n2868) );
  INV_X1 U3364 ( .A(n2865), .ZN(n4909) );
  NAND2_X1 U3365 ( .A1(n3704), .A2(REG2_REG_31__SCAN_IN), .ZN(n2867) );
  AND2_X2 U3366 ( .A1(n2865), .A2(n2864), .ZN(n2931) );
  NAND2_X1 U3367 ( .A1(n2931), .A2(REG0_REG_31__SCAN_IN), .ZN(n2866) );
  NAND2_X1 U3368 ( .A1(n4914), .A2(n4915), .ZN(n3424) );
  INV_X1 U3369 ( .A(B_REG_SCAN_IN), .ZN(n2871) );
  OR2_X1 U3370 ( .A1(n2870), .A2(n2871), .ZN(n2872) );
  NAND2_X1 U3371 ( .A1(n5283), .A2(n2872), .ZN(n3708) );
  NOR2_X1 U3372 ( .A1(n4453), .A2(n3708), .ZN(n5329) );
  AOI21_X1 U3373 ( .B1(n4456), .B2(n5282), .A(n5329), .ZN(n5347) );
  INV_X1 U3374 ( .A(n5347), .ZN(n2873) );
  AOI21_X1 U3375 ( .B1(n5345), .B2(n5335), .A(n2873), .ZN(n2904) );
  NAND2_X1 U3376 ( .A1(n2874), .A2(IR_REG_31__SCAN_IN), .ZN(n2880) );
  NAND2_X1 U3377 ( .A1(n2533), .A2(IR_REG_31__SCAN_IN), .ZN(n2879) );
  OR2_X1 U3378 ( .A1(n2880), .A2(n3965), .ZN(n2881) );
  NAND2_X1 U3379 ( .A1(n4866), .A2(n4592), .ZN(n2883) );
  NAND2_X1 U3380 ( .A1(n3298), .A2(n2883), .ZN(n3277) );
  INV_X1 U3381 ( .A(n4912), .ZN(n3294) );
  NAND2_X1 U3382 ( .A1(n3295), .A2(n3294), .ZN(n2884) );
  MUX2_X1 U3383 ( .A(n3295), .B(n2884), .S(B_REG_SCAN_IN), .Z(n2885) );
  NOR4_X1 U3384 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2886) );
  INV_X1 U3385 ( .A(D_REG_8__SCAN_IN), .ZN(n4934) );
  INV_X1 U3386 ( .A(D_REG_14__SCAN_IN), .ZN(n4939) );
  NAND3_X1 U3387 ( .A1(n2886), .A2(n4934), .A3(n4939), .ZN(n2892) );
  NOR4_X1 U3388 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_27__SCAN_IN), .ZN(n2890) );
  NOR4_X1 U3389 ( .A1(D_REG_19__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2889) );
  NOR4_X1 U3390 ( .A1(D_REG_21__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2888) );
  NOR4_X1 U3391 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_31__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2887) );
  NAND4_X1 U3392 ( .A1(n2890), .A2(n2889), .A3(n2888), .A4(n2887), .ZN(n2891)
         );
  NOR4_X1 U3393 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(n2892), 
        .A4(n2891), .ZN(n2895) );
  INV_X1 U3394 ( .A(D_REG_12__SCAN_IN), .ZN(n4937) );
  INV_X1 U3395 ( .A(D_REG_23__SCAN_IN), .ZN(n4947) );
  INV_X1 U3396 ( .A(D_REG_22__SCAN_IN), .ZN(n4946) );
  INV_X1 U3397 ( .A(D_REG_16__SCAN_IN), .ZN(n4941) );
  NAND4_X1 U3398 ( .A1(n4937), .A2(n4947), .A3(n4946), .A4(n4941), .ZN(n2893)
         );
  NOR3_X1 U3399 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(n2893), 
        .ZN(n2894) );
  NAND2_X1 U3400 ( .A1(n2895), .A2(n2894), .ZN(n2896) );
  OAI22_X1 U3401 ( .A1(n3292), .A2(D_REG_1__SCAN_IN), .B1(n4911), .B2(n4912), 
        .ZN(n3259) );
  NAND2_X1 U3402 ( .A1(n3259), .A2(n3267), .ZN(n2897) );
  INV_X1 U3403 ( .A(D_REG_0__SCAN_IN), .ZN(n4173) );
  INV_X1 U3404 ( .A(n4911), .ZN(n2898) );
  NOR2_X1 U3405 ( .A1(n5339), .A2(REG1_REG_31__SCAN_IN), .ZN(n2901) );
  AOI21_X1 U3406 ( .B1(n2904), .B2(n5339), .A(n2901), .ZN(U3549) );
  NOR2_X1 U3407 ( .A1(n5343), .A2(REG0_REG_31__SCAN_IN), .ZN(n2903) );
  AOI21_X1 U3408 ( .B1(n2904), .B2(n5343), .A(n2903), .ZN(U3517) );
  NAND2_X1 U3409 ( .A1(n2945), .A2(REG3_REG_1__SCAN_IN), .ZN(n2908) );
  NAND2_X1 U3410 ( .A1(n2931), .A2(REG0_REG_1__SCAN_IN), .ZN(n2905) );
  NAND2_X1 U3411 ( .A1(n4915), .A2(n4866), .ZN(n2913) );
  INV_X1 U3412 ( .A(n2913), .ZN(n2909) );
  NAND2_X1 U3413 ( .A1(n3417), .A2(n3004), .ZN(n2911) );
  NAND2_X1 U3414 ( .A1(n3804), .A2(n2959), .ZN(n2910) );
  NAND2_X1 U3415 ( .A1(n2911), .A2(n2910), .ZN(n2914) );
  NAND2_X1 U3416 ( .A1(n4914), .A2(n4592), .ZN(n2912) );
  NAND2_X1 U3417 ( .A1(n3804), .A2(n3004), .ZN(n2915) );
  XNOR2_X1 U3418 ( .A(n2928), .B(n2929), .ZN(n3802) );
  NAND2_X1 U3419 ( .A1(n2917), .A2(REG2_REG_0__SCAN_IN), .ZN(n2921) );
  NAND2_X1 U3420 ( .A1(n2945), .A2(REG3_REG_0__SCAN_IN), .ZN(n2920) );
  NAND2_X1 U3421 ( .A1(n2931), .A2(REG0_REG_0__SCAN_IN), .ZN(n2919) );
  NAND2_X1 U3422 ( .A1(n2932), .A2(REG1_REG_0__SCAN_IN), .ZN(n2918) );
  INV_X1 U3423 ( .A(n2926), .ZN(n2927) );
  NAND2_X1 U3424 ( .A1(n5015), .A2(n3004), .ZN(n2922) );
  INV_X1 U3425 ( .A(n3288), .ZN(n2924) );
  NAND2_X1 U3426 ( .A1(n2924), .A2(REG1_REG_0__SCAN_IN), .ZN(n2925) );
  NAND2_X1 U3427 ( .A1(n2926), .A2(n2925), .ZN(n3372) );
  NAND2_X1 U3428 ( .A1(n3371), .A2(n3372), .ZN(n3370) );
  OAI21_X1 U3429 ( .B1(n2927), .B2(n3727), .A(n3370), .ZN(n3801) );
  NAND2_X1 U3430 ( .A1(n3802), .A2(n3801), .ZN(n3800) );
  NAND2_X1 U3431 ( .A1(n3800), .A2(n2930), .ZN(n3394) );
  INV_X1 U3432 ( .A(n3394), .ZN(n2939) );
  NAND2_X1 U3433 ( .A1(n2917), .A2(REG2_REG_2__SCAN_IN), .ZN(n2936) );
  NAND2_X1 U3434 ( .A1(n2945), .A2(REG3_REG_2__SCAN_IN), .ZN(n2935) );
  NAND2_X1 U3435 ( .A1(n2931), .A2(REG0_REG_2__SCAN_IN), .ZN(n2934) );
  NAND2_X1 U3436 ( .A1(n2932), .A2(REG1_REG_2__SCAN_IN), .ZN(n2933) );
  INV_X2 U3437 ( .A(n2959), .ZN(n3725) );
  OAI22_X1 U3438 ( .A1(n3488), .A2(n3726), .B1(n3725), .B2(n3487), .ZN(n2937)
         );
  XNOR2_X1 U3439 ( .A(n2937), .B(n3727), .ZN(n2940) );
  OAI22_X1 U3440 ( .A1(n3488), .A2(n2951), .B1(n3726), .B2(n3487), .ZN(n2941)
         );
  XNOR2_X1 U3441 ( .A(n2940), .B(n2941), .ZN(n3393) );
  INV_X1 U3442 ( .A(n3393), .ZN(n2938) );
  NAND2_X1 U3443 ( .A1(n2939), .A2(n2938), .ZN(n3395) );
  INV_X1 U3444 ( .A(n2940), .ZN(n2943) );
  INV_X1 U3445 ( .A(n2941), .ZN(n2942) );
  NAND2_X1 U3446 ( .A1(n3040), .A2(REG1_REG_3__SCAN_IN), .ZN(n2949) );
  NAND2_X1 U3447 ( .A1(n3044), .A2(REG0_REG_3__SCAN_IN), .ZN(n2948) );
  NAND2_X1 U3448 ( .A1(n3704), .A2(REG2_REG_3__SCAN_IN), .ZN(n2947) );
  CLKBUF_X3 U3449 ( .A(n2945), .Z(n3685) );
  INV_X1 U3450 ( .A(REG3_REG_3__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U3451 ( .A1(n3685), .A2(n5066), .ZN(n2946) );
  INV_X1 U3452 ( .A(n5048), .ZN(n5057) );
  OAI22_X1 U3453 ( .A1(n3482), .A2(n3726), .B1(n3725), .B2(n5057), .ZN(n2950)
         );
  XNOR2_X1 U3454 ( .A(n2950), .B(n3727), .ZN(n2953) );
  OAI22_X1 U3455 ( .A1(n3482), .A2(n2951), .B1(n3726), .B2(n5057), .ZN(n2952)
         );
  XNOR2_X1 U3456 ( .A(n2953), .B(n2952), .ZN(n3469) );
  OAI22_X1 U3457 ( .A1(n3470), .A2(n3469), .B1(n2953), .B2(n2952), .ZN(n3531)
         );
  NAND2_X1 U34580 ( .A1(n3704), .A2(REG2_REG_4__SCAN_IN), .ZN(n2958) );
  NAND2_X1 U34590 ( .A1(n3040), .A2(REG1_REG_4__SCAN_IN), .ZN(n2957) );
  NOR2_X1 U3460 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2954) );
  NOR2_X1 U3461 ( .A1(n2967), .A2(n2954), .ZN(n3534) );
  NAND2_X1 U3462 ( .A1(n3685), .A2(n3534), .ZN(n2956) );
  NAND2_X1 U3463 ( .A1(n3044), .A2(REG0_REG_4__SCAN_IN), .ZN(n2955) );
  INV_X1 U3464 ( .A(n3493), .ZN(n3536) );
  AOI22_X1 U3465 ( .A1(n5053), .A2(n3253), .B1(n3004), .B2(n3536), .ZN(n2964)
         );
  NAND2_X1 U3466 ( .A1(n5053), .A2(n3004), .ZN(n2961) );
  XOR2_X1 U34670 ( .A(n2964), .B(n2963), .Z(n3533) );
  NOR2_X1 U3468 ( .A1(n3531), .A2(n3533), .ZN(n3532) );
  INV_X1 U34690 ( .A(n2963), .ZN(n2965) );
  NOR2_X1 U3470 ( .A1(n2965), .A2(n2964), .ZN(n2966) );
  NOR2_X1 U34710 ( .A1(n3532), .A2(n2966), .ZN(n3543) );
  NAND2_X1 U3472 ( .A1(n3704), .A2(REG2_REG_5__SCAN_IN), .ZN(n2972) );
  NAND2_X1 U34730 ( .A1(n3040), .A2(REG1_REG_5__SCAN_IN), .ZN(n2971) );
  NAND2_X1 U3474 ( .A1(n2967), .A2(REG3_REG_5__SCAN_IN), .ZN(n2985) );
  OAI21_X1 U34750 ( .B1(n2967), .B2(REG3_REG_5__SCAN_IN), .A(n2985), .ZN(n3549) );
  INV_X1 U3476 ( .A(n3549), .ZN(n2968) );
  NAND2_X1 U34770 ( .A1(n3685), .A2(n2968), .ZN(n2970) );
  NAND2_X1 U3478 ( .A1(n3044), .A2(REG0_REG_5__SCAN_IN), .ZN(n2969) );
  INV_X1 U34790 ( .A(n3545), .ZN(n3522) );
  OAI22_X1 U3480 ( .A1(n3504), .A2(n2951), .B1(n3726), .B2(n3522), .ZN(n2974)
         );
  OAI22_X1 U34810 ( .A1(n3504), .A2(n3726), .B1(n3725), .B2(n3522), .ZN(n2973)
         );
  XNOR2_X1 U3482 ( .A(n2973), .B(n3727), .ZN(n2975) );
  XOR2_X1 U34830 ( .A(n2974), .B(n2975), .Z(n3544) );
  NAND2_X1 U3484 ( .A1(n3543), .A2(n3544), .ZN(n3542) );
  OR2_X1 U34850 ( .A1(n2975), .A2(n2974), .ZN(n2976) );
  NAND2_X1 U3486 ( .A1(n3542), .A2(n2976), .ZN(n3572) );
  NAND2_X1 U34870 ( .A1(n3704), .A2(REG2_REG_6__SCAN_IN), .ZN(n2980) );
  NAND2_X1 U3488 ( .A1(n3040), .A2(REG1_REG_6__SCAN_IN), .ZN(n2979) );
  XNOR2_X1 U34890 ( .A(n2985), .B(REG3_REG_6__SCAN_IN), .ZN(n3508) );
  NAND2_X1 U3490 ( .A1(n3685), .A2(n3508), .ZN(n2978) );
  NAND2_X1 U34910 ( .A1(n3044), .A2(REG0_REG_6__SCAN_IN), .ZN(n2977) );
  NAND4_X1 U3492 ( .A1(n2980), .A2(n2979), .A3(n2978), .A4(n2977), .ZN(n4483)
         );
  INV_X1 U34930 ( .A(n4483), .ZN(n3499) );
  OAI22_X1 U3494 ( .A1(n3499), .A2(n3726), .B1(n3725), .B2(n3501), .ZN(n2981)
         );
  XNOR2_X1 U34950 ( .A(n2981), .B(n3727), .ZN(n3569) );
  OAI22_X1 U3496 ( .A1(n3499), .A2(n2951), .B1(n3726), .B2(n3501), .ZN(n3570)
         );
  NAND2_X1 U34970 ( .A1(n3569), .A2(n3570), .ZN(n2982) );
  NAND2_X1 U3498 ( .A1(n3040), .A2(REG1_REG_7__SCAN_IN), .ZN(n2991) );
  NAND2_X1 U34990 ( .A1(n3704), .A2(REG2_REG_7__SCAN_IN), .ZN(n2990) );
  INV_X1 U3500 ( .A(n2985), .ZN(n2983) );
  AOI21_X1 U35010 ( .B1(n2983), .B2(REG3_REG_6__SCAN_IN), .A(
        REG3_REG_7__SCAN_IN), .ZN(n2986) );
  NAND2_X1 U3502 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n2984) );
  NOR2_X1 U35030 ( .A1(n2985), .A2(n2984), .ZN(n2997) );
  OR2_X1 U3504 ( .A1(n2986), .A2(n2997), .ZN(n3748) );
  INV_X1 U35050 ( .A(n3748), .ZN(n2987) );
  NAND2_X1 U35060 ( .A1(n3685), .A2(n2987), .ZN(n2989) );
  NAND2_X1 U35070 ( .A1(n3044), .A2(REG0_REG_7__SCAN_IN), .ZN(n2988) );
  OR2_X1 U35080 ( .A1(n3596), .A2(n2951), .ZN(n2993) );
  NAND2_X1 U35090 ( .A1(n3745), .A2(n3004), .ZN(n2992) );
  NAND2_X1 U35100 ( .A1(n2993), .A2(n2992), .ZN(n2996) );
  OAI22_X1 U35110 ( .A1(n3596), .A2(n3726), .B1(n3725), .B2(n3554), .ZN(n2994)
         );
  XNOR2_X1 U35120 ( .A(n2994), .B(n3727), .ZN(n2995) );
  XOR2_X1 U35130 ( .A(n2996), .B(n2995), .Z(n3743) );
  NAND2_X1 U35140 ( .A1(n3040), .A2(REG1_REG_8__SCAN_IN), .ZN(n3003) );
  NAND2_X1 U35150 ( .A1(n3044), .A2(REG0_REG_8__SCAN_IN), .ZN(n3002) );
  NOR2_X1 U35160 ( .A1(n2997), .A2(REG3_REG_8__SCAN_IN), .ZN(n2998) );
  OR2_X1 U35170 ( .A1(n3012), .A2(n2998), .ZN(n3799) );
  INV_X1 U35180 ( .A(n3799), .ZN(n2999) );
  NAND2_X1 U35190 ( .A1(n3685), .A2(n2999), .ZN(n3001) );
  NAND2_X1 U35200 ( .A1(n3704), .A2(REG2_REG_8__SCAN_IN), .ZN(n3000) );
  NAND4_X1 U35210 ( .A1(n3003), .A2(n3002), .A3(n3001), .A4(n3000), .ZN(n4480)
         );
  NAND2_X1 U35220 ( .A1(n4480), .A2(n3004), .ZN(n3006) );
  OR2_X1 U35230 ( .A1(n3613), .A2(n3725), .ZN(n3005) );
  NAND2_X1 U35240 ( .A1(n3006), .A2(n3005), .ZN(n3007) );
  XNOR2_X1 U35250 ( .A(n3007), .B(n3250), .ZN(n3009) );
  INV_X1 U35260 ( .A(n3613), .ZN(n3796) );
  AOI22_X1 U35270 ( .A1(n4480), .A2(n3253), .B1(n3004), .B2(n3796), .ZN(n3008)
         );
  NAND2_X1 U35280 ( .A1(n3009), .A2(n3008), .ZN(n3011) );
  OAI21_X1 U35290 ( .B1(n3009), .B2(n3008), .A(n3011), .ZN(n3010) );
  INV_X1 U35300 ( .A(n3010), .ZN(n3788) );
  NAND2_X1 U35310 ( .A1(n3787), .A2(n3011), .ZN(n4266) );
  NOR2_X1 U35320 ( .A1(n3012), .A2(REG3_REG_9__SCAN_IN), .ZN(n3013) );
  OR2_X1 U35330 ( .A1(n3022), .A2(n3013), .ZN(n5132) );
  INV_X1 U35340 ( .A(n5132), .ZN(n3014) );
  NAND2_X1 U35350 ( .A1(n3685), .A2(n3014), .ZN(n3018) );
  NAND2_X1 U35360 ( .A1(n3040), .A2(REG1_REG_9__SCAN_IN), .ZN(n3017) );
  NAND2_X1 U35370 ( .A1(n3044), .A2(REG0_REG_9__SCAN_IN), .ZN(n3016) );
  NAND2_X1 U35380 ( .A1(n3704), .A2(REG2_REG_9__SCAN_IN), .ZN(n3015) );
  NAND4_X1 U35390 ( .A1(n3018), .A2(n3017), .A3(n3016), .A4(n3015), .ZN(n4479)
         );
  INV_X1 U35400 ( .A(n4479), .ZN(n3612) );
  OAI22_X1 U35410 ( .A1(n3612), .A2(n2951), .B1(n3726), .B2(n5105), .ZN(n3032)
         );
  NAND2_X1 U35420 ( .A1(n4479), .A2(n3004), .ZN(n3020) );
  OR2_X1 U35430 ( .A1(n5105), .A2(n3725), .ZN(n3019) );
  NAND2_X1 U35440 ( .A1(n3020), .A2(n3019), .ZN(n3021) );
  XNOR2_X1 U35450 ( .A(n3021), .B(n3727), .ZN(n3031) );
  XOR2_X1 U35460 ( .A(n3032), .B(n3031), .Z(n4267) );
  NAND2_X1 U35470 ( .A1(n4266), .A2(n4267), .ZN(n3775) );
  NAND2_X1 U35480 ( .A1(n3704), .A2(REG2_REG_10__SCAN_IN), .ZN(n3027) );
  NAND2_X1 U35490 ( .A1(n3040), .A2(REG1_REG_10__SCAN_IN), .ZN(n3026) );
  NAND2_X1 U35500 ( .A1(n3022), .A2(REG3_REG_10__SCAN_IN), .ZN(n3042) );
  OR2_X1 U35510 ( .A1(n3022), .A2(REG3_REG_10__SCAN_IN), .ZN(n3023) );
  AND2_X1 U35520 ( .A1(n3042), .A2(n3023), .ZN(n3621) );
  NAND2_X1 U35530 ( .A1(n3685), .A2(n3621), .ZN(n3025) );
  NAND2_X1 U35540 ( .A1(n3044), .A2(REG0_REG_10__SCAN_IN), .ZN(n3024) );
  OR2_X1 U35550 ( .A1(n5108), .A2(n2951), .ZN(n3029) );
  NAND2_X1 U35560 ( .A1(n3782), .A2(n3004), .ZN(n3028) );
  NAND2_X1 U35570 ( .A1(n3029), .A2(n3028), .ZN(n3037) );
  INV_X1 U35580 ( .A(n3782), .ZN(n3626) );
  OAI22_X1 U35590 ( .A1(n5108), .A2(n3726), .B1(n3725), .B2(n3626), .ZN(n3030)
         );
  XNOR2_X1 U35600 ( .A(n3030), .B(n3727), .ZN(n3036) );
  XOR2_X1 U35610 ( .A(n3037), .B(n3036), .Z(n3778) );
  INV_X1 U35620 ( .A(n3031), .ZN(n3034) );
  INV_X1 U35630 ( .A(n3032), .ZN(n3033) );
  NAND2_X1 U35640 ( .A1(n3034), .A2(n3033), .ZN(n3776) );
  INV_X1 U35650 ( .A(n3036), .ZN(n3039) );
  INV_X1 U35660 ( .A(n3037), .ZN(n3038) );
  NAND2_X1 U35670 ( .A1(n3704), .A2(REG2_REG_11__SCAN_IN), .ZN(n3048) );
  NAND2_X1 U35680 ( .A1(n3040), .A2(REG1_REG_11__SCAN_IN), .ZN(n3047) );
  NAND2_X1 U35690 ( .A1(n3042), .A2(n3041), .ZN(n3043) );
  AND2_X1 U35700 ( .A1(n3055), .A2(n3043), .ZN(n4860) );
  NAND2_X1 U35710 ( .A1(n3685), .A2(n4860), .ZN(n3046) );
  NAND2_X1 U35720 ( .A1(n3044), .A2(REG0_REG_11__SCAN_IN), .ZN(n3045) );
  OAI22_X1 U35730 ( .A1(n3809), .A2(n3726), .B1(n3725), .B2(n4858), .ZN(n3049)
         );
  XNOR2_X1 U35740 ( .A(n3049), .B(n3250), .ZN(n3053) );
  OR2_X1 U35750 ( .A1(n3809), .A2(n2951), .ZN(n3051) );
  NAND2_X1 U35760 ( .A1(n4846), .A2(n3004), .ZN(n3050) );
  AND2_X1 U35770 ( .A1(n3051), .A2(n3050), .ZN(n3052) );
  NAND2_X1 U35780 ( .A1(n3053), .A2(n3052), .ZN(n3817) );
  OAI21_X1 U35790 ( .B1(n3053), .B2(n3052), .A(n3817), .ZN(n4297) );
  INV_X1 U35800 ( .A(n4297), .ZN(n3054) );
  NAND2_X1 U35810 ( .A1(n3814), .A2(n3817), .ZN(n3068) );
  NAND2_X1 U3582 ( .A1(n3704), .A2(REG2_REG_12__SCAN_IN), .ZN(n3059) );
  NAND2_X1 U3583 ( .A1(n3040), .A2(REG1_REG_12__SCAN_IN), .ZN(n3058) );
  AOI21_X1 U3584 ( .B1(n3055), .B2(n3586), .A(n3070), .ZN(n4834) );
  NAND2_X1 U3585 ( .A1(n3685), .A2(n4834), .ZN(n3057) );
  NAND2_X1 U3586 ( .A1(n3044), .A2(REG0_REG_12__SCAN_IN), .ZN(n3056) );
  OAI22_X1 U3587 ( .A1(n4849), .A2(n3726), .B1(n3725), .B2(n4832), .ZN(n3060)
         );
  XNOR2_X1 U3588 ( .A(n3060), .B(n3250), .ZN(n3063) );
  OR2_X1 U3589 ( .A1(n4849), .A2(n2951), .ZN(n3062) );
  NAND2_X1 U3590 ( .A1(n4829), .A2(n3004), .ZN(n3061) );
  AND2_X1 U3591 ( .A1(n3062), .A2(n3061), .ZN(n3064) );
  NAND2_X1 U3592 ( .A1(n3063), .A2(n3064), .ZN(n3069) );
  INV_X1 U3593 ( .A(n3063), .ZN(n3066) );
  INV_X1 U3594 ( .A(n3064), .ZN(n3065) );
  NAND2_X1 U3595 ( .A1(n3066), .A2(n3065), .ZN(n3067) );
  AND2_X1 U3596 ( .A1(n3069), .A2(n3067), .ZN(n3815) );
  NAND2_X1 U3597 ( .A1(n3819), .A2(n3069), .ZN(n4275) );
  NAND2_X1 U3598 ( .A1(n3070), .A2(REG3_REG_13__SCAN_IN), .ZN(n3083) );
  OAI21_X1 U3599 ( .B1(n3070), .B2(REG3_REG_13__SCAN_IN), .A(n3083), .ZN(n4280) );
  INV_X1 U3600 ( .A(n4280), .ZN(n5179) );
  NAND2_X1 U3601 ( .A1(n3685), .A2(n5179), .ZN(n3074) );
  NAND2_X1 U3602 ( .A1(n3040), .A2(REG1_REG_13__SCAN_IN), .ZN(n3073) );
  NAND2_X1 U3603 ( .A1(n3044), .A2(REG0_REG_13__SCAN_IN), .ZN(n3072) );
  NAND2_X1 U3604 ( .A1(n3704), .A2(REG2_REG_13__SCAN_IN), .ZN(n3071) );
  NAND4_X1 U3605 ( .A1(n3074), .A2(n3073), .A3(n3072), .A4(n3071), .ZN(n4475)
         );
  INV_X1 U3606 ( .A(n4475), .ZN(n3660) );
  OAI22_X1 U3607 ( .A1(n3660), .A2(n2951), .B1(n3726), .B2(n5160), .ZN(n3079)
         );
  NAND2_X1 U3608 ( .A1(n4475), .A2(n3004), .ZN(n3076) );
  OR2_X1 U3609 ( .A1(n5160), .A2(n3725), .ZN(n3075) );
  NAND2_X1 U3610 ( .A1(n3076), .A2(n3075), .ZN(n3077) );
  XNOR2_X1 U3611 ( .A(n3077), .B(n3727), .ZN(n3078) );
  XOR2_X1 U3612 ( .A(n3079), .B(n3078), .Z(n4276) );
  INV_X1 U3613 ( .A(n3078), .ZN(n3081) );
  INV_X1 U3614 ( .A(n3079), .ZN(n3080) );
  NAND2_X1 U3615 ( .A1(n3081), .A2(n3080), .ZN(n3082) );
  NAND2_X1 U3616 ( .A1(n3040), .A2(REG1_REG_14__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U3617 ( .A1(n3704), .A2(REG2_REG_14__SCAN_IN), .ZN(n3086) );
  NAND2_X1 U3618 ( .A1(n3044), .A2(REG0_REG_14__SCAN_IN), .ZN(n3085) );
  AOI21_X1 U3619 ( .B1(n3083), .B2(n4514), .A(n3092), .ZN(n4820) );
  NAND2_X1 U3620 ( .A1(n3685), .A2(n4820), .ZN(n3084) );
  OAI22_X1 U3621 ( .A1(n4792), .A2(n3726), .B1(n3725), .B2(n4818), .ZN(n3088)
         );
  XNOR2_X1 U3622 ( .A(n3088), .B(n3250), .ZN(n3091) );
  INV_X1 U3623 ( .A(n4792), .ZN(n4474) );
  NOR2_X1 U3624 ( .A1(n4818), .A2(n3726), .ZN(n3089) );
  AOI21_X1 U3625 ( .B1(n4474), .B2(n3253), .A(n3089), .ZN(n3090) );
  AND2_X1 U3626 ( .A1(n3091), .A2(n3090), .ZN(n3752) );
  NAND2_X1 U3627 ( .A1(n2932), .A2(REG1_REG_15__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U3628 ( .A1(n2931), .A2(REG0_REG_15__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U3629 ( .A1(n3704), .A2(REG2_REG_15__SCAN_IN), .ZN(n3095) );
  NAND2_X1 U3630 ( .A1(n3092), .A2(REG3_REG_15__SCAN_IN), .ZN(n3101) );
  OAI21_X1 U3631 ( .B1(n3092), .B2(REG3_REG_15__SCAN_IN), .A(n3101), .ZN(n5197) );
  INV_X1 U3632 ( .A(n5197), .ZN(n3093) );
  NAND2_X1 U3633 ( .A1(n3685), .A2(n3093), .ZN(n3094) );
  OAI22_X1 U3634 ( .A1(n4774), .A2(n3726), .B1(n3725), .B2(n4796), .ZN(n3098)
         );
  XNOR2_X1 U3635 ( .A(n3098), .B(n3250), .ZN(n5191) );
  OR2_X1 U3636 ( .A1(n4774), .A2(n2951), .ZN(n3100) );
  OR2_X1 U3637 ( .A1(n4796), .A2(n3726), .ZN(n3099) );
  NAND2_X1 U3638 ( .A1(n3704), .A2(REG2_REG_16__SCAN_IN), .ZN(n3105) );
  NAND2_X1 U3639 ( .A1(n3040), .A2(REG1_REG_16__SCAN_IN), .ZN(n3104) );
  AOI21_X1 U3640 ( .B1(n3101), .B2(n3840), .A(n3113), .ZN(n4785) );
  NAND2_X1 U3641 ( .A1(n3685), .A2(n4785), .ZN(n3103) );
  NAND2_X1 U3642 ( .A1(n2931), .A2(REG0_REG_16__SCAN_IN), .ZN(n3102) );
  NAND4_X1 U3643 ( .A1(n3105), .A2(n3104), .A3(n3103), .A4(n3102), .ZN(n4756)
         );
  NAND2_X1 U3644 ( .A1(n4756), .A2(n3004), .ZN(n3107) );
  OR2_X1 U3645 ( .A1(n4779), .A2(n3725), .ZN(n3106) );
  NAND2_X1 U3646 ( .A1(n3107), .A2(n3106), .ZN(n3108) );
  XNOR2_X1 U3647 ( .A(n3108), .B(n3250), .ZN(n3110) );
  INV_X1 U3648 ( .A(n4779), .ZN(n3631) );
  AOI22_X1 U3649 ( .A1(n4756), .A2(n3253), .B1(n3004), .B2(n3631), .ZN(n3109)
         );
  OR2_X1 U3650 ( .A1(n3110), .A2(n3109), .ZN(n3832) );
  OAI21_X1 U3651 ( .B1(n5191), .B2(n5190), .A(n3832), .ZN(n3112) );
  NAND2_X1 U3652 ( .A1(n3110), .A2(n3109), .ZN(n3849) );
  NAND3_X1 U3653 ( .A1(n5191), .A2(n5190), .A3(n3832), .ZN(n3111) );
  NAND2_X1 U3654 ( .A1(n3704), .A2(REG2_REG_17__SCAN_IN), .ZN(n3118) );
  NAND2_X1 U3655 ( .A1(n2932), .A2(REG1_REG_17__SCAN_IN), .ZN(n3117) );
  INV_X1 U3656 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3925) );
  INV_X1 U3657 ( .A(n3113), .ZN(n3114) );
  NAND2_X1 U3658 ( .A1(n3113), .A2(REG3_REG_17__SCAN_IN), .ZN(n3127) );
  INV_X1 U3659 ( .A(n3127), .ZN(n3129) );
  AOI21_X1 U3660 ( .B1(n3925), .B2(n3114), .A(n3129), .ZN(n4763) );
  NAND2_X1 U3661 ( .A1(n3685), .A2(n4763), .ZN(n3116) );
  NAND2_X1 U3662 ( .A1(n2931), .A2(REG0_REG_17__SCAN_IN), .ZN(n3115) );
  INV_X1 U3663 ( .A(n4761), .ZN(n3635) );
  OAI22_X1 U3664 ( .A1(n4775), .A2(n3726), .B1(n3725), .B2(n3635), .ZN(n3119)
         );
  XNOR2_X1 U3665 ( .A(n3119), .B(n3250), .ZN(n3123) );
  OR2_X1 U3666 ( .A1(n4775), .A2(n2951), .ZN(n3121) );
  NAND2_X1 U3667 ( .A1(n4761), .A2(n3004), .ZN(n3120) );
  NAND2_X1 U3668 ( .A1(n3121), .A2(n3120), .ZN(n3124) );
  XNOR2_X1 U3669 ( .A(n3123), .B(n3124), .ZN(n3847) );
  NAND2_X1 U3670 ( .A1(n3122), .A2(n3847), .ZN(n3851) );
  NAND2_X1 U3671 ( .A1(n3851), .A2(n3126), .ZN(n5222) );
  NAND2_X1 U3672 ( .A1(n3704), .A2(REG2_REG_18__SCAN_IN), .ZN(n3134) );
  NAND2_X1 U3673 ( .A1(n2932), .A2(REG1_REG_18__SCAN_IN), .ZN(n3133) );
  INV_X1 U3674 ( .A(n3140), .ZN(n3128) );
  OAI21_X1 U3675 ( .B1(REG3_REG_18__SCAN_IN), .B2(n3129), .A(n3128), .ZN(n5232) );
  INV_X1 U3676 ( .A(n5232), .ZN(n3130) );
  NAND2_X1 U3677 ( .A1(n3685), .A2(n3130), .ZN(n3132) );
  NAND2_X1 U3678 ( .A1(n2931), .A2(REG0_REG_18__SCAN_IN), .ZN(n3131) );
  NAND4_X1 U3679 ( .A1(n3134), .A2(n3133), .A3(n3132), .A4(n3131), .ZN(n4724)
         );
  NAND2_X1 U3680 ( .A1(n4724), .A2(n3004), .ZN(n3136) );
  OR2_X1 U3681 ( .A1(n4747), .A2(n3725), .ZN(n3135) );
  NAND2_X1 U3682 ( .A1(n3136), .A2(n3135), .ZN(n3137) );
  XNOR2_X1 U3683 ( .A(n3137), .B(n3250), .ZN(n3139) );
  AOI22_X1 U3684 ( .A1(n4724), .A2(n3253), .B1(n3004), .B2(n5227), .ZN(n3138)
         );
  OR2_X1 U3685 ( .A1(n3139), .A2(n3138), .ZN(n5221) );
  NAND2_X1 U3686 ( .A1(n3139), .A2(n3138), .ZN(n5225) );
  NAND2_X1 U3687 ( .A1(n3140), .A2(REG3_REG_19__SCAN_IN), .ZN(n3150) );
  OAI21_X1 U3688 ( .B1(REG3_REG_19__SCAN_IN), .B2(n3140), .A(n3150), .ZN(n5250) );
  INV_X1 U3689 ( .A(n5250), .ZN(n4731) );
  NAND2_X1 U3690 ( .A1(n3685), .A2(n4731), .ZN(n3144) );
  NAND2_X1 U3691 ( .A1(n3040), .A2(REG1_REG_19__SCAN_IN), .ZN(n3143) );
  NAND2_X1 U3692 ( .A1(n3044), .A2(REG0_REG_19__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U3693 ( .A1(n3704), .A2(REG2_REG_19__SCAN_IN), .ZN(n3141) );
  NAND4_X1 U3694 ( .A1(n3144), .A2(n3143), .A3(n3142), .A4(n3141), .ZN(n5265)
         );
  INV_X1 U3695 ( .A(n5265), .ZN(n5287) );
  OAI22_X1 U3696 ( .A1(n5287), .A2(n2951), .B1(n3726), .B2(n4729), .ZN(n3148)
         );
  NAND2_X1 U3697 ( .A1(n5265), .A2(n3004), .ZN(n3146) );
  OR2_X1 U3698 ( .A1(n4729), .A2(n3725), .ZN(n3145) );
  NAND2_X1 U3699 ( .A1(n3146), .A2(n3145), .ZN(n3147) );
  XNOR2_X1 U3700 ( .A(n3147), .B(n3727), .ZN(n3149) );
  XOR2_X1 U3701 ( .A(n3148), .B(n3149), .Z(n5245) );
  NAND2_X1 U3702 ( .A1(n2932), .A2(REG1_REG_20__SCAN_IN), .ZN(n3156) );
  NAND2_X1 U3703 ( .A1(n2931), .A2(REG0_REG_20__SCAN_IN), .ZN(n3155) );
  OAI21_X1 U3704 ( .B1(REG3_REG_20__SCAN_IN), .B2(n3151), .A(n3178), .ZN(n5301) );
  INV_X1 U3705 ( .A(n5301), .ZN(n3152) );
  NAND2_X1 U3706 ( .A1(n3685), .A2(n3152), .ZN(n3154) );
  NAND2_X1 U3707 ( .A1(n3704), .A2(REG2_REG_20__SCAN_IN), .ZN(n3153) );
  NAND4_X1 U3708 ( .A1(n3156), .A2(n3155), .A3(n3154), .A4(n3153), .ZN(n5312)
         );
  NAND2_X1 U3709 ( .A1(n5312), .A2(n3004), .ZN(n3158) );
  OR2_X1 U3710 ( .A1(n5276), .A2(n3725), .ZN(n3157) );
  NAND2_X1 U3711 ( .A1(n3158), .A2(n3157), .ZN(n3159) );
  XNOR2_X1 U3712 ( .A(n3159), .B(n3250), .ZN(n3162) );
  NOR2_X1 U3713 ( .A1(n5276), .A2(n3726), .ZN(n3160) );
  AOI21_X1 U3714 ( .B1(n5312), .B2(n3253), .A(n3160), .ZN(n3161) );
  OR2_X1 U3715 ( .A1(n3162), .A2(n3161), .ZN(n5260) );
  AND2_X1 U3716 ( .A1(n3162), .A2(n3161), .ZN(n5261) );
  INV_X1 U3717 ( .A(REG3_REG_21__SCAN_IN), .ZN(n5313) );
  XNOR2_X1 U3718 ( .A(n3178), .B(n5313), .ZN(n5325) );
  INV_X1 U3719 ( .A(n5325), .ZN(n4714) );
  NAND2_X1 U3720 ( .A1(n3685), .A2(n4714), .ZN(n3166) );
  NAND2_X1 U3721 ( .A1(n2932), .A2(REG1_REG_21__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U3722 ( .A1(n2931), .A2(REG0_REG_21__SCAN_IN), .ZN(n3164) );
  NAND2_X1 U3723 ( .A1(n3704), .A2(REG2_REG_21__SCAN_IN), .ZN(n3163) );
  NAND4_X1 U3724 ( .A1(n3166), .A2(n3165), .A3(n3164), .A4(n3163), .ZN(n5284)
         );
  NAND2_X1 U3725 ( .A1(n5284), .A2(n3004), .ZN(n3168) );
  OR2_X1 U3726 ( .A1(n5318), .A2(n3725), .ZN(n3167) );
  NAND2_X1 U3727 ( .A1(n3168), .A2(n3167), .ZN(n3169) );
  XNOR2_X1 U3728 ( .A(n3169), .B(n3250), .ZN(n3171) );
  NOR2_X1 U3729 ( .A1(n5318), .A2(n3726), .ZN(n3170) );
  AOI21_X1 U3730 ( .B1(n5284), .B2(n3253), .A(n3170), .ZN(n3172) );
  NAND2_X1 U3731 ( .A1(n3171), .A2(n3172), .ZN(n5309) );
  NAND2_X1 U3732 ( .A1(n5308), .A2(n5309), .ZN(n3175) );
  INV_X1 U3733 ( .A(n3171), .ZN(n3174) );
  INV_X1 U3734 ( .A(n3172), .ZN(n3173) );
  NAND2_X1 U3735 ( .A1(n3174), .A2(n3173), .ZN(n5310) );
  NAND2_X1 U3736 ( .A1(n3175), .A2(n5310), .ZN(n4285) );
  INV_X1 U3737 ( .A(n4285), .ZN(n3186) );
  NAND2_X1 U3738 ( .A1(n3704), .A2(REG2_REG_22__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U3739 ( .A1(n2932), .A2(REG1_REG_22__SCAN_IN), .ZN(n3182) );
  INV_X1 U3740 ( .A(n3178), .ZN(n3176) );
  AOI21_X1 U3741 ( .B1(n3176), .B2(REG3_REG_21__SCAN_IN), .A(
        REG3_REG_22__SCAN_IN), .ZN(n3179) );
  NAND2_X1 U3742 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n3177) );
  OR2_X1 U3743 ( .A1(n3179), .A2(n3187), .ZN(n4695) );
  INV_X1 U3744 ( .A(n4695), .ZN(n4293) );
  NAND2_X1 U3745 ( .A1(n3685), .A2(n4293), .ZN(n3181) );
  NAND2_X1 U3746 ( .A1(n2931), .A2(REG0_REG_22__SCAN_IN), .ZN(n3180) );
  INV_X1 U3747 ( .A(n4694), .ZN(n4290) );
  OAI22_X1 U3748 ( .A1(n5316), .A2(n3726), .B1(n3725), .B2(n4290), .ZN(n3184)
         );
  XNOR2_X1 U3749 ( .A(n3184), .B(n3727), .ZN(n3197) );
  OAI22_X1 U3750 ( .A1(n5316), .A2(n2951), .B1(n3726), .B2(n4290), .ZN(n3196)
         );
  XNOR2_X1 U3751 ( .A(n3197), .B(n3196), .ZN(n4287) );
  NAND2_X1 U3752 ( .A1(n3186), .A2(n3185), .ZN(n3764) );
  NAND2_X1 U3753 ( .A1(n3704), .A2(REG2_REG_23__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U3754 ( .A1(n3040), .A2(REG1_REG_23__SCAN_IN), .ZN(n3191) );
  NAND2_X1 U3755 ( .A1(n3187), .A2(REG3_REG_23__SCAN_IN), .ZN(n3199) );
  OR2_X1 U3756 ( .A1(n3187), .A2(REG3_REG_23__SCAN_IN), .ZN(n3188) );
  AND2_X1 U3757 ( .A1(n3199), .A2(n3188), .ZN(n3770) );
  NAND2_X1 U3758 ( .A1(n3685), .A2(n3770), .ZN(n3190) );
  NAND2_X1 U3759 ( .A1(n3044), .A2(REG0_REG_23__SCAN_IN), .ZN(n3189) );
  OAI22_X1 U3760 ( .A1(n4692), .A2(n3726), .B1(n3725), .B2(n4671), .ZN(n3193)
         );
  XNOR2_X1 U3761 ( .A(n3193), .B(n3727), .ZN(n3209) );
  OR2_X1 U3762 ( .A1(n4692), .A2(n2951), .ZN(n3195) );
  NAND2_X1 U3763 ( .A1(n3769), .A2(n3004), .ZN(n3194) );
  NAND2_X1 U3764 ( .A1(n3195), .A2(n3194), .ZN(n3208) );
  XNOR2_X1 U3765 ( .A(n3209), .B(n3208), .ZN(n3765) );
  NOR2_X1 U3766 ( .A1(n3197), .A2(n3196), .ZN(n3766) );
  NOR2_X1 U3767 ( .A1(n3765), .A2(n3766), .ZN(n3198) );
  NAND2_X1 U3768 ( .A1(n3040), .A2(REG1_REG_24__SCAN_IN), .ZN(n3204) );
  NAND2_X1 U3769 ( .A1(n3044), .A2(REG0_REG_24__SCAN_IN), .ZN(n3203) );
  NAND2_X1 U3770 ( .A1(n3199), .A2(n4258), .ZN(n3200) );
  AND2_X1 U3771 ( .A1(n3213), .A2(n3200), .ZN(n4657) );
  NAND2_X1 U3772 ( .A1(n3685), .A2(n4657), .ZN(n3202) );
  NAND2_X1 U3773 ( .A1(n3704), .A2(REG2_REG_24__SCAN_IN), .ZN(n3201) );
  NAND4_X1 U3774 ( .A1(n3204), .A2(n3203), .A3(n3202), .A4(n3201), .ZN(n4668)
         );
  NAND2_X1 U3775 ( .A1(n4668), .A2(n3004), .ZN(n3206) );
  OR2_X1 U3776 ( .A1(n4656), .A2(n3725), .ZN(n3205) );
  NAND2_X1 U3777 ( .A1(n3206), .A2(n3205), .ZN(n3207) );
  XNOR2_X1 U3778 ( .A(n3207), .B(n3250), .ZN(n3211) );
  NAND2_X1 U3779 ( .A1(n3209), .A2(n3208), .ZN(n3210) );
  INV_X1 U3780 ( .A(n4668), .ZN(n3827) );
  INV_X1 U3781 ( .A(n3211), .ZN(n3212) );
  INV_X1 U3782 ( .A(n3823), .ZN(n3225) );
  NAND2_X1 U3783 ( .A1(n3040), .A2(REG1_REG_25__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U3784 ( .A1(n3044), .A2(REG0_REG_25__SCAN_IN), .ZN(n3217) );
  INV_X1 U3785 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3918) );
  NAND2_X1 U3786 ( .A1(n3213), .A2(n3918), .ZN(n3214) );
  AND2_X1 U3787 ( .A1(n3227), .A2(n3214), .ZN(n4640) );
  NAND2_X1 U3788 ( .A1(n3685), .A2(n4640), .ZN(n3216) );
  NAND2_X1 U3789 ( .A1(n3704), .A2(REG2_REG_25__SCAN_IN), .ZN(n3215) );
  INV_X1 U3790 ( .A(n4632), .ZN(n4638) );
  OAI22_X1 U3791 ( .A1(n4651), .A2(n3726), .B1(n3725), .B2(n4638), .ZN(n3219)
         );
  XNOR2_X1 U3792 ( .A(n3219), .B(n3250), .ZN(n3223) );
  OR2_X1 U3793 ( .A1(n4651), .A2(n2951), .ZN(n3221) );
  NAND2_X1 U3794 ( .A1(n4632), .A2(n3004), .ZN(n3220) );
  AND2_X1 U3795 ( .A1(n3221), .A2(n3220), .ZN(n3222) );
  NAND2_X1 U3796 ( .A1(n3223), .A2(n3222), .ZN(n3226) );
  OAI21_X1 U3797 ( .B1(n3223), .B2(n3222), .A(n3226), .ZN(n3826) );
  INV_X1 U3798 ( .A(n3826), .ZN(n3224) );
  NAND2_X1 U3799 ( .A1(n3704), .A2(REG2_REG_26__SCAN_IN), .ZN(n3232) );
  NAND2_X1 U3800 ( .A1(n3040), .A2(REG1_REG_26__SCAN_IN), .ZN(n3231) );
  INV_X1 U3801 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4310) );
  AND2_X1 U3802 ( .A1(n3227), .A2(n4310), .ZN(n3228) );
  NOR2_X1 U3803 ( .A1(n3241), .A2(n3228), .ZN(n4624) );
  NAND2_X1 U3804 ( .A1(n3685), .A2(n4624), .ZN(n3230) );
  NAND2_X1 U3805 ( .A1(n3044), .A2(REG0_REG_26__SCAN_IN), .ZN(n3229) );
  INV_X1 U3806 ( .A(n4621), .ZN(n3656) );
  OAI22_X1 U3807 ( .A1(n4634), .A2(n3726), .B1(n3725), .B2(n3656), .ZN(n3233)
         );
  XNOR2_X1 U3808 ( .A(n3233), .B(n3250), .ZN(n3236) );
  OR2_X1 U3809 ( .A1(n4634), .A2(n2951), .ZN(n3235) );
  NAND2_X1 U3810 ( .A1(n4621), .A2(n3004), .ZN(n3234) );
  AND2_X1 U3811 ( .A1(n3235), .A2(n3234), .ZN(n3237) );
  AND2_X1 U3812 ( .A1(n3236), .A2(n3237), .ZN(n4306) );
  INV_X1 U3813 ( .A(n3236), .ZN(n3239) );
  INV_X1 U3814 ( .A(n3237), .ZN(n3238) );
  NAND2_X1 U3815 ( .A1(n3239), .A2(n3238), .ZN(n4305) );
  NAND2_X1 U3816 ( .A1(n3240), .A2(n4305), .ZN(n3266) );
  NAND2_X1 U3817 ( .A1(n3040), .A2(REG1_REG_27__SCAN_IN), .ZN(n3247) );
  NAND2_X1 U3818 ( .A1(n3044), .A2(REG0_REG_27__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U3819 ( .A1(n3241), .A2(REG3_REG_27__SCAN_IN), .ZN(n3270) );
  INV_X1 U3820 ( .A(n3241), .ZN(n3242) );
  INV_X1 U3821 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4098) );
  NAND2_X1 U3822 ( .A1(n3242), .A2(n4098), .ZN(n3243) );
  NAND2_X1 U3823 ( .A1(n3685), .A2(n4595), .ZN(n3245) );
  NAND2_X1 U3824 ( .A1(n3704), .A2(REG2_REG_27__SCAN_IN), .ZN(n3244) );
  NAND4_X1 U3825 ( .A1(n3247), .A2(n3246), .A3(n3245), .A4(n3244), .ZN(n4470)
         );
  NAND2_X1 U3826 ( .A1(n4470), .A2(n3004), .ZN(n3249) );
  OR2_X1 U3827 ( .A1(n3657), .A2(n3725), .ZN(n3248) );
  NAND2_X1 U3828 ( .A1(n3249), .A2(n3248), .ZN(n3251) );
  XNOR2_X1 U3829 ( .A(n3251), .B(n3250), .ZN(n3255) );
  NOR2_X1 U3830 ( .A1(n3657), .A2(n3726), .ZN(n3252) );
  AOI21_X1 U3831 ( .B1(n4470), .B2(n3253), .A(n3252), .ZN(n3254) );
  NOR2_X1 U3832 ( .A1(n3255), .A2(n3254), .ZN(n3719) );
  AOI21_X1 U3833 ( .B1(n3255), .B2(n3254), .A(n3719), .ZN(n3265) );
  INV_X1 U3834 ( .A(n3265), .ZN(n3257) );
  OR2_X1 U3835 ( .A1(n4306), .A2(n3257), .ZN(n3256) );
  OR2_X1 U3836 ( .A1(n3257), .A2(n4305), .ZN(n3721) );
  INV_X1 U3837 ( .A(n3259), .ZN(n3432) );
  NAND3_X1 U3838 ( .A1(n3432), .A2(n3261), .A3(n3260), .ZN(n3281) );
  INV_X1 U3839 ( .A(n3269), .ZN(n3263) );
  NAND2_X1 U3840 ( .A1(n5014), .A2(n5173), .ZN(n3262) );
  AND3_X1 U3841 ( .A1(n5327), .A2(n3424), .A3(n3262), .ZN(n3276) );
  OAI211_X1 U3842 ( .C1(n3266), .C2(n3265), .A(n3264), .B(n5322), .ZN(n3287)
         );
  NAND2_X1 U3843 ( .A1(n4462), .A2(n3298), .ZN(n3279) );
  INV_X1 U3844 ( .A(n2869), .ZN(n4981) );
  NOR2_X2 U3845 ( .A1(n3793), .A2(n4981), .ZN(n5258) );
  NAND2_X1 U3846 ( .A1(n3704), .A2(REG2_REG_28__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U3847 ( .A1(n3040), .A2(REG1_REG_28__SCAN_IN), .ZN(n3274) );
  INV_X1 U3848 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3910) );
  OR2_X1 U3849 ( .A1(n3270), .A2(n3910), .ZN(n3684) );
  NAND2_X1 U3850 ( .A1(n3270), .A2(n3910), .ZN(n3271) );
  NAND2_X1 U3851 ( .A1(n3685), .A2(n3733), .ZN(n3273) );
  NAND2_X1 U3852 ( .A1(n3044), .A2(REG0_REG_28__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U3853 ( .A1(n4603), .A2(n5246), .B1(n5258), .B2(n4469), .ZN(n3286)
         );
  NOR2_X2 U3854 ( .A1(n3793), .A2(n2869), .ZN(n5264) );
  AOI22_X1 U3855 ( .A1(n5264), .A2(n4604), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3284) );
  NAND2_X1 U3856 ( .A1(n3281), .A2(n3276), .ZN(n3373) );
  NAND4_X1 U3857 ( .A1(n3373), .A2(n3288), .A3(n3301), .A4(n3277), .ZN(n3278)
         );
  NAND2_X1 U3858 ( .A1(n3278), .A2(STATE_REG_SCAN_IN), .ZN(n3282) );
  OAI21_X1 U3859 ( .B1(n5327), .B2(U3149), .A(n3279), .ZN(n3280) );
  NAND2_X1 U3860 ( .A1(n3281), .A2(n3280), .ZN(n3374) );
  NAND2_X1 U3861 ( .A1(n4301), .A2(n4595), .ZN(n3283) );
  AND2_X1 U3862 ( .A1(n3284), .A2(n3283), .ZN(n3285) );
  NAND3_X1 U3863 ( .A1(n3287), .A2(n3286), .A3(n3285), .ZN(U3211) );
  INV_X1 U3864 ( .A(DATAI_27_), .ZN(n3289) );
  MUX2_X1 U3865 ( .A(n3289), .B(n2870), .S(STATE_REG_SCAN_IN), .Z(n3290) );
  INV_X1 U3866 ( .A(n3290), .ZN(U3325) );
  INV_X1 U3867 ( .A(D_REG_1__SCAN_IN), .ZN(n3973) );
  NOR2_X1 U3868 ( .A1(n4911), .A2(n3293), .ZN(n3296) );
  AOI22_X1 U3869 ( .A1(n4954), .A2(n3973), .B1(n3296), .B2(n3294), .ZN(U3459)
         );
  AOI22_X1 U3870 ( .A1(n4954), .A2(n4173), .B1(n3296), .B2(n3295), .ZN(U3458)
         );
  NAND2_X1 U3871 ( .A1(n4485), .A2(DATAO_REG_31__SCAN_IN), .ZN(n3297) );
  OAI21_X1 U3872 ( .B1(n4453), .B2(n4485), .A(n3297), .ZN(U3581) );
  NAND2_X1 U3873 ( .A1(n3298), .A2(n3301), .ZN(n3299) );
  AND2_X1 U3874 ( .A1(n3300), .A2(n3299), .ZN(n3317) );
  INV_X1 U3875 ( .A(n3317), .ZN(n3303) );
  OR2_X1 U3876 ( .A1(n3301), .A2(U3149), .ZN(n4465) );
  NAND2_X1 U3877 ( .A1(n3302), .A2(n4465), .ZN(n3318) );
  NOR2_X1 U3878 ( .A1(n4998), .A2(n4481), .ZN(U3148) );
  INV_X1 U3879 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3604) );
  INV_X1 U3880 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3509) );
  NAND2_X1 U3881 ( .A1(n4958), .A2(REG2_REG_0__SCAN_IN), .ZN(n4978) );
  INV_X1 U3882 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U3883 ( .A1(n4989), .A2(n3305), .B1(REG2_REG_2__SCAN_IN), .B2(n5039), .ZN(n4988) );
  NAND2_X1 U3884 ( .A1(n4989), .A2(REG2_REG_2__SCAN_IN), .ZN(n3306) );
  INV_X1 U3885 ( .A(REG2_REG_3__SCAN_IN), .ZN(n5069) );
  OAI21_X1 U3886 ( .B1(n3309), .B2(n5002), .A(n3310), .ZN(n5001) );
  INV_X1 U3887 ( .A(REG2_REG_4__SCAN_IN), .ZN(n5000) );
  INV_X1 U3888 ( .A(n3310), .ZN(n3311) );
  INV_X1 U3889 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3312) );
  MUX2_X1 U3890 ( .A(n3312), .B(REG2_REG_5__SCAN_IN), .S(n4928), .Z(n3365) );
  NAND2_X1 U3891 ( .A1(n4926), .A2(REG2_REG_7__SCAN_IN), .ZN(n3315) );
  OAI21_X1 U3892 ( .B1(n4926), .B2(REG2_REG_7__SCAN_IN), .A(n3315), .ZN(n3332)
         );
  XNOR2_X1 U3893 ( .A(n3383), .B(n3384), .ZN(n3320) );
  NOR2_X1 U3894 ( .A1(n3604), .A2(n3320), .ZN(n3385) );
  NAND2_X1 U3895 ( .A1(n3318), .A2(n3317), .ZN(n4966) );
  OR2_X1 U3896 ( .A1(n2869), .A2(n2870), .ZN(n3319) );
  AOI211_X1 U3897 ( .C1(n3604), .C2(n3320), .A(n3385), .B(n4968), .ZN(n3330)
         );
  NAND2_X1 U3898 ( .A1(n4926), .A2(REG1_REG_7__SCAN_IN), .ZN(n3324) );
  INV_X1 U3899 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3321) );
  MUX2_X1 U3900 ( .A(REG1_REG_7__SCAN_IN), .B(n3321), .S(n4926), .Z(n3336) );
  INV_X1 U3901 ( .A(REG1_REG_2__SCAN_IN), .ZN(n5043) );
  MUX2_X1 U3902 ( .A(REG1_REG_2__SCAN_IN), .B(n5043), .S(n4989), .Z(n4993) );
  INV_X1 U3903 ( .A(REG1_REG_1__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U3904 ( .A1(n4993), .A2(n4994), .ZN(n4992) );
  INV_X1 U3905 ( .A(REG1_REG_5__SCAN_IN), .ZN(n5080) );
  MUX2_X1 U3906 ( .A(n5080), .B(REG1_REG_5__SCAN_IN), .S(n4928), .Z(n3360) );
  XNOR2_X1 U3907 ( .A(n3322), .B(n4927), .ZN(n3351) );
  INV_X1 U3908 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3323) );
  OAI22_X1 U3909 ( .A1(n3351), .A2(n3323), .B1(n3322), .B2(n4927), .ZN(n3335)
         );
  NAND2_X1 U3910 ( .A1(n3336), .A2(n3335), .ZN(n3334) );
  NAND2_X1 U3911 ( .A1(n3324), .A2(n3334), .ZN(n3377) );
  XNOR2_X1 U3912 ( .A(n3377), .B(n3383), .ZN(n3325) );
  INV_X1 U3913 ( .A(n2870), .ZN(n4979) );
  NAND2_X1 U3914 ( .A1(REG1_REG_8__SCAN_IN), .A2(n3325), .ZN(n3378) );
  OAI211_X1 U3915 ( .C1(n3325), .C2(REG1_REG_8__SCAN_IN), .A(n5010), .B(n3378), 
        .ZN(n3328) );
  INV_X1 U3916 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3326) );
  NOR2_X1 U3917 ( .A1(n3326), .A2(STATE_REG_SCAN_IN), .ZN(n3791) );
  AOI21_X1 U3918 ( .B1(n4998), .B2(ADDR_REG_8__SCAN_IN), .A(n3791), .ZN(n3327)
         );
  OAI211_X1 U3919 ( .C1(n4591), .C2(n3383), .A(n3328), .B(n3327), .ZN(n3329)
         );
  OR2_X1 U3920 ( .A1(n3330), .A2(n3329), .ZN(U3248) );
  AOI211_X1 U3921 ( .C1(n3333), .C2(n3332), .A(n3331), .B(n4968), .ZN(n3343)
         );
  INV_X1 U3922 ( .A(n4926), .ZN(n3341) );
  OAI211_X1 U3923 ( .C1(n3336), .C2(n3335), .A(n5010), .B(n3334), .ZN(n3340)
         );
  INV_X1 U3924 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3337) );
  NOR2_X1 U3925 ( .A1(STATE_REG_SCAN_IN), .A2(n3337), .ZN(n3338) );
  AOI21_X1 U3926 ( .B1(n4998), .B2(ADDR_REG_7__SCAN_IN), .A(n3338), .ZN(n3339)
         );
  OAI211_X1 U3927 ( .C1(n4591), .C2(n3341), .A(n3340), .B(n3339), .ZN(n3342)
         );
  OR2_X1 U3928 ( .A1(n3343), .A2(n3342), .ZN(U3247) );
  INV_X1 U3929 ( .A(n4591), .ZN(n5003) );
  XOR2_X1 U3930 ( .A(REG1_REG_3__SCAN_IN), .B(n3344), .Z(n3346) );
  NOR2_X1 U3931 ( .A1(STATE_REG_SCAN_IN), .A2(n5066), .ZN(n3472) );
  AOI21_X1 U3932 ( .B1(n4998), .B2(ADDR_REG_3__SCAN_IN), .A(n3472), .ZN(n3345)
         );
  OAI21_X1 U3933 ( .B1(n3346), .B2(n4550), .A(n3345), .ZN(n3349) );
  AOI211_X1 U3934 ( .C1(n5003), .C2(n4929), .A(n3349), .B(n3348), .ZN(n3350)
         );
  INV_X1 U3935 ( .A(n3350), .ZN(U3243) );
  XNOR2_X1 U3936 ( .A(n3351), .B(REG1_REG_6__SCAN_IN), .ZN(n3357) );
  AND2_X1 U3937 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3574) );
  AOI21_X1 U3938 ( .B1(n4998), .B2(ADDR_REG_6__SCAN_IN), .A(n3574), .ZN(n3352)
         );
  OAI21_X1 U3939 ( .B1(n4927), .B2(n4591), .A(n3352), .ZN(n3356) );
  AOI211_X1 U3940 ( .C1(n3509), .C2(n3354), .A(n3353), .B(n4968), .ZN(n3355)
         );
  AOI211_X1 U3941 ( .C1(n5010), .C2(n3357), .A(n3356), .B(n3355), .ZN(n3358)
         );
  INV_X1 U3942 ( .A(n3358), .ZN(U3246) );
  INV_X1 U3943 ( .A(n4928), .ZN(n3369) );
  AOI211_X1 U3944 ( .C1(n3361), .C2(n3360), .A(n3359), .B(n4550), .ZN(n3362)
         );
  INV_X1 U3945 ( .A(n3362), .ZN(n3368) );
  INV_X1 U3946 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3363) );
  NOR2_X1 U3947 ( .A1(STATE_REG_SCAN_IN), .A2(n3363), .ZN(n3546) );
  AOI211_X1 U3948 ( .C1(n2555), .C2(n3365), .A(n3364), .B(n4968), .ZN(n3366)
         );
  AOI211_X1 U3949 ( .C1(n4998), .C2(ADDR_REG_5__SCAN_IN), .A(n3546), .B(n3366), 
        .ZN(n3367) );
  OAI211_X1 U3950 ( .C1(n4591), .C2(n3369), .A(n3368), .B(n3367), .ZN(U3245)
         );
  OAI21_X1 U3951 ( .B1(n3372), .B2(n3371), .A(n3370), .ZN(n4980) );
  NAND3_X1 U3952 ( .A1(n3374), .A2(n3373), .A3(n4462), .ZN(n3803) );
  AOI22_X1 U3953 ( .A1(n5267), .A2(n5015), .B1(n3803), .B2(REG3_REG_0__SCAN_IN), .ZN(n3376) );
  NAND2_X1 U3954 ( .A1(n5258), .A2(n3417), .ZN(n3375) );
  OAI211_X1 U3955 ( .C1(n4980), .C2(n5226), .A(n3376), .B(n3375), .ZN(U3229)
         );
  NAND2_X1 U3956 ( .A1(n4925), .A2(n3377), .ZN(n3379) );
  AND2_X1 U3957 ( .A1(n3379), .A2(n3378), .ZN(n3381) );
  INV_X1 U3958 ( .A(REG1_REG_9__SCAN_IN), .ZN(n5121) );
  MUX2_X1 U3959 ( .A(REG1_REG_9__SCAN_IN), .B(n5121), .S(n3405), .Z(n3380) );
  AOI211_X1 U3960 ( .C1(n3381), .C2(n3380), .A(n4550), .B(n3400), .ZN(n3382)
         );
  INV_X1 U3961 ( .A(n3382), .ZN(n3392) );
  AND2_X1 U3962 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4268) );
  NOR2_X1 U3963 ( .A1(n3384), .A2(n3383), .ZN(n3386) );
  NOR2_X1 U3964 ( .A1(n3386), .A2(n3385), .ZN(n3389) );
  INV_X1 U3965 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3404) );
  MUX2_X1 U3966 ( .A(REG2_REG_9__SCAN_IN), .B(n3404), .S(n3405), .Z(n3388) );
  INV_X1 U3967 ( .A(n3407), .ZN(n3387) );
  AOI211_X1 U3968 ( .C1(n3389), .C2(n3388), .A(n3387), .B(n4968), .ZN(n3390)
         );
  AOI211_X1 U3969 ( .C1(n4998), .C2(ADDR_REG_9__SCAN_IN), .A(n4268), .B(n3390), 
        .ZN(n3391) );
  OAI211_X1 U3970 ( .C1(n4591), .C2(n3405), .A(n3392), .B(n3391), .ZN(U3249)
         );
  INV_X1 U3971 ( .A(n3395), .ZN(n3396) );
  AOI21_X1 U3972 ( .B1(n3393), .B2(n3394), .A(n3396), .ZN(n3399) );
  AOI22_X1 U3973 ( .A1(n5258), .A2(n4486), .B1(n5264), .B2(n3417), .ZN(n3398)
         );
  AOI22_X1 U3974 ( .A1(n5267), .A2(n3416), .B1(n3803), .B2(REG3_REG_2__SCAN_IN), .ZN(n3397) );
  OAI211_X1 U3975 ( .C1(n3399), .C2(n5226), .A(n3398), .B(n3397), .ZN(U3234)
         );
  INV_X1 U3976 ( .A(n3405), .ZN(n4924) );
  XNOR2_X1 U3977 ( .A(n3459), .B(REG1_REG_10__SCAN_IN), .ZN(n3412) );
  INV_X1 U3978 ( .A(n4923), .ZN(n3460) );
  INV_X1 U3979 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3401) );
  NOR2_X1 U3980 ( .A1(STATE_REG_SCAN_IN), .A2(n3401), .ZN(n3402) );
  AOI21_X1 U3981 ( .B1(n4998), .B2(ADDR_REG_10__SCAN_IN), .A(n3402), .ZN(n3403) );
  OAI21_X1 U3982 ( .B1(n3460), .B2(n4591), .A(n3403), .ZN(n3411) );
  OR2_X1 U3983 ( .A1(n3405), .A2(n3404), .ZN(n3406) );
  AOI211_X1 U3984 ( .C1(n3622), .C2(n3409), .A(n3455), .B(n4968), .ZN(n3410)
         );
  AOI211_X1 U3985 ( .C1(n5010), .C2(n3412), .A(n3411), .B(n3410), .ZN(n3413)
         );
  INV_X1 U3986 ( .A(n3413), .ZN(U3250) );
  NAND2_X1 U3987 ( .A1(n4914), .A2(n5173), .ZN(n3415) );
  NAND2_X1 U3988 ( .A1(n4915), .A2(n4916), .ZN(n3414) );
  INV_X1 U3989 ( .A(n3488), .ZN(n3471) );
  NAND2_X1 U3990 ( .A1(n3488), .A2(n3416), .ZN(n5050) );
  INV_X1 U3991 ( .A(n3478), .ZN(n4396) );
  NAND2_X1 U3992 ( .A1(n3439), .A2(n5015), .ZN(n4399) );
  XNOR2_X1 U3993 ( .A(n4396), .B(n3479), .ZN(n3429) );
  AND2_X1 U3994 ( .A1(n3418), .A2(n5015), .ZN(n3440) );
  NAND2_X1 U3995 ( .A1(n3419), .A2(n3440), .ZN(n3442) );
  NAND2_X1 U3996 ( .A1(n3417), .A2(n3804), .ZN(n3420) );
  NAND2_X1 U3997 ( .A1(n3442), .A2(n3420), .ZN(n3422) );
  INV_X1 U3998 ( .A(n3422), .ZN(n3421) );
  NAND2_X1 U3999 ( .A1(n3421), .A2(n4396), .ZN(n3490) );
  NAND2_X1 U4000 ( .A1(n3422), .A2(n3478), .ZN(n3423) );
  NAND2_X1 U4001 ( .A1(n3490), .A2(n3423), .ZN(n3427) );
  INV_X1 U4002 ( .A(n4869), .ZN(n5177) );
  NOR2_X2 U4003 ( .A1(n2869), .A2(n3424), .ZN(n5054) );
  AOI22_X1 U4004 ( .A1(n5283), .A2(n4486), .B1(n3417), .B2(n5054), .ZN(n3425)
         );
  OAI21_X1 U4005 ( .B1(n3487), .B2(n5327), .A(n3425), .ZN(n3426) );
  AOI21_X1 U4006 ( .B1(n3427), .B2(n5177), .A(n3426), .ZN(n3428) );
  OAI21_X1 U4007 ( .B1(n5115), .B2(n3429), .A(n3428), .ZN(n5042) );
  INV_X1 U4008 ( .A(n5042), .ZN(n3438) );
  INV_X1 U4009 ( .A(n3430), .ZN(n3433) );
  NAND3_X1 U4010 ( .A1(n3433), .A2(n3432), .A3(n3431), .ZN(n3434) );
  OAI21_X1 U4011 ( .B1(n2518), .B2(n3487), .A(n5047), .ZN(n5040) );
  AOI22_X1 U4012 ( .A1(n5348), .A2(REG2_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(n5178), .ZN(n3435) );
  OAI21_X1 U4013 ( .B1(n5302), .B2(n5040), .A(n3435), .ZN(n3436) );
  INV_X1 U4014 ( .A(n3436), .ZN(n3437) );
  OAI21_X1 U4015 ( .B1(n3438), .B2(n5348), .A(n3437), .ZN(U3288) );
  INV_X1 U4016 ( .A(n4399), .ZN(n4342) );
  XNOR2_X1 U4017 ( .A(n3419), .B(n4342), .ZN(n3447) );
  OAI22_X1 U4018 ( .A1(n3439), .A2(n5286), .B1(n3488), .B2(n5107), .ZN(n3445)
         );
  OR2_X1 U4019 ( .A1(n3419), .A2(n3440), .ZN(n3441) );
  NAND2_X1 U4020 ( .A1(n3442), .A2(n3441), .ZN(n3443) );
  NOR2_X1 U4021 ( .A1(n3443), .A2(n4869), .ZN(n3444) );
  AOI211_X1 U4022 ( .C1(n5282), .C2(n3804), .A(n3445), .B(n3444), .ZN(n3446)
         );
  OAI21_X1 U4023 ( .B1(n5115), .B2(n3447), .A(n3446), .ZN(n5033) );
  NOR2_X1 U4024 ( .A1(n3448), .A2(n4340), .ZN(n5032) );
  NOR3_X1 U4025 ( .A1(n5302), .A2(n2518), .A3(n5032), .ZN(n3451) );
  AOI22_X1 U4026 ( .A1(n5348), .A2(REG2_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(n5178), .ZN(n3449) );
  INV_X1 U4027 ( .A(n3449), .ZN(n3450) );
  AOI211_X1 U4028 ( .C1(n5033), .C2(n5305), .A(n3451), .B(n3450), .ZN(n3452)
         );
  INV_X1 U4029 ( .A(n3452), .ZN(U3289) );
  NAND2_X1 U4030 ( .A1(n5139), .A2(REG2_REG_11__SCAN_IN), .ZN(n3456) );
  OAI21_X1 U4031 ( .B1(n5139), .B2(REG2_REG_11__SCAN_IN), .A(n3456), .ZN(n3457) );
  AOI211_X1 U4032 ( .C1(n2551), .C2(n3457), .A(n3581), .B(n4968), .ZN(n3468)
         );
  INV_X1 U4033 ( .A(n5139), .ZN(n3466) );
  INV_X1 U4034 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3458) );
  INV_X1 U4035 ( .A(REG1_REG_11__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U4036 ( .A1(n5139), .A2(REG1_REG_11__SCAN_IN), .ZN(n3584) );
  INV_X1 U4037 ( .A(n3584), .ZN(n3461) );
  AOI21_X1 U4038 ( .B1(n5145), .B2(n3466), .A(n3461), .ZN(n3462) );
  OAI211_X1 U4039 ( .C1(n3463), .C2(n3462), .A(n5010), .B(n3583), .ZN(n3465)
         );
  AND2_X1 U4040 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4300) );
  AOI21_X1 U4041 ( .B1(n4998), .B2(ADDR_REG_11__SCAN_IN), .A(n4300), .ZN(n3464) );
  OAI211_X1 U4042 ( .C1(n4591), .C2(n3466), .A(n3465), .B(n3464), .ZN(n3467)
         );
  OR2_X1 U40430 ( .A1(n3468), .A2(n3467), .ZN(U3251) );
  XNOR2_X1 U4044 ( .A(n3470), .B(n3469), .ZN(n3476) );
  AOI22_X1 U4045 ( .A1(n5048), .A2(n5246), .B1(n5264), .B2(n3471), .ZN(n3474)
         );
  AOI21_X1 U4046 ( .B1(n5258), .B2(n5053), .A(n3472), .ZN(n3473) );
  OAI211_X1 U4047 ( .C1(REG3_REG_3__SCAN_IN), .C2(n5326), .A(n3474), .B(n3473), 
        .ZN(n3475) );
  AOI21_X1 U4048 ( .B1(n3476), .B2(n5322), .A(n3475), .ZN(n3477) );
  INV_X1 U4049 ( .A(n3477), .ZN(U3215) );
  NAND2_X1 U4050 ( .A1(n5053), .A2(n3493), .ZN(n4350) );
  NAND2_X1 U4051 ( .A1(n2768), .A2(n4350), .ZN(n4395) );
  NAND2_X1 U4052 ( .A1(n3482), .A2(n5048), .ZN(n4398) );
  AND2_X1 U4053 ( .A1(n4398), .A2(n5050), .ZN(n3480) );
  NAND2_X1 U4054 ( .A1(n4486), .A2(n5057), .ZN(n4397) );
  INV_X1 U4055 ( .A(n3498), .ZN(n3481) );
  XOR2_X1 U4056 ( .A(n4395), .B(n3481), .Z(n3486) );
  NOR2_X1 U4057 ( .A1(n3493), .A2(n5327), .ZN(n3485) );
  OR2_X1 U4058 ( .A1(n3504), .A2(n5107), .ZN(n3484) );
  OR2_X1 U4059 ( .A1(n3482), .A2(n5286), .ZN(n3483) );
  NAND2_X1 U4060 ( .A1(n3484), .A2(n3483), .ZN(n3535) );
  AOI211_X1 U4061 ( .C1(n3486), .C2(n5289), .A(n3485), .B(n3535), .ZN(n5072)
         );
  NAND2_X1 U4062 ( .A1(n3488), .A2(n3487), .ZN(n3489) );
  NAND2_X1 U4063 ( .A1(n3490), .A2(n3489), .ZN(n5059) );
  NOR2_X1 U4064 ( .A1(n4486), .A2(n5048), .ZN(n3492) );
  NAND2_X1 U4065 ( .A1(n4486), .A2(n5048), .ZN(n3491) );
  OAI21_X1 U4066 ( .B1(n5059), .B2(n3492), .A(n3491), .ZN(n3511) );
  XNOR2_X1 U4067 ( .A(n3511), .B(n4395), .ZN(n5073) );
  INV_X1 U4068 ( .A(n5073), .ZN(n3496) );
  OAI211_X1 U4069 ( .C1(n5046), .C2(n3493), .A(n5335), .B(n3525), .ZN(n5071)
         );
  AOI22_X1 U4070 ( .A1(n5348), .A2(REG2_REG_4__SCAN_IN), .B1(n3534), .B2(n5178), .ZN(n3494) );
  OAI21_X1 U4071 ( .B1(n5071), .B2(n4733), .A(n3494), .ZN(n3495) );
  AOI21_X1 U4072 ( .B1(n3496), .B2(n4863), .A(n3495), .ZN(n3497) );
  OAI21_X1 U4073 ( .B1(n5072), .B2(n5348), .A(n3497), .ZN(U3286) );
  AND2_X1 U4074 ( .A1(n4484), .A2(n3522), .ZN(n3517) );
  NAND2_X1 U4075 ( .A1(n3504), .A2(n3545), .ZN(n4328) );
  NAND2_X1 U4076 ( .A1(n3499), .A2(n3573), .ZN(n3592) );
  NAND2_X1 U4077 ( .A1(n4483), .A2(n3501), .ZN(n4348) );
  NAND2_X1 U4078 ( .A1(n3592), .A2(n4348), .ZN(n4401) );
  INV_X1 U4079 ( .A(n4401), .ZN(n3500) );
  XNOR2_X1 U4080 ( .A(n3553), .B(n3500), .ZN(n3506) );
  OR2_X1 U4081 ( .A1(n3596), .A2(n5107), .ZN(n3503) );
  OR2_X1 U4082 ( .A1(n3501), .A2(n5327), .ZN(n3502) );
  OAI211_X1 U4083 ( .C1(n3504), .C2(n5286), .A(n3503), .B(n3502), .ZN(n3505)
         );
  AOI21_X1 U4084 ( .B1(n3506), .B2(n5289), .A(n3505), .ZN(n5087) );
  AND2_X1 U4085 ( .A1(n3523), .A2(n3573), .ZN(n3507) );
  NOR2_X1 U4086 ( .A1(n3560), .A2(n3507), .ZN(n5084) );
  INV_X1 U4087 ( .A(n3508), .ZN(n3577) );
  OAI22_X1 U4088 ( .A1(n5305), .A2(n3509), .B1(n3577), .B2(n5300), .ZN(n3510)
         );
  AOI21_X1 U4089 ( .B1(n5084), .B2(n5344), .A(n3510), .ZN(n3516) );
  NAND2_X1 U4090 ( .A1(n3511), .A2(n4395), .ZN(n3513) );
  NAND2_X1 U4091 ( .A1(n5053), .A2(n3536), .ZN(n3512) );
  NAND2_X1 U4092 ( .A1(n3513), .A2(n3512), .ZN(n3527) );
  AND2_X1 U4093 ( .A1(n4484), .A2(n3545), .ZN(n3514) );
  XNOR2_X1 U4094 ( .A(n3565), .B(n4401), .ZN(n5083) );
  NAND2_X1 U4095 ( .A1(n5083), .A2(n4863), .ZN(n3515) );
  OAI211_X1 U4096 ( .C1(n5087), .C2(n5348), .A(n3516), .B(n3515), .ZN(U3284)
         );
  INV_X1 U4097 ( .A(n3517), .ZN(n4349) );
  NAND2_X1 U4098 ( .A1(n4349), .A2(n4328), .ZN(n4392) );
  XNOR2_X1 U4099 ( .A(n3518), .B(n4392), .ZN(n3519) );
  NAND2_X1 U4100 ( .A1(n3519), .A2(n5289), .ZN(n3521) );
  AOI22_X1 U4101 ( .A1(n5054), .A2(n5053), .B1(n4483), .B2(n5283), .ZN(n3520)
         );
  OAI211_X1 U4102 ( .C1(n5327), .C2(n3522), .A(n3521), .B(n3520), .ZN(n5077)
         );
  INV_X1 U4103 ( .A(n5077), .ZN(n3530) );
  AOI211_X1 U4104 ( .C1(n3545), .C2(n3525), .A(n5291), .B(n3524), .ZN(n5078)
         );
  OAI22_X1 U4105 ( .A1(n5305), .A2(n3312), .B1(n3549), .B2(n5300), .ZN(n3526)
         );
  AOI21_X1 U4106 ( .B1(n5078), .B2(n4838), .A(n3526), .ZN(n3529) );
  XOR2_X1 U4107 ( .A(n4392), .B(n3527), .Z(n5079) );
  NAND2_X1 U4108 ( .A1(n5079), .A2(n4863), .ZN(n3528) );
  OAI211_X1 U4109 ( .C1(n3530), .C2(n5348), .A(n3529), .B(n3528), .ZN(U3285)
         );
  AOI211_X1 U4110 ( .C1(n3533), .C2(n3531), .A(n5226), .B(n3532), .ZN(n3541)
         );
  INV_X1 U4111 ( .A(n3534), .ZN(n3539) );
  AOI22_X1 U4112 ( .A1(n3535), .A2(n5243), .B1(REG3_REG_4__SCAN_IN), .B2(U3149), .ZN(n3538) );
  NAND2_X1 U4113 ( .A1(n5267), .A2(n3536), .ZN(n3537) );
  OAI211_X1 U4114 ( .C1(n5326), .C2(n3539), .A(n3538), .B(n3537), .ZN(n3540)
         );
  OR2_X1 U4115 ( .A1(n3541), .A2(n3540), .ZN(U3227) );
  OAI21_X1 U4116 ( .B1(n3544), .B2(n3543), .A(n3542), .ZN(n3551) );
  AOI22_X1 U4117 ( .A1(n3545), .A2(n5246), .B1(n5264), .B2(n5053), .ZN(n3548)
         );
  AOI21_X1 U4118 ( .B1(n5258), .B2(n4483), .A(n3546), .ZN(n3547) );
  OAI211_X1 U4119 ( .C1(n5326), .C2(n3549), .A(n3548), .B(n3547), .ZN(n3550)
         );
  AOI21_X1 U4120 ( .B1(n3551), .B2(n5322), .A(n3550), .ZN(n3552) );
  INV_X1 U4121 ( .A(n3552), .ZN(U3224) );
  NAND2_X1 U4122 ( .A1(n3593), .A2(n3592), .ZN(n3555) );
  NAND2_X1 U4123 ( .A1(n3596), .A2(n3745), .ZN(n3591) );
  NAND2_X1 U4124 ( .A1(n4482), .A2(n3554), .ZN(n4326) );
  NAND2_X1 U4125 ( .A1(n3591), .A2(n4326), .ZN(n4394) );
  XNOR2_X1 U4126 ( .A(n3555), .B(n4394), .ZN(n3559) );
  NAND2_X1 U4127 ( .A1(n4480), .A2(n5283), .ZN(n3557) );
  NAND2_X1 U4128 ( .A1(n4483), .A2(n5054), .ZN(n3556) );
  NAND2_X1 U4129 ( .A1(n3557), .A2(n3556), .ZN(n3744) );
  AOI21_X1 U4130 ( .B1(n3745), .B2(n5282), .A(n3744), .ZN(n3558) );
  OAI21_X1 U4131 ( .B1(n3559), .B2(n5115), .A(n3558), .ZN(n5090) );
  INV_X1 U4132 ( .A(n5090), .ZN(n3568) );
  INV_X1 U4133 ( .A(n3560), .ZN(n3561) );
  AOI211_X1 U4134 ( .C1(n3745), .C2(n3561), .A(n5291), .B(n3603), .ZN(n5091)
         );
  INV_X1 U4135 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3562) );
  OAI22_X1 U4136 ( .A1(n5305), .A2(n3562), .B1(n3748), .B2(n5300), .ZN(n3563)
         );
  AOI21_X1 U4137 ( .B1(n5091), .B2(n4838), .A(n3563), .ZN(n3567) );
  NOR2_X1 U4138 ( .A1(n4483), .A2(n3573), .ZN(n3564) );
  XOR2_X1 U4139 ( .A(n3601), .B(n4394), .Z(n5092) );
  NAND2_X1 U4140 ( .A1(n5092), .A2(n4863), .ZN(n3566) );
  OAI211_X1 U4141 ( .C1(n3568), .C2(n5348), .A(n3567), .B(n3566), .ZN(U3283)
         );
  XOR2_X1 U4142 ( .A(n3570), .B(n3569), .Z(n3571) );
  XNOR2_X1 U4143 ( .A(n3572), .B(n3571), .ZN(n3579) );
  AOI22_X1 U4144 ( .A1(n3573), .A2(n5246), .B1(n5264), .B2(n4484), .ZN(n3576)
         );
  AOI21_X1 U4145 ( .B1(n5258), .B2(n4482), .A(n3574), .ZN(n3575) );
  OAI211_X1 U4146 ( .C1(n5326), .C2(n3577), .A(n3576), .B(n3575), .ZN(n3578)
         );
  AOI21_X1 U4147 ( .B1(n3579), .B2(n5322), .A(n3578), .ZN(n3580) );
  INV_X1 U4148 ( .A(n3580), .ZN(U3236) );
  INV_X1 U4149 ( .A(REG2_REG_12__SCAN_IN), .ZN(n4836) );
  INV_X1 U4150 ( .A(n4922), .ZN(n4494) );
  AOI211_X1 U4151 ( .C1(n4836), .C2(n3582), .A(n4497), .B(n4968), .ZN(n3590)
         );
  OAI211_X1 U4152 ( .C1(n3585), .C2(REG1_REG_12__SCAN_IN), .A(n5010), .B(n4488), .ZN(n3588) );
  NOR2_X1 U4153 ( .A1(n3586), .A2(STATE_REG_SCAN_IN), .ZN(n3808) );
  AOI21_X1 U4154 ( .B1(n4998), .B2(ADDR_REG_12__SCAN_IN), .A(n3808), .ZN(n3587) );
  OAI211_X1 U4155 ( .C1(n4591), .C2(n4494), .A(n3588), .B(n3587), .ZN(n3589)
         );
  OR2_X1 U4156 ( .A1(n3590), .A2(n3589), .ZN(U3252) );
  AND2_X1 U4157 ( .A1(n3592), .A2(n3591), .ZN(n4353) );
  NAND2_X1 U4158 ( .A1(n3593), .A2(n4353), .ZN(n3594) );
  NAND2_X1 U4159 ( .A1(n3594), .A2(n4326), .ZN(n3614) );
  AND2_X1 U4160 ( .A1(n4480), .A2(n3796), .ZN(n3610) );
  INV_X1 U4161 ( .A(n3610), .ZN(n3595) );
  INV_X1 U4162 ( .A(n4480), .ZN(n5109) );
  NAND2_X1 U4163 ( .A1(n5109), .A2(n3613), .ZN(n3609) );
  XNOR2_X1 U4164 ( .A(n3614), .B(n4421), .ZN(n3600) );
  OR2_X1 U4165 ( .A1(n3596), .A2(n5286), .ZN(n3598) );
  NAND2_X1 U4166 ( .A1(n4479), .A2(n5283), .ZN(n3597) );
  AND2_X1 U4167 ( .A1(n3598), .A2(n3597), .ZN(n3794) );
  OAI21_X1 U4168 ( .B1(n3613), .B2(n5327), .A(n3794), .ZN(n3599) );
  AOI21_X1 U4169 ( .B1(n3600), .B2(n5289), .A(n3599), .ZN(n5095) );
  NAND2_X1 U4170 ( .A1(n4482), .A2(n3745), .ZN(n3602) );
  XOR2_X1 U4171 ( .A(n4421), .B(n3611), .Z(n5098) );
  NAND2_X1 U4172 ( .A1(n5098), .A2(n4863), .ZN(n3608) );
  OAI21_X1 U4173 ( .B1(n3603), .B2(n3613), .A(n5103), .ZN(n5096) );
  INV_X1 U4174 ( .A(n5096), .ZN(n3606) );
  OAI22_X1 U4175 ( .A1(n5305), .A2(n3604), .B1(n3799), .B2(n5300), .ZN(n3605)
         );
  AOI21_X1 U4176 ( .B1(n3606), .B2(n5344), .A(n3605), .ZN(n3607) );
  OAI211_X1 U4177 ( .C1(n5348), .C2(n5095), .A(n3608), .B(n3607), .ZN(U3282)
         );
  NAND2_X1 U4178 ( .A1(n4479), .A2(n5119), .ZN(n4418) );
  NAND2_X1 U4179 ( .A1(n3612), .A2(n5105), .ZN(n4419) );
  NAND2_X1 U4180 ( .A1(n5108), .A2(n3782), .ZN(n4334) );
  INV_X1 U4181 ( .A(n5108), .ZN(n4478) );
  NAND2_X1 U4182 ( .A1(n4478), .A2(n3626), .ZN(n4331) );
  XNOR2_X1 U4183 ( .A(n3627), .B(n4393), .ZN(n5133) );
  AND2_X1 U4184 ( .A1(n4480), .A2(n3613), .ZN(n4325) );
  NAND2_X1 U4185 ( .A1(n5109), .A2(n3796), .ZN(n4355) );
  NOR2_X1 U4186 ( .A1(n4479), .A2(n5105), .ZN(n5111) );
  NAND2_X1 U4187 ( .A1(n4479), .A2(n5105), .ZN(n4358) );
  OAI211_X1 U4188 ( .C1(n3615), .C2(n4393), .A(n3658), .B(n5289), .ZN(n3619)
         );
  OR2_X1 U4189 ( .A1(n3809), .A2(n5107), .ZN(n3617) );
  NAND2_X1 U4190 ( .A1(n4479), .A2(n5054), .ZN(n3616) );
  NAND2_X1 U4191 ( .A1(n3617), .A2(n3616), .ZN(n3780) );
  INV_X1 U4192 ( .A(n3780), .ZN(n3618) );
  OAI211_X1 U4193 ( .C1(n5327), .C2(n3626), .A(n3619), .B(n3618), .ZN(n5135)
         );
  NAND2_X1 U4194 ( .A1(n5135), .A2(n5305), .ZN(n3625) );
  AND2_X1 U4195 ( .A1(n5104), .A2(n3782), .ZN(n3620) );
  NOR2_X1 U4196 ( .A1(n4859), .A2(n3620), .ZN(n5136) );
  INV_X1 U4197 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3622) );
  INV_X1 U4198 ( .A(n3621), .ZN(n3781) );
  OAI22_X1 U4199 ( .A1(n5305), .A2(n3622), .B1(n3781), .B2(n5300), .ZN(n3623)
         );
  AOI21_X1 U4200 ( .B1(n5136), .B2(n5344), .A(n3623), .ZN(n3624) );
  OAI211_X1 U4201 ( .C1(n5133), .C2(n4841), .A(n3625), .B(n3624), .ZN(U3280)
         );
  NAND2_X1 U4202 ( .A1(n3809), .A2(n4846), .ZN(n4320) );
  INV_X1 U4203 ( .A(n3809), .ZN(n4477) );
  NAND2_X1 U4204 ( .A1(n4477), .A2(n4858), .ZN(n4332) );
  NAND2_X1 U4205 ( .A1(n4855), .A2(n4854), .ZN(n4853) );
  NAND2_X1 U4206 ( .A1(n3809), .A2(n4858), .ZN(n3628) );
  NAND2_X1 U4207 ( .A1(n4849), .A2(n4829), .ZN(n4321) );
  INV_X1 U4208 ( .A(n4849), .ZN(n4476) );
  NAND2_X1 U4209 ( .A1(n4476), .A2(n4832), .ZN(n5155) );
  NAND2_X1 U4210 ( .A1(n4321), .A2(n5155), .ZN(n4826) );
  NOR2_X1 U4211 ( .A1(n4475), .A2(n5163), .ZN(n4797) );
  NAND2_X1 U4212 ( .A1(n4475), .A2(n5163), .ZN(n4391) );
  NAND2_X1 U4213 ( .A1(n4792), .A2(n3757), .ZN(n4323) );
  NAND2_X1 U4214 ( .A1(n4474), .A2(n4818), .ZN(n4318) );
  NAND2_X1 U4215 ( .A1(n4792), .A2(n4818), .ZN(n4801) );
  NAND2_X1 U4216 ( .A1(n4774), .A2(n4796), .ZN(n3663) );
  NAND3_X1 U4217 ( .A1(n3629), .A2(n4801), .A3(n3663), .ZN(n3630) );
  INV_X1 U4218 ( .A(n4774), .ZN(n4473) );
  NAND2_X1 U4219 ( .A1(n4473), .A2(n5193), .ZN(n3662) );
  NAND2_X1 U4220 ( .A1(n3630), .A2(n3662), .ZN(n4783) );
  AND2_X1 U4221 ( .A1(n4756), .A2(n4779), .ZN(n4754) );
  NOR2_X1 U4222 ( .A1(n4756), .A2(n4779), .ZN(n4436) );
  NAND2_X1 U4223 ( .A1(n4783), .A2(n4782), .ZN(n4784) );
  NAND2_X1 U4224 ( .A1(n4756), .A2(n3631), .ZN(n3632) );
  NAND2_X1 U4225 ( .A1(n4784), .A2(n3632), .ZN(n4753) );
  INV_X1 U4226 ( .A(n4753), .ZN(n3634) );
  NAND2_X1 U4227 ( .A1(n4775), .A2(n4761), .ZN(n4738) );
  INV_X1 U4228 ( .A(n4775), .ZN(n4472) );
  NAND2_X1 U4229 ( .A1(n4472), .A2(n3635), .ZN(n3665) );
  INV_X1 U4230 ( .A(n4752), .ZN(n3633) );
  NAND2_X1 U4231 ( .A1(n3634), .A2(n3633), .ZN(n3637) );
  NAND2_X1 U4232 ( .A1(n4775), .A2(n3635), .ZN(n3636) );
  NAND2_X1 U4233 ( .A1(n3637), .A2(n3636), .ZN(n4719) );
  INV_X1 U4234 ( .A(n4724), .ZN(n4757) );
  NAND2_X1 U4235 ( .A1(n4757), .A2(n5227), .ZN(n3667) );
  AND2_X1 U4236 ( .A1(n4724), .A2(n4747), .ZN(n4743) );
  INV_X1 U4237 ( .A(n4743), .ZN(n3638) );
  NAND2_X1 U4238 ( .A1(n3667), .A2(n3638), .ZN(n4739) );
  INV_X1 U4239 ( .A(n5276), .ZN(n5281) );
  NOR2_X1 U4240 ( .A1(n5312), .A2(n5281), .ZN(n3645) );
  NAND2_X1 U4241 ( .A1(n5287), .A2(n4729), .ZN(n3644) );
  INV_X1 U4242 ( .A(n3644), .ZN(n3640) );
  NOR2_X1 U4243 ( .A1(n5265), .A2(n4729), .ZN(n3672) );
  INV_X1 U4244 ( .A(n3672), .ZN(n3669) );
  AND2_X1 U4245 ( .A1(n5265), .A2(n4729), .ZN(n3668) );
  INV_X1 U4246 ( .A(n3668), .ZN(n3639) );
  NAND2_X1 U4247 ( .A1(n3669), .A2(n3639), .ZN(n4722) );
  OR2_X1 U4248 ( .A1(n3640), .A2(n4722), .ZN(n5272) );
  OR2_X1 U4249 ( .A1(n3645), .A2(n5272), .ZN(n3643) );
  AND2_X1 U4250 ( .A1(n4739), .A2(n3643), .ZN(n3641) );
  NAND2_X1 U4251 ( .A1(n5312), .A2(n5281), .ZN(n3642) );
  AND2_X1 U4252 ( .A1(n3641), .A2(n3642), .ZN(n3651) );
  INV_X1 U4253 ( .A(n3642), .ZN(n3650) );
  INV_X1 U4254 ( .A(n3643), .ZN(n3648) );
  NAND2_X1 U4255 ( .A1(n4757), .A2(n4747), .ZN(n4720) );
  AND2_X1 U4256 ( .A1(n4720), .A2(n3644), .ZN(n5270) );
  INV_X1 U4257 ( .A(n3645), .ZN(n3646) );
  AND2_X1 U4258 ( .A1(n5270), .A2(n3646), .ZN(n3647) );
  OR2_X1 U4259 ( .A1(n3648), .A2(n3647), .ZN(n3649) );
  AND2_X1 U4260 ( .A1(n5284), .A2(n4711), .ZN(n3652) );
  INV_X1 U4261 ( .A(n5284), .ZN(n4289) );
  NAND2_X1 U4262 ( .A1(n4289), .A2(n5318), .ZN(n3653) );
  NAND2_X1 U4263 ( .A1(n5316), .A2(n4694), .ZN(n4663) );
  NAND2_X1 U4264 ( .A1(n4710), .A2(n4290), .ZN(n3678) );
  NAND2_X1 U4265 ( .A1(n4710), .A2(n4694), .ZN(n3654) );
  NAND2_X1 U4266 ( .A1(n4682), .A2(n3654), .ZN(n4677) );
  INV_X1 U4267 ( .A(n4692), .ZN(n4471) );
  XNOR2_X1 U4268 ( .A(n4471), .B(n4671), .ZN(n4676) );
  NAND2_X1 U4269 ( .A1(n4677), .A2(n4676), .ZN(n4678) );
  NAND2_X1 U4270 ( .A1(n4678), .A2(n2541), .ZN(n4645) );
  NAND2_X1 U4271 ( .A1(n3827), .A2(n4656), .ZN(n3655) );
  INV_X1 U4272 ( .A(n4656), .ZN(n4257) );
  NOR2_X1 U4273 ( .A1(n4616), .A2(n4632), .ZN(n4408) );
  NAND2_X1 U4274 ( .A1(n4616), .A2(n4632), .ZN(n4407) );
  INV_X1 U4275 ( .A(n4470), .ZN(n4618) );
  NAND2_X1 U4276 ( .A1(n4618), .A2(n4603), .ZN(n4383) );
  NAND2_X1 U4277 ( .A1(n4470), .A2(n3657), .ZN(n4375) );
  NAND2_X1 U4278 ( .A1(n4607), .A2(n3734), .ZN(n4382) );
  NAND2_X1 U4279 ( .A1(n4469), .A2(n3724), .ZN(n4374) );
  NAND2_X1 U4280 ( .A1(n4382), .A2(n4374), .ZN(n4410) );
  XNOR2_X1 U4281 ( .A(n3699), .B(n4410), .ZN(n4874) );
  NAND2_X1 U4282 ( .A1(n4845), .A2(n4844), .ZN(n4843) );
  NAND2_X1 U4283 ( .A1(n4475), .A2(n5160), .ZN(n3659) );
  AND2_X1 U4284 ( .A1(n5155), .A2(n3659), .ZN(n4339) );
  NAND2_X1 U4285 ( .A1(n3660), .A2(n5163), .ZN(n4324) );
  NAND2_X1 U4286 ( .A1(n4791), .A2(n3664), .ZN(n4790) );
  OR2_X1 U4287 ( .A1(n4774), .A2(n5193), .ZN(n4319) );
  NAND2_X1 U4288 ( .A1(n4790), .A2(n4319), .ZN(n4771) );
  INV_X1 U4289 ( .A(n4782), .ZN(n4770) );
  INV_X1 U4290 ( .A(n4754), .ZN(n3666) );
  NAND2_X1 U4291 ( .A1(n3666), .A2(n3665), .ZN(n4364) );
  NAND2_X1 U4292 ( .A1(n4738), .A2(n3667), .ZN(n3674) );
  NOR2_X1 U4293 ( .A1(n4743), .A2(n3668), .ZN(n3675) );
  INV_X1 U4294 ( .A(n3675), .ZN(n4366) );
  NOR2_X1 U4295 ( .A1(n5312), .A2(n5276), .ZN(n3673) );
  INV_X1 U4296 ( .A(n3673), .ZN(n3671) );
  AND2_X1 U4297 ( .A1(n5312), .A2(n5276), .ZN(n4365) );
  INV_X1 U4298 ( .A(n4365), .ZN(n3670) );
  AOI211_X1 U4299 ( .C1(n3675), .C2(n3674), .A(n3673), .B(n3672), .ZN(n3676)
         );
  NOR2_X1 U4300 ( .A1(n3676), .A2(n4365), .ZN(n4662) );
  INV_X1 U4301 ( .A(n4663), .ZN(n3677) );
  NOR2_X1 U4302 ( .A1(n5284), .A2(n5318), .ZN(n4415) );
  NOR3_X1 U4303 ( .A1(n4662), .A2(n3677), .A3(n4415), .ZN(n4439) );
  NAND2_X1 U4304 ( .A1(n5284), .A2(n5318), .ZN(n4687) );
  NAND2_X1 U4305 ( .A1(n4687), .A2(n3678), .ZN(n3679) );
  NAND2_X1 U4306 ( .A1(n4663), .A2(n3679), .ZN(n3681) );
  OR2_X1 U4307 ( .A1(n4692), .A2(n3769), .ZN(n3680) );
  NAND2_X1 U4308 ( .A1(n3681), .A2(n3680), .ZN(n4438) );
  NAND2_X1 U4309 ( .A1(n3827), .A2(n4257), .ZN(n4413) );
  NAND2_X1 U4310 ( .A1(n4692), .A2(n3769), .ZN(n4646) );
  NAND2_X1 U4311 ( .A1(n4413), .A2(n4646), .ZN(n4442) );
  AND2_X1 U4312 ( .A1(n4668), .A2(n4656), .ZN(n4369) );
  INV_X1 U4313 ( .A(n4369), .ZN(n4414) );
  NOR2_X1 U4314 ( .A1(n4651), .A2(n4632), .ZN(n4370) );
  NAND2_X1 U4315 ( .A1(n4634), .A2(n4621), .ZN(n4420) );
  NAND2_X1 U4316 ( .A1(n4651), .A2(n4632), .ZN(n4611) );
  NAND2_X1 U4317 ( .A1(n4420), .A2(n4611), .ZN(n4444) );
  OR2_X1 U4318 ( .A1(n4634), .A2(n4621), .ZN(n4600) );
  NAND2_X1 U4319 ( .A1(n4599), .A2(n4600), .ZN(n4446) );
  NAND2_X1 U4320 ( .A1(n3040), .A2(REG1_REG_29__SCAN_IN), .ZN(n3689) );
  NAND2_X1 U4321 ( .A1(n3044), .A2(REG0_REG_29__SCAN_IN), .ZN(n3688) );
  INV_X1 U4322 ( .A(n3684), .ZN(n3714) );
  NAND2_X1 U4323 ( .A1(n3685), .A2(n3714), .ZN(n3687) );
  NAND2_X1 U4324 ( .A1(n3704), .A2(REG2_REG_29__SCAN_IN), .ZN(n3686) );
  NAND4_X1 U4325 ( .A1(n3689), .A2(n3688), .A3(n3687), .A4(n3686), .ZN(n4468)
         );
  NAND2_X1 U4326 ( .A1(n4468), .A2(n5283), .ZN(n3690) );
  OAI21_X1 U4327 ( .B1(n5327), .B2(n3724), .A(n3690), .ZN(n3692) );
  AND2_X1 U4328 ( .A1(n4470), .A2(n5054), .ZN(n3691) );
  INV_X1 U4329 ( .A(n4873), .ZN(n3697) );
  OAI211_X1 U4330 ( .C1(n4594), .C2(n3724), .A(n3712), .B(n5335), .ZN(n4872)
         );
  AOI22_X1 U4331 ( .A1(n5348), .A2(REG2_REG_28__SCAN_IN), .B1(n3733), .B2(
        n5178), .ZN(n3695) );
  OAI21_X1 U4332 ( .B1(n4872), .B2(n4733), .A(n3695), .ZN(n3696) );
  AOI21_X1 U4333 ( .B1(n3697), .B2(n5305), .A(n3696), .ZN(n3698) );
  OAI21_X1 U4334 ( .B1(n4874), .B2(n4841), .A(n3698), .ZN(U3262) );
  AOI22_X1 U4335 ( .A1(n3699), .A2(n4410), .B1(n3734), .B2(n4469), .ZN(n3700)
         );
  XOR2_X1 U4336 ( .A(n4468), .B(n4372), .Z(n4426) );
  XNOR2_X1 U4337 ( .A(n3700), .B(n4426), .ZN(n4871) );
  INV_X1 U4338 ( .A(n4382), .ZN(n3701) );
  NAND2_X1 U4339 ( .A1(n3040), .A2(REG1_REG_30__SCAN_IN), .ZN(n3707) );
  NAND2_X1 U4340 ( .A1(n3704), .A2(REG2_REG_30__SCAN_IN), .ZN(n3706) );
  NAND2_X1 U4341 ( .A1(n3044), .A2(REG0_REG_30__SCAN_IN), .ZN(n3705) );
  AND3_X1 U4342 ( .A1(n3707), .A2(n3706), .A3(n3705), .ZN(n4376) );
  OAI22_X1 U4343 ( .A1(n4376), .A2(n3708), .B1(n5327), .B2(n4372), .ZN(n3709)
         );
  AOI21_X1 U4344 ( .B1(n3712), .B2(n4378), .A(n5291), .ZN(n3713) );
  NAND2_X1 U4345 ( .A1(n3713), .A2(n5331), .ZN(n4870) );
  AOI22_X1 U4346 ( .A1(n5348), .A2(REG2_REG_29__SCAN_IN), .B1(n3714), .B2(
        n5178), .ZN(n3715) );
  OAI21_X1 U4347 ( .B1(n4870), .B2(n4733), .A(n3715), .ZN(n3716) );
  AOI21_X1 U4348 ( .B1(n3711), .B2(n5305), .A(n3716), .ZN(n3717) );
  OAI21_X1 U4349 ( .B1(n4871), .B2(n4841), .A(n3717), .ZN(U3354) );
  INV_X1 U4350 ( .A(n3719), .ZN(n3720) );
  AND2_X1 U4351 ( .A1(n3721), .A2(n3720), .ZN(n3722) );
  NAND2_X1 U4352 ( .A1(n3723), .A2(n3722), .ZN(n3732) );
  OAI22_X1 U4353 ( .A1(n4607), .A2(n2951), .B1(n3726), .B2(n3724), .ZN(n3730)
         );
  OAI22_X1 U4354 ( .A1(n4607), .A2(n3726), .B1(n3725), .B2(n3724), .ZN(n3728)
         );
  XNOR2_X1 U4355 ( .A(n3728), .B(n3727), .ZN(n3729) );
  XNOR2_X1 U4356 ( .A(n3732), .B(n3731), .ZN(n3741) );
  INV_X1 U4357 ( .A(n3733), .ZN(n3738) );
  AOI22_X1 U4358 ( .A1(n3734), .A2(n5246), .B1(n5264), .B2(n4470), .ZN(n3737)
         );
  NOR2_X1 U4359 ( .A1(n3910), .A2(STATE_REG_SCAN_IN), .ZN(n3735) );
  AOI21_X1 U4360 ( .B1(n5258), .B2(n4468), .A(n3735), .ZN(n3736) );
  OAI211_X1 U4361 ( .C1(n5326), .C2(n3738), .A(n3737), .B(n3736), .ZN(n3739)
         );
  INV_X1 U4362 ( .A(n3739), .ZN(n3740) );
  OAI21_X1 U4363 ( .B1(n3741), .B2(n5226), .A(n3740), .ZN(U3217) );
  XOR2_X1 U4364 ( .A(n3743), .B(n3742), .Z(n3750) );
  AOI22_X1 U4365 ( .A1(n3744), .A2(n5243), .B1(REG3_REG_7__SCAN_IN), .B2(U3149), .ZN(n3747) );
  NAND2_X1 U4366 ( .A1(n5246), .A2(n3745), .ZN(n3746) );
  OAI211_X1 U4367 ( .C1(n5326), .C2(n3748), .A(n3747), .B(n3746), .ZN(n3749)
         );
  AOI21_X1 U4368 ( .B1(n3750), .B2(n5322), .A(n3749), .ZN(n3751) );
  INV_X1 U4369 ( .A(n3751), .ZN(U3210) );
  NOR2_X1 U4370 ( .A1(n2553), .A2(n3752), .ZN(n3753) );
  XNOR2_X1 U4371 ( .A(n3754), .B(n3753), .ZN(n3762) );
  INV_X1 U4372 ( .A(n4820), .ZN(n3760) );
  OR2_X1 U4373 ( .A1(n4774), .A2(n5107), .ZN(n3756) );
  NAND2_X1 U4374 ( .A1(n4475), .A2(n5054), .ZN(n3755) );
  NAND2_X1 U4375 ( .A1(n3756), .A2(n3755), .ZN(n4811) );
  AOI22_X1 U4376 ( .A1(n4811), .A2(n5243), .B1(REG3_REG_14__SCAN_IN), .B2(
        U3149), .ZN(n3759) );
  NAND2_X1 U4377 ( .A1(n5267), .A2(n3757), .ZN(n3758) );
  OAI211_X1 U4378 ( .C1(n5326), .C2(n3760), .A(n3759), .B(n3758), .ZN(n3761)
         );
  AOI21_X1 U4379 ( .B1(n3762), .B2(n5322), .A(n3761), .ZN(n3763) );
  INV_X1 U4380 ( .A(n3763), .ZN(U3212) );
  INV_X1 U4381 ( .A(n3764), .ZN(n4286) );
  OAI21_X1 U4382 ( .B1(n4286), .B2(n3766), .A(n3765), .ZN(n3768) );
  NAND3_X1 U4383 ( .A1(n3768), .A2(n5322), .A3(n3767), .ZN(n3774) );
  AOI22_X1 U4384 ( .A1(n5264), .A2(n4710), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3773) );
  AOI22_X1 U4385 ( .A1(n3769), .A2(n5267), .B1(n5258), .B2(n4668), .ZN(n3772)
         );
  INV_X1 U4386 ( .A(n3770), .ZN(n4672) );
  OR2_X1 U4387 ( .A1(n5326), .A2(n4672), .ZN(n3771) );
  NAND4_X1 U4388 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(U3213)
         );
  AND2_X1 U4389 ( .A1(n3775), .A2(n3776), .ZN(n3779) );
  OAI211_X1 U4390 ( .C1(n3779), .C2(n3778), .A(n5322), .B(n3777), .ZN(n3786)
         );
  AOI22_X1 U4391 ( .A1(n3780), .A2(n5243), .B1(REG3_REG_10__SCAN_IN), .B2(
        U3149), .ZN(n3785) );
  OR2_X1 U4392 ( .A1(n5326), .A2(n3781), .ZN(n3784) );
  NAND2_X1 U4393 ( .A1(n5267), .A2(n3782), .ZN(n3783) );
  NAND4_X1 U4394 ( .A1(n3786), .A2(n3785), .A3(n3784), .A4(n3783), .ZN(U3214)
         );
  OAI21_X1 U4395 ( .B1(n3789), .B2(n3788), .A(n3787), .ZN(n3790) );
  NAND2_X1 U4396 ( .A1(n3790), .A2(n5322), .ZN(n3798) );
  INV_X1 U4397 ( .A(n3791), .ZN(n3792) );
  OAI21_X1 U4398 ( .B1(n3794), .B2(n3793), .A(n3792), .ZN(n3795) );
  AOI21_X1 U4399 ( .B1(n3796), .B2(n5267), .A(n3795), .ZN(n3797) );
  OAI211_X1 U4400 ( .C1(n5326), .C2(n3799), .A(n3798), .B(n3797), .ZN(U3218)
         );
  OAI211_X1 U4401 ( .C1(n3802), .C2(n3801), .A(n3800), .B(n5322), .ZN(n3807)
         );
  AOI22_X1 U4402 ( .A1(n5264), .A2(n3418), .B1(n5258), .B2(n3471), .ZN(n3806)
         );
  AOI22_X1 U4403 ( .A1(n5267), .A2(n3804), .B1(n3803), .B2(REG3_REG_1__SCAN_IN), .ZN(n3805) );
  NAND3_X1 U4404 ( .A1(n3807), .A2(n3806), .A3(n3805), .ZN(U3219) );
  INV_X1 U4405 ( .A(n3808), .ZN(n3813) );
  OR2_X1 U4406 ( .A1(n3809), .A2(n5286), .ZN(n3811) );
  NAND2_X1 U4407 ( .A1(n4475), .A2(n5283), .ZN(n3810) );
  NAND2_X1 U4408 ( .A1(n3811), .A2(n3810), .ZN(n4828) );
  NAND2_X1 U4409 ( .A1(n4828), .A2(n5243), .ZN(n3812) );
  OAI211_X1 U4410 ( .C1(n5319), .C2(n4832), .A(n3813), .B(n3812), .ZN(n3821)
         );
  INV_X1 U4411 ( .A(n3815), .ZN(n3816) );
  NAND3_X1 U4412 ( .A1(n3814), .A2(n3817), .A3(n3816), .ZN(n3818) );
  AOI21_X1 U4413 ( .B1(n3819), .B2(n3818), .A(n5226), .ZN(n3820) );
  AOI211_X1 U4414 ( .C1(n4834), .C2(n4301), .A(n3821), .B(n3820), .ZN(n3822)
         );
  INV_X1 U4415 ( .A(n3822), .ZN(U3221) );
  INV_X1 U4416 ( .A(n3824), .ZN(n3825) );
  AOI21_X1 U4417 ( .B1(n3826), .B2(n3823), .A(n3825), .ZN(n3831) );
  INV_X1 U4418 ( .A(n5264), .ZN(n5315) );
  OAI22_X1 U4419 ( .A1(n5315), .A2(n3827), .B1(STATE_REG_SCAN_IN), .B2(n3918), 
        .ZN(n3829) );
  INV_X1 U4420 ( .A(n5258), .ZN(n5317) );
  OAI22_X1 U4421 ( .A1(n5319), .A2(n4638), .B1(n5317), .B2(n4634), .ZN(n3828)
         );
  AOI211_X1 U4422 ( .C1(n4640), .C2(n4301), .A(n3829), .B(n3828), .ZN(n3830)
         );
  OAI21_X1 U4423 ( .B1(n3831), .B2(n5226), .A(n3830), .ZN(U3222) );
  INV_X1 U4424 ( .A(n4785), .ZN(n3844) );
  AND2_X1 U4425 ( .A1(n3832), .A2(n3849), .ZN(n3838) );
  INV_X1 U4426 ( .A(n5191), .ZN(n3836) );
  INV_X1 U4427 ( .A(n3833), .ZN(n3834) );
  AOI21_X1 U4428 ( .B1(n3834), .B2(n5191), .A(n5190), .ZN(n3835) );
  AOI21_X1 U4429 ( .B1(n3833), .B2(n3836), .A(n3835), .ZN(n3837) );
  NAND2_X1 U4430 ( .A1(n3837), .A2(n3838), .ZN(n3850) );
  OAI21_X1 U4431 ( .B1(n3838), .B2(n3837), .A(n3850), .ZN(n3839) );
  NAND2_X1 U4432 ( .A1(n3839), .A2(n5322), .ZN(n3843) );
  NOR2_X1 U4433 ( .A1(STATE_REG_SCAN_IN), .A2(n3840), .ZN(n4547) );
  OAI22_X1 U4434 ( .A1(n5319), .A2(n4779), .B1(n5315), .B2(n4774), .ZN(n3841)
         );
  AOI211_X1 U4435 ( .C1(n5258), .C2(n4472), .A(n4547), .B(n3841), .ZN(n3842)
         );
  OAI211_X1 U4436 ( .C1(n5326), .C2(n3844), .A(n3843), .B(n3842), .ZN(U3223)
         );
  AOI22_X1 U4437 ( .A1(n4761), .A2(n5246), .B1(n5264), .B2(n4756), .ZN(n3846)
         );
  NOR2_X1 U4438 ( .A1(STATE_REG_SCAN_IN), .A2(n3925), .ZN(n4564) );
  INV_X1 U4439 ( .A(n4564), .ZN(n3845) );
  OAI211_X1 U4440 ( .C1(n4757), .C2(n5317), .A(n3846), .B(n3845), .ZN(n3854)
         );
  INV_X1 U4441 ( .A(n3847), .ZN(n3848) );
  NAND3_X1 U4442 ( .A1(n3850), .A2(n3849), .A3(n3848), .ZN(n3852) );
  AOI21_X1 U4443 ( .B1(n3852), .B2(n3851), .A(n5226), .ZN(n3853) );
  AOI211_X1 U4444 ( .C1(n4763), .C2(n4301), .A(n3854), .B(n3853), .ZN(n4252)
         );
  XOR2_X1 U4445 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_126), .Z(n4250) );
  XOR2_X1 U4446 ( .A(DATAI_30_), .B(keyinput_1), .Z(n3857) );
  XOR2_X1 U4447 ( .A(DATAI_31_), .B(keyinput_0), .Z(n3856) );
  XNOR2_X1 U4448 ( .A(DATAI_29_), .B(keyinput_2), .ZN(n3855) );
  NAND3_X1 U4449 ( .A1(n3857), .A2(n3856), .A3(n3855), .ZN(n3861) );
  XOR2_X1 U4450 ( .A(DATAI_28_), .B(keyinput_3), .Z(n3860) );
  XNOR2_X1 U4451 ( .A(DATAI_26_), .B(keyinput_5), .ZN(n3859) );
  XNOR2_X1 U4452 ( .A(DATAI_27_), .B(keyinput_4), .ZN(n3858) );
  AOI211_X1 U4453 ( .C1(n3861), .C2(n3860), .A(n3859), .B(n3858), .ZN(n3868)
         );
  XOR2_X1 U4454 ( .A(DATAI_23_), .B(keyinput_8), .Z(n3865) );
  XNOR2_X1 U4455 ( .A(DATAI_22_), .B(keyinput_9), .ZN(n3864) );
  XNOR2_X1 U4456 ( .A(DATAI_24_), .B(keyinput_7), .ZN(n3863) );
  XNOR2_X1 U4457 ( .A(DATAI_25_), .B(keyinput_6), .ZN(n3862) );
  NAND4_X1 U4458 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3867)
         );
  XOR2_X1 U4459 ( .A(DATAI_21_), .B(keyinput_10), .Z(n3866) );
  OAI21_X1 U4460 ( .B1(n3868), .B2(n3867), .A(n3866), .ZN(n3871) );
  XNOR2_X1 U4461 ( .A(DATAI_20_), .B(keyinput_11), .ZN(n3870) );
  XNOR2_X1 U4462 ( .A(DATAI_19_), .B(keyinput_12), .ZN(n3869) );
  AOI21_X1 U4463 ( .B1(n3871), .B2(n3870), .A(n3869), .ZN(n3879) );
  XNOR2_X1 U4464 ( .A(n4062), .B(keyinput_17), .ZN(n3878) );
  XNOR2_X1 U4465 ( .A(DATAI_17_), .B(keyinput_14), .ZN(n3877) );
  XNOR2_X1 U4466 ( .A(n3872), .B(keyinput_15), .ZN(n3875) );
  XNOR2_X1 U4467 ( .A(DATAI_15_), .B(keyinput_16), .ZN(n3874) );
  XNOR2_X1 U4468 ( .A(DATAI_18_), .B(keyinput_13), .ZN(n3873) );
  NAND3_X1 U4469 ( .A1(n3875), .A2(n3874), .A3(n3873), .ZN(n3876) );
  NOR4_X1 U4470 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3888)
         );
  XNOR2_X1 U4471 ( .A(DATAI_13_), .B(keyinput_18), .ZN(n3887) );
  XOR2_X1 U4472 ( .A(DATAI_11_), .B(keyinput_20), .Z(n3882) );
  XNOR2_X1 U4473 ( .A(DATAI_12_), .B(keyinput_19), .ZN(n3881) );
  XNOR2_X1 U4474 ( .A(DATAI_9_), .B(keyinput_22), .ZN(n3880) );
  NAND3_X1 U4475 ( .A1(n3882), .A2(n3881), .A3(n3880), .ZN(n3885) );
  XNOR2_X1 U4476 ( .A(DATAI_8_), .B(keyinput_23), .ZN(n3884) );
  XNOR2_X1 U4477 ( .A(DATAI_10_), .B(keyinput_21), .ZN(n3883) );
  NOR3_X1 U4478 ( .A1(n3885), .A2(n3884), .A3(n3883), .ZN(n3886) );
  OAI21_X1 U4479 ( .B1(n3888), .B2(n3887), .A(n3886), .ZN(n3891) );
  XOR2_X1 U4480 ( .A(DATAI_7_), .B(keyinput_24), .Z(n3890) );
  XNOR2_X1 U4481 ( .A(DATAI_6_), .B(keyinput_25), .ZN(n3889) );
  NAND3_X1 U4482 ( .A1(n3891), .A2(n3890), .A3(n3889), .ZN(n3894) );
  XNOR2_X1 U4483 ( .A(DATAI_5_), .B(keyinput_26), .ZN(n3893) );
  XNOR2_X1 U4484 ( .A(DATAI_4_), .B(keyinput_27), .ZN(n3892) );
  AOI21_X1 U4485 ( .B1(n3894), .B2(n3893), .A(n3892), .ZN(n3900) );
  XOR2_X1 U4486 ( .A(DATAI_3_), .B(keyinput_28), .Z(n3899) );
  XNOR2_X1 U4487 ( .A(n2721), .B(keyinput_31), .ZN(n3897) );
  XNOR2_X1 U4488 ( .A(DATAI_2_), .B(keyinput_29), .ZN(n3896) );
  XNOR2_X1 U4489 ( .A(DATAI_1_), .B(keyinput_30), .ZN(n3895) );
  NOR3_X1 U4490 ( .A1(n3897), .A2(n3896), .A3(n3895), .ZN(n3898) );
  OAI21_X1 U4491 ( .B1(n3900), .B2(n3899), .A(n3898), .ZN(n3903) );
  XNOR2_X1 U4492 ( .A(U3149), .B(keyinput_32), .ZN(n3902) );
  XNOR2_X1 U4493 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_33), .ZN(n3901) );
  NAND3_X1 U4494 ( .A1(n3903), .A2(n3902), .A3(n3901), .ZN(n3906) );
  XNOR2_X1 U4495 ( .A(n4098), .B(keyinput_34), .ZN(n3905) );
  XOR2_X1 U4496 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_35), .Z(n3904) );
  NAND3_X1 U4497 ( .A1(n3906), .A2(n3905), .A3(n3904), .ZN(n3909) );
  XOR2_X1 U4498 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_36), .Z(n3908) );
  XNOR2_X1 U4499 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_37), .ZN(n3907) );
  AOI21_X1 U4500 ( .B1(n3909), .B2(n3908), .A(n3907), .ZN(n3914) );
  XNOR2_X1 U4501 ( .A(n5066), .B(keyinput_38), .ZN(n3913) );
  XNOR2_X1 U4502 ( .A(n3910), .B(keyinput_40), .ZN(n3912) );
  XNOR2_X1 U4503 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_39), .ZN(n3911) );
  OAI211_X1 U4504 ( .C1(n3914), .C2(n3913), .A(n3912), .B(n3911), .ZN(n3917)
         );
  XNOR2_X1 U4505 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_41), .ZN(n3916) );
  XNOR2_X1 U4506 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .ZN(n3915) );
  NAND3_X1 U4507 ( .A1(n3917), .A2(n3916), .A3(n3915), .ZN(n3924) );
  XNOR2_X1 U4508 ( .A(n5313), .B(keyinput_43), .ZN(n3923) );
  XNOR2_X1 U4509 ( .A(n3918), .B(keyinput_45), .ZN(n3921) );
  XNOR2_X1 U4510 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput_46), .ZN(n3920) );
  XNOR2_X1 U4511 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_44), .ZN(n3919) );
  NAND3_X1 U4512 ( .A1(n3921), .A2(n3920), .A3(n3919), .ZN(n3922) );
  AOI21_X1 U4513 ( .B1(n3924), .B2(n3923), .A(n3922), .ZN(n3929) );
  XOR2_X1 U4514 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_47), .Z(n3928) );
  XNOR2_X1 U4515 ( .A(n3925), .B(keyinput_48), .ZN(n3927) );
  XNOR2_X1 U4516 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_49), .ZN(n3926) );
  OAI211_X1 U4517 ( .C1(n3929), .C2(n3928), .A(n3927), .B(n3926), .ZN(n3936)
         );
  XOR2_X1 U4518 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput_51), .Z(n3935) );
  XOR2_X1 U4519 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_52), .Z(n3932) );
  XOR2_X1 U4520 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_53), .Z(n3931) );
  XNOR2_X1 U4521 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_50), .ZN(n3930) );
  NOR3_X1 U4522 ( .A1(n3932), .A2(n3931), .A3(n3930), .ZN(n3934) );
  XNOR2_X1 U4523 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_54), .ZN(n3933) );
  NAND4_X1 U4524 ( .A1(n3936), .A2(n3935), .A3(n3934), .A4(n3933), .ZN(n3939)
         );
  XNOR2_X1 U4525 ( .A(n4958), .B(keyinput_55), .ZN(n3938) );
  XOR2_X1 U4526 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_56), .Z(n3937) );
  AOI21_X1 U4527 ( .B1(n3939), .B2(n3938), .A(n3937), .ZN(n3946) );
  XNOR2_X1 U4528 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n3943) );
  XNOR2_X1 U4529 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_58), .ZN(n3942) );
  XNOR2_X1 U4530 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_57), .ZN(n3941) );
  XNOR2_X1 U4531 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_59), .ZN(n3940) );
  NAND4_X1 U4532 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3945)
         );
  XNOR2_X1 U4533 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_61), .ZN(n3944) );
  OAI21_X1 U4534 ( .B1(n3946), .B2(n3945), .A(n3944), .ZN(n3951) );
  OAI22_X1 U4535 ( .A1(n4141), .A2(keyinput_63), .B1(keyinput_62), .B2(
        IR_REG_7__SCAN_IN), .ZN(n3947) );
  AOI21_X1 U4536 ( .B1(IR_REG_7__SCAN_IN), .B2(keyinput_62), .A(n3947), .ZN(
        n3950) );
  XNOR2_X1 U4537 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_64), .ZN(n3949) );
  NAND2_X1 U4538 ( .A1(n4141), .A2(keyinput_63), .ZN(n3948) );
  NAND4_X1 U4539 ( .A1(n3951), .A2(n3950), .A3(n3949), .A4(n3948), .ZN(n3958)
         );
  XOR2_X1 U4540 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_65), .Z(n3957) );
  XOR2_X1 U4541 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_67), .Z(n3955) );
  XNOR2_X1 U4542 ( .A(n4147), .B(keyinput_69), .ZN(n3954) );
  XNOR2_X1 U4543 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_68), .ZN(n3953) );
  XNOR2_X1 U4544 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_66), .ZN(n3952) );
  NAND4_X1 U4545 ( .A1(n3955), .A2(n3954), .A3(n3953), .A4(n3952), .ZN(n3956)
         );
  AOI21_X1 U4546 ( .B1(n3958), .B2(n3957), .A(n3956), .ZN(n3961) );
  XNOR2_X1 U4547 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_70), .ZN(n3960) );
  XNOR2_X1 U4548 ( .A(n4155), .B(keyinput_71), .ZN(n3959) );
  OAI21_X1 U4549 ( .B1(n3961), .B2(n3960), .A(n3959), .ZN(n3964) );
  XNOR2_X1 U4550 ( .A(n4159), .B(keyinput_72), .ZN(n3963) );
  XNOR2_X1 U4551 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_73), .ZN(n3962) );
  AOI21_X1 U4552 ( .B1(n3964), .B2(n3963), .A(n3962), .ZN(n3972) );
  XNOR2_X1 U4553 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_74), .ZN(n3971) );
  XOR2_X1 U4554 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_76), .Z(n3969) );
  XNOR2_X1 U4555 ( .A(n3965), .B(keyinput_78), .ZN(n3968) );
  XNOR2_X1 U4556 ( .A(IR_REG_20__SCAN_IN), .B(keyinput_75), .ZN(n3967) );
  XNOR2_X1 U4557 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_77), .ZN(n3966) );
  NOR4_X1 U4558 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3970)
         );
  OAI21_X1 U4559 ( .B1(n3972), .B2(n3971), .A(n3970), .ZN(n3988) );
  XNOR2_X1 U4560 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_79), .ZN(n3987) );
  XOR2_X1 U4561 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_86), .Z(n3977) );
  XNOR2_X1 U4562 ( .A(n4172), .B(keyinput_84), .ZN(n3976) );
  XNOR2_X1 U4563 ( .A(n4173), .B(keyinput_87), .ZN(n3975) );
  XNOR2_X1 U4564 ( .A(keyinput_88), .B(n3973), .ZN(n3974) );
  NOR4_X1 U4565 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(n3985)
         );
  XNOR2_X1 U4566 ( .A(n4174), .B(keyinput_85), .ZN(n3984) );
  XOR2_X1 U4567 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_80), .Z(n3983) );
  XNOR2_X1 U4568 ( .A(n2683), .B(keyinput_83), .ZN(n3981) );
  XNOR2_X1 U4569 ( .A(n3978), .B(keyinput_82), .ZN(n3980) );
  XNOR2_X1 U4570 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_81), .ZN(n3979) );
  NOR3_X1 U4571 ( .A1(n3981), .A2(n3980), .A3(n3979), .ZN(n3982) );
  NAND4_X1 U4572 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3986)
         );
  AOI21_X1 U4573 ( .B1(n3988), .B2(n3987), .A(n3986), .ZN(n3995) );
  XNOR2_X1 U4574 ( .A(D_REG_2__SCAN_IN), .B(keyinput_89), .ZN(n3994) );
  INV_X1 U4575 ( .A(D_REG_4__SCAN_IN), .ZN(n4932) );
  XNOR2_X1 U4576 ( .A(n4932), .B(keyinput_91), .ZN(n3992) );
  XNOR2_X1 U4577 ( .A(D_REG_5__SCAN_IN), .B(keyinput_92), .ZN(n3991) );
  XNOR2_X1 U4578 ( .A(D_REG_6__SCAN_IN), .B(keyinput_93), .ZN(n3990) );
  XNOR2_X1 U4579 ( .A(D_REG_3__SCAN_IN), .B(keyinput_90), .ZN(n3989) );
  NOR4_X1 U4580 ( .A1(n3992), .A2(n3991), .A3(n3990), .A4(n3989), .ZN(n3993)
         );
  OAI21_X1 U4581 ( .B1(n3995), .B2(n3994), .A(n3993), .ZN(n3998) );
  XNOR2_X1 U4582 ( .A(D_REG_7__SCAN_IN), .B(keyinput_94), .ZN(n3997) );
  XOR2_X1 U4583 ( .A(D_REG_8__SCAN_IN), .B(keyinput_95), .Z(n3996) );
  AOI21_X1 U4584 ( .B1(n3998), .B2(n3997), .A(n3996), .ZN(n4007) );
  INV_X1 U4585 ( .A(D_REG_11__SCAN_IN), .ZN(n4003) );
  INV_X1 U4586 ( .A(keyinput_98), .ZN(n4002) );
  XNOR2_X1 U4587 ( .A(D_REG_10__SCAN_IN), .B(keyinput_97), .ZN(n4001) );
  OAI22_X1 U4588 ( .A1(D_REG_9__SCAN_IN), .A2(keyinput_96), .B1(
        D_REG_11__SCAN_IN), .B2(keyinput_98), .ZN(n3999) );
  AOI21_X1 U4589 ( .B1(D_REG_9__SCAN_IN), .B2(keyinput_96), .A(n3999), .ZN(
        n4000) );
  OAI211_X1 U4590 ( .C1(n4003), .C2(n4002), .A(n4001), .B(n4000), .ZN(n4006)
         );
  XNOR2_X1 U4591 ( .A(D_REG_13__SCAN_IN), .B(keyinput_100), .ZN(n4005) );
  XNOR2_X1 U4592 ( .A(D_REG_12__SCAN_IN), .B(keyinput_99), .ZN(n4004) );
  OAI211_X1 U4593 ( .C1(n4007), .C2(n4006), .A(n4005), .B(n4004), .ZN(n4010)
         );
  XNOR2_X1 U4594 ( .A(D_REG_14__SCAN_IN), .B(keyinput_101), .ZN(n4009) );
  INV_X1 U4595 ( .A(D_REG_15__SCAN_IN), .ZN(n4940) );
  XNOR2_X1 U4596 ( .A(n4940), .B(keyinput_102), .ZN(n4008) );
  AOI21_X1 U4597 ( .B1(n4010), .B2(n4009), .A(n4008), .ZN(n4013) );
  XOR2_X1 U4598 ( .A(D_REG_16__SCAN_IN), .B(keyinput_103), .Z(n4012) );
  INV_X1 U4599 ( .A(D_REG_17__SCAN_IN), .ZN(n4942) );
  XNOR2_X1 U4600 ( .A(n4942), .B(keyinput_104), .ZN(n4011) );
  NOR3_X1 U4601 ( .A1(n4013), .A2(n4012), .A3(n4011), .ZN(n4016) );
  INV_X1 U4602 ( .A(D_REG_18__SCAN_IN), .ZN(n4943) );
  XNOR2_X1 U4603 ( .A(n4943), .B(keyinput_105), .ZN(n4015) );
  INV_X1 U4604 ( .A(D_REG_19__SCAN_IN), .ZN(n4944) );
  XNOR2_X1 U4605 ( .A(n4944), .B(keyinput_106), .ZN(n4014) );
  OAI21_X1 U4606 ( .B1(n4016), .B2(n4015), .A(n4014), .ZN(n4020) );
  INV_X1 U4607 ( .A(D_REG_20__SCAN_IN), .ZN(n4945) );
  XNOR2_X1 U4608 ( .A(n4945), .B(keyinput_107), .ZN(n4019) );
  XNOR2_X1 U4609 ( .A(D_REG_22__SCAN_IN), .B(keyinput_109), .ZN(n4018) );
  XNOR2_X1 U4610 ( .A(D_REG_21__SCAN_IN), .B(keyinput_108), .ZN(n4017) );
  AOI211_X1 U4611 ( .C1(n4020), .C2(n4019), .A(n4018), .B(n4017), .ZN(n4023)
         );
  XNOR2_X1 U4612 ( .A(D_REG_23__SCAN_IN), .B(keyinput_110), .ZN(n4022) );
  XNOR2_X1 U4613 ( .A(D_REG_24__SCAN_IN), .B(keyinput_111), .ZN(n4021) );
  OAI21_X1 U4614 ( .B1(n4023), .B2(n4022), .A(n4021), .ZN(n4026) );
  INV_X1 U4615 ( .A(D_REG_25__SCAN_IN), .ZN(n4949) );
  XNOR2_X1 U4616 ( .A(n4949), .B(keyinput_112), .ZN(n4025) );
  XNOR2_X1 U4617 ( .A(D_REG_26__SCAN_IN), .B(keyinput_113), .ZN(n4024) );
  AOI21_X1 U4618 ( .B1(n4026), .B2(n4025), .A(n4024), .ZN(n4029) );
  INV_X1 U4619 ( .A(D_REG_28__SCAN_IN), .ZN(n4952) );
  XNOR2_X1 U4620 ( .A(n4952), .B(keyinput_115), .ZN(n4028) );
  XNOR2_X1 U4621 ( .A(D_REG_27__SCAN_IN), .B(keyinput_114), .ZN(n4027) );
  NOR3_X1 U4622 ( .A1(n4029), .A2(n4028), .A3(n4027), .ZN(n4032) );
  INV_X1 U4623 ( .A(D_REG_29__SCAN_IN), .ZN(n4953) );
  XNOR2_X1 U4624 ( .A(n4953), .B(keyinput_116), .ZN(n4031) );
  XNOR2_X1 U4625 ( .A(D_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n4030) );
  NOR3_X1 U4626 ( .A1(n4032), .A2(n4031), .A3(n4030), .ZN(n4038) );
  XNOR2_X1 U4627 ( .A(D_REG_31__SCAN_IN), .B(keyinput_118), .ZN(n4037) );
  XOR2_X1 U4628 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_119), .Z(n4035) );
  XNOR2_X1 U4629 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_121), .ZN(n4034) );
  XNOR2_X1 U4630 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_120), .ZN(n4033) );
  NOR3_X1 U4631 ( .A1(n4035), .A2(n4034), .A3(n4033), .ZN(n4036) );
  OAI21_X1 U4632 ( .B1(n4038), .B2(n4037), .A(n4036), .ZN(n4041) );
  XNOR2_X1 U4633 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_122), .ZN(n4040) );
  XNOR2_X1 U4634 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_123), .ZN(n4039) );
  AOI21_X1 U4635 ( .B1(n4041), .B2(n4040), .A(n4039), .ZN(n4044) );
  XOR2_X1 U4636 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_124), .Z(n4043) );
  XOR2_X1 U4637 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_125), .Z(n4042) );
  OAI21_X1 U4638 ( .B1(n4044), .B2(n4043), .A(n4042), .ZN(n4249) );
  XOR2_X1 U4639 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_127), .Z(n4248) );
  XOR2_X1 U4640 ( .A(DATAI_28_), .B(keyinput_131), .Z(n4051) );
  XOR2_X1 U4641 ( .A(DATAI_31_), .B(keyinput_128), .Z(n4047) );
  XOR2_X1 U4642 ( .A(DATAI_30_), .B(keyinput_129), .Z(n4046) );
  XOR2_X1 U4643 ( .A(DATAI_29_), .B(keyinput_130), .Z(n4045) );
  NAND3_X1 U4644 ( .A1(n4047), .A2(n4046), .A3(n4045), .ZN(n4050) );
  XNOR2_X1 U4645 ( .A(DATAI_26_), .B(keyinput_133), .ZN(n4049) );
  XOR2_X1 U4646 ( .A(DATAI_27_), .B(keyinput_132), .Z(n4048) );
  AOI211_X1 U4647 ( .C1(n4051), .C2(n4050), .A(n4049), .B(n4048), .ZN(n4058)
         );
  XOR2_X1 U4648 ( .A(DATAI_23_), .B(keyinput_136), .Z(n4055) );
  XOR2_X1 U4649 ( .A(DATAI_25_), .B(keyinput_134), .Z(n4054) );
  XOR2_X1 U4650 ( .A(DATAI_24_), .B(keyinput_135), .Z(n4053) );
  XNOR2_X1 U4651 ( .A(DATAI_22_), .B(keyinput_137), .ZN(n4052) );
  NAND4_X1 U4652 ( .A1(n4055), .A2(n4054), .A3(n4053), .A4(n4052), .ZN(n4057)
         );
  XOR2_X1 U4653 ( .A(DATAI_21_), .B(keyinput_138), .Z(n4056) );
  OAI21_X1 U4654 ( .B1(n4058), .B2(n4057), .A(n4056), .ZN(n4061) );
  XNOR2_X1 U4655 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n4060) );
  XNOR2_X1 U4656 ( .A(DATAI_19_), .B(keyinput_140), .ZN(n4059) );
  AOI21_X1 U4657 ( .B1(n4061), .B2(n4060), .A(n4059), .ZN(n4069) );
  XNOR2_X1 U4658 ( .A(DATAI_18_), .B(keyinput_141), .ZN(n4068) );
  XNOR2_X1 U4659 ( .A(DATAI_17_), .B(keyinput_142), .ZN(n4067) );
  XNOR2_X1 U4660 ( .A(n4062), .B(keyinput_145), .ZN(n4065) );
  XNOR2_X1 U4661 ( .A(DATAI_16_), .B(keyinput_143), .ZN(n4064) );
  XNOR2_X1 U4662 ( .A(DATAI_15_), .B(keyinput_144), .ZN(n4063) );
  NAND3_X1 U4663 ( .A1(n4065), .A2(n4064), .A3(n4063), .ZN(n4066) );
  NOR4_X1 U4664 ( .A1(n4069), .A2(n4068), .A3(n4067), .A4(n4066), .ZN(n4080)
         );
  XNOR2_X1 U4665 ( .A(n4070), .B(keyinput_146), .ZN(n4079) );
  XOR2_X1 U4666 ( .A(DATAI_12_), .B(keyinput_147), .Z(n4074) );
  XNOR2_X1 U4667 ( .A(n4071), .B(keyinput_150), .ZN(n4073) );
  XNOR2_X1 U4668 ( .A(DATAI_8_), .B(keyinput_151), .ZN(n4072) );
  NAND3_X1 U4669 ( .A1(n4074), .A2(n4073), .A3(n4072), .ZN(n4077) );
  XNOR2_X1 U4670 ( .A(DATAI_11_), .B(keyinput_148), .ZN(n4076) );
  XNOR2_X1 U4671 ( .A(DATAI_10_), .B(keyinput_149), .ZN(n4075) );
  NOR3_X1 U4672 ( .A1(n4077), .A2(n4076), .A3(n4075), .ZN(n4078) );
  OAI21_X1 U4673 ( .B1(n4080), .B2(n4079), .A(n4078), .ZN(n4084) );
  XNOR2_X1 U4674 ( .A(n4081), .B(keyinput_153), .ZN(n4083) );
  XNOR2_X1 U4675 ( .A(DATAI_7_), .B(keyinput_152), .ZN(n4082) );
  NAND3_X1 U4676 ( .A1(n4084), .A2(n4083), .A3(n4082), .ZN(n4088) );
  XNOR2_X1 U4677 ( .A(DATAI_5_), .B(keyinput_154), .ZN(n4087) );
  XNOR2_X1 U4678 ( .A(n4085), .B(keyinput_155), .ZN(n4086) );
  AOI21_X1 U4679 ( .B1(n4088), .B2(n4087), .A(n4086), .ZN(n4094) );
  XNOR2_X1 U4680 ( .A(DATAI_3_), .B(keyinput_156), .ZN(n4093) );
  INV_X1 U4681 ( .A(DATAI_2_), .ZN(n5038) );
  XNOR2_X1 U4682 ( .A(n5038), .B(keyinput_157), .ZN(n4091) );
  INV_X1 U4683 ( .A(DATAI_1_), .ZN(n5030) );
  XNOR2_X1 U4684 ( .A(n5030), .B(keyinput_158), .ZN(n4090) );
  XNOR2_X1 U4685 ( .A(DATAI_0_), .B(keyinput_159), .ZN(n4089) );
  NOR3_X1 U4686 ( .A1(n4091), .A2(n4090), .A3(n4089), .ZN(n4092) );
  OAI21_X1 U4687 ( .B1(n4094), .B2(n4093), .A(n4092), .ZN(n4097) );
  XNOR2_X1 U4688 ( .A(STATE_REG_SCAN_IN), .B(keyinput_160), .ZN(n4096) );
  XNOR2_X1 U4689 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_161), .ZN(n4095) );
  NAND3_X1 U4690 ( .A1(n4097), .A2(n4096), .A3(n4095), .ZN(n4101) );
  XNOR2_X1 U4691 ( .A(n4098), .B(keyinput_162), .ZN(n4100) );
  XOR2_X1 U4692 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_163), .Z(n4099) );
  NAND3_X1 U4693 ( .A1(n4101), .A2(n4100), .A3(n4099), .ZN(n4104) );
  XNOR2_X1 U4694 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_164), .ZN(n4103) );
  XNOR2_X1 U4695 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_165), .ZN(n4102) );
  AOI21_X1 U4696 ( .B1(n4104), .B2(n4103), .A(n4102), .ZN(n4108) );
  XNOR2_X1 U4697 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_166), .ZN(n4107) );
  XOR2_X1 U4698 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_167), .Z(n4106) );
  XNOR2_X1 U4699 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput_168), .ZN(n4105) );
  OAI211_X1 U4700 ( .C1(n4108), .C2(n4107), .A(n4106), .B(n4105), .ZN(n4111)
         );
  XOR2_X1 U4701 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_170), .Z(n4110) );
  XNOR2_X1 U4702 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_169), .ZN(n4109) );
  NAND3_X1 U4703 ( .A1(n4111), .A2(n4110), .A3(n4109), .ZN(n4117) );
  XNOR2_X1 U4704 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_171), .ZN(n4116) );
  XNOR2_X1 U4705 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput_174), .ZN(n4114) );
  XNOR2_X1 U4706 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_173), .ZN(n4113) );
  XNOR2_X1 U4707 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_172), .ZN(n4112) );
  NAND3_X1 U4708 ( .A1(n4114), .A2(n4113), .A3(n4112), .ZN(n4115) );
  AOI21_X1 U4709 ( .B1(n4117), .B2(n4116), .A(n4115), .ZN(n4121) );
  XNOR2_X1 U4710 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_175), .ZN(n4120) );
  XNOR2_X1 U4711 ( .A(n4258), .B(keyinput_177), .ZN(n4119) );
  XNOR2_X1 U4712 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_176), .ZN(n4118) );
  OAI211_X1 U4713 ( .C1(n4121), .C2(n4120), .A(n4119), .B(n4118), .ZN(n4130)
         );
  XOR2_X1 U4714 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_181), .Z(n4127) );
  XNOR2_X1 U4715 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_178), .ZN(n4123) );
  XNOR2_X1 U4716 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_182), .ZN(n4122) );
  NAND2_X1 U4717 ( .A1(n4123), .A2(n4122), .ZN(n4126) );
  XNOR2_X1 U4718 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput_179), .ZN(n4125) );
  XNOR2_X1 U4719 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_180), .ZN(n4124) );
  NOR4_X1 U4720 ( .A1(n4127), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n4129)
         );
  XOR2_X1 U4721 ( .A(n4958), .B(keyinput_183), .Z(n4128) );
  AOI21_X1 U4722 ( .B1(n4130), .B2(n4129), .A(n4128), .ZN(n4137) );
  XOR2_X1 U4723 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_184), .Z(n4136) );
  XNOR2_X1 U4724 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_188), .ZN(n4134) );
  XNOR2_X1 U4725 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_187), .ZN(n4133) );
  XNOR2_X1 U4726 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_185), .ZN(n4132) );
  XNOR2_X1 U4727 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_186), .ZN(n4131) );
  NOR4_X1 U4728 ( .A1(n4134), .A2(n4133), .A3(n4132), .A4(n4131), .ZN(n4135)
         );
  OAI21_X1 U4729 ( .B1(n4137), .B2(n4136), .A(n4135), .ZN(n4139) );
  XNOR2_X1 U4730 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n4138) );
  NAND2_X1 U4731 ( .A1(n4139), .A2(n4138), .ZN(n4145) );
  XNOR2_X1 U4732 ( .A(n4140), .B(keyinput_190), .ZN(n4144) );
  XNOR2_X1 U4733 ( .A(n4141), .B(keyinput_191), .ZN(n4143) );
  XNOR2_X1 U4734 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_192), .ZN(n4142) );
  NAND4_X1 U4735 ( .A1(n4145), .A2(n4144), .A3(n4143), .A4(n4142), .ZN(n4154)
         );
  XOR2_X1 U4736 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_193), .Z(n4153) );
  XNOR2_X1 U4737 ( .A(n4146), .B(keyinput_194), .ZN(n4151) );
  XNOR2_X1 U4738 ( .A(n4147), .B(keyinput_197), .ZN(n4150) );
  XNOR2_X1 U4739 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_196), .ZN(n4149) );
  XNOR2_X1 U4740 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_195), .ZN(n4148) );
  NAND4_X1 U4741 ( .A1(n4151), .A2(n4150), .A3(n4149), .A4(n4148), .ZN(n4152)
         );
  AOI21_X1 U4742 ( .B1(n4154), .B2(n4153), .A(n4152), .ZN(n4158) );
  XNOR2_X1 U4743 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_198), .ZN(n4157) );
  XNOR2_X1 U4744 ( .A(n4155), .B(keyinput_199), .ZN(n4156) );
  OAI21_X1 U4745 ( .B1(n4158), .B2(n4157), .A(n4156), .ZN(n4163) );
  XNOR2_X1 U4746 ( .A(n4159), .B(keyinput_200), .ZN(n4162) );
  XNOR2_X1 U4747 ( .A(n4160), .B(keyinput_201), .ZN(n4161) );
  AOI21_X1 U4748 ( .B1(n4163), .B2(n4162), .A(n4161), .ZN(n4171) );
  XNOR2_X1 U4749 ( .A(n2777), .B(keyinput_202), .ZN(n4170) );
  XNOR2_X1 U4750 ( .A(n4164), .B(keyinput_205), .ZN(n4168) );
  XNOR2_X1 U4751 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_206), .ZN(n4167) );
  XNOR2_X1 U4752 ( .A(IR_REG_20__SCAN_IN), .B(keyinput_203), .ZN(n4166) );
  XNOR2_X1 U4753 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_204), .ZN(n4165) );
  NOR4_X1 U4754 ( .A1(n4168), .A2(n4167), .A3(n4166), .A4(n4165), .ZN(n4169)
         );
  OAI21_X1 U4755 ( .B1(n4171), .B2(n4170), .A(n4169), .ZN(n4189) );
  XNOR2_X1 U4756 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_207), .ZN(n4188) );
  XNOR2_X1 U4757 ( .A(n4172), .B(keyinput_212), .ZN(n4178) );
  XNOR2_X1 U4758 ( .A(n4173), .B(keyinput_215), .ZN(n4177) );
  XNOR2_X1 U4759 ( .A(n4174), .B(keyinput_213), .ZN(n4176) );
  XNOR2_X1 U4760 ( .A(D_REG_1__SCAN_IN), .B(keyinput_216), .ZN(n4175) );
  NOR4_X1 U4761 ( .A1(n4178), .A2(n4177), .A3(n4176), .A4(n4175), .ZN(n4186)
         );
  XOR2_X1 U4762 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_214), .Z(n4185) );
  XOR2_X1 U4763 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_208), .Z(n4184) );
  XNOR2_X1 U4764 ( .A(n2683), .B(keyinput_211), .ZN(n4182) );
  XNOR2_X1 U4765 ( .A(n4179), .B(keyinput_209), .ZN(n4181) );
  XNOR2_X1 U4766 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_210), .ZN(n4180) );
  NOR3_X1 U4767 ( .A1(n4182), .A2(n4181), .A3(n4180), .ZN(n4183) );
  NAND4_X1 U4768 ( .A1(n4186), .A2(n4185), .A3(n4184), .A4(n4183), .ZN(n4187)
         );
  AOI21_X1 U4769 ( .B1(n4189), .B2(n4188), .A(n4187), .ZN(n4196) );
  XNOR2_X1 U4770 ( .A(D_REG_2__SCAN_IN), .B(keyinput_217), .ZN(n4195) );
  XNOR2_X1 U4771 ( .A(D_REG_5__SCAN_IN), .B(keyinput_220), .ZN(n4193) );
  XNOR2_X1 U4772 ( .A(D_REG_3__SCAN_IN), .B(keyinput_218), .ZN(n4192) );
  XNOR2_X1 U4773 ( .A(D_REG_4__SCAN_IN), .B(keyinput_219), .ZN(n4191) );
  XNOR2_X1 U4774 ( .A(D_REG_6__SCAN_IN), .B(keyinput_221), .ZN(n4190) );
  NOR4_X1 U4775 ( .A1(n4193), .A2(n4192), .A3(n4191), .A4(n4190), .ZN(n4194)
         );
  OAI21_X1 U4776 ( .B1(n4196), .B2(n4195), .A(n4194), .ZN(n4199) );
  XNOR2_X1 U4777 ( .A(D_REG_7__SCAN_IN), .B(keyinput_222), .ZN(n4198) );
  XOR2_X1 U4778 ( .A(D_REG_8__SCAN_IN), .B(keyinput_223), .Z(n4197) );
  AOI21_X1 U4779 ( .B1(n4199), .B2(n4198), .A(n4197), .ZN(n4206) );
  XOR2_X1 U4780 ( .A(D_REG_11__SCAN_IN), .B(keyinput_226), .Z(n4202) );
  INV_X1 U4781 ( .A(D_REG_10__SCAN_IN), .ZN(n4936) );
  XNOR2_X1 U4782 ( .A(n4936), .B(keyinput_225), .ZN(n4201) );
  XNOR2_X1 U4783 ( .A(D_REG_9__SCAN_IN), .B(keyinput_224), .ZN(n4200) );
  NAND3_X1 U4784 ( .A1(n4202), .A2(n4201), .A3(n4200), .ZN(n4205) );
  INV_X1 U4785 ( .A(D_REG_13__SCAN_IN), .ZN(n4938) );
  XNOR2_X1 U4786 ( .A(n4938), .B(keyinput_228), .ZN(n4204) );
  XNOR2_X1 U4787 ( .A(D_REG_12__SCAN_IN), .B(keyinput_227), .ZN(n4203) );
  OAI211_X1 U4788 ( .C1(n4206), .C2(n4205), .A(n4204), .B(n4203), .ZN(n4209)
         );
  XOR2_X1 U4789 ( .A(D_REG_14__SCAN_IN), .B(keyinput_229), .Z(n4208) );
  XNOR2_X1 U4790 ( .A(n4940), .B(keyinput_230), .ZN(n4207) );
  AOI21_X1 U4791 ( .B1(n4209), .B2(n4208), .A(n4207), .ZN(n4212) );
  XNOR2_X1 U4792 ( .A(D_REG_17__SCAN_IN), .B(keyinput_232), .ZN(n4211) );
  XNOR2_X1 U4793 ( .A(D_REG_16__SCAN_IN), .B(keyinput_231), .ZN(n4210) );
  NOR3_X1 U4794 ( .A1(n4212), .A2(n4211), .A3(n4210), .ZN(n4215) );
  XNOR2_X1 U4795 ( .A(D_REG_18__SCAN_IN), .B(keyinput_233), .ZN(n4214) );
  XNOR2_X1 U4796 ( .A(D_REG_19__SCAN_IN), .B(keyinput_234), .ZN(n4213) );
  OAI21_X1 U4797 ( .B1(n4215), .B2(n4214), .A(n4213), .ZN(n4219) );
  XNOR2_X1 U4798 ( .A(D_REG_20__SCAN_IN), .B(keyinput_235), .ZN(n4218) );
  XOR2_X1 U4799 ( .A(D_REG_22__SCAN_IN), .B(keyinput_237), .Z(n4217) );
  XNOR2_X1 U4800 ( .A(D_REG_21__SCAN_IN), .B(keyinput_236), .ZN(n4216) );
  AOI211_X1 U4801 ( .C1(n4219), .C2(n4218), .A(n4217), .B(n4216), .ZN(n4222)
         );
  XOR2_X1 U4802 ( .A(D_REG_23__SCAN_IN), .B(keyinput_238), .Z(n4221) );
  XNOR2_X1 U4803 ( .A(D_REG_24__SCAN_IN), .B(keyinput_239), .ZN(n4220) );
  OAI21_X1 U4804 ( .B1(n4222), .B2(n4221), .A(n4220), .ZN(n4225) );
  XNOR2_X1 U4805 ( .A(n4949), .B(keyinput_240), .ZN(n4224) );
  XNOR2_X1 U4806 ( .A(D_REG_26__SCAN_IN), .B(keyinput_241), .ZN(n4223) );
  AOI21_X1 U4807 ( .B1(n4225), .B2(n4224), .A(n4223), .ZN(n4228) );
  INV_X1 U4808 ( .A(D_REG_27__SCAN_IN), .ZN(n4951) );
  XNOR2_X1 U4809 ( .A(n4951), .B(keyinput_242), .ZN(n4227) );
  XNOR2_X1 U4810 ( .A(D_REG_28__SCAN_IN), .B(keyinput_243), .ZN(n4226) );
  NOR3_X1 U4811 ( .A1(n4228), .A2(n4227), .A3(n4226), .ZN(n4231) );
  XNOR2_X1 U4812 ( .A(D_REG_29__SCAN_IN), .B(keyinput_244), .ZN(n4230) );
  XNOR2_X1 U4813 ( .A(D_REG_30__SCAN_IN), .B(keyinput_245), .ZN(n4229) );
  NOR3_X1 U4814 ( .A1(n4231), .A2(n4230), .A3(n4229), .ZN(n4237) );
  INV_X1 U4815 ( .A(D_REG_31__SCAN_IN), .ZN(n4955) );
  XNOR2_X1 U4816 ( .A(n4955), .B(keyinput_246), .ZN(n4236) );
  XOR2_X1 U4817 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_247), .Z(n4234) );
  XOR2_X1 U4818 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_249), .Z(n4233) );
  XNOR2_X1 U4819 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_248), .ZN(n4232) );
  NOR3_X1 U4820 ( .A1(n4234), .A2(n4233), .A3(n4232), .ZN(n4235) );
  OAI21_X1 U4821 ( .B1(n4237), .B2(n4236), .A(n4235), .ZN(n4240) );
  XNOR2_X1 U4822 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_250), .ZN(n4239) );
  XNOR2_X1 U4823 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_251), .ZN(n4238) );
  AOI21_X1 U4824 ( .B1(n4240), .B2(n4239), .A(n4238), .ZN(n4243) );
  XNOR2_X1 U4825 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_252), .ZN(n4242) );
  XNOR2_X1 U4826 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_253), .ZN(n4241) );
  OAI21_X1 U4827 ( .B1(n4243), .B2(n4242), .A(n4241), .ZN(n4246) );
  XOR2_X1 U4828 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_254), .Z(n4245) );
  XOR2_X1 U4829 ( .A(keyinput_127), .B(keyinput_255), .Z(n4244) );
  AOI21_X1 U4830 ( .B1(n4246), .B2(n4245), .A(n4244), .ZN(n4247) );
  AOI211_X1 U4831 ( .C1(n4250), .C2(n4249), .A(n4248), .B(n4247), .ZN(n4251)
         );
  XNOR2_X1 U4832 ( .A(n4252), .B(n4251), .ZN(U3225) );
  NAND2_X1 U4833 ( .A1(n4253), .A2(n4254), .ZN(n4256) );
  XNOR2_X1 U4834 ( .A(n4256), .B(n4255), .ZN(n4264) );
  INV_X1 U4835 ( .A(n4657), .ZN(n4262) );
  AOI22_X1 U4836 ( .A1(n4257), .A2(n5246), .B1(n5258), .B2(n4616), .ZN(n4261)
         );
  NOR2_X1 U4837 ( .A1(n4258), .A2(STATE_REG_SCAN_IN), .ZN(n4259) );
  AOI21_X1 U4838 ( .B1(n5264), .B2(n4471), .A(n4259), .ZN(n4260) );
  OAI211_X1 U4839 ( .C1(n5326), .C2(n4262), .A(n4261), .B(n4260), .ZN(n4263)
         );
  AOI21_X1 U4840 ( .B1(n4264), .B2(n5322), .A(n4263), .ZN(n4265) );
  INV_X1 U4841 ( .A(n4265), .ZN(U3226) );
  OAI21_X1 U4842 ( .B1(n4267), .B2(n4266), .A(n3775), .ZN(n4272) );
  AOI22_X1 U4843 ( .A1(n5119), .A2(n5246), .B1(n5264), .B2(n4480), .ZN(n4270)
         );
  AOI21_X1 U4844 ( .B1(n5258), .B2(n4478), .A(n4268), .ZN(n4269) );
  OAI211_X1 U4845 ( .C1(n5326), .C2(n5132), .A(n4270), .B(n4269), .ZN(n4271)
         );
  AOI21_X1 U4846 ( .B1(n4272), .B2(n5322), .A(n4271), .ZN(n4273) );
  INV_X1 U4847 ( .A(n4273), .ZN(U3228) );
  OAI21_X1 U4848 ( .B1(n4276), .B2(n4275), .A(n4274), .ZN(n4277) );
  NAND2_X1 U4849 ( .A1(n4277), .A2(n5322), .ZN(n4284) );
  OR2_X1 U4850 ( .A1(n4792), .A2(n5107), .ZN(n4279) );
  OR2_X1 U4851 ( .A1(n4849), .A2(n5286), .ZN(n4278) );
  NAND2_X1 U4852 ( .A1(n4279), .A2(n4278), .ZN(n5158) );
  AOI22_X1 U4853 ( .A1(n5158), .A2(n5243), .B1(REG3_REG_13__SCAN_IN), .B2(
        U3149), .ZN(n4283) );
  OR2_X1 U4854 ( .A1(n5326), .A2(n4280), .ZN(n4282) );
  NAND2_X1 U4855 ( .A1(n5267), .A2(n5163), .ZN(n4281) );
  NAND4_X1 U4856 ( .A1(n4284), .A2(n4283), .A3(n4282), .A4(n4281), .ZN(U3231)
         );
  AOI21_X1 U4857 ( .B1(n4287), .B2(n4285), .A(n4286), .ZN(n4295) );
  INV_X1 U4858 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4288) );
  OAI22_X1 U4859 ( .A1(n5315), .A2(n4289), .B1(STATE_REG_SCAN_IN), .B2(n4288), 
        .ZN(n4292) );
  OAI22_X1 U4860 ( .A1(n5319), .A2(n4290), .B1(n5317), .B2(n4692), .ZN(n4291)
         );
  AOI211_X1 U4861 ( .C1(n4293), .C2(n4301), .A(n4292), .B(n4291), .ZN(n4294)
         );
  OAI21_X1 U4862 ( .B1(n4295), .B2(n5226), .A(n4294), .ZN(U3232) );
  INV_X1 U4863 ( .A(n3814), .ZN(n4296) );
  AOI21_X1 U4864 ( .B1(n4298), .B2(n4297), .A(n4296), .ZN(n4304) );
  OAI22_X1 U4865 ( .A1(n5319), .A2(n4858), .B1(n5315), .B2(n5108), .ZN(n4299)
         );
  AOI211_X1 U4866 ( .C1(n5258), .C2(n4476), .A(n4300), .B(n4299), .ZN(n4303)
         );
  NAND2_X1 U4867 ( .A1(n4301), .A2(n4860), .ZN(n4302) );
  OAI211_X1 U4868 ( .C1(n4304), .C2(n5226), .A(n4303), .B(n4302), .ZN(U3233)
         );
  INV_X1 U4869 ( .A(n4305), .ZN(n4307) );
  NOR2_X1 U4870 ( .A1(n4307), .A2(n4306), .ZN(n4308) );
  XNOR2_X1 U4871 ( .A(n4309), .B(n4308), .ZN(n4316) );
  INV_X1 U4872 ( .A(n4624), .ZN(n4314) );
  AOI22_X1 U4873 ( .A1(n4621), .A2(n5246), .B1(n5258), .B2(n4470), .ZN(n4313)
         );
  NOR2_X1 U4874 ( .A1(n4310), .A2(STATE_REG_SCAN_IN), .ZN(n4311) );
  AOI21_X1 U4875 ( .B1(n5264), .B2(n4616), .A(n4311), .ZN(n4312) );
  OAI211_X1 U4876 ( .C1(n5326), .C2(n4314), .A(n4313), .B(n4312), .ZN(n4315)
         );
  AOI21_X1 U4877 ( .B1(n4316), .B2(n5322), .A(n4315), .ZN(n4317) );
  INV_X1 U4878 ( .A(n4317), .ZN(U3237) );
  NAND2_X1 U4879 ( .A1(n4319), .A2(n4318), .ZN(n4360) );
  NAND2_X1 U4880 ( .A1(n4774), .A2(n5193), .ZN(n4322) );
  AND2_X1 U4881 ( .A1(n4360), .A2(n4322), .ZN(n4432) );
  NAND2_X1 U4882 ( .A1(n4321), .A2(n4320), .ZN(n4338) );
  AND2_X1 U4883 ( .A1(n4323), .A2(n4322), .ZN(n4433) );
  NAND2_X1 U4884 ( .A1(n4433), .A2(n4324), .ZN(n4337) );
  INV_X1 U4885 ( .A(n4325), .ZN(n4327) );
  NAND2_X1 U4886 ( .A1(n4327), .A2(n4326), .ZN(n4352) );
  INV_X1 U4887 ( .A(n4352), .ZN(n4330) );
  INV_X1 U4888 ( .A(n4328), .ZN(n4329) );
  NAND4_X1 U4889 ( .A1(n4330), .A2(n4329), .A3(n4358), .A4(n4348), .ZN(n4335)
         );
  AND2_X1 U4890 ( .A1(n4332), .A2(n4331), .ZN(n4333) );
  NAND2_X1 U4891 ( .A1(n4339), .A2(n4333), .ZN(n4359) );
  AOI21_X1 U4892 ( .B1(n4335), .B2(n4334), .A(n4359), .ZN(n4336) );
  AOI211_X1 U4893 ( .C1(n4339), .C2(n4338), .A(n4337), .B(n4336), .ZN(n4363)
         );
  NAND2_X1 U4894 ( .A1(n3418), .A2(n4340), .ZN(n4400) );
  OAI211_X1 U4895 ( .C1(n4342), .C2(n4915), .A(n4400), .B(n4341), .ZN(n4344)
         );
  NAND3_X1 U4896 ( .A1(n4344), .A2(n5050), .A3(n4343), .ZN(n4346) );
  NAND3_X1 U4897 ( .A1(n4346), .A2(n4345), .A3(n4397), .ZN(n4347) );
  NAND3_X1 U4898 ( .A1(n4347), .A2(n2768), .A3(n4398), .ZN(n4351) );
  NAND4_X1 U4899 ( .A1(n4351), .A2(n4350), .A3(n4349), .A4(n4348), .ZN(n4354)
         );
  AOI21_X1 U4900 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(n4357) );
  INV_X1 U4901 ( .A(n4355), .ZN(n4356) );
  NOR3_X1 U4902 ( .A1(n4357), .A2(n5111), .A3(n4356), .ZN(n4361) );
  INV_X1 U4903 ( .A(n4358), .ZN(n5110) );
  OR4_X1 U4904 ( .A1(n4361), .A2(n5110), .A3(n4360), .A4(n4359), .ZN(n4362) );
  OAI21_X1 U4905 ( .B1(n4432), .B2(n4363), .A(n4362), .ZN(n4367) );
  NOR3_X1 U4906 ( .A1(n4366), .A2(n4365), .A3(n4364), .ZN(n4435) );
  OAI21_X1 U4907 ( .B1(n4436), .B2(n4367), .A(n4435), .ZN(n4368) );
  AOI21_X1 U4908 ( .B1(n4439), .B2(n4368), .A(n4438), .ZN(n4371) );
  NOR2_X1 U4909 ( .A1(n4370), .A2(n4369), .ZN(n4441) );
  AOI221_X1 U4910 ( .B1(n4371), .B2(n4441), .C1(n4442), .C2(n4441), .A(n4444), 
        .ZN(n4390) );
  INV_X1 U4911 ( .A(n4376), .ZN(n4467) );
  AOI22_X1 U4912 ( .A1(n4467), .A2(n5330), .B1(n4453), .B2(n4456), .ZN(n4430)
         );
  NAND2_X1 U4913 ( .A1(n4468), .A2(n4372), .ZN(n4373) );
  AND2_X1 U4914 ( .A1(n4374), .A2(n4373), .ZN(n4445) );
  NAND4_X1 U4915 ( .A1(n4430), .A2(n4445), .A3(n4600), .A4(n4375), .ZN(n4389)
         );
  NOR2_X1 U4916 ( .A1(n4453), .A2(n4456), .ZN(n4387) );
  AND2_X1 U4917 ( .A1(n4376), .A2(n4452), .ZN(n4377) );
  OR2_X1 U4918 ( .A1(n4387), .A2(n4377), .ZN(n4417) );
  INV_X1 U4919 ( .A(n4417), .ZN(n4381) );
  INV_X1 U4920 ( .A(n4468), .ZN(n4379) );
  NAND2_X1 U4921 ( .A1(n4379), .A2(n4378), .ZN(n4380) );
  NAND2_X1 U4922 ( .A1(n4381), .A2(n4380), .ZN(n4386) );
  NAND2_X1 U4923 ( .A1(n4383), .A2(n4382), .ZN(n4384) );
  AND2_X1 U4924 ( .A1(n4384), .A2(n4445), .ZN(n4385) );
  OR2_X1 U4925 ( .A1(n4386), .A2(n4385), .ZN(n4451) );
  OAI21_X1 U4926 ( .B1(n4387), .B2(n4430), .A(n4451), .ZN(n4388) );
  OAI21_X1 U4927 ( .B1(n4390), .B2(n4389), .A(n4388), .ZN(n4460) );
  INV_X1 U4928 ( .A(n4391), .ZN(n4799) );
  NOR4_X1 U4929 ( .A1(n3633), .A2(n2765), .A3(n4392), .A4(n4722), .ZN(n4406)
         );
  INV_X1 U4930 ( .A(n4844), .ZN(n4854) );
  NOR4_X1 U4931 ( .A1(n4854), .A2(n2681), .A3(n4826), .A4(n4394), .ZN(n4405)
         );
  NOR4_X1 U4932 ( .A1(n4396), .A2(n4815), .A3(n4395), .A4(n3419), .ZN(n4404)
         );
  INV_X1 U4933 ( .A(n5058), .ZN(n4402) );
  NAND2_X1 U4934 ( .A1(n4400), .A2(n4399), .ZN(n5016) );
  NOR4_X1 U4935 ( .A1(n4402), .A2(n5016), .A3(n4739), .A4(n4401), .ZN(n4403)
         );
  NAND4_X1 U4936 ( .A1(n4406), .A2(n4405), .A3(n4404), .A4(n4403), .ZN(n4429)
         );
  INV_X1 U4937 ( .A(n4407), .ZN(n4409) );
  OR2_X1 U4938 ( .A1(n4409), .A2(n4408), .ZN(n4631) );
  INV_X1 U4939 ( .A(n4410), .ZN(n4411) );
  NAND4_X1 U4940 ( .A1(n4631), .A2(n5280), .A3(n4411), .A4(n4430), .ZN(n4412)
         );
  NOR3_X1 U4941 ( .A1(n4412), .A2(n4803), .A3(n4782), .ZN(n4425) );
  INV_X1 U4942 ( .A(n4686), .ZN(n4683) );
  NAND2_X1 U4943 ( .A1(n4414), .A2(n4413), .ZN(n4649) );
  INV_X1 U4944 ( .A(n4687), .ZN(n4416) );
  NOR4_X1 U4945 ( .A1(n4683), .A2(n4649), .A3(n4417), .A4(n4701), .ZN(n4424)
         );
  INV_X1 U4946 ( .A(n4599), .ZN(n4422) );
  AND2_X1 U4947 ( .A1(n4419), .A2(n4418), .ZN(n5113) );
  NAND2_X1 U4948 ( .A1(n4600), .A2(n4420), .ZN(n4614) );
  NOR4_X1 U4949 ( .A1(n4422), .A2(n4421), .A3(n5113), .A4(n4614), .ZN(n4423)
         );
  NAND3_X1 U4950 ( .A1(n4425), .A2(n4424), .A3(n4423), .ZN(n4428) );
  INV_X1 U4951 ( .A(n4426), .ZN(n4427) );
  NOR4_X1 U4952 ( .A1(n4429), .A2(n4428), .A3(n4427), .A4(n4676), .ZN(n4458)
         );
  INV_X1 U4953 ( .A(n4430), .ZN(n4455) );
  INV_X1 U4954 ( .A(n4431), .ZN(n4434) );
  AOI21_X1 U4955 ( .B1(n4434), .B2(n4433), .A(n4432), .ZN(n4437) );
  OAI21_X1 U4956 ( .B1(n4437), .B2(n4436), .A(n4435), .ZN(n4440) );
  AOI21_X1 U4957 ( .B1(n4440), .B2(n4439), .A(n4438), .ZN(n4443) );
  OAI21_X1 U4958 ( .B1(n4443), .B2(n4442), .A(n4441), .ZN(n4449) );
  INV_X1 U4959 ( .A(n4444), .ZN(n4448) );
  INV_X1 U4960 ( .A(n4445), .ZN(n4447) );
  AOI211_X1 U4961 ( .C1(n4449), .C2(n4448), .A(n4447), .B(n4446), .ZN(n4450)
         );
  AOI211_X1 U4962 ( .C1(n4453), .C2(n4452), .A(n4451), .B(n4450), .ZN(n4454)
         );
  AOI21_X1 U4963 ( .B1(n4456), .B2(n4455), .A(n4454), .ZN(n4457) );
  MUX2_X1 U4964 ( .A(n4458), .B(n4457), .S(n4915), .Z(n4459) );
  MUX2_X1 U4965 ( .A(n4460), .B(n4459), .S(n4916), .Z(n4461) );
  XNOR2_X1 U4966 ( .A(n4461), .B(n5173), .ZN(n4466) );
  NAND3_X1 U4967 ( .A1(n4462), .A2(n4979), .A3(n5054), .ZN(n4463) );
  OAI211_X1 U4968 ( .C1(n4914), .C2(n4465), .A(n4463), .B(B_REG_SCAN_IN), .ZN(
        n4464) );
  OAI21_X1 U4969 ( .B1(n4466), .B2(n4465), .A(n4464), .ZN(U3239) );
  MUX2_X1 U4970 ( .A(DATAO_REG_30__SCAN_IN), .B(n4467), .S(n4481), .Z(U3580)
         );
  MUX2_X1 U4971 ( .A(n4468), .B(DATAO_REG_29__SCAN_IN), .S(n4485), .Z(U3579)
         );
  MUX2_X1 U4972 ( .A(DATAO_REG_28__SCAN_IN), .B(n4469), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4973 ( .A(n4470), .B(DATAO_REG_27__SCAN_IN), .S(n4485), .Z(U3577)
         );
  MUX2_X1 U4974 ( .A(DATAO_REG_26__SCAN_IN), .B(n4604), .S(n4481), .Z(U3576)
         );
  MUX2_X1 U4975 ( .A(DATAO_REG_25__SCAN_IN), .B(n4616), .S(n4481), .Z(U3575)
         );
  MUX2_X1 U4976 ( .A(n4668), .B(DATAO_REG_24__SCAN_IN), .S(n4485), .Z(U3574)
         );
  MUX2_X1 U4977 ( .A(DATAO_REG_23__SCAN_IN), .B(n4471), .S(n4481), .Z(U3573)
         );
  MUX2_X1 U4978 ( .A(DATAO_REG_22__SCAN_IN), .B(n4710), .S(n4481), .Z(U3572)
         );
  MUX2_X1 U4979 ( .A(n5284), .B(DATAO_REG_21__SCAN_IN), .S(n4485), .Z(U3571)
         );
  MUX2_X1 U4980 ( .A(n5312), .B(DATAO_REG_20__SCAN_IN), .S(n4485), .Z(U3570)
         );
  MUX2_X1 U4981 ( .A(n5265), .B(DATAO_REG_19__SCAN_IN), .S(n4485), .Z(U3569)
         );
  MUX2_X1 U4982 ( .A(n4724), .B(DATAO_REG_18__SCAN_IN), .S(n4485), .Z(U3568)
         );
  MUX2_X1 U4983 ( .A(DATAO_REG_17__SCAN_IN), .B(n4472), .S(n4481), .Z(U3567)
         );
  MUX2_X1 U4984 ( .A(n4756), .B(DATAO_REG_16__SCAN_IN), .S(n4485), .Z(U3566)
         );
  MUX2_X1 U4985 ( .A(DATAO_REG_15__SCAN_IN), .B(n4473), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4986 ( .A(DATAO_REG_14__SCAN_IN), .B(n4474), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4987 ( .A(n4475), .B(DATAO_REG_13__SCAN_IN), .S(n4485), .Z(U3563)
         );
  MUX2_X1 U4988 ( .A(DATAO_REG_12__SCAN_IN), .B(n4476), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4989 ( .A(DATAO_REG_11__SCAN_IN), .B(n4477), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4990 ( .A(DATAO_REG_10__SCAN_IN), .B(n4478), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4991 ( .A(n4479), .B(DATAO_REG_9__SCAN_IN), .S(n4485), .Z(U3559) );
  MUX2_X1 U4992 ( .A(n4480), .B(DATAO_REG_8__SCAN_IN), .S(n4485), .Z(U3558) );
  MUX2_X1 U4993 ( .A(DATAO_REG_7__SCAN_IN), .B(n4482), .S(n4481), .Z(U3557) );
  MUX2_X1 U4994 ( .A(n4483), .B(DATAO_REG_6__SCAN_IN), .S(n4485), .Z(U3556) );
  MUX2_X1 U4995 ( .A(DATAO_REG_5__SCAN_IN), .B(n4484), .S(U4043), .Z(U3555) );
  MUX2_X1 U4996 ( .A(n5053), .B(DATAO_REG_4__SCAN_IN), .S(n4485), .Z(U3554) );
  MUX2_X1 U4997 ( .A(DATAO_REG_3__SCAN_IN), .B(n4486), .S(n4481), .Z(U3553) );
  MUX2_X1 U4998 ( .A(DATAO_REG_2__SCAN_IN), .B(n3471), .S(n4481), .Z(U3552) );
  MUX2_X1 U4999 ( .A(DATAO_REG_1__SCAN_IN), .B(n3417), .S(U4043), .Z(U3551) );
  MUX2_X1 U5000 ( .A(DATAO_REG_0__SCAN_IN), .B(n3418), .S(n4481), .Z(U3550) );
  NAND2_X1 U5001 ( .A1(n4922), .A2(n4487), .ZN(n4489) );
  INV_X1 U5002 ( .A(n4507), .ZN(n4921) );
  INV_X1 U5003 ( .A(REG1_REG_13__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U5004 ( .A1(n4507), .A2(n5169), .ZN(n4491) );
  INV_X1 U5005 ( .A(n4491), .ZN(n4490) );
  AOI21_X1 U5006 ( .B1(REG1_REG_13__SCAN_IN), .B2(n4921), .A(n4490), .ZN(n4492) );
  NAND2_X1 U5007 ( .A1(n4921), .A2(REG1_REG_13__SCAN_IN), .ZN(n4512) );
  OAI211_X1 U5008 ( .C1(n4493), .C2(n4492), .A(n4511), .B(n5010), .ZN(n4506)
         );
  NOR2_X1 U5009 ( .A1(n4495), .A2(n4494), .ZN(n4496) );
  INV_X1 U5010 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4498) );
  OR2_X1 U5011 ( .A1(n4507), .A2(n4498), .ZN(n4508) );
  NAND2_X1 U5012 ( .A1(n4507), .A2(n4498), .ZN(n4499) );
  NAND2_X1 U5013 ( .A1(n4508), .A2(n4499), .ZN(n4500) );
  AOI211_X1 U5014 ( .C1(n4501), .C2(n4500), .A(n2543), .B(n4968), .ZN(n4504)
         );
  INV_X1 U5015 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4502) );
  NOR2_X1 U5016 ( .A1(STATE_REG_SCAN_IN), .A2(n4502), .ZN(n4503) );
  AOI211_X1 U5017 ( .C1(n4998), .C2(ADDR_REG_13__SCAN_IN), .A(n4504), .B(n4503), .ZN(n4505) );
  OAI211_X1 U5018 ( .C1(n4591), .C2(n4507), .A(n4506), .B(n4505), .ZN(U3253)
         );
  INV_X1 U5019 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4510) );
  AOI211_X1 U5020 ( .C1(n4510), .C2(n4509), .A(n4523), .B(n4968), .ZN(n4519)
         );
  NAND2_X1 U5021 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4513), .ZN(n4528) );
  OAI211_X1 U5022 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4513), .A(n5010), .B(n4528), .ZN(n4517) );
  NOR2_X1 U5023 ( .A1(STATE_REG_SCAN_IN), .A2(n4514), .ZN(n4515) );
  AOI21_X1 U5024 ( .B1(n4998), .B2(ADDR_REG_14__SCAN_IN), .A(n4515), .ZN(n4516) );
  OAI211_X1 U5025 ( .C1(n4591), .C2(n4521), .A(n4517), .B(n4516), .ZN(n4518)
         );
  OR2_X1 U5026 ( .A1(n4519), .A2(n4518), .ZN(U3254) );
  INV_X1 U5027 ( .A(n4520), .ZN(n4522) );
  NOR2_X1 U5028 ( .A1(n4522), .A2(n4521), .ZN(n4524) );
  NAND2_X1 U5029 ( .A1(n4919), .A2(REG2_REG_15__SCAN_IN), .ZN(n4525) );
  OAI21_X1 U5030 ( .B1(n4919), .B2(REG2_REG_15__SCAN_IN), .A(n4525), .ZN(n4526) );
  AOI211_X1 U5031 ( .C1(n2547), .C2(n4526), .A(n4542), .B(n4968), .ZN(n4538)
         );
  NAND2_X1 U5032 ( .A1(n4920), .A2(n4527), .ZN(n4529) );
  NAND2_X1 U5033 ( .A1(n4529), .A2(n4528), .ZN(n4532) );
  INV_X1 U5034 ( .A(REG1_REG_15__SCAN_IN), .ZN(n5201) );
  NAND2_X1 U5035 ( .A1(n4919), .A2(REG1_REG_15__SCAN_IN), .ZN(n4540) );
  INV_X1 U5036 ( .A(n4540), .ZN(n4530) );
  AOI21_X1 U5037 ( .B1(n5201), .B2(n4536), .A(n4530), .ZN(n4531) );
  OAI211_X1 U5038 ( .C1(n4532), .C2(n4531), .A(n5010), .B(n4539), .ZN(n4535)
         );
  AND2_X1 U5039 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4533) );
  AOI21_X1 U5040 ( .B1(n4998), .B2(ADDR_REG_15__SCAN_IN), .A(n4533), .ZN(n4534) );
  OAI211_X1 U5041 ( .C1(n4591), .C2(n4536), .A(n4535), .B(n4534), .ZN(n4537)
         );
  OR2_X1 U5042 ( .A1(n4538), .A2(n4537), .ZN(U3255) );
  AOI21_X1 U5043 ( .B1(n4541), .B2(REG1_REG_16__SCAN_IN), .A(n4559), .ZN(n4551) );
  INV_X1 U5044 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4543) );
  AOI221_X1 U5045 ( .B1(n4544), .B2(n4555), .C1(n4543), .C2(n4555), .A(n4968), 
        .ZN(n4545) );
  INV_X1 U5046 ( .A(n4545), .ZN(n4549) );
  NOR2_X1 U5047 ( .A1(n4591), .A2(n4552), .ZN(n4546) );
  AOI211_X1 U5048 ( .C1(n4998), .C2(ADDR_REG_16__SCAN_IN), .A(n4547), .B(n4546), .ZN(n4548) );
  OAI211_X1 U5049 ( .C1(n4551), .C2(n4550), .A(n4549), .B(n4548), .ZN(U3256)
         );
  INV_X1 U5050 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4765) );
  AOI22_X1 U5051 ( .A1(n4570), .A2(n4765), .B1(REG2_REG_17__SCAN_IN), .B2(
        n5213), .ZN(n4557) );
  NAND2_X1 U5052 ( .A1(n4553), .A2(n4552), .ZN(n4554) );
  AOI211_X1 U5053 ( .C1(n4557), .C2(n4556), .A(n4569), .B(n4968), .ZN(n4568)
         );
  NOR2_X1 U5054 ( .A1(n4918), .A2(n4558), .ZN(n4560) );
  INV_X1 U5055 ( .A(REG1_REG_17__SCAN_IN), .ZN(n5217) );
  NOR2_X1 U5056 ( .A1(n5213), .A2(n5217), .ZN(n4561) );
  AOI21_X1 U5057 ( .B1(n5217), .B2(n5213), .A(n4561), .ZN(n4562) );
  NAND2_X1 U5058 ( .A1(n4562), .A2(n4563), .ZN(n4574) );
  OAI211_X1 U5059 ( .C1(n4563), .C2(n4562), .A(n4574), .B(n5010), .ZN(n4566)
         );
  AOI21_X1 U5060 ( .B1(n4998), .B2(ADDR_REG_17__SCAN_IN), .A(n4564), .ZN(n4565) );
  OAI211_X1 U5061 ( .C1(n4591), .C2(n5213), .A(n4566), .B(n4565), .ZN(n4567)
         );
  OR2_X1 U5062 ( .A1(n4568), .A2(n4567), .ZN(U3257) );
  INV_X1 U5063 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4571) );
  AOI22_X1 U5064 ( .A1(n4917), .A2(n4571), .B1(REG2_REG_18__SCAN_IN), .B2(
        n4581), .ZN(n4572) );
  AOI211_X1 U5065 ( .C1(n2528), .C2(n4572), .A(n4584), .B(n4968), .ZN(n4583)
         );
  NOR2_X1 U5066 ( .A1(n4917), .A2(REG1_REG_18__SCAN_IN), .ZN(n4573) );
  AOI21_X1 U5067 ( .B1(REG1_REG_18__SCAN_IN), .B2(n4917), .A(n4573), .ZN(n4576) );
  OAI21_X1 U5068 ( .B1(n5213), .B2(n5217), .A(n4574), .ZN(n4575) );
  OAI211_X1 U5069 ( .C1(n4576), .C2(n4575), .A(n5010), .B(n4587), .ZN(n4580)
         );
  NOR2_X1 U5070 ( .A1(STATE_REG_SCAN_IN), .A2(n4577), .ZN(n4578) );
  AOI21_X1 U5071 ( .B1(n4998), .B2(ADDR_REG_18__SCAN_IN), .A(n4578), .ZN(n4579) );
  OAI211_X1 U5072 ( .C1(n4591), .C2(n4581), .A(n4580), .B(n4579), .ZN(n4582)
         );
  OR2_X1 U5073 ( .A1(n4583), .A2(n4582), .ZN(U3258) );
  INV_X1 U5074 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4585) );
  MUX2_X1 U5075 ( .A(REG2_REG_19__SCAN_IN), .B(n4585), .S(n4592), .Z(n4586) );
  INV_X1 U5076 ( .A(n4968), .ZN(n5005) );
  INV_X1 U5077 ( .A(REG1_REG_19__SCAN_IN), .ZN(n5255) );
  MUX2_X1 U5078 ( .A(n5255), .B(REG1_REG_19__SCAN_IN), .S(n4592), .Z(n4588) );
  AOI22_X1 U5079 ( .A1(n4998), .A2(ADDR_REG_19__SCAN_IN), .B1(
        REG3_REG_19__SCAN_IN), .B2(U3149), .ZN(n4590) );
  XNOR2_X1 U5080 ( .A(n4593), .B(n4599), .ZN(n4878) );
  AOI21_X1 U5081 ( .B1(n4603), .B2(n4622), .A(n4594), .ZN(n4876) );
  INV_X1 U5082 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4597) );
  INV_X1 U5083 ( .A(n4595), .ZN(n4596) );
  OAI22_X1 U5084 ( .A1(n5305), .A2(n4597), .B1(n4596), .B2(n5300), .ZN(n4598)
         );
  AOI21_X1 U5085 ( .B1(n4876), .B2(n5344), .A(n4598), .ZN(n4609) );
  AOI21_X1 U5086 ( .B1(n2531), .B2(n4600), .A(n4599), .ZN(n4602) );
  OAI21_X1 U5087 ( .B1(n4602), .B2(n4601), .A(n5289), .ZN(n4606) );
  AOI22_X1 U5088 ( .A1(n4604), .A2(n5054), .B1(n4603), .B2(n5282), .ZN(n4605)
         );
  OAI211_X1 U5089 ( .C1(n4607), .C2(n5107), .A(n4606), .B(n4605), .ZN(n4875)
         );
  NAND2_X1 U5090 ( .A1(n4875), .A2(n5305), .ZN(n4608) );
  OAI211_X1 U5091 ( .C1(n4878), .C2(n4841), .A(n4609), .B(n4608), .ZN(U3263)
         );
  XNOR2_X1 U5092 ( .A(n4610), .B(n4614), .ZN(n4881) );
  INV_X1 U5093 ( .A(n4611), .ZN(n4612) );
  NOR2_X1 U5094 ( .A1(n4613), .A2(n4612), .ZN(n4615) );
  XNOR2_X1 U5095 ( .A(n4615), .B(n4614), .ZN(n4620) );
  AOI22_X1 U5096 ( .A1(n4616), .A2(n5054), .B1(n4621), .B2(n5282), .ZN(n4617)
         );
  OAI21_X1 U5097 ( .B1(n4618), .B2(n5107), .A(n4617), .ZN(n4619) );
  AOI21_X1 U5098 ( .B1(n4620), .B2(n5289), .A(n4619), .ZN(n4880) );
  INV_X1 U5099 ( .A(n4880), .ZN(n4627) );
  AOI21_X1 U5100 ( .B1(n4637), .B2(n4621), .A(n5291), .ZN(n4623) );
  NAND2_X1 U5101 ( .A1(n4623), .A2(n4622), .ZN(n4879) );
  AOI22_X1 U5102 ( .A1(n5348), .A2(REG2_REG_26__SCAN_IN), .B1(n4624), .B2(
        n5178), .ZN(n4625) );
  OAI21_X1 U5103 ( .B1(n4879), .B2(n4733), .A(n4625), .ZN(n4626) );
  AOI21_X1 U5104 ( .B1(n4627), .B2(n5305), .A(n4626), .ZN(n4628) );
  OAI21_X1 U5105 ( .B1(n4881), .B2(n4841), .A(n4628), .ZN(U3264) );
  XNOR2_X1 U5106 ( .A(n4629), .B(n4631), .ZN(n4884) );
  XOR2_X1 U5107 ( .A(n4631), .B(n4630), .Z(n4636) );
  AOI22_X1 U5108 ( .A1(n4668), .A2(n5054), .B1(n4632), .B2(n5282), .ZN(n4633)
         );
  OAI21_X1 U5109 ( .B1(n4634), .B2(n5107), .A(n4633), .ZN(n4635) );
  AOI21_X1 U5110 ( .B1(n4636), .B2(n5289), .A(n4635), .ZN(n4883) );
  INV_X1 U5111 ( .A(n4883), .ZN(n4643) );
  INV_X1 U5112 ( .A(n4655), .ZN(n4639) );
  OAI211_X1 U5113 ( .C1(n4639), .C2(n4638), .A(n5335), .B(n4637), .ZN(n4882)
         );
  AOI22_X1 U5114 ( .A1(n5348), .A2(REG2_REG_25__SCAN_IN), .B1(n4640), .B2(
        n5178), .ZN(n4641) );
  OAI21_X1 U5115 ( .B1(n4882), .B2(n4733), .A(n4641), .ZN(n4642) );
  AOI21_X1 U5116 ( .B1(n4643), .B2(n5305), .A(n4642), .ZN(n4644) );
  OAI21_X1 U5117 ( .B1(n4884), .B2(n4841), .A(n4644), .ZN(U3265) );
  XNOR2_X1 U5118 ( .A(n4645), .B(n4649), .ZN(n4887) );
  INV_X1 U5119 ( .A(n4646), .ZN(n4647) );
  NOR2_X1 U5120 ( .A1(n4648), .A2(n4647), .ZN(n4650) );
  XNOR2_X1 U5121 ( .A(n4650), .B(n4649), .ZN(n4654) );
  NOR2_X1 U5122 ( .A1(n4651), .A2(n5107), .ZN(n4653) );
  OAI22_X1 U5123 ( .A1(n4692), .A2(n5286), .B1(n4656), .B2(n5327), .ZN(n4652)
         );
  AOI211_X1 U5124 ( .C1(n4654), .C2(n5289), .A(n4653), .B(n4652), .ZN(n4886)
         );
  INV_X1 U5125 ( .A(n4886), .ZN(n4660) );
  OAI211_X1 U5126 ( .C1(n4669), .C2(n4656), .A(n5335), .B(n4655), .ZN(n4885)
         );
  AOI22_X1 U5127 ( .A1(n5348), .A2(REG2_REG_24__SCAN_IN), .B1(n4657), .B2(
        n5178), .ZN(n4658) );
  OAI21_X1 U5128 ( .B1(n4885), .B2(n4733), .A(n4658), .ZN(n4659) );
  AOI21_X1 U5129 ( .B1(n4660), .B2(n5305), .A(n4659), .ZN(n4661) );
  OAI21_X1 U5130 ( .B1(n4841), .B2(n4887), .A(n4661), .ZN(U3266) );
  OAI22_X1 U5131 ( .A1(n5316), .A2(n5286), .B1(n5327), .B2(n4671), .ZN(n4667)
         );
  INV_X1 U5132 ( .A(n4701), .ZN(n4704) );
  INV_X1 U5133 ( .A(n4662), .ZN(n4705) );
  NAND3_X1 U5134 ( .A1(n5278), .A2(n4704), .A3(n4705), .ZN(n4703) );
  NAND3_X1 U5135 ( .A1(n4703), .A2(n4686), .A3(n4687), .ZN(n4685) );
  NAND2_X1 U5136 ( .A1(n4685), .A2(n4663), .ZN(n4664) );
  XNOR2_X1 U5137 ( .A(n4664), .B(n4676), .ZN(n4665) );
  NOR2_X1 U5138 ( .A1(n4665), .A2(n5115), .ZN(n4666) );
  AOI211_X1 U5139 ( .C1(n5283), .C2(n4668), .A(n4667), .B(n4666), .ZN(n4890)
         );
  INV_X1 U5140 ( .A(n4669), .ZN(n4670) );
  OAI21_X1 U5141 ( .B1(n4693), .B2(n4671), .A(n4670), .ZN(n4891) );
  INV_X1 U5142 ( .A(n4891), .ZN(n4675) );
  INV_X1 U5143 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4673) );
  OAI22_X1 U5144 ( .A1(n5305), .A2(n4673), .B1(n4672), .B2(n5300), .ZN(n4674)
         );
  AOI21_X1 U5145 ( .B1(n4675), .B2(n5344), .A(n4674), .ZN(n4680) );
  OR2_X1 U5146 ( .A1(n4677), .A2(n4676), .ZN(n4888) );
  NAND3_X1 U5147 ( .A1(n4888), .A2(n4863), .A3(n4678), .ZN(n4679) );
  OAI211_X1 U5148 ( .C1(n4890), .C2(n5348), .A(n4680), .B(n4679), .ZN(U3267)
         );
  INV_X1 U5149 ( .A(n4681), .ZN(n4684) );
  OAI21_X1 U5150 ( .B1(n4684), .B2(n4683), .A(n4682), .ZN(n4895) );
  INV_X1 U5151 ( .A(n4685), .ZN(n4689) );
  AOI21_X1 U5152 ( .B1(n4703), .B2(n4687), .A(n4686), .ZN(n4688) );
  OAI21_X1 U5153 ( .B1(n4689), .B2(n4688), .A(n5289), .ZN(n4691) );
  AOI22_X1 U5154 ( .A1(n5284), .A2(n5054), .B1(n4694), .B2(n5282), .ZN(n4690)
         );
  OAI211_X1 U5155 ( .C1(n4692), .C2(n5107), .A(n4691), .B(n4690), .ZN(n4892)
         );
  NAND2_X1 U5156 ( .A1(n4892), .A2(n5305), .ZN(n4699) );
  AOI21_X1 U5157 ( .B1(n4694), .B2(n4712), .A(n4693), .ZN(n4893) );
  INV_X1 U5158 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4696) );
  OAI22_X1 U5159 ( .A1(n5305), .A2(n4696), .B1(n4695), .B2(n5300), .ZN(n4697)
         );
  AOI21_X1 U5160 ( .B1(n4893), .B2(n5344), .A(n4697), .ZN(n4698) );
  OAI211_X1 U5161 ( .C1(n4895), .C2(n4841), .A(n4699), .B(n4698), .ZN(U3268)
         );
  XNOR2_X1 U5162 ( .A(n4700), .B(n4701), .ZN(n4898) );
  NAND2_X1 U5163 ( .A1(n5312), .A2(n5054), .ZN(n4702) );
  OAI21_X1 U5164 ( .B1(n5327), .B2(n5318), .A(n4702), .ZN(n4709) );
  INV_X1 U5165 ( .A(n4703), .ZN(n4707) );
  AOI21_X1 U5166 ( .B1(n5278), .B2(n4705), .A(n4704), .ZN(n4706) );
  NOR3_X1 U5167 ( .A1(n4707), .A2(n4706), .A3(n5115), .ZN(n4708) );
  AOI211_X1 U5168 ( .C1(n5283), .C2(n4710), .A(n4709), .B(n4708), .ZN(n4897)
         );
  INV_X1 U5169 ( .A(n4897), .ZN(n4717) );
  AOI21_X1 U5170 ( .B1(n5275), .B2(n4711), .A(n5291), .ZN(n4713) );
  NAND2_X1 U5171 ( .A1(n4713), .A2(n4712), .ZN(n4896) );
  AOI22_X1 U5172 ( .A1(n5348), .A2(REG2_REG_21__SCAN_IN), .B1(n4714), .B2(
        n5178), .ZN(n4715) );
  OAI21_X1 U5173 ( .B1(n4896), .B2(n4733), .A(n4715), .ZN(n4716) );
  AOI21_X1 U5174 ( .B1(n4717), .B2(n5305), .A(n4716), .ZN(n4718) );
  OAI21_X1 U5175 ( .B1(n4841), .B2(n4898), .A(n4718), .ZN(U3269) );
  NAND2_X1 U5176 ( .A1(n4719), .A2(n4739), .ZN(n5271) );
  NAND2_X1 U5177 ( .A1(n5271), .A2(n4720), .ZN(n4721) );
  XNOR2_X1 U5178 ( .A(n4721), .B(n4722), .ZN(n5254) );
  INV_X1 U5179 ( .A(n5254), .ZN(n4736) );
  NOR2_X1 U5180 ( .A1(n4737), .A2(n4743), .ZN(n4723) );
  XNOR2_X1 U5181 ( .A(n4723), .B(n4722), .ZN(n4728) );
  NAND2_X1 U5182 ( .A1(n5312), .A2(n5283), .ZN(n4726) );
  NAND2_X1 U5183 ( .A1(n4724), .A2(n5054), .ZN(n4725) );
  NAND2_X1 U5184 ( .A1(n4726), .A2(n4725), .ZN(n5242) );
  AOI21_X1 U5185 ( .B1(n2630), .B2(n5282), .A(n5242), .ZN(n4727) );
  OAI21_X1 U5186 ( .B1(n4728), .B2(n5115), .A(n4727), .ZN(n5252) );
  OAI21_X1 U5187 ( .B1(n4748), .B2(n4729), .A(n5335), .ZN(n4730) );
  OR2_X1 U5188 ( .A1(n4730), .A2(n5277), .ZN(n5251) );
  AOI22_X1 U5189 ( .A1(n5348), .A2(REG2_REG_19__SCAN_IN), .B1(n4731), .B2(
        n5178), .ZN(n4732) );
  OAI21_X1 U5190 ( .B1(n5251), .B2(n4733), .A(n4732), .ZN(n4734) );
  AOI21_X1 U5191 ( .B1(n5252), .B2(n5305), .A(n4734), .ZN(n4735) );
  OAI21_X1 U5192 ( .B1(n4736), .B2(n4841), .A(n4735), .ZN(U3271) );
  XOR2_X1 U5193 ( .A(n4739), .B(n4719), .Z(n5234) );
  INV_X1 U5194 ( .A(n4737), .ZN(n4744) );
  INV_X1 U5195 ( .A(n4738), .ZN(n4740) );
  OAI21_X1 U5196 ( .B1(n4741), .B2(n4740), .A(n4739), .ZN(n4742) );
  OAI211_X1 U5197 ( .C1(n4744), .C2(n4743), .A(n4742), .B(n5289), .ZN(n4746)
         );
  OAI22_X1 U5198 ( .A1(n5287), .A2(n5107), .B1(n4775), .B2(n5286), .ZN(n5220)
         );
  INV_X1 U5199 ( .A(n5220), .ZN(n4745) );
  OAI211_X1 U5200 ( .C1(n5327), .C2(n4747), .A(n4746), .B(n4745), .ZN(n5236)
         );
  NAND2_X1 U5201 ( .A1(n5236), .A2(n5305), .ZN(n4751) );
  AOI21_X1 U5202 ( .B1(n5227), .B2(n2769), .A(n4748), .ZN(n5237) );
  OAI22_X1 U5203 ( .A1(n5305), .A2(n4571), .B1(n5232), .B2(n5300), .ZN(n4749)
         );
  AOI21_X1 U5204 ( .B1(n5237), .B2(n5344), .A(n4749), .ZN(n4750) );
  OAI211_X1 U5205 ( .C1(n5234), .C2(n4841), .A(n4751), .B(n4750), .ZN(U3272)
         );
  XNOR2_X1 U5206 ( .A(n4753), .B(n4752), .ZN(n5216) );
  INV_X1 U5207 ( .A(n5216), .ZN(n4769) );
  NOR2_X1 U5208 ( .A1(n4773), .A2(n4754), .ZN(n4755) );
  XNOR2_X1 U5209 ( .A(n4755), .B(n3633), .ZN(n4760) );
  INV_X1 U5210 ( .A(n4756), .ZN(n4793) );
  OAI22_X1 U5211 ( .A1(n4793), .A2(n5286), .B1(n4757), .B2(n5107), .ZN(n4758)
         );
  AOI21_X1 U5212 ( .B1(n4761), .B2(n5282), .A(n4758), .ZN(n4759) );
  OAI21_X1 U5213 ( .B1(n4760), .B2(n5115), .A(n4759), .ZN(n5214) );
  NAND2_X1 U5214 ( .A1(n5214), .A2(n5305), .ZN(n4768) );
  AOI21_X1 U5215 ( .B1(n4781), .B2(n4761), .A(n5291), .ZN(n4762) );
  AND2_X1 U5216 ( .A1(n4762), .A2(n2769), .ZN(n5215) );
  INV_X1 U5217 ( .A(n4763), .ZN(n4764) );
  OAI22_X1 U5218 ( .A1(n5305), .A2(n4765), .B1(n4764), .B2(n5300), .ZN(n4766)
         );
  AOI21_X1 U5219 ( .B1(n5215), .B2(n4838), .A(n4766), .ZN(n4767) );
  OAI211_X1 U5220 ( .C1(n4769), .C2(n4841), .A(n4768), .B(n4767), .ZN(U3273)
         );
  OAI21_X1 U5221 ( .B1(n4771), .B2(n4770), .A(n5289), .ZN(n4772) );
  OR2_X1 U5222 ( .A1(n4773), .A2(n4772), .ZN(n4778) );
  OAI22_X1 U5223 ( .A1(n4775), .A2(n5107), .B1(n4774), .B2(n5286), .ZN(n4776)
         );
  INV_X1 U5224 ( .A(n4776), .ZN(n4777) );
  OAI211_X1 U5225 ( .C1(n5327), .C2(n4779), .A(n4778), .B(n4777), .ZN(n5208)
         );
  OR2_X1 U5226 ( .A1(n4804), .A2(n4779), .ZN(n4780) );
  NAND2_X1 U5227 ( .A1(n4781), .A2(n4780), .ZN(n5206) );
  OR2_X1 U5228 ( .A1(n4783), .A2(n4782), .ZN(n5204) );
  NAND3_X1 U5229 ( .A1(n5204), .A2(n4784), .A3(n4863), .ZN(n4787) );
  AOI22_X1 U5230 ( .A1(n5348), .A2(REG2_REG_16__SCAN_IN), .B1(n4785), .B2(
        n5178), .ZN(n4786) );
  OAI211_X1 U5231 ( .C1(n5302), .C2(n5206), .A(n4787), .B(n4786), .ZN(n4788)
         );
  AOI21_X1 U5232 ( .B1(n5305), .B2(n5208), .A(n4788), .ZN(n4789) );
  INV_X1 U5233 ( .A(n4789), .ZN(U3274) );
  OAI211_X1 U5234 ( .C1(n4791), .C2(n3664), .A(n5289), .B(n4790), .ZN(n4795)
         );
  OAI22_X1 U5235 ( .A1(n4793), .A2(n5107), .B1(n4792), .B2(n5286), .ZN(n5189)
         );
  INV_X1 U5236 ( .A(n5189), .ZN(n4794) );
  OAI211_X1 U5237 ( .C1(n5327), .C2(n4796), .A(n4795), .B(n4794), .ZN(n5198)
         );
  INV_X1 U5238 ( .A(n5198), .ZN(n4809) );
  INV_X1 U5239 ( .A(n5154), .ZN(n4800) );
  INV_X1 U5240 ( .A(n4797), .ZN(n4798) );
  OAI21_X1 U5241 ( .B1(n4800), .B2(n4799), .A(n4798), .ZN(n4816) );
  NAND2_X1 U5242 ( .A1(n4816), .A2(n4815), .ZN(n4814) );
  NAND2_X1 U5243 ( .A1(n4801), .A2(n4814), .ZN(n4802) );
  XNOR2_X1 U5244 ( .A(n4803), .B(n4802), .ZN(n5200) );
  NAND2_X1 U5245 ( .A1(n5200), .A2(n4863), .ZN(n4808) );
  AOI211_X1 U5246 ( .C1(n5193), .C2(n4817), .A(n5291), .B(n4804), .ZN(n5199)
         );
  INV_X1 U5247 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4805) );
  OAI22_X1 U5248 ( .A1(n5305), .A2(n4805), .B1(n5197), .B2(n5300), .ZN(n4806)
         );
  AOI21_X1 U5249 ( .B1(n5199), .B2(n4838), .A(n4806), .ZN(n4807) );
  OAI211_X1 U5250 ( .C1(n5348), .C2(n4809), .A(n4808), .B(n4807), .ZN(U3275)
         );
  XNOR2_X1 U5251 ( .A(n4431), .B(n4810), .ZN(n4813) );
  NOR2_X1 U5252 ( .A1(n4818), .A2(n5327), .ZN(n4812) );
  AOI211_X1 U5253 ( .C1(n4813), .C2(n5289), .A(n4812), .B(n4811), .ZN(n5182)
         );
  OAI21_X1 U5254 ( .B1(n4816), .B2(n4815), .A(n4814), .ZN(n5185) );
  INV_X1 U5255 ( .A(n5166), .ZN(n4819) );
  OAI21_X1 U5256 ( .B1(n4819), .B2(n4818), .A(n4817), .ZN(n5183) );
  AOI22_X1 U5257 ( .A1(n5348), .A2(REG2_REG_14__SCAN_IN), .B1(n5178), .B2(
        n4820), .ZN(n4821) );
  OAI21_X1 U5258 ( .B1(n5183), .B2(n5302), .A(n4821), .ZN(n4822) );
  AOI21_X1 U5259 ( .B1(n5185), .B2(n4863), .A(n4822), .ZN(n4823) );
  OAI21_X1 U5260 ( .B1(n5348), .B2(n5182), .A(n4823), .ZN(U3276) );
  OAI21_X1 U5261 ( .B1(n4825), .B2(n4826), .A(n4824), .ZN(n5150) );
  INV_X1 U5262 ( .A(n5150), .ZN(n4842) );
  XOR2_X1 U5263 ( .A(n4827), .B(n4826), .Z(n4831) );
  AOI21_X1 U5264 ( .B1(n4829), .B2(n5282), .A(n4828), .ZN(n4830) );
  OAI21_X1 U5265 ( .B1(n4831), .B2(n5115), .A(n4830), .ZN(n5148) );
  NAND2_X1 U5266 ( .A1(n5148), .A2(n5305), .ZN(n4840) );
  OR2_X1 U5267 ( .A1(n4856), .A2(n4832), .ZN(n4833) );
  AND3_X1 U5268 ( .A1(n5164), .A2(n4833), .A3(n5335), .ZN(n5149) );
  INV_X1 U5269 ( .A(n4834), .ZN(n4835) );
  OAI22_X1 U5270 ( .A1(n5305), .A2(n4836), .B1(n4835), .B2(n5300), .ZN(n4837)
         );
  AOI21_X1 U5271 ( .B1(n5149), .B2(n4838), .A(n4837), .ZN(n4839) );
  OAI211_X1 U5272 ( .C1(n4842), .C2(n4841), .A(n4840), .B(n4839), .ZN(U3278)
         );
  OAI211_X1 U5273 ( .C1(n4845), .C2(n4844), .A(n4843), .B(n5289), .ZN(n4852)
         );
  OR2_X1 U5274 ( .A1(n5108), .A2(n5286), .ZN(n4848) );
  NAND2_X1 U5275 ( .A1(n4846), .A2(n5282), .ZN(n4847) );
  OAI211_X1 U5276 ( .C1(n4849), .C2(n5107), .A(n4848), .B(n4847), .ZN(n4850)
         );
  INV_X1 U5277 ( .A(n4850), .ZN(n4851) );
  NAND2_X1 U5278 ( .A1(n4852), .A2(n4851), .ZN(n5142) );
  INV_X1 U5279 ( .A(n5142), .ZN(n4865) );
  OAI21_X1 U5280 ( .B1(n4855), .B2(n4854), .A(n4853), .ZN(n5144) );
  INV_X1 U5281 ( .A(n4856), .ZN(n4857) );
  OAI21_X1 U5282 ( .B1(n4859), .B2(n4858), .A(n4857), .ZN(n5141) );
  AOI22_X1 U5283 ( .A1(n5348), .A2(REG2_REG_11__SCAN_IN), .B1(n4860), .B2(
        n5178), .ZN(n4861) );
  OAI21_X1 U5284 ( .B1(n5141), .B2(n5302), .A(n4861), .ZN(n4862) );
  AOI21_X1 U5285 ( .B1(n5144), .B2(n4863), .A(n4862), .ZN(n4864) );
  OAI21_X1 U5286 ( .B1(n5348), .B2(n4865), .A(n4864), .ZN(U3279) );
  AND2_X1 U5287 ( .A1(n4866), .A2(n5173), .ZN(n5022) );
  INV_X1 U5288 ( .A(n4914), .ZN(n4867) );
  NAND2_X1 U5289 ( .A1(n5022), .A2(n4867), .ZN(n4868) );
  MUX2_X1 U5290 ( .A(REG1_REG_29__SCAN_IN), .B(n4899), .S(n5339), .Z(U3547) );
  OAI211_X1 U5291 ( .C1(n5233), .C2(n4874), .A(n4873), .B(n4872), .ZN(n4900)
         );
  MUX2_X1 U5292 ( .A(REG1_REG_28__SCAN_IN), .B(n4900), .S(n5339), .Z(U3546) );
  AOI21_X1 U5293 ( .B1(n5335), .B2(n4876), .A(n4875), .ZN(n4877) );
  OAI21_X1 U5294 ( .B1(n4878), .B2(n5233), .A(n4877), .ZN(n4901) );
  MUX2_X1 U5295 ( .A(REG1_REG_27__SCAN_IN), .B(n4901), .S(n5339), .Z(U3545) );
  OAI211_X1 U5296 ( .C1(n4881), .C2(n5233), .A(n4880), .B(n4879), .ZN(n4902)
         );
  MUX2_X1 U5297 ( .A(REG1_REG_26__SCAN_IN), .B(n4902), .S(n5339), .Z(U3544) );
  OAI211_X1 U5298 ( .C1(n4884), .C2(n5233), .A(n4883), .B(n4882), .ZN(n4903)
         );
  MUX2_X1 U5299 ( .A(REG1_REG_25__SCAN_IN), .B(n4903), .S(n5339), .Z(U3543) );
  OAI211_X1 U5300 ( .C1(n4887), .C2(n5233), .A(n4886), .B(n4885), .ZN(n4904)
         );
  MUX2_X1 U5301 ( .A(REG1_REG_24__SCAN_IN), .B(n4904), .S(n5339), .Z(U3542) );
  NAND3_X1 U5302 ( .A1(n4888), .A2(n4678), .A3(n5293), .ZN(n4889) );
  OAI211_X1 U5303 ( .C1(n5291), .C2(n4891), .A(n4890), .B(n4889), .ZN(n4905)
         );
  MUX2_X1 U5304 ( .A(REG1_REG_23__SCAN_IN), .B(n4905), .S(n5339), .Z(U3541) );
  AOI21_X1 U5305 ( .B1(n5335), .B2(n4893), .A(n4892), .ZN(n4894) );
  OAI21_X1 U5306 ( .B1(n5233), .B2(n4895), .A(n4894), .ZN(n4906) );
  MUX2_X1 U5307 ( .A(REG1_REG_22__SCAN_IN), .B(n4906), .S(n5339), .Z(U3540) );
  OAI211_X1 U5308 ( .C1(n5233), .C2(n4898), .A(n4897), .B(n4896), .ZN(n4907)
         );
  MUX2_X1 U5309 ( .A(REG1_REG_21__SCAN_IN), .B(n4907), .S(n5339), .Z(U3539) );
  MUX2_X1 U5310 ( .A(REG0_REG_29__SCAN_IN), .B(n4899), .S(n5343), .Z(U3515) );
  MUX2_X1 U5311 ( .A(REG0_REG_28__SCAN_IN), .B(n4900), .S(n5343), .Z(U3514) );
  MUX2_X1 U5312 ( .A(REG0_REG_27__SCAN_IN), .B(n4901), .S(n5343), .Z(U3513) );
  MUX2_X1 U5313 ( .A(REG0_REG_26__SCAN_IN), .B(n4902), .S(n5343), .Z(U3512) );
  MUX2_X1 U5314 ( .A(REG0_REG_25__SCAN_IN), .B(n4903), .S(n5343), .Z(U3511) );
  MUX2_X1 U5315 ( .A(REG0_REG_24__SCAN_IN), .B(n4904), .S(n5343), .Z(U3510) );
  MUX2_X1 U5316 ( .A(REG0_REG_23__SCAN_IN), .B(n4905), .S(n5343), .Z(U3509) );
  MUX2_X1 U5317 ( .A(REG0_REG_22__SCAN_IN), .B(n4906), .S(n5343), .Z(U3508) );
  MUX2_X1 U5318 ( .A(REG0_REG_21__SCAN_IN), .B(n4907), .S(n5343), .Z(U3507) );
  NOR3_X1 U5319 ( .A1(n2863), .A2(IR_REG_30__SCAN_IN), .A3(n2841), .ZN(n4908)
         );
  MUX2_X1 U5320 ( .A(DATAI_31_), .B(n4908), .S(STATE_REG_SCAN_IN), .Z(U3321)
         );
  MUX2_X1 U5321 ( .A(DATAI_30_), .B(n4909), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5322 ( .A(n4910), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5323 ( .A(n4981), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U5324 ( .A(n4911), .B(DATAI_26_), .S(U3149), .Z(U3326) );
  MUX2_X1 U5325 ( .A(n4912), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5326 ( .A(DATAI_24_), .B(n4913), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5327 ( .A(n4914), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5328 ( .A(n4915), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5329 ( .A(DATAI_20_), .B(n4916), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5330 ( .A(DATAI_19_), .B(n5173), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5331 ( .A(n4917), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U5332 ( .A(DATAI_16_), .B(n4918), .S(STATE_REG_SCAN_IN), .Z(U3336)
         );
  MUX2_X1 U5333 ( .A(n4919), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5334 ( .A(n4920), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5335 ( .A(DATAI_13_), .B(n4921), .S(STATE_REG_SCAN_IN), .Z(U3339)
         );
  MUX2_X1 U5336 ( .A(n4922), .B(DATAI_12_), .S(U3149), .Z(U3340) );
  MUX2_X1 U5337 ( .A(n4923), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5338 ( .A(DATAI_9_), .B(n4924), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5339 ( .A(n4925), .B(DATAI_8_), .S(U3149), .Z(U3344) );
  MUX2_X1 U5340 ( .A(n4926), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5341 ( .A(DATAI_6_), .B(n2561), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U5342 ( .A(DATAI_5_), .B(n4928), .S(STATE_REG_SCAN_IN), .Z(U3347) );
  MUX2_X1 U5343 ( .A(n5002), .B(DATAI_4_), .S(U3149), .Z(U3348) );
  MUX2_X1 U5344 ( .A(n4929), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  INV_X1 U5345 ( .A(DATAI_23_), .ZN(n4931) );
  AOI21_X1 U5346 ( .B1(U3149), .B2(n4931), .A(n4930), .ZN(U3329) );
  AND2_X1 U5347 ( .A1(n4954), .A2(D_REG_2__SCAN_IN), .ZN(U3320) );
  AND2_X1 U5348 ( .A1(n4954), .A2(D_REG_3__SCAN_IN), .ZN(U3319) );
  NOR2_X1 U5349 ( .A1(n4956), .A2(n4932), .ZN(U3318) );
  AND2_X1 U5350 ( .A1(n4954), .A2(D_REG_5__SCAN_IN), .ZN(U3317) );
  AND2_X1 U5351 ( .A1(n4954), .A2(D_REG_6__SCAN_IN), .ZN(U3316) );
  INV_X1 U5352 ( .A(D_REG_7__SCAN_IN), .ZN(n4933) );
  NOR2_X1 U5353 ( .A1(n4956), .A2(n4933), .ZN(U3315) );
  NOR2_X1 U5354 ( .A1(n4956), .A2(n4934), .ZN(U3314) );
  INV_X1 U5355 ( .A(D_REG_9__SCAN_IN), .ZN(n4935) );
  NOR2_X1 U5356 ( .A1(n4956), .A2(n4935), .ZN(U3313) );
  NOR2_X1 U5357 ( .A1(n4956), .A2(n4936), .ZN(U3312) );
  AND2_X1 U5358 ( .A1(n4954), .A2(D_REG_11__SCAN_IN), .ZN(U3311) );
  NOR2_X1 U5359 ( .A1(n4956), .A2(n4937), .ZN(U3310) );
  NOR2_X1 U5360 ( .A1(n4956), .A2(n4938), .ZN(U3309) );
  NOR2_X1 U5361 ( .A1(n4956), .A2(n4939), .ZN(U3308) );
  NOR2_X1 U5362 ( .A1(n4956), .A2(n4940), .ZN(U3307) );
  NOR2_X1 U5363 ( .A1(n4956), .A2(n4941), .ZN(U3306) );
  NOR2_X1 U5364 ( .A1(n4956), .A2(n4942), .ZN(U3305) );
  NOR2_X1 U5365 ( .A1(n4956), .A2(n4943), .ZN(U3304) );
  NOR2_X1 U5366 ( .A1(n4956), .A2(n4944), .ZN(U3303) );
  NOR2_X1 U5367 ( .A1(n4956), .A2(n4945), .ZN(U3302) );
  AND2_X1 U5368 ( .A1(n4954), .A2(D_REG_21__SCAN_IN), .ZN(U3301) );
  NOR2_X1 U5369 ( .A1(n4956), .A2(n4946), .ZN(U3300) );
  NOR2_X1 U5370 ( .A1(n4956), .A2(n4947), .ZN(U3299) );
  INV_X1 U5371 ( .A(D_REG_24__SCAN_IN), .ZN(n4948) );
  NOR2_X1 U5372 ( .A1(n4956), .A2(n4948), .ZN(U3298) );
  NOR2_X1 U5373 ( .A1(n4956), .A2(n4949), .ZN(U3297) );
  INV_X1 U5374 ( .A(D_REG_26__SCAN_IN), .ZN(n4950) );
  NOR2_X1 U5375 ( .A1(n4956), .A2(n4950), .ZN(U3296) );
  NOR2_X1 U5376 ( .A1(n4956), .A2(n4951), .ZN(U3295) );
  NOR2_X1 U5377 ( .A1(n4956), .A2(n4952), .ZN(U3294) );
  NOR2_X1 U5378 ( .A1(n4956), .A2(n4953), .ZN(U3293) );
  AND2_X1 U5379 ( .A1(n4954), .A2(D_REG_30__SCAN_IN), .ZN(U3292) );
  NOR2_X1 U5380 ( .A1(n4956), .A2(n4955), .ZN(U3291) );
  INV_X1 U5381 ( .A(REG1_REG_0__SCAN_IN), .ZN(n5019) );
  AND2_X1 U5382 ( .A1(n2870), .A2(n5019), .ZN(n4960) );
  OR2_X1 U5383 ( .A1(n2870), .A2(REG2_REG_0__SCAN_IN), .ZN(n4957) );
  NAND2_X1 U5384 ( .A1(n4957), .A2(n4981), .ZN(n4961) );
  NOR2_X1 U5385 ( .A1(n4961), .A2(n4960), .ZN(n4959) );
  MUX2_X1 U5386 ( .A(n4960), .B(n4959), .S(n4958), .Z(n4963) );
  NAND2_X1 U5387 ( .A1(n4961), .A2(n2566), .ZN(n4983) );
  INV_X1 U5388 ( .A(n4983), .ZN(n4962) );
  OR2_X1 U5389 ( .A1(n4963), .A2(n4962), .ZN(n4965) );
  AOI22_X1 U5390 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4998), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4964) );
  OAI21_X1 U5391 ( .B1(n4966), .B2(n4965), .A(n4964), .ZN(U3240) );
  AOI22_X1 U5392 ( .A1(ADDR_REG_1__SCAN_IN), .A2(n4998), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4977) );
  INV_X1 U5393 ( .A(n4967), .ZN(n4969) );
  AOI211_X1 U5394 ( .C1(n4978), .C2(n4970), .A(n4969), .B(n4968), .ZN(n4971)
         );
  NOR2_X1 U5395 ( .A1(n2566), .A2(n5019), .ZN(n4974) );
  OAI211_X1 U5396 ( .C1(n4974), .C2(n4973), .A(n5010), .B(n4972), .ZN(n4975)
         );
  NAND3_X1 U5397 ( .A1(n4977), .A2(n4976), .A3(n4975), .ZN(U3241) );
  AOI22_X1 U5398 ( .A1(STATE_REG_SCAN_IN), .A2(n2566), .B1(n2721), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5399 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4998), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4997) );
  MUX2_X1 U5400 ( .A(n4980), .B(n2567), .S(n4979), .Z(n4982) );
  NAND2_X1 U5401 ( .A1(n4982), .A2(n4981), .ZN(n4985) );
  AND2_X1 U5402 ( .A1(n4983), .A2(U4043), .ZN(n4984) );
  NAND2_X1 U5403 ( .A1(n4985), .A2(n4984), .ZN(n5007) );
  AOI21_X1 U5404 ( .B1(n4988), .B2(n4987), .A(n4986), .ZN(n4990) );
  AOI22_X1 U5405 ( .A1(n5005), .A2(n4990), .B1(n5003), .B2(n4989), .ZN(n4991)
         );
  AND2_X1 U5406 ( .A1(n5007), .A2(n4991), .ZN(n4996) );
  OAI211_X1 U5407 ( .C1(n4994), .C2(n4993), .A(n5010), .B(n4992), .ZN(n4995)
         );
  NAND3_X1 U5408 ( .A1(n4997), .A2(n4996), .A3(n4995), .ZN(U3242) );
  AOI22_X1 U5409 ( .A1(ADDR_REG_4__SCAN_IN), .A2(n4998), .B1(
        REG3_REG_4__SCAN_IN), .B2(U3149), .ZN(n5013) );
  AOI21_X1 U5410 ( .B1(n5001), .B2(n5000), .A(n4999), .ZN(n5004) );
  AOI22_X1 U5411 ( .A1(n5005), .A2(n5004), .B1(n5003), .B2(n5002), .ZN(n5006)
         );
  AND2_X1 U5412 ( .A1(n5007), .A2(n5006), .ZN(n5012) );
  XOR2_X1 U5413 ( .A(REG1_REG_4__SCAN_IN), .B(n5008), .Z(n5009) );
  NAND2_X1 U5414 ( .A1(n5010), .A2(n5009), .ZN(n5011) );
  NAND3_X1 U5415 ( .A1(n5013), .A2(n5012), .A3(n5011), .ZN(U3244) );
  AND2_X1 U5416 ( .A1(n5015), .A2(n5014), .ZN(n5024) );
  OAI21_X1 U5417 ( .B1(n5177), .B2(n5289), .A(n5016), .ZN(n5017) );
  OAI21_X1 U5418 ( .B1(n5018), .B2(n5107), .A(n5017), .ZN(n5026) );
  NOR2_X1 U5419 ( .A1(n5024), .A2(n5026), .ZN(n5021) );
  AOI22_X1 U5420 ( .A1(n5339), .A2(n5021), .B1(n5019), .B2(n5337), .ZN(U3518)
         );
  INV_X1 U5421 ( .A(REG0_REG_0__SCAN_IN), .ZN(n5020) );
  AOI22_X1 U5422 ( .A1(n5343), .A2(n5021), .B1(n5020), .B2(n5340), .ZN(U3467)
         );
  INV_X1 U5423 ( .A(REG2_REG_0__SCAN_IN), .ZN(n5029) );
  INV_X1 U5424 ( .A(n5022), .ZN(n5023) );
  AOI22_X1 U5425 ( .A1(n5024), .A2(n5023), .B1(REG3_REG_0__SCAN_IN), .B2(n5178), .ZN(n5025) );
  INV_X1 U5426 ( .A(n5025), .ZN(n5027) );
  NOR2_X1 U5427 ( .A1(n5027), .A2(n5026), .ZN(n5028) );
  AOI22_X1 U5428 ( .A1(n5348), .A2(n5029), .B1(n5028), .B2(n5305), .ZN(U3290)
         );
  AOI22_X1 U5429 ( .A1(STATE_REG_SCAN_IN), .A2(n5031), .B1(n5030), .B2(U3149), 
        .ZN(U3351) );
  NOR3_X1 U5430 ( .A1(n5032), .A2(n2518), .A3(n5291), .ZN(n5034) );
  NOR2_X1 U5431 ( .A1(n5034), .A2(n5033), .ZN(n5037) );
  AOI22_X1 U5432 ( .A1(n5339), .A2(n5037), .B1(n5035), .B2(n5337), .ZN(U3519)
         );
  INV_X1 U5433 ( .A(REG0_REG_1__SCAN_IN), .ZN(n5036) );
  AOI22_X1 U5434 ( .A1(n5343), .A2(n5037), .B1(n5036), .B2(n5340), .ZN(U3469)
         );
  AOI22_X1 U5435 ( .A1(STATE_REG_SCAN_IN), .A2(n5039), .B1(n5038), .B2(U3149), 
        .ZN(U3350) );
  NOR2_X1 U5436 ( .A1(n5291), .A2(n5040), .ZN(n5041) );
  NOR2_X1 U5437 ( .A1(n5042), .A2(n5041), .ZN(n5045) );
  AOI22_X1 U5438 ( .A1(n5339), .A2(n5045), .B1(n5043), .B2(n5337), .ZN(U3520)
         );
  INV_X1 U5439 ( .A(REG0_REG_2__SCAN_IN), .ZN(n5044) );
  AOI22_X1 U5440 ( .A1(n5343), .A2(n5045), .B1(n5044), .B2(n5340), .ZN(U3471)
         );
  AOI21_X1 U5441 ( .B1(n5048), .B2(n5047), .A(n5046), .ZN(n5067) );
  NAND2_X1 U5442 ( .A1(n5049), .A2(n5050), .ZN(n5051) );
  XNOR2_X1 U5443 ( .A(n5051), .B(n5058), .ZN(n5052) );
  NAND2_X1 U5444 ( .A1(n5052), .A2(n5289), .ZN(n5056) );
  AOI22_X1 U5445 ( .A1(n3471), .A2(n5054), .B1(n5283), .B2(n5053), .ZN(n5055)
         );
  OAI211_X1 U5446 ( .C1(n5327), .C2(n5057), .A(n5056), .B(n5055), .ZN(n5064)
         );
  XNOR2_X1 U5447 ( .A(n5059), .B(n5058), .ZN(n5063) );
  NOR2_X1 U5448 ( .A1(n5063), .A2(n5233), .ZN(n5060) );
  AOI211_X1 U5449 ( .C1(n5335), .C2(n5067), .A(n5064), .B(n5060), .ZN(n5062)
         );
  AOI22_X1 U5450 ( .A1(n5339), .A2(n5062), .B1(n2691), .B2(n5337), .ZN(U3521)
         );
  INV_X1 U5451 ( .A(REG0_REG_3__SCAN_IN), .ZN(n5061) );
  AOI22_X1 U5452 ( .A1(n5343), .A2(n5062), .B1(n5061), .B2(n5340), .ZN(U3473)
         );
  INV_X1 U5453 ( .A(n5063), .ZN(n5065) );
  AOI21_X1 U5454 ( .B1(n5177), .B2(n5065), .A(n5064), .ZN(n5070) );
  AOI22_X1 U5455 ( .A1(n5067), .A2(n5344), .B1(n5178), .B2(n5066), .ZN(n5068)
         );
  OAI221_X1 U5456 ( .B1(n5348), .B2(n5070), .C1(n5305), .C2(n5069), .A(n5068), 
        .ZN(U3287) );
  OAI211_X1 U5457 ( .C1(n5233), .C2(n5073), .A(n5072), .B(n5071), .ZN(n5074)
         );
  INV_X1 U5458 ( .A(n5074), .ZN(n5076) );
  AOI22_X1 U5459 ( .A1(n5339), .A2(n5076), .B1(n2594), .B2(n5337), .ZN(U3522)
         );
  INV_X1 U5460 ( .A(REG0_REG_4__SCAN_IN), .ZN(n5075) );
  AOI22_X1 U5461 ( .A1(n5343), .A2(n5076), .B1(n5075), .B2(n5340), .ZN(U3475)
         );
  AOI211_X1 U5462 ( .C1(n5079), .C2(n5293), .A(n5078), .B(n5077), .ZN(n5082)
         );
  AOI22_X1 U5463 ( .A1(n5339), .A2(n5082), .B1(n5080), .B2(n5337), .ZN(U3523)
         );
  INV_X1 U5464 ( .A(REG0_REG_5__SCAN_IN), .ZN(n5081) );
  AOI22_X1 U5465 ( .A1(n5343), .A2(n5082), .B1(n5081), .B2(n5340), .ZN(U3477)
         );
  NAND2_X1 U5466 ( .A1(n5083), .A2(n5293), .ZN(n5086) );
  NAND2_X1 U5467 ( .A1(n5084), .A2(n5335), .ZN(n5085) );
  AOI22_X1 U5468 ( .A1(n5339), .A2(n5089), .B1(n3323), .B2(n5337), .ZN(U3524)
         );
  INV_X1 U5469 ( .A(REG0_REG_6__SCAN_IN), .ZN(n5088) );
  AOI22_X1 U5470 ( .A1(n5343), .A2(n5089), .B1(n5088), .B2(n5340), .ZN(U3479)
         );
  AOI211_X1 U5471 ( .C1(n5092), .C2(n5293), .A(n5091), .B(n5090), .ZN(n5094)
         );
  AOI22_X1 U5472 ( .A1(n5339), .A2(n5094), .B1(n3321), .B2(n5337), .ZN(U3525)
         );
  INV_X1 U5473 ( .A(REG0_REG_7__SCAN_IN), .ZN(n5093) );
  AOI22_X1 U5474 ( .A1(n5343), .A2(n5094), .B1(n5093), .B2(n5340), .ZN(U3481)
         );
  OAI21_X1 U5475 ( .B1(n5291), .B2(n5096), .A(n5095), .ZN(n5097) );
  AOI21_X1 U5476 ( .B1(n5098), .B2(n5293), .A(n5097), .ZN(n5101) );
  INV_X1 U5477 ( .A(REG1_REG_8__SCAN_IN), .ZN(n5099) );
  AOI22_X1 U5478 ( .A1(n5339), .A2(n5101), .B1(n5099), .B2(n5337), .ZN(U3526)
         );
  INV_X1 U5479 ( .A(REG0_REG_8__SCAN_IN), .ZN(n5100) );
  AOI22_X1 U5480 ( .A1(n5343), .A2(n5101), .B1(n5100), .B2(n5340), .ZN(U3483)
         );
  XNOR2_X1 U5481 ( .A(n5102), .B(n5113), .ZN(n5126) );
  INV_X1 U5482 ( .A(n5103), .ZN(n5106) );
  OAI21_X1 U5483 ( .B1(n5106), .B2(n5105), .A(n5104), .ZN(n5124) );
  OAI22_X1 U5484 ( .A1(n5109), .A2(n5286), .B1(n5108), .B2(n5107), .ZN(n5118)
         );
  NOR2_X1 U5485 ( .A1(n5111), .A2(n5110), .ZN(n5114) );
  MUX2_X1 U5486 ( .A(n5114), .B(n5113), .S(n5112), .Z(n5116) );
  NOR2_X1 U5487 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  AOI211_X1 U5488 ( .C1(n5282), .C2(n5119), .A(n5118), .B(n5117), .ZN(n5127)
         );
  OAI21_X1 U5489 ( .B1(n5291), .B2(n5124), .A(n5127), .ZN(n5120) );
  AOI21_X1 U5490 ( .B1(n5126), .B2(n5293), .A(n5120), .ZN(n5123) );
  AOI22_X1 U5491 ( .A1(n5339), .A2(n5123), .B1(n5121), .B2(n5337), .ZN(U3527)
         );
  INV_X1 U5492 ( .A(REG0_REG_9__SCAN_IN), .ZN(n5122) );
  AOI22_X1 U5493 ( .A1(n5343), .A2(n5123), .B1(n5122), .B2(n5340), .ZN(U3485)
         );
  INV_X1 U5494 ( .A(n5124), .ZN(n5125) );
  AOI22_X1 U5495 ( .A1(n5125), .A2(n5344), .B1(REG2_REG_9__SCAN_IN), .B2(n5348), .ZN(n5131) );
  INV_X1 U5496 ( .A(n5126), .ZN(n5128) );
  OAI21_X1 U5497 ( .B1(n4869), .B2(n5128), .A(n5127), .ZN(n5129) );
  NAND2_X1 U5498 ( .A1(n5129), .A2(n5305), .ZN(n5130) );
  OAI211_X1 U5499 ( .C1(n5300), .C2(n5132), .A(n5131), .B(n5130), .ZN(U3281)
         );
  NOR2_X1 U5500 ( .A1(n5133), .A2(n5233), .ZN(n5134) );
  AOI211_X1 U5501 ( .C1(n5335), .C2(n5136), .A(n5135), .B(n5134), .ZN(n5138)
         );
  AOI22_X1 U5502 ( .A1(n5339), .A2(n5138), .B1(n3458), .B2(n5337), .ZN(U3528)
         );
  INV_X1 U5503 ( .A(REG0_REG_10__SCAN_IN), .ZN(n5137) );
  AOI22_X1 U5504 ( .A1(n5343), .A2(n5138), .B1(n5137), .B2(n5340), .ZN(U3487)
         );
  OAI22_X1 U5505 ( .A1(U3149), .A2(n5139), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n5140) );
  INV_X1 U5506 ( .A(n5140), .ZN(U3341) );
  NOR2_X1 U5507 ( .A1(n5141), .A2(n5291), .ZN(n5143) );
  AOI211_X1 U5508 ( .C1(n5144), .C2(n5293), .A(n5143), .B(n5142), .ZN(n5147)
         );
  AOI22_X1 U5509 ( .A1(n5339), .A2(n5147), .B1(n5145), .B2(n5337), .ZN(U3529)
         );
  INV_X1 U5510 ( .A(REG0_REG_11__SCAN_IN), .ZN(n5146) );
  AOI22_X1 U5511 ( .A1(n5343), .A2(n5147), .B1(n5146), .B2(n5340), .ZN(U3489)
         );
  AOI211_X1 U5512 ( .C1(n5293), .C2(n5150), .A(n5149), .B(n5148), .ZN(n5153)
         );
  INV_X1 U5513 ( .A(REG1_REG_12__SCAN_IN), .ZN(n5151) );
  AOI22_X1 U5514 ( .A1(n5339), .A2(n5153), .B1(n5151), .B2(n5337), .ZN(U3530)
         );
  INV_X1 U5515 ( .A(REG0_REG_12__SCAN_IN), .ZN(n5152) );
  AOI22_X1 U5516 ( .A1(n5343), .A2(n5153), .B1(n5152), .B2(n5340), .ZN(U3491)
         );
  XNOR2_X1 U5517 ( .A(n5154), .B(n2765), .ZN(n5176) );
  NAND2_X1 U5518 ( .A1(n5156), .A2(n5155), .ZN(n5157) );
  XNOR2_X1 U5519 ( .A(n5157), .B(n2765), .ZN(n5162) );
  INV_X1 U5520 ( .A(n5158), .ZN(n5159) );
  OAI21_X1 U5521 ( .B1(n5160), .B2(n5327), .A(n5159), .ZN(n5161) );
  AOI21_X1 U5522 ( .B1(n5162), .B2(n5289), .A(n5161), .ZN(n5174) );
  NAND2_X1 U5523 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  NAND3_X1 U5524 ( .A1(n5166), .A2(n5335), .A3(n5165), .ZN(n5167) );
  INV_X1 U5525 ( .A(n5172), .ZN(n5168) );
  AOI21_X1 U5526 ( .B1(n5176), .B2(n5293), .A(n5168), .ZN(n5171) );
  AOI22_X1 U5527 ( .A1(n5339), .A2(n5171), .B1(n5169), .B2(n5337), .ZN(U3531)
         );
  INV_X1 U5528 ( .A(REG0_REG_13__SCAN_IN), .ZN(n5170) );
  AOI22_X1 U5529 ( .A1(n5343), .A2(n5171), .B1(n5170), .B2(n5340), .ZN(U3493)
         );
  AOI21_X1 U5530 ( .B1(n5174), .B2(n5173), .A(n5172), .ZN(n5175) );
  AOI21_X1 U5531 ( .B1(n5177), .B2(n5176), .A(n5175), .ZN(n5181) );
  NAND2_X1 U5532 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  OAI221_X1 U5533 ( .B1(n5348), .B2(n5181), .C1(n5305), .C2(n4498), .A(n5180), 
        .ZN(U3277) );
  OAI21_X1 U5534 ( .B1(n5291), .B2(n5183), .A(n5182), .ZN(n5184) );
  AOI21_X1 U5535 ( .B1(n5293), .B2(n5185), .A(n5184), .ZN(n5188) );
  INV_X1 U5536 ( .A(REG1_REG_14__SCAN_IN), .ZN(n5186) );
  AOI22_X1 U5537 ( .A1(n5339), .A2(n5188), .B1(n5186), .B2(n5337), .ZN(U3532)
         );
  INV_X1 U5538 ( .A(REG0_REG_14__SCAN_IN), .ZN(n5187) );
  AOI22_X1 U5539 ( .A1(n5343), .A2(n5188), .B1(n5187), .B2(n5340), .ZN(U3495)
         );
  AOI22_X1 U5540 ( .A1(n5243), .A2(n5189), .B1(REG3_REG_15__SCAN_IN), .B2(
        U3149), .ZN(n5196) );
  XNOR2_X1 U5541 ( .A(n5191), .B(n5190), .ZN(n5192) );
  XNOR2_X1 U5542 ( .A(n3833), .B(n5192), .ZN(n5194) );
  AOI22_X1 U5543 ( .A1(n5194), .A2(n5322), .B1(n5193), .B2(n5246), .ZN(n5195)
         );
  OAI211_X1 U5544 ( .C1(n5326), .C2(n5197), .A(n5196), .B(n5195), .ZN(U3238)
         );
  AOI211_X1 U5545 ( .C1(n5200), .C2(n5293), .A(n5199), .B(n5198), .ZN(n5203)
         );
  AOI22_X1 U5546 ( .A1(n5339), .A2(n5203), .B1(n5201), .B2(n5337), .ZN(U3533)
         );
  INV_X1 U5547 ( .A(REG0_REG_15__SCAN_IN), .ZN(n5202) );
  AOI22_X1 U5548 ( .A1(n5343), .A2(n5203), .B1(n5202), .B2(n5340), .ZN(U3497)
         );
  NAND3_X1 U5549 ( .A1(n5204), .A2(n4784), .A3(n5293), .ZN(n5205) );
  OAI21_X1 U5550 ( .B1(n5206), .B2(n5291), .A(n5205), .ZN(n5207) );
  NOR2_X1 U5551 ( .A1(n5208), .A2(n5207), .ZN(n5211) );
  INV_X1 U5552 ( .A(REG1_REG_16__SCAN_IN), .ZN(n5209) );
  AOI22_X1 U5553 ( .A1(n5339), .A2(n5211), .B1(n5209), .B2(n5337), .ZN(U3534)
         );
  INV_X1 U5554 ( .A(REG0_REG_16__SCAN_IN), .ZN(n5210) );
  AOI22_X1 U5555 ( .A1(n5343), .A2(n5211), .B1(n5210), .B2(n5340), .ZN(U3499)
         );
  INV_X1 U5556 ( .A(DATAI_17_), .ZN(n5212) );
  AOI22_X1 U5557 ( .A1(STATE_REG_SCAN_IN), .A2(n5213), .B1(n5212), .B2(U3149), 
        .ZN(U3335) );
  AOI211_X1 U5558 ( .C1(n5216), .C2(n5293), .A(n5215), .B(n5214), .ZN(n5219)
         );
  AOI22_X1 U5559 ( .A1(n5339), .A2(n5219), .B1(n5217), .B2(n5337), .ZN(U3535)
         );
  INV_X1 U5560 ( .A(REG0_REG_17__SCAN_IN), .ZN(n5218) );
  AOI22_X1 U5561 ( .A1(n5343), .A2(n5219), .B1(n5218), .B2(n5340), .ZN(U3501)
         );
  AOI22_X1 U5562 ( .A1(n5243), .A2(n5220), .B1(REG3_REG_18__SCAN_IN), .B2(
        U3149), .ZN(n5231) );
  AND2_X1 U5563 ( .A1(n5221), .A2(n5225), .ZN(n5224) );
  OAI21_X1 U5564 ( .B1(n5224), .B2(n5222), .A(n5223), .ZN(n5229) );
  AOI21_X1 U5565 ( .B1(n5222), .B2(n2738), .A(n5226), .ZN(n5228) );
  AOI22_X1 U5566 ( .A1(n5229), .A2(n5228), .B1(n5227), .B2(n5246), .ZN(n5230)
         );
  OAI211_X1 U5567 ( .C1(n5326), .C2(n5232), .A(n5231), .B(n5230), .ZN(U3235)
         );
  NOR2_X1 U5568 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  AOI211_X1 U5569 ( .C1(n5335), .C2(n5237), .A(n5236), .B(n5235), .ZN(n5240)
         );
  INV_X1 U5570 ( .A(REG1_REG_18__SCAN_IN), .ZN(n5238) );
  AOI22_X1 U5571 ( .A1(n5339), .A2(n5240), .B1(n5238), .B2(n5337), .ZN(U3536)
         );
  INV_X1 U5572 ( .A(REG0_REG_18__SCAN_IN), .ZN(n5239) );
  AOI22_X1 U5573 ( .A1(n5343), .A2(n5240), .B1(n5239), .B2(n5340), .ZN(U3503)
         );
  AOI22_X1 U5574 ( .A1(n5243), .A2(n5242), .B1(REG3_REG_19__SCAN_IN), .B2(
        U3149), .ZN(n5249) );
  XNOR2_X1 U5575 ( .A(n5244), .B(n5245), .ZN(n5247) );
  AOI22_X1 U5576 ( .A1(n5247), .A2(n5322), .B1(n2630), .B2(n5246), .ZN(n5248)
         );
  OAI211_X1 U5577 ( .C1(n5326), .C2(n5250), .A(n5249), .B(n5248), .ZN(U3216)
         );
  INV_X1 U5578 ( .A(n5251), .ZN(n5253) );
  AOI211_X1 U5579 ( .C1(n5293), .C2(n5254), .A(n5253), .B(n5252), .ZN(n5257)
         );
  AOI22_X1 U5580 ( .A1(n5339), .A2(n5257), .B1(n5255), .B2(n5337), .ZN(U3537)
         );
  INV_X1 U5581 ( .A(REG0_REG_19__SCAN_IN), .ZN(n5256) );
  AOI22_X1 U5582 ( .A1(n5343), .A2(n5257), .B1(n5256), .B2(n5340), .ZN(U3505)
         );
  AOI22_X1 U5583 ( .A1(n5258), .A2(n5284), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n5269) );
  INV_X1 U5584 ( .A(n5260), .ZN(n5262) );
  NOR2_X1 U5585 ( .A1(n5262), .A2(n5261), .ZN(n5263) );
  XNOR2_X1 U5586 ( .A(n5259), .B(n5263), .ZN(n5266) );
  AOI222_X1 U5587 ( .A1(n5267), .A2(n5281), .B1(n5322), .B2(n5266), .C1(n5265), 
        .C2(n5264), .ZN(n5268) );
  OAI211_X1 U5588 ( .C1(n5326), .C2(n5301), .A(n5269), .B(n5268), .ZN(U3230)
         );
  NAND2_X1 U5589 ( .A1(n5271), .A2(n5270), .ZN(n5273) );
  AND2_X1 U5590 ( .A1(n5273), .A2(n5272), .ZN(n5274) );
  XOR2_X1 U5591 ( .A(n5280), .B(n5274), .Z(n5297) );
  OAI21_X1 U5592 ( .B1(n5277), .B2(n5276), .A(n5275), .ZN(n5303) );
  OAI21_X1 U5593 ( .B1(n5280), .B2(n5279), .A(n5278), .ZN(n5290) );
  AOI22_X1 U5594 ( .A1(n5284), .A2(n5283), .B1(n5282), .B2(n5281), .ZN(n5285)
         );
  OAI21_X1 U5595 ( .B1(n5287), .B2(n5286), .A(n5285), .ZN(n5288) );
  AOI21_X1 U5596 ( .B1(n5290), .B2(n5289), .A(n5288), .ZN(n5298) );
  OAI21_X1 U5597 ( .B1(n5291), .B2(n5303), .A(n5298), .ZN(n5292) );
  AOI21_X1 U5598 ( .B1(n5293), .B2(n5297), .A(n5292), .ZN(n5296) );
  INV_X1 U5599 ( .A(REG1_REG_20__SCAN_IN), .ZN(n5294) );
  AOI22_X1 U5600 ( .A1(n5339), .A2(n5296), .B1(n5294), .B2(n5337), .ZN(U3538)
         );
  INV_X1 U5601 ( .A(REG0_REG_20__SCAN_IN), .ZN(n5295) );
  AOI22_X1 U5602 ( .A1(n5343), .A2(n5296), .B1(n5295), .B2(n5340), .ZN(U3506)
         );
  INV_X1 U5603 ( .A(n5297), .ZN(n5299) );
  OAI21_X1 U5604 ( .B1(n5299), .B2(n4869), .A(n5298), .ZN(n5306) );
  OAI22_X1 U5605 ( .A1(n5303), .A2(n5302), .B1(n5301), .B2(n5300), .ZN(n5304)
         );
  AOI221_X1 U5606 ( .B1(REG2_REG_20__SCAN_IN), .B2(n5348), .C1(n5306), .C2(
        n5305), .A(n5304), .ZN(n5307) );
  INV_X1 U5607 ( .A(n5307), .ZN(U3270) );
  NAND2_X1 U5608 ( .A1(n5310), .A2(n5309), .ZN(n5311) );
  XNOR2_X1 U5609 ( .A(n5308), .B(n5311), .ZN(n5323) );
  INV_X1 U5610 ( .A(n5312), .ZN(n5314) );
  OAI22_X1 U5611 ( .A1(n5315), .A2(n5314), .B1(STATE_REG_SCAN_IN), .B2(n5313), 
        .ZN(n5321) );
  OAI22_X1 U5612 ( .A1(n5319), .A2(n5318), .B1(n5317), .B2(n5316), .ZN(n5320)
         );
  AOI211_X1 U5613 ( .C1(n5323), .C2(n5322), .A(n5321), .B(n5320), .ZN(n5324)
         );
  OAI21_X1 U5614 ( .B1(n5326), .B2(n5325), .A(n5324), .ZN(U3220) );
  NOR2_X1 U5615 ( .A1(n5330), .A2(n5327), .ZN(n5328) );
  NOR2_X1 U5616 ( .A1(n5329), .A2(n5328), .ZN(n5333) );
  XNOR2_X1 U5617 ( .A(n5331), .B(n5330), .ZN(n5336) );
  AOI22_X1 U5618 ( .A1(n5336), .A2(n5344), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5348), .ZN(n5332) );
  OAI21_X1 U5619 ( .B1(n5348), .B2(n5333), .A(n5332), .ZN(U3261) );
  INV_X1 U5620 ( .A(n5333), .ZN(n5334) );
  AOI21_X1 U5621 ( .B1(n5336), .B2(n5335), .A(n5334), .ZN(n5342) );
  INV_X1 U5622 ( .A(REG1_REG_30__SCAN_IN), .ZN(n5338) );
  AOI22_X1 U5623 ( .A1(n5339), .A2(n5342), .B1(n5338), .B2(n5337), .ZN(U3548)
         );
  INV_X1 U5624 ( .A(REG0_REG_30__SCAN_IN), .ZN(n5341) );
  AOI22_X1 U5625 ( .A1(n5343), .A2(n5342), .B1(n5341), .B2(n5340), .ZN(U3516)
         );
  AOI22_X1 U5626 ( .A1(n5345), .A2(n5344), .B1(n5348), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n5346) );
  OAI21_X1 U5627 ( .B1(n5348), .B2(n5347), .A(n5346), .ZN(U3260) );
  INV_X2 U2553 ( .A(n2951), .ZN(n3253) );
endmodule

