

module b20_C_SARLock_k_64_10 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226,
         n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
         n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
         n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
         n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296,
         n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306,
         n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316,
         n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326,
         n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336,
         n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346,
         n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356,
         n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366,
         n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396,
         n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406,
         n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416,
         n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426,
         n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436,
         n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446,
         n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
         n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466,
         n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476,
         n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486,
         n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536,
         n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546,
         n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556,
         n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566,
         n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576,
         n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586,
         n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606,
         n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616,
         n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626,
         n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636,
         n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656,
         n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666,
         n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
         n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686,
         n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696,
         n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706,
         n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716,
         n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726,
         n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736,
         n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746,
         n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756,
         n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766,
         n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776,
         n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786,
         n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796,
         n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806,
         n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816,
         n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826,
         n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
         n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846,
         n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856,
         n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866,
         n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876,
         n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886,
         n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896,
         n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906,
         n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916,
         n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
         n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936,
         n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946,
         n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966,
         n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976,
         n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986,
         n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996,
         n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178;

  CLKBUF_X2 U4784 ( .A(n6095), .Z(n4278) );
  CLKBUF_X2 U4785 ( .A(n6095), .Z(n4279) );
  INV_X4 U4786 ( .A(n5642), .ZN(n4429) );
  AOI21_X1 U4787 ( .B1(n9808), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9803), .ZN(
        n9266) );
  NAND2_X1 U4788 ( .A1(n5007), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5425) );
  OR2_X1 U4789 ( .A1(n6285), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6296) );
  OAI21_X1 U4790 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9264), .A(n9263), .ZN(
        n9793) );
  INV_X1 U4791 ( .A(n4388), .ZN(n6530) );
  NAND2_X1 U4792 ( .A1(n8250), .A2(n7957), .ZN(n8296) );
  AND2_X1 U4793 ( .A1(n6400), .A2(n6399), .ZN(n8464) );
  NAND3_X1 U4794 ( .A1(n5685), .A2(n5689), .A3(n5671), .ZN(n6529) );
  INV_X1 U4795 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4975) );
  INV_X2 U4796 ( .A(n8420), .ZN(n8391) );
  BUF_X1 U4797 ( .A(n5001), .Z(n4281) );
  XNOR2_X1 U4798 ( .A(n4976), .B(n4975), .ZN(n9410) );
  NAND2_X1 U4799 ( .A1(n9659), .A2(n4281), .ZN(n6095) );
  AND2_X1 U4800 ( .A1(n6326), .A2(n6325), .ZN(n4277) );
  NAND4_X2 U4801 ( .A1(n6137), .A2(n6136), .A3(n6135), .A4(n6134), .ZN(n8344)
         );
  NOR2_X2 U4802 ( .A1(n6296), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6306) );
  OAI21_X2 U4803 ( .B1(n7497), .B2(n7496), .A(n7495), .ZN(n7586) );
  NOR2_X2 U4804 ( .A1(n6964), .A2(n6963), .ZN(n6962) );
  XNOR2_X2 U4805 ( .A(n4476), .B(n6007), .ZN(n6908) );
  AOI21_X2 U4806 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9669), .A(n9664), .ZN(
        n9771) );
  NAND2_X1 U4807 ( .A1(n5016), .A2(n5014), .ZN(n4280) );
  AOI21_X2 U4808 ( .B1(n6609), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9245), .ZN(
        n9744) );
  AND2_X1 U4809 ( .A1(n8874), .A2(n5649), .ZN(n5731) );
  INV_X1 U4810 ( .A(n9111), .ZN(n9104) );
  INV_X1 U4811 ( .A(n8345), .ZN(n7109) );
  NAND2_X1 U4812 ( .A1(n8773), .A2(n6112), .ZN(n7724) );
  XNOR2_X1 U4813 ( .A(n4998), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5001) );
  NAND2_X2 U4814 ( .A1(n5995), .A2(n5703), .ZN(n6567) );
  CLKBUF_X1 U4815 ( .A(n5823), .Z(n5830) );
  CLKBUF_X3 U4816 ( .A(n6537), .Z(n4388) );
  INV_X4 U4817 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AND2_X1 U4818 ( .A1(n4437), .A2(n4432), .ZN(n9187) );
  NAND2_X1 U4819 ( .A1(n4526), .A2(n4525), .ZN(n8874) );
  AOI21_X1 U4820 ( .B1(n8772), .B2(n5986), .A(n5980), .ZN(n9606) );
  AND2_X1 U4821 ( .A1(n9091), .A2(n9095), .ZN(n9342) );
  NAND2_X1 U4822 ( .A1(n5652), .A2(n5651), .ZN(n9354) );
  NAND2_X1 U4823 ( .A1(n5631), .A2(n5630), .ZN(n9543) );
  XNOR2_X1 U4824 ( .A(n5355), .B(n5356), .ZN(n8885) );
  XNOR2_X1 U4825 ( .A(n5650), .B(n5963), .ZN(n7600) );
  AND2_X1 U4826 ( .A1(n9283), .A2(n9282), .ZN(n9284) );
  AND2_X1 U4827 ( .A1(n5663), .A2(n5662), .ZN(n6058) );
  NOR2_X1 U4828 ( .A1(n7828), .A2(n5890), .ZN(n7811) );
  NAND2_X1 U4829 ( .A1(n4532), .A2(n4531), .ZN(n4530) );
  AOI22_X1 U4830 ( .A1(n7228), .A2(n7227), .B1(n5177), .B2(n5176), .ZN(n7552)
         );
  INV_X2 U4831 ( .A(n9716), .ZN(n9719) );
  AOI21_X1 U4832 ( .B1(n5090), .B2(n5089), .A(n6770), .ZN(n6952) );
  NAND2_X1 U4833 ( .A1(n6295), .A2(n6294), .ZN(n7589) );
  NAND2_X1 U4834 ( .A1(n6816), .A2(n6815), .ZN(n6997) );
  NAND2_X1 U4835 ( .A1(n5234), .A2(n5233), .ZN(n9841) );
  AOI21_X1 U4836 ( .B1(n6840), .B2(n6839), .A(n6812), .ZN(n6816) );
  NAND2_X1 U4837 ( .A1(n5294), .A2(n5293), .ZN(n9005) );
  OAI21_X1 U4838 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6870), .A(n6863), .ZN(
        n9666) );
  OAI21_X1 U4839 ( .B1(n6846), .B2(n6845), .A(n6810), .ZN(n6840) );
  NAND2_X1 U4840 ( .A1(n5248), .A2(n5247), .ZN(n7574) );
  AND2_X1 U4841 ( .A1(n5879), .A2(n4574), .ZN(n7905) );
  OR2_X1 U4842 ( .A1(n5878), .A2(n6554), .ZN(n4573) );
  NAND2_X1 U4843 ( .A1(n5187), .A2(n5186), .ZN(n5189) );
  OR2_X1 U4844 ( .A1(n6729), .A2(n5877), .ZN(n5878) );
  AND2_X1 U4845 ( .A1(n6352), .A2(n8287), .ZN(n6361) );
  AND4_X1 U4846 ( .A1(n5024), .A2(n5023), .A3(n5022), .A4(n5021), .ZN(n7209)
         );
  NAND3_X4 U4847 ( .A1(n6529), .A2(n9180), .A3(n9179), .ZN(n5014) );
  AND3_X1 U4848 ( .A1(n5101), .A2(n5100), .A3(n5099), .ZN(n9921) );
  NAND4_X1 U4849 ( .A1(n5075), .A2(n5074), .A3(n5073), .A4(n5072), .ZN(n9212)
         );
  BUF_X2 U4850 ( .A(n6308), .Z(n6299) );
  NAND2_X1 U4851 ( .A1(n6155), .A2(n6530), .ZN(n8001) );
  AND3_X2 U4852 ( .A1(n5067), .A2(n5066), .A3(n5065), .ZN(n4476) );
  CLKBUF_X2 U4853 ( .A(n5093), .Z(n5704) );
  NAND2_X1 U4854 ( .A1(n4997), .A2(n9652), .ZN(n9659) );
  OAI21_X1 U4855 ( .B1(n4998), .B2(n4993), .A(n4992), .ZN(n4997) );
  AND2_X1 U4856 ( .A1(n4972), .A2(n4967), .ZN(n5671) );
  MUX2_X1 U4857 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6111), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n6112) );
  XNOR2_X1 U4858 ( .A(n5778), .B(n5777), .ZN(n8223) );
  XNOR2_X1 U4859 ( .A(n4968), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U4860 ( .A1(n4990), .A2(n4989), .ZN(n4998) );
  INV_X2 U4861 ( .A(n8775), .ZN(n7747) );
  NAND2_X2 U4862 ( .A1(n6537), .A2(P1_U3086), .ZN(n7993) );
  XNOR2_X1 U4863 ( .A(n5819), .B(n5818), .ZN(n6718) );
  OR2_X1 U4864 ( .A1(n6201), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6212) );
  NAND2_X2 U4865 ( .A1(n4407), .A2(n4405), .ZN(n6536) );
  AND2_X1 U4866 ( .A1(n4939), .A2(n4343), .ZN(n4744) );
  XNOR2_X1 U4867 ( .A(n5042), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6832) );
  AND2_X1 U4868 ( .A1(n4746), .A2(n4940), .ZN(n4745) );
  NAND2_X1 U4869 ( .A1(n5810), .A2(n5809), .ZN(n6691) );
  INV_X1 U4870 ( .A(n5025), .ZN(n4936) );
  NAND2_X1 U4871 ( .A1(n5041), .A2(n4572), .ZN(n5025) );
  NAND2_X1 U4872 ( .A1(n4844), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n4993) );
  NAND4_X1 U4873 ( .A1(n5739), .A2(n4813), .A3(n4814), .A4(n4815), .ZN(n5817)
         );
  AND3_X1 U4874 ( .A1(n4973), .A2(n5230), .A3(n4964), .ZN(n4939) );
  AND2_X1 U4875 ( .A1(n4938), .A2(n5316), .ZN(n4746) );
  AND4_X1 U4876 ( .A1(n4956), .A2(n4955), .A3(n4957), .A4(n4975), .ZN(n4940)
         );
  INV_X1 U4877 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n4957) );
  INV_X1 U4878 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4956) );
  INV_X4 U4879 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U4880 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4955) );
  NOR2_X2 U4881 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5867) );
  NOR2_X1 U4882 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6185) );
  NOR2_X1 U4883 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4947) );
  NOR2_X2 U4884 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5041) );
  NOR2_X1 U4885 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5316) );
  INV_X1 U4886 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4813) );
  INV_X1 U4887 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5230) );
  NOR2_X1 U4888 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n4938) );
  INV_X1 U4889 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4814) );
  INV_X1 U4890 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4815) );
  NAND2_X1 U4891 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5129) );
  NOR2_X1 U4892 ( .A1(n7790), .A2(n7789), .ZN(n7788) );
  AOI21_X4 U4893 ( .B1(n8296), .B2(n7960), .A(n7959), .ZN(n8267) );
  AOI21_X2 U4894 ( .B1(n6612), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9743), .ZN(
        n9759) );
  AOI21_X2 U4895 ( .B1(n9796), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9791), .ZN(
        n9805) );
  NOR2_X1 U4896 ( .A1(n4896), .A2(n4639), .ZN(n4638) );
  INV_X1 U4897 ( .A(n4892), .ZN(n4639) );
  INV_X1 U4898 ( .A(n5245), .ZN(n4896) );
  OR2_X1 U4899 ( .A1(n8273), .A2(n8464), .ZN(n8160) );
  NOR2_X1 U4900 ( .A1(n6262), .A2(n4715), .ZN(n4714) );
  INV_X1 U4901 ( .A(n4717), .ZN(n4715) );
  INV_X1 U4902 ( .A(n5118), .ZN(n4950) );
  AND2_X1 U4903 ( .A1(n6529), .A2(n6937), .ZN(n4988) );
  OR2_X1 U4904 ( .A1(n5695), .A2(n9184), .ZN(n4987) );
  NAND2_X1 U4905 ( .A1(n9097), .A2(n9098), .ZN(n8950) );
  AOI21_X1 U4906 ( .B1(n5484), .B2(n4623), .A(n4621), .ZN(n4620) );
  INV_X1 U4907 ( .A(n5511), .ZN(n4621) );
  INV_X1 U4908 ( .A(n6058), .ZN(n9368) );
  MUX2_X1 U4909 ( .A(n9080), .B(n9079), .S(n9104), .Z(n9084) );
  OR2_X1 U4910 ( .A1(n8179), .A2(n8015), .ZN(n8017) );
  OR2_X1 U4911 ( .A1(n8245), .A2(n8288), .ZN(n8151) );
  AND2_X1 U4912 ( .A1(n5471), .A2(n4548), .ZN(n4547) );
  NAND2_X1 U4913 ( .A1(n8790), .A2(n8794), .ZN(n4548) );
  INV_X1 U4914 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4788) );
  INV_X1 U4915 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4943) );
  INV_X1 U4916 ( .A(n7983), .ZN(n4802) );
  NAND2_X1 U4917 ( .A1(n4369), .A2(n6554), .ZN(n5834) );
  OR2_X1 U4918 ( .A1(n8278), .A2(n8488), .ZN(n8144) );
  OR2_X1 U4919 ( .A1(n7688), .A2(n7731), .ZN(n8129) );
  OR2_X1 U4920 ( .A1(n7274), .A2(n6225), .ZN(n6229) );
  AND2_X1 U4921 ( .A1(n6183), .A2(n6182), .ZN(n7119) );
  OR2_X1 U4922 ( .A1(n6149), .A2(n6148), .ZN(n6183) );
  NAND2_X1 U4923 ( .A1(n5797), .A2(n5754), .ZN(n5787) );
  INV_X1 U4924 ( .A(n4420), .ZN(n4418) );
  AOI21_X1 U4925 ( .B1(n4550), .B2(n4551), .A(n4322), .ZN(n4549) );
  INV_X1 U4926 ( .A(n9205), .ZN(n7069) );
  INV_X1 U4927 ( .A(n4786), .ZN(n4784) );
  NAND2_X1 U4928 ( .A1(n5971), .A2(n5970), .ZN(n5982) );
  OR2_X1 U4929 ( .A1(n5985), .A2(n5967), .ZN(n5971) );
  NAND2_X1 U4930 ( .A1(n5600), .A2(n5599), .ZN(n5622) );
  NAND2_X1 U4931 ( .A1(n5571), .A2(n5570), .ZN(n5594) );
  NAND2_X1 U4932 ( .A1(n4626), .A2(n5480), .ZN(n4625) );
  INV_X1 U4933 ( .A(n5485), .ZN(n4626) );
  AND2_X1 U4934 ( .A1(n5457), .A2(n5442), .ZN(n5455) );
  INV_X1 U4935 ( .A(n5411), .ZN(n4612) );
  INV_X1 U4936 ( .A(n4611), .ZN(n4610) );
  OAI21_X1 U4937 ( .B1(n4614), .B2(n4292), .A(n5436), .ZN(n4611) );
  AND2_X1 U4938 ( .A1(n4923), .A2(n4922), .ZN(n5361) );
  OR2_X1 U4939 ( .A1(n4919), .A2(n5335), .ZN(n4923) );
  XNOR2_X1 U4940 ( .A(n4920), .B(SI_15_), .ZN(n5337) );
  AOI21_X1 U4941 ( .B1(n4631), .B2(n4633), .A(n4329), .ZN(n4630) );
  INV_X1 U4942 ( .A(n5189), .ZN(n4627) );
  NAND2_X1 U4943 ( .A1(n4897), .A2(n8682), .ZN(n4900) );
  NAND2_X1 U4944 ( .A1(n5189), .A2(n4638), .ZN(n4629) );
  NAND2_X1 U4945 ( .A1(n4889), .A2(n4888), .ZN(n4892) );
  OAI21_X1 U4946 ( .B1(n6536), .B2(n4857), .A(n4431), .ZN(n4860) );
  NAND2_X1 U4947 ( .A1(n6536), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4431) );
  NAND2_X1 U4948 ( .A1(n7969), .A2(n8455), .ZN(n4809) );
  NAND2_X1 U4949 ( .A1(n4603), .A2(n4310), .ZN(n4602) );
  AND2_X1 U4950 ( .A1(n6115), .A2(n6117), .ZN(n6211) );
  INV_X1 U4951 ( .A(n5874), .ZN(n4577) );
  NAND2_X1 U4952 ( .A1(n4649), .A2(n4648), .ZN(n7801) );
  NAND2_X1 U4953 ( .A1(n4653), .A2(n4652), .ZN(n4648) );
  OR2_X1 U4954 ( .A1(n8352), .A2(n4650), .ZN(n4649) );
  OAI211_X1 U4955 ( .C1(n7801), .C2(n4363), .A(n4362), .B(n4361), .ZN(n7776)
         );
  NAND2_X1 U4956 ( .A1(n4365), .A2(n4364), .ZN(n4362) );
  OR2_X1 U4957 ( .A1(n4365), .A2(n4364), .ZN(n4363) );
  NAND2_X1 U4958 ( .A1(n7801), .A2(n4364), .ZN(n4361) );
  OR2_X1 U4959 ( .A1(n7776), .A2(n7775), .ZN(n4663) );
  XNOR2_X1 U4960 ( .A(n8399), .B(n8404), .ZN(n8395) );
  OR2_X1 U4961 ( .A1(n6468), .A2(n6467), .ZN(n6469) );
  AOI22_X1 U4962 ( .A1(n8418), .A2(n6410), .B1(n8405), .B2(n8426), .ZN(n8403)
         );
  OR2_X1 U4963 ( .A1(n8442), .A2(n8455), .ZN(n8427) );
  NOR2_X1 U4964 ( .A1(n4294), .A2(n4727), .ZN(n4726) );
  OR2_X1 U4965 ( .A1(n8137), .A2(n8389), .ZN(n9710) );
  NAND2_X1 U4966 ( .A1(n6155), .A2(n6537), .ZN(n6207) );
  NOR2_X1 U4967 ( .A1(n5779), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5775) );
  AND2_X1 U4968 ( .A1(n5147), .A2(n5146), .ZN(n7207) );
  INV_X1 U4969 ( .A(n5092), .ZN(n5501) );
  INV_X1 U4970 ( .A(n5500), .ZN(n6094) );
  OR2_X1 U4971 ( .A1(n9659), .A2(n4281), .ZN(n5093) );
  OR2_X1 U4972 ( .A1(n9358), .A2(n9354), .ZN(n9349) );
  NOR2_X1 U4973 ( .A1(n9335), .A2(n9083), .ZN(n4793) );
  AOI21_X1 U4974 ( .B1(n4498), .B2(n4496), .A(n4325), .ZN(n4495) );
  INV_X1 U4975 ( .A(n4502), .ZN(n4496) );
  AOI21_X1 U4976 ( .B1(n4502), .B2(n4282), .A(n4302), .ZN(n4501) );
  OR2_X1 U4977 ( .A1(n9973), .A2(n6076), .ZN(n9137) );
  NAND2_X1 U4978 ( .A1(n6567), .A2(n6530), .ZN(n5064) );
  OR2_X1 U4979 ( .A1(n9410), .A2(n9179), .ZN(n6937) );
  INV_X1 U4982 ( .A(n5987), .ZN(n5419) );
  INV_X1 U4983 ( .A(n6567), .ZN(n5418) );
  XNOR2_X1 U4984 ( .A(n4946), .B(n4945), .ZN(n5995) );
  OAI21_X1 U4985 ( .B1(n4969), .B2(n4786), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4946) );
  INV_X1 U4986 ( .A(n4620), .ZN(n4619) );
  AND2_X1 U4987 ( .A1(n4618), .A2(n5518), .ZN(n4617) );
  NAND2_X1 U4988 ( .A1(n4963), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U4989 ( .A1(n5388), .A2(n4934), .ZN(n5413) );
  XNOR2_X1 U4990 ( .A(n4870), .B(SI_4_), .ZN(n5030) );
  NAND2_X1 U4991 ( .A1(n5044), .A2(n5043), .ZN(n4865) );
  INV_X1 U4992 ( .A(n9190), .ZN(n9409) );
  INV_X1 U4993 ( .A(n4516), .ZN(n6060) );
  OAI21_X1 U4994 ( .B1(n6056), .B2(n4512), .A(n4511), .ZN(n4516) );
  AOI21_X1 U4995 ( .B1(n4513), .B2(n9366), .A(n6059), .ZN(n4511) );
  OAI21_X1 U4996 ( .B1(n8974), .B2(n9111), .A(n4452), .ZN(n4451) );
  OAI21_X1 U4997 ( .B1(n8975), .B2(n9104), .A(n9850), .ZN(n4453) );
  OR2_X1 U4998 ( .A1(n8959), .A2(n9500), .ZN(n8957) );
  AND2_X1 U4999 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  NAND2_X1 U5000 ( .A1(n8347), .A2(n6168), .ZN(n8038) );
  AND2_X1 U5001 ( .A1(n5742), .A2(n5741), .ZN(n5743) );
  OAI21_X1 U5002 ( .B1(n9084), .B2(n9083), .A(n9082), .ZN(n9089) );
  INV_X1 U5003 ( .A(n6029), .ZN(n4487) );
  NOR2_X1 U5004 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4954) );
  AND2_X1 U5005 ( .A1(n5358), .A2(n4910), .ZN(n4906) );
  AND2_X1 U5006 ( .A1(n5334), .A2(n5337), .ZN(n5358) );
  OAI21_X1 U5007 ( .B1(n4388), .B2(P2_DATAO_REG_16__SCAN_IN), .A(n4397), .ZN(
        n4907) );
  NAND2_X1 U5008 ( .A1(n4388), .A2(n6657), .ZN(n4397) );
  OAI21_X1 U5009 ( .B1(n4388), .B2(P2_DATAO_REG_14__SCAN_IN), .A(n4390), .ZN(
        n4912) );
  NAND2_X1 U5010 ( .A1(n6537), .A2(n6664), .ZN(n4390) );
  OAI21_X1 U5011 ( .B1(n4388), .B2(n4395), .A(n4394), .ZN(n4911) );
  NAND2_X1 U5012 ( .A1(n4388), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n4394) );
  OAI21_X1 U5013 ( .B1(n4388), .B2(P2_DATAO_REG_10__SCAN_IN), .A(n4392), .ZN(
        n4893) );
  NAND2_X1 U5014 ( .A1(n4388), .A2(n6577), .ZN(n4392) );
  NAND2_X1 U5015 ( .A1(n4884), .A2(n4883), .ZN(n4887) );
  AND2_X1 U5016 ( .A1(n4299), .A2(n7966), .ZN(n4798) );
  INV_X1 U5017 ( .A(n7974), .ZN(n7961) );
  OR2_X1 U5018 ( .A1(n5871), .A2(n6538), .ZN(n4589) );
  INV_X1 U5019 ( .A(n5825), .ZN(n5827) );
  OR2_X1 U5020 ( .A1(n7903), .A2(n5881), .ZN(n5882) );
  NOR2_X1 U5021 ( .A1(n7857), .A2(n4371), .ZN(n5849) );
  NOR2_X1 U5022 ( .A1(n7862), .A2(n4372), .ZN(n4371) );
  OR2_X1 U5023 ( .A1(n7809), .A2(n5892), .ZN(n5894) );
  INV_X1 U5024 ( .A(n4696), .ZN(n4695) );
  OAI21_X1 U5025 ( .B1(n8410), .B2(n4697), .A(n6471), .ZN(n4696) );
  INV_X1 U5026 ( .A(n8020), .ZN(n4697) );
  OR2_X1 U5027 ( .A1(n8426), .A2(n8438), .ZN(n8022) );
  OR2_X1 U5028 ( .A1(n7498), .A2(n9711), .ZN(n8118) );
  INV_X1 U5029 ( .A(n4716), .ZN(n4708) );
  NAND2_X1 U5030 ( .A1(n7108), .A2(n7223), .ZN(n8040) );
  AND2_X1 U5031 ( .A1(n8038), .A2(n8040), .ZN(n6449) );
  NOR2_X1 U5032 ( .A1(n4685), .A2(n4684), .ZN(n4683) );
  INV_X1 U5033 ( .A(n8145), .ZN(n4685) );
  NAND2_X1 U5034 ( .A1(n4702), .A2(n4701), .ZN(n5779) );
  INV_X1 U5035 ( .A(n5774), .ZN(n4702) );
  INV_X1 U5036 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4408) );
  INV_X1 U5037 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4409) );
  AND2_X1 U5038 ( .A1(n5746), .A2(n4823), .ZN(n4822) );
  AND2_X1 U5039 ( .A1(n5743), .A2(n4838), .ZN(n4837) );
  INV_X1 U5040 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4838) );
  AND2_X1 U5041 ( .A1(n5821), .A2(n5740), .ZN(n5823) );
  INV_X1 U5042 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5740) );
  AND2_X1 U5043 ( .A1(n5592), .A2(n5730), .ZN(n4524) );
  AND2_X1 U5044 ( .A1(n4539), .A2(n4535), .ZN(n4531) );
  INV_X1 U5045 ( .A(n7602), .ZN(n4535) );
  INV_X1 U5046 ( .A(n4547), .ZN(n4546) );
  INV_X1 U5047 ( .A(n4544), .ZN(n4415) );
  AOI21_X1 U5048 ( .B1(n4547), .B2(n4545), .A(n4327), .ZN(n4544) );
  INV_X1 U5049 ( .A(n8794), .ZN(n4545) );
  NAND2_X1 U5050 ( .A1(n4528), .A2(n4530), .ZN(n4412) );
  NOR2_X1 U5051 ( .A1(n4529), .A2(n5333), .ZN(n4528) );
  INV_X1 U5052 ( .A(n4533), .ZN(n4529) );
  INV_X1 U5053 ( .A(n9101), .ZN(n9176) );
  OR2_X1 U5054 ( .A1(n9383), .A2(n6088), .ZN(n9077) );
  NOR2_X1 U5055 ( .A1(n9406), .A2(n9060), .ZN(n4769) );
  INV_X1 U5056 ( .A(n9068), .ZN(n4766) );
  NOR2_X1 U5057 ( .A1(n4499), .A2(n6047), .ZN(n4498) );
  INV_X1 U5058 ( .A(n4501), .ZN(n4499) );
  AOI21_X1 U5059 ( .B1(n6086), .B2(n8960), .A(n9440), .ZN(n4736) );
  AND2_X1 U5060 ( .A1(n6081), .A2(n4755), .ZN(n4754) );
  NAND2_X1 U5061 ( .A1(n8943), .A2(n4756), .ZN(n4755) );
  INV_X1 U5062 ( .A(n8943), .ZN(n4757) );
  OR2_X1 U5063 ( .A1(n7701), .A2(n8940), .ZN(n6078) );
  INV_X1 U5064 ( .A(n9137), .ZN(n4742) );
  INV_X1 U5065 ( .A(n8931), .ZN(n4776) );
  INV_X1 U5066 ( .A(n8993), .ZN(n4778) );
  NAND2_X1 U5067 ( .A1(n4456), .A2(n4311), .ZN(n6070) );
  INV_X1 U5068 ( .A(n9865), .ZN(n4456) );
  NAND2_X1 U5069 ( .A1(n9117), .A2(n6068), .ZN(n4762) );
  NOR2_X1 U5070 ( .A1(n6069), .A2(n4764), .ZN(n4763) );
  INV_X1 U5071 ( .A(n6068), .ZN(n4764) );
  INV_X1 U5072 ( .A(n9890), .ZN(n6017) );
  AOI21_X1 U5073 ( .B1(n8923), .B2(n6907), .A(n6064), .ZN(n6979) );
  AOI21_X1 U5074 ( .B1(n4791), .B2(n4793), .A(n4790), .ZN(n4789) );
  INV_X1 U5075 ( .A(n9095), .ZN(n4790) );
  INV_X1 U5076 ( .A(n6089), .ZN(n4791) );
  NAND2_X1 U5077 ( .A1(n4994), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4990) );
  INV_X1 U5078 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4787) );
  INV_X1 U5079 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4945) );
  NAND2_X1 U5080 ( .A1(n5628), .A2(n5627), .ZN(n5966) );
  NAND2_X1 U5081 ( .A1(n4640), .A2(n5563), .ZN(n5571) );
  NAND2_X1 U5082 ( .A1(n5561), .A2(n5562), .ZN(n4640) );
  NAND2_X1 U5083 ( .A1(n5538), .A2(n5537), .ZN(n5561) );
  AND3_X1 U5084 ( .A1(n4935), .A2(n4954), .A3(n4947), .ZN(n4937) );
  NOR2_X1 U5085 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4935) );
  NOR2_X1 U5086 ( .A1(n5412), .A2(n4615), .ZN(n4614) );
  INV_X1 U5087 ( .A(n4934), .ZN(n4615) );
  AND2_X1 U5088 ( .A1(n4924), .A2(n5361), .ZN(n5360) );
  XNOR2_X1 U5089 ( .A(n4893), .B(SI_10_), .ZN(n5245) );
  OAI21_X1 U5090 ( .B1(n5198), .B2(n5197), .A(n4887), .ZN(n5187) );
  AND2_X1 U5091 ( .A1(n4892), .A2(n4891), .ZN(n5186) );
  INV_X1 U5092 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4949) );
  AND2_X1 U5093 ( .A1(n4572), .A2(n4948), .ZN(n4570) );
  NAND2_X1 U5094 ( .A1(n4808), .A2(n8438), .ZN(n4807) );
  OR2_X1 U5095 ( .A1(n8319), .A2(n4809), .ZN(n4806) );
  INV_X1 U5096 ( .A(n7970), .ZN(n4808) );
  NOR2_X1 U5097 ( .A1(n4800), .A2(n8319), .ZN(n4799) );
  INV_X1 U5098 ( .A(n4804), .ZN(n4800) );
  NAND2_X1 U5099 ( .A1(n7041), .A2(n4834), .ZN(n7097) );
  AND2_X1 U5100 ( .A1(n7043), .A2(n7040), .ZN(n4834) );
  NAND2_X1 U5101 ( .A1(n6132), .A2(n6131), .ZN(n8442) );
  NAND2_X1 U5102 ( .A1(n4833), .A2(n6997), .ZN(n7011) );
  AND2_X1 U5103 ( .A1(n6998), .A2(n6996), .ZN(n4833) );
  NAND2_X1 U5104 ( .A1(n7305), .A2(n7304), .ZN(n7382) );
  NOR2_X1 U5105 ( .A1(n8308), .A2(n4828), .ZN(n4827) );
  INV_X1 U5106 ( .A(n4830), .ZN(n4828) );
  OR2_X1 U5107 ( .A1(n6795), .A2(n8225), .ZN(n6801) );
  AND4_X1 U5108 ( .A1(n8010), .A2(n8009), .A3(n8008), .A4(n8007), .ZN(n8373)
         );
  AND2_X1 U5109 ( .A1(n4375), .A2(n6700), .ZN(n4374) );
  OR2_X1 U5110 ( .A1(n6538), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4375) );
  NAND2_X1 U5111 ( .A1(n5875), .A2(n4580), .ZN(n4576) );
  NAND2_X1 U5112 ( .A1(n4578), .A2(n4581), .ZN(n4579) );
  AND2_X1 U5113 ( .A1(n5873), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4578) );
  OAI22_X1 U5114 ( .A1(n7927), .A2(n7926), .B1(n5913), .B2(n6554), .ZN(n7908)
         );
  NAND2_X1 U5115 ( .A1(n7908), .A2(n7907), .ZN(n7906) );
  OAI21_X1 U5116 ( .B1(n5882), .B2(n6571), .A(n5883), .ZN(n6964) );
  AOI21_X1 U5117 ( .B1(n5835), .B2(n4666), .A(n4347), .ZN(n4665) );
  OAI21_X1 U5118 ( .B1(n7877), .B2(n4668), .A(n4667), .ZN(n7857) );
  NAND2_X1 U5119 ( .A1(n4669), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4668) );
  NAND2_X1 U5120 ( .A1(n5847), .A2(n4669), .ZN(n4667) );
  INV_X1 U5121 ( .A(n7858), .ZN(n4669) );
  XNOR2_X1 U5122 ( .A(n5849), .B(n7843), .ZN(n7839) );
  OR2_X1 U5123 ( .A1(n7839), .A2(n9724), .ZN(n4370) );
  OR2_X1 U5124 ( .A1(n7846), .A2(n4584), .ZN(n4583) );
  NOR2_X1 U5125 ( .A1(n7862), .A2(n4585), .ZN(n4584) );
  AOI21_X1 U5126 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n6655), .A(n7788), .ZN(
        n5896) );
  NAND2_X1 U5127 ( .A1(n4663), .A2(n4296), .ZN(n4662) );
  NOR2_X1 U5128 ( .A1(n7801), .A2(n4365), .ZN(n5855) );
  NAND2_X1 U5129 ( .A1(n4595), .A2(n4594), .ZN(n4593) );
  INV_X1 U5130 ( .A(n5897), .ZN(n4594) );
  NAND2_X1 U5131 ( .A1(n5950), .A2(n8240), .ZN(n4384) );
  NAND2_X1 U5132 ( .A1(n8411), .A2(n8410), .ZN(n8409) );
  AND2_X1 U5133 ( .A1(n8022), .A2(n8023), .ZN(n8428) );
  OAI21_X1 U5134 ( .B1(n8459), .B2(n6463), .A(n8160), .ZN(n8448) );
  AOI21_X1 U5135 ( .B1(n4720), .B2(n4719), .A(n4321), .ZN(n4718) );
  INV_X1 U5136 ( .A(n6387), .ZN(n4719) );
  NAND2_X1 U5137 ( .A1(n8462), .A2(n6387), .ZN(n4723) );
  AND2_X1 U5138 ( .A1(n8498), .A2(n6349), .ZN(n4732) );
  NAND2_X1 U5139 ( .A1(n4300), .A2(n6348), .ZN(n8509) );
  OR2_X1 U5140 ( .A1(n8312), .A2(n7942), .ZN(n8517) );
  OAI21_X1 U5141 ( .B1(n7425), .B2(n4689), .A(n4688), .ZN(n7614) );
  NAND2_X1 U5142 ( .A1(n8124), .A2(n8129), .ZN(n4689) );
  NAND2_X1 U5143 ( .A1(n4691), .A2(n8129), .ZN(n4688) );
  OAI21_X1 U5144 ( .B1(n4731), .B2(n4730), .A(n4330), .ZN(n4729) );
  INV_X1 U5145 ( .A(n6315), .ZN(n4730) );
  INV_X1 U5146 ( .A(n7610), .ZN(n6459) );
  NAND2_X1 U5147 ( .A1(n7425), .A2(n8121), .ZN(n7427) );
  OR2_X1 U5148 ( .A1(n7315), .A2(n9709), .ZN(n8109) );
  INV_X1 U5149 ( .A(n4681), .ZN(n4680) );
  OAI21_X1 U5150 ( .B1(n8203), .B2(n4682), .A(n9707), .ZN(n4681) );
  INV_X1 U5151 ( .A(n8109), .ZN(n4682) );
  NAND2_X1 U5152 ( .A1(n6272), .A2(n6271), .ZN(n8113) );
  OR2_X1 U5153 ( .A1(n7315), .A2(n8337), .ZN(n4716) );
  NAND2_X1 U5154 ( .A1(n4710), .A2(n4288), .ZN(n4709) );
  AOI21_X1 U5155 ( .B1(n8197), .B2(n8091), .A(n4700), .ZN(n4699) );
  OR2_X1 U5156 ( .A1(n7440), .A2(n8197), .ZN(n7438) );
  NAND2_X1 U5157 ( .A1(n6232), .A2(n6231), .ZN(n4728) );
  INV_X1 U5158 ( .A(n8340), .ZN(n7278) );
  AND4_X1 U5159 ( .A1(n6218), .A2(n6217), .A3(n6216), .A4(n6215), .ZN(n6222)
         );
  AND3_X1 U5160 ( .A1(n6193), .A2(n6192), .A3(n6191), .ZN(n7005) );
  INV_X1 U5161 ( .A(n8069), .ZN(n4676) );
  INV_X1 U5162 ( .A(n4675), .ZN(n4674) );
  OAI21_X1 U5163 ( .B1(n8067), .B2(n4676), .A(n8060), .ZN(n4675) );
  INV_X1 U5164 ( .A(n9710), .ZN(n8512) );
  NAND2_X1 U5165 ( .A1(n7215), .A2(n8040), .ZN(n7104) );
  AND3_X1 U5166 ( .A1(n6178), .A2(n6177), .A3(n6176), .ZN(n8049) );
  NAND2_X1 U5167 ( .A1(n6427), .A2(n6426), .ZN(n8179) );
  INV_X1 U5168 ( .A(n8414), .ZN(n8537) );
  NAND2_X1 U5169 ( .A1(n6379), .A2(n6378), .ZN(n7962) );
  NAND2_X1 U5170 ( .A1(n6369), .A2(n6368), .ZN(n8029) );
  NAND2_X1 U5171 ( .A1(n8479), .A2(n8478), .ZN(n8560) );
  NAND2_X1 U5172 ( .A1(n6351), .A2(n6350), .ZN(n8278) );
  NAND2_X1 U5173 ( .A1(n6339), .A2(n6338), .ZN(n8236) );
  NAND2_X1 U5174 ( .A1(n6317), .A2(n6316), .ZN(n8582) );
  NAND2_X1 U5175 ( .A1(n6305), .A2(n6304), .ZN(n7688) );
  INV_X1 U5176 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6108) );
  AND2_X1 U5177 ( .A1(n5758), .A2(n4706), .ZN(n4705) );
  NOR2_X1 U5178 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n4706) );
  XNOR2_X1 U5179 ( .A(n5748), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U5180 ( .A1(n4818), .A2(n4817), .ZN(n5748) );
  AOI21_X1 U5181 ( .B1(n4820), .B2(n6109), .A(n6109), .ZN(n4817) );
  INV_X1 U5182 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4599) );
  INV_X1 U5183 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5739) );
  AOI21_X1 U5184 ( .B1(n6951), .B2(n4562), .A(n4312), .ZN(n4561) );
  NOR2_X1 U5185 ( .A1(n5591), .A2(n4287), .ZN(n4525) );
  OR2_X1 U5186 ( .A1(n5208), .A2(n5178), .ZN(n5250) );
  AOI21_X1 U5187 ( .B1(n4549), .B2(n4421), .A(n4305), .ZN(n4420) );
  INV_X1 U5188 ( .A(n4550), .ZN(n4421) );
  AOI22_X1 U5189 ( .A1(n9212), .A2(n4429), .B1(n6904), .B2(n4280), .ZN(n5080)
         );
  INV_X1 U5190 ( .A(n5547), .ZN(n5545) );
  NOR2_X1 U5191 ( .A1(n7087), .A2(n4563), .ZN(n4562) );
  INV_X1 U5192 ( .A(n4565), .ZN(n4563) );
  NAND2_X1 U5193 ( .A1(n5105), .A2(n4566), .ZN(n4565) );
  INV_X1 U5194 ( .A(n5106), .ZN(n4566) );
  NAND2_X1 U5195 ( .A1(n5461), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5498) );
  OAI21_X1 U5196 ( .B1(n7553), .B2(n5223), .A(n5222), .ZN(n5224) );
  XNOR2_X1 U5197 ( .A(n4567), .B(n5014), .ZN(n5084) );
  NAND2_X1 U5198 ( .A1(n5068), .A2(n4568), .ZN(n4567) );
  NAND2_X1 U5199 ( .A1(n4280), .A2(n6903), .ZN(n4568) );
  NAND2_X1 U5200 ( .A1(n5002), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5131) );
  INV_X1 U5201 ( .A(n5129), .ZN(n5002) );
  NAND2_X1 U5202 ( .A1(n9175), .A2(n9308), .ZN(n4441) );
  NAND2_X1 U5203 ( .A1(n9107), .A2(n4443), .ZN(n4442) );
  OAI21_X1 U5204 ( .B1(n9103), .B2(n9610), .A(n4454), .ZN(n9106) );
  AND4_X1 U5205 ( .A1(n5117), .A2(n5116), .A3(n5115), .A4(n5114), .ZN(n7230)
         );
  OR2_X1 U5206 ( .A1(n9659), .A2(n5052), .ZN(n5092) );
  NOR2_X1 U5207 ( .A1(n9323), .A2(n4471), .ZN(n4470) );
  OR2_X1 U5208 ( .A1(n4472), .A2(n9543), .ZN(n4471) );
  AND2_X1 U5209 ( .A1(n9618), .A2(n9396), .ZN(n9381) );
  AND2_X1 U5210 ( .A1(n9077), .A2(n9365), .ZN(n9375) );
  AND2_X1 U5211 ( .A1(n9416), .A2(n9432), .ZN(n6049) );
  NOR2_X1 U5212 ( .A1(n9421), .A2(n9416), .ZN(n9405) );
  NAND2_X1 U5213 ( .A1(n6087), .A2(n9427), .ZN(n9430) );
  INV_X1 U5214 ( .A(n4498), .ZN(n4497) );
  NOR2_X1 U5215 ( .A1(n6046), .A2(n4503), .ZN(n4502) );
  INV_X1 U5216 ( .A(n6045), .ZN(n4503) );
  INV_X1 U5217 ( .A(n5396), .ZN(n5007) );
  NAND2_X1 U5218 ( .A1(n4743), .A2(n6077), .ZN(n7645) );
  INV_X1 U5219 ( .A(n7643), .ZN(n4743) );
  OR2_X1 U5220 ( .A1(n9841), .A2(n9201), .ZN(n8995) );
  NAND2_X1 U5221 ( .A1(n4508), .A2(n4506), .ZN(n7397) );
  NAND2_X1 U5222 ( .A1(n4507), .A2(n9841), .ZN(n4506) );
  NAND2_X1 U5223 ( .A1(n6028), .A2(n4504), .ZN(n4508) );
  NOR2_X1 U5224 ( .A1(n4509), .A2(n4505), .ZN(n4504) );
  OR2_X1 U5225 ( .A1(n7398), .A2(n7523), .ZN(n7417) );
  NAND2_X1 U5226 ( .A1(n5004), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5252) );
  INV_X1 U5227 ( .A(n5250), .ZN(n5004) );
  AOI21_X1 U5228 ( .B1(n9847), .B2(n4490), .A(n4320), .ZN(n4489) );
  NAND2_X1 U5229 ( .A1(n6017), .A2(n6016), .ZN(n4484) );
  NAND2_X1 U5230 ( .A1(n5574), .A2(n5573), .ZN(n9553) );
  INV_X1 U5231 ( .A(n7363), .ZN(n9940) );
  AND3_X1 U5232 ( .A1(n5142), .A2(n5141), .A3(n5140), .ZN(n9934) );
  XNOR2_X1 U5233 ( .A(n5979), .B(n5978), .ZN(n8772) );
  OAI21_X1 U5234 ( .B1(n5982), .B2(n5981), .A(n5976), .ZN(n5979) );
  XNOR2_X1 U5235 ( .A(n5982), .B(n5981), .ZN(n7996) );
  XNOR2_X1 U5236 ( .A(n5561), .B(n5562), .ZN(n7299) );
  NAND2_X1 U5237 ( .A1(n5458), .A2(n5457), .ZN(n5485) );
  AOI21_X1 U5238 ( .B1(n4610), .B2(n4292), .A(n4609), .ZN(n4608) );
  INV_X1 U5239 ( .A(n5483), .ZN(n4624) );
  INV_X1 U5240 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4964) );
  XNOR2_X1 U5241 ( .A(n5338), .B(n5337), .ZN(n6665) );
  NAND2_X1 U5242 ( .A1(n4635), .A2(n4900), .ZN(n5267) );
  NAND2_X1 U5243 ( .A1(n4629), .A2(n4636), .ZN(n4635) );
  NAND2_X1 U5244 ( .A1(n4426), .A2(n4878), .ZN(n5168) );
  XNOR2_X1 U5245 ( .A(n4873), .B(SI_5_), .ZN(n5136) );
  XNOR2_X1 U5246 ( .A(n4866), .B(SI_3_), .ZN(n5094) );
  OAI21_X1 U5247 ( .B1(n5063), .B2(n4449), .A(n4861), .ZN(n5044) );
  XNOR2_X1 U5248 ( .A(n4862), .B(SI_2_), .ZN(n5043) );
  AND4_X1 U5250 ( .A1(n6303), .A2(n6302), .A3(n6301), .A4(n6300), .ZN(n7693)
         );
  INV_X1 U5251 ( .A(n8341), .ZN(n7442) );
  AND3_X1 U5252 ( .A1(n6365), .A2(n6364), .A3(n6363), .ZN(n8288) );
  NAND2_X1 U5253 ( .A1(n4810), .A2(n4809), .ZN(n4359) );
  NAND2_X1 U5254 ( .A1(n4801), .A2(n4804), .ZN(n4810) );
  AND2_X1 U5255 ( .A1(n6130), .A2(n6129), .ZN(n8455) );
  NOR2_X1 U5256 ( .A1(n6959), .A2(n10113), .ZN(n6958) );
  XNOR2_X1 U5257 ( .A(n4583), .B(n6636), .ZN(n7829) );
  NOR2_X1 U5258 ( .A1(n7829), .A2(n9718), .ZN(n7828) );
  OR2_X1 U5259 ( .A1(n8352), .A2(n8351), .ZN(n4651) );
  NAND2_X1 U5260 ( .A1(n4662), .A2(n4661), .ZN(n7762) );
  OR2_X1 U5261 ( .A1(n4662), .A2(n4661), .ZN(n4660) );
  INV_X1 U5262 ( .A(n4593), .ZN(n7753) );
  NAND2_X1 U5263 ( .A1(n4657), .A2(n4656), .ZN(n4655) );
  INV_X1 U5264 ( .A(n7763), .ZN(n4657) );
  NAND2_X1 U5265 ( .A1(n7764), .A2(n7765), .ZN(n4656) );
  INV_X1 U5266 ( .A(n8586), .ZN(n8376) );
  OR2_X1 U5267 ( .A1(n8387), .A2(n7526), .ZN(n6477) );
  AND2_X1 U5268 ( .A1(n6414), .A2(n6413), .ZN(n8399) );
  AND2_X1 U5269 ( .A1(n6402), .A2(n6401), .ZN(n8743) );
  NAND4_X1 U5270 ( .A1(n5759), .A2(n5775), .A3(n4705), .A4(n6108), .ZN(n8773)
         );
  NAND2_X1 U5271 ( .A1(n5784), .A2(n4316), .ZN(n4378) );
  AND2_X1 U5272 ( .A1(n6107), .A2(n4346), .ZN(n4376) );
  NAND2_X1 U5273 ( .A1(n5323), .A2(n5322), .ZN(n9973) );
  NAND2_X1 U5274 ( .A1(n5521), .A2(n5520), .ZN(n9563) );
  NOR2_X1 U5275 ( .A1(n6854), .A2(n6855), .ZN(n6853) );
  OAI211_X1 U5276 ( .C1(n5064), .C2(n6541), .A(n5032), .B(n4314), .ZN(n9927)
         );
  NAND2_X1 U5277 ( .A1(n4966), .A2(n4965), .ZN(n9520) );
  NAND2_X1 U5278 ( .A1(n8885), .A2(n8886), .ZN(n8884) );
  NAND2_X1 U5279 ( .A1(n5585), .A2(n5584), .ZN(n9190) );
  NAND2_X1 U5280 ( .A1(n5530), .A2(n5529), .ZN(n9065) );
  OR2_X1 U5281 ( .A1(n5303), .A2(n5302), .ZN(n9199) );
  INV_X1 U5282 ( .A(n7539), .ZN(n9200) );
  NAND2_X1 U5283 ( .A1(n4794), .A2(n4793), .ZN(n9338) );
  NOR2_X1 U5284 ( .A1(n9345), .A2(n9344), .ZN(n9539) );
  AND2_X1 U5285 ( .A1(n4515), .A2(n4513), .ZN(n9345) );
  AND2_X1 U5286 ( .A1(n9343), .A2(n9342), .ZN(n9344) );
  NAND2_X1 U5287 ( .A1(n4515), .A2(n6057), .ZN(n9343) );
  OR2_X1 U5288 ( .A1(n9900), .A2(n6887), .ZN(n9526) );
  INV_X1 U5289 ( .A(n9351), .ZN(n9896) );
  NOR2_X1 U5290 ( .A1(n9330), .A2(n4773), .ZN(n4772) );
  INV_X1 U5291 ( .A(n6100), .ZN(n4773) );
  NAND2_X1 U5292 ( .A1(n4557), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4976) );
  INV_X1 U5293 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U5294 ( .A1(n4450), .A2(n8984), .ZN(n8992) );
  NOR2_X1 U5295 ( .A1(n4448), .A2(n9055), .ZN(n4446) );
  AND2_X1 U5296 ( .A1(n9046), .A2(n9057), .ZN(n4445) );
  OR2_X1 U5297 ( .A1(n9064), .A2(n9104), .ZN(n4355) );
  OR2_X1 U5298 ( .A1(n6464), .A2(n8428), .ZN(n6466) );
  INV_X1 U5299 ( .A(n8152), .ZN(n4684) );
  AND2_X1 U5300 ( .A1(n7551), .A2(n7453), .ZN(n5221) );
  NOR2_X1 U5301 ( .A1(n9500), .A2(n9484), .ZN(n4466) );
  INV_X1 U5302 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n4748) );
  AOI21_X1 U5303 ( .B1(n5966), .B2(n5965), .A(n4853), .ZN(n5969) );
  OAI21_X1 U5304 ( .B1(n4388), .B2(P2_DATAO_REG_25__SCAN_IN), .A(n4404), .ZN(
        n5565) );
  NAND2_X1 U5305 ( .A1(n4388), .A2(n7751), .ZN(n4404) );
  OAI21_X1 U5306 ( .B1(n4388), .B2(P2_DATAO_REG_22__SCAN_IN), .A(n4402), .ZN(
        n5487) );
  NAND2_X1 U5307 ( .A1(n4388), .A2(n7082), .ZN(n4402) );
  OAI21_X1 U5308 ( .B1(n4388), .B2(P2_DATAO_REG_21__SCAN_IN), .A(n4401), .ZN(
        n5481) );
  NAND2_X1 U5309 ( .A1(n4388), .A2(n6948), .ZN(n4401) );
  OAI21_X1 U5310 ( .B1(n4388), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n4403), .ZN(
        n5440) );
  NAND2_X1 U5311 ( .A1(n4388), .A2(n6916), .ZN(n4403) );
  OAI21_X1 U5312 ( .B1(n4388), .B2(P2_DATAO_REG_19__SCAN_IN), .A(n4399), .ZN(
        n5415) );
  NAND2_X1 U5313 ( .A1(n4388), .A2(n6899), .ZN(n4399) );
  OAI21_X1 U5314 ( .B1(n4388), .B2(P2_DATAO_REG_18__SCAN_IN), .A(n4398), .ZN(
        n5409) );
  NAND2_X1 U5315 ( .A1(n4388), .A2(n6693), .ZN(n4398) );
  OAI21_X1 U5316 ( .B1(n4388), .B2(P2_DATAO_REG_17__SCAN_IN), .A(n4400), .ZN(
        n4929) );
  NAND2_X1 U5317 ( .A1(n4388), .A2(n6652), .ZN(n4400) );
  OAI21_X1 U5318 ( .B1(n4388), .B2(P2_DATAO_REG_15__SCAN_IN), .A(n4393), .ZN(
        n4920) );
  NAND2_X1 U5319 ( .A1(n4388), .A2(n6666), .ZN(n4393) );
  INV_X1 U5320 ( .A(n4638), .ZN(n4628) );
  INV_X1 U5321 ( .A(n4633), .ZN(n4632) );
  NOR2_X1 U5322 ( .A1(n4903), .A2(n4634), .ZN(n4633) );
  INV_X1 U5323 ( .A(n4900), .ZN(n4634) );
  INV_X1 U5324 ( .A(n5268), .ZN(n4903) );
  INV_X1 U5325 ( .A(n4636), .ZN(n4631) );
  OAI21_X1 U5326 ( .B1(n4388), .B2(P2_DATAO_REG_12__SCAN_IN), .A(n4391), .ZN(
        n4901) );
  NAND2_X1 U5327 ( .A1(n4388), .A2(n6631), .ZN(n4391) );
  OAI21_X1 U5328 ( .B1(n4388), .B2(P2_DATAO_REG_11__SCAN_IN), .A(n4396), .ZN(
        n4897) );
  NAND2_X1 U5329 ( .A1(n4388), .A2(n8631), .ZN(n4396) );
  OR2_X1 U5330 ( .A1(n6804), .A2(n8183), .ZN(n6807) );
  NOR2_X1 U5331 ( .A1(n6394), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U5332 ( .A1(n8182), .A2(n8176), .ZN(n4606) );
  OR2_X1 U5333 ( .A1(n8181), .A2(n4605), .ZN(n4604) );
  NAND2_X1 U5334 ( .A1(n8217), .A2(n8137), .ZN(n4605) );
  OAI21_X1 U5335 ( .B1(n6675), .B2(n7583), .A(n4377), .ZN(n5901) );
  NAND2_X1 U5336 ( .A1(n7583), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4377) );
  NAND2_X1 U5337 ( .A1(n4367), .A2(n4366), .ZN(n4369) );
  AOI21_X1 U5338 ( .B1(n5827), .B2(n4368), .A(n4333), .ZN(n4366) );
  INV_X1 U5339 ( .A(n6722), .ZN(n4368) );
  INV_X1 U5340 ( .A(n7914), .ZN(n4666) );
  AOI21_X1 U5341 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n6578), .A(n7889), .ZN(
        n5846) );
  NOR2_X1 U5342 ( .A1(n7868), .A2(n5923), .ZN(n7851) );
  NOR2_X1 U5343 ( .A1(n7851), .A2(n7852), .ZN(n7850) );
  INV_X1 U5344 ( .A(n7802), .ZN(n4652) );
  NAND2_X1 U5345 ( .A1(n4652), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4650) );
  AND2_X1 U5346 ( .A1(n6655), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4365) );
  NAND2_X1 U5347 ( .A1(n4592), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4591) );
  OR2_X1 U5348 ( .A1(n8236), .A2(n8286), .ZN(n8033) );
  AND2_X1 U5349 ( .A1(n8207), .A2(n6293), .ZN(n4731) );
  INV_X1 U5350 ( .A(n8103), .ZN(n4700) );
  AOI21_X1 U5351 ( .B1(n4713), .B2(n4712), .A(n4306), .ZN(n4711) );
  INV_X1 U5352 ( .A(n6262), .ZN(n4713) );
  AND2_X1 U5353 ( .A1(n6253), .A2(n4717), .ZN(n4712) );
  INV_X1 U5354 ( .A(n6233), .ZN(n4727) );
  AND2_X1 U5355 ( .A1(n7155), .A2(n6229), .ZN(n6226) );
  OR2_X1 U5356 ( .A1(n7551), .A2(n7453), .ZN(n5217) );
  AND2_X1 U5357 ( .A1(n9606), .A2(n8916), .ZN(n9101) );
  NAND2_X1 U5358 ( .A1(n9094), .A2(n9093), .ZN(n4455) );
  OR2_X1 U5359 ( .A1(n9323), .A2(n9104), .ZN(n4454) );
  OR2_X1 U5360 ( .A1(n5093), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6015) );
  OR2_X1 U5361 ( .A1(n6105), .A2(n9339), .ZN(n9097) );
  NAND2_X1 U5362 ( .A1(n4474), .A2(n4473), .ZN(n4472) );
  OR2_X1 U5363 ( .A1(n9354), .A2(n6058), .ZN(n9091) );
  NAND2_X1 U5364 ( .A1(n9553), .A2(n9409), .ZN(n9074) );
  INV_X1 U5365 ( .A(n6027), .ZN(n4505) );
  NOR2_X1 U5366 ( .A1(n9841), .A2(n4510), .ZN(n4509) );
  NOR2_X1 U5367 ( .A1(n7324), .A2(n7574), .ZN(n7293) );
  AND2_X1 U5368 ( .A1(n4284), .A2(n9953), .ZN(n4469) );
  INV_X1 U5369 ( .A(n6022), .ZN(n4490) );
  NAND2_X1 U5370 ( .A1(n6943), .A2(n9208), .ZN(n4477) );
  OR2_X1 U5371 ( .A1(n9893), .A2(n9927), .ZN(n6942) );
  AND2_X1 U5372 ( .A1(n9405), .A2(n9401), .ZN(n9396) );
  NAND2_X1 U5373 ( .A1(n9518), .A2(n4466), .ZN(n9482) );
  NAND2_X1 U5374 ( .A1(n7648), .A2(n4283), .ZN(n7707) );
  NAND2_X1 U5375 ( .A1(n4485), .A2(n6032), .ZN(n7647) );
  NOR2_X1 U5376 ( .A1(n6031), .A2(n4487), .ZN(n4486) );
  XNOR2_X1 U5377 ( .A(n5969), .B(n5968), .ZN(n5985) );
  NAND2_X1 U5378 ( .A1(n5622), .A2(n5621), .ZN(n5628) );
  NAND2_X1 U5379 ( .A1(n5594), .A2(n5593), .ZN(n5600) );
  NAND2_X1 U5380 ( .A1(n4943), .A2(n4788), .ZN(n4785) );
  NAND2_X1 U5381 ( .A1(n4620), .A2(n4622), .ZN(n4618) );
  INV_X1 U5382 ( .A(n5455), .ZN(n4609) );
  OR2_X1 U5383 ( .A1(n4925), .A2(n5360), .ZN(n4926) );
  OR2_X1 U5384 ( .A1(n4918), .A2(n4917), .ZN(n5335) );
  AND2_X1 U5385 ( .A1(n5311), .A2(n4916), .ZN(n4917) );
  AND2_X1 U5386 ( .A1(n5310), .A2(n4915), .ZN(n5334) );
  NOR2_X1 U5387 ( .A1(n5227), .A2(n4637), .ZN(n4636) );
  INV_X1 U5388 ( .A(n4895), .ZN(n4637) );
  INV_X1 U5389 ( .A(n4425), .ZN(n4424) );
  OAI21_X1 U5390 ( .B1(n4878), .B2(n5167), .A(n4881), .ZN(n4425) );
  NAND2_X1 U5391 ( .A1(n4887), .A2(n4886), .ZN(n5197) );
  OAI21_X1 U5392 ( .B1(n4388), .B2(P2_DATAO_REG_6__SCAN_IN), .A(n4389), .ZN(
        n4876) );
  NAND2_X1 U5393 ( .A1(n6537), .A2(n6549), .ZN(n4389) );
  AND2_X1 U5394 ( .A1(n7951), .A2(n8279), .ZN(n8238) );
  NAND2_X1 U5395 ( .A1(n4797), .A2(n4795), .ZN(n7982) );
  NAND2_X1 U5396 ( .A1(n4299), .A2(n4796), .ZN(n4795) );
  INV_X1 U5397 ( .A(n4799), .ZN(n4796) );
  AND2_X1 U5398 ( .A1(n6213), .A2(n7098), .ZN(n6237) );
  NAND2_X1 U5399 ( .A1(n6237), .A2(n6236), .ZN(n6247) );
  NAND2_X1 U5400 ( .A1(n8238), .A2(n8286), .ZN(n8237) );
  NOR2_X1 U5401 ( .A1(n6265), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6274) );
  INV_X1 U5402 ( .A(n8338), .ZN(n7385) );
  OR2_X1 U5403 ( .A1(n6256), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U5404 ( .A1(n7940), .A2(n8332), .ZN(n4830) );
  NAND2_X1 U5405 ( .A1(n4832), .A2(n8311), .ZN(n4831) );
  INV_X1 U5406 ( .A(n7940), .ZN(n4832) );
  OR2_X1 U5407 ( .A1(n6329), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6343) );
  AND2_X1 U5408 ( .A1(n8259), .A2(n4805), .ZN(n4804) );
  NAND2_X1 U5409 ( .A1(n7967), .A2(n7966), .ZN(n4805) );
  AND4_X1 U5410 ( .A1(n6334), .A2(n6333), .A3(n6332), .A4(n6331), .ZN(n7942)
         );
  AND4_X1 U5411 ( .A1(n6190), .A2(n6189), .A3(n6188), .A4(n6187), .ZN(n7025)
         );
  OAI21_X1 U5412 ( .B1(n6679), .B2(n10097), .A(n5812), .ZN(n10017) );
  OR2_X1 U5413 ( .A1(n5816), .A2(n6538), .ZN(n4670) );
  NAND2_X1 U5414 ( .A1(n4589), .A2(n6706), .ZN(n6747) );
  NAND2_X1 U5415 ( .A1(n4586), .A2(n6706), .ZN(n6745) );
  INV_X1 U5416 ( .A(n4587), .ZN(n4586) );
  NOR2_X1 U5417 ( .A1(n6759), .A2(n10105), .ZN(n6758) );
  NOR2_X1 U5418 ( .A1(n6758), .A2(n5827), .ZN(n6723) );
  NOR2_X1 U5419 ( .A1(n6719), .A2(n4379), .ZN(n7927) );
  AND2_X1 U5420 ( .A1(n5912), .A2(n6734), .ZN(n4379) );
  NAND2_X1 U5421 ( .A1(n7906), .A2(n5915), .ZN(n6971) );
  CLKBUF_X1 U5422 ( .A(n5805), .Z(n5806) );
  NOR2_X1 U5423 ( .A1(n6958), .A2(n5845), .ZN(n7891) );
  XNOR2_X1 U5424 ( .A(n5846), .B(n7881), .ZN(n7877) );
  NOR2_X1 U5425 ( .A1(n7896), .A2(n5920), .ZN(n7869) );
  NOR2_X1 U5426 ( .A1(n7869), .A2(n7870), .ZN(n7868) );
  OAI21_X1 U5427 ( .B1(n6962), .B2(n4597), .A(n4596), .ZN(n5886) );
  NAND2_X1 U5428 ( .A1(n7884), .A2(n4598), .ZN(n4596) );
  NAND2_X1 U5429 ( .A1(n5883), .A2(n4598), .ZN(n4597) );
  NAND2_X1 U5430 ( .A1(n6578), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4598) );
  NOR2_X1 U5431 ( .A1(n7877), .A2(n10117), .ZN(n7876) );
  AND2_X1 U5432 ( .A1(n5830), .A2(n4836), .ZN(n5797) );
  AND2_X1 U5433 ( .A1(n4837), .A2(n4338), .ZN(n4836) );
  AND2_X1 U5434 ( .A1(n4308), .A2(n4370), .ZN(n7821) );
  NOR2_X1 U5435 ( .A1(n7831), .A2(n5931), .ZN(n7813) );
  NOR2_X1 U5436 ( .A1(n7813), .A2(n7814), .ZN(n7812) );
  NOR2_X1 U5437 ( .A1(n7812), .A2(n5935), .ZN(n8355) );
  NOR2_X1 U5438 ( .A1(n8355), .A2(n8356), .ZN(n8354) );
  OR2_X1 U5439 ( .A1(n7769), .A2(n7770), .ZN(n4595) );
  INV_X1 U5440 ( .A(n7761), .ZN(n4661) );
  AOI21_X1 U5441 ( .B1(n4695), .B2(n4697), .A(n4323), .ZN(n4694) );
  AOI21_X1 U5442 ( .B1(n6424), .B2(n6423), .A(n4845), .ZN(n6432) );
  NOR2_X1 U5443 ( .A1(n6380), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6392) );
  AND2_X1 U5444 ( .A1(n6376), .A2(n6375), .ZN(n8489) );
  NOR2_X1 U5445 ( .A1(n6343), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6352) );
  AND2_X1 U5446 ( .A1(n8033), .A2(n8141), .ZN(n8519) );
  NAND2_X1 U5447 ( .A1(n4277), .A2(n6335), .ZN(n7676) );
  NAND2_X1 U5448 ( .A1(n6319), .A2(n6318), .ZN(n6329) );
  NAND2_X1 U5449 ( .A1(n7485), .A2(n4731), .ZN(n7506) );
  AND2_X1 U5450 ( .A1(n7485), .A2(n6293), .ZN(n7428) );
  NAND2_X1 U5451 ( .A1(n4679), .A2(n4677), .ZN(n7490) );
  AOI21_X1 U5452 ( .B1(n4680), .B2(n4682), .A(n4678), .ZN(n4677) );
  INV_X1 U5453 ( .A(n8114), .ZN(n4678) );
  AND2_X1 U5454 ( .A1(n8118), .A2(n8119), .ZN(n8205) );
  NAND2_X1 U5455 ( .A1(n4709), .A2(n4707), .ZN(n6282) );
  NOR2_X1 U5456 ( .A1(n6280), .A2(n4708), .ZN(n4707) );
  NAND2_X1 U5457 ( .A1(n6292), .A2(n6291), .ZN(n7485) );
  AND4_X1 U5458 ( .A1(n6290), .A2(n6289), .A3(n6288), .A4(n6287), .ZN(n9711)
         );
  NAND2_X1 U5459 ( .A1(n4710), .A2(n4711), .ZN(n7252) );
  NAND2_X1 U5460 ( .A1(n4733), .A2(n6224), .ZN(n7274) );
  NOR2_X1 U5461 ( .A1(n6212), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6213) );
  INV_X1 U5462 ( .A(n4855), .ZN(n8194) );
  AND3_X1 U5463 ( .A1(n6210), .A2(n6209), .A3(n6208), .ZN(n6454) );
  NAND2_X1 U5464 ( .A1(n4673), .A2(n4671), .ZN(n7260) );
  AOI21_X1 U5465 ( .B1(n4674), .B2(n4676), .A(n4672), .ZN(n4671) );
  INV_X1 U5466 ( .A(n8068), .ZN(n4672) );
  XNOR2_X1 U5467 ( .A(n8346), .B(n8049), .ZN(n7107) );
  NAND2_X1 U5468 ( .A1(n6448), .A2(n6449), .ZN(n7215) );
  INV_X1 U5469 ( .A(n6449), .ZN(n8043) );
  INV_X1 U5470 ( .A(n8399), .ZN(n8533) );
  NAND2_X1 U5471 ( .A1(n6390), .A2(n6389), .ZN(n8273) );
  NAND2_X1 U5472 ( .A1(n6359), .A2(n6358), .ZN(n8245) );
  NAND2_X1 U5473 ( .A1(n6284), .A2(n6283), .ZN(n7498) );
  INV_X1 U5474 ( .A(n10068), .ZN(n10028) );
  CLKBUF_X1 U5475 ( .A(n6487), .Z(n6509) );
  AND2_X1 U5476 ( .A1(n5758), .A2(n5780), .ZN(n4704) );
  AND2_X1 U5477 ( .A1(n5781), .A2(n5780), .ZN(n5782) );
  INV_X1 U5478 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4406) );
  INV_X1 U5479 ( .A(n4821), .ZN(n4820) );
  OAI21_X1 U5480 ( .B1(n4822), .B2(n6109), .A(n5747), .ZN(n4821) );
  NOR2_X1 U5481 ( .A1(n5867), .A2(n6109), .ZN(n4600) );
  INV_X1 U5482 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U5483 ( .A1(n4517), .A2(n4518), .ZN(n4521) );
  INV_X1 U5484 ( .A(n4522), .ZN(n4518) );
  OAI21_X1 U5485 ( .B1(n4525), .B2(n4523), .A(n5648), .ZN(n4522) );
  AOI21_X1 U5486 ( .B1(n4531), .B2(n4534), .A(n4326), .ZN(n4533) );
  INV_X1 U5487 ( .A(n4537), .ZN(n4534) );
  NAND2_X1 U5488 ( .A1(n4416), .A2(n4414), .ZN(n5509) );
  AOI21_X1 U5489 ( .B1(n4417), .B2(n4422), .A(n4415), .ZN(n4414) );
  NOR2_X1 U5490 ( .A1(n4546), .A2(n4418), .ZN(n4417) );
  INV_X1 U5491 ( .A(n4549), .ZN(n4422) );
  INV_X1 U5492 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5205) );
  AND2_X1 U5493 ( .A1(n5265), .A2(n5264), .ZN(n4543) );
  INV_X1 U5494 ( .A(n5078), .ZN(n5079) );
  OAI22_X1 U5495 ( .A1(n6891), .A2(n5642), .B1(n6529), .B2(n9730), .ZN(n5078)
         );
  NAND2_X1 U5496 ( .A1(n5005), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5298) );
  INV_X1 U5497 ( .A(n5276), .ZN(n5005) );
  OR2_X1 U5498 ( .A1(n4541), .A2(n4334), .ZN(n4539) );
  AOI21_X1 U5499 ( .B1(n4543), .B2(n5266), .A(n4542), .ZN(n4541) );
  INV_X1 U5500 ( .A(n7517), .ZN(n4542) );
  NOR2_X1 U5501 ( .A1(n4538), .A2(n4334), .ZN(n4537) );
  INV_X1 U5502 ( .A(n4543), .ZN(n4538) );
  NAND2_X1 U5503 ( .A1(n5496), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5522) );
  XNOR2_X1 U5504 ( .A(n5509), .B(n5507), .ZN(n8851) );
  XNOR2_X1 U5505 ( .A(n4427), .B(n5666), .ZN(n7625) );
  NAND2_X1 U5506 ( .A1(n4430), .A2(n4428), .ZN(n4427) );
  NAND2_X1 U5507 ( .A1(n4510), .A2(n4429), .ZN(n4428) );
  NAND2_X1 U5508 ( .A1(n9841), .A2(n5047), .ZN(n4430) );
  NAND2_X1 U5509 ( .A1(n4556), .A2(n5385), .ZN(n4551) );
  OR2_X1 U5510 ( .A1(n4553), .A2(n4850), .ZN(n4550) );
  AND2_X1 U5511 ( .A1(n8829), .A2(n4554), .ZN(n4553) );
  OR2_X1 U5512 ( .A1(n4555), .A2(n8819), .ZN(n4554) );
  NAND2_X1 U5513 ( .A1(n5003), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5159) );
  INV_X1 U5514 ( .A(n5131), .ZN(n5003) );
  NAND2_X1 U5515 ( .A1(n4413), .A2(n4410), .ZN(n5355) );
  NAND2_X1 U5516 ( .A1(n4412), .A2(n4411), .ZN(n4410) );
  NAND2_X1 U5517 ( .A1(n7636), .A2(n5333), .ZN(n4413) );
  INV_X1 U5518 ( .A(n7633), .ZN(n4411) );
  INV_X1 U5519 ( .A(n5016), .ZN(n5612) );
  OR2_X1 U5520 ( .A1(n9173), .A2(n9172), .ZN(n4434) );
  INV_X1 U5521 ( .A(n9177), .ZN(n4439) );
  INV_X1 U5522 ( .A(n5704), .ZN(n5632) );
  AND4_X1 U5523 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n7287)
         );
  OR2_X1 U5524 ( .A1(n5093), .A2(n5034), .ZN(n5040) );
  AND2_X1 U5525 ( .A1(n9247), .A2(n9248), .ZN(n9245) );
  AOI21_X1 U5526 ( .B1(n6613), .B2(P1_REG2_REG_6__SCAN_IN), .A(n9758), .ZN(
        n9680) );
  AOI21_X1 U5527 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n9683), .A(n9678), .ZN(
        n9693) );
  AND2_X1 U5528 ( .A1(n9688), .A2(n9687), .ZN(n9690) );
  NOR2_X1 U5529 ( .A1(n9267), .A2(n9815), .ZN(n9269) );
  AND2_X1 U5530 ( .A1(n4960), .A2(n4949), .ZN(n4569) );
  AND2_X1 U5531 ( .A1(n9294), .A2(n9293), .ZN(n9830) );
  AND2_X1 U5532 ( .A1(n9354), .A2(n9368), .ZN(n6059) );
  INV_X1 U5533 ( .A(n4513), .ZN(n4512) );
  NOR2_X1 U5534 ( .A1(n9358), .A2(n4472), .ZN(n9319) );
  NAND2_X1 U5535 ( .A1(n4794), .A2(n9090), .ZN(n9336) );
  NOR2_X1 U5536 ( .A1(n9342), .A2(n4514), .ZN(n4513) );
  INV_X1 U5537 ( .A(n6057), .ZN(n4514) );
  AOI21_X1 U5538 ( .B1(n4769), .B2(n4767), .A(n4766), .ZN(n4765) );
  INV_X1 U5539 ( .A(n4769), .ZN(n4768) );
  AND2_X1 U5540 ( .A1(n5604), .A2(n5577), .ZN(n9398) );
  AND2_X1 U5541 ( .A1(n9073), .A2(n9074), .ZN(n9393) );
  NAND2_X1 U5542 ( .A1(n4494), .A2(n4492), .ZN(n9412) );
  AND2_X1 U5543 ( .A1(n4493), .A2(n6048), .ZN(n4492) );
  AND2_X1 U5544 ( .A1(n9518), .A2(n4462), .ZN(n9449) );
  NOR2_X1 U5545 ( .A1(n4464), .A2(n9450), .ZN(n4462) );
  NAND2_X1 U5546 ( .A1(n9449), .A2(n9426), .ZN(n9421) );
  NAND2_X1 U5547 ( .A1(n4735), .A2(n4734), .ZN(n9443) );
  AOI21_X1 U5548 ( .B1(n4736), .B2(n4737), .A(n9052), .ZN(n4734) );
  INV_X1 U5549 ( .A(n6086), .ZN(n4737) );
  NAND2_X1 U5550 ( .A1(n6084), .A2(n8905), .ZN(n9460) );
  NAND2_X1 U5551 ( .A1(n4753), .A2(n4751), .ZN(n9491) );
  AOI21_X1 U5552 ( .B1(n4754), .B2(n4757), .A(n4752), .ZN(n4751) );
  INV_X1 U5553 ( .A(n9148), .ZN(n4752) );
  AND2_X1 U5554 ( .A1(n9517), .A2(n9640), .ZN(n9518) );
  NAND2_X1 U5555 ( .A1(n9518), .A2(n9636), .ZN(n9497) );
  OR2_X1 U5556 ( .A1(n5373), .A2(n5372), .ZN(n5396) );
  NAND2_X1 U5557 ( .A1(n6078), .A2(n9141), .ZN(n7742) );
  NAND2_X1 U5558 ( .A1(n7742), .A2(n8943), .ZN(n9511) );
  AND2_X1 U5559 ( .A1(n7648), .A2(n4459), .ZN(n9517) );
  AND2_X1 U5560 ( .A1(n4285), .A2(n4460), .ZN(n4459) );
  NAND2_X1 U5561 ( .A1(n7648), .A2(n4285), .ZN(n7739) );
  AOI21_X1 U5562 ( .B1(n8938), .B2(n4741), .A(n4740), .ZN(n4739) );
  INV_X1 U5563 ( .A(n8962), .ZN(n4740) );
  NAND2_X1 U5564 ( .A1(n5006), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5373) );
  INV_X1 U5565 ( .A(n5346), .ZN(n5006) );
  AND2_X1 U5566 ( .A1(n7648), .A2(n7650), .ZN(n7659) );
  NOR2_X1 U5567 ( .A1(n7417), .A2(n9005), .ZN(n7648) );
  NOR2_X1 U5568 ( .A1(n6071), .A2(n4780), .ZN(n4779) );
  NAND2_X1 U5569 ( .A1(n8966), .A2(n8993), .ZN(n4780) );
  NAND2_X1 U5570 ( .A1(n4781), .A2(n6070), .ZN(n9128) );
  NOR2_X1 U5571 ( .A1(n6071), .A2(n4782), .ZN(n4781) );
  NAND3_X1 U5572 ( .A1(n9873), .A2(n4468), .A3(n4469), .ZN(n7324) );
  NAND2_X1 U5573 ( .A1(n9873), .A2(n4469), .ZN(n7322) );
  AND4_X1 U5574 ( .A1(n5257), .A2(n5256), .A3(n5255), .A4(n5254), .ZN(n7540)
         );
  NAND2_X1 U5575 ( .A1(n9873), .A2(n4284), .ZN(n9859) );
  NAND2_X1 U5576 ( .A1(n4491), .A2(n6022), .ZN(n9849) );
  NAND2_X1 U5577 ( .A1(n7072), .A2(n7073), .ZN(n4491) );
  AND2_X1 U5578 ( .A1(n9873), .A2(n9940), .ZN(n9860) );
  NAND2_X1 U5579 ( .A1(n4758), .A2(n4760), .ZN(n9865) );
  INV_X1 U5580 ( .A(n4761), .ZN(n4760) );
  OAI21_X1 U5581 ( .B1(n6069), .B2(n4762), .A(n9121), .ZN(n4761) );
  NOR2_X1 U5582 ( .A1(n6942), .A2(n9870), .ZN(n9873) );
  CLKBUF_X1 U5583 ( .A(n9879), .Z(n9880) );
  CLKBUF_X1 U5584 ( .A(n6979), .Z(n6980) );
  AND2_X1 U5585 ( .A1(n9182), .A2(n8918), .ZN(n9433) );
  AND2_X1 U5586 ( .A1(n7620), .A2(n8918), .ZN(n9431) );
  INV_X1 U5587 ( .A(n4793), .ZN(n4792) );
  NAND2_X1 U5588 ( .A1(n5603), .A2(n5602), .ZN(n9383) );
  AND2_X1 U5589 ( .A1(n5170), .A2(n5169), .ZN(n9946) );
  NOR2_X1 U5590 ( .A1(n4783), .A2(n4458), .ZN(n4457) );
  INV_X1 U5591 ( .A(n4942), .ZN(n4458) );
  NAND2_X1 U5592 ( .A1(n4784), .A2(n4945), .ZN(n4783) );
  XNOR2_X1 U5593 ( .A(n5985), .B(SI_29_), .ZN(n7722) );
  INV_X1 U5594 ( .A(n5571), .ZN(n5568) );
  NAND2_X1 U5595 ( .A1(n4625), .A2(n4623), .ZN(n5512) );
  NAND2_X1 U5596 ( .A1(n4625), .A2(n5483), .ZN(n5491) );
  NOR2_X1 U5597 ( .A1(n4750), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4747) );
  INV_X1 U5598 ( .A(n5190), .ZN(n4749) );
  OAI21_X1 U5599 ( .B1(n5388), .B2(n4292), .A(n4610), .ZN(n5456) );
  NOR2_X1 U5600 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4558) );
  NAND2_X1 U5601 ( .A1(n4613), .A2(n5411), .ZN(n5438) );
  NAND2_X1 U5602 ( .A1(n5388), .A2(n4614), .ZN(n4613) );
  NAND2_X1 U5603 ( .A1(n5366), .A2(n5365), .ZN(n6653) );
  NAND2_X1 U5604 ( .A1(n4629), .A2(n4895), .ZN(n5228) );
  NAND2_X1 U5605 ( .A1(n5189), .A2(n4892), .ZN(n5246) );
  NOR2_X1 U5606 ( .A1(n4571), .A2(n5025), .ZN(n5138) );
  INV_X1 U5607 ( .A(n4947), .ZN(n4571) );
  AND2_X1 U5608 ( .A1(n7041), .A2(n7040), .ZN(n7044) );
  NAND2_X1 U5609 ( .A1(n4803), .A2(n4295), .ZN(n7984) );
  NAND2_X1 U5610 ( .A1(n4801), .A2(n4799), .ZN(n4803) );
  AND3_X1 U5611 ( .A1(n6356), .A2(n6355), .A3(n6354), .ZN(n8488) );
  INV_X1 U5612 ( .A(n8442), .ZN(n8261) );
  OAI21_X1 U5613 ( .B1(n8267), .B2(n7967), .A(n7966), .ZN(n8258) );
  AND4_X1 U5614 ( .A1(n6206), .A2(n6205), .A3(n6204), .A4(n6203), .ZN(n7154)
         );
  NAND2_X1 U5615 ( .A1(n6997), .A2(n6996), .ZN(n7013) );
  NOR2_X1 U5616 ( .A1(n7140), .A2(n4812), .ZN(n4811) );
  INV_X1 U5617 ( .A(n7136), .ZN(n4812) );
  NAND2_X1 U5618 ( .A1(n4829), .A2(n4830), .ZN(n8307) );
  AND4_X1 U5619 ( .A1(n6312), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(n7731)
         );
  OR2_X1 U5620 ( .A1(n6801), .A2(n6796), .ZN(n8299) );
  INV_X1 U5621 ( .A(n7003), .ZN(n8291) );
  NAND2_X1 U5622 ( .A1(n4602), .A2(n4601), .ZN(n8220) );
  NAND2_X1 U5623 ( .A1(n4303), .A2(n4286), .ZN(n4601) );
  INV_X1 U5624 ( .A(n7154), .ZN(n6453) );
  INV_X1 U5625 ( .A(n7025), .ZN(n8343) );
  NAND2_X1 U5626 ( .A1(n6437), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6137) );
  OR2_X1 U5627 ( .A1(n6340), .A2(n6140), .ZN(n6141) );
  OR2_X1 U5628 ( .A1(n6676), .A2(n6675), .ZN(n6678) );
  NAND2_X1 U5629 ( .A1(n4670), .A2(n6701), .ZN(n6744) );
  NOR2_X1 U5630 ( .A1(n6737), .A2(n4381), .ZN(n6699) );
  AND2_X1 U5631 ( .A1(n5907), .A2(n6752), .ZN(n4381) );
  NAND2_X1 U5632 ( .A1(n6699), .A2(n6698), .ZN(n6697) );
  NAND2_X1 U5633 ( .A1(n6697), .A2(n4380), .ZN(n6757) );
  NAND2_X1 U5634 ( .A1(n5908), .A2(n6718), .ZN(n4380) );
  NAND2_X1 U5635 ( .A1(n6757), .A2(n6756), .ZN(n6755) );
  NAND2_X1 U5636 ( .A1(n4581), .A2(n5873), .ZN(n6762) );
  INV_X1 U5637 ( .A(n4579), .ZN(n6760) );
  NAND2_X1 U5638 ( .A1(n4573), .A2(n5879), .ZN(n7925) );
  NOR2_X1 U5639 ( .A1(n7915), .A2(n7914), .ZN(n7913) );
  NOR2_X1 U5640 ( .A1(n7931), .A2(n5835), .ZN(n7915) );
  NAND2_X1 U5641 ( .A1(n5843), .A2(n4360), .ZN(n6959) );
  NOR2_X1 U5642 ( .A1(n6962), .A2(n5884), .ZN(n7885) );
  INV_X1 U5643 ( .A(n4370), .ZN(n7838) );
  INV_X1 U5644 ( .A(n4583), .ZN(n5889) );
  NOR2_X1 U5645 ( .A1(n5895), .A2(n8362), .ZN(n7790) );
  INV_X1 U5646 ( .A(n4663), .ZN(n7774) );
  XNOR2_X1 U5647 ( .A(n5948), .B(n5947), .ZN(n4385) );
  NAND2_X1 U5648 ( .A1(n8409), .A2(n8020), .ZN(n8396) );
  AOI211_X1 U5649 ( .C1(n8394), .C2(n8510), .A(n8393), .B(n8392), .ZN(n8536)
         );
  AND2_X1 U5650 ( .A1(n8390), .A2(n8389), .ZN(n8393) );
  AND2_X1 U5651 ( .A1(n4647), .A2(n6106), .ZN(n8414) );
  NAND2_X1 U5652 ( .A1(n7582), .A2(n6219), .ZN(n4647) );
  AOI21_X1 U5653 ( .B1(n8408), .B2(n8510), .A(n8407), .ZN(n8539) );
  OAI21_X1 U5654 ( .B1(n6472), .B2(n9712), .A(n8406), .ZN(n8407) );
  NAND2_X1 U5655 ( .A1(n8405), .A2(n8512), .ZN(n8406) );
  AND2_X1 U5656 ( .A1(n8431), .A2(n8430), .ZN(n8542) );
  INV_X1 U5657 ( .A(n8743), .ZN(n8426) );
  NAND2_X1 U5658 ( .A1(n4723), .A2(n4720), .ZN(n8452) );
  NAND2_X1 U5659 ( .A1(n8560), .A2(n8027), .ZN(n8465) );
  AND2_X1 U5660 ( .A1(n8509), .A2(n6349), .ZN(n8499) );
  NAND2_X1 U5661 ( .A1(n7613), .A2(n4687), .ZN(n8578) );
  AND2_X1 U5662 ( .A1(n8210), .A2(n8034), .ZN(n4687) );
  NAND2_X1 U5663 ( .A1(n7613), .A2(n8034), .ZN(n7681) );
  NAND2_X1 U5664 ( .A1(n6328), .A2(n6327), .ZN(n8312) );
  OAI21_X1 U5665 ( .B1(n7425), .B2(n4692), .A(n4690), .ZN(n7509) );
  NAND2_X1 U5666 ( .A1(n7427), .A2(n8124), .ZN(n7510) );
  OAI21_X1 U5667 ( .B1(n7250), .B2(n4682), .A(n4680), .ZN(n9700) );
  NAND2_X1 U5668 ( .A1(n7249), .A2(n8109), .ZN(n9701) );
  NAND2_X1 U5669 ( .A1(n6264), .A2(n6263), .ZN(n7315) );
  OAI21_X1 U5670 ( .B1(n7172), .B2(n6253), .A(n4717), .ZN(n7344) );
  NAND2_X1 U5671 ( .A1(n7438), .A2(n8091), .ZN(n7346) );
  NAND2_X1 U5672 ( .A1(n4728), .A2(n6233), .ZN(n7437) );
  NAND2_X1 U5673 ( .A1(n6221), .A2(n6220), .ZN(n7166) );
  AOI22_X1 U5674 ( .A1(n6425), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6337), .B2(
        n7936), .ZN(n6221) );
  INV_X1 U5675 ( .A(n6454), .ZN(n7268) );
  OAI21_X1 U5676 ( .B1(n6452), .B2(n4676), .A(n4674), .ZN(n7118) );
  OR2_X1 U5677 ( .A1(n6926), .A2(n6925), .ZN(n9703) );
  OR2_X1 U5678 ( .A1(n6929), .A2(n9705), .ZN(n8523) );
  NAND2_X1 U5679 ( .A1(n8003), .A2(n8002), .ZN(n8586) );
  NAND2_X1 U5680 ( .A1(n7999), .A2(n7998), .ZN(n8591) );
  OR2_X1 U5681 ( .A1(n8550), .A2(n8549), .ZN(n8744) );
  INV_X1 U5682 ( .A(n7962), .ZN(n8752) );
  INV_X1 U5683 ( .A(n8029), .ZN(n8756) );
  AND2_X1 U5684 ( .A1(n6779), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6588) );
  OR2_X1 U5685 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  OR2_X1 U5686 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  NAND2_X1 U5687 ( .A1(n6434), .A2(n6433), .ZN(n8183) );
  NAND2_X1 U5688 ( .A1(n4816), .A2(n4820), .ZN(n6433) );
  NAND2_X1 U5689 ( .A1(n4297), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6434) );
  OR2_X1 U5690 ( .A1(n5856), .A2(n6109), .ZN(n4816) );
  INV_X1 U5691 ( .A(n7936), .ZN(n6554) );
  INV_X1 U5692 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6549) );
  OR2_X1 U5693 ( .A1(n5832), .A2(n5831), .ZN(n6548) );
  INV_X1 U5694 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6547) );
  INV_X1 U5695 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6542) );
  INV_X1 U5696 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6540) );
  XNOR2_X1 U5697 ( .A(n5815), .B(n5739), .ZN(n6538) );
  INV_X1 U5698 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6544) );
  INV_X1 U5699 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4857) );
  NAND2_X1 U5700 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5808) );
  NAND2_X1 U5701 ( .A1(n5155), .A2(n5154), .ZN(n7228) );
  NAND2_X1 U5702 ( .A1(n4521), .A2(n4520), .ZN(n4519) );
  INV_X1 U5703 ( .A(n5649), .ZN(n4520) );
  NAND2_X1 U5704 ( .A1(n4530), .A2(n4533), .ZN(n7636) );
  NAND2_X1 U5705 ( .A1(n4419), .A2(n4420), .ZN(n8793) );
  OR2_X1 U5706 ( .A1(n8820), .A2(n4422), .ZN(n4419) );
  NAND2_X1 U5707 ( .A1(n5724), .A2(n5723), .ZN(n5725) );
  NAND2_X1 U5708 ( .A1(n4540), .A2(n4543), .ZN(n7516) );
  OR2_X1 U5709 ( .A1(n7622), .A2(n5266), .ZN(n4540) );
  INV_X1 U5710 ( .A(n4387), .ZN(n8871) );
  INV_X1 U5711 ( .A(n7207), .ZN(n5148) );
  NAND2_X1 U5712 ( .A1(n4552), .A2(n5385), .ZN(n8828) );
  NAND2_X1 U5713 ( .A1(n8820), .A2(n8819), .ZN(n4552) );
  NAND2_X1 U5714 ( .A1(n4564), .A2(n4565), .ZN(n7086) );
  AND2_X1 U5715 ( .A1(n4564), .A2(n4562), .ZN(n7085) );
  OR2_X1 U5716 ( .A1(n6952), .A2(n6951), .ZN(n4564) );
  NAND2_X1 U5717 ( .A1(n4536), .A2(n4539), .ZN(n7603) );
  NAND2_X1 U5718 ( .A1(n7622), .A2(n4537), .ZN(n4536) );
  AOI21_X1 U5719 ( .B1(n5086), .B2(n5085), .A(n6853), .ZN(n6772) );
  NOR2_X1 U5720 ( .A1(n6772), .A2(n6771), .ZN(n6770) );
  OAI211_X1 U5721 ( .C1(n6567), .C2(n6534), .A(n5046), .B(n5045), .ZN(n6989)
         );
  OAI21_X1 U5722 ( .B1(n8820), .B2(n4551), .A(n4550), .ZN(n8861) );
  AND2_X1 U5723 ( .A1(n5720), .A2(n9501), .ZN(n8883) );
  OAI21_X1 U5724 ( .B1(n4387), .B2(n8873), .A(n8872), .ZN(n4386) );
  AND2_X1 U5725 ( .A1(n5657), .A2(n5605), .ZN(n9384) );
  OAI21_X1 U5726 ( .B1(n4442), .B2(n4435), .A(n4433), .ZN(n4432) );
  NAND2_X1 U5727 ( .A1(n4436), .A2(n6091), .ZN(n4435) );
  NOR2_X1 U5728 ( .A1(n4434), .A2(n9174), .ZN(n4433) );
  INV_X1 U5729 ( .A(n9112), .ZN(n4436) );
  NAND2_X1 U5730 ( .A1(n4440), .A2(n4309), .ZN(n4437) );
  NAND2_X1 U5731 ( .A1(n4442), .A2(n4441), .ZN(n4440) );
  NAND2_X1 U5732 ( .A1(n4439), .A2(n7084), .ZN(n4438) );
  INV_X1 U5733 ( .A(n9377), .ZN(n9189) );
  NAND2_X1 U5734 ( .A1(n5553), .A2(n5552), .ZN(n9432) );
  OR2_X1 U5735 ( .A1(n5429), .A2(n5428), .ZN(n9193) );
  OR2_X1 U5736 ( .A1(n5010), .A2(n5009), .ZN(n9194) );
  OR2_X1 U5737 ( .A1(n5401), .A2(n5400), .ZN(n9195) );
  INV_X1 U5738 ( .A(n7665), .ZN(n9196) );
  OR2_X1 U5739 ( .A1(n5331), .A2(n5330), .ZN(n9198) );
  OR2_X1 U5740 ( .A1(n5212), .A2(n5211), .ZN(n9204) );
  OR2_X1 U5741 ( .A1(n5164), .A2(n5163), .ZN(n9205) );
  OR2_X1 U5742 ( .A1(n5135), .A2(n5134), .ZN(n9207) );
  OR2_X1 U5743 ( .A1(n5093), .A2(n5070), .ZN(n5074) );
  OR2_X1 U5744 ( .A1(n4279), .A2(n5069), .ZN(n5075) );
  OR2_X1 U5745 ( .A1(n9269), .A2(n9268), .ZN(n9283) );
  NOR2_X1 U5746 ( .A1(n5990), .A2(n9909), .ZN(n9314) );
  NAND2_X1 U5747 ( .A1(n6101), .A2(n6100), .ZN(n9331) );
  AOI211_X1 U5748 ( .C1(n6105), .C2(n9349), .A(n9909), .B(n9319), .ZN(n9330)
         );
  NAND2_X1 U5749 ( .A1(n9430), .A2(n9059), .ZN(n9407) );
  NAND2_X1 U5750 ( .A1(n5544), .A2(n5543), .ZN(n9416) );
  INV_X1 U5751 ( .A(n9563), .ZN(n9426) );
  OAI21_X1 U5752 ( .B1(n9477), .B2(n4497), .A(n4495), .ZN(n9420) );
  NAND2_X1 U5753 ( .A1(n4500), .A2(n4501), .ZN(n9439) );
  NAND2_X1 U5754 ( .A1(n9477), .A2(n4502), .ZN(n4500) );
  OAI21_X1 U5755 ( .B1(n9477), .B2(n4282), .A(n6045), .ZN(n9458) );
  NAND2_X1 U5756 ( .A1(n7645), .A2(n9137), .ZN(n7663) );
  NAND2_X1 U5757 ( .A1(n5342), .A2(n5341), .ZN(n9011) );
  NAND2_X1 U5758 ( .A1(n6030), .A2(n6029), .ZN(n7416) );
  NAND2_X1 U5759 ( .A1(n7536), .A2(n8921), .ZN(n7535) );
  NAND2_X1 U5760 ( .A1(n6028), .A2(n6027), .ZN(n7536) );
  INV_X1 U5761 ( .A(n9927), .ZN(n6943) );
  AND2_X1 U5762 ( .A1(n4482), .A2(n4484), .ZN(n6936) );
  NAND2_X1 U5763 ( .A1(n9889), .A2(n6018), .ZN(n4482) );
  NOR2_X1 U5764 ( .A1(n6103), .A2(n6880), .ZN(n9994) );
  INV_X1 U5765 ( .A(n9994), .ZN(n9996) );
  INV_X1 U5766 ( .A(n9996), .ZN(n9998) );
  AOI21_X1 U5767 ( .B1(n9539), .B2(n9971), .A(n9538), .ZN(n9611) );
  AOI211_X1 U5768 ( .C1(n9549), .C2(n9971), .A(n9548), .B(n9547), .ZN(n9615)
         );
  NAND2_X1 U5769 ( .A1(n5274), .A2(n5273), .ZN(n7523) );
  INV_X1 U5770 ( .A(n9841), .ZN(n7546) );
  CLKBUF_X1 U5771 ( .A(n5995), .Z(n9728) );
  NAND2_X1 U5772 ( .A1(n5485), .A2(n4623), .ZN(n4616) );
  NAND2_X1 U5773 ( .A1(n4559), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4974) );
  NAND2_X1 U5774 ( .A1(n5390), .A2(n4964), .ZN(n4559) );
  INV_X1 U5775 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6545) );
  AND2_X1 U5776 ( .A1(n4725), .A2(n4293), .ZN(n5137) );
  INV_X1 U5777 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6535) );
  XNOR2_X1 U5778 ( .A(n5031), .B(n5030), .ZN(n6541) );
  INV_X1 U5779 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6532) );
  INV_X1 U5780 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6533) );
  XNOR2_X1 U5781 ( .A(n4359), .B(n8319), .ZN(n8329) );
  INV_X1 U5782 ( .A(n4651), .ZN(n8350) );
  AOI21_X1 U5783 ( .B1(n4659), .B2(n4658), .A(n4655), .ZN(n7766) );
  NAND2_X1 U5784 ( .A1(n4660), .A2(n7762), .ZN(n4659) );
  MUX2_X1 U5785 ( .A(n6522), .B(n6521), .S(n10121), .Z(n6523) );
  MUX2_X1 U5786 ( .A(n6506), .B(n6521), .S(n10094), .Z(n6507) );
  MUX2_X1 U5787 ( .A(n9310), .B(n9309), .S(n9308), .Z(n9312) );
  AOI211_X1 U5788 ( .C1(n9542), .C2(n9896), .A(n9371), .B(n9370), .ZN(n9372)
         );
  NAND2_X1 U5789 ( .A1(n4475), .A2(n6906), .ZN(n6913) );
  OAI21_X1 U5790 ( .B1(n6524), .B2(n9982), .A(n4774), .ZN(P1_U3519) );
  NOR2_X1 U5791 ( .A1(n4348), .A2(n4775), .ZN(n4774) );
  NOR2_X1 U5792 ( .A1(n9983), .A2(n6104), .ZN(n4775) );
  NAND2_X2 U5793 ( .A1(n5016), .A2(n5014), .ZN(n5047) );
  INV_X1 U5794 ( .A(n6211), .ZN(n6397) );
  INV_X1 U5795 ( .A(n5014), .ZN(n5666) );
  NAND2_X1 U5796 ( .A1(n4749), .A2(n4747), .ZN(n4977) );
  AND2_X1 U5797 ( .A1(n9484), .A2(n9192), .ZN(n4282) );
  AND2_X1 U5798 ( .A1(n7721), .A2(n7650), .ZN(n4283) );
  XNOR2_X1 U5799 ( .A(n4880), .B(SI_7_), .ZN(n5167) );
  AND2_X1 U5800 ( .A1(n9940), .A2(n9946), .ZN(n4284) );
  AND2_X1 U5801 ( .A1(n4283), .A2(n4461), .ZN(n4285) );
  INV_X1 U5802 ( .A(n8921), .ZN(n4507) );
  OR2_X1 U5803 ( .A1(n8586), .A2(n8373), .ZN(n4286) );
  OR2_X1 U5804 ( .A1(n8872), .A2(n8873), .ZN(n4287) );
  AND2_X1 U5805 ( .A1(n4332), .A2(n4711), .ZN(n4288) );
  INV_X1 U5806 ( .A(n9450), .ZN(n9628) );
  NAND2_X1 U5807 ( .A1(n5495), .A2(n5494), .ZN(n9450) );
  AND2_X1 U5808 ( .A1(n4651), .A2(n4654), .ZN(n4289) );
  OR2_X1 U5809 ( .A1(n5589), .A2(n8810), .ZN(n5590) );
  OR2_X1 U5810 ( .A1(n9416), .A2(n8784), .ZN(n9068) );
  AND2_X1 U5811 ( .A1(n7592), .A2(n7588), .ZN(n4290) );
  INV_X1 U5812 ( .A(n9354), .ZN(n4473) );
  NAND2_X1 U5813 ( .A1(n4577), .A2(n4582), .ZN(n4581) );
  INV_X1 U5814 ( .A(n7752), .ZN(n4592) );
  INV_X2 U5815 ( .A(n6536), .ZN(n6537) );
  AND2_X1 U5816 ( .A1(n9121), .A2(n8965), .ZN(n4291) );
  INV_X1 U5817 ( .A(n6170), .ZN(n6340) );
  AND2_X2 U5818 ( .A1(n6117), .A2(n7724), .ZN(n6170) );
  OR2_X1 U5819 ( .A1(n5437), .A2(n4612), .ZN(n4292) );
  INV_X2 U5820 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6109) );
  OR2_X1 U5821 ( .A1(n4969), .A2(n4785), .ZN(n4967) );
  OR2_X1 U5822 ( .A1(n4871), .A2(n5030), .ZN(n4293) );
  NOR2_X1 U5823 ( .A1(n7138), .A2(n8340), .ZN(n4294) );
  AND2_X1 U5824 ( .A1(n4806), .A2(n4807), .ZN(n4295) );
  OR2_X1 U5825 ( .A1(n7780), .A2(n5855), .ZN(n4296) );
  AND2_X1 U5826 ( .A1(n4819), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4297) );
  INV_X1 U5827 ( .A(n6769), .ZN(n4582) );
  OR2_X1 U5828 ( .A1(n9563), .A2(n9065), .ZN(n4298) );
  AND2_X1 U5829 ( .A1(n4295), .A2(n4802), .ZN(n4299) );
  AND2_X1 U5830 ( .A1(n7676), .A2(n6336), .ZN(n4300) );
  AND2_X1 U5831 ( .A1(n8874), .A2(n8895), .ZN(n4301) );
  AND2_X1 U5832 ( .A1(n9574), .A2(n9191), .ZN(n4302) );
  INV_X1 U5833 ( .A(n5730), .ZN(n4523) );
  AND4_X1 U5834 ( .A1(n8219), .A2(n8218), .A3(n8217), .A4(n8216), .ZN(n4303)
         );
  XNOR2_X1 U5835 ( .A(n6114), .B(n6113), .ZN(n6117) );
  AND2_X1 U5836 ( .A1(n7073), .A2(n9847), .ZN(n4304) );
  AND2_X1 U5837 ( .A1(n8858), .A2(n8859), .ZN(n4305) );
  NAND2_X1 U5838 ( .A1(n5421), .A2(n5420), .ZN(n9500) );
  NAND2_X1 U5839 ( .A1(n5984), .A2(n5983), .ZN(n9323) );
  NAND2_X1 U5840 ( .A1(n4950), .A2(n4949), .ZN(n5165) );
  AND2_X1 U5841 ( .A1(n7390), .A2(n8338), .ZN(n4306) );
  NOR2_X1 U5842 ( .A1(n8793), .A2(n8790), .ZN(n4307) );
  OR2_X1 U5843 ( .A1(n7843), .A2(n5849), .ZN(n4308) );
  AND2_X1 U5844 ( .A1(n9090), .A2(n9085), .ZN(n9366) );
  NAND2_X1 U5845 ( .A1(n5867), .A2(n4599), .ZN(n5814) );
  OR2_X1 U5846 ( .A1(n9543), .A2(n9377), .ZN(n9090) );
  INV_X1 U5847 ( .A(n9323), .ZN(n9610) );
  NOR2_X1 U5848 ( .A1(n9178), .A2(n4438), .ZN(n4309) );
  OR2_X1 U5849 ( .A1(n8014), .A2(n8183), .ZN(n4310) );
  AND2_X1 U5850 ( .A1(n8752), .A2(n8475), .ZN(n8186) );
  NAND2_X1 U5851 ( .A1(n9207), .A2(n9934), .ZN(n4311) );
  INV_X1 U5852 ( .A(n5385), .ZN(n4555) );
  AND2_X1 U5853 ( .A1(n5108), .A2(n5109), .ZN(n4312) );
  AND2_X1 U5854 ( .A1(n4616), .A2(n4620), .ZN(n4313) );
  OR2_X1 U5855 ( .A1(n6567), .A2(n9240), .ZN(n4314) );
  INV_X1 U5856 ( .A(n4654), .ZN(n4653) );
  NAND2_X1 U5857 ( .A1(n5854), .A2(n6667), .ZN(n4654) );
  AND2_X1 U5858 ( .A1(n4593), .A2(n4592), .ZN(n4315) );
  AND2_X1 U5859 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4316) );
  NAND2_X1 U5860 ( .A1(n5745), .A2(n5744), .ZN(n4317) );
  AND2_X1 U5861 ( .A1(n4723), .A2(n6388), .ZN(n4318) );
  INV_X1 U5862 ( .A(n4464), .ZN(n4463) );
  NAND2_X1 U5863 ( .A1(n4466), .A2(n4465), .ZN(n4464) );
  OR2_X1 U5864 ( .A1(n5767), .A2(n5774), .ZN(n4319) );
  INV_X1 U5865 ( .A(n6730), .ZN(n4580) );
  XNOR2_X1 U5866 ( .A(n6060), .B(n8950), .ZN(n9325) );
  AND2_X1 U5867 ( .A1(n7069), .A2(n9946), .ZN(n4320) );
  INV_X1 U5868 ( .A(n5590), .ZN(n5591) );
  AND2_X1 U5869 ( .A1(n8273), .A2(n8331), .ZN(n4321) );
  NOR2_X1 U5870 ( .A1(n8858), .A2(n8859), .ZN(n4322) );
  NOR2_X1 U5871 ( .A1(n8533), .A2(n6472), .ZN(n4323) );
  OR2_X1 U5872 ( .A1(n5190), .A2(n4750), .ZN(n4324) );
  NOR2_X1 U5873 ( .A1(n9450), .A2(n9434), .ZN(n4325) );
  NOR2_X1 U5874 ( .A1(n5309), .A2(n5308), .ZN(n4326) );
  INV_X1 U5875 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4973) );
  OR2_X1 U5876 ( .A1(n4851), .A2(n4841), .ZN(n4327) );
  AND2_X1 U5877 ( .A1(n6538), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4328) );
  INV_X1 U5878 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4941) );
  INV_X1 U5879 ( .A(n8966), .ZN(n4782) );
  AND2_X1 U5880 ( .A1(n4902), .A2(SI_12_), .ZN(n4329) );
  NAND2_X1 U5881 ( .A1(n9460), .A2(n6086), .ZN(n9442) );
  OR2_X1 U5882 ( .A1(n6314), .A2(n8208), .ZN(n4330) );
  OR2_X1 U5883 ( .A1(n4632), .A2(n4628), .ZN(n4331) );
  NAND2_X1 U5884 ( .A1(n7315), .A2(n8337), .ZN(n4332) );
  INV_X1 U5885 ( .A(n4691), .ZN(n4690) );
  OAI21_X1 U5886 ( .B1(n8121), .B2(n4692), .A(n8126), .ZN(n4691) );
  INV_X1 U5887 ( .A(n8124), .ZN(n4692) );
  OR2_X1 U5888 ( .A1(n7589), .A2(n7693), .ZN(n8124) );
  NAND2_X1 U5889 ( .A1(n5882), .A2(n6571), .ZN(n5883) );
  AND2_X1 U5890 ( .A1(n6548), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4333) );
  AND2_X1 U5891 ( .A1(n5289), .A2(n5288), .ZN(n4334) );
  OR2_X1 U5892 ( .A1(n8591), .A2(n8004), .ZN(n8217) );
  NAND2_X1 U5893 ( .A1(n5536), .A2(n8780), .ZN(n8809) );
  AND2_X1 U5894 ( .A1(n4495), .A2(n4298), .ZN(n4335) );
  AND2_X1 U5895 ( .A1(n8216), .A2(n8177), .ZN(n4336) );
  INV_X1 U5896 ( .A(n9953), .ZN(n7457) );
  AND2_X1 U5897 ( .A1(n5202), .A2(n5201), .ZN(n9953) );
  AND4_X1 U5898 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n8420)
         );
  AND2_X1 U5899 ( .A1(n6291), .A2(n6315), .ZN(n4337) );
  AND2_X1 U5900 ( .A1(n5800), .A2(n5802), .ZN(n4338) );
  AND2_X1 U5901 ( .A1(n4293), .A2(n5136), .ZN(n4339) );
  INV_X1 U5902 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5229) );
  NOR2_X1 U5903 ( .A1(n7662), .A2(n4742), .ZN(n4741) );
  AND2_X1 U5904 ( .A1(n8157), .A2(n8027), .ZN(n4340) );
  AND2_X1 U5905 ( .A1(n5151), .A2(n5150), .ZN(n4341) );
  AND2_X1 U5906 ( .A1(n4286), .A2(n8183), .ZN(n4342) );
  AND2_X1 U5907 ( .A1(n4941), .A2(n4748), .ZN(n4343) );
  NOR2_X1 U5908 ( .A1(n8172), .A2(n8171), .ZN(n4344) );
  NAND2_X1 U5909 ( .A1(n5878), .A2(n6554), .ZN(n5879) );
  OR2_X1 U5910 ( .A1(n4969), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4345) );
  OR2_X1 U5911 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4346) );
  INV_X1 U5912 ( .A(n4721), .ZN(n4720) );
  NAND2_X1 U5913 ( .A1(n4722), .A2(n6388), .ZN(n4721) );
  INV_X1 U5914 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4703) );
  INV_X1 U5915 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4823) );
  NAND2_X1 U5916 ( .A1(n5989), .A2(n5988), .ZN(n6105) );
  INV_X1 U5917 ( .A(n6105), .ZN(n4474) );
  AND2_X1 U5918 ( .A1(n8517), .A2(n8133), .ZN(n8210) );
  AND2_X1 U5919 ( .A1(n6559), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4347) );
  OAI21_X1 U5920 ( .B1(n7738), .B2(n9029), .A(n9027), .ZN(n9509) );
  NAND2_X1 U5921 ( .A1(n4686), .A2(n8145), .ZN(n8490) );
  INV_X1 U5922 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4701) );
  AND4_X1 U5923 ( .A1(n6324), .A2(n6323), .A3(n6322), .A4(n6321), .ZN(n8311)
         );
  NAND2_X1 U5924 ( .A1(n4936), .A2(n4937), .ZN(n5190) );
  OR2_X1 U5925 ( .A1(n8825), .A2(n7665), .ZN(n9141) );
  INV_X1 U5926 ( .A(n9141), .ZN(n4756) );
  NAND2_X1 U5927 ( .A1(n4824), .A2(n7588), .ZN(n7590) );
  INV_X1 U5928 ( .A(n4623), .ZN(n4622) );
  NOR2_X1 U5929 ( .A1(n5490), .A2(n4624), .ZN(n4623) );
  NOR2_X1 U5930 ( .A1(n4474), .A2(n9645), .ZN(n4348) );
  INV_X1 U5931 ( .A(n8438), .ZN(n8405) );
  AND4_X1 U5932 ( .A1(n6409), .A2(n6408), .A3(n6407), .A4(n6406), .ZN(n8438)
         );
  INV_X1 U5933 ( .A(n5047), .ZN(n5243) );
  AND2_X1 U5934 ( .A1(n8899), .A2(n9059), .ZN(n9427) );
  INV_X1 U5935 ( .A(n9427), .ZN(n4767) );
  NAND2_X1 U5936 ( .A1(n9518), .A2(n4463), .ZN(n4467) );
  INV_X1 U5937 ( .A(n8458), .ZN(n4722) );
  AND3_X1 U5938 ( .A1(n6347), .A2(n6346), .A3(n6345), .ZN(n8286) );
  INV_X1 U5939 ( .A(n9346), .ZN(n9900) );
  NAND2_X1 U5940 ( .A1(n9410), .A2(n8955), .ZN(n5695) );
  NAND2_X1 U5941 ( .A1(n5370), .A2(n5369), .ZN(n8825) );
  INV_X1 U5942 ( .A(n8825), .ZN(n4461) );
  AND2_X1 U5943 ( .A1(n4560), .A2(n4561), .ZN(n4349) );
  NAND2_X1 U5944 ( .A1(n5392), .A2(n5391), .ZN(n9594) );
  INV_X1 U5945 ( .A(n9594), .ZN(n4460) );
  NAND2_X1 U5946 ( .A1(n6452), .A2(n8067), .ZN(n7189) );
  NAND2_X1 U5947 ( .A1(n9128), .A2(n9125), .ZN(n7286) );
  NAND2_X1 U5948 ( .A1(n4709), .A2(n4716), .ZN(n9706) );
  NAND2_X1 U5949 ( .A1(n5460), .A2(n5459), .ZN(n9574) );
  INV_X1 U5950 ( .A(n9574), .ZN(n4465) );
  NAND2_X1 U5951 ( .A1(n7137), .A2(n7136), .ZN(n7139) );
  NAND2_X1 U5952 ( .A1(n7250), .A2(n8203), .ZN(n7249) );
  NOR2_X1 U5953 ( .A1(n7876), .A2(n5847), .ZN(n4350) );
  NOR2_X1 U5954 ( .A1(n7885), .A2(n7884), .ZN(n4351) );
  NOR2_X1 U5955 ( .A1(n5955), .A2(n4384), .ZN(n4352) );
  INV_X1 U5956 ( .A(n10014), .ZN(n4658) );
  AND4_X1 U5957 ( .A1(n5040), .A2(n5039), .A3(n5038), .A4(n5037), .ZN(n6011)
         );
  INV_X1 U5958 ( .A(n5873), .ZN(n5875) );
  NAND2_X1 U5959 ( .A1(n5874), .A2(n6769), .ZN(n5873) );
  XNOR2_X1 U5960 ( .A(n5862), .B(n4823), .ZN(n8221) );
  NAND2_X1 U5961 ( .A1(n5193), .A2(n5192), .ZN(n9959) );
  INV_X1 U5962 ( .A(n9959), .ZN(n4468) );
  AND2_X1 U5963 ( .A1(n4579), .A2(n5873), .ZN(n4353) );
  AND4_X1 U5964 ( .A1(n5242), .A2(n5241), .A3(n5240), .A4(n5239), .ZN(n9201)
         );
  INV_X1 U5965 ( .A(n9201), .ZN(n4510) );
  NOR2_X1 U5966 ( .A1(n6723), .A2(n6722), .ZN(n4354) );
  NAND2_X1 U5967 ( .A1(n5816), .A2(n6538), .ZN(n6701) );
  INV_X1 U5968 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4395) );
  INV_X1 U5969 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n4585) );
  INV_X1 U5970 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n4372) );
  AOI21_X1 U5971 ( .B1(n9341), .B2(n9882), .A(n9340), .ZN(n9537) );
  INV_X1 U5972 ( .A(n7780), .ZN(n4364) );
  XNOR2_X1 U5973 ( .A(n5896), .B(n7780), .ZN(n7769) );
  NOR2_X1 U5974 ( .A1(n7780), .A2(n5896), .ZN(n5897) );
  OAI211_X1 U5975 ( .C1(n8874), .C2(n4527), .A(n8895), .B(n4519), .ZN(n5738)
         );
  XNOR2_X1 U5976 ( .A(n5886), .B(n7881), .ZN(n7866) );
  INV_X1 U5977 ( .A(n5957), .ZN(n5958) );
  NOR2_X1 U5978 ( .A1(n7848), .A2(n7847), .ZN(n7846) );
  INV_X1 U5979 ( .A(n4383), .ZN(n4382) );
  NAND4_X1 U5980 ( .A1(n4356), .A2(n9066), .A3(n9411), .A4(n4355), .ZN(n9070)
         );
  OR2_X1 U5981 ( .A1(n9063), .A2(n9111), .ZN(n4356) );
  MUX2_X2 U5982 ( .A(n9103), .B(n9111), .S(n9323), .Z(n9109) );
  INV_X1 U5983 ( .A(n4357), .ZN(n9024) );
  AOI21_X1 U5984 ( .B1(n9008), .B2(n9007), .A(n4358), .ZN(n4357) );
  NAND3_X1 U5985 ( .A1(n9023), .A2(n9022), .A3(n9021), .ZN(n4358) );
  NAND2_X1 U5986 ( .A1(n4451), .A2(n8981), .ZN(n4450) );
  INV_X1 U5987 ( .A(n4453), .ZN(n4452) );
  INV_X1 U5988 ( .A(n4444), .ZN(n4443) );
  OAI21_X1 U5989 ( .B1(n4385), .B2(n8357), .A(n4382), .ZN(n5957) );
  OAI211_X1 U5990 ( .C1(n7769), .C2(n4591), .A(n4590), .B(n5898), .ZN(n5899)
         );
  OAI21_X1 U5991 ( .B1(n5956), .B2(n9999), .A(n4352), .ZN(n4383) );
  NAND2_X1 U5992 ( .A1(n4576), .A2(n4575), .ZN(n6729) );
  NOR2_X1 U5993 ( .A1(n7811), .A2(n7810), .ZN(n7809) );
  NOR2_X1 U5994 ( .A1(n5887), .A2(n7865), .ZN(n7848) );
  OAI21_X1 U5995 ( .B1(n5894), .B2(n6667), .A(n5893), .ZN(n8364) );
  NAND2_X1 U5996 ( .A1(n7134), .A2(n7133), .ZN(n7137) );
  NAND2_X1 U5997 ( .A1(n7311), .A2(n7310), .ZN(n7373) );
  NAND2_X1 U5998 ( .A1(n4829), .A2(n4827), .ZN(n8305) );
  NAND2_X1 U5999 ( .A1(n4825), .A2(n8280), .ZN(n8246) );
  NAND2_X1 U6000 ( .A1(n7941), .A2(n4831), .ZN(n4829) );
  NAND2_X1 U6001 ( .A1(n4835), .A2(n7031), .ZN(n7041) );
  OAI21_X4 U6002 ( .B1(n6806), .B2(n6807), .A(n6805), .ZN(n6813) );
  NAND2_X2 U6003 ( .A1(n6486), .A2(n6586), .ZN(n6806) );
  INV_X2 U6004 ( .A(n5805), .ZN(n5759) );
  NAND2_X1 U6005 ( .A1(n7690), .A2(n7689), .ZN(n7728) );
  NAND2_X1 U6006 ( .A1(n4824), .A2(n4290), .ZN(n7687) );
  NAND2_X1 U6007 ( .A1(n4826), .A2(n8279), .ZN(n4825) );
  OR2_X1 U6008 ( .A1(n5844), .A2(n6571), .ZN(n4360) );
  NAND2_X1 U6009 ( .A1(n5844), .A2(n6571), .ZN(n5843) );
  NAND2_X1 U6010 ( .A1(n6758), .A2(n4368), .ZN(n4367) );
  OAI21_X1 U6011 ( .B1(n6554), .B2(n4369), .A(n5834), .ZN(n7932) );
  OR2_X1 U6012 ( .A1(n5816), .A2(n4328), .ZN(n4373) );
  NAND2_X1 U6013 ( .A1(n4374), .A2(n4373), .ZN(n6704) );
  NAND3_X1 U6014 ( .A1(n4670), .A2(n6701), .A3(P2_REG1_REG_3__SCAN_IN), .ZN(
        n6742) );
  NAND2_X4 U6015 ( .A1(n4378), .A2(n4376), .ZN(n7583) );
  NAND2_X1 U6016 ( .A1(n4386), .A2(n4301), .ZN(n8882) );
  NAND2_X1 U6017 ( .A1(n4526), .A2(n5590), .ZN(n4387) );
  NAND3_X1 U6018 ( .A1(n4406), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4405) );
  NAND3_X1 U6019 ( .A1(n4409), .A2(n9313), .A3(n4408), .ZN(n4407) );
  NAND2_X1 U6020 ( .A1(n8820), .A2(n4417), .ZN(n4416) );
  NAND2_X1 U6021 ( .A1(n5121), .A2(n5120), .ZN(n4426) );
  NAND2_X1 U6022 ( .A1(n4424), .A2(n4423), .ZN(n5198) );
  NAND3_X1 U6023 ( .A1(n5121), .A2(n5120), .A3(n4879), .ZN(n4423) );
  OAI21_X2 U6024 ( .B1(n9109), .B2(n9108), .A(n9165), .ZN(n4444) );
  AOI21_X1 U6025 ( .B1(n9045), .B2(n4445), .A(n4446), .ZN(n4447) );
  NAND2_X1 U6026 ( .A1(n9045), .A2(n9046), .ZN(n9056) );
  NAND2_X1 U6027 ( .A1(n4447), .A2(n9441), .ZN(n9062) );
  INV_X1 U6028 ( .A(n9057), .ZN(n4448) );
  INV_X1 U6029 ( .A(n5062), .ZN(n4449) );
  AOI21_X2 U6030 ( .B1(n4455), .B2(n4843), .A(n9100), .ZN(n9103) );
  NAND2_X1 U6031 ( .A1(n6070), .A2(n8966), .ZN(n8973) );
  NAND2_X1 U6032 ( .A1(n4981), .A2(n4942), .ZN(n4969) );
  NAND2_X1 U6033 ( .A1(n4981), .A2(n4457), .ZN(n4994) );
  INV_X1 U6034 ( .A(n4467), .ZN(n9470) );
  NAND2_X1 U6035 ( .A1(n9381), .A2(n4470), .ZN(n9318) );
  NAND2_X1 U6036 ( .A1(n9381), .A2(n9363), .ZN(n9358) );
  INV_X1 U6037 ( .A(n4476), .ZN(n6903) );
  NAND2_X1 U6038 ( .A1(n4476), .A2(n6891), .ZN(n6986) );
  NAND2_X1 U6039 ( .A1(n6892), .A2(n4476), .ZN(n6008) );
  OAI22_X1 U6040 ( .A1(n6892), .A2(n5016), .B1(n4476), .B2(n5642), .ZN(n5083)
         );
  NOR2_X1 U6041 ( .A1(n9210), .A2(n4476), .ZN(n6064) );
  AOI21_X1 U6042 ( .B1(n9210), .B2(n4476), .A(n9118), .ZN(n9120) );
  OAI22_X1 U6043 ( .A1(n9910), .A2(n9909), .B1(n4476), .B2(n9967), .ZN(n9912)
         );
  OR2_X1 U6044 ( .A1(n9526), .A2(n4476), .ZN(n4475) );
  INV_X1 U6045 ( .A(n6977), .ZN(n4480) );
  NAND2_X1 U6046 ( .A1(n4477), .A2(n8965), .ZN(n4478) );
  NAND3_X1 U6047 ( .A1(n4484), .A2(n4479), .A3(n4478), .ZN(n4483) );
  OAI21_X1 U6048 ( .B1(n4481), .B2(n4480), .A(n6018), .ZN(n4479) );
  INV_X1 U6049 ( .A(n6978), .ZN(n4481) );
  NAND2_X1 U6050 ( .A1(n6943), .A2(n9208), .ZN(n9121) );
  NAND2_X1 U6051 ( .A1(n6978), .A2(n6977), .ZN(n9889) );
  NAND2_X1 U6052 ( .A1(n4483), .A2(n6019), .ZN(n9871) );
  NAND2_X1 U6053 ( .A1(n6030), .A2(n4486), .ZN(n4485) );
  NAND2_X1 U6054 ( .A1(n7072), .A2(n4304), .ZN(n4488) );
  NAND2_X1 U6055 ( .A1(n4488), .A2(n4489), .ZN(n7235) );
  NAND2_X1 U6056 ( .A1(n9477), .A2(n4335), .ZN(n4494) );
  NAND3_X1 U6057 ( .A1(n4495), .A2(n4497), .A3(n4298), .ZN(n4493) );
  NAND2_X1 U6058 ( .A1(n6056), .A2(n6055), .ZN(n4515) );
  NAND2_X1 U6059 ( .A1(n8809), .A2(n4524), .ZN(n4517) );
  INV_X1 U6060 ( .A(n4521), .ZN(n4527) );
  NAND2_X1 U6061 ( .A1(n8809), .A2(n5592), .ZN(n4526) );
  INV_X1 U6062 ( .A(n7622), .ZN(n4532) );
  OAI21_X1 U6063 ( .B1(n8793), .B2(n8790), .A(n8794), .ZN(n8800) );
  INV_X1 U6064 ( .A(n4850), .ZN(n4556) );
  NAND2_X1 U6065 ( .A1(n5390), .A2(n4558), .ZN(n4557) );
  NAND2_X1 U6066 ( .A1(n6952), .A2(n4562), .ZN(n4560) );
  NAND3_X1 U6067 ( .A1(n4560), .A2(n4561), .A3(n4341), .ZN(n5155) );
  NAND2_X1 U6068 ( .A1(n4950), .A2(n4569), .ZN(n5367) );
  INV_X1 U6069 ( .A(n5367), .ZN(n4962) );
  NAND3_X1 U6070 ( .A1(n4947), .A2(n5041), .A3(n4570), .ZN(n5118) );
  INV_X1 U6071 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4572) );
  NAND3_X1 U6072 ( .A1(n4573), .A2(n5879), .A3(P2_REG2_REG_7__SCAN_IN), .ZN(
        n4574) );
  INV_X1 U6073 ( .A(n4574), .ZN(n7923) );
  NAND4_X1 U6074 ( .A1(n4581), .A2(n5873), .A3(P2_REG2_REG_5__SCAN_IN), .A4(
        n4580), .ZN(n4575) );
  NAND2_X1 U6075 ( .A1(n4589), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4587) );
  NAND2_X1 U6076 ( .A1(n4587), .A2(n6706), .ZN(n4588) );
  NAND2_X1 U6077 ( .A1(n4588), .A2(n6705), .ZN(n6709) );
  NAND2_X1 U6078 ( .A1(n5897), .A2(n4592), .ZN(n4590) );
  INV_X1 U6079 ( .A(n4595), .ZN(n7768) );
  XNOR2_X2 U6080 ( .A(n4600), .B(n4599), .ZN(n6175) );
  NAND2_X2 U6081 ( .A1(n4988), .A2(n4987), .ZN(n5016) );
  NAND3_X1 U6082 ( .A1(n4606), .A2(n4604), .A3(n4342), .ZN(n4603) );
  NAND2_X1 U6083 ( .A1(n5388), .A2(n4610), .ZN(n4607) );
  NAND2_X1 U6084 ( .A1(n4607), .A2(n4608), .ZN(n5458) );
  OAI21_X1 U6085 ( .B1(n5485), .B2(n4619), .A(n4617), .ZN(n5538) );
  OAI21_X2 U6086 ( .B1(n4627), .B2(n4331), .A(n4630), .ZN(n5359) );
  NAND3_X1 U6087 ( .A1(n4645), .A2(n4643), .A3(n4641), .ZN(n8180) );
  NOR2_X1 U6088 ( .A1(n4642), .A2(n4344), .ZN(n4641) );
  NOR2_X1 U6089 ( .A1(n8179), .A2(n8018), .ZN(n4642) );
  NAND2_X1 U6090 ( .A1(n4644), .A2(n8176), .ZN(n4643) );
  OAI21_X1 U6091 ( .B1(n8178), .B2(n8533), .A(n8217), .ZN(n4644) );
  NAND2_X1 U6092 ( .A1(n4646), .A2(n8137), .ZN(n4645) );
  OAI21_X1 U6093 ( .B1(n8178), .B2(n8404), .A(n4336), .ZN(n4646) );
  NAND2_X1 U6094 ( .A1(n8414), .A2(n8391), .ZN(n8020) );
  XNOR2_X1 U6095 ( .A(n5853), .B(n8368), .ZN(n8352) );
  NAND2_X1 U6096 ( .A1(n4664), .A2(n4665), .ZN(n5844) );
  NAND2_X1 U6097 ( .A1(n7931), .A2(n4666), .ZN(n4664) );
  NAND2_X1 U6098 ( .A1(n6452), .A2(n4674), .ZN(n4673) );
  NAND2_X1 U6099 ( .A1(n7250), .A2(n4680), .ZN(n4679) );
  NAND2_X1 U6100 ( .A1(n8503), .A2(n8144), .ZN(n4686) );
  NAND2_X1 U6101 ( .A1(n4686), .A2(n4683), .ZN(n6461) );
  NAND2_X1 U6102 ( .A1(n8578), .A2(n8138), .ZN(n6460) );
  NAND2_X1 U6103 ( .A1(n8411), .A2(n4695), .ZN(n4693) );
  NAND2_X1 U6104 ( .A1(n4693), .A2(n4694), .ZN(n7995) );
  NAND2_X1 U6105 ( .A1(n4698), .A2(n4699), .ZN(n6457) );
  NAND2_X1 U6106 ( .A1(n7440), .A2(n8091), .ZN(n4698) );
  NAND2_X1 U6107 ( .A1(n8560), .A2(n4340), .ZN(n6462) );
  NAND3_X1 U6108 ( .A1(n5771), .A2(n4703), .A3(n5763), .ZN(n5774) );
  AND3_X1 U6109 ( .A1(n5759), .A2(n5775), .A3(n4705), .ZN(n6110) );
  NAND2_X1 U6110 ( .A1(n5759), .A2(n5758), .ZN(n5776) );
  NAND3_X1 U6111 ( .A1(n5759), .A2(n5775), .A3(n4704), .ZN(n6107) );
  NAND2_X1 U6112 ( .A1(n7172), .A2(n4714), .ZN(n4710) );
  OR2_X1 U6113 ( .A1(n7336), .A2(n8339), .ZN(n4717) );
  OAI21_X1 U6114 ( .B1(n8462), .B2(n4721), .A(n4718), .ZN(n8437) );
  NAND2_X1 U6115 ( .A1(n4724), .A2(n4875), .ZN(n5121) );
  NAND2_X1 U6116 ( .A1(n4339), .A2(n4725), .ZN(n4724) );
  NAND2_X1 U6117 ( .A1(n5029), .A2(n4872), .ZN(n4725) );
  NAND2_X1 U6118 ( .A1(n4728), .A2(n4726), .ZN(n6244) );
  AOI21_X1 U6119 ( .B1(n6292), .B2(n4337), .A(n4729), .ZN(n7611) );
  NAND2_X1 U6120 ( .A1(n8509), .A2(n4732), .ZN(n8497) );
  NAND3_X1 U6121 ( .A1(n7271), .A2(n6223), .A3(n8078), .ZN(n4733) );
  NAND2_X1 U6122 ( .A1(n6084), .A2(n4736), .ZN(n4735) );
  NAND2_X1 U6123 ( .A1(n7643), .A2(n4741), .ZN(n4738) );
  NAND2_X1 U6124 ( .A1(n4738), .A2(n4739), .ZN(n7701) );
  AND4_X2 U6125 ( .A1(n4937), .A2(n4745), .A3(n4744), .A4(n4936), .ZN(n4981)
         );
  NAND3_X1 U6126 ( .A1(n4940), .A2(n4746), .A3(n4939), .ZN(n4750) );
  NAND2_X1 U6127 ( .A1(n6078), .A2(n4754), .ZN(n4753) );
  NAND2_X1 U6128 ( .A1(n9880), .A2(n4763), .ZN(n4758) );
  NAND2_X1 U6129 ( .A1(n4759), .A2(n6068), .ZN(n8964) );
  OR2_X1 U6130 ( .A1(n9879), .A2(n9117), .ZN(n4759) );
  OAI21_X1 U6131 ( .B1(n6087), .B2(n4768), .A(n4765), .ZN(n4770) );
  INV_X1 U6132 ( .A(n4770), .ZN(n9392) );
  NAND2_X1 U6133 ( .A1(n6101), .A2(n4772), .ZN(n4771) );
  AOI21_X1 U6134 ( .B1(n9325), .B2(n9971), .A(n4771), .ZN(n6524) );
  AOI21_X1 U6135 ( .B1(n9125), .B2(n4776), .A(n4778), .ZN(n4777) );
  AOI21_X1 U6136 ( .B1(n6070), .B2(n4779), .A(n4777), .ZN(n7542) );
  NAND3_X1 U6137 ( .A1(n4943), .A2(n4788), .A3(n4787), .ZN(n4786) );
  OAI21_X1 U6138 ( .B1(n9364), .B2(n4792), .A(n4789), .ZN(n6090) );
  NAND2_X1 U6139 ( .A1(n9364), .A2(n6089), .ZN(n4794) );
  NAND2_X1 U6140 ( .A1(n8267), .A2(n4798), .ZN(n4797) );
  NAND2_X1 U6141 ( .A1(n8267), .A2(n7966), .ZN(n4801) );
  NAND2_X1 U6142 ( .A1(n7137), .A2(n4811), .ZN(n7305) );
  NAND2_X1 U6143 ( .A1(n5856), .A2(n4820), .ZN(n4818) );
  NAND2_X1 U6144 ( .A1(n5856), .A2(n4822), .ZN(n4819) );
  NAND2_X1 U6145 ( .A1(n5856), .A2(n5746), .ZN(n5859) );
  NAND2_X1 U6146 ( .A1(n7586), .A2(n7585), .ZN(n4824) );
  NAND2_X1 U6147 ( .A1(n7951), .A2(n8286), .ZN(n4826) );
  INV_X1 U6148 ( .A(n7029), .ZN(n4835) );
  NAND2_X1 U6149 ( .A1(n5823), .A2(n5743), .ZN(n5805) );
  NAND2_X1 U6150 ( .A1(n5823), .A2(n4837), .ZN(n5799) );
  INV_X1 U6151 ( .A(n6175), .ZN(n10012) );
  NAND2_X1 U6152 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  NAND2_X1 U6153 ( .A1(n9089), .A2(n9088), .ZN(n9094) );
  NAND2_X1 U6154 ( .A1(n5783), .A2(n5782), .ZN(n5784) );
  OAI21_X1 U6155 ( .B1(n8455), .B2(n8261), .A(n8435), .ZN(n8418) );
  INV_X1 U6156 ( .A(n5064), .ZN(n5199) );
  OR2_X1 U6157 ( .A1(n5093), .A2(n5050), .ZN(n5057) );
  NAND2_X1 U6158 ( .A1(n7948), .A2(n7947), .ZN(n7951) );
  INV_X2 U6159 ( .A(n6155), .ZN(n6337) );
  AND2_X4 U6160 ( .A1(n6118), .A2(n7724), .ZN(n6159) );
  INV_X1 U6161 ( .A(n5001), .ZN(n5052) );
  INV_X1 U6162 ( .A(n7982), .ZN(n7986) );
  INV_X2 U6163 ( .A(n8001), .ZN(n6425) );
  AOI21_X1 U6164 ( .B1(n7984), .B2(n7983), .A(n8328), .ZN(n7985) );
  OR2_X1 U6165 ( .A1(n5865), .A2(n10014), .ZN(n4839) );
  AND2_X1 U6166 ( .A1(n6888), .A2(n9501), .ZN(n9523) );
  AND2_X1 U6167 ( .A1(n6480), .A2(n10072), .ZN(n4840) );
  INV_X1 U6168 ( .A(n6472), .ZN(n8404) );
  AND2_X1 U6169 ( .A1(n5479), .A2(n5478), .ZN(n4841) );
  OR2_X1 U6170 ( .A1(n8381), .A2(n8768), .ZN(n4842) );
  AND2_X1 U6171 ( .A1(n9096), .A2(n4854), .ZN(n4843) );
  NAND2_X1 U6172 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .ZN(n4844) );
  AND2_X1 U6173 ( .A1(n8533), .A2(n8404), .ZN(n4845) );
  AND2_X1 U6174 ( .A1(n5699), .A2(n5698), .ZN(n4846) );
  OR2_X1 U6175 ( .A1(n8381), .A2(n8576), .ZN(n4847) );
  OR2_X1 U6176 ( .A1(n4474), .A2(n9602), .ZN(n4848) );
  OR2_X1 U6177 ( .A1(n8376), .A2(n8330), .ZN(n4849) );
  AND2_X1 U6178 ( .A1(n5407), .A2(n5406), .ZN(n4850) );
  NOR2_X1 U6179 ( .A1(n5476), .A2(n8801), .ZN(n4851) );
  NOR2_X1 U6180 ( .A1(n5757), .A2(n5756), .ZN(n5758) );
  INV_X1 U6181 ( .A(n9602), .ZN(n6004) );
  INV_X1 U6182 ( .A(n8369), .ZN(n5954) );
  AND2_X1 U6183 ( .A1(n8176), .A2(n8389), .ZN(n8513) );
  INV_X1 U6184 ( .A(n8513), .ZN(n9712) );
  NAND2_X1 U6185 ( .A1(n7154), .A2(n6454), .ZN(n4852) );
  NOR2_X1 U6186 ( .A1(n5964), .A2(n5963), .ZN(n4853) );
  OR2_X1 U6187 ( .A1(n9095), .A2(n9104), .ZN(n4854) );
  NAND2_X1 U6188 ( .A1(n7271), .A2(n8078), .ZN(n4855) );
  OR2_X1 U6189 ( .A1(n5357), .A2(n5356), .ZN(n4856) );
  INV_X1 U6190 ( .A(n5337), .ZN(n4919) );
  XNOR2_X1 U6191 ( .A(n6067), .B(n9921), .ZN(n9890) );
  AOI21_X1 U6192 ( .B1(n8175), .B2(n8174), .A(n8173), .ZN(n8178) );
  NAND2_X1 U6193 ( .A1(n7156), .A2(n6228), .ZN(n6230) );
  AND2_X1 U6194 ( .A1(n8998), .A2(n8995), .ZN(n9131) );
  NAND2_X1 U6195 ( .A1(n8399), .A2(n6472), .ZN(n6423) );
  INV_X1 U6196 ( .A(n8205), .ZN(n6291) );
  INV_X1 U6197 ( .A(n8519), .ZN(n6348) );
  INV_X1 U6198 ( .A(n8895), .ZN(n5697) );
  INV_X1 U6199 ( .A(n5498), .ZN(n5496) );
  OR2_X1 U6200 ( .A1(n5522), .A2(n8783), .ZN(n5547) );
  NAND2_X1 U6201 ( .A1(n5359), .A2(n4906), .ZN(n4927) );
  INV_X1 U6202 ( .A(n5290), .ZN(n5310) );
  INV_X1 U6203 ( .A(n5167), .ZN(n4879) );
  INV_X1 U6204 ( .A(n7591), .ZN(n7592) );
  INV_X1 U6205 ( .A(n7014), .ZN(n6998) );
  INV_X1 U6206 ( .A(n7030), .ZN(n7031) );
  NOR2_X1 U6207 ( .A1(n5954), .A2(n8221), .ZN(n5955) );
  INV_X1 U6208 ( .A(n8210), .ZN(n6335) );
  INV_X1 U6209 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6184) );
  OR2_X1 U6210 ( .A1(n8137), .A2(n6475), .ZN(n6483) );
  NAND2_X1 U6211 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  NOR2_X1 U6212 ( .A1(n5701), .A2(n5697), .ZN(n5698) );
  OR2_X1 U6213 ( .A1(n5576), .A2(n5575), .ZN(n5604) );
  OR2_X1 U6214 ( .A1(n9675), .A2(n6617), .ZN(n9688) );
  INV_X1 U6215 ( .A(n9342), .ZN(n9335) );
  NAND2_X1 U6216 ( .A1(n5545), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U6217 ( .A1(n6567), .A2(n6537), .ZN(n5096) );
  INV_X1 U6218 ( .A(n9646), .ZN(n5999) );
  OR2_X1 U6219 ( .A1(n5969), .A2(n5968), .ZN(n5970) );
  OR2_X1 U6220 ( .A1(n6247), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U6221 ( .A1(n6361), .A2(n6360), .ZN(n6370) );
  AND2_X1 U6222 ( .A1(n6306), .A2(n7691), .ZN(n6319) );
  OR2_X1 U6223 ( .A1(n6370), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6380) );
  INV_X1 U6224 ( .A(n8297), .ZN(n8322) );
  AOI21_X1 U6225 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n6662), .A(n7819), .ZN(
        n5853) );
  NAND2_X1 U6226 ( .A1(n8017), .A2(n8177), .ZN(n6473) );
  AND2_X1 U6227 ( .A1(n8160), .A2(n8161), .ZN(n8458) );
  AND2_X1 U6228 ( .A1(n8109), .A2(n8108), .ZN(n8203) );
  NAND2_X1 U6229 ( .A1(n6455), .A2(n8194), .ZN(n7272) );
  INV_X1 U6230 ( .A(n8179), .ZN(n8381) );
  INV_X1 U6231 ( .A(n8337), .ZN(n9709) );
  INV_X1 U6232 ( .A(n8510), .ZN(n10024) );
  NAND2_X1 U6233 ( .A1(n8773), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6114) );
  AND2_X1 U6234 ( .A1(n5153), .A2(n5152), .ZN(n5154) );
  OR2_X1 U6235 ( .A1(n5384), .A2(n5383), .ZN(n5385) );
  AND2_X1 U6236 ( .A1(n5196), .A2(n5195), .ZN(n7553) );
  OR2_X1 U6237 ( .A1(n5710), .A2(n5694), .ZN(n5716) );
  OR2_X1 U6238 ( .A1(n9348), .A2(n5704), .ZN(n5663) );
  INV_X1 U6239 ( .A(n5994), .ZN(n5500) );
  AND2_X1 U6240 ( .A1(n9674), .A2(n9673), .ZN(n9675) );
  INV_X1 U6241 ( .A(n9543), .ZN(n9363) );
  INV_X1 U6242 ( .A(n9065), .ZN(n9447) );
  AND2_X1 U6243 ( .A1(n9152), .A2(n9156), .ZN(n9495) );
  NAND2_X1 U6244 ( .A1(n7299), .A2(n5986), .ZN(n5544) );
  NAND2_X1 U6245 ( .A1(n4991), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4992) );
  XNOR2_X1 U6246 ( .A(n4860), .B(SI_1_), .ZN(n5063) );
  AND4_X1 U6247 ( .A1(n6422), .A2(n6421), .A3(n6420), .A4(n6419), .ZN(n6472)
         );
  INV_X1 U6248 ( .A(n6473), .ZN(n8219) );
  AND2_X1 U6249 ( .A1(n9716), .A2(n9714), .ZN(n8525) );
  AND2_X1 U6250 ( .A1(n6519), .A2(n6518), .ZN(n6920) );
  AND2_X1 U6251 ( .A1(n8445), .A2(n7081), .ZN(n10072) );
  OAI21_X1 U6252 ( .B1(n9363), .B2(n8883), .A(n5735), .ZN(n5736) );
  OAI21_X1 U6253 ( .B1(n6857), .B2(n5016), .A(n5079), .ZN(n6821) );
  INV_X1 U6254 ( .A(n8883), .ZN(n8887) );
  OR2_X1 U6255 ( .A1(n9414), .A2(n5704), .ZN(n5553) );
  AND4_X1 U6256 ( .A1(n5378), .A2(n5377), .A3(n5376), .A4(n5375), .ZN(n7665)
         );
  AND4_X1 U6257 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n7539)
         );
  AND2_X1 U6258 ( .A1(n9510), .A2(n9147), .ZN(n8943) );
  INV_X1 U6259 ( .A(n9934), .ZN(n9870) );
  INV_X1 U6260 ( .A(n9526), .ZN(n9884) );
  INV_X1 U6261 ( .A(n9484), .ZN(n6085) );
  NAND2_X1 U6262 ( .A1(n9851), .A2(n9977), .ZN(n9971) );
  AND2_X1 U6263 ( .A1(n4986), .A2(n5691), .ZN(n9184) );
  XNOR2_X1 U6264 ( .A(n4876), .B(SI_6_), .ZN(n5120) );
  NAND2_X1 U6265 ( .A1(n7986), .A2(n7985), .ZN(n7990) );
  OR3_X1 U6266 ( .A1(n6793), .A2(n6792), .A3(n6925), .ZN(n8328) );
  AND4_X1 U6267 ( .A1(n8010), .A2(n6431), .A3(n6430), .A4(n6429), .ZN(n8015)
         );
  OR2_X1 U6268 ( .A1(P2_U3150), .A2(n5949), .ZN(n10021) );
  OR2_X1 U6269 ( .A1(n6642), .A2(n8224), .ZN(n10014) );
  OR2_X1 U6270 ( .A1(n6642), .A2(n7583), .ZN(n9999) );
  XNOR2_X1 U6271 ( .A(n7995), .B(n8219), .ZN(n8387) );
  INV_X1 U6272 ( .A(n10121), .ZN(n10119) );
  AND2_X1 U6273 ( .A1(n6505), .A2(n6504), .ZN(n10092) );
  INV_X1 U6274 ( .A(n6569), .ZN(n6580) );
  NAND2_X1 U6275 ( .A1(n5700), .A2(n4846), .ZN(n5728) );
  AND2_X1 U6276 ( .A1(n5709), .A2(n5708), .ZN(n9339) );
  OAI211_X1 U6277 ( .C1(n4278), .C2(n9626), .A(n5503), .B(n5502), .ZN(n9434)
         );
  OR2_X1 U6278 ( .A1(n5351), .A2(n5350), .ZN(n9197) );
  OR2_X1 U6279 ( .A1(n9900), .A2(n6938), .ZN(n9530) );
  NAND2_X1 U6280 ( .A1(n9105), .A2(n6004), .ZN(n6005) );
  INV_X1 U6281 ( .A(n9383), .ZN(n9618) );
  OR2_X1 U6282 ( .A1(n6103), .A2(n6102), .ZN(n9982) );
  INV_X1 U6283 ( .A(n9906), .ZN(n9907) );
  INV_X1 U6284 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n8651) );
  INV_X1 U6285 ( .A(n8348), .ZN(P2_U3893) );
  AND2_X1 U6286 ( .A1(n6536), .A2(SI_0_), .ZN(n5077) );
  NAND2_X1 U6287 ( .A1(n5077), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4859) );
  AND2_X1 U6288 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4858) );
  NAND2_X1 U6289 ( .A1(n6537), .A2(n4858), .ZN(n6166) );
  NAND2_X1 U6290 ( .A1(n4859), .A2(n6166), .ZN(n5062) );
  NAND2_X1 U6291 ( .A1(n4860), .A2(SI_1_), .ZN(n4861) );
  MUX2_X1 U6292 ( .A(n6544), .B(n6533), .S(n6536), .Z(n4862) );
  INV_X1 U6293 ( .A(n4862), .ZN(n4863) );
  NAND2_X1 U6294 ( .A1(n4863), .A2(SI_2_), .ZN(n4864) );
  NAND2_X1 U6295 ( .A1(n4865), .A2(n4864), .ZN(n5095) );
  MUX2_X1 U6296 ( .A(n6540), .B(n6532), .S(n6536), .Z(n4866) );
  NAND2_X1 U6297 ( .A1(n5095), .A2(n5094), .ZN(n5029) );
  INV_X1 U6298 ( .A(n4866), .ZN(n4867) );
  NAND2_X1 U6299 ( .A1(n4867), .A2(SI_3_), .ZN(n5028) );
  MUX2_X1 U6300 ( .A(n6542), .B(n6535), .S(n6536), .Z(n4870) );
  INV_X1 U6301 ( .A(n4870), .ZN(n4868) );
  NAND2_X1 U6302 ( .A1(n4868), .A2(SI_4_), .ZN(n4869) );
  AND2_X1 U6303 ( .A1(n5028), .A2(n4869), .ZN(n4872) );
  INV_X1 U6304 ( .A(n4869), .ZN(n4871) );
  MUX2_X1 U6305 ( .A(n6547), .B(n6545), .S(n6536), .Z(n4873) );
  INV_X1 U6306 ( .A(n4873), .ZN(n4874) );
  NAND2_X1 U6307 ( .A1(n4874), .A2(SI_5_), .ZN(n4875) );
  INV_X1 U6308 ( .A(n4876), .ZN(n4877) );
  NAND2_X1 U6309 ( .A1(n4877), .A2(SI_6_), .ZN(n4878) );
  MUX2_X1 U6310 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6536), .Z(n4880) );
  NAND2_X1 U6311 ( .A1(n4880), .A2(SI_7_), .ZN(n4881) );
  INV_X1 U6312 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6561) );
  INV_X1 U6313 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n4882) );
  MUX2_X1 U6314 ( .A(n6561), .B(n4882), .S(n6536), .Z(n4884) );
  INV_X1 U6315 ( .A(SI_8_), .ZN(n4883) );
  INV_X1 U6316 ( .A(n4884), .ZN(n4885) );
  NAND2_X1 U6317 ( .A1(n4885), .A2(SI_8_), .ZN(n4886) );
  INV_X1 U6318 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6572) );
  INV_X1 U6319 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6574) );
  MUX2_X1 U6320 ( .A(n6572), .B(n6574), .S(n6536), .Z(n4889) );
  INV_X1 U6321 ( .A(SI_9_), .ZN(n4888) );
  INV_X1 U6322 ( .A(n4889), .ZN(n4890) );
  NAND2_X1 U6323 ( .A1(n4890), .A2(SI_9_), .ZN(n4891) );
  INV_X1 U6324 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6577) );
  INV_X1 U6325 ( .A(n4893), .ZN(n4894) );
  NAND2_X1 U6326 ( .A1(n4894), .A2(SI_10_), .ZN(n4895) );
  INV_X1 U6327 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n8631) );
  INV_X1 U6328 ( .A(SI_11_), .ZN(n8682) );
  INV_X1 U6329 ( .A(n4897), .ZN(n4898) );
  NAND2_X1 U6330 ( .A1(n4898), .A2(SI_11_), .ZN(n4899) );
  NAND2_X1 U6331 ( .A1(n4900), .A2(n4899), .ZN(n5227) );
  INV_X1 U6332 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6631) );
  INV_X1 U6333 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6634) );
  XNOR2_X1 U6334 ( .A(n4901), .B(SI_12_), .ZN(n5268) );
  INV_X1 U6335 ( .A(n4901), .ZN(n4902) );
  XNOR2_X1 U6336 ( .A(n4911), .B(SI_13_), .ZN(n5290) );
  INV_X1 U6337 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6664) );
  INV_X1 U6338 ( .A(SI_14_), .ZN(n4904) );
  NAND2_X1 U6339 ( .A1(n4912), .A2(n4904), .ZN(n4915) );
  INV_X1 U6340 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6666) );
  INV_X1 U6341 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6670) );
  INV_X1 U6342 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6657) );
  INV_X1 U6343 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6654) );
  INV_X1 U6344 ( .A(SI_16_), .ZN(n4905) );
  NAND2_X1 U6345 ( .A1(n4907), .A2(n4905), .ZN(n4910) );
  INV_X1 U6346 ( .A(n4910), .ZN(n4925) );
  INV_X1 U6347 ( .A(n4907), .ZN(n4908) );
  NAND2_X1 U6348 ( .A1(n4908), .A2(SI_16_), .ZN(n4909) );
  NAND2_X1 U6349 ( .A1(n4910), .A2(n4909), .ZN(n5363) );
  INV_X1 U6350 ( .A(n5363), .ZN(n4924) );
  INV_X1 U6351 ( .A(n4915), .ZN(n4918) );
  NAND2_X1 U6352 ( .A1(n4911), .A2(SI_13_), .ZN(n5311) );
  INV_X1 U6353 ( .A(n4912), .ZN(n4913) );
  NAND2_X1 U6354 ( .A1(n4913), .A2(SI_14_), .ZN(n4914) );
  NAND2_X1 U6355 ( .A1(n4915), .A2(n4914), .ZN(n5313) );
  INV_X1 U6356 ( .A(n5313), .ZN(n4916) );
  INV_X1 U6357 ( .A(n4920), .ZN(n4921) );
  NAND2_X1 U6358 ( .A1(n4921), .A2(SI_15_), .ZN(n4922) );
  NAND2_X1 U6359 ( .A1(n4927), .A2(n4926), .ZN(n5387) );
  INV_X1 U6360 ( .A(n5387), .ZN(n4933) );
  INV_X1 U6361 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6652) );
  INV_X1 U6362 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6650) );
  INV_X1 U6363 ( .A(SI_17_), .ZN(n4928) );
  NAND2_X1 U6364 ( .A1(n4929), .A2(n4928), .ZN(n4934) );
  INV_X1 U6365 ( .A(n4929), .ZN(n4930) );
  NAND2_X1 U6366 ( .A1(n4930), .A2(SI_17_), .ZN(n4931) );
  NAND2_X1 U6367 ( .A1(n4934), .A2(n4931), .ZN(n5386) );
  INV_X1 U6368 ( .A(n5386), .ZN(n4932) );
  NAND2_X1 U6369 ( .A1(n4933), .A2(n4932), .ZN(n5388) );
  INV_X1 U6370 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6693) );
  XNOR2_X1 U6371 ( .A(n5409), .B(SI_18_), .ZN(n5408) );
  XNOR2_X1 U6372 ( .A(n5413), .B(n5408), .ZN(n6672) );
  NOR2_X1 U6373 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n4942) );
  INV_X1 U6374 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4944) );
  XNOR2_X1 U6375 ( .A(n4990), .B(n4944), .ZN(n5703) );
  NAND2_X1 U6376 ( .A1(n6672), .A2(n5986), .ZN(n4966) );
  INV_X1 U6377 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4948) );
  INV_X1 U6378 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4951) );
  NAND2_X1 U6379 ( .A1(n5230), .A2(n4951), .ZN(n5269) );
  INV_X1 U6380 ( .A(n5269), .ZN(n4953) );
  INV_X1 U6381 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n4952) );
  NAND3_X1 U6382 ( .A1(n4954), .A2(n4953), .A3(n4952), .ZN(n4959) );
  INV_X1 U6383 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5272) );
  NAND4_X1 U6384 ( .A1(n4957), .A2(n4956), .A3(n5272), .A4(n4955), .ZN(n4958)
         );
  NOR2_X1 U6385 ( .A1(n4959), .A2(n4958), .ZN(n4960) );
  INV_X1 U6386 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4961) );
  NAND2_X1 U6387 ( .A1(n4962), .A2(n4961), .ZN(n4963) );
  XNOR2_X1 U6388 ( .A(n4974), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9834) );
  AOI22_X1 U6389 ( .A1(n5419), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5418), .B2(
        n9834), .ZN(n4965) );
  NAND2_X1 U6390 ( .A1(n4967), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4968) );
  NAND2_X1 U6391 ( .A1(n4969), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4970) );
  XNOR2_X1 U6392 ( .A(n4970), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U6393 ( .A1(n4345), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4971) );
  MUX2_X1 U6394 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4971), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n4972) );
  NAND2_X1 U6395 ( .A1(n4977), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4978) );
  XNOR2_X1 U6396 ( .A(n4978), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U6397 ( .A1(n4324), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4979) );
  MUX2_X1 U6398 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4979), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n4980) );
  NAND2_X1 U6399 ( .A1(n4980), .A2(n4977), .ZN(n8955) );
  NAND2_X1 U6400 ( .A1(n6091), .A2(n8955), .ZN(n9179) );
  INV_X1 U6401 ( .A(n4981), .ZN(n4982) );
  NAND2_X1 U6402 ( .A1(n4982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4985) );
  INV_X1 U6403 ( .A(n4985), .ZN(n4983) );
  NAND2_X1 U6404 ( .A1(n4983), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n4986) );
  INV_X1 U6405 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4984) );
  NAND2_X1 U6406 ( .A1(n4985), .A2(n4984), .ZN(n5691) );
  NAND2_X1 U6407 ( .A1(n9410), .A2(n9184), .ZN(n9180) );
  NAND2_X1 U6408 ( .A1(n9520), .A2(n5047), .ZN(n5013) );
  NAND2_X1 U6409 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n4989) );
  INV_X1 U6410 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4991) );
  INV_X1 U6411 ( .A(n4994), .ZN(n4996) );
  NOR3_X1 U6412 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .A3(
        P1_IR_REG_30__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U6413 ( .A1(n4996), .A2(n4995), .ZN(n9652) );
  INV_X1 U6414 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n5000) );
  NAND2_X2 U6415 ( .A1(n5052), .A2(n9659), .ZN(n5994) );
  INV_X1 U6416 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9590) );
  OR2_X1 U6417 ( .A1(n6094), .A2(n9590), .ZN(n4999) );
  OAI21_X1 U6418 ( .B1(n5637), .B2(n5000), .A(n4999), .ZN(n5010) );
  OR2_X2 U6419 ( .A1(n5159), .A2(n5158), .ZN(n5206) );
  OR2_X2 U6420 ( .A1(n5206), .A2(n5205), .ZN(n5208) );
  INV_X1 U6421 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5178) );
  INV_X1 U6422 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5236) );
  OR2_X2 U6423 ( .A1(n5252), .A2(n5236), .ZN(n5276) );
  INV_X1 U6424 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5297) );
  OR2_X2 U6425 ( .A1(n5298), .A2(n5297), .ZN(n5326) );
  INV_X1 U6426 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5325) );
  OR2_X2 U6427 ( .A1(n5326), .A2(n5325), .ZN(n5346) );
  INV_X1 U6428 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5372) );
  INV_X1 U6429 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8865) );
  XNOR2_X1 U6430 ( .A(n5425), .B(n8865), .ZN(n9521) );
  INV_X1 U6431 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9638) );
  OR2_X1 U6432 ( .A1(n4278), .A2(n9638), .ZN(n5008) );
  OAI21_X1 U6433 ( .B1(n5704), .B2(n9521), .A(n5008), .ZN(n5009) );
  INV_X1 U6434 ( .A(n9179), .ZN(n5011) );
  NAND2_X2 U6435 ( .A1(n6529), .A2(n5011), .ZN(n5642) );
  NAND2_X1 U6436 ( .A1(n9194), .A2(n4429), .ZN(n5012) );
  NAND2_X1 U6437 ( .A1(n5013), .A2(n5012), .ZN(n5015) );
  XNOR2_X1 U6438 ( .A(n5015), .B(n5014), .ZN(n8858) );
  NAND2_X1 U6439 ( .A1(n9520), .A2(n4429), .ZN(n5018) );
  NAND2_X1 U6440 ( .A1(n9194), .A2(n5612), .ZN(n5017) );
  NAND2_X1 U6441 ( .A1(n5018), .A2(n5017), .ZN(n8859) );
  INV_X2 U6442 ( .A(n5501), .ZN(n5637) );
  INV_X1 U6443 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6941) );
  OR2_X1 U6444 ( .A1(n5637), .A2(n6941), .ZN(n5024) );
  OAI21_X1 U6445 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5129), .ZN(n7093) );
  OR2_X1 U6446 ( .A1(n5704), .A2(n7093), .ZN(n5023) );
  INV_X1 U6447 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5019) );
  OR2_X1 U6448 ( .A1(n5994), .A2(n5019), .ZN(n5022) );
  INV_X1 U6449 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5020) );
  OR2_X1 U6450 ( .A1(n4279), .A2(n5020), .ZN(n5021) );
  NAND2_X1 U6451 ( .A1(n5025), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5098) );
  INV_X1 U6452 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6453 ( .A1(n5098), .A2(n5097), .ZN(n5026) );
  NAND2_X1 U6454 ( .A1(n5026), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5027) );
  XNOR2_X1 U6455 ( .A(n5027), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6609) );
  INV_X1 U6456 ( .A(n6609), .ZN(n9240) );
  NAND2_X1 U6457 ( .A1(n5029), .A2(n5028), .ZN(n5031) );
  OR2_X1 U6458 ( .A1(n5987), .A2(n6535), .ZN(n5032) );
  OAI22_X1 U6459 ( .A1(n7209), .A2(n5016), .B1(n6943), .B2(n5642), .ZN(n5109)
         );
  INV_X1 U6460 ( .A(n7209), .ZN(n9208) );
  AOI22_X1 U6461 ( .A1(n9208), .A2(n4429), .B1(n9927), .B2(n5047), .ZN(n5033)
         );
  XNOR2_X1 U6462 ( .A(n5033), .B(n5014), .ZN(n5107) );
  INV_X1 U6463 ( .A(n5107), .ZN(n5108) );
  INV_X1 U6464 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n5034) );
  INV_X1 U6465 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5035) );
  OR2_X1 U6466 ( .A1(n5092), .A2(n5035), .ZN(n5039) );
  INV_X1 U6467 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5036) );
  OR2_X1 U6468 ( .A1(n4278), .A2(n5036), .ZN(n5038) );
  INV_X1 U6469 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9985) );
  OR2_X1 U6470 ( .A1(n5994), .A2(n9985), .ZN(n5037) );
  OR2_X1 U6471 ( .A1(n5041), .A2(n5229), .ZN(n5042) );
  INV_X1 U6472 ( .A(n6832), .ZN(n6534) );
  XNOR2_X1 U6473 ( .A(n5044), .B(n5043), .ZN(n6543) );
  OR2_X1 U6474 ( .A1(n5064), .A2(n6543), .ZN(n5046) );
  OR2_X1 U6475 ( .A1(n5096), .A2(n6533), .ZN(n5045) );
  INV_X1 U6476 ( .A(n6989), .ZN(n9917) );
  OAI22_X1 U6477 ( .A1(n6011), .A2(n5016), .B1(n9917), .B2(n5642), .ZN(n5087)
         );
  INV_X1 U6478 ( .A(n5087), .ZN(n5090) );
  OAI22_X1 U6479 ( .A1(n6011), .A2(n5642), .B1(n9917), .B2(n5243), .ZN(n5048)
         );
  XNOR2_X1 U6480 ( .A(n5048), .B(n5014), .ZN(n5088) );
  INV_X1 U6481 ( .A(n5088), .ZN(n5089) );
  INV_X1 U6482 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5049) );
  OR2_X1 U6483 ( .A1(n6095), .A2(n5049), .ZN(n5058) );
  INV_X1 U6484 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n5050) );
  INV_X1 U6485 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5051) );
  OR2_X1 U6486 ( .A1(n9659), .A2(n5051), .ZN(n5053) );
  OR2_X1 U6487 ( .A1(n5053), .A2(n5052), .ZN(n5056) );
  INV_X1 U6488 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5054) );
  OR2_X1 U6489 ( .A1(n5994), .A2(n5054), .ZN(n5055) );
  NAND4_X2 U6490 ( .A1(n5058), .A2(n5057), .A3(n5056), .A4(n5055), .ZN(n6007)
         );
  INV_X1 U6491 ( .A(n6007), .ZN(n6892) );
  INV_X1 U6492 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6531) );
  OR2_X1 U6493 ( .A1(n5096), .A2(n6531), .ZN(n5067) );
  NAND2_X1 U6494 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5059) );
  MUX2_X1 U6495 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5059), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5061) );
  INV_X1 U6496 ( .A(n5041), .ZN(n5060) );
  NAND2_X1 U6497 ( .A1(n5061), .A2(n5060), .ZN(n6604) );
  OR2_X1 U6498 ( .A1(n6567), .A2(n6604), .ZN(n5066) );
  XNOR2_X1 U6499 ( .A(n5063), .B(n5062), .ZN(n6154) );
  INV_X1 U6500 ( .A(n6154), .ZN(n6553) );
  OR2_X1 U6501 ( .A1(n5064), .A2(n6553), .ZN(n5065) );
  INV_X1 U6502 ( .A(n5083), .ZN(n5086) );
  NAND2_X1 U6503 ( .A1(n6007), .A2(n4429), .ZN(n5068) );
  INV_X1 U6504 ( .A(n5084), .ZN(n5085) );
  INV_X1 U6505 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5069) );
  INV_X1 U6506 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5070) );
  INV_X1 U6507 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5071) );
  OR2_X1 U6508 ( .A1(n5092), .A2(n5071), .ZN(n5073) );
  INV_X1 U6509 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5081) );
  OR2_X1 U6510 ( .A1(n5994), .A2(n5081), .ZN(n5072) );
  INV_X1 U6511 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5076) );
  XNOR2_X1 U6512 ( .A(n5077), .B(n5076), .ZN(n9660) );
  MUX2_X1 U6513 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9660), .S(n6567), .Z(n6904) );
  INV_X1 U6514 ( .A(n5080), .ZN(n5082) );
  INV_X1 U6515 ( .A(n9212), .ZN(n6857) );
  INV_X1 U6516 ( .A(n6904), .ZN(n6891) );
  INV_X1 U6517 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9730) );
  OAI21_X1 U6518 ( .B1(n6529), .B2(n5081), .A(n5080), .ZN(n6820) );
  NAND2_X1 U6519 ( .A1(n6821), .A2(n6820), .ZN(n6819) );
  OAI21_X1 U6520 ( .B1(n5082), .B2(n5014), .A(n6819), .ZN(n6854) );
  XNOR2_X1 U6521 ( .A(n5084), .B(n5083), .ZN(n6855) );
  XNOR2_X1 U6522 ( .A(n5088), .B(n5087), .ZN(n6771) );
  INV_X1 U6523 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5091) );
  OR2_X1 U6524 ( .A1(n4278), .A2(n5091), .ZN(n6013) );
  INV_X1 U6525 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6596) );
  OR2_X1 U6526 ( .A1(n5092), .A2(n6596), .ZN(n6014) );
  INV_X1 U6527 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6607) );
  OR2_X1 U6528 ( .A1(n5994), .A2(n6607), .ZN(n6012) );
  NAND4_X1 U6529 ( .A1(n6013), .A2(n6014), .A3(n6015), .A4(n6012), .ZN(n6067)
         );
  NAND2_X1 U6530 ( .A1(n6067), .A2(n5612), .ZN(n5103) );
  XNOR2_X1 U6531 ( .A(n5095), .B(n5094), .ZN(n6539) );
  OR2_X1 U6532 ( .A1(n5064), .A2(n6539), .ZN(n5101) );
  OR2_X1 U6533 ( .A1(n5096), .A2(n6532), .ZN(n5100) );
  XNOR2_X1 U6534 ( .A(n5098), .B(n5097), .ZN(n9224) );
  OR2_X1 U6535 ( .A1(n6567), .A2(n9224), .ZN(n5099) );
  OR2_X1 U6536 ( .A1(n9921), .A2(n5642), .ZN(n5102) );
  NAND2_X1 U6537 ( .A1(n5103), .A2(n5102), .ZN(n5106) );
  INV_X1 U6538 ( .A(n9921), .ZN(n9885) );
  AOI22_X1 U6539 ( .A1(n4429), .A2(n6067), .B1(n9885), .B2(n5047), .ZN(n5104)
         );
  XNOR2_X1 U6540 ( .A(n5104), .B(n5014), .ZN(n5105) );
  XOR2_X1 U6541 ( .A(n5106), .B(n5105), .Z(n6951) );
  XOR2_X1 U6542 ( .A(n5109), .B(n5107), .Z(n7087) );
  INV_X1 U6543 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7075) );
  OR2_X1 U6544 ( .A1(n5637), .A2(n7075), .ZN(n5117) );
  INV_X1 U6545 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6546 ( .A1(n5131), .A2(n5110), .ZN(n5111) );
  NAND2_X1 U6547 ( .A1(n5159), .A2(n5111), .ZN(n7361) );
  OR2_X1 U6548 ( .A1(n5704), .A2(n7361), .ZN(n5116) );
  INV_X1 U6549 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5112) );
  OR2_X1 U6550 ( .A1(n4278), .A2(n5112), .ZN(n5115) );
  INV_X1 U6551 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5113) );
  OR2_X1 U6552 ( .A1(n5994), .A2(n5113), .ZN(n5114) );
  NAND2_X1 U6553 ( .A1(n5118), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5119) );
  XNOR2_X1 U6554 ( .A(n5119), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6613) );
  INV_X1 U6555 ( .A(n6613), .ZN(n9764) );
  XNOR2_X1 U6556 ( .A(n5121), .B(n5120), .ZN(n6550) );
  OR2_X1 U6557 ( .A1(n5064), .A2(n6550), .ZN(n5123) );
  OR2_X1 U6558 ( .A1(n5987), .A2(n8651), .ZN(n5122) );
  OAI211_X1 U6559 ( .C1(n6567), .C2(n9764), .A(n5123), .B(n5122), .ZN(n7363)
         );
  OAI22_X1 U6560 ( .A1(n7230), .A2(n5642), .B1(n9940), .B2(n5243), .ZN(n5124)
         );
  XNOR2_X1 U6561 ( .A(n5124), .B(n5014), .ZN(n7355) );
  OAI22_X1 U6562 ( .A1(n7230), .A2(n5016), .B1(n9940), .B2(n5642), .ZN(n7356)
         );
  NAND2_X1 U6563 ( .A1(n7355), .A2(n7356), .ZN(n5151) );
  INV_X1 U6564 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5127) );
  INV_X1 U6565 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5125) );
  OR2_X1 U6566 ( .A1(n5994), .A2(n5125), .ZN(n5126) );
  OAI21_X1 U6567 ( .B1(n5637), .B2(n5127), .A(n5126), .ZN(n5135) );
  INV_X1 U6568 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5128) );
  NAND2_X1 U6569 ( .A1(n5129), .A2(n5128), .ZN(n5130) );
  NAND2_X1 U6570 ( .A1(n5131), .A2(n5130), .ZN(n9868) );
  INV_X1 U6571 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5132) );
  OR2_X1 U6572 ( .A1(n4279), .A2(n5132), .ZN(n5133) );
  OAI21_X1 U6573 ( .B1(n5704), .B2(n9868), .A(n5133), .ZN(n5134) );
  NAND2_X1 U6574 ( .A1(n9207), .A2(n4429), .ZN(n5144) );
  XNOR2_X1 U6575 ( .A(n5137), .B(n5136), .ZN(n6546) );
  OR2_X1 U6576 ( .A1(n5064), .A2(n6546), .ZN(n5142) );
  OR2_X1 U6577 ( .A1(n5987), .A2(n6545), .ZN(n5141) );
  OR2_X1 U6578 ( .A1(n5138), .A2(n5229), .ZN(n5139) );
  XNOR2_X1 U6579 ( .A(n5139), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6612) );
  INV_X1 U6580 ( .A(n6612), .ZN(n9749) );
  OR2_X1 U6581 ( .A1(n6567), .A2(n9749), .ZN(n5140) );
  OR2_X1 U6582 ( .A1(n9934), .A2(n5243), .ZN(n5143) );
  NAND2_X1 U6583 ( .A1(n5144), .A2(n5143), .ZN(n5145) );
  XNOR2_X1 U6584 ( .A(n5145), .B(n5666), .ZN(n7354) );
  INV_X1 U6585 ( .A(n7354), .ZN(n5149) );
  NAND2_X1 U6586 ( .A1(n9207), .A2(n5612), .ZN(n5147) );
  OR2_X1 U6587 ( .A1(n9934), .A2(n5642), .ZN(n5146) );
  NAND3_X1 U6588 ( .A1(n5151), .A2(n7354), .A3(n7207), .ZN(n5153) );
  OR2_X1 U6589 ( .A1(n7355), .A2(n7356), .ZN(n5152) );
  INV_X1 U6590 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5157) );
  INV_X1 U6591 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6603) );
  OR2_X1 U6592 ( .A1(n5994), .A2(n6603), .ZN(n5156) );
  OAI21_X1 U6593 ( .B1(n5637), .B2(n5157), .A(n5156), .ZN(n5164) );
  NAND2_X1 U6594 ( .A1(n5159), .A2(n5158), .ZN(n5160) );
  NAND2_X1 U6595 ( .A1(n5206), .A2(n5160), .ZN(n9855) );
  INV_X1 U6596 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5161) );
  OR2_X1 U6597 ( .A1(n4279), .A2(n5161), .ZN(n5162) );
  OAI21_X1 U6598 ( .B1(n5704), .B2(n9855), .A(n5162), .ZN(n5163) );
  NAND2_X1 U6599 ( .A1(n5165), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5166) );
  XNOR2_X1 U6600 ( .A(n5166), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9683) );
  AOI22_X1 U6601 ( .A1(n5419), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5418), .B2(
        n9683), .ZN(n5170) );
  XNOR2_X1 U6602 ( .A(n5168), .B(n5167), .ZN(n6551) );
  NAND2_X1 U6603 ( .A1(n6551), .A2(n5199), .ZN(n5169) );
  OAI22_X1 U6604 ( .A1(n7069), .A2(n5016), .B1(n9946), .B2(n5642), .ZN(n5175)
         );
  NAND2_X1 U6605 ( .A1(n9205), .A2(n4429), .ZN(n5172) );
  OR2_X1 U6606 ( .A1(n9946), .A2(n5243), .ZN(n5171) );
  NAND2_X1 U6607 ( .A1(n5172), .A2(n5171), .ZN(n5173) );
  XNOR2_X1 U6608 ( .A(n5173), .B(n5014), .ZN(n5174) );
  XOR2_X1 U6609 ( .A(n5175), .B(n5174), .Z(n7227) );
  INV_X1 U6610 ( .A(n5174), .ZN(n5177) );
  INV_X1 U6611 ( .A(n5175), .ZN(n5176) );
  INV_X1 U6612 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7331) );
  OR2_X1 U6613 ( .A1(n5637), .A2(n7331), .ZN(n5185) );
  NAND2_X1 U6614 ( .A1(n5208), .A2(n5178), .ZN(n5179) );
  NAND2_X1 U6615 ( .A1(n5250), .A2(n5179), .ZN(n7557) );
  OR2_X1 U6616 ( .A1(n5704), .A2(n7557), .ZN(n5184) );
  INV_X1 U6617 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5180) );
  OR2_X1 U6618 ( .A1(n5994), .A2(n5180), .ZN(n5183) );
  INV_X1 U6619 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5181) );
  OR2_X1 U6620 ( .A1(n4278), .A2(n5181), .ZN(n5182) );
  INV_X1 U6621 ( .A(n7287), .ZN(n9203) );
  OR2_X1 U6622 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  NAND2_X1 U6623 ( .A1(n5189), .A2(n5188), .ZN(n6570) );
  NAND2_X1 U6624 ( .A1(n6570), .A2(n5199), .ZN(n5193) );
  NAND2_X1 U6625 ( .A1(n5190), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5191) );
  XNOR2_X1 U6626 ( .A(n5191), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6870) );
  AOI22_X1 U6627 ( .A1(n5419), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5418), .B2(
        n6870), .ZN(n5192) );
  AOI22_X1 U6628 ( .A1(n4429), .A2(n9203), .B1(n9959), .B2(n5047), .ZN(n5194)
         );
  XNOR2_X1 U6629 ( .A(n5194), .B(n5014), .ZN(n7554) );
  OR2_X1 U6630 ( .A1(n7287), .A2(n5016), .ZN(n5196) );
  NAND2_X1 U6631 ( .A1(n9959), .A2(n4429), .ZN(n5195) );
  NAND2_X1 U6632 ( .A1(n7554), .A2(n7553), .ZN(n5218) );
  XNOR2_X1 U6633 ( .A(n5198), .B(n5197), .ZN(n6557) );
  NAND2_X1 U6634 ( .A1(n6557), .A2(n5199), .ZN(n5202) );
  OAI21_X1 U6635 ( .B1(n5165), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5200) );
  XNOR2_X1 U6636 ( .A(n5200), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9696) );
  AOI22_X1 U6637 ( .A1(n5419), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5418), .B2(
        n9696), .ZN(n5201) );
  INV_X1 U6638 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7242) );
  INV_X1 U6639 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5203) );
  OR2_X1 U6640 ( .A1(n4278), .A2(n5203), .ZN(n5204) );
  OAI21_X1 U6641 ( .B1(n5637), .B2(n7242), .A(n5204), .ZN(n5212) );
  NAND2_X1 U6642 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  NAND2_X1 U6643 ( .A1(n5208), .A2(n5207), .ZN(n7460) );
  INV_X1 U6644 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5209) );
  OR2_X1 U6645 ( .A1(n5994), .A2(n5209), .ZN(n5210) );
  OAI21_X1 U6646 ( .B1(n5704), .B2(n7460), .A(n5210), .ZN(n5211) );
  NAND2_X1 U6647 ( .A1(n9204), .A2(n4429), .ZN(n5213) );
  OAI21_X1 U6648 ( .B1(n9953), .B2(n5243), .A(n5213), .ZN(n5214) );
  XNOR2_X1 U6649 ( .A(n5214), .B(n5014), .ZN(n7551) );
  OR2_X1 U6650 ( .A1(n9953), .A2(n5642), .ZN(n5216) );
  NAND2_X1 U6651 ( .A1(n9204), .A2(n5612), .ZN(n5215) );
  NAND2_X1 U6652 ( .A1(n5216), .A2(n5215), .ZN(n7453) );
  NAND3_X1 U6653 ( .A1(n7552), .A2(n5218), .A3(n5217), .ZN(n5226) );
  INV_X1 U6654 ( .A(n5221), .ZN(n5223) );
  INV_X1 U6655 ( .A(n7553), .ZN(n5220) );
  INV_X1 U6656 ( .A(n7554), .ZN(n5219) );
  OAI21_X1 U6657 ( .B1(n5221), .B2(n5220), .A(n5219), .ZN(n5222) );
  INV_X1 U6658 ( .A(n5224), .ZN(n5225) );
  NAND2_X1 U6659 ( .A1(n5226), .A2(n5225), .ZN(n7622) );
  XNOR2_X1 U6660 ( .A(n5228), .B(n5227), .ZN(n6581) );
  NAND2_X1 U6661 ( .A1(n6581), .A2(n5986), .ZN(n5234) );
  NOR2_X1 U6662 ( .A1(n5190), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5318) );
  OR2_X1 U6663 ( .A1(n5318), .A2(n5229), .ZN(n5271) );
  NAND2_X1 U6664 ( .A1(n5271), .A2(n5230), .ZN(n5231) );
  NAND2_X1 U6665 ( .A1(n5231), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5232) );
  XNOR2_X1 U6666 ( .A(n5232), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9769) );
  AOI22_X1 U6667 ( .A1(n5419), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5418), .B2(
        n9769), .ZN(n5233) );
  INV_X1 U6668 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5235) );
  OR2_X1 U6669 ( .A1(n5637), .A2(n5235), .ZN(n5242) );
  NAND2_X1 U6670 ( .A1(n5252), .A2(n5236), .ZN(n5237) );
  NAND2_X1 U6671 ( .A1(n5276), .A2(n5237), .ZN(n9839) );
  OR2_X1 U6672 ( .A1(n5704), .A2(n9839), .ZN(n5241) );
  INV_X1 U6673 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5238) );
  OR2_X1 U6674 ( .A1(n4278), .A2(n5238), .ZN(n5240) );
  INV_X1 U6675 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6871) );
  OR2_X1 U6676 ( .A1(n6094), .A2(n6871), .ZN(n5239) );
  NOR2_X1 U6677 ( .A1(n9201), .A2(n5016), .ZN(n5244) );
  AOI21_X1 U6678 ( .B1(n9841), .B2(n4429), .A(n5244), .ZN(n7624) );
  XNOR2_X1 U6679 ( .A(n5246), .B(n5245), .ZN(n6575) );
  NAND2_X1 U6680 ( .A1(n6575), .A2(n5986), .ZN(n5248) );
  XNOR2_X1 U6681 ( .A(n5271), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9669) );
  AOI22_X1 U6682 ( .A1(n5419), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5418), .B2(
        n9669), .ZN(n5247) );
  INV_X1 U6683 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6684 ( .A1(n5250), .A2(n5249), .ZN(n5251) );
  NAND2_X1 U6685 ( .A1(n5252), .A2(n5251), .ZN(n7578) );
  OR2_X1 U6686 ( .A1(n5704), .A2(n7578), .ZN(n5257) );
  INV_X1 U6687 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7292) );
  OR2_X1 U6688 ( .A1(n5637), .A2(n7292), .ZN(n5256) );
  INV_X1 U6689 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5253) );
  OR2_X1 U6690 ( .A1(n4278), .A2(n5253), .ZN(n5255) );
  INV_X1 U6691 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6868) );
  OR2_X1 U6692 ( .A1(n5994), .A2(n6868), .ZN(n5254) );
  NOR2_X1 U6693 ( .A1(n7540), .A2(n5016), .ZN(n5258) );
  AOI21_X1 U6694 ( .B1(n7574), .B2(n4429), .A(n5258), .ZN(n7573) );
  NAND2_X1 U6695 ( .A1(n7574), .A2(n5047), .ZN(n5260) );
  INV_X1 U6696 ( .A(n7540), .ZN(n9202) );
  NAND2_X1 U6697 ( .A1(n9202), .A2(n4429), .ZN(n5259) );
  NAND2_X1 U6698 ( .A1(n5260), .A2(n5259), .ZN(n5261) );
  XNOR2_X1 U6699 ( .A(n5261), .B(n5666), .ZN(n7571) );
  OAI22_X1 U6700 ( .A1(n7625), .A2(n7624), .B1(n7573), .B2(n7571), .ZN(n5266)
         );
  NAND3_X1 U6701 ( .A1(n7624), .A2(n7573), .A3(n7571), .ZN(n5265) );
  INV_X1 U6702 ( .A(n7571), .ZN(n7623) );
  INV_X1 U6703 ( .A(n7573), .ZN(n5262) );
  NOR2_X1 U6704 ( .A1(n7623), .A2(n5262), .ZN(n5263) );
  OAI21_X1 U6705 ( .B1(n7624), .B2(n5263), .A(n7625), .ZN(n5264) );
  XNOR2_X1 U6706 ( .A(n5267), .B(n5268), .ZN(n6630) );
  NAND2_X1 U6707 ( .A1(n6630), .A2(n5986), .ZN(n5274) );
  NAND2_X1 U6708 ( .A1(n5269), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6709 ( .A1(n5271), .A2(n5270), .ZN(n5291) );
  XNOR2_X1 U6710 ( .A(n5291), .B(n5272), .ZN(n9264) );
  AOI22_X1 U6711 ( .A1(n5419), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5418), .B2(
        n9264), .ZN(n5273) );
  NAND2_X1 U6712 ( .A1(n7523), .A2(n5047), .ZN(n5285) );
  INV_X1 U6713 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7401) );
  OR2_X1 U6714 ( .A1(n5637), .A2(n7401), .ZN(n5283) );
  INV_X1 U6715 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5275) );
  NAND2_X1 U6716 ( .A1(n5276), .A2(n5275), .ZN(n5277) );
  NAND2_X1 U6717 ( .A1(n5298), .A2(n5277), .ZN(n7518) );
  OR2_X1 U6718 ( .A1(n5704), .A2(n7518), .ZN(n5282) );
  INV_X1 U6719 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5278) );
  OR2_X1 U6720 ( .A1(n4279), .A2(n5278), .ZN(n5281) );
  INV_X1 U6721 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5279) );
  OR2_X1 U6722 ( .A1(n6094), .A2(n5279), .ZN(n5280) );
  NAND2_X1 U6723 ( .A1(n9200), .A2(n4429), .ZN(n5284) );
  NAND2_X1 U6724 ( .A1(n5285), .A2(n5284), .ZN(n5286) );
  XNOR2_X1 U6725 ( .A(n5286), .B(n5014), .ZN(n5287) );
  AOI22_X1 U6726 ( .A1(n7523), .A2(n4429), .B1(n5612), .B2(n9200), .ZN(n5288)
         );
  XNOR2_X1 U6727 ( .A(n5287), .B(n5288), .ZN(n7517) );
  INV_X1 U6728 ( .A(n5287), .ZN(n5289) );
  XNOR2_X1 U6729 ( .A(n5359), .B(n5290), .ZN(n6635) );
  NAND2_X1 U6730 ( .A1(n6635), .A2(n5986), .ZN(n5294) );
  OAI21_X1 U6731 ( .B1(n5291), .B2(P1_IR_REG_12__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5292) );
  XNOR2_X1 U6732 ( .A(n5292), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9796) );
  AOI22_X1 U6733 ( .A1(n5419), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5418), .B2(
        n9796), .ZN(n5293) );
  INV_X1 U6734 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7419) );
  INV_X1 U6735 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5295) );
  OR2_X1 U6736 ( .A1(n6094), .A2(n5295), .ZN(n5296) );
  OAI21_X1 U6737 ( .B1(n5637), .B2(n7419), .A(n5296), .ZN(n5303) );
  NAND2_X1 U6738 ( .A1(n5298), .A2(n5297), .ZN(n5299) );
  NAND2_X1 U6739 ( .A1(n5326), .A2(n5299), .ZN(n7606) );
  INV_X1 U6740 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5300) );
  OR2_X1 U6741 ( .A1(n4279), .A2(n5300), .ZN(n5301) );
  OAI21_X1 U6742 ( .B1(n5704), .B2(n7606), .A(n5301), .ZN(n5302) );
  AOI22_X1 U6743 ( .A1(n9005), .A2(n4429), .B1(n5612), .B2(n9199), .ZN(n5307)
         );
  NAND2_X1 U6744 ( .A1(n9005), .A2(n5047), .ZN(n5305) );
  NAND2_X1 U6745 ( .A1(n9199), .A2(n4429), .ZN(n5304) );
  NAND2_X1 U6746 ( .A1(n5305), .A2(n5304), .ZN(n5306) );
  XNOR2_X1 U6747 ( .A(n5306), .B(n5014), .ZN(n5309) );
  XOR2_X1 U6748 ( .A(n5307), .B(n5309), .Z(n7602) );
  INV_X1 U6749 ( .A(n5307), .ZN(n5308) );
  NAND2_X1 U6750 ( .A1(n5359), .A2(n5310), .ZN(n5312) );
  NAND2_X1 U6751 ( .A1(n5312), .A2(n5311), .ZN(n5314) );
  XNOR2_X1 U6752 ( .A(n5314), .B(n5313), .ZN(n6639) );
  NAND2_X1 U6753 ( .A1(n6639), .A2(n5986), .ZN(n5323) );
  NOR2_X1 U6754 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5315) );
  AND2_X1 U6755 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  NAND2_X1 U6756 ( .A1(n5318), .A2(n5317), .ZN(n5320) );
  NAND2_X1 U6757 ( .A1(n5320), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5319) );
  MUX2_X1 U6758 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5319), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5321) );
  OR2_X1 U6759 ( .A1(n5320), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5339) );
  AND2_X1 U6760 ( .A1(n5321), .A2(n5339), .ZN(n9808) );
  AOI22_X1 U6761 ( .A1(n5419), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5418), .B2(
        n9808), .ZN(n5322) );
  INV_X1 U6762 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9260) );
  INV_X1 U6763 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9253) );
  OR2_X1 U6764 ( .A1(n6094), .A2(n9253), .ZN(n5324) );
  OAI21_X1 U6765 ( .B1(n5637), .B2(n9260), .A(n5324), .ZN(n5331) );
  NAND2_X1 U6766 ( .A1(n5326), .A2(n5325), .ZN(n5327) );
  NAND2_X1 U6767 ( .A1(n5346), .A2(n5327), .ZN(n7651) );
  INV_X1 U6768 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5328) );
  OR2_X1 U6769 ( .A1(n4279), .A2(n5328), .ZN(n5329) );
  OAI21_X1 U6770 ( .B1(n5704), .B2(n7651), .A(n5329), .ZN(n5330) );
  AOI22_X1 U6771 ( .A1(n9973), .A2(n5047), .B1(n4429), .B2(n9198), .ZN(n5332)
         );
  XNOR2_X1 U6772 ( .A(n5332), .B(n5014), .ZN(n5333) );
  INV_X1 U6773 ( .A(n9973), .ZN(n7650) );
  INV_X1 U6774 ( .A(n9198), .ZN(n6076) );
  OAI22_X1 U6775 ( .A1(n7650), .A2(n5642), .B1(n6076), .B2(n5016), .ZN(n7633)
         );
  INV_X1 U6776 ( .A(n5333), .ZN(n7634) );
  NAND2_X1 U6777 ( .A1(n5359), .A2(n5334), .ZN(n5336) );
  AND2_X1 U6778 ( .A1(n5336), .A2(n5335), .ZN(n5338) );
  NAND2_X1 U6779 ( .A1(n6665), .A2(n5986), .ZN(n5342) );
  NAND2_X1 U6780 ( .A1(n5339), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5340) );
  XNOR2_X1 U6781 ( .A(n5340), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9819) );
  AOI22_X1 U6782 ( .A1(n5419), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5418), .B2(
        n9819), .ZN(n5341) );
  NAND2_X1 U6783 ( .A1(n9011), .A2(n5047), .ZN(n5353) );
  INV_X1 U6784 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7658) );
  INV_X1 U6785 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5343) );
  OR2_X1 U6786 ( .A1(n4279), .A2(n5343), .ZN(n5344) );
  OAI21_X1 U6787 ( .B1(n5637), .B2(n7658), .A(n5344), .ZN(n5351) );
  INV_X1 U6788 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U6789 ( .A1(n5346), .A2(n5345), .ZN(n5347) );
  NAND2_X1 U6790 ( .A1(n5373), .A2(n5347), .ZN(n8892) );
  INV_X1 U6791 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5348) );
  OR2_X1 U6792 ( .A1(n6094), .A2(n5348), .ZN(n5349) );
  OAI21_X1 U6793 ( .B1(n5704), .B2(n8892), .A(n5349), .ZN(n5350) );
  NAND2_X1 U6794 ( .A1(n9197), .A2(n4429), .ZN(n5352) );
  NAND2_X1 U6795 ( .A1(n5353), .A2(n5352), .ZN(n5354) );
  XNOR2_X1 U6796 ( .A(n5354), .B(n5014), .ZN(n5356) );
  AOI22_X1 U6797 ( .A1(n9011), .A2(n4429), .B1(n5612), .B2(n9197), .ZN(n8886)
         );
  INV_X1 U6798 ( .A(n5355), .ZN(n5357) );
  NAND2_X1 U6799 ( .A1(n8884), .A2(n4856), .ZN(n8820) );
  NAND2_X1 U6800 ( .A1(n5359), .A2(n5358), .ZN(n5362) );
  NAND2_X1 U6801 ( .A1(n5362), .A2(n5360), .ZN(n5366) );
  NAND2_X1 U6802 ( .A1(n5362), .A2(n5361), .ZN(n5364) );
  NAND2_X1 U6803 ( .A1(n5364), .A2(n5363), .ZN(n5365) );
  NAND2_X1 U6804 ( .A1(n6653), .A2(n5986), .ZN(n5370) );
  NAND2_X1 U6805 ( .A1(n5367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5368) );
  XNOR2_X1 U6806 ( .A(n5368), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9281) );
  AOI22_X1 U6807 ( .A1(n5419), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5418), .B2(
        n9281), .ZN(n5369) );
  NAND2_X1 U6808 ( .A1(n8825), .A2(n5047), .ZN(n5380) );
  INV_X1 U6809 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5371) );
  OR2_X1 U6810 ( .A1(n5637), .A2(n5371), .ZN(n5378) );
  NAND2_X1 U6811 ( .A1(n5373), .A2(n5372), .ZN(n5374) );
  NAND2_X1 U6812 ( .A1(n5396), .A2(n5374), .ZN(n8821) );
  OR2_X1 U6813 ( .A1(n5704), .A2(n8821), .ZN(n5377) );
  INV_X1 U6814 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9643) );
  OR2_X1 U6815 ( .A1(n4279), .A2(n9643), .ZN(n5376) );
  INV_X1 U6816 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9600) );
  OR2_X1 U6817 ( .A1(n6094), .A2(n9600), .ZN(n5375) );
  NAND2_X1 U6818 ( .A1(n9196), .A2(n4429), .ZN(n5379) );
  NAND2_X1 U6819 ( .A1(n5380), .A2(n5379), .ZN(n5381) );
  XNOR2_X1 U6820 ( .A(n5381), .B(n5014), .ZN(n5384) );
  AOI22_X1 U6821 ( .A1(n8825), .A2(n4429), .B1(n5612), .B2(n9196), .ZN(n5382)
         );
  XNOR2_X1 U6822 ( .A(n5384), .B(n5382), .ZN(n8819) );
  INV_X1 U6823 ( .A(n5382), .ZN(n5383) );
  NAND2_X1 U6824 ( .A1(n5387), .A2(n5386), .ZN(n5389) );
  NAND2_X1 U6825 ( .A1(n5389), .A2(n5388), .ZN(n6649) );
  NAND2_X1 U6826 ( .A1(n6649), .A2(n5986), .ZN(n5392) );
  XNOR2_X1 U6827 ( .A(n5390), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9298) );
  AOI22_X1 U6828 ( .A1(n5419), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5418), .B2(
        n9298), .ZN(n5391) );
  NAND2_X1 U6829 ( .A1(n9594), .A2(n5047), .ZN(n5403) );
  INV_X1 U6830 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9280) );
  INV_X1 U6831 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n5393) );
  OR2_X1 U6832 ( .A1(n4278), .A2(n5393), .ZN(n5394) );
  OAI21_X1 U6833 ( .B1(n5637), .B2(n9280), .A(n5394), .ZN(n5401) );
  INV_X1 U6834 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5395) );
  NAND2_X1 U6835 ( .A1(n5396), .A2(n5395), .ZN(n5397) );
  NAND2_X1 U6836 ( .A1(n5425), .A2(n5397), .ZN(n8830) );
  INV_X1 U6837 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n5398) );
  OR2_X1 U6838 ( .A1(n6094), .A2(n5398), .ZN(n5399) );
  OAI21_X1 U6839 ( .B1(n5704), .B2(n8830), .A(n5399), .ZN(n5400) );
  NAND2_X1 U6840 ( .A1(n9195), .A2(n4429), .ZN(n5402) );
  NAND2_X1 U6841 ( .A1(n5403), .A2(n5402), .ZN(n5404) );
  XNOR2_X1 U6842 ( .A(n5404), .B(n5014), .ZN(n5405) );
  AOI22_X1 U6843 ( .A1(n9594), .A2(n4429), .B1(n5612), .B2(n9195), .ZN(n5406)
         );
  XNOR2_X1 U6844 ( .A(n5405), .B(n5406), .ZN(n8829) );
  INV_X1 U6845 ( .A(n5405), .ZN(n5407) );
  INV_X1 U6846 ( .A(n5408), .ZN(n5412) );
  INV_X1 U6847 ( .A(n5409), .ZN(n5410) );
  NAND2_X1 U6848 ( .A1(n5410), .A2(SI_18_), .ZN(n5411) );
  INV_X1 U6849 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6899) );
  INV_X1 U6850 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6949) );
  INV_X1 U6851 ( .A(SI_19_), .ZN(n5414) );
  NAND2_X1 U6852 ( .A1(n5415), .A2(n5414), .ZN(n5436) );
  INV_X1 U6853 ( .A(n5415), .ZN(n5416) );
  NAND2_X1 U6854 ( .A1(n5416), .A2(SI_19_), .ZN(n5417) );
  NAND2_X1 U6855 ( .A1(n5436), .A2(n5417), .ZN(n5437) );
  XNOR2_X1 U6856 ( .A(n5438), .B(n5437), .ZN(n6898) );
  NAND2_X1 U6857 ( .A1(n6898), .A2(n5986), .ZN(n5421) );
  INV_X1 U6858 ( .A(n9410), .ZN(n9308) );
  AOI22_X1 U6859 ( .A1(n5419), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9308), .B2(
        n5418), .ZN(n5420) );
  NAND2_X1 U6860 ( .A1(n9500), .A2(n5047), .ZN(n5431) );
  INV_X1 U6861 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9503) );
  INV_X1 U6862 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9585) );
  OR2_X1 U6863 ( .A1(n6094), .A2(n9585), .ZN(n5422) );
  OAI21_X1 U6864 ( .B1(n5637), .B2(n9503), .A(n5422), .ZN(n5429) );
  INV_X1 U6865 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5423) );
  OAI21_X1 U6866 ( .B1(n5425), .B2(n8865), .A(n5423), .ZN(n5426) );
  NAND2_X1 U6867 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5424) );
  OR2_X2 U6868 ( .A1(n5425), .A2(n5424), .ZN(n5445) );
  NAND2_X1 U6869 ( .A1(n5426), .A2(n5445), .ZN(n9502) );
  INV_X1 U6870 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9634) );
  OR2_X1 U6871 ( .A1(n4279), .A2(n9634), .ZN(n5427) );
  OAI21_X1 U6872 ( .B1(n5704), .B2(n9502), .A(n5427), .ZN(n5428) );
  NAND2_X1 U6873 ( .A1(n9193), .A2(n4429), .ZN(n5430) );
  NAND2_X1 U6874 ( .A1(n5431), .A2(n5430), .ZN(n5432) );
  XNOR2_X1 U6875 ( .A(n5432), .B(n5666), .ZN(n5435) );
  AND2_X1 U6876 ( .A1(n9193), .A2(n5612), .ZN(n5433) );
  AOI21_X1 U6877 ( .B1(n9500), .B2(n4429), .A(n5433), .ZN(n5434) );
  NOR2_X1 U6878 ( .A1(n5435), .A2(n5434), .ZN(n8790) );
  NAND2_X1 U6879 ( .A1(n5435), .A2(n5434), .ZN(n8794) );
  INV_X1 U6880 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6916) );
  INV_X1 U6881 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6917) );
  INV_X1 U6882 ( .A(SI_20_), .ZN(n5439) );
  NAND2_X1 U6883 ( .A1(n5440), .A2(n5439), .ZN(n5457) );
  INV_X1 U6884 ( .A(n5440), .ZN(n5441) );
  NAND2_X1 U6885 ( .A1(n5441), .A2(SI_20_), .ZN(n5442) );
  XNOR2_X1 U6886 ( .A(n5456), .B(n5455), .ZN(n6915) );
  NAND2_X1 U6887 ( .A1(n6915), .A2(n5986), .ZN(n5444) );
  OR2_X1 U6888 ( .A1(n5987), .A2(n6917), .ZN(n5443) );
  NAND2_X2 U6889 ( .A1(n5444), .A2(n5443), .ZN(n9484) );
  INV_X1 U6890 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8846) );
  OR2_X2 U6891 ( .A1(n5445), .A2(n8846), .ZN(n5462) );
  NAND2_X1 U6892 ( .A1(n5445), .A2(n8846), .ZN(n5446) );
  AND2_X1 U6893 ( .A1(n5462), .A2(n5446), .ZN(n9485) );
  NAND2_X1 U6894 ( .A1(n9485), .A2(n5632), .ZN(n5451) );
  INV_X1 U6895 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5447) );
  OR2_X1 U6896 ( .A1(n5637), .A2(n5447), .ZN(n5450) );
  INV_X1 U6897 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9580) );
  OR2_X1 U6898 ( .A1(n6094), .A2(n9580), .ZN(n5449) );
  INV_X1 U6899 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9631) );
  OR2_X1 U6900 ( .A1(n4279), .A2(n9631), .ZN(n5448) );
  NAND4_X1 U6901 ( .A1(n5451), .A2(n5450), .A3(n5449), .A4(n5448), .ZN(n9192)
         );
  INV_X1 U6902 ( .A(n9192), .ZN(n9468) );
  OAI22_X1 U6903 ( .A1(n6085), .A2(n5642), .B1(n9468), .B2(n5016), .ZN(n5473)
         );
  NAND2_X1 U6904 ( .A1(n9484), .A2(n5047), .ZN(n5453) );
  NAND2_X1 U6905 ( .A1(n9192), .A2(n4429), .ZN(n5452) );
  NAND2_X1 U6906 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  XNOR2_X1 U6907 ( .A(n5454), .B(n5014), .ZN(n5472) );
  XOR2_X1 U6908 ( .A(n5473), .B(n5472), .Z(n8844) );
  INV_X1 U6909 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6948) );
  INV_X1 U6910 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6956) );
  XNOR2_X1 U6911 ( .A(n5481), .B(SI_21_), .ZN(n5480) );
  XNOR2_X1 U6912 ( .A(n5485), .B(n5480), .ZN(n6947) );
  NAND2_X1 U6913 ( .A1(n6947), .A2(n5986), .ZN(n5460) );
  OR2_X1 U6914 ( .A1(n5987), .A2(n6956), .ZN(n5459) );
  NAND2_X1 U6915 ( .A1(n9574), .A2(n5047), .ZN(n5469) );
  INV_X1 U6916 ( .A(n5462), .ZN(n5461) );
  INV_X1 U6917 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8804) );
  NAND2_X1 U6918 ( .A1(n5462), .A2(n8804), .ZN(n5463) );
  NAND2_X1 U6919 ( .A1(n5498), .A2(n5463), .ZN(n9471) );
  INV_X1 U6920 ( .A(n4278), .ZN(n5464) );
  AOI22_X1 U6921 ( .A1(n5501), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n5464), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n5467) );
  INV_X1 U6922 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5465) );
  OR2_X1 U6923 ( .A1(n6094), .A2(n5465), .ZN(n5466) );
  OAI211_X1 U6924 ( .C1(n9471), .C2(n5704), .A(n5467), .B(n5466), .ZN(n9191)
         );
  NAND2_X1 U6925 ( .A1(n9191), .A2(n4429), .ZN(n5468) );
  NAND2_X1 U6926 ( .A1(n5469), .A2(n5468), .ZN(n5470) );
  XNOR2_X1 U6927 ( .A(n5470), .B(n5014), .ZN(n5477) );
  AOI22_X1 U6928 ( .A1(n9574), .A2(n4429), .B1(n5612), .B2(n9191), .ZN(n5478)
         );
  XNOR2_X1 U6929 ( .A(n5477), .B(n5478), .ZN(n8803) );
  AND2_X1 U6930 ( .A1(n8844), .A2(n8803), .ZN(n5471) );
  INV_X1 U6931 ( .A(n8803), .ZN(n5476) );
  INV_X1 U6932 ( .A(n5472), .ZN(n5475) );
  INV_X1 U6933 ( .A(n5473), .ZN(n5474) );
  NAND2_X1 U6934 ( .A1(n5475), .A2(n5474), .ZN(n8801) );
  INV_X1 U6935 ( .A(n5477), .ZN(n5479) );
  INV_X1 U6936 ( .A(n5480), .ZN(n5484) );
  INV_X1 U6937 ( .A(n5481), .ZN(n5482) );
  NAND2_X1 U6938 ( .A1(n5482), .A2(SI_21_), .ZN(n5483) );
  INV_X1 U6939 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7082) );
  INV_X1 U6940 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n5493) );
  INV_X1 U6941 ( .A(SI_22_), .ZN(n5486) );
  NAND2_X1 U6942 ( .A1(n5487), .A2(n5486), .ZN(n5511) );
  INV_X1 U6943 ( .A(n5487), .ZN(n5488) );
  NAND2_X1 U6944 ( .A1(n5488), .A2(SI_22_), .ZN(n5489) );
  NAND2_X1 U6945 ( .A1(n5511), .A2(n5489), .ZN(n5490) );
  NAND2_X1 U6946 ( .A1(n5491), .A2(n5490), .ZN(n5492) );
  NAND2_X1 U6947 ( .A1(n5512), .A2(n5492), .ZN(n7080) );
  NAND2_X1 U6948 ( .A1(n7080), .A2(n5986), .ZN(n5495) );
  OR2_X1 U6949 ( .A1(n5987), .A2(n5493), .ZN(n5494) );
  NAND2_X1 U6950 ( .A1(n9450), .A2(n5047), .ZN(n5505) );
  INV_X1 U6951 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9626) );
  INV_X1 U6952 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U6953 ( .A1(n5498), .A2(n5497), .ZN(n5499) );
  NAND2_X1 U6954 ( .A1(n5522), .A2(n5499), .ZN(n9451) );
  OR2_X1 U6955 ( .A1(n9451), .A2(n5704), .ZN(n5503) );
  AOI22_X1 U6956 ( .A1(n5501), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n5500), .B2(
        P1_REG1_REG_22__SCAN_IN), .ZN(n5502) );
  NAND2_X1 U6957 ( .A1(n9434), .A2(n4429), .ZN(n5504) );
  NAND2_X1 U6958 ( .A1(n5505), .A2(n5504), .ZN(n5506) );
  XNOR2_X1 U6959 ( .A(n5506), .B(n5014), .ZN(n5507) );
  AOI22_X1 U6960 ( .A1(n9450), .A2(n4429), .B1(n5612), .B2(n9434), .ZN(n8852)
         );
  NAND2_X1 U6961 ( .A1(n8851), .A2(n8852), .ZN(n8850) );
  INV_X1 U6962 ( .A(n5507), .ZN(n5508) );
  NAND2_X1 U6963 ( .A1(n5509), .A2(n5508), .ZN(n5510) );
  NAND2_X1 U6964 ( .A1(n8850), .A2(n5510), .ZN(n8779) );
  INV_X1 U6965 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5513) );
  INV_X1 U6966 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7150) );
  MUX2_X1 U6967 ( .A(n5513), .B(n7150), .S(n6530), .Z(n5514) );
  INV_X1 U6968 ( .A(SI_23_), .ZN(n8693) );
  NAND2_X1 U6969 ( .A1(n5514), .A2(n8693), .ZN(n5537) );
  INV_X1 U6970 ( .A(n5514), .ZN(n5515) );
  NAND2_X1 U6971 ( .A1(n5515), .A2(SI_23_), .ZN(n5516) );
  NAND2_X1 U6972 ( .A1(n5537), .A2(n5516), .ZN(n5517) );
  NAND2_X1 U6973 ( .A1(n4313), .A2(n5517), .ZN(n5519) );
  INV_X1 U6974 ( .A(n5517), .ZN(n5518) );
  NAND2_X1 U6975 ( .A1(n5519), .A2(n5538), .ZN(n7148) );
  NAND2_X1 U6976 ( .A1(n7148), .A2(n5986), .ZN(n5521) );
  OR2_X1 U6977 ( .A1(n5987), .A2(n7150), .ZN(n5520) );
  INV_X1 U6978 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8783) );
  NAND2_X1 U6979 ( .A1(n5522), .A2(n8783), .ZN(n5523) );
  AND2_X1 U6980 ( .A1(n5547), .A2(n5523), .ZN(n9424) );
  NAND2_X1 U6981 ( .A1(n9424), .A2(n5632), .ZN(n5530) );
  INV_X1 U6982 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5527) );
  INV_X1 U6983 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n8695) );
  OR2_X1 U6984 ( .A1(n6094), .A2(n8695), .ZN(n5526) );
  INV_X1 U6985 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n5524) );
  OR2_X1 U6986 ( .A1(n4279), .A2(n5524), .ZN(n5525) );
  OAI211_X1 U6987 ( .C1(n5637), .C2(n5527), .A(n5526), .B(n5525), .ZN(n5528)
         );
  INV_X1 U6988 ( .A(n5528), .ZN(n5529) );
  AOI22_X1 U6989 ( .A1(n9563), .A2(n5047), .B1(n4429), .B2(n9065), .ZN(n5531)
         );
  XOR2_X1 U6990 ( .A(n5014), .B(n5531), .Z(n5532) );
  OAI22_X1 U6991 ( .A1(n9426), .A2(n5642), .B1(n9447), .B2(n5016), .ZN(n5533)
         );
  NAND2_X1 U6992 ( .A1(n5532), .A2(n5533), .ZN(n8781) );
  NAND2_X1 U6993 ( .A1(n8779), .A2(n8781), .ZN(n5536) );
  INV_X1 U6994 ( .A(n5532), .ZN(n5535) );
  INV_X1 U6995 ( .A(n5533), .ZN(n5534) );
  NAND2_X1 U6996 ( .A1(n5535), .A2(n5534), .ZN(n8780) );
  INV_X1 U6997 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7369) );
  INV_X1 U6998 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7300) );
  MUX2_X1 U6999 ( .A(n7369), .B(n7300), .S(n6530), .Z(n5540) );
  INV_X1 U7000 ( .A(SI_24_), .ZN(n5539) );
  NAND2_X1 U7001 ( .A1(n5540), .A2(n5539), .ZN(n5563) );
  INV_X1 U7002 ( .A(n5540), .ZN(n5541) );
  NAND2_X1 U7003 ( .A1(n5541), .A2(SI_24_), .ZN(n5542) );
  AND2_X1 U7004 ( .A1(n5563), .A2(n5542), .ZN(n5562) );
  OR2_X1 U7005 ( .A1(n5987), .A2(n7300), .ZN(n5543) );
  NAND2_X1 U7006 ( .A1(n9416), .A2(n5047), .ZN(n5555) );
  INV_X1 U7007 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7008 ( .A1(n5547), .A2(n5546), .ZN(n5548) );
  NAND2_X1 U7009 ( .A1(n5576), .A2(n5548), .ZN(n9414) );
  INV_X1 U7010 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9413) );
  INV_X1 U7011 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9560) );
  OR2_X1 U7012 ( .A1(n6094), .A2(n9560), .ZN(n5550) );
  INV_X1 U7013 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9621) );
  OR2_X1 U7014 ( .A1(n4279), .A2(n9621), .ZN(n5549) );
  OAI211_X1 U7015 ( .C1(n5637), .C2(n9413), .A(n5550), .B(n5549), .ZN(n5551)
         );
  INV_X1 U7016 ( .A(n5551), .ZN(n5552) );
  NAND2_X1 U7017 ( .A1(n9432), .A2(n4429), .ZN(n5554) );
  NAND2_X1 U7018 ( .A1(n5555), .A2(n5554), .ZN(n5556) );
  XNOR2_X1 U7019 ( .A(n5556), .B(n5014), .ZN(n5560) );
  NAND2_X1 U7020 ( .A1(n9416), .A2(n4429), .ZN(n5558) );
  NAND2_X1 U7021 ( .A1(n9432), .A2(n5612), .ZN(n5557) );
  NAND2_X1 U7022 ( .A1(n5558), .A2(n5557), .ZN(n5559) );
  NOR2_X1 U7023 ( .A1(n5560), .A2(n5559), .ZN(n5588) );
  AOI21_X1 U7024 ( .B1(n5560), .B2(n5559), .A(n5588), .ZN(n8837) );
  INV_X1 U7025 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7751) );
  INV_X1 U7026 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7367) );
  INV_X1 U7027 ( .A(SI_25_), .ZN(n5564) );
  NAND2_X1 U7028 ( .A1(n5565), .A2(n5564), .ZN(n5593) );
  INV_X1 U7029 ( .A(n5565), .ZN(n5566) );
  NAND2_X1 U7030 ( .A1(n5566), .A2(SI_25_), .ZN(n5567) );
  NAND2_X1 U7031 ( .A1(n5593), .A2(n5567), .ZN(n5569) );
  NAND2_X1 U7032 ( .A1(n5568), .A2(n5569), .ZN(n5572) );
  INV_X1 U7033 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7034 ( .A1(n5572), .A2(n5594), .ZN(n7366) );
  NAND2_X1 U7035 ( .A1(n7366), .A2(n5986), .ZN(n5574) );
  OR2_X1 U7036 ( .A1(n5987), .A2(n7367), .ZN(n5573) );
  INV_X1 U7037 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7038 ( .A1(n5576), .A2(n5575), .ZN(n5577) );
  NAND2_X1 U7039 ( .A1(n9398), .A2(n5632), .ZN(n5585) );
  INV_X1 U7040 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n5582) );
  INV_X1 U7041 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5578) );
  OR2_X1 U7042 ( .A1(n6094), .A2(n5578), .ZN(n5581) );
  INV_X1 U7043 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5579) );
  OR2_X1 U7044 ( .A1(n4278), .A2(n5579), .ZN(n5580) );
  OAI211_X1 U7045 ( .C1(n5637), .C2(n5582), .A(n5581), .B(n5580), .ZN(n5583)
         );
  INV_X1 U7046 ( .A(n5583), .ZN(n5584) );
  AND2_X1 U7047 ( .A1(n9190), .A2(n5612), .ZN(n5586) );
  AOI21_X1 U7048 ( .B1(n9553), .B2(n4429), .A(n5586), .ZN(n5618) );
  AOI22_X1 U7049 ( .A1(n9553), .A2(n5047), .B1(n4429), .B2(n9190), .ZN(n5587)
         );
  XNOR2_X1 U7050 ( .A(n5587), .B(n5014), .ZN(n5617) );
  XOR2_X1 U7051 ( .A(n5618), .B(n5617), .Z(n8812) );
  AND2_X1 U7052 ( .A1(n8837), .A2(n8812), .ZN(n5592) );
  INV_X1 U7053 ( .A(n8812), .ZN(n5589) );
  INV_X1 U7054 ( .A(n5588), .ZN(n8810) );
  INV_X1 U7055 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7476) );
  INV_X1 U7056 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7472) );
  MUX2_X1 U7057 ( .A(n7476), .B(n7472), .S(n6530), .Z(n5596) );
  INV_X1 U7058 ( .A(SI_26_), .ZN(n5595) );
  NAND2_X1 U7059 ( .A1(n5596), .A2(n5595), .ZN(n5621) );
  INV_X1 U7060 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U7061 ( .A1(n5597), .A2(SI_26_), .ZN(n5598) );
  AND2_X1 U7062 ( .A1(n5621), .A2(n5598), .ZN(n5599) );
  OR2_X1 U7063 ( .A1(n5600), .A2(n5599), .ZN(n5601) );
  NAND2_X1 U7064 ( .A1(n5622), .A2(n5601), .ZN(n7471) );
  NAND2_X1 U7065 ( .A1(n7471), .A2(n5986), .ZN(n5603) );
  OR2_X1 U7066 ( .A1(n5987), .A2(n7472), .ZN(n5602) );
  INV_X1 U7067 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8875) );
  OR2_X2 U7068 ( .A1(n5604), .A2(n8875), .ZN(n5657) );
  NAND2_X1 U7069 ( .A1(n5604), .A2(n8875), .ZN(n5605) );
  NAND2_X1 U7070 ( .A1(n9384), .A2(n5632), .ZN(n5611) );
  INV_X1 U7071 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5608) );
  INV_X1 U7072 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9550) );
  OR2_X1 U7073 ( .A1(n6094), .A2(n9550), .ZN(n5607) );
  INV_X1 U7074 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9616) );
  OR2_X1 U7075 ( .A1(n4279), .A2(n9616), .ZN(n5606) );
  OAI211_X1 U7076 ( .C1(n5637), .C2(n5608), .A(n5607), .B(n5606), .ZN(n5609)
         );
  INV_X1 U7077 ( .A(n5609), .ZN(n5610) );
  NAND2_X2 U7078 ( .A1(n5611), .A2(n5610), .ZN(n9394) );
  AND2_X1 U7079 ( .A1(n9394), .A2(n5612), .ZN(n5613) );
  AOI21_X1 U7080 ( .B1(n9383), .B2(n4429), .A(n5613), .ZN(n5645) );
  NAND2_X1 U7081 ( .A1(n9383), .A2(n5047), .ZN(n5615) );
  NAND2_X1 U7082 ( .A1(n9394), .A2(n4429), .ZN(n5614) );
  NAND2_X1 U7083 ( .A1(n5615), .A2(n5614), .ZN(n5616) );
  XNOR2_X1 U7084 ( .A(n5616), .B(n5014), .ZN(n5647) );
  XOR2_X1 U7085 ( .A(n5645), .B(n5647), .Z(n8872) );
  INV_X1 U7086 ( .A(n5617), .ZN(n5620) );
  INV_X1 U7087 ( .A(n5618), .ZN(n5619) );
  NOR2_X1 U7088 ( .A1(n5620), .A2(n5619), .ZN(n8873) );
  INV_X1 U7089 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7584) );
  INV_X1 U7090 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8684) );
  MUX2_X1 U7091 ( .A(n7584), .B(n8684), .S(n6530), .Z(n5624) );
  INV_X1 U7092 ( .A(SI_27_), .ZN(n5623) );
  NAND2_X1 U7093 ( .A1(n5624), .A2(n5623), .ZN(n5961) );
  INV_X1 U7094 ( .A(n5624), .ZN(n5625) );
  NAND2_X1 U7095 ( .A1(n5625), .A2(SI_27_), .ZN(n5626) );
  AND2_X1 U7096 ( .A1(n5961), .A2(n5626), .ZN(n5627) );
  OR2_X1 U7097 ( .A1(n5628), .A2(n5627), .ZN(n5629) );
  NAND2_X1 U7098 ( .A1(n5966), .A2(n5629), .ZN(n7582) );
  NAND2_X1 U7099 ( .A1(n7582), .A2(n5986), .ZN(n5631) );
  OR2_X1 U7100 ( .A1(n5987), .A2(n8684), .ZN(n5630) );
  XNOR2_X1 U7101 ( .A(n5657), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9361) );
  NAND2_X1 U7102 ( .A1(n9361), .A2(n5632), .ZN(n5640) );
  INV_X1 U7103 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5636) );
  INV_X1 U7104 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8680) );
  OR2_X1 U7105 ( .A1(n6094), .A2(n8680), .ZN(n5635) );
  INV_X1 U7106 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5633) );
  OR2_X1 U7107 ( .A1(n4278), .A2(n5633), .ZN(n5634) );
  OAI211_X1 U7108 ( .C1(n5637), .C2(n5636), .A(n5635), .B(n5634), .ZN(n5638)
         );
  INV_X1 U7109 ( .A(n5638), .ZN(n5639) );
  AND2_X2 U7110 ( .A1(n5640), .A2(n5639), .ZN(n9377) );
  AOI22_X1 U7111 ( .A1(n9543), .A2(n5047), .B1(n4429), .B2(n9189), .ZN(n5641)
         );
  XOR2_X1 U7112 ( .A(n5014), .B(n5641), .Z(n5644) );
  OAI22_X1 U7113 ( .A1(n9363), .A2(n5642), .B1(n9377), .B2(n5016), .ZN(n5643)
         );
  NOR2_X1 U7114 ( .A1(n5644), .A2(n5643), .ZN(n5701) );
  AOI21_X1 U7115 ( .B1(n5644), .B2(n5643), .A(n5701), .ZN(n5729) );
  INV_X1 U7116 ( .A(n5729), .ZN(n5648) );
  INV_X1 U7117 ( .A(n5645), .ZN(n5646) );
  NAND2_X1 U7118 ( .A1(n5647), .A2(n5646), .ZN(n5730) );
  NOR2_X1 U7119 ( .A1(n5648), .A2(n4523), .ZN(n5649) );
  INV_X1 U7120 ( .A(n5731), .ZN(n5700) );
  NAND2_X1 U7121 ( .A1(n5966), .A2(n5961), .ZN(n5650) );
  INV_X1 U7122 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7601) );
  INV_X1 U7123 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7618) );
  MUX2_X1 U7124 ( .A(n7601), .B(n7618), .S(n6530), .Z(n5960) );
  XNOR2_X1 U7125 ( .A(n5960), .B(SI_28_), .ZN(n5963) );
  NAND2_X1 U7126 ( .A1(n7600), .A2(n5986), .ZN(n5652) );
  OR2_X1 U7127 ( .A1(n5987), .A2(n7618), .ZN(n5651) );
  NAND2_X1 U7128 ( .A1(n9354), .A2(n5047), .ZN(n5665) );
  INV_X1 U7129 ( .A(n5657), .ZN(n5654) );
  AND2_X1 U7130 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5653) );
  NAND2_X1 U7131 ( .A1(n5654), .A2(n5653), .ZN(n9327) );
  INV_X1 U7132 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5656) );
  INV_X1 U7133 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5655) );
  OAI21_X1 U7134 ( .B1(n5657), .B2(n5656), .A(n5655), .ZN(n5658) );
  NAND2_X1 U7135 ( .A1(n9327), .A2(n5658), .ZN(n9348) );
  INV_X1 U7136 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9347) );
  INV_X1 U7137 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9612) );
  OR2_X1 U7138 ( .A1(n4279), .A2(n9612), .ZN(n5660) );
  INV_X1 U7139 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9540) );
  OR2_X1 U7140 ( .A1(n5994), .A2(n9540), .ZN(n5659) );
  OAI211_X1 U7141 ( .C1(n5637), .C2(n9347), .A(n5660), .B(n5659), .ZN(n5661)
         );
  INV_X1 U7142 ( .A(n5661), .ZN(n5662) );
  NAND2_X1 U7143 ( .A1(n9368), .A2(n4429), .ZN(n5664) );
  NAND2_X1 U7144 ( .A1(n5665), .A2(n5664), .ZN(n5667) );
  XNOR2_X1 U7145 ( .A(n5667), .B(n5666), .ZN(n5670) );
  NAND2_X1 U7146 ( .A1(n9354), .A2(n4429), .ZN(n5668) );
  OAI21_X1 U7147 ( .B1(n6058), .B2(n5016), .A(n5668), .ZN(n5669) );
  XNOR2_X1 U7148 ( .A(n5670), .B(n5669), .ZN(n5702) );
  INV_X1 U7149 ( .A(n5702), .ZN(n5699) );
  INV_X1 U7150 ( .A(n5671), .ZN(n7368) );
  NAND2_X1 U7151 ( .A1(n7368), .A2(P1_B_REG_SCAN_IN), .ZN(n5672) );
  MUX2_X1 U7152 ( .A(n5672), .B(P1_B_REG_SCAN_IN), .S(n5689), .Z(n5673) );
  NAND2_X1 U7153 ( .A1(n5673), .A2(n5685), .ZN(n9646) );
  NOR4_X1 U7154 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5677) );
  NOR4_X1 U7155 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n5676) );
  NOR4_X1 U7156 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5675) );
  NOR4_X1 U7157 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5674) );
  AND4_X1 U7158 ( .A1(n5677), .A2(n5676), .A3(n5675), .A4(n5674), .ZN(n5683)
         );
  NOR2_X1 U7159 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .ZN(
        n5681) );
  NOR4_X1 U7160 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_30__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5680) );
  NOR4_X1 U7161 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5679) );
  NOR4_X1 U7162 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5678) );
  AND4_X1 U7163 ( .A1(n5681), .A2(n5680), .A3(n5679), .A4(n5678), .ZN(n5682)
         );
  NAND2_X1 U7164 ( .A1(n5683), .A2(n5682), .ZN(n5998) );
  INV_X1 U7165 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5684) );
  OR2_X1 U7166 ( .A1(n5998), .A2(n5684), .ZN(n5687) );
  INV_X1 U7167 ( .A(n5685), .ZN(n7473) );
  NAND2_X1 U7168 ( .A1(n7473), .A2(n7368), .ZN(n9648) );
  INV_X1 U7169 ( .A(n9648), .ZN(n5686) );
  AOI21_X1 U7170 ( .B1(n5999), .B2(n5687), .A(n5686), .ZN(n6882) );
  INV_X1 U7171 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7172 ( .A1(n5999), .A2(n5688), .ZN(n5690) );
  INV_X1 U7173 ( .A(n5689), .ZN(n7301) );
  NAND2_X1 U7174 ( .A1(n7473), .A2(n7301), .ZN(n9649) );
  NAND2_X1 U7175 ( .A1(n5690), .A2(n9649), .ZN(n6880) );
  INV_X1 U7176 ( .A(n6880), .ZN(n6102) );
  NAND2_X1 U7177 ( .A1(n6882), .A2(n6102), .ZN(n5710) );
  NAND2_X1 U7178 ( .A1(n5691), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5693) );
  INV_X1 U7179 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5692) );
  XNOR2_X1 U7180 ( .A(n5693), .B(n5692), .ZN(n6565) );
  AND2_X1 U7181 ( .A1(n6565), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6527) );
  AND2_X1 U7182 ( .A1(n6529), .A2(n6527), .ZN(n9647) );
  INV_X1 U7183 ( .A(n9647), .ZN(n5694) );
  INV_X1 U7184 ( .A(n9184), .ZN(n7084) );
  INV_X1 U7185 ( .A(n6091), .ZN(n9118) );
  AND2_X1 U7186 ( .A1(n7084), .A2(n9118), .ZN(n6061) );
  AND2_X1 U7187 ( .A1(n5695), .A2(n6061), .ZN(n9974) );
  AND2_X1 U7188 ( .A1(n9184), .A2(n6091), .ZN(n8918) );
  OR2_X1 U7189 ( .A1(n9974), .A2(n8918), .ZN(n5696) );
  NOR2_X1 U7190 ( .A1(n5716), .A2(n5696), .ZN(n8895) );
  AND2_X1 U7191 ( .A1(n5702), .A2(n8895), .ZN(n5726) );
  NAND3_X1 U7192 ( .A1(n5702), .A2(n5701), .A3(n8895), .ZN(n5724) );
  NOR2_X2 U7193 ( .A1(n5716), .A2(n5695), .ZN(n8888) );
  INV_X1 U7194 ( .A(n5703), .ZN(n9182) );
  AND2_X1 U7195 ( .A1(n8888), .A2(n9433), .ZN(n8832) );
  OR2_X1 U7196 ( .A1(n9327), .A2(n5704), .ZN(n5709) );
  INV_X1 U7197 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9326) );
  INV_X1 U7198 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6525) );
  OR2_X1 U7199 ( .A1(n5994), .A2(n6525), .ZN(n5706) );
  INV_X1 U7200 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6104) );
  OR2_X1 U7201 ( .A1(n4278), .A2(n6104), .ZN(n5705) );
  OAI211_X1 U7202 ( .C1(n5092), .C2(n9326), .A(n5706), .B(n5705), .ZN(n5707)
         );
  INV_X1 U7203 ( .A(n5707), .ZN(n5708) );
  INV_X1 U7204 ( .A(n9182), .ZN(n7620) );
  AND2_X1 U7205 ( .A1(n8888), .A2(n9431), .ZN(n8813) );
  INV_X1 U7206 ( .A(n8813), .ZN(n8877) );
  INV_X1 U7207 ( .A(n9348), .ZN(n5714) );
  AND2_X1 U7208 ( .A1(n6061), .A2(n8955), .ZN(n9892) );
  NAND2_X1 U7209 ( .A1(n9308), .A2(n9892), .ZN(n6000) );
  NAND2_X1 U7210 ( .A1(n5710), .A2(n6000), .ZN(n5712) );
  NAND2_X1 U7211 ( .A1(n5695), .A2(n8918), .ZN(n5997) );
  AND2_X1 U7212 ( .A1(n5997), .A2(n6529), .ZN(n5711) );
  NAND2_X1 U7213 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  OR2_X1 U7214 ( .A1(n6565), .A2(P1_U3086), .ZN(n9186) );
  INV_X1 U7215 ( .A(n9186), .ZN(n6564) );
  AOI21_X1 U7216 ( .B1(n5713), .B2(P1_STATE_REG_SCAN_IN), .A(n6564), .ZN(n8862) );
  INV_X1 U7217 ( .A(n8862), .ZN(n8880) );
  AOI22_X1 U7218 ( .A1(n5714), .A2(n8880), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5715) );
  OAI21_X1 U7219 ( .B1(n9339), .B2(n8877), .A(n5715), .ZN(n5722) );
  INV_X1 U7220 ( .A(n5716), .ZN(n5718) );
  INV_X1 U7221 ( .A(n8955), .ZN(n9114) );
  NAND2_X1 U7222 ( .A1(n6061), .A2(n9114), .ZN(n6887) );
  INV_X1 U7223 ( .A(n6887), .ZN(n5717) );
  NAND2_X1 U7224 ( .A1(n5718), .A2(n5717), .ZN(n5720) );
  INV_X1 U7225 ( .A(n6000), .ZN(n5719) );
  NAND2_X1 U7226 ( .A1(n9647), .A2(n5719), .ZN(n9501) );
  NOR2_X1 U7227 ( .A1(n4473), .A2(n8883), .ZN(n5721) );
  AOI211_X1 U7228 ( .C1(n8832), .C2(n9189), .A(n5722), .B(n5721), .ZN(n5723)
         );
  AOI21_X1 U7229 ( .B1(n5731), .B2(n5726), .A(n5725), .ZN(n5727) );
  NAND2_X1 U7230 ( .A1(n5728), .A2(n5727), .ZN(P1_U3220) );
  INV_X1 U7231 ( .A(n8880), .ZN(n8893) );
  INV_X1 U7232 ( .A(n9361), .ZN(n5733) );
  AOI22_X1 U7233 ( .A1(n9394), .A2(n8832), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n5732) );
  OAI21_X1 U7234 ( .B1(n8893), .B2(n5733), .A(n5732), .ZN(n5734) );
  AOI21_X1 U7235 ( .B1(n8813), .B2(n9368), .A(n5734), .ZN(n5735) );
  INV_X1 U7236 ( .A(n5736), .ZN(n5737) );
  NAND2_X1 U7237 ( .A1(n5738), .A2(n5737), .ZN(P1_U3214) );
  NOR2_X2 U7238 ( .A1(n5817), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5821) );
  NOR2_X1 U7239 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5742) );
  NOR2_X1 U7240 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5741) );
  INV_X1 U7241 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5800) );
  INV_X1 U7242 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5802) );
  INV_X1 U7243 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5754) );
  INV_X1 U7244 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5794) );
  INV_X1 U7245 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5755) );
  NAND2_X1 U7246 ( .A1(n5794), .A2(n5755), .ZN(n5788) );
  INV_X1 U7247 ( .A(n5788), .ZN(n5745) );
  NOR2_X1 U7248 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5744) );
  NOR2_X2 U7249 ( .A1(n5787), .A2(n4317), .ZN(n5856) );
  INV_X1 U7250 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5746) );
  INV_X1 U7251 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5747) );
  NOR2_X1 U7252 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5752) );
  NOR2_X1 U7253 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5751) );
  NOR2_X1 U7254 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5750) );
  NOR2_X1 U7255 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5749) );
  NAND4_X1 U7256 ( .A1(n5752), .A2(n5751), .A3(n5750), .A4(n5749), .ZN(n5757)
         );
  INV_X1 U7257 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5753) );
  NAND4_X1 U7258 ( .A1(n5755), .A2(n5794), .A3(n5754), .A4(n5753), .ZN(n5756)
         );
  NAND2_X1 U7259 ( .A1(n5776), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5760) );
  XNOR2_X1 U7260 ( .A(n5760), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8226) );
  AND2_X2 U7261 ( .A1(n6804), .A2(n8226), .ZN(n8176) );
  INV_X2 U7262 ( .A(n8176), .ZN(n8137) );
  INV_X1 U7263 ( .A(n5776), .ZN(n5783) );
  INV_X1 U7264 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7265 ( .A1(n5783), .A2(n5780), .ZN(n5767) );
  NAND2_X1 U7266 ( .A1(n5767), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5772) );
  INV_X1 U7267 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U7268 ( .A1(n5772), .A2(n5771), .ZN(n5761) );
  NAND2_X1 U7269 ( .A1(n5761), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5764) );
  INV_X1 U7270 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U7271 ( .A1(n5764), .A2(n5763), .ZN(n5766) );
  NAND2_X1 U7272 ( .A1(n5766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5762) );
  XNOR2_X1 U7273 ( .A(n5762), .B(n4703), .ZN(n7748) );
  INV_X1 U7274 ( .A(n7748), .ZN(n5770) );
  NAND2_X1 U7275 ( .A1(n5766), .A2(n5765), .ZN(n7370) );
  NAND2_X1 U7276 ( .A1(n4319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5768) );
  XNOR2_X1 U7277 ( .A(n5768), .B(n4701), .ZN(n7474) );
  NOR2_X1 U7278 ( .A1(n7370), .A2(n7474), .ZN(n5769) );
  NAND2_X1 U7279 ( .A1(n5770), .A2(n5769), .ZN(n6780) );
  NAND2_X1 U7280 ( .A1(n8137), .A2(n6780), .ZN(n5773) );
  XNOR2_X1 U7281 ( .A(n5772), .B(n5771), .ZN(n6779) );
  NAND2_X1 U7282 ( .A1(n5773), .A2(n6779), .ZN(n5864) );
  NAND2_X1 U7283 ( .A1(n6107), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5778) );
  INV_X1 U7284 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5777) );
  INV_X1 U7285 ( .A(n5779), .ZN(n5781) );
  NAND2_X2 U7286 ( .A1(n8223), .A2(n7583), .ZN(n6155) );
  NAND2_X1 U7287 ( .A1(n5864), .A2(n6443), .ZN(n5785) );
  NAND2_X1 U7288 ( .A1(n5785), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7289 ( .A(n6588), .ZN(n5786) );
  OR2_X2 U7290 ( .A1(n6780), .A2(n5786), .ZN(n8348) );
  INV_X1 U7291 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U7292 ( .A1(n5787), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U7293 ( .A1(n5788), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5789) );
  NAND2_X1 U7294 ( .A1(n5795), .A2(n5789), .ZN(n5791) );
  OR2_X1 U7295 ( .A1(n5791), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7296 ( .A1(n5793), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5790) );
  XNOR2_X1 U7297 ( .A(n5790), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7780) );
  NAND2_X1 U7298 ( .A1(n5791), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5792) );
  AND2_X1 U7299 ( .A1(n5793), .A2(n5792), .ZN(n7796) );
  INV_X1 U7300 ( .A(n7796), .ZN(n6655) );
  NAND2_X1 U7301 ( .A1(n5795), .A2(n5794), .ZN(n5851) );
  OR2_X1 U7302 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  NAND2_X1 U7303 ( .A1(n5851), .A2(n5796), .ZN(n6662) );
  OR2_X1 U7304 ( .A1(n5797), .A2(n6109), .ZN(n5798) );
  XNOR2_X1 U7305 ( .A(n5798), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7843) );
  NAND2_X1 U7306 ( .A1(n5799), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7307 ( .A1(n5804), .A2(n5800), .ZN(n5801) );
  NAND2_X1 U7308 ( .A1(n5801), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5803) );
  XNOR2_X1 U7309 ( .A(n5803), .B(n5802), .ZN(n6632) );
  XNOR2_X1 U7310 ( .A(n5804), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7881) );
  NAND2_X1 U7311 ( .A1(n5806), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5807) );
  XNOR2_X1 U7312 ( .A(n5807), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7895) );
  INV_X1 U7313 ( .A(n7895), .ZN(n6578) );
  MUX2_X1 U7314 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5808), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5810) );
  INV_X1 U7315 ( .A(n5867), .ZN(n5809) );
  INV_X1 U7316 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5866) );
  AND2_X1 U7317 ( .A1(n5866), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7318 ( .A1(n5867), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5812) );
  OAI21_X1 U7319 ( .B1(n6691), .B2(n5811), .A(n5812), .ZN(n6679) );
  INV_X1 U7320 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10097) );
  XNOR2_X1 U7321 ( .A(n6175), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n10015) );
  NAND2_X1 U7322 ( .A1(n10017), .A2(n10015), .ZN(n10016) );
  NAND2_X1 U7323 ( .A1(n10012), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7324 ( .A1(n10016), .A2(n5813), .ZN(n5816) );
  NAND2_X1 U7325 ( .A1(n5814), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5815) );
  INV_X1 U7326 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10101) );
  INV_X1 U7327 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10103) );
  NAND2_X1 U7328 ( .A1(n5817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5819) );
  INV_X1 U7329 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5818) );
  MUX2_X1 U7330 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10103), .S(n6718), .Z(n6700)
         );
  NAND2_X1 U7331 ( .A1(n6718), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U7332 ( .A1(n6704), .A2(n5820), .ZN(n5826) );
  NOR2_X1 U7333 ( .A1(n5821), .A2(n6109), .ZN(n5822) );
  MUX2_X1 U7334 ( .A(n6109), .B(n5822), .S(P2_IR_REG_5__SCAN_IN), .Z(n5824) );
  OR2_X1 U7335 ( .A1(n5824), .A2(n5830), .ZN(n6769) );
  NAND2_X1 U7336 ( .A1(n5826), .A2(n6769), .ZN(n5825) );
  INV_X1 U7337 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10105) );
  OAI21_X1 U7338 ( .B1(n5826), .B2(n6769), .A(n5825), .ZN(n6759) );
  NOR2_X1 U7339 ( .A1(n5830), .A2(n6109), .ZN(n5828) );
  MUX2_X1 U7340 ( .A(n6109), .B(n5828), .S(P2_IR_REG_6__SCAN_IN), .Z(n5832) );
  INV_X1 U7341 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U7342 ( .A1(n5830), .A2(n5829), .ZN(n5836) );
  INV_X1 U7343 ( .A(n5836), .ZN(n5831) );
  INV_X1 U7344 ( .A(n6548), .ZN(n6734) );
  INV_X1 U7345 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U7346 ( .A1(n6734), .A2(P2_REG1_REG_6__SCAN_IN), .B1(n10107), .B2(
        n6548), .ZN(n6722) );
  NAND2_X1 U7347 ( .A1(n5836), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5833) );
  XNOR2_X1 U7348 ( .A(n5833), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7936) );
  INV_X1 U7349 ( .A(n5834), .ZN(n5835) );
  INV_X1 U7350 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10109) );
  NOR2_X1 U7351 ( .A1(n10109), .A2(n7932), .ZN(n7931) );
  OR2_X1 U7352 ( .A1(n5836), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7353 ( .A1(n5840), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5838) );
  INV_X1 U7354 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5837) );
  XNOR2_X1 U7355 ( .A(n5838), .B(n5837), .ZN(n6559) );
  NAND2_X1 U7356 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n6559), .ZN(n5839) );
  OAI21_X1 U7357 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n6559), .A(n5839), .ZN(
        n7914) );
  OAI21_X1 U7358 ( .B1(n5840), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5841) );
  MUX2_X1 U7359 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5841), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5842) );
  AND2_X1 U7360 ( .A1(n5842), .A2(n5806), .ZN(n6968) );
  INV_X1 U7361 ( .A(n6968), .ZN(n6571) );
  INV_X1 U7362 ( .A(n5843), .ZN(n5845) );
  INV_X1 U7363 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10113) );
  INV_X1 U7364 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10115) );
  AOI22_X1 U7365 ( .A1(n7895), .A2(P2_REG1_REG_10__SCAN_IN), .B1(n10115), .B2(
        n6578), .ZN(n7890) );
  NOR2_X1 U7366 ( .A1(n7891), .A2(n7890), .ZN(n7889) );
  NOR2_X1 U7367 ( .A1(n7881), .A2(n5846), .ZN(n5847) );
  INV_X1 U7368 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10117) );
  NAND2_X1 U7369 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n6632), .ZN(n5848) );
  OAI21_X1 U7370 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n6632), .A(n5848), .ZN(
        n7858) );
  INV_X1 U7371 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9724) );
  INV_X1 U7372 ( .A(n7843), .ZN(n6636) );
  NAND2_X1 U7373 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n6662), .ZN(n5850) );
  OAI21_X1 U7374 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n6662), .A(n5850), .ZN(
        n7820) );
  NOR2_X1 U7375 ( .A1(n7821), .A2(n7820), .ZN(n7819) );
  INV_X1 U7376 ( .A(n5853), .ZN(n5854) );
  NAND2_X1 U7377 ( .A1(n5851), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5852) );
  XNOR2_X1 U7378 ( .A(n5852), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8368) );
  INV_X1 U7379 ( .A(n8368), .ZN(n6667) );
  INV_X1 U7380 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8351) );
  XNOR2_X1 U7381 ( .A(n6655), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n7802) );
  INV_X1 U7382 ( .A(n5856), .ZN(n5857) );
  NAND2_X1 U7383 ( .A1(n5857), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5858) );
  MUX2_X1 U7384 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5858), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n5860) );
  NAND2_X1 U7385 ( .A1(n5860), .A2(n5859), .ZN(n7757) );
  NAND2_X1 U7386 ( .A1(n7757), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5861) );
  OAI21_X1 U7387 ( .B1(n7757), .B2(P2_REG1_REG_18__SCAN_IN), .A(n5861), .ZN(
        n7761) );
  NAND2_X1 U7388 ( .A1(n7762), .A2(n5861), .ZN(n5863) );
  NAND2_X1 U7389 ( .A1(n5859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5862) );
  XNOR2_X1 U7390 ( .A(n8221), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n5946) );
  XNOR2_X1 U7391 ( .A(n5863), .B(n5946), .ZN(n5865) );
  NAND2_X1 U7392 ( .A1(n5864), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5951) );
  OR2_X1 U7393 ( .A1(n5951), .A2(n8223), .ZN(n6642) );
  INV_X1 U7394 ( .A(n7583), .ZN(n8224) );
  INV_X1 U7395 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7924) );
  AND2_X1 U7396 ( .A1(n5866), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7397 ( .A1(n5867), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5869) );
  OAI21_X1 U7398 ( .B1(n6691), .B2(n5868), .A(n5869), .ZN(n6676) );
  INV_X1 U7399 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U7400 ( .A1(n6678), .A2(n5869), .ZN(n10001) );
  XNOR2_X1 U7401 ( .A(n6175), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U7402 ( .A1(n10001), .A2(n10002), .ZN(n10000) );
  NAND2_X1 U7403 ( .A1(n10012), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U7404 ( .A1(n10000), .A2(n5870), .ZN(n5871) );
  NAND2_X1 U7405 ( .A1(n5871), .A2(n6538), .ZN(n6706) );
  INV_X1 U7406 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7204) );
  INV_X1 U7407 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7195) );
  MUX2_X1 U7408 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7195), .S(n6718), .Z(n6705)
         );
  NAND2_X1 U7409 ( .A1(n6718), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U7410 ( .A1(n6709), .A2(n5872), .ZN(n5874) );
  INV_X1 U7411 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U7412 ( .A1(P2_REG2_REG_6__SCAN_IN), .A2(n6548), .ZN(n5876) );
  OAI21_X1 U7413 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n6548), .A(n5876), .ZN(
        n6730) );
  INV_X1 U7414 ( .A(n5876), .ZN(n5877) );
  NAND2_X1 U7415 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n6559), .ZN(n5880) );
  OAI21_X1 U7416 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n6559), .A(n5880), .ZN(
        n7904) );
  NOR2_X1 U7417 ( .A1(n7905), .A2(n7904), .ZN(n7903) );
  AND2_X1 U7418 ( .A1(n6559), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5881) );
  INV_X1 U7419 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6963) );
  INV_X1 U7420 ( .A(n5883), .ZN(n5884) );
  INV_X1 U7421 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5885) );
  AOI22_X1 U7422 ( .A1(n7895), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n5885), .B2(
        n6578), .ZN(n7884) );
  NOR2_X1 U7423 ( .A1(n7881), .A2(n5886), .ZN(n5887) );
  INV_X1 U7424 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7867) );
  NOR2_X1 U7425 ( .A1(n7867), .A2(n7866), .ZN(n7865) );
  NAND2_X1 U7426 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n6632), .ZN(n5888) );
  OAI21_X1 U7427 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n6632), .A(n5888), .ZN(
        n7847) );
  NOR2_X1 U7428 ( .A1(n7843), .A2(n5889), .ZN(n5890) );
  INV_X1 U7429 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U7430 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n6662), .ZN(n5891) );
  OAI21_X1 U7431 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n6662), .A(n5891), .ZN(
        n7810) );
  AND2_X1 U7432 ( .A1(n6662), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7433 ( .A1(n5894), .A2(n6667), .ZN(n5893) );
  INV_X1 U7434 ( .A(n5893), .ZN(n5895) );
  INV_X1 U7435 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8363) );
  NOR2_X1 U7436 ( .A1(n8363), .A2(n8364), .ZN(n8362) );
  INV_X1 U7437 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5900) );
  AOI22_X1 U7438 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n7796), .B1(n6655), .B2(
        n5900), .ZN(n7789) );
  INV_X1 U7439 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U7440 ( .A1(n7757), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5898) );
  OAI21_X1 U7441 ( .B1(n7757), .B2(P2_REG2_REG_18__SCAN_IN), .A(n5898), .ZN(
        n7752) );
  INV_X1 U7442 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8692) );
  MUX2_X1 U7443 ( .A(n8692), .B(P2_REG2_REG_19__SCAN_IN), .S(n8221), .Z(n5945)
         );
  XNOR2_X1 U7444 ( .A(n5899), .B(n5945), .ZN(n5956) );
  MUX2_X1 U7445 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n7583), .Z(n5941) );
  XNOR2_X1 U7446 ( .A(n5941), .B(n7780), .ZN(n7782) );
  INV_X1 U7447 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7671) );
  MUX2_X1 U7448 ( .A(n5900), .B(n7671), .S(n7583), .Z(n5940) );
  NOR2_X1 U7449 ( .A1(n5940), .A2(n7796), .ZN(n7791) );
  MUX2_X1 U7450 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n7583), .Z(n5936) );
  NOR2_X1 U7451 ( .A1(n5936), .A2(n6667), .ZN(n5939) );
  MUX2_X1 U7452 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n7583), .Z(n5932) );
  NOR2_X1 U7453 ( .A1(n5932), .A2(n6662), .ZN(n5935) );
  MUX2_X1 U7454 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n7583), .Z(n5928) );
  NOR2_X1 U7455 ( .A1(n5928), .A2(n6636), .ZN(n5931) );
  MUX2_X1 U7456 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n7583), .Z(n5924) );
  NOR2_X1 U7457 ( .A1(n5924), .A2(n6632), .ZN(n5927) );
  MUX2_X1 U7458 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n7583), .Z(n5921) );
  INV_X1 U7459 ( .A(n7881), .ZN(n6583) );
  NOR2_X1 U7460 ( .A1(n5921), .A2(n6583), .ZN(n5923) );
  MUX2_X1 U7461 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n7583), .Z(n5918) );
  NOR2_X1 U7462 ( .A1(n5918), .A2(n6578), .ZN(n5920) );
  MUX2_X1 U7463 ( .A(n6963), .B(n10113), .S(n7583), .Z(n5916) );
  NOR2_X1 U7464 ( .A1(n5916), .A2(n6968), .ZN(n6969) );
  INV_X1 U7465 ( .A(n6969), .ZN(n5917) );
  MUX2_X1 U7466 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n7583), .Z(n5914) );
  OR2_X1 U7467 ( .A1(n5914), .A2(n6559), .ZN(n5915) );
  MUX2_X1 U7468 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n7583), .Z(n5911) );
  INV_X1 U7469 ( .A(n5911), .ZN(n5912) );
  MUX2_X1 U7470 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n7583), .Z(n5909) );
  INV_X1 U7471 ( .A(n5909), .ZN(n5910) );
  MUX2_X1 U7472 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n7583), .Z(n5908) );
  INV_X1 U7473 ( .A(n6538), .ZN(n6752) );
  MUX2_X1 U7474 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n7583), .Z(n5906) );
  INV_X1 U7475 ( .A(n5906), .ZN(n5907) );
  MUX2_X1 U7476 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n7583), .Z(n5904) );
  INV_X1 U7477 ( .A(n5904), .ZN(n5905) );
  INV_X1 U7478 ( .A(n6691), .ZN(n5903) );
  INV_X1 U7479 ( .A(n5901), .ZN(n5902) );
  XNOR2_X1 U7480 ( .A(n5901), .B(n5903), .ZN(n6682) );
  INV_X1 U7481 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6935) );
  INV_X1 U7482 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10095) );
  MUX2_X1 U7483 ( .A(n6935), .B(n10095), .S(n7583), .Z(n6643) );
  NAND2_X1 U7484 ( .A1(n6643), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6681) );
  NAND2_X1 U7485 ( .A1(n6682), .A2(n6681), .ZN(n6680) );
  OAI21_X1 U7486 ( .B1(n5903), .B2(n5902), .A(n6680), .ZN(n10009) );
  XNOR2_X1 U7487 ( .A(n5904), .B(n6175), .ZN(n10008) );
  NAND2_X1 U7488 ( .A1(n10009), .A2(n10008), .ZN(n10007) );
  OAI21_X1 U7489 ( .B1(n6175), .B2(n5905), .A(n10007), .ZN(n6738) );
  XNOR2_X1 U7490 ( .A(n5906), .B(n6538), .ZN(n6739) );
  NOR2_X1 U7491 ( .A1(n6738), .A2(n6739), .ZN(n6737) );
  XOR2_X1 U7492 ( .A(n6718), .B(n5908), .Z(n6698) );
  XNOR2_X1 U7493 ( .A(n5909), .B(n4582), .ZN(n6756) );
  OAI21_X1 U7494 ( .B1(n4582), .B2(n5910), .A(n6755), .ZN(n6720) );
  XNOR2_X1 U7495 ( .A(n5911), .B(n6548), .ZN(n6721) );
  NOR2_X1 U7496 ( .A1(n6720), .A2(n6721), .ZN(n6719) );
  MUX2_X1 U7497 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n7583), .Z(n5913) );
  XOR2_X1 U7498 ( .A(n7936), .B(n5913), .Z(n7926) );
  INV_X1 U7499 ( .A(n6559), .ZN(n7919) );
  XNOR2_X1 U7500 ( .A(n5914), .B(n7919), .ZN(n7907) );
  AND2_X1 U7501 ( .A1(n5916), .A2(n6968), .ZN(n6970) );
  AOI21_X1 U7502 ( .B1(n5917), .B2(n6971), .A(n6970), .ZN(n7898) );
  AOI21_X1 U7503 ( .B1(n5918), .B2(n6578), .A(n5920), .ZN(n5919) );
  INV_X1 U7504 ( .A(n5919), .ZN(n7897) );
  NOR2_X1 U7505 ( .A1(n7898), .A2(n7897), .ZN(n7896) );
  AOI21_X1 U7506 ( .B1(n5921), .B2(n6583), .A(n5923), .ZN(n5922) );
  INV_X1 U7507 ( .A(n5922), .ZN(n7870) );
  INV_X1 U7508 ( .A(n6632), .ZN(n7862) );
  INV_X1 U7509 ( .A(n5924), .ZN(n5926) );
  INV_X1 U7510 ( .A(n5927), .ZN(n5925) );
  OAI21_X1 U7511 ( .B1(n7862), .B2(n5926), .A(n5925), .ZN(n7852) );
  NOR2_X1 U7512 ( .A1(n5927), .A2(n7850), .ZN(n7832) );
  INV_X1 U7513 ( .A(n5928), .ZN(n5930) );
  INV_X1 U7514 ( .A(n5931), .ZN(n5929) );
  OAI21_X1 U7515 ( .B1(n7843), .B2(n5930), .A(n5929), .ZN(n7833) );
  NOR2_X1 U7516 ( .A1(n7832), .A2(n7833), .ZN(n7831) );
  INV_X1 U7517 ( .A(n6662), .ZN(n7825) );
  INV_X1 U7518 ( .A(n5932), .ZN(n5934) );
  INV_X1 U7519 ( .A(n5935), .ZN(n5933) );
  OAI21_X1 U7520 ( .B1(n7825), .B2(n5934), .A(n5933), .ZN(n7814) );
  INV_X1 U7521 ( .A(n5936), .ZN(n5938) );
  INV_X1 U7522 ( .A(n5939), .ZN(n5937) );
  OAI21_X1 U7523 ( .B1(n8368), .B2(n5938), .A(n5937), .ZN(n8356) );
  NOR2_X1 U7524 ( .A1(n5939), .A2(n8354), .ZN(n7795) );
  NAND2_X1 U7525 ( .A1(n5940), .A2(n7796), .ZN(n7793) );
  OAI21_X1 U7526 ( .B1(n7791), .B2(n7795), .A(n7793), .ZN(n7783) );
  NAND2_X1 U7527 ( .A1(n7782), .A2(n7783), .ZN(n7781) );
  OAI21_X1 U7528 ( .B1(n5941), .B2(n4364), .A(n7781), .ZN(n5944) );
  INV_X1 U7529 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n7679) );
  INV_X1 U7530 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n5942) );
  MUX2_X1 U7531 ( .A(n7679), .B(n5942), .S(n7583), .Z(n5943) );
  NAND2_X1 U7532 ( .A1(n5944), .A2(n5943), .ZN(n7755) );
  NOR2_X1 U7533 ( .A1(n5944), .A2(n5943), .ZN(n7754) );
  AOI21_X1 U7534 ( .B1(n7757), .B2(n7755), .A(n7754), .ZN(n5948) );
  MUX2_X1 U7535 ( .A(n5946), .B(n5945), .S(n8224), .Z(n5947) );
  INV_X1 U7536 ( .A(n8223), .ZN(n6441) );
  OR2_X1 U7537 ( .A1(n8348), .A2(n6441), .ZN(n8357) );
  INV_X1 U7538 ( .A(n6779), .ZN(n7130) );
  NOR2_X1 U7539 ( .A1(n6780), .A2(n7130), .ZN(n5949) );
  INV_X1 U7540 ( .A(n10021), .ZN(n6766) );
  NAND2_X1 U7541 ( .A1(n6766), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U7542 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8240) );
  INV_X1 U7543 ( .A(n5951), .ZN(n5952) );
  MUX2_X1 U7544 ( .A(P2_U3893), .B(n5952), .S(n8223), .Z(n5953) );
  AND2_X1 U7545 ( .A1(n5953), .A2(n6443), .ZN(n8369) );
  INV_X1 U7546 ( .A(n8221), .ZN(n6479) );
  NAND2_X1 U7547 ( .A1(n4839), .A2(n5958), .ZN(P2_U3201) );
  INV_X1 U7548 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6003) );
  INV_X1 U7549 ( .A(SI_28_), .ZN(n5959) );
  NAND2_X1 U7550 ( .A1(n5960), .A2(n5959), .ZN(n5962) );
  AND2_X1 U7551 ( .A1(n5961), .A2(n5962), .ZN(n5965) );
  INV_X1 U7552 ( .A(n5962), .ZN(n5964) );
  INV_X1 U7553 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7723) );
  INV_X1 U7554 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7992) );
  MUX2_X1 U7555 ( .A(n7723), .B(n7992), .S(n6530), .Z(n5968) );
  INV_X1 U7556 ( .A(SI_29_), .ZN(n5967) );
  INV_X1 U7557 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7997) );
  INV_X1 U7558 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9656) );
  MUX2_X1 U7559 ( .A(n7997), .B(n9656), .S(n6530), .Z(n5973) );
  INV_X1 U7560 ( .A(SI_30_), .ZN(n5972) );
  NAND2_X1 U7561 ( .A1(n5973), .A2(n5972), .ZN(n5976) );
  INV_X1 U7562 ( .A(n5973), .ZN(n5974) );
  NAND2_X1 U7563 ( .A1(n5974), .A2(SI_30_), .ZN(n5975) );
  NAND2_X1 U7564 ( .A1(n5976), .A2(n5975), .ZN(n5981) );
  INV_X1 U7565 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8000) );
  INV_X1 U7566 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9650) );
  MUX2_X1 U7567 ( .A(n8000), .B(n9650), .S(n6530), .Z(n5977) );
  XNOR2_X1 U7568 ( .A(n5977), .B(SI_31_), .ZN(n5978) );
  NOR2_X1 U7569 ( .A1(n5987), .A2(n9650), .ZN(n5980) );
  INV_X1 U7570 ( .A(n9606), .ZN(n9105) );
  NAND2_X1 U7571 ( .A1(n7996), .A2(n5986), .ZN(n5984) );
  OR2_X1 U7572 ( .A1(n5987), .A2(n9656), .ZN(n5983) );
  NAND2_X1 U7573 ( .A1(n7722), .A2(n5986), .ZN(n5989) );
  OR2_X1 U7574 ( .A1(n5987), .A2(n7992), .ZN(n5988) );
  NOR2_X1 U7575 ( .A1(n6986), .A2(n6989), .ZN(n9894) );
  NAND2_X1 U7576 ( .A1(n9894), .A2(n9921), .ZN(n9893) );
  NAND2_X1 U7577 ( .A1(n7293), .A2(n7546), .ZN(n7398) );
  INV_X1 U7578 ( .A(n9011), .ZN(n7721) );
  INV_X1 U7579 ( .A(n9520), .ZN(n9640) );
  INV_X1 U7580 ( .A(n9500), .ZN(n9636) );
  INV_X1 U7581 ( .A(n9553), .ZN(n9401) );
  XNOR2_X1 U7582 ( .A(n9105), .B(n9318), .ZN(n5990) );
  INV_X1 U7583 ( .A(n9892), .ZN(n9909) );
  INV_X1 U7584 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n5991) );
  OR2_X1 U7585 ( .A1(n5092), .A2(n5991), .ZN(n5993) );
  INV_X1 U7586 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9604) );
  OR2_X1 U7587 ( .A1(n4278), .A2(n9604), .ZN(n5992) );
  OAI211_X1 U7588 ( .C1(n5994), .C2(n6003), .A(n5993), .B(n5992), .ZN(n8916)
         );
  INV_X1 U7589 ( .A(n9728), .ZN(n6622) );
  NAND2_X1 U7590 ( .A1(n6622), .A2(P1_B_REG_SCAN_IN), .ZN(n5996) );
  AND2_X1 U7591 ( .A1(n9431), .A2(n5996), .ZN(n6099) );
  AND2_X1 U7592 ( .A1(n8916), .A2(n6099), .ZN(n9315) );
  NOR2_X1 U7593 ( .A1(n9314), .A2(n9315), .ZN(n9603) );
  AND2_X1 U7594 ( .A1(n9647), .A2(n5997), .ZN(n6881) );
  OAI21_X1 U7595 ( .B1(n9646), .B2(P1_D_REG_1__SCAN_IN), .A(n9648), .ZN(n6002)
         );
  NAND2_X1 U7596 ( .A1(n5999), .A2(n5998), .ZN(n6001) );
  NAND4_X1 U7597 ( .A1(n6881), .A2(n6002), .A3(n6001), .A4(n6000), .ZN(n6103)
         );
  MUX2_X1 U7598 ( .A(n6003), .B(n9603), .S(n9998), .Z(n6006) );
  NAND2_X1 U7599 ( .A1(n9998), .A2(n9974), .ZN(n9602) );
  NAND2_X1 U7600 ( .A1(n6006), .A2(n6005), .ZN(P1_U3553) );
  NAND2_X1 U7601 ( .A1(n9212), .A2(n6904), .ZN(n6901) );
  NAND2_X1 U7602 ( .A1(n6908), .A2(n6901), .ZN(n6009) );
  NAND2_X1 U7603 ( .A1(n6009), .A2(n6008), .ZN(n6978) );
  NAND2_X1 U7604 ( .A1(n6011), .A2(n6989), .ZN(n6065) );
  INV_X1 U7605 ( .A(n6011), .ZN(n6010) );
  NAND2_X1 U7606 ( .A1(n6010), .A2(n9917), .ZN(n9119) );
  NAND2_X1 U7607 ( .A1(n6065), .A2(n9119), .ZN(n6977) );
  NAND2_X1 U7608 ( .A1(n6011), .A2(n9917), .ZN(n9888) );
  AND4_X1 U7609 ( .A1(n6015), .A2(n6014), .A3(n6013), .A4(n6012), .ZN(n6773)
         );
  NAND2_X1 U7610 ( .A1(n6773), .A2(n9921), .ZN(n6016) );
  AND2_X1 U7611 ( .A1(n9888), .A2(n6016), .ZN(n6018) );
  NAND2_X1 U7612 ( .A1(n7209), .A2(n9927), .ZN(n8965) );
  NAND2_X1 U7613 ( .A1(n7209), .A2(n6943), .ZN(n6019) );
  XNOR2_X1 U7614 ( .A(n9207), .B(n9934), .ZN(n9872) );
  NAND2_X1 U7615 ( .A1(n9871), .A2(n9872), .ZN(n6021) );
  INV_X1 U7616 ( .A(n9207), .ZN(n7070) );
  NAND2_X1 U7617 ( .A1(n7070), .A2(n9934), .ZN(n6020) );
  NAND2_X1 U7618 ( .A1(n6021), .A2(n6020), .ZN(n7072) );
  NAND2_X1 U7619 ( .A1(n7230), .A2(n7363), .ZN(n8969) );
  INV_X1 U7620 ( .A(n7230), .ZN(n9206) );
  NAND2_X1 U7621 ( .A1(n9206), .A2(n9940), .ZN(n8971) );
  NAND2_X1 U7622 ( .A1(n8969), .A2(n8971), .ZN(n7073) );
  NAND2_X1 U7623 ( .A1(n7230), .A2(n9940), .ZN(n6022) );
  XNOR2_X1 U7624 ( .A(n9205), .B(n9946), .ZN(n9847) );
  NAND2_X1 U7625 ( .A1(n9953), .A2(n9204), .ZN(n8977) );
  INV_X1 U7626 ( .A(n9204), .ZN(n7558) );
  NAND2_X1 U7627 ( .A1(n7558), .A2(n7457), .ZN(n8982) );
  NAND2_X1 U7628 ( .A1(n8977), .A2(n8982), .ZN(n7237) );
  NAND2_X1 U7629 ( .A1(n7235), .A2(n7237), .ZN(n6024) );
  NAND2_X1 U7630 ( .A1(n9953), .A2(n7558), .ZN(n6023) );
  NAND2_X1 U7631 ( .A1(n6024), .A2(n6023), .ZN(n7321) );
  OR2_X1 U7632 ( .A1(n7287), .A2(n9959), .ZN(n8990) );
  NAND2_X1 U7633 ( .A1(n9959), .A2(n7287), .ZN(n8985) );
  NAND2_X1 U7634 ( .A1(n8990), .A2(n8985), .ZN(n7327) );
  NAND2_X1 U7635 ( .A1(n7321), .A2(n7327), .ZN(n6026) );
  OR2_X1 U7636 ( .A1(n9959), .A2(n9203), .ZN(n6025) );
  NAND2_X1 U7637 ( .A1(n6026), .A2(n6025), .ZN(n7291) );
  OR2_X1 U7638 ( .A1(n7574), .A2(n7540), .ZN(n9124) );
  NAND2_X1 U7639 ( .A1(n7574), .A2(n7540), .ZN(n8993) );
  NAND2_X1 U7640 ( .A1(n9124), .A2(n8993), .ZN(n8931) );
  NAND2_X1 U7641 ( .A1(n7291), .A2(n8931), .ZN(n6028) );
  OR2_X1 U7642 ( .A1(n7574), .A2(n9202), .ZN(n6027) );
  NAND2_X1 U7643 ( .A1(n9841), .A2(n9201), .ZN(n8997) );
  NAND2_X1 U7644 ( .A1(n8995), .A2(n8997), .ZN(n8921) );
  OR2_X1 U7645 ( .A1(n7523), .A2(n7539), .ZN(n8998) );
  NAND2_X1 U7646 ( .A1(n7523), .A2(n7539), .ZN(n9134) );
  NAND2_X1 U7647 ( .A1(n8998), .A2(n9134), .ZN(n7396) );
  NAND2_X1 U7648 ( .A1(n7397), .A2(n7396), .ZN(n6030) );
  NAND2_X1 U7649 ( .A1(n7523), .A2(n9200), .ZN(n6029) );
  AND2_X1 U7650 ( .A1(n9005), .A2(n9199), .ZN(n6031) );
  OR2_X1 U7651 ( .A1(n9005), .A2(n9199), .ZN(n6032) );
  NAND2_X1 U7652 ( .A1(n9973), .A2(n9198), .ZN(n6033) );
  NAND2_X1 U7653 ( .A1(n7647), .A2(n6033), .ZN(n6035) );
  OR2_X1 U7654 ( .A1(n9973), .A2(n9198), .ZN(n6034) );
  NAND2_X1 U7655 ( .A1(n6035), .A2(n6034), .ZN(n7657) );
  NOR2_X1 U7656 ( .A1(n9011), .A2(n9197), .ZN(n6037) );
  NAND2_X1 U7657 ( .A1(n9011), .A2(n9197), .ZN(n6036) );
  OAI21_X1 U7658 ( .B1(n7657), .B2(n6037), .A(n6036), .ZN(n7699) );
  NAND2_X1 U7659 ( .A1(n8825), .A2(n7665), .ZN(n9143) );
  NAND2_X1 U7660 ( .A1(n9141), .A2(n9143), .ZN(n8940) );
  NAND2_X1 U7661 ( .A1(n7699), .A2(n8940), .ZN(n6039) );
  NAND2_X1 U7662 ( .A1(n8825), .A2(n9196), .ZN(n6038) );
  NAND2_X1 U7663 ( .A1(n6039), .A2(n6038), .ZN(n7738) );
  AND2_X1 U7664 ( .A1(n9594), .A2(n9195), .ZN(n9029) );
  OR2_X1 U7665 ( .A1(n9594), .A2(n9195), .ZN(n9027) );
  NOR2_X1 U7666 ( .A1(n9520), .A2(n9194), .ZN(n6041) );
  NAND2_X1 U7667 ( .A1(n9520), .A2(n9194), .ZN(n6040) );
  OAI21_X1 U7668 ( .B1(n9509), .B2(n6041), .A(n6040), .ZN(n9496) );
  OR2_X1 U7669 ( .A1(n9500), .A2(n9193), .ZN(n6042) );
  NAND2_X1 U7670 ( .A1(n9496), .A2(n6042), .ZN(n6044) );
  NAND2_X1 U7671 ( .A1(n9500), .A2(n9193), .ZN(n6043) );
  NAND2_X1 U7672 ( .A1(n6044), .A2(n6043), .ZN(n9477) );
  OR2_X1 U7673 ( .A1(n9484), .A2(n9192), .ZN(n6045) );
  NOR2_X1 U7674 ( .A1(n9574), .A2(n9191), .ZN(n6046) );
  AND2_X1 U7675 ( .A1(n9450), .A2(n9434), .ZN(n6047) );
  NAND2_X1 U7676 ( .A1(n9563), .A2(n9065), .ZN(n6048) );
  OAI22_X1 U7677 ( .A1(n9412), .A2(n6049), .B1(n9432), .B2(n9416), .ZN(n9390)
         );
  NOR2_X1 U7678 ( .A1(n9553), .A2(n9190), .ZN(n6051) );
  NAND2_X1 U7679 ( .A1(n9553), .A2(n9190), .ZN(n6050) );
  OAI21_X1 U7680 ( .B1(n9390), .B2(n6051), .A(n6050), .ZN(n9373) );
  OR2_X1 U7681 ( .A1(n9383), .A2(n9394), .ZN(n6052) );
  NAND2_X1 U7682 ( .A1(n9373), .A2(n6052), .ZN(n6054) );
  NAND2_X1 U7683 ( .A1(n9383), .A2(n9394), .ZN(n6053) );
  NAND2_X1 U7684 ( .A1(n6054), .A2(n6053), .ZN(n9357) );
  INV_X1 U7685 ( .A(n9357), .ZN(n6056) );
  NAND2_X1 U7686 ( .A1(n9543), .A2(n9377), .ZN(n9085) );
  INV_X1 U7687 ( .A(n9366), .ZN(n6055) );
  OR2_X1 U7688 ( .A1(n9543), .A2(n9189), .ZN(n6057) );
  NAND2_X1 U7689 ( .A1(n9354), .A2(n6058), .ZN(n9095) );
  NAND2_X1 U7690 ( .A1(n6105), .A2(n9339), .ZN(n9098) );
  OR2_X1 U7691 ( .A1(n9180), .A2(n9179), .ZN(n6062) );
  INV_X1 U7692 ( .A(n6061), .ZN(n6660) );
  NAND2_X1 U7693 ( .A1(n6062), .A2(n6660), .ZN(n6885) );
  AND2_X1 U7694 ( .A1(n9180), .A2(n5695), .ZN(n6063) );
  OR2_X1 U7695 ( .A1(n6885), .A2(n6063), .ZN(n9851) );
  NAND2_X1 U7696 ( .A1(n9308), .A2(n7084), .ZN(n9111) );
  OR2_X1 U7697 ( .A1(n9111), .A2(n9114), .ZN(n9977) );
  INV_X1 U7698 ( .A(n6908), .ZN(n8923) );
  NOR2_X1 U7699 ( .A1(n9212), .A2(n6891), .ZN(n6907) );
  INV_X1 U7700 ( .A(n6892), .ZN(n9210) );
  NAND2_X1 U7701 ( .A1(n6979), .A2(n6065), .ZN(n6066) );
  NAND2_X1 U7702 ( .A1(n6066), .A2(n9119), .ZN(n9879) );
  AND2_X1 U7703 ( .A1(n6067), .A2(n9921), .ZN(n9117) );
  NAND2_X1 U7704 ( .A1(n6773), .A2(n9885), .ZN(n6068) );
  INV_X1 U7705 ( .A(n8965), .ZN(n6069) );
  NAND2_X1 U7706 ( .A1(n7070), .A2(n9870), .ZN(n8966) );
  AND2_X1 U7707 ( .A1(n8990), .A2(n8977), .ZN(n8983) );
  INV_X1 U7708 ( .A(n9946), .ZN(n9857) );
  NAND2_X1 U7709 ( .A1(n7069), .A2(n9857), .ZN(n7236) );
  NAND2_X1 U7710 ( .A1(n8982), .A2(n7236), .ZN(n8979) );
  INV_X1 U7711 ( .A(n8985), .ZN(n8991) );
  AOI21_X1 U7712 ( .B1(n8983), .B2(n8979), .A(n8991), .ZN(n8928) );
  NAND2_X1 U7713 ( .A1(n8928), .A2(n8969), .ZN(n6071) );
  NAND2_X1 U7714 ( .A1(n9205), .A2(n9946), .ZN(n8976) );
  AND2_X1 U7715 ( .A1(n8971), .A2(n8976), .ZN(n6072) );
  NAND2_X1 U7716 ( .A1(n8983), .A2(n6072), .ZN(n8926) );
  NAND2_X1 U7717 ( .A1(n8928), .A2(n8926), .ZN(n9125) );
  INV_X1 U7718 ( .A(n7542), .ZN(n6073) );
  NAND2_X1 U7719 ( .A1(n6073), .A2(n4507), .ZN(n7404) );
  NAND2_X1 U7720 ( .A1(n7404), .A2(n9131), .ZN(n6074) );
  NAND2_X1 U7721 ( .A1(n6074), .A2(n9134), .ZN(n7410) );
  XNOR2_X1 U7722 ( .A(n9005), .B(n9199), .ZN(n8935) );
  NAND2_X1 U7723 ( .A1(n7410), .A2(n8935), .ZN(n6075) );
  INV_X1 U7724 ( .A(n9199), .ZN(n9004) );
  NAND2_X1 U7725 ( .A1(n9005), .A2(n9004), .ZN(n9133) );
  NAND2_X1 U7726 ( .A1(n6075), .A2(n9133), .ZN(n7643) );
  NAND2_X1 U7727 ( .A1(n9973), .A2(n6076), .ZN(n9014) );
  NAND2_X1 U7728 ( .A1(n9137), .A2(n9014), .ZN(n8938) );
  INV_X1 U7729 ( .A(n8938), .ZN(n6077) );
  INV_X1 U7730 ( .A(n9197), .ZN(n9010) );
  XNOR2_X1 U7731 ( .A(n9011), .B(n9010), .ZN(n7662) );
  NAND2_X1 U7732 ( .A1(n9011), .A2(n9010), .ZN(n8962) );
  INV_X1 U7733 ( .A(n9195), .ZN(n6079) );
  OR2_X1 U7734 ( .A1(n9594), .A2(n6079), .ZN(n9510) );
  NAND2_X1 U7735 ( .A1(n9594), .A2(n6079), .ZN(n9147) );
  INV_X1 U7736 ( .A(n9194), .ZN(n9036) );
  OR2_X1 U7737 ( .A1(n9520), .A2(n9036), .ZN(n9151) );
  NAND2_X1 U7738 ( .A1(n9520), .A2(n9036), .ZN(n9148) );
  NAND2_X1 U7739 ( .A1(n9151), .A2(n9148), .ZN(n9512) );
  INV_X1 U7740 ( .A(n9510), .ZN(n6080) );
  NOR2_X1 U7741 ( .A1(n9512), .A2(n6080), .ZN(n6081) );
  INV_X1 U7742 ( .A(n9193), .ZN(n6082) );
  OR2_X1 U7743 ( .A1(n9500), .A2(n6082), .ZN(n9152) );
  NAND2_X1 U7744 ( .A1(n9500), .A2(n6082), .ZN(n9156) );
  NAND2_X1 U7745 ( .A1(n9491), .A2(n9495), .ZN(n6083) );
  NAND2_X1 U7746 ( .A1(n6083), .A2(n9156), .ZN(n8903) );
  INV_X1 U7747 ( .A(n8903), .ZN(n6084) );
  AND2_X1 U7748 ( .A1(n9484), .A2(n9468), .ZN(n8960) );
  INV_X1 U7749 ( .A(n9191), .ZN(n9448) );
  OR2_X1 U7750 ( .A1(n9574), .A2(n9448), .ZN(n9057) );
  NAND2_X1 U7751 ( .A1(n9574), .A2(n9448), .ZN(n9048) );
  NAND2_X1 U7752 ( .A1(n9057), .A2(n9048), .ZN(n9463) );
  AND2_X1 U7753 ( .A1(n6085), .A2(n9192), .ZN(n8959) );
  NOR2_X1 U7754 ( .A1(n9463), .A2(n8959), .ZN(n6086) );
  XNOR2_X1 U7755 ( .A(n9450), .B(n9434), .ZN(n9441) );
  INV_X1 U7756 ( .A(n9434), .ZN(n9466) );
  NAND2_X1 U7757 ( .A1(n9450), .A2(n9466), .ZN(n9428) );
  NAND2_X1 U7758 ( .A1(n9443), .A2(n9428), .ZN(n6087) );
  NAND2_X1 U7759 ( .A1(n9426), .A2(n9065), .ZN(n8899) );
  NAND2_X1 U7760 ( .A1(n9563), .A2(n9447), .ZN(n9059) );
  INV_X1 U7761 ( .A(n9432), .ZN(n8784) );
  NAND2_X1 U7762 ( .A1(n9416), .A2(n8784), .ZN(n9067) );
  NAND2_X1 U7763 ( .A1(n9068), .A2(n9067), .ZN(n9406) );
  OR2_X1 U7764 ( .A1(n9553), .A2(n9409), .ZN(n9073) );
  NAND2_X1 U7765 ( .A1(n9392), .A2(n9393), .ZN(n9391) );
  NAND2_X1 U7766 ( .A1(n9391), .A2(n9074), .ZN(n9374) );
  INV_X1 U7767 ( .A(n9394), .ZN(n6088) );
  NAND2_X1 U7768 ( .A1(n9383), .A2(n6088), .ZN(n9365) );
  NAND2_X1 U7769 ( .A1(n9374), .A2(n9375), .ZN(n9364) );
  INV_X1 U7770 ( .A(n9365), .ZN(n9159) );
  NOR2_X1 U7771 ( .A1(n6055), .A2(n9159), .ZN(n6089) );
  INV_X1 U7772 ( .A(n8950), .ZN(n9096) );
  XNOR2_X1 U7773 ( .A(n6090), .B(n9096), .ZN(n6093) );
  NAND2_X1 U7774 ( .A1(n9308), .A2(n9184), .ZN(n6092) );
  NAND2_X1 U7775 ( .A1(n6091), .A2(n9114), .ZN(n9177) );
  NAND2_X1 U7776 ( .A1(n6092), .A2(n9177), .ZN(n9882) );
  NAND2_X1 U7777 ( .A1(n6093), .A2(n9882), .ZN(n6101) );
  INV_X1 U7778 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9320) );
  NOR2_X1 U7779 ( .A1(n5637), .A2(n9320), .ZN(n6098) );
  INV_X1 U7780 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9534) );
  NOR2_X1 U7781 ( .A1(n6094), .A2(n9534), .ZN(n6097) );
  INV_X1 U7782 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9608) );
  NOR2_X1 U7783 ( .A1(n4279), .A2(n9608), .ZN(n6096) );
  OR3_X1 U7784 ( .A1(n6098), .A2(n6097), .A3(n6096), .ZN(n9188) );
  AOI22_X1 U7785 ( .A1(n9368), .A2(n9433), .B1(n6099), .B2(n9188), .ZN(n6100)
         );
  INV_X2 U7786 ( .A(n9982), .ZN(n9983) );
  NAND2_X1 U7787 ( .A1(n9983), .A2(n9974), .ZN(n9645) );
  INV_X1 U7788 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6506) );
  INV_X2 U7789 ( .A(n6207), .ZN(n6219) );
  NAND2_X1 U7790 ( .A1(n6425), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6106) );
  INV_X1 U7791 ( .A(n7724), .ZN(n6115) );
  INV_X1 U7792 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6113) );
  INV_X2 U7793 ( .A(n6397), .ZN(n6437) );
  NAND2_X1 U7794 ( .A1(n6437), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6122) );
  INV_X1 U7795 ( .A(n6117), .ZN(n6118) );
  AND2_X2 U7796 ( .A1(n6115), .A2(n6118), .ZN(n6308) );
  INV_X1 U7797 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U7798 ( .A1(n6185), .A2(n6184), .ZN(n6201) );
  INV_X1 U7799 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7098) );
  INV_X1 U7800 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6236) );
  INV_X1 U7801 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7802 ( .A1(n6274), .A2(n6273), .ZN(n6285) );
  INV_X1 U7803 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7691) );
  INV_X1 U7804 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6318) );
  INV_X1 U7805 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8287) );
  INV_X1 U7806 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6360) );
  INV_X1 U7807 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U7808 ( .A1(n6392), .A2(n6391), .ZN(n6394) );
  NAND2_X1 U7809 ( .A1(n8638), .A2(n6123), .ZN(n6404) );
  NAND2_X1 U7810 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(n6404), .ZN(n6116) );
  NOR2_X1 U7811 ( .A1(n6404), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6415) );
  INV_X1 U7812 ( .A(n6415), .ZN(n6417) );
  NAND2_X1 U7813 ( .A1(n6116), .A2(n6417), .ZN(n8412) );
  NAND2_X1 U7814 ( .A1(n6308), .A2(n8412), .ZN(n6121) );
  INV_X2 U7815 ( .A(n6340), .ZN(n6436) );
  NAND2_X1 U7816 ( .A1(n6436), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7817 ( .A1(n6159), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6119) );
  OR2_X1 U7818 ( .A1(n8420), .A2(n8414), .ZN(n6411) );
  NAND2_X1 U7819 ( .A1(n6394), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6124) );
  INV_X1 U7820 ( .A(n6123), .ZN(n6403) );
  NAND2_X1 U7821 ( .A1(n6124), .A2(n6403), .ZN(n8443) );
  NAND2_X1 U7822 ( .A1(n8443), .A2(n6299), .ZN(n6130) );
  INV_X1 U7823 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7824 ( .A1(n6437), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U7825 ( .A1(n6159), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6125) );
  OAI211_X1 U7826 ( .C1(n6340), .C2(n6127), .A(n6126), .B(n6125), .ZN(n6128)
         );
  INV_X1 U7827 ( .A(n6128), .ZN(n6129) );
  NAND2_X1 U7828 ( .A1(n7366), .A2(n6219), .ZN(n6132) );
  NAND2_X1 U7829 ( .A1(n6425), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6131) );
  AND2_X1 U7830 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6133) );
  OR2_X1 U7831 ( .A1(n6133), .A2(n6185), .ZN(n7192) );
  NAND2_X1 U7832 ( .A1(n6299), .A2(n7192), .ZN(n6136) );
  NAND2_X1 U7833 ( .A1(n6436), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7834 ( .A1(n6159), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6134) );
  OR2_X1 U7835 ( .A1(n8001), .A2(n6542), .ZN(n6139) );
  OR2_X1 U7836 ( .A1(n6207), .A2(n6541), .ZN(n6138) );
  OAI211_X1 U7837 ( .C1(n6443), .C2(n6718), .A(n6139), .B(n6138), .ZN(n7193)
         );
  NAND2_X1 U7838 ( .A1(n8344), .A2(n7193), .ZN(n6180) );
  INV_X1 U7839 ( .A(n6180), .ZN(n6149) );
  NAND2_X1 U7840 ( .A1(n6211), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6144) );
  INV_X1 U7841 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7201) );
  NAND2_X1 U7842 ( .A1(n6299), .A2(n7201), .ZN(n6143) );
  NAND2_X1 U7843 ( .A1(n6159), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6142) );
  INV_X1 U7844 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6140) );
  NAND4_X1 U7845 ( .A1(n6144), .A2(n6143), .A3(n6142), .A4(n6141), .ZN(n8345)
         );
  OR2_X1 U7846 ( .A1(n6207), .A2(n6539), .ZN(n6146) );
  OR2_X1 U7847 ( .A1(n8001), .A2(n6540), .ZN(n6145) );
  OAI211_X1 U7848 ( .C1(n6443), .C2(n6538), .A(n6146), .B(n6145), .ZN(n7202)
         );
  INV_X1 U7849 ( .A(n7202), .ZN(n8048) );
  NAND2_X1 U7850 ( .A1(n7109), .A2(n8048), .ZN(n7185) );
  OR2_X1 U7851 ( .A1(n8344), .A2(n7193), .ZN(n6147) );
  AND2_X1 U7852 ( .A1(n7185), .A2(n6147), .ZN(n6148) );
  NAND2_X1 U7853 ( .A1(n6211), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7854 ( .A1(n6308), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7855 ( .A1(n6170), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7856 ( .A1(n6159), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6150) );
  AND4_X2 U7857 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(n7108)
         );
  INV_X1 U7858 ( .A(n7108), .ZN(n8347) );
  OR2_X1 U7859 ( .A1(n8001), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6158) );
  OR2_X1 U7860 ( .A1(n6207), .A2(n6154), .ZN(n6157) );
  NAND2_X1 U7861 ( .A1(n6337), .A2(n6691), .ZN(n6156) );
  AND3_X2 U7862 ( .A1(n6158), .A2(n6157), .A3(n6156), .ZN(n7223) );
  INV_X1 U7863 ( .A(n7223), .ZN(n6168) );
  NAND2_X1 U7864 ( .A1(n6308), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6163) );
  NAND2_X1 U7865 ( .A1(n6211), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7866 ( .A1(n6159), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7867 ( .A1(n6170), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6160) );
  NAND4_X1 U7868 ( .A1(n6163), .A2(n6162), .A3(n6161), .A4(n6160), .ZN(n8349)
         );
  NAND2_X1 U7869 ( .A1(n6537), .A2(SI_0_), .ZN(n6165) );
  INV_X1 U7870 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6164) );
  NAND2_X1 U7871 ( .A1(n6165), .A2(n6164), .ZN(n6167) );
  AND2_X1 U7872 ( .A1(n6167), .A2(n6166), .ZN(n8778) );
  MUX2_X1 U7873 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8778), .S(n6443), .Z(n10027)
         );
  NAND2_X1 U7874 ( .A1(n8349), .A2(n10027), .ZN(n7217) );
  NAND2_X1 U7875 ( .A1(n8043), .A2(n7217), .ZN(n7216) );
  NAND2_X1 U7876 ( .A1(n7108), .A2(n6168), .ZN(n6169) );
  NAND2_X1 U7877 ( .A1(n7216), .A2(n6169), .ZN(n7106) );
  NAND2_X1 U7878 ( .A1(n6211), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7879 ( .A1(n6308), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7880 ( .A1(n6170), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7881 ( .A1(n6159), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6171) );
  NAND4_X1 U7882 ( .A1(n6174), .A2(n6173), .A3(n6172), .A4(n6171), .ZN(n8346)
         );
  OR2_X1 U7883 ( .A1(n6207), .A2(n6543), .ZN(n6178) );
  OR2_X1 U7884 ( .A1(n8001), .A2(n6544), .ZN(n6177) );
  NAND2_X1 U7885 ( .A1(n6337), .A2(n6175), .ZN(n6176) );
  NAND2_X1 U7886 ( .A1(n7106), .A2(n7107), .ZN(n7105) );
  INV_X1 U7887 ( .A(n8346), .ZN(n6848) );
  NAND2_X1 U7888 ( .A1(n6848), .A2(n8049), .ZN(n6179) );
  NAND2_X1 U7889 ( .A1(n7105), .A2(n6179), .ZN(n7198) );
  NAND2_X1 U7890 ( .A1(n8345), .A2(n7202), .ZN(n7184) );
  AND2_X1 U7891 ( .A1(n7184), .A2(n6180), .ZN(n6181) );
  NAND2_X1 U7892 ( .A1(n7198), .A2(n6181), .ZN(n6182) );
  NAND2_X1 U7893 ( .A1(n6211), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6190) );
  OR2_X1 U7894 ( .A1(n6185), .A2(n6184), .ZN(n6186) );
  NAND2_X1 U7895 ( .A1(n6201), .A2(n6186), .ZN(n7125) );
  NAND2_X1 U7896 ( .A1(n6299), .A2(n7125), .ZN(n6189) );
  NAND2_X1 U7897 ( .A1(n6436), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7898 ( .A1(n6159), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6187) );
  OR2_X1 U7899 ( .A1(n6207), .A2(n6546), .ZN(n6193) );
  OR2_X1 U7900 ( .A1(n8001), .A2(n6547), .ZN(n6192) );
  NAND2_X1 U7901 ( .A1(n6337), .A2(n4582), .ZN(n6191) );
  NAND2_X1 U7902 ( .A1(n7025), .A2(n7005), .ZN(n7155) );
  NAND2_X1 U7903 ( .A1(n6437), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6198) );
  NOR2_X1 U7904 ( .A1(n6213), .A2(n7098), .ZN(n6194) );
  OR2_X1 U7905 ( .A1(n6237), .A2(n6194), .ZN(n7279) );
  NAND2_X1 U7906 ( .A1(n6299), .A2(n7279), .ZN(n6197) );
  NAND2_X1 U7907 ( .A1(n6436), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7908 ( .A1(n6159), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6195) );
  NAND4_X1 U7909 ( .A1(n6198), .A2(n6197), .A3(n6196), .A4(n6195), .ZN(n8341)
         );
  NAND2_X1 U7910 ( .A1(n6557), .A2(n6219), .ZN(n6200) );
  AOI22_X1 U7911 ( .A1(n6425), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6337), .B2(
        n7919), .ZN(n6199) );
  NAND2_X1 U7912 ( .A1(n6200), .A2(n6199), .ZN(n7283) );
  NAND2_X1 U7913 ( .A1(n8341), .A2(n7283), .ZN(n6228) );
  INV_X1 U7914 ( .A(n6228), .ZN(n6225) );
  NAND2_X1 U7915 ( .A1(n6437), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7916 ( .A1(n6201), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U7917 ( .A1(n6212), .A2(n6202), .ZN(n7267) );
  NAND2_X1 U7918 ( .A1(n6308), .A2(n7267), .ZN(n6205) );
  NAND2_X1 U7919 ( .A1(n6159), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7920 ( .A1(n6436), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6203) );
  OR2_X1 U7921 ( .A1(n6207), .A2(n6550), .ZN(n6210) );
  OR2_X1 U7922 ( .A1(n8001), .A2(n6549), .ZN(n6209) );
  NAND2_X1 U7923 ( .A1(n6337), .A2(n6734), .ZN(n6208) );
  NAND2_X1 U7924 ( .A1(n6211), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6218) );
  AND2_X1 U7925 ( .A1(n6212), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6214) );
  OR2_X1 U7926 ( .A1(n6214), .A2(n6213), .ZN(n7165) );
  NAND2_X1 U7927 ( .A1(n6308), .A2(n7165), .ZN(n6217) );
  NAND2_X1 U7928 ( .A1(n6170), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7929 ( .A1(n6159), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7930 ( .A1(n6551), .A2(n6219), .ZN(n6220) );
  INV_X1 U7931 ( .A(n7166), .ZN(n7042) );
  NAND2_X1 U7932 ( .A1(n6222), .A2(n7042), .ZN(n6223) );
  NAND2_X1 U7933 ( .A1(n4852), .A2(n6223), .ZN(n6224) );
  INV_X1 U7934 ( .A(n6222), .ZN(n8342) );
  NAND2_X1 U7935 ( .A1(n8342), .A2(n7042), .ZN(n7271) );
  NAND2_X1 U7936 ( .A1(n6222), .A2(n7166), .ZN(n8078) );
  NAND2_X1 U7937 ( .A1(n7119), .A2(n6226), .ZN(n6232) );
  INV_X1 U7938 ( .A(n7005), .ZN(n7126) );
  NAND2_X1 U7939 ( .A1(n8343), .A2(n7126), .ZN(n7262) );
  NAND2_X1 U7940 ( .A1(n6453), .A2(n7268), .ZN(n6227) );
  AND2_X1 U7941 ( .A1(n7262), .A2(n6227), .ZN(n7158) );
  AND2_X1 U7942 ( .A1(n7158), .A2(n4855), .ZN(n7156) );
  INV_X1 U7943 ( .A(n7283), .ZN(n10063) );
  NAND2_X1 U7944 ( .A1(n7442), .A2(n10063), .ZN(n6233) );
  NAND2_X1 U7945 ( .A1(n6570), .A2(n6219), .ZN(n6235) );
  AOI22_X1 U7946 ( .A1(n6425), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6337), .B2(
        n6968), .ZN(n6234) );
  NAND2_X1 U7947 ( .A1(n6235), .A2(n6234), .ZN(n7138) );
  NAND2_X1 U7948 ( .A1(n6437), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6242) );
  OR2_X1 U7949 ( .A1(n6237), .A2(n6236), .ZN(n6238) );
  NAND2_X1 U7950 ( .A1(n6247), .A2(n6238), .ZN(n7447) );
  NAND2_X1 U7951 ( .A1(n6299), .A2(n7447), .ZN(n6241) );
  NAND2_X1 U7952 ( .A1(n6436), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7953 ( .A1(n6159), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6239) );
  NAND4_X1 U7954 ( .A1(n6242), .A2(n6241), .A3(n6240), .A4(n6239), .ZN(n8340)
         );
  NAND2_X1 U7955 ( .A1(n7138), .A2(n8340), .ZN(n6243) );
  NAND2_X1 U7956 ( .A1(n6244), .A2(n6243), .ZN(n7172) );
  NAND2_X1 U7957 ( .A1(n6575), .A2(n6219), .ZN(n6246) );
  AOI22_X1 U7958 ( .A1(n6425), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6337), .B2(
        n7895), .ZN(n6245) );
  NAND2_X1 U7959 ( .A1(n6246), .A2(n6245), .ZN(n7336) );
  NAND2_X1 U7960 ( .A1(n6437), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7961 ( .A1(n6247), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7962 ( .A1(n6256), .A2(n6248), .ZN(n7341) );
  NAND2_X1 U7963 ( .A1(n6299), .A2(n7341), .ZN(n6251) );
  NAND2_X1 U7964 ( .A1(n6436), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6250) );
  NAND2_X1 U7965 ( .A1(n6159), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6249) );
  NAND4_X1 U7966 ( .A1(n6252), .A2(n6251), .A3(n6250), .A4(n6249), .ZN(n8339)
         );
  AND2_X1 U7967 ( .A1(n7336), .A2(n8339), .ZN(n6253) );
  NAND2_X1 U7968 ( .A1(n6581), .A2(n6219), .ZN(n6255) );
  AOI22_X1 U7969 ( .A1(n6425), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6337), .B2(
        n7881), .ZN(n6254) );
  NAND2_X1 U7970 ( .A1(n6255), .A2(n6254), .ZN(n7390) );
  NAND2_X1 U7971 ( .A1(n6437), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6261) );
  NAND2_X1 U7972 ( .A1(n6256), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6257) );
  NAND2_X1 U7973 ( .A1(n6265), .A2(n6257), .ZN(n7393) );
  NAND2_X1 U7974 ( .A1(n6299), .A2(n7393), .ZN(n6260) );
  NAND2_X1 U7975 ( .A1(n6436), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U7976 ( .A1(n6159), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6258) );
  NAND4_X1 U7977 ( .A1(n6261), .A2(n6260), .A3(n6259), .A4(n6258), .ZN(n8338)
         );
  NOR2_X1 U7978 ( .A1(n7390), .A2(n8338), .ZN(n6262) );
  NAND2_X1 U7979 ( .A1(n6630), .A2(n6219), .ZN(n6264) );
  AOI22_X1 U7980 ( .A1(n6425), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6337), .B2(
        n7862), .ZN(n6263) );
  NAND2_X1 U7981 ( .A1(n6437), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6270) );
  AND2_X1 U7982 ( .A1(n6265), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6266) );
  OR2_X1 U7983 ( .A1(n6266), .A2(n6274), .ZN(n7318) );
  NAND2_X1 U7984 ( .A1(n6308), .A2(n7318), .ZN(n6269) );
  NAND2_X1 U7985 ( .A1(n6436), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6268) );
  NAND2_X1 U7986 ( .A1(n6159), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6267) );
  NAND4_X1 U7987 ( .A1(n6270), .A2(n6269), .A3(n6268), .A4(n6267), .ZN(n8337)
         );
  NAND2_X1 U7988 ( .A1(n6635), .A2(n6219), .ZN(n6272) );
  AOI22_X1 U7989 ( .A1(n6425), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6337), .B2(
        n7843), .ZN(n6271) );
  OR2_X1 U7990 ( .A1(n6274), .A2(n6273), .ZN(n6275) );
  NAND2_X1 U7991 ( .A1(n6285), .A2(n6275), .ZN(n9702) );
  NAND2_X1 U7992 ( .A1(n6308), .A2(n9702), .ZN(n6279) );
  NAND2_X1 U7993 ( .A1(n6437), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7994 ( .A1(n6159), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7995 ( .A1(n6436), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6276) );
  NAND4_X1 U7996 ( .A1(n6279), .A2(n6278), .A3(n6277), .A4(n6276), .ZN(n8336)
         );
  NOR2_X1 U7997 ( .A1(n8113), .A2(n8336), .ZN(n6280) );
  NAND2_X1 U7998 ( .A1(n8113), .A2(n8336), .ZN(n6281) );
  NAND2_X1 U7999 ( .A1(n6282), .A2(n6281), .ZN(n7487) );
  INV_X1 U8000 ( .A(n7487), .ZN(n6292) );
  NAND2_X1 U8001 ( .A1(n6639), .A2(n6219), .ZN(n6284) );
  AOI22_X1 U8002 ( .A1(n6425), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6337), .B2(
        n7825), .ZN(n6283) );
  NAND2_X1 U8003 ( .A1(n6437), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U8004 ( .A1(n6285), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U8005 ( .A1(n6296), .A2(n6286), .ZN(n7502) );
  NAND2_X1 U8006 ( .A1(n6308), .A2(n7502), .ZN(n6289) );
  NAND2_X1 U8007 ( .A1(n6436), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U8008 ( .A1(n6159), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U8009 ( .A1(n7498), .A2(n9711), .ZN(n8119) );
  INV_X1 U8010 ( .A(n9711), .ZN(n8335) );
  OR2_X1 U8011 ( .A1(n7498), .A2(n8335), .ZN(n6293) );
  NAND2_X1 U8012 ( .A1(n6665), .A2(n6219), .ZN(n6295) );
  AOI22_X1 U8013 ( .A1(n6425), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6337), .B2(
        n8368), .ZN(n6294) );
  NAND2_X1 U8014 ( .A1(n6437), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6303) );
  INV_X1 U8015 ( .A(n6306), .ZN(n6298) );
  NAND2_X1 U8016 ( .A1(n6296), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U8017 ( .A1(n6298), .A2(n6297), .ZN(n7596) );
  NAND2_X1 U8018 ( .A1(n6299), .A2(n7596), .ZN(n6302) );
  NAND2_X1 U8019 ( .A1(n6436), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U8020 ( .A1(n6159), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6300) );
  NAND2_X1 U8021 ( .A1(n7589), .A2(n7693), .ZN(n8123) );
  NAND2_X1 U8022 ( .A1(n8124), .A2(n8123), .ZN(n8207) );
  INV_X1 U8023 ( .A(n7693), .ZN(n8334) );
  NAND2_X1 U8024 ( .A1(n7589), .A2(n8334), .ZN(n7505) );
  NAND2_X1 U8025 ( .A1(n6653), .A2(n6219), .ZN(n6305) );
  AOI22_X1 U8026 ( .A1(n6425), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6337), .B2(
        n7796), .ZN(n6304) );
  NAND2_X1 U8027 ( .A1(n6437), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6312) );
  NOR2_X1 U8028 ( .A1(n6306), .A2(n7691), .ZN(n6307) );
  OR2_X1 U8029 ( .A1(n6319), .A2(n6307), .ZN(n7695) );
  NAND2_X1 U8030 ( .A1(n6308), .A2(n7695), .ZN(n6311) );
  NAND2_X1 U8031 ( .A1(n6159), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U8032 ( .A1(n6436), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6309) );
  INV_X1 U8033 ( .A(n7731), .ZN(n8333) );
  NAND2_X1 U8034 ( .A1(n7688), .A2(n8333), .ZN(n6313) );
  AND2_X1 U8035 ( .A1(n7505), .A2(n6313), .ZN(n6315) );
  INV_X1 U8036 ( .A(n6313), .ZN(n6314) );
  NAND2_X1 U8037 ( .A1(n7688), .A2(n7731), .ZN(n8128) );
  NAND2_X1 U8038 ( .A1(n8129), .A2(n8128), .ZN(n8208) );
  NAND2_X1 U8039 ( .A1(n6649), .A2(n6219), .ZN(n6317) );
  AOI22_X1 U8040 ( .A1(n6425), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6337), .B2(
        n7780), .ZN(n6316) );
  NAND2_X1 U8041 ( .A1(n6437), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6324) );
  OR2_X1 U8042 ( .A1(n6319), .A2(n6318), .ZN(n6320) );
  NAND2_X1 U8043 ( .A1(n6329), .A2(n6320), .ZN(n7735) );
  NAND2_X1 U8044 ( .A1(n6308), .A2(n7735), .ZN(n6323) );
  NAND2_X1 U8045 ( .A1(n6170), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U8046 ( .A1(n6159), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6321) );
  XNOR2_X1 U8047 ( .A(n8582), .B(n8311), .ZN(n7610) );
  NAND2_X1 U8048 ( .A1(n7611), .A2(n7610), .ZN(n6326) );
  INV_X1 U8049 ( .A(n8311), .ZN(n8332) );
  NAND2_X1 U8050 ( .A1(n8582), .A2(n8332), .ZN(n6325) );
  NAND2_X1 U8051 ( .A1(n6672), .A2(n6219), .ZN(n6328) );
  INV_X1 U8052 ( .A(n7757), .ZN(n7765) );
  AOI22_X1 U8053 ( .A1(n6425), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6337), .B2(
        n7765), .ZN(n6327) );
  NAND2_X1 U8054 ( .A1(n6437), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U8055 ( .A1(n6329), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U8056 ( .A1(n6343), .A2(n6330), .ZN(n8316) );
  NAND2_X1 U8057 ( .A1(n6299), .A2(n8316), .ZN(n6333) );
  NAND2_X1 U8058 ( .A1(n6436), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6332) );
  NAND2_X1 U8059 ( .A1(n6159), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U8060 ( .A1(n8312), .A2(n7942), .ZN(n8133) );
  INV_X1 U8061 ( .A(n7942), .ZN(n8511) );
  OR2_X1 U8062 ( .A1(n8312), .A2(n8511), .ZN(n6336) );
  NAND2_X1 U8063 ( .A1(n6898), .A2(n6219), .ZN(n6339) );
  AOI22_X1 U8064 ( .A1(n6425), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6479), .B2(
        n6337), .ZN(n6338) );
  NAND2_X1 U8065 ( .A1(n6437), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U8066 ( .A1(n6436), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6341) );
  AND2_X1 U8067 ( .A1(n6342), .A2(n6341), .ZN(n6347) );
  AND2_X1 U8068 ( .A1(n6343), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6344) );
  OR2_X1 U8069 ( .A1(n6344), .A2(n6352), .ZN(n8520) );
  NAND2_X1 U8070 ( .A1(n8520), .A2(n6299), .ZN(n6346) );
  NAND2_X1 U8071 ( .A1(n6159), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6345) );
  NAND2_X1 U8072 ( .A1(n8236), .A2(n8286), .ZN(n8141) );
  INV_X1 U8073 ( .A(n8286), .ZN(n8500) );
  NAND2_X1 U8074 ( .A1(n8236), .A2(n8500), .ZN(n6349) );
  NAND2_X1 U8075 ( .A1(n6915), .A2(n6219), .ZN(n6351) );
  NAND2_X1 U8076 ( .A1(n6425), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6350) );
  NOR2_X1 U8077 ( .A1(n6352), .A2(n8287), .ZN(n6353) );
  OR2_X1 U8078 ( .A1(n6361), .A2(n6353), .ZN(n8505) );
  NAND2_X1 U8079 ( .A1(n8505), .A2(n6299), .ZN(n6356) );
  AOI22_X1 U8080 ( .A1(n6437), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6436), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8081 ( .A1(n6159), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U8082 ( .A1(n8278), .A2(n8488), .ZN(n8145) );
  NAND2_X1 U8083 ( .A1(n8144), .A2(n8145), .ZN(n8498) );
  INV_X1 U8084 ( .A(n8488), .ZN(n8514) );
  OR2_X1 U8085 ( .A1(n8278), .A2(n8514), .ZN(n6357) );
  NAND2_X1 U8086 ( .A1(n8497), .A2(n6357), .ZN(n8486) );
  NAND2_X1 U8087 ( .A1(n6947), .A2(n6219), .ZN(n6359) );
  NAND2_X1 U8088 ( .A1(n6425), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6358) );
  OR2_X1 U8089 ( .A1(n6361), .A2(n6360), .ZN(n6362) );
  NAND2_X1 U8090 ( .A1(n6370), .A2(n6362), .ZN(n8492) );
  NAND2_X1 U8091 ( .A1(n8492), .A2(n6299), .ZN(n6365) );
  AOI22_X1 U8092 ( .A1(n6437), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n6436), .B2(
        P2_REG0_REG_21__SCAN_IN), .ZN(n6364) );
  NAND2_X1 U8093 ( .A1(n6159), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8094 ( .A1(n8245), .A2(n8288), .ZN(n8152) );
  NAND2_X1 U8095 ( .A1(n8151), .A2(n8152), .ZN(n8187) );
  NAND2_X1 U8096 ( .A1(n8486), .A2(n8187), .ZN(n6367) );
  INV_X1 U8097 ( .A(n8288), .ZN(n8501) );
  OR2_X1 U8098 ( .A1(n8245), .A2(n8501), .ZN(n6366) );
  NAND2_X1 U8099 ( .A1(n6367), .A2(n6366), .ZN(n8473) );
  NAND2_X1 U8100 ( .A1(n7080), .A2(n6219), .ZN(n6369) );
  NAND2_X1 U8101 ( .A1(n6425), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6368) );
  NAND2_X1 U8102 ( .A1(n6370), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U8103 ( .A1(n6380), .A2(n6371), .ZN(n8481) );
  NAND2_X1 U8104 ( .A1(n8481), .A2(n6299), .ZN(n6376) );
  INV_X1 U8105 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U8106 ( .A1(n6170), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8107 ( .A1(n6159), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6372) );
  OAI211_X1 U8108 ( .C1(n6397), .C2(n8630), .A(n6373), .B(n6372), .ZN(n6374)
         );
  INV_X1 U8109 ( .A(n6374), .ZN(n6375) );
  XNOR2_X1 U8110 ( .A(n8029), .B(n8489), .ZN(n8474) );
  NAND2_X1 U8111 ( .A1(n8473), .A2(n8474), .ZN(n8472) );
  NAND2_X1 U8112 ( .A1(n8756), .A2(n8489), .ZN(n6377) );
  NAND2_X1 U8113 ( .A1(n8472), .A2(n6377), .ZN(n8462) );
  NAND2_X1 U8114 ( .A1(n7148), .A2(n6219), .ZN(n6379) );
  NAND2_X1 U8115 ( .A1(n6425), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6378) );
  AND2_X1 U8116 ( .A1(n6380), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6381) );
  OR2_X1 U8117 ( .A1(n6381), .A2(n6392), .ZN(n8467) );
  NAND2_X1 U8118 ( .A1(n8467), .A2(n6299), .ZN(n6386) );
  INV_X1 U8119 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8685) );
  NAND2_X1 U8120 ( .A1(n6436), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U8121 ( .A1(n6159), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6382) );
  OAI211_X1 U8122 ( .C1(n6397), .C2(n8685), .A(n6383), .B(n6382), .ZN(n6384)
         );
  INV_X1 U8123 ( .A(n6384), .ZN(n6385) );
  NAND2_X1 U8124 ( .A1(n6386), .A2(n6385), .ZN(n8475) );
  NAND2_X1 U8125 ( .A1(n7962), .A2(n8475), .ZN(n6387) );
  INV_X1 U8126 ( .A(n8475), .ZN(n8300) );
  NAND2_X1 U8127 ( .A1(n8752), .A2(n8300), .ZN(n6388) );
  NAND2_X1 U8128 ( .A1(n7299), .A2(n6219), .ZN(n6390) );
  NAND2_X1 U8129 ( .A1(n6425), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6389) );
  OR2_X1 U8130 ( .A1(n6392), .A2(n6391), .ZN(n6393) );
  NAND2_X1 U8131 ( .A1(n6394), .A2(n6393), .ZN(n8457) );
  NAND2_X1 U8132 ( .A1(n8457), .A2(n6299), .ZN(n6400) );
  INV_X1 U8133 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U8134 ( .A1(n6170), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U8135 ( .A1(n6159), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6395) );
  OAI211_X1 U8136 ( .C1(n6397), .C2(n8553), .A(n6396), .B(n6395), .ZN(n6398)
         );
  INV_X1 U8137 ( .A(n6398), .ZN(n6399) );
  NAND2_X1 U8138 ( .A1(n8273), .A2(n8464), .ZN(n8161) );
  INV_X1 U8139 ( .A(n8464), .ZN(n8331) );
  NAND2_X1 U8140 ( .A1(n8442), .A2(n8455), .ZN(n8165) );
  NAND2_X1 U8141 ( .A1(n8427), .A2(n8165), .ZN(n8436) );
  NAND2_X1 U8142 ( .A1(n8437), .A2(n8436), .ZN(n8435) );
  NAND2_X1 U8143 ( .A1(n7471), .A2(n6219), .ZN(n6402) );
  NAND2_X1 U8144 ( .A1(n6425), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6401) );
  NAND2_X1 U8145 ( .A1(n6437), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U8146 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(n6403), .ZN(n6405) );
  NAND2_X1 U8147 ( .A1(n6405), .A2(n6404), .ZN(n8421) );
  NAND2_X1 U8148 ( .A1(n6308), .A2(n8421), .ZN(n6408) );
  NAND2_X1 U8149 ( .A1(n6159), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8150 ( .A1(n6170), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U8151 ( .A1(n8743), .A2(n8438), .ZN(n6410) );
  NAND2_X1 U8152 ( .A1(n6411), .A2(n8403), .ZN(n6412) );
  OAI21_X1 U8153 ( .B1(n8537), .B2(n8391), .A(n6412), .ZN(n8388) );
  INV_X1 U8154 ( .A(n8388), .ZN(n6424) );
  NAND2_X1 U8155 ( .A1(n7600), .A2(n6219), .ZN(n6414) );
  NAND2_X1 U8156 ( .A1(n6425), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U8157 ( .A1(n6437), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6422) );
  INV_X1 U8158 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8159 ( .A1(n6416), .A2(n6415), .ZN(n8374) );
  NAND2_X1 U8160 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n6417), .ZN(n6418) );
  NAND2_X1 U8161 ( .A1(n8374), .A2(n6418), .ZN(n8397) );
  NAND2_X1 U8162 ( .A1(n6299), .A2(n8397), .ZN(n6421) );
  NAND2_X1 U8163 ( .A1(n6170), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6420) );
  NAND2_X1 U8164 ( .A1(n6159), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U8165 ( .A1(n7722), .A2(n6219), .ZN(n6427) );
  NAND2_X1 U8166 ( .A1(n6425), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6426) );
  INV_X1 U8167 ( .A(n8374), .ZN(n6428) );
  NAND2_X1 U8168 ( .A1(n6299), .A2(n6428), .ZN(n8010) );
  NAND2_X1 U8169 ( .A1(n6437), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U8170 ( .A1(n6159), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U8171 ( .A1(n6170), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6429) );
  NAND2_X1 U8172 ( .A1(n8179), .A2(n8015), .ZN(n8177) );
  XNOR2_X1 U8173 ( .A(n6432), .B(n6473), .ZN(n6446) );
  INV_X1 U8174 ( .A(n8183), .ZN(n6514) );
  NAND2_X1 U8175 ( .A1(n6804), .A2(n6514), .ZN(n6435) );
  NAND2_X1 U8176 ( .A1(n6479), .A2(n8226), .ZN(n6481) );
  NAND2_X1 U8177 ( .A1(n6435), .A2(n6481), .ZN(n8510) );
  NAND2_X1 U8178 ( .A1(n6436), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8179 ( .A1(n6437), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8180 ( .A1(n6159), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6438) );
  AND4_X1 U8181 ( .A1(n8010), .A2(n6440), .A3(n6439), .A4(n6438), .ZN(n8004)
         );
  NAND2_X1 U8182 ( .A1(n6441), .A2(n8224), .ZN(n6442) );
  NAND2_X1 U8183 ( .A1(n6443), .A2(n6442), .ZN(n8389) );
  NAND2_X1 U8184 ( .A1(n6443), .A2(P2_B_REG_SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8185 ( .A1(n8513), .A2(n6444), .ZN(n8372) );
  OAI22_X1 U8186 ( .A1(n8004), .A2(n8372), .B1(n6472), .B2(n9710), .ZN(n6445)
         );
  AOI21_X1 U8187 ( .B1(n6446), .B2(n8510), .A(n6445), .ZN(n6478) );
  INV_X1 U8188 ( .A(n8349), .ZN(n6447) );
  NAND2_X1 U8189 ( .A1(n6447), .A2(n10027), .ZN(n8036) );
  INV_X1 U8190 ( .A(n8036), .ZN(n6448) );
  INV_X1 U8191 ( .A(n7107), .ZN(n8042) );
  NAND2_X1 U8192 ( .A1(n7104), .A2(n8042), .ZN(n6451) );
  INV_X1 U8193 ( .A(n8049), .ZN(n6450) );
  NAND2_X1 U8194 ( .A1(n6848), .A2(n6450), .ZN(n8051) );
  NAND2_X1 U8195 ( .A1(n6451), .A2(n8051), .ZN(n7200) );
  XNOR2_X1 U8196 ( .A(n8345), .B(n7202), .ZN(n8190) );
  NAND2_X1 U8197 ( .A1(n7200), .A2(n8190), .ZN(n6452) );
  NAND2_X1 U8198 ( .A1(n7109), .A2(n7202), .ZN(n8067) );
  INV_X1 U8199 ( .A(n7193), .ZN(n7015) );
  NAND2_X1 U8200 ( .A1(n8344), .A2(n7015), .ZN(n8069) );
  INV_X1 U8201 ( .A(n8344), .ZN(n7000) );
  NAND2_X1 U8202 ( .A1(n7000), .A2(n7193), .ZN(n8060) );
  NAND2_X1 U8203 ( .A1(n8343), .A2(n7005), .ZN(n8068) );
  NAND2_X1 U8204 ( .A1(n7154), .A2(n7268), .ZN(n8063) );
  NAND2_X1 U8205 ( .A1(n7025), .A2(n7126), .ZN(n8059) );
  AND2_X1 U8206 ( .A1(n8063), .A2(n8059), .ZN(n8073) );
  NAND2_X1 U8207 ( .A1(n7260), .A2(n8073), .ZN(n7152) );
  NAND2_X1 U8208 ( .A1(n6453), .A2(n6454), .ZN(n8062) );
  NAND2_X1 U8209 ( .A1(n7152), .A2(n8062), .ZN(n6455) );
  NAND2_X1 U8210 ( .A1(n10063), .A2(n8341), .ZN(n8083) );
  AND2_X1 U8211 ( .A1(n8083), .A2(n7271), .ZN(n8080) );
  NAND2_X1 U8212 ( .A1(n7272), .A2(n8080), .ZN(n6456) );
  NAND2_X1 U8213 ( .A1(n7442), .A2(n7283), .ZN(n8085) );
  NAND2_X1 U8214 ( .A1(n6456), .A2(n8085), .ZN(n7440) );
  OR2_X1 U8215 ( .A1(n7278), .A2(n7138), .ZN(n8084) );
  NAND2_X1 U8216 ( .A1(n7138), .A2(n7278), .ZN(n8089) );
  NAND2_X1 U8217 ( .A1(n8084), .A2(n8089), .ZN(n8197) );
  INV_X1 U8218 ( .A(n8339), .ZN(n7441) );
  OR2_X1 U8219 ( .A1(n7336), .A2(n7441), .ZN(n8097) );
  AND2_X1 U8220 ( .A1(n8097), .A2(n8084), .ZN(n8091) );
  NAND2_X1 U8221 ( .A1(n7390), .A2(n7385), .ZN(n8099) );
  NAND2_X1 U8222 ( .A1(n7336), .A2(n7441), .ZN(n8090) );
  AND2_X1 U8223 ( .A1(n8099), .A2(n8090), .ZN(n8103) );
  OR2_X1 U8224 ( .A1(n7390), .A2(n7385), .ZN(n8101) );
  NAND2_X1 U8225 ( .A1(n6457), .A2(n8101), .ZN(n7250) );
  NAND2_X1 U8226 ( .A1(n7315), .A2(n9709), .ZN(n8108) );
  XNOR2_X1 U8227 ( .A(n8113), .B(n8336), .ZN(n9707) );
  INV_X1 U8228 ( .A(n8336), .ZN(n8112) );
  OR2_X1 U8229 ( .A1(n8113), .A2(n8112), .ZN(n8114) );
  NAND2_X1 U8230 ( .A1(n7490), .A2(n8205), .ZN(n6458) );
  NAND2_X1 U8231 ( .A1(n6458), .A2(n8118), .ZN(n7425) );
  INV_X1 U8232 ( .A(n8207), .ZN(n8121) );
  INV_X1 U8233 ( .A(n8208), .ZN(n8126) );
  NAND2_X1 U8234 ( .A1(n7614), .A2(n6459), .ZN(n7613) );
  NAND2_X1 U8235 ( .A1(n8582), .A2(n8311), .ZN(n8034) );
  AND2_X1 U8236 ( .A1(n8033), .A2(n8517), .ZN(n8138) );
  NAND2_X1 U8237 ( .A1(n6460), .A2(n8141), .ZN(n8503) );
  NAND2_X1 U8238 ( .A1(n6461), .A2(n8151), .ZN(n8479) );
  INV_X1 U8239 ( .A(n8474), .ZN(n8478) );
  INV_X1 U8240 ( .A(n8489), .ZN(n8253) );
  NAND2_X1 U8241 ( .A1(n8756), .A2(n8253), .ZN(n8027) );
  NAND2_X1 U8242 ( .A1(n7962), .A2(n8300), .ZN(n8184) );
  NAND2_X1 U8243 ( .A1(n6462), .A2(n8184), .ZN(n8459) );
  INV_X1 U8244 ( .A(n8161), .ZN(n6463) );
  INV_X1 U8245 ( .A(n8436), .ZN(n8447) );
  INV_X1 U8246 ( .A(n8022), .ZN(n6464) );
  NAND2_X1 U8247 ( .A1(n8426), .A2(n8438), .ZN(n8023) );
  AND2_X1 U8248 ( .A1(n8447), .A2(n6466), .ZN(n6465) );
  NAND2_X1 U8249 ( .A1(n8448), .A2(n6465), .ZN(n6470) );
  INV_X1 U8250 ( .A(n6466), .ZN(n6468) );
  AND2_X1 U8251 ( .A1(n8427), .A2(n8022), .ZN(n6467) );
  NAND2_X1 U8252 ( .A1(n6470), .A2(n6469), .ZN(n8411) );
  XNOR2_X2 U8253 ( .A(n8537), .B(n8391), .ZN(n8410) );
  NAND2_X1 U8254 ( .A1(n8533), .A2(n6472), .ZN(n6471) );
  INV_X1 U8255 ( .A(n6804), .ZN(n8011) );
  INV_X1 U8256 ( .A(n8226), .ZN(n7081) );
  NAND2_X1 U8257 ( .A1(n8011), .A2(n7081), .ZN(n10068) );
  AOI21_X1 U8258 ( .B1(n6514), .B2(n7081), .A(n6479), .ZN(n6474) );
  AND2_X1 U8259 ( .A1(n10068), .A2(n6474), .ZN(n6476) );
  AND2_X1 U8260 ( .A1(n8183), .A2(n8221), .ZN(n6508) );
  INV_X1 U8261 ( .A(n6508), .ZN(n6475) );
  NAND2_X1 U8262 ( .A1(n6476), .A2(n6483), .ZN(n7526) );
  NAND2_X1 U8263 ( .A1(n6478), .A2(n6477), .ZN(n8380) );
  INV_X1 U8264 ( .A(n8387), .ZN(n6480) );
  AND2_X1 U8265 ( .A1(n8183), .A2(n6479), .ZN(n8445) );
  NOR2_X1 U8266 ( .A1(n8380), .A2(n4840), .ZN(n6521) );
  NAND2_X1 U8267 ( .A1(n6780), .A2(n6588), .ZN(n6925) );
  INV_X1 U8268 ( .A(n6807), .ZN(n8188) );
  INV_X1 U8269 ( .A(n6481), .ZN(n6482) );
  NAND2_X1 U8270 ( .A1(n8188), .A2(n6482), .ZN(n6788) );
  INV_X1 U8271 ( .A(n6483), .ZN(n6927) );
  INV_X1 U8272 ( .A(n6925), .ZN(n6786) );
  NAND2_X1 U8273 ( .A1(n6927), .A2(n6786), .ZN(n8225) );
  OAI21_X1 U8274 ( .B1(n6925), .B2(n6788), .A(n8225), .ZN(n6500) );
  XNOR2_X1 U8275 ( .A(n7370), .B(P2_B_REG_SCAN_IN), .ZN(n6484) );
  AOI21_X1 U8276 ( .B1(n7748), .B2(n6484), .A(n7474), .ZN(n6487) );
  INV_X1 U8277 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U8278 ( .A1(n6487), .A2(n6485), .ZN(n6486) );
  NAND2_X1 U8279 ( .A1(n7370), .A2(n7474), .ZN(n6586) );
  INV_X1 U8280 ( .A(n6509), .ZN(n6488) );
  OR2_X1 U8281 ( .A1(n6488), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6490) );
  NAND2_X1 U8282 ( .A1(n7748), .A2(n7474), .ZN(n6489) );
  NAND2_X1 U8283 ( .A1(n6490), .A2(n6489), .ZN(n6563) );
  NOR2_X1 U8284 ( .A1(n6806), .A2(n6563), .ZN(n6921) );
  NOR4_X1 U8285 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6499) );
  OR4_X1 U8286 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6496) );
  NOR4_X1 U8287 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6494) );
  NOR4_X1 U8288 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6493) );
  NOR4_X1 U8289 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6492) );
  NOR4_X1 U8290 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6491) );
  NAND4_X1 U8291 ( .A1(n6494), .A2(n6493), .A3(n6492), .A4(n6491), .ZN(n6495)
         );
  NOR4_X1 U8292 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6496), .A4(n6495), .ZN(n6498) );
  NOR4_X1 U8293 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6497) );
  NAND3_X1 U8294 ( .A1(n6499), .A2(n6498), .A3(n6497), .ZN(n6510) );
  NAND2_X1 U8295 ( .A1(n6509), .A2(n6510), .ZN(n6502) );
  AND2_X1 U8296 ( .A1(n6921), .A2(n6502), .ZN(n6790) );
  NAND2_X1 U8297 ( .A1(n6500), .A2(n6790), .ZN(n6505) );
  AND2_X1 U8298 ( .A1(n8137), .A2(n10068), .ZN(n6791) );
  NAND2_X1 U8299 ( .A1(n6788), .A2(n6791), .ZN(n6501) );
  OR2_X1 U8300 ( .A1(n10068), .A2(n8445), .ZN(n9705) );
  NAND2_X1 U8301 ( .A1(n6501), .A2(n9705), .ZN(n6784) );
  NAND2_X1 U8302 ( .A1(n6806), .A2(n6563), .ZN(n6512) );
  INV_X1 U8303 ( .A(n6502), .ZN(n6503) );
  NOR2_X1 U8304 ( .A1(n6512), .A2(n6503), .ZN(n6794) );
  NAND3_X1 U8305 ( .A1(n6784), .A2(n6786), .A3(n6794), .ZN(n6504) );
  INV_X2 U8306 ( .A(n10092), .ZN(n10094) );
  OR2_X1 U8307 ( .A1(n10092), .A2(n10068), .ZN(n8768) );
  NAND2_X1 U8308 ( .A1(n6507), .A2(n4842), .ZN(P2_U3456) );
  INV_X1 U8309 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6522) );
  OR2_X1 U8310 ( .A1(n8137), .A2(n6508), .ZN(n6781) );
  OR2_X1 U8311 ( .A1(n6509), .A2(n6925), .ZN(n6569) );
  OAI21_X1 U8312 ( .B1(n6510), .B2(n6925), .A(n6569), .ZN(n6511) );
  NAND2_X1 U8313 ( .A1(n6781), .A2(n6511), .ZN(n6922) );
  NAND2_X1 U8314 ( .A1(n10072), .A2(n8011), .ZN(n6926) );
  NAND2_X1 U8315 ( .A1(n6926), .A2(n6512), .ZN(n6513) );
  NOR2_X1 U8316 ( .A1(n6922), .A2(n6513), .ZN(n6520) );
  NAND3_X1 U8317 ( .A1(n6514), .A2(n8226), .A3(n8221), .ZN(n6515) );
  NAND2_X1 U8318 ( .A1(n8137), .A2(n6515), .ZN(n6517) );
  OR2_X1 U8319 ( .A1(n6563), .A2(n6517), .ZN(n6519) );
  INV_X1 U8320 ( .A(n6806), .ZN(n6516) );
  NAND2_X1 U8321 ( .A1(n6517), .A2(n6516), .ZN(n6518) );
  AND2_X2 U8322 ( .A1(n6520), .A2(n6920), .ZN(n10121) );
  NAND2_X1 U8323 ( .A1(n10121), .A2(n10028), .ZN(n8576) );
  NAND2_X1 U8324 ( .A1(n6523), .A2(n4847), .ZN(P2_U3488) );
  MUX2_X1 U8325 ( .A(n6525), .B(n6524), .S(n9998), .Z(n6526) );
  NAND2_X1 U8326 ( .A1(n6526), .A2(n4848), .ZN(P1_U3551) );
  INV_X1 U8327 ( .A(n6527), .ZN(n6528) );
  OR2_X2 U8328 ( .A1(n6529), .A2(n6528), .ZN(n9211) );
  INV_X1 U8329 ( .A(n9211), .ZN(P1_U3973) );
  AND2_X1 U8330 ( .A1(n6530), .A2(P1_U3086), .ZN(n7147) );
  INV_X2 U8331 ( .A(n7147), .ZN(n9658) );
  OAI222_X1 U8332 ( .A1(n6604), .A2(P1_U3086), .B1(n9658), .B2(n6553), .C1(
        n6531), .C2(n7993), .ZN(P1_U3354) );
  OAI222_X1 U8333 ( .A1(n9224), .A2(P1_U3086), .B1(n9658), .B2(n6539), .C1(
        n6532), .C2(n7993), .ZN(P1_U3352) );
  OAI222_X1 U8334 ( .A1(n6534), .A2(P1_U3086), .B1(n9658), .B2(n6543), .C1(
        n6533), .C2(n7993), .ZN(P1_U3353) );
  OAI222_X1 U8335 ( .A1(n9240), .A2(P1_U3086), .B1(n9658), .B2(n6541), .C1(
        n6535), .C2(n7993), .ZN(P1_U3351) );
  AND2_X1 U8336 ( .A1(n6536), .A2(P2_U3151), .ZN(n8775) );
  NAND2_X1 U8337 ( .A1(n6537), .A2(P2_U3151), .ZN(n8777) );
  OAI222_X1 U8338 ( .A1(n7747), .A2(n6540), .B1(n8777), .B2(n6539), .C1(
        P2_U3151), .C2(n6538), .ZN(P2_U3292) );
  CLKBUF_X1 U8339 ( .A(n8777), .Z(n7750) );
  OAI222_X1 U8340 ( .A1(n7747), .A2(n6542), .B1(n7750), .B2(n6541), .C1(
        P2_U3151), .C2(n6718), .ZN(P2_U3291) );
  OAI222_X1 U8341 ( .A1(n7747), .A2(n6544), .B1(n7750), .B2(n6543), .C1(
        P2_U3151), .C2(n10012), .ZN(P2_U3293) );
  OAI222_X1 U8342 ( .A1(n9749), .A2(P1_U3086), .B1(n9658), .B2(n6546), .C1(
        n6545), .C2(n7993), .ZN(P1_U3350) );
  OAI222_X1 U8343 ( .A1(n7747), .A2(n6547), .B1(n8777), .B2(n6546), .C1(
        P2_U3151), .C2(n6769), .ZN(P2_U3290) );
  OAI222_X1 U8344 ( .A1(n7747), .A2(n6549), .B1(n7750), .B2(n6550), .C1(
        P2_U3151), .C2(n6548), .ZN(P2_U3289) );
  OAI222_X1 U8345 ( .A1(n9764), .A2(P1_U3086), .B1(n9658), .B2(n6550), .C1(
        n8651), .C2(n7993), .ZN(P1_U3349) );
  INV_X1 U8346 ( .A(n6551), .ZN(n6555) );
  INV_X1 U8347 ( .A(n7993), .ZN(n6673) );
  AOI22_X1 U8348 ( .A1(n9683), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n6673), .ZN(n6552) );
  OAI21_X1 U8349 ( .B1(n6555), .B2(n9658), .A(n6552), .ZN(P1_U3348) );
  OAI222_X1 U8350 ( .A1(n7747), .A2(n4857), .B1(n7750), .B2(n6553), .C1(
        P2_U3151), .C2(n6691), .ZN(P2_U3294) );
  INV_X1 U8351 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6556) );
  OAI222_X1 U8352 ( .A1(n7747), .A2(n6556), .B1(n7750), .B2(n6555), .C1(
        P2_U3151), .C2(n6554), .ZN(P2_U3288) );
  INV_X1 U8353 ( .A(n6557), .ZN(n6560) );
  AOI22_X1 U8354 ( .A1(n9696), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n6673), .ZN(n6558) );
  OAI21_X1 U8355 ( .B1(n6560), .B2(n9658), .A(n6558), .ZN(P1_U3347) );
  OAI222_X1 U8356 ( .A1(n7747), .A2(n6561), .B1(n7750), .B2(n6560), .C1(
        P2_U3151), .C2(n6559), .ZN(P2_U3287) );
  NAND2_X1 U8357 ( .A1(n6925), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6562) );
  OAI21_X1 U8358 ( .B1(n6563), .B2(n6925), .A(n6562), .ZN(P2_U3377) );
  NOR2_X1 U8359 ( .A1(n9647), .A2(n6564), .ZN(n6589) );
  INV_X1 U8360 ( .A(n6589), .ZN(n6568) );
  NAND2_X1 U8361 ( .A1(n8918), .A2(n6565), .ZN(n6566) );
  NAND2_X1 U8362 ( .A1(n6567), .A2(n6566), .ZN(n6590) );
  AND2_X1 U8363 ( .A1(n6568), .A2(n6590), .ZN(n9735) );
  NOR2_X1 U8364 ( .A1(n9735), .A2(P1_U3973), .ZN(P1_U3085) );
  AND2_X1 U8365 ( .A1(n6569), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8366 ( .A1(n6569), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8367 ( .A1(n6569), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8368 ( .A1(n6569), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8369 ( .A1(n6569), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8370 ( .A1(n6569), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8371 ( .A1(n6569), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8372 ( .A1(n6569), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8373 ( .A1(n6569), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8374 ( .A1(n6569), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8375 ( .A1(n6569), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  INV_X1 U8376 ( .A(n6570), .ZN(n6573) );
  OAI222_X1 U8377 ( .A1(n7747), .A2(n6572), .B1(n7750), .B2(n6573), .C1(
        P2_U3151), .C2(n6571), .ZN(P2_U3286) );
  INV_X1 U8378 ( .A(n6870), .ZN(n6626) );
  OAI222_X1 U8379 ( .A1(n7993), .A2(n6574), .B1(n9658), .B2(n6573), .C1(n6626), 
        .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U8380 ( .A(n6575), .ZN(n6579) );
  AOI22_X1 U8381 ( .A1(n9669), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n6673), .ZN(n6576) );
  OAI21_X1 U8382 ( .B1(n6579), .B2(n9658), .A(n6576), .ZN(P1_U3345) );
  OAI222_X1 U8383 ( .A1(n7750), .A2(n6579), .B1(n6578), .B2(P2_U3151), .C1(
        n6577), .C2(n7747), .ZN(P2_U3285) );
  INV_X1 U8384 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n8690) );
  NOR2_X1 U8385 ( .A1(n6580), .A2(n8690), .ZN(P2_U3259) );
  INV_X1 U8386 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n8672) );
  NOR2_X1 U8387 ( .A1(n6580), .A2(n8672), .ZN(P2_U3255) );
  INV_X1 U8388 ( .A(n6581), .ZN(n6584) );
  AOI22_X1 U8389 ( .A1(n9769), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n6673), .ZN(n6582) );
  OAI21_X1 U8390 ( .B1(n6584), .B2(n9658), .A(n6582), .ZN(P1_U3344) );
  OAI222_X1 U8391 ( .A1(n7747), .A2(n8631), .B1(n7750), .B2(n6584), .C1(
        P2_U3151), .C2(n6583), .ZN(P2_U3284) );
  NAND2_X1 U8392 ( .A1(n8916), .A2(P1_U3973), .ZN(n6585) );
  OAI21_X1 U8393 ( .B1(P1_U3973), .B2(n8000), .A(n6585), .ZN(P1_U3585) );
  INV_X1 U8394 ( .A(n6586), .ZN(n6587) );
  AOI22_X1 U8395 ( .A1(n6569), .A2(n6485), .B1(n6588), .B2(n6587), .ZN(
        P2_U3376) );
  OR2_X1 U8396 ( .A1(n6590), .A2(n6589), .ZN(n9738) );
  OR2_X1 U8397 ( .A1(n7620), .A2(n9728), .ZN(n6591) );
  OR2_X1 U8398 ( .A1(n9738), .A2(n6591), .ZN(n9814) );
  INV_X1 U8399 ( .A(n9814), .ZN(n9827) );
  NOR2_X1 U8400 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6870), .ZN(n6592) );
  AOI21_X1 U8401 ( .B1(n6870), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6592), .ZN(
        n6602) );
  XNOR2_X1 U8402 ( .A(n9683), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n9679) );
  MUX2_X1 U8403 ( .A(n5051), .B(P1_REG2_REG_1__SCAN_IN), .S(n6604), .Z(n9218)
         );
  NAND2_X1 U8404 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6823) );
  INV_X1 U8405 ( .A(n6823), .ZN(n9217) );
  NAND2_X1 U8406 ( .A1(n9218), .A2(n9217), .ZN(n9216) );
  INV_X1 U8407 ( .A(n6604), .ZN(n9219) );
  NAND2_X1 U8408 ( .A1(n9219), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U8409 ( .A1(n9216), .A2(n6593), .ZN(n6827) );
  NAND2_X1 U8410 ( .A1(n6832), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6595) );
  OAI21_X1 U8411 ( .B1(n6832), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6595), .ZN(
        n6594) );
  INV_X1 U8412 ( .A(n6594), .ZN(n6828) );
  NAND2_X1 U8413 ( .A1(n6827), .A2(n6828), .ZN(n6826) );
  NAND2_X1 U8414 ( .A1(n6826), .A2(n6595), .ZN(n9230) );
  XNOR2_X1 U8415 ( .A(n9224), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9231) );
  NAND2_X1 U8416 ( .A1(n9230), .A2(n9231), .ZN(n9229) );
  OR2_X1 U8417 ( .A1(n9224), .A2(n6596), .ZN(n6597) );
  NAND2_X1 U8418 ( .A1(n9229), .A2(n6597), .ZN(n9247) );
  MUX2_X1 U8419 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6941), .S(n6609), .Z(n9248)
         );
  NAND2_X1 U8420 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6612), .ZN(n6598) );
  OAI21_X1 U8421 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6612), .A(n6598), .ZN(
        n9745) );
  NOR2_X1 U8422 ( .A1(n9744), .A2(n9745), .ZN(n9743) );
  NAND2_X1 U8423 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n6613), .ZN(n6599) );
  OAI21_X1 U8424 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6613), .A(n6599), .ZN(
        n9760) );
  NOR2_X1 U8425 ( .A1(n9759), .A2(n9760), .ZN(n9758) );
  NOR2_X1 U8426 ( .A1(n9679), .A2(n9680), .ZN(n9678) );
  NAND2_X1 U8427 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n9696), .ZN(n6600) );
  OAI21_X1 U8428 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9696), .A(n6600), .ZN(
        n9692) );
  NOR2_X1 U8429 ( .A1(n9693), .A2(n9692), .ZN(n9691) );
  AOI21_X1 U8430 ( .B1(n9696), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9691), .ZN(
        n6601) );
  NAND2_X1 U8431 ( .A1(n6602), .A2(n6601), .ZN(n6863) );
  OAI21_X1 U8432 ( .B1(n6602), .B2(n6601), .A(n6863), .ZN(n6628) );
  OR2_X1 U8433 ( .A1(n9738), .A2(n9182), .ZN(n9782) );
  AOI22_X1 U8434 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n6870), .B1(n6626), .B2(
        n5180), .ZN(n6621) );
  XNOR2_X1 U8435 ( .A(n9683), .B(n6603), .ZN(n9674) );
  NAND2_X1 U8436 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(n6613), .ZN(n6616) );
  MUX2_X1 U8437 ( .A(n5054), .B(P1_REG1_REG_1__SCAN_IN), .S(n6604), .Z(n9215)
         );
  AND2_X1 U8438 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9214) );
  NAND2_X1 U8439 ( .A1(n9215), .A2(n9214), .ZN(n9213) );
  NAND2_X1 U8440 ( .A1(n9219), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U8441 ( .A1(n9213), .A2(n6605), .ZN(n6830) );
  XNOR2_X1 U8442 ( .A(n6832), .B(n9985), .ZN(n6831) );
  NAND2_X1 U8443 ( .A1(n6830), .A2(n6831), .ZN(n6829) );
  NAND2_X1 U8444 ( .A1(n6832), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U8445 ( .A1(n6829), .A2(n6606), .ZN(n9233) );
  XNOR2_X1 U8446 ( .A(n9224), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9234) );
  NAND2_X1 U8447 ( .A1(n9233), .A2(n9234), .ZN(n9232) );
  OR2_X1 U8448 ( .A1(n9224), .A2(n6607), .ZN(n6608) );
  NAND2_X1 U8449 ( .A1(n9232), .A2(n6608), .ZN(n9243) );
  MUX2_X1 U8450 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n5019), .S(n6609), .Z(n9244)
         );
  NAND2_X1 U8451 ( .A1(n9243), .A2(n9244), .ZN(n9242) );
  NAND2_X1 U8452 ( .A1(n6609), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6610) );
  AND2_X1 U8453 ( .A1(n9242), .A2(n6610), .ZN(n9741) );
  NAND2_X1 U8454 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6612), .ZN(n6611) );
  OAI21_X1 U8455 ( .B1(n6612), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6611), .ZN(
        n9740) );
  NOR2_X1 U8456 ( .A1(n9741), .A2(n9740), .ZN(n9739) );
  AOI21_X1 U8457 ( .B1(n6612), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9739), .ZN(
        n9755) );
  OR2_X1 U8458 ( .A1(n6613), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U8459 ( .A1(n6614), .A2(n6616), .ZN(n9756) );
  NOR2_X1 U8460 ( .A1(n9755), .A2(n9756), .ZN(n9754) );
  INV_X1 U8461 ( .A(n9754), .ZN(n6615) );
  NAND2_X1 U8462 ( .A1(n6616), .A2(n6615), .ZN(n9673) );
  AND2_X1 U8463 ( .A1(n9683), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6617) );
  OR2_X1 U8464 ( .A1(n9696), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6619) );
  NAND2_X1 U8465 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n9696), .ZN(n6618) );
  AND2_X1 U8466 ( .A1(n6619), .A2(n6618), .ZN(n9687) );
  AOI21_X1 U8467 ( .B1(n9696), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9690), .ZN(
        n6620) );
  NAND2_X1 U8468 ( .A1(n6621), .A2(n6620), .ZN(n6869) );
  OAI21_X1 U8469 ( .B1(n6621), .B2(n6620), .A(n6869), .ZN(n6623) );
  OR2_X1 U8470 ( .A1(n9738), .A2(n6622), .ZN(n9824) );
  INV_X1 U8471 ( .A(n9824), .ZN(n9778) );
  NAND2_X1 U8472 ( .A1(n6623), .A2(n9778), .ZN(n6625) );
  AND2_X1 U8473 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7560) );
  AOI21_X1 U8474 ( .B1(n9735), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7560), .ZN(
        n6624) );
  OAI211_X1 U8475 ( .C1(n9782), .C2(n6626), .A(n6625), .B(n6624), .ZN(n6627)
         );
  AOI21_X1 U8476 ( .B1(n9827), .B2(n6628), .A(n6627), .ZN(n6629) );
  INV_X1 U8477 ( .A(n6629), .ZN(P1_U3252) );
  AND2_X1 U8478 ( .A1(n6569), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8479 ( .A1(n6569), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8480 ( .A1(n6569), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8481 ( .A1(n6569), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8482 ( .A1(n6569), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8483 ( .A1(n6569), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8484 ( .A1(n6569), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8485 ( .A1(n6569), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8486 ( .A1(n6569), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8487 ( .A1(n6569), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8488 ( .A1(n6569), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8489 ( .A1(n6569), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8490 ( .A1(n6569), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8491 ( .A1(n6569), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8492 ( .A1(n6569), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8493 ( .A1(n6569), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8494 ( .A1(n6569), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  INV_X1 U8495 ( .A(n6630), .ZN(n6633) );
  OAI222_X1 U8496 ( .A1(n7750), .A2(n6633), .B1(n6632), .B2(P2_U3151), .C1(
        n6631), .C2(n7747), .ZN(P2_U3283) );
  INV_X1 U8497 ( .A(n9264), .ZN(n6875) );
  OAI222_X1 U8498 ( .A1(n7993), .A2(n6634), .B1(P1_U3086), .B2(n6875), .C1(
        n6633), .C2(n9658), .ZN(P1_U3343) );
  INV_X1 U8499 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6637) );
  INV_X1 U8500 ( .A(n6635), .ZN(n6638) );
  OAI222_X1 U8501 ( .A1(n7747), .A2(n6637), .B1(n7750), .B2(n6638), .C1(
        P2_U3151), .C2(n6636), .ZN(P2_U3282) );
  INV_X1 U8502 ( .A(n9796), .ZN(n9256) );
  OAI222_X1 U8503 ( .A1(n9256), .A2(P1_U3086), .B1(n9658), .B2(n6638), .C1(
        n4395), .C2(n7993), .ZN(P1_U3342) );
  INV_X1 U8504 ( .A(n6639), .ZN(n6663) );
  AOI22_X1 U8505 ( .A1(n9808), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n6673), .ZN(n6640) );
  OAI21_X1 U8506 ( .B1(n6663), .B2(n9658), .A(n6640), .ZN(P1_U3341) );
  NAND2_X1 U8507 ( .A1(n8253), .A2(P2_U3893), .ZN(n6641) );
  OAI21_X1 U8508 ( .B1(P2_U3893), .B2(n5493), .A(n6641), .ZN(P2_U3513) );
  INV_X1 U8509 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U8510 ( .A1(n8369), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U8511 ( .A1(n6642), .A2(n8357), .ZN(n6645) );
  OAI21_X1 U8512 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6643), .A(n6681), .ZN(n6644) );
  AOI22_X1 U8513 ( .A1(n6645), .A2(n6644), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6646) );
  OAI211_X1 U8514 ( .C1(n10021), .C2(n6648), .A(n6647), .B(n6646), .ZN(
        P2_U3182) );
  INV_X1 U8515 ( .A(n6649), .ZN(n6651) );
  INV_X1 U8516 ( .A(n9298), .ZN(n9287) );
  OAI222_X1 U8517 ( .A1(n7993), .A2(n6650), .B1(n9658), .B2(n6651), .C1(n9287), 
        .C2(P1_U3086), .ZN(P1_U3338) );
  OAI222_X1 U8518 ( .A1(n7747), .A2(n6652), .B1(n7750), .B2(n6651), .C1(
        P2_U3151), .C2(n4364), .ZN(P2_U3278) );
  INV_X1 U8519 ( .A(n6653), .ZN(n6656) );
  INV_X1 U8520 ( .A(n9281), .ZN(n9277) );
  OAI222_X1 U8521 ( .A1(n7993), .A2(n6654), .B1(n9658), .B2(n6656), .C1(n9277), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  OAI222_X1 U8522 ( .A1(n7747), .A2(n6657), .B1(n7750), .B2(n6656), .C1(
        P2_U3151), .C2(n6655), .ZN(P2_U3279) );
  AND2_X1 U8523 ( .A1(n9212), .A2(n6891), .ZN(n9116) );
  NOR2_X1 U8524 ( .A1(n6907), .A2(n9116), .ZN(n8922) );
  INV_X1 U8525 ( .A(n8922), .ZN(n6658) );
  OAI21_X1 U8526 ( .B1(n9971), .B2(n9882), .A(n6658), .ZN(n6659) );
  NAND2_X1 U8527 ( .A1(n9210), .A2(n9431), .ZN(n6884) );
  OAI211_X1 U8528 ( .C1(n6660), .C2(n6891), .A(n6659), .B(n6884), .ZN(n6694)
         );
  NAND2_X1 U8529 ( .A1(n6694), .A2(n9983), .ZN(n6661) );
  OAI21_X1 U8530 ( .B1(n9983), .B2(n5069), .A(n6661), .ZN(P1_U3453) );
  OAI222_X1 U8531 ( .A1(n7747), .A2(n6664), .B1(n7750), .B2(n6663), .C1(
        P2_U3151), .C2(n6662), .ZN(P2_U3281) );
  INV_X1 U8532 ( .A(n6665), .ZN(n6671) );
  OAI222_X1 U8533 ( .A1(n7750), .A2(n6671), .B1(n6667), .B2(P2_U3151), .C1(
        n6666), .C2(n7747), .ZN(P2_U3280) );
  NAND2_X1 U8534 ( .A1(n9065), .A2(P1_U3973), .ZN(n6668) );
  OAI21_X1 U8535 ( .B1(P1_U3973), .B2(n5513), .A(n6668), .ZN(P1_U3577) );
  NAND2_X1 U8536 ( .A1(n8475), .A2(P2_U3893), .ZN(n6669) );
  OAI21_X1 U8537 ( .B1(P2_U3893), .B2(n7150), .A(n6669), .ZN(P2_U3514) );
  INV_X1 U8538 ( .A(n9819), .ZN(n9265) );
  OAI222_X1 U8539 ( .A1(P1_U3086), .A2(n9265), .B1(n9658), .B2(n6671), .C1(
        n6670), .C2(n7993), .ZN(P1_U3340) );
  INV_X1 U8540 ( .A(n6672), .ZN(n6692) );
  AOI22_X1 U8541 ( .A1(n9834), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n6673), .ZN(n6674) );
  OAI21_X1 U8542 ( .B1(n6692), .B2(n9658), .A(n6674), .ZN(P1_U3337) );
  NAND2_X1 U8543 ( .A1(n6676), .A2(n6675), .ZN(n6677) );
  AOI21_X1 U8544 ( .B1(n6678), .B2(n6677), .A(n9999), .ZN(n6689) );
  XOR2_X1 U8545 ( .A(n10097), .B(n6679), .Z(n6684) );
  INV_X1 U8546 ( .A(n8357), .ZN(n10006) );
  OAI211_X1 U8547 ( .C1(n6682), .C2(n6681), .A(n6680), .B(n10006), .ZN(n6683)
         );
  OAI21_X1 U8548 ( .B1(n10014), .B2(n6684), .A(n6683), .ZN(n6688) );
  INV_X1 U8549 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6686) );
  INV_X1 U8550 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6685) );
  OAI22_X1 U8551 ( .A1(n10021), .A2(n6686), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6685), .ZN(n6687) );
  NOR3_X1 U8552 ( .A1(n6689), .A2(n6688), .A3(n6687), .ZN(n6690) );
  OAI21_X1 U8553 ( .B1(n6691), .B2(n5954), .A(n6690), .ZN(P2_U3183) );
  OAI222_X1 U8554 ( .A1(n7747), .A2(n6693), .B1(n7757), .B2(P2_U3151), .C1(
        n7750), .C2(n6692), .ZN(P2_U3277) );
  NAND2_X1 U8555 ( .A1(n6694), .A2(n9998), .ZN(n6695) );
  OAI21_X1 U8556 ( .B1(n9998), .B2(n5081), .A(n6695), .ZN(P1_U3522) );
  NAND2_X1 U8557 ( .A1(n8348), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6696) );
  OAI21_X1 U8558 ( .B1(n8455), .B2(n8348), .A(n6696), .ZN(P2_U3516) );
  OAI211_X1 U8559 ( .C1(n6699), .C2(n6698), .A(n6697), .B(n10006), .ZN(n6717)
         );
  INV_X1 U8560 ( .A(n6700), .ZN(n6702) );
  NAND3_X1 U8561 ( .A1(n6742), .A2(n6702), .A3(n6701), .ZN(n6703) );
  AOI21_X1 U8562 ( .B1(n6704), .B2(n6703), .A(n10014), .ZN(n6715) );
  INV_X1 U8563 ( .A(n6705), .ZN(n6707) );
  NAND3_X1 U8564 ( .A1(n6745), .A2(n6707), .A3(n6706), .ZN(n6708) );
  AOI21_X1 U8565 ( .B1(n6709), .B2(n6708), .A(n9999), .ZN(n6714) );
  INV_X1 U8566 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6712) );
  INV_X1 U8567 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6710) );
  NOR2_X1 U8568 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6710), .ZN(n7017) );
  INV_X1 U8569 ( .A(n7017), .ZN(n6711) );
  OAI21_X1 U8570 ( .B1(n10021), .B2(n6712), .A(n6711), .ZN(n6713) );
  NOR3_X1 U8571 ( .A1(n6715), .A2(n6714), .A3(n6713), .ZN(n6716) );
  OAI211_X1 U8572 ( .C1(n5954), .C2(n6718), .A(n6717), .B(n6716), .ZN(P2_U3186) );
  AOI21_X1 U8573 ( .B1(n6721), .B2(n6720), .A(n6719), .ZN(n6736) );
  AOI21_X1 U8574 ( .B1(n6723), .B2(n6722), .A(n4354), .ZN(n6728) );
  INV_X1 U8575 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6724) );
  NOR2_X1 U8576 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6724), .ZN(n7033) );
  INV_X1 U8577 ( .A(n7033), .ZN(n6727) );
  INV_X1 U8578 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6725) );
  OR2_X1 U8579 ( .A1(n10021), .A2(n6725), .ZN(n6726) );
  OAI211_X1 U8580 ( .C1(n6728), .C2(n10014), .A(n6727), .B(n6726), .ZN(n6733)
         );
  AOI21_X1 U8581 ( .B1(n4353), .B2(n6730), .A(n6729), .ZN(n6731) );
  NOR2_X1 U8582 ( .A1(n9999), .A2(n6731), .ZN(n6732) );
  AOI211_X1 U8583 ( .C1(n8369), .C2(n6734), .A(n6733), .B(n6732), .ZN(n6735)
         );
  OAI21_X1 U8584 ( .B1(n6736), .B2(n8357), .A(n6735), .ZN(P2_U3188) );
  AOI21_X1 U8585 ( .B1(n6739), .B2(n6738), .A(n6737), .ZN(n6754) );
  INV_X1 U8586 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6741) );
  NOR2_X1 U8587 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7201), .ZN(n6803) );
  INV_X1 U8588 ( .A(n6803), .ZN(n6740) );
  OAI21_X1 U8589 ( .B1(n10021), .B2(n6741), .A(n6740), .ZN(n6751) );
  INV_X1 U8590 ( .A(n6742), .ZN(n6743) );
  AOI21_X1 U8591 ( .B1(n10101), .B2(n6744), .A(n6743), .ZN(n6749) );
  INV_X1 U8592 ( .A(n6745), .ZN(n6746) );
  AOI21_X1 U8593 ( .B1(n7204), .B2(n6747), .A(n6746), .ZN(n6748) );
  OAI22_X1 U8594 ( .A1(n6749), .A2(n10014), .B1(n9999), .B2(n6748), .ZN(n6750)
         );
  AOI211_X1 U8595 ( .C1(n6752), .C2(n8369), .A(n6751), .B(n6750), .ZN(n6753)
         );
  OAI21_X1 U8596 ( .B1(n6754), .B2(n8357), .A(n6753), .ZN(P2_U3185) );
  OAI211_X1 U8597 ( .C1(n6757), .C2(n6756), .A(n6755), .B(n10006), .ZN(n6768)
         );
  AND2_X1 U8598 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7004) );
  AOI21_X1 U8599 ( .B1(n6759), .B2(n10105), .A(n6758), .ZN(n6764) );
  AOI21_X1 U8600 ( .B1(n6762), .B2(n6761), .A(n6760), .ZN(n6763) );
  OAI22_X1 U8601 ( .A1(n6764), .A2(n10014), .B1(n9999), .B2(n6763), .ZN(n6765)
         );
  AOI211_X1 U8602 ( .C1(n6766), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7004), .B(
        n6765), .ZN(n6767) );
  OAI211_X1 U8603 ( .C1(n5954), .C2(n6769), .A(n6768), .B(n6767), .ZN(P2_U3187) );
  AOI21_X1 U8604 ( .B1(n6772), .B2(n6771), .A(n6770), .ZN(n6778) );
  INV_X1 U8605 ( .A(n6773), .ZN(n9209) );
  NAND2_X1 U8606 ( .A1(n9209), .A2(n9431), .ZN(n6775) );
  NAND2_X1 U8607 ( .A1(n9210), .A2(n9433), .ZN(n6774) );
  NAND2_X1 U8608 ( .A1(n6775), .A2(n6774), .ZN(n6982) );
  AOI22_X1 U8609 ( .A1(n8887), .A2(n6989), .B1(n6982), .B2(n8888), .ZN(n6777)
         );
  NAND2_X1 U8610 ( .A1(n8893), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6894) );
  NAND2_X1 U8611 ( .A1(n6894), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6776) );
  OAI211_X1 U8612 ( .C1(n6778), .C2(n5697), .A(n6777), .B(n6776), .ZN(P1_U3237) );
  INV_X1 U8613 ( .A(n6790), .ZN(n6783) );
  NAND3_X1 U8614 ( .A1(n6781), .A2(n6780), .A3(n6779), .ZN(n6782) );
  NOR2_X1 U8615 ( .A1(n6794), .A2(n6788), .ZN(n6792) );
  AOI211_X1 U8616 ( .C1(n6784), .C2(n6783), .A(n6782), .B(n6792), .ZN(n6785)
         );
  OAI22_X1 U8617 ( .A1(n6785), .A2(P2_U3151), .B1(n6794), .B2(n8225), .ZN(
        n8326) );
  INV_X1 U8618 ( .A(n8326), .ZN(n7003) );
  NAND2_X1 U8619 ( .A1(n7003), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6850) );
  INV_X1 U8620 ( .A(n6850), .ZN(n6800) );
  INV_X1 U8621 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6930) );
  OR2_X1 U8622 ( .A1(n6790), .A2(n8445), .ZN(n6787) );
  AND2_X1 U8623 ( .A1(n6787), .A2(n6786), .ZN(n7021) );
  NAND2_X1 U8624 ( .A1(n7021), .A2(n10028), .ZN(n8323) );
  INV_X1 U8625 ( .A(n8323), .ZN(n6798) );
  INV_X1 U8626 ( .A(n10027), .ZN(n6931) );
  NAND2_X1 U8627 ( .A1(n8349), .A2(n6931), .ZN(n8045) );
  AND2_X1 U8628 ( .A1(n8036), .A2(n8045), .ZN(n10023) );
  INV_X1 U8629 ( .A(n6788), .ZN(n6789) );
  AOI21_X1 U8630 ( .B1(n6791), .B2(n6790), .A(n6789), .ZN(n6793) );
  INV_X1 U8631 ( .A(n6794), .ZN(n6795) );
  INV_X1 U8632 ( .A(n8389), .ZN(n6796) );
  OAI22_X1 U8633 ( .A1(n10023), .A2(n8328), .B1(n8299), .B2(n7108), .ZN(n6797)
         );
  AOI21_X1 U8634 ( .B1(n10027), .B2(n6798), .A(n6797), .ZN(n6799) );
  OAI21_X1 U8635 ( .B1(n6800), .B2(n6930), .A(n6799), .ZN(P2_U3172) );
  NOR2_X1 U8636 ( .A1(n8048), .A2(n10068), .ZN(n10041) );
  NOR2_X2 U8637 ( .A1(n6801), .A2(n8389), .ZN(n8297) );
  OAI22_X1 U8638 ( .A1(n8322), .A2(n6848), .B1(n7000), .B2(n8299), .ZN(n6802)
         );
  AOI211_X1 U8639 ( .C1(n7021), .C2(n10041), .A(n6803), .B(n6802), .ZN(n6818)
         );
  OAI21_X1 U8640 ( .B1(n6804), .B2(n8221), .A(n8183), .ZN(n6805) );
  XNOR2_X1 U8641 ( .A(n6813), .B(n7223), .ZN(n6809) );
  XNOR2_X1 U8642 ( .A(n6809), .B(n7108), .ZN(n6846) );
  OR2_X1 U8643 ( .A1(n6813), .A2(n10027), .ZN(n6808) );
  AND2_X1 U8644 ( .A1(n8036), .A2(n6808), .ZN(n6845) );
  NAND2_X1 U8645 ( .A1(n6809), .A2(n7108), .ZN(n6810) );
  XNOR2_X1 U8646 ( .A(n6813), .B(n8049), .ZN(n6811) );
  XNOR2_X1 U8647 ( .A(n6811), .B(n6848), .ZN(n6839) );
  NOR2_X1 U8648 ( .A1(n6811), .A2(n8346), .ZN(n6812) );
  INV_X2 U8649 ( .A(n6813), .ZN(n6814) );
  INV_X8 U8650 ( .A(n6814), .ZN(n7974) );
  XNOR2_X1 U8651 ( .A(n7974), .B(n8048), .ZN(n6995) );
  XNOR2_X1 U8652 ( .A(n6995), .B(n7109), .ZN(n6815) );
  INV_X1 U8653 ( .A(n8328), .ZN(n8283) );
  OAI211_X1 U8654 ( .C1(n6816), .C2(n6815), .A(n6997), .B(n8283), .ZN(n6817)
         );
  OAI211_X1 U8655 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7003), .A(n6818), .B(
        n6817), .ZN(P2_U3158) );
  OAI21_X1 U8656 ( .B1(n6821), .B2(n6820), .A(n6819), .ZN(n6896) );
  INV_X1 U8657 ( .A(n6896), .ZN(n6822) );
  MUX2_X1 U8658 ( .A(n6823), .B(n6822), .S(n9728), .Z(n6825) );
  NOR2_X1 U8659 ( .A1(n9728), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6824) );
  OR2_X1 U8660 ( .A1(n7620), .A2(n6824), .ZN(n9727) );
  NAND2_X1 U8661 ( .A1(n9727), .A2(n9730), .ZN(n9733) );
  OAI211_X1 U8662 ( .C1(n6825), .C2(n7620), .A(P1_U3973), .B(n9733), .ZN(n9252) );
  INV_X1 U8663 ( .A(n9252), .ZN(n6838) );
  OAI211_X1 U8664 ( .C1(n6828), .C2(n6827), .A(n9827), .B(n6826), .ZN(n6836)
         );
  OAI211_X1 U8665 ( .C1(n6831), .C2(n6830), .A(n9778), .B(n6829), .ZN(n6835)
         );
  AOI22_X1 U8666 ( .A1(n9735), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6834) );
  INV_X1 U8667 ( .A(n9782), .ZN(n9835) );
  NAND2_X1 U8668 ( .A1(n9835), .A2(n6832), .ZN(n6833) );
  NAND4_X1 U8669 ( .A1(n6836), .A2(n6835), .A3(n6834), .A4(n6833), .ZN(n6837)
         );
  OR2_X1 U8670 ( .A1(n6838), .A2(n6837), .ZN(P1_U3245) );
  XOR2_X1 U8671 ( .A(n6840), .B(n6839), .Z(n6844) );
  NOR2_X1 U8672 ( .A1(n8049), .A2(n10068), .ZN(n10036) );
  AOI22_X1 U8673 ( .A1(n8297), .A2(n8347), .B1(n10036), .B2(n7021), .ZN(n6841)
         );
  OAI21_X1 U8674 ( .B1(n7109), .B2(n8299), .A(n6841), .ZN(n6842) );
  AOI21_X1 U8675 ( .B1(n6850), .B2(P2_REG3_REG_2__SCAN_IN), .A(n6842), .ZN(
        n6843) );
  OAI21_X1 U8676 ( .B1(n6844), .B2(n8328), .A(n6843), .ZN(P2_U3177) );
  XOR2_X1 U8677 ( .A(n6846), .B(n6845), .Z(n6852) );
  AND2_X1 U8678 ( .A1(n7223), .A2(n10028), .ZN(n10031) );
  AOI22_X1 U8679 ( .A1(n8297), .A2(n8349), .B1(n10031), .B2(n7021), .ZN(n6847)
         );
  OAI21_X1 U8680 ( .B1(n6848), .B2(n8299), .A(n6847), .ZN(n6849) );
  AOI21_X1 U8681 ( .B1(n6850), .B2(P2_REG3_REG_1__SCAN_IN), .A(n6849), .ZN(
        n6851) );
  OAI21_X1 U8682 ( .B1(n8328), .B2(n6852), .A(n6851), .ZN(P2_U3162) );
  AOI21_X1 U8683 ( .B1(n6855), .B2(n6854), .A(n6853), .ZN(n6860) );
  INV_X1 U8684 ( .A(n8832), .ZN(n8876) );
  AOI22_X1 U8685 ( .A1(n6903), .A2(n8887), .B1(n8813), .B2(n6010), .ZN(n6856)
         );
  OAI21_X1 U8686 ( .B1(n6857), .B2(n8876), .A(n6856), .ZN(n6858) );
  AOI21_X1 U8687 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n6894), .A(n6858), .ZN(
        n6859) );
  OAI21_X1 U8688 ( .B1(n6860), .B2(n5697), .A(n6859), .ZN(P1_U3222) );
  NOR2_X1 U8689 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9264), .ZN(n6861) );
  AOI21_X1 U8690 ( .B1(n9264), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6861), .ZN(
        n6866) );
  NAND2_X1 U8691 ( .A1(n9669), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6862) );
  OAI21_X1 U8692 ( .B1(n9669), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6862), .ZN(
        n9665) );
  NOR2_X1 U8693 ( .A1(n9665), .A2(n9666), .ZN(n9664) );
  NAND2_X1 U8694 ( .A1(n9769), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6864) );
  OAI21_X1 U8695 ( .B1(n9769), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6864), .ZN(
        n9772) );
  NOR2_X1 U8696 ( .A1(n9771), .A2(n9772), .ZN(n9770) );
  AOI21_X1 U8697 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9769), .A(n9770), .ZN(
        n6865) );
  NAND2_X1 U8698 ( .A1(n6866), .A2(n6865), .ZN(n9263) );
  OAI21_X1 U8699 ( .B1(n6866), .B2(n6865), .A(n9263), .ZN(n6867) );
  NAND2_X1 U8700 ( .A1(n6867), .A2(n9827), .ZN(n6879) );
  MUX2_X1 U8701 ( .A(n6868), .B(P1_REG1_REG_10__SCAN_IN), .S(n9669), .Z(n9662)
         );
  OAI21_X1 U8702 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n6870), .A(n6869), .ZN(
        n9663) );
  NOR2_X1 U8703 ( .A1(n9662), .A2(n9663), .ZN(n9661) );
  AOI21_X1 U8704 ( .B1(n9669), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9661), .ZN(
        n9775) );
  MUX2_X1 U8705 ( .A(n6871), .B(P1_REG1_REG_11__SCAN_IN), .S(n9769), .Z(n9776)
         );
  NOR2_X1 U8706 ( .A1(n9775), .A2(n9776), .ZN(n9774) );
  AOI21_X1 U8707 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9769), .A(n9774), .ZN(
        n6873) );
  AOI22_X1 U8708 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n9264), .B1(n6875), .B2(
        n5279), .ZN(n6872) );
  NAND2_X1 U8709 ( .A1(n6873), .A2(n6872), .ZN(n9257) );
  OAI21_X1 U8710 ( .B1(n6873), .B2(n6872), .A(n9257), .ZN(n6877) );
  NAND2_X1 U8711 ( .A1(n9735), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6874) );
  NAND2_X1 U8712 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7520) );
  OAI211_X1 U8713 ( .C1(n9782), .C2(n6875), .A(n6874), .B(n7520), .ZN(n6876)
         );
  AOI21_X1 U8714 ( .B1(n6877), .B2(n9778), .A(n6876), .ZN(n6878) );
  NAND2_X1 U8715 ( .A1(n6879), .A2(n6878), .ZN(P1_U3255) );
  NAND3_X1 U8716 ( .A1(n6882), .A2(n6881), .A3(n6880), .ZN(n6888) );
  INV_X1 U8717 ( .A(n9523), .ZN(n9528) );
  INV_X1 U8718 ( .A(n9501), .ZN(n9886) );
  NAND2_X1 U8719 ( .A1(n9886), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6883) );
  OAI211_X1 U8720 ( .C1(n8922), .C2(n6885), .A(n6884), .B(n6883), .ZN(n6886)
         );
  INV_X1 U8721 ( .A(n9523), .ZN(n9346) );
  NAND2_X1 U8722 ( .A1(n6886), .A2(n9346), .ZN(n6890) );
  OR2_X1 U8723 ( .A1(n6888), .A2(n9308), .ZN(n9351) );
  NOR2_X1 U8724 ( .A1(n9351), .A2(n9909), .ZN(n6905) );
  OAI21_X1 U8725 ( .B1(n9884), .B2(n6905), .A(n6904), .ZN(n6889) );
  OAI211_X1 U8726 ( .C1(n5071), .C2(n9528), .A(n6890), .B(n6889), .ZN(P1_U3293) );
  OAI22_X1 U8727 ( .A1(n8877), .A2(n6892), .B1(n8883), .B2(n6891), .ZN(n6893)
         );
  AOI21_X1 U8728 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6894), .A(n6893), .ZN(
        n6895) );
  OAI21_X1 U8729 ( .B1(n6896), .B2(n5697), .A(n6895), .ZN(P1_U3232) );
  NAND2_X1 U8730 ( .A1(n8348), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6897) );
  OAI21_X1 U8731 ( .B1(n8004), .B2(n8348), .A(n6897), .ZN(P2_U3521) );
  INV_X1 U8732 ( .A(n6898), .ZN(n6950) );
  OAI222_X1 U8733 ( .A1(n7747), .A2(n6899), .B1(n7750), .B2(n6950), .C1(n8221), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  NAND2_X1 U8734 ( .A1(n8348), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6900) );
  OAI21_X1 U8735 ( .B1(n8015), .B2(n8348), .A(n6900), .ZN(P2_U3520) );
  XNOR2_X1 U8736 ( .A(n6908), .B(n6901), .ZN(n9913) );
  NOR2_X1 U8737 ( .A1(n9900), .A2(n6937), .ZN(n9862) );
  INV_X1 U8738 ( .A(n6986), .ZN(n6902) );
  AOI21_X1 U8739 ( .B1(n6904), .B2(n6903), .A(n6902), .ZN(n9908) );
  AOI22_X1 U8740 ( .A1(n9908), .A2(n6905), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9886), .ZN(n6906) );
  XNOR2_X1 U8741 ( .A(n6908), .B(n6907), .ZN(n6911) );
  INV_X1 U8742 ( .A(n9882), .ZN(n9465) );
  INV_X1 U8743 ( .A(n9851), .ZN(n9981) );
  NAND2_X1 U8744 ( .A1(n9913), .A2(n9981), .ZN(n6910) );
  AOI22_X1 U8745 ( .A1(n6010), .A2(n9431), .B1(n9433), .B2(n9212), .ZN(n6909)
         );
  OAI211_X1 U8746 ( .C1(n6911), .C2(n9465), .A(n6910), .B(n6909), .ZN(n9911)
         );
  MUX2_X1 U8747 ( .A(n9911), .B(P1_REG2_REG_1__SCAN_IN), .S(n9523), .Z(n6912)
         );
  AOI211_X1 U8748 ( .C1(n9913), .C2(n9862), .A(n6913), .B(n6912), .ZN(n6914)
         );
  INV_X1 U8749 ( .A(n6914), .ZN(P1_U3292) );
  INV_X1 U8750 ( .A(n6915), .ZN(n6918) );
  OAI222_X1 U8751 ( .A1(n8777), .A2(n6918), .B1(P2_U3151), .B2(n8183), .C1(
        n6916), .C2(n7747), .ZN(P2_U3275) );
  OAI222_X1 U8752 ( .A1(n8955), .A2(P1_U3086), .B1(n9658), .B2(n6918), .C1(
        n6917), .C2(n7993), .ZN(P1_U3335) );
  NAND2_X1 U8753 ( .A1(n9211), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6919) );
  OAI21_X1 U8754 ( .B1(n9339), .B2(n9211), .A(n6919), .ZN(P1_U3583) );
  INV_X1 U8755 ( .A(n6920), .ZN(n6924) );
  NOR2_X1 U8756 ( .A1(n6922), .A2(n6921), .ZN(n6923) );
  NAND2_X1 U8757 ( .A1(n6924), .A2(n6923), .ZN(n6929) );
  NAND2_X2 U8758 ( .A1(n6929), .A2(n9703), .ZN(n9716) );
  NOR3_X1 U8759 ( .A1(n10023), .A2(n6927), .A3(n10028), .ZN(n6928) );
  NOR2_X1 U8760 ( .A1(n7108), .A2(n9712), .ZN(n10026) );
  OAI21_X1 U8761 ( .B1(n6928), .B2(n10026), .A(n9716), .ZN(n6934) );
  OAI22_X1 U8762 ( .A1(n8523), .A2(n6931), .B1(n6930), .B2(n9703), .ZN(n6932)
         );
  INV_X1 U8763 ( .A(n6932), .ZN(n6933) );
  OAI211_X1 U8764 ( .C1(n6935), .C2(n9716), .A(n6934), .B(n6933), .ZN(P2_U3233) );
  XNOR2_X1 U8765 ( .A(n6936), .B(n4291), .ZN(n9930) );
  AND2_X1 U8766 ( .A1(n9851), .A2(n6937), .ZN(n6938) );
  XNOR2_X1 U8767 ( .A(n8964), .B(n4291), .ZN(n6940) );
  AOI22_X1 U8768 ( .A1(n9431), .A2(n9207), .B1(n9209), .B2(n9433), .ZN(n7089)
         );
  INV_X1 U8769 ( .A(n7089), .ZN(n6939) );
  AOI21_X1 U8770 ( .B1(n6940), .B2(n9882), .A(n6939), .ZN(n9929) );
  MUX2_X1 U8771 ( .A(n9929), .B(n6941), .S(n9523), .Z(n6946) );
  INV_X1 U8772 ( .A(n6942), .ZN(n9875) );
  AOI211_X1 U8773 ( .C1(n9927), .C2(n9893), .A(n9909), .B(n9875), .ZN(n9926)
         );
  OAI22_X1 U8774 ( .A1(n9526), .A2(n6943), .B1(n9501), .B2(n7093), .ZN(n6944)
         );
  AOI21_X1 U8775 ( .B1(n9926), .B2(n9896), .A(n6944), .ZN(n6945) );
  OAI211_X1 U8776 ( .C1(n9930), .C2(n9530), .A(n6946), .B(n6945), .ZN(P1_U3289) );
  INV_X1 U8777 ( .A(n6947), .ZN(n6957) );
  OAI222_X1 U8778 ( .A1(n7750), .A2(n6957), .B1(P2_U3151), .B2(n8011), .C1(
        n6948), .C2(n7747), .ZN(P2_U3274) );
  OAI222_X1 U8779 ( .A1(P1_U3086), .A2(n9410), .B1(n9658), .B2(n6950), .C1(
        n6949), .C2(n7993), .ZN(P1_U3336) );
  XOR2_X1 U8780 ( .A(n6952), .B(n6951), .Z(n6955) );
  INV_X1 U8781 ( .A(n9431), .ZN(n9467) );
  INV_X1 U8782 ( .A(n9433), .ZN(n9469) );
  OAI22_X1 U8783 ( .A1(n7209), .A2(n9467), .B1(n6011), .B2(n9469), .ZN(n9881)
         );
  AOI22_X1 U8784 ( .A1(n9881), .A2(n8888), .B1(n9885), .B2(n8887), .ZN(n6954)
         );
  INV_X1 U8785 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9887) );
  MUX2_X1 U8786 ( .A(P1_STATE_REG_SCAN_IN), .B(n8862), .S(n9887), .Z(n6953) );
  OAI211_X1 U8787 ( .C1(n6955), .C2(n5697), .A(n6954), .B(n6953), .ZN(P1_U3218) );
  OAI222_X1 U8788 ( .A1(n9118), .A2(P1_U3086), .B1(n9658), .B2(n6957), .C1(
        n6956), .C2(n7993), .ZN(P1_U3334) );
  AOI21_X1 U8789 ( .B1(n10113), .B2(n6959), .A(n6958), .ZN(n6976) );
  INV_X1 U8790 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6961) );
  AND2_X1 U8791 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7142) );
  INV_X1 U8792 ( .A(n7142), .ZN(n6960) );
  OAI21_X1 U8793 ( .B1(n10021), .B2(n6961), .A(n6960), .ZN(n6967) );
  AOI21_X1 U8794 ( .B1(n6964), .B2(n6963), .A(n6962), .ZN(n6965) );
  NOR2_X1 U8795 ( .A1(n6965), .A2(n9999), .ZN(n6966) );
  AOI211_X1 U8796 ( .C1(n8369), .C2(n6968), .A(n6967), .B(n6966), .ZN(n6975)
         );
  NOR2_X1 U8797 ( .A1(n6970), .A2(n6969), .ZN(n6972) );
  XNOR2_X1 U8798 ( .A(n6972), .B(n6971), .ZN(n6973) );
  NAND2_X1 U8799 ( .A1(n6973), .A2(n10006), .ZN(n6974) );
  OAI211_X1 U8800 ( .C1(n6976), .C2(n10014), .A(n6975), .B(n6974), .ZN(
        P2_U3191) );
  XNOR2_X1 U8801 ( .A(n6978), .B(n6977), .ZN(n9914) );
  NAND2_X1 U8802 ( .A1(n9914), .A2(n9981), .ZN(n6985) );
  XNOR2_X1 U8803 ( .A(n6980), .B(n6977), .ZN(n6981) );
  NAND2_X1 U8804 ( .A1(n6981), .A2(n9882), .ZN(n6984) );
  INV_X1 U8805 ( .A(n6982), .ZN(n6983) );
  NAND3_X1 U8806 ( .A1(n6985), .A2(n6984), .A3(n6983), .ZN(n9919) );
  INV_X1 U8807 ( .A(n9919), .ZN(n6994) );
  NAND2_X1 U8808 ( .A1(n6986), .A2(n6989), .ZN(n6987) );
  NAND2_X1 U8809 ( .A1(n6987), .A2(n9892), .ZN(n6988) );
  OR2_X1 U8810 ( .A1(n6988), .A2(n9894), .ZN(n9915) );
  AOI22_X1 U8811 ( .A1(n9523), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9886), .ZN(n6991) );
  NAND2_X1 U8812 ( .A1(n9884), .A2(n6989), .ZN(n6990) );
  OAI211_X1 U8813 ( .C1(n9915), .C2(n9351), .A(n6991), .B(n6990), .ZN(n6992)
         );
  AOI21_X1 U8814 ( .B1(n9914), .B2(n9862), .A(n6992), .ZN(n6993) );
  OAI21_X1 U8815 ( .B1(n6994), .B2(n9523), .A(n6993), .ZN(P1_U3291) );
  NAND2_X1 U8816 ( .A1(n6995), .A2(n8345), .ZN(n6996) );
  XNOR2_X1 U8817 ( .A(n7974), .B(n7015), .ZN(n6999) );
  XNOR2_X1 U8818 ( .A(n6999), .B(n8344), .ZN(n7014) );
  INV_X1 U8819 ( .A(n6999), .ZN(n7001) );
  NAND2_X1 U8820 ( .A1(n7001), .A2(n7000), .ZN(n7002) );
  NAND2_X1 U8821 ( .A1(n7011), .A2(n7002), .ZN(n7023) );
  XNOR2_X1 U8822 ( .A(n7974), .B(n7005), .ZN(n7024) );
  XNOR2_X1 U8823 ( .A(n7024), .B(n7025), .ZN(n7022) );
  XOR2_X1 U8824 ( .A(n7023), .B(n7022), .Z(n7010) );
  AOI21_X1 U8825 ( .B1(n8297), .B2(n8344), .A(n7004), .ZN(n7007) );
  NOR2_X1 U8826 ( .A1(n7005), .A2(n10068), .ZN(n10049) );
  NAND2_X1 U8827 ( .A1(n7021), .A2(n10049), .ZN(n7006) );
  OAI211_X1 U8828 ( .C1(n7154), .C2(n8299), .A(n7007), .B(n7006), .ZN(n7008)
         );
  AOI21_X1 U8829 ( .B1(n8291), .B2(n7125), .A(n7008), .ZN(n7009) );
  OAI21_X1 U8830 ( .B1(n7010), .B2(n8328), .A(n7009), .ZN(P2_U3167) );
  INV_X1 U8831 ( .A(n7011), .ZN(n7012) );
  AOI21_X1 U8832 ( .B1(n7014), .B2(n7013), .A(n7012), .ZN(n7020) );
  NOR2_X1 U8833 ( .A1(n7015), .A2(n10068), .ZN(n10045) );
  OAI22_X1 U8834 ( .A1(n8322), .A2(n7109), .B1(n7025), .B2(n8299), .ZN(n7016)
         );
  AOI211_X1 U8835 ( .C1(n7021), .C2(n10045), .A(n7017), .B(n7016), .ZN(n7019)
         );
  NAND2_X1 U8836 ( .A1(n8291), .A2(n7192), .ZN(n7018) );
  OAI211_X1 U8837 ( .C1(n7020), .C2(n8328), .A(n7019), .B(n7018), .ZN(P2_U3170) );
  INV_X1 U8838 ( .A(n7021), .ZN(n8313) );
  NAND2_X1 U8839 ( .A1(n7268), .A2(n10028), .ZN(n10053) );
  NAND2_X1 U8840 ( .A1(n7023), .A2(n7022), .ZN(n7028) );
  INV_X1 U8841 ( .A(n7024), .ZN(n7026) );
  NAND2_X1 U8842 ( .A1(n7026), .A2(n7025), .ZN(n7027) );
  NAND2_X1 U8843 ( .A1(n7028), .A2(n7027), .ZN(n7029) );
  XNOR2_X1 U8844 ( .A(n7974), .B(n7268), .ZN(n7038) );
  XNOR2_X1 U8845 ( .A(n7038), .B(n7154), .ZN(n7030) );
  AOI21_X1 U8846 ( .B1(n7029), .B2(n7030), .A(n8328), .ZN(n7032) );
  NAND2_X1 U8847 ( .A1(n7032), .A2(n7041), .ZN(n7037) );
  AOI21_X1 U8848 ( .B1(n8297), .B2(n8343), .A(n7033), .ZN(n7034) );
  OAI21_X1 U8849 ( .B1(n6222), .B2(n8299), .A(n7034), .ZN(n7035) );
  AOI21_X1 U8850 ( .B1(n8291), .B2(n7267), .A(n7035), .ZN(n7036) );
  OAI211_X1 U8851 ( .C1(n8313), .C2(n10053), .A(n7037), .B(n7036), .ZN(
        P2_U3179) );
  AND2_X1 U8852 ( .A1(n7166), .A2(n10028), .ZN(n10060) );
  INV_X1 U8853 ( .A(n10060), .ZN(n7051) );
  INV_X1 U8854 ( .A(n7038), .ZN(n7039) );
  NAND2_X1 U8855 ( .A1(n6453), .A2(n7039), .ZN(n7040) );
  XNOR2_X1 U8856 ( .A(n7042), .B(n7974), .ZN(n7094) );
  XNOR2_X1 U8857 ( .A(n7094), .B(n6222), .ZN(n7043) );
  OAI21_X1 U8858 ( .B1(n7044), .B2(n7043), .A(n7097), .ZN(n7045) );
  NAND2_X1 U8859 ( .A1(n7045), .A2(n8283), .ZN(n7050) );
  NAND2_X1 U8860 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7929) );
  INV_X1 U8861 ( .A(n7929), .ZN(n7046) );
  AOI21_X1 U8862 ( .B1(n8297), .B2(n6453), .A(n7046), .ZN(n7047) );
  OAI21_X1 U8863 ( .B1(n7442), .B2(n8299), .A(n7047), .ZN(n7048) );
  AOI21_X1 U8864 ( .B1(n8291), .B2(n7165), .A(n7048), .ZN(n7049) );
  OAI211_X1 U8865 ( .C1(n8313), .C2(n7051), .A(n7050), .B(n7049), .ZN(P2_U3153) );
  INV_X1 U8866 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10127) );
  NOR2_X1 U8867 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7052) );
  AOI21_X1 U8868 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7052), .ZN(n10133) );
  NOR2_X1 U8869 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7053) );
  AOI21_X1 U8870 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7053), .ZN(n10136) );
  INV_X1 U8871 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8361) );
  INV_X1 U8872 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U8873 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .B1(n8361), .B2(n9822), .ZN(n10139) );
  NOR2_X1 U8874 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7054) );
  AOI21_X1 U8875 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7054), .ZN(n10142) );
  INV_X1 U8876 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7837) );
  INV_X1 U8877 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U8878 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .B1(n7837), .B2(n9799), .ZN(n10145) );
  NOR2_X1 U8879 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7055) );
  AOI21_X1 U8880 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7055), .ZN(n10148) );
  NOR2_X1 U8881 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7056) );
  AOI21_X1 U8882 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7056), .ZN(n10151) );
  INV_X1 U8883 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7888) );
  INV_X1 U8884 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9672) );
  AOI22_X1 U8885 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .B1(n7888), .B2(n9672), .ZN(n10154) );
  NOR2_X1 U8886 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7057) );
  AOI21_X1 U8887 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7057), .ZN(n10163) );
  NOR2_X1 U8888 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7058) );
  AOI21_X1 U8889 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7058), .ZN(n10169) );
  NOR2_X1 U8890 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7059) );
  AOI21_X1 U8891 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7059), .ZN(n10166) );
  NOR2_X1 U8892 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7060) );
  AOI21_X1 U8893 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7060), .ZN(n10157) );
  NOR2_X1 U8894 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7061) );
  AOI21_X1 U8895 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7061), .ZN(n10160) );
  AND2_X1 U8896 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7062) );
  NOR2_X1 U8897 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7062), .ZN(n10123) );
  INV_X1 U8898 ( .A(n10123), .ZN(n10124) );
  NAND3_X1 U8899 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U8900 ( .A1(n6686), .A2(n10125), .ZN(n10122) );
  NAND2_X1 U8901 ( .A1(n10124), .A2(n10122), .ZN(n10172) );
  NAND2_X1 U8902 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7063) );
  OAI21_X1 U8903 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7063), .ZN(n10171) );
  NOR2_X1 U8904 ( .A1(n10172), .A2(n10171), .ZN(n10170) );
  AOI21_X1 U8905 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10170), .ZN(n10175) );
  NAND2_X1 U8906 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7064) );
  OAI21_X1 U8907 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7064), .ZN(n10174) );
  NOR2_X1 U8908 ( .A1(n10175), .A2(n10174), .ZN(n10173) );
  AOI21_X1 U8909 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10173), .ZN(n10178) );
  NOR2_X1 U8910 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7065) );
  AOI21_X1 U8911 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7065), .ZN(n10177) );
  NAND2_X1 U8912 ( .A1(n10178), .A2(n10177), .ZN(n10176) );
  OAI21_X1 U8913 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10176), .ZN(n10159) );
  NAND2_X1 U8914 ( .A1(n10160), .A2(n10159), .ZN(n10158) );
  OAI21_X1 U8915 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10158), .ZN(n10156) );
  NAND2_X1 U8916 ( .A1(n10157), .A2(n10156), .ZN(n10155) );
  OAI21_X1 U8917 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10155), .ZN(n10165) );
  NAND2_X1 U8918 ( .A1(n10166), .A2(n10165), .ZN(n10164) );
  OAI21_X1 U8919 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10164), .ZN(n10168) );
  NAND2_X1 U8920 ( .A1(n10169), .A2(n10168), .ZN(n10167) );
  OAI21_X1 U8921 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10167), .ZN(n10162) );
  NAND2_X1 U8922 ( .A1(n10163), .A2(n10162), .ZN(n10161) );
  OAI21_X1 U8923 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10161), .ZN(n10153) );
  NAND2_X1 U8924 ( .A1(n10154), .A2(n10153), .ZN(n10152) );
  OAI21_X1 U8925 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10152), .ZN(n10150) );
  NAND2_X1 U8926 ( .A1(n10151), .A2(n10150), .ZN(n10149) );
  OAI21_X1 U8927 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10149), .ZN(n10147) );
  NAND2_X1 U8928 ( .A1(n10148), .A2(n10147), .ZN(n10146) );
  OAI21_X1 U8929 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10146), .ZN(n10144) );
  NAND2_X1 U8930 ( .A1(n10145), .A2(n10144), .ZN(n10143) );
  OAI21_X1 U8931 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10143), .ZN(n10141) );
  NAND2_X1 U8932 ( .A1(n10142), .A2(n10141), .ZN(n10140) );
  OAI21_X1 U8933 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10140), .ZN(n10138) );
  NAND2_X1 U8934 ( .A1(n10139), .A2(n10138), .ZN(n10137) );
  OAI21_X1 U8935 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10137), .ZN(n10135) );
  NAND2_X1 U8936 ( .A1(n10136), .A2(n10135), .ZN(n10134) );
  OAI21_X1 U8937 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10134), .ZN(n10132) );
  NAND2_X1 U8938 ( .A1(n10133), .A2(n10132), .ZN(n10131) );
  OAI21_X1 U8939 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10131), .ZN(n10128) );
  NAND2_X1 U8940 ( .A1(n10127), .A2(n10128), .ZN(n7066) );
  NOR2_X1 U8941 ( .A1(n10127), .A2(n10128), .ZN(n10126) );
  AOI21_X1 U8942 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7066), .A(n10126), .ZN(
        n7068) );
  XNOR2_X1 U8943 ( .A(n9313), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7067) );
  XNOR2_X1 U8944 ( .A(n7068), .B(n7067), .ZN(ADD_1068_U4) );
  XOR2_X1 U8945 ( .A(n8973), .B(n7073), .Z(n7071) );
  OAI22_X1 U8946 ( .A1(n7070), .A2(n9469), .B1(n7069), .B2(n9467), .ZN(n7359)
         );
  AOI21_X1 U8947 ( .B1(n7071), .B2(n9882), .A(n7359), .ZN(n9941) );
  XNOR2_X1 U8948 ( .A(n7072), .B(n7073), .ZN(n9944) );
  INV_X1 U8949 ( .A(n9530), .ZN(n9897) );
  INV_X1 U8950 ( .A(n9860), .ZN(n7074) );
  OAI211_X1 U8951 ( .C1(n9940), .C2(n9873), .A(n7074), .B(n9892), .ZN(n9939)
         );
  OAI22_X1 U8952 ( .A1(n9528), .A2(n7075), .B1(n7361), .B2(n9501), .ZN(n7076)
         );
  AOI21_X1 U8953 ( .B1(n9884), .B2(n7363), .A(n7076), .ZN(n7077) );
  OAI21_X1 U8954 ( .B1(n9939), .B2(n9351), .A(n7077), .ZN(n7078) );
  AOI21_X1 U8955 ( .B1(n9944), .B2(n9897), .A(n7078), .ZN(n7079) );
  OAI21_X1 U8956 ( .B1(n9941), .B2(n9523), .A(n7079), .ZN(P1_U3287) );
  INV_X1 U8957 ( .A(n7080), .ZN(n7083) );
  OAI222_X1 U8958 ( .A1(n7747), .A2(n7082), .B1(n7750), .B2(n7083), .C1(n7081), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  OAI222_X1 U8959 ( .A1(P1_U3086), .A2(n7084), .B1(n9658), .B2(n7083), .C1(
        n7993), .C2(n5493), .ZN(P1_U3333) );
  AOI211_X1 U8960 ( .C1(n7087), .C2(n7086), .A(n5697), .B(n7085), .ZN(n7088)
         );
  INV_X1 U8961 ( .A(n7088), .ZN(n7092) );
  INV_X1 U8962 ( .A(n8888), .ZN(n8866) );
  NAND2_X1 U8963 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9239) );
  OAI21_X1 U8964 ( .B1(n7089), .B2(n8866), .A(n9239), .ZN(n7090) );
  AOI21_X1 U8965 ( .B1(n9927), .B2(n8887), .A(n7090), .ZN(n7091) );
  OAI211_X1 U8966 ( .C1(n8893), .C2(n7093), .A(n7092), .B(n7091), .ZN(P1_U3230) );
  INV_X1 U8967 ( .A(n7094), .ZN(n7095) );
  NAND2_X1 U8968 ( .A1(n7095), .A2(n6222), .ZN(n7096) );
  NAND2_X1 U8969 ( .A1(n7097), .A2(n7096), .ZN(n7134) );
  XNOR2_X1 U8970 ( .A(n7283), .B(n7974), .ZN(n7135) );
  XNOR2_X1 U8971 ( .A(n7135), .B(n8341), .ZN(n7133) );
  XOR2_X1 U8972 ( .A(n7134), .B(n7133), .Z(n7103) );
  NOR2_X1 U8973 ( .A1(n8323), .A2(n10063), .ZN(n7101) );
  NOR2_X1 U8974 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7098), .ZN(n7910) );
  AOI21_X1 U8975 ( .B1(n8297), .B2(n8342), .A(n7910), .ZN(n7099) );
  OAI21_X1 U8976 ( .B1(n7278), .B2(n8299), .A(n7099), .ZN(n7100) );
  AOI211_X1 U8977 ( .C1(n8291), .C2(n7279), .A(n7101), .B(n7100), .ZN(n7102)
         );
  OAI21_X1 U8978 ( .B1(n7103), .B2(n8328), .A(n7102), .ZN(P2_U3161) );
  XNOR2_X1 U8979 ( .A(n7104), .B(n7107), .ZN(n10034) );
  AND2_X1 U8980 ( .A1(n6804), .A2(n8445), .ZN(n7190) );
  NAND2_X1 U8981 ( .A1(n9716), .A2(n7190), .ZN(n8386) );
  INV_X1 U8982 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7116) );
  OAI21_X1 U8983 ( .B1(n7107), .B2(n7106), .A(n7105), .ZN(n7111) );
  OAI22_X1 U8984 ( .A1(n7109), .A2(n9712), .B1(n7108), .B2(n9710), .ZN(n7110)
         );
  AOI21_X1 U8985 ( .B1(n7111), .B2(n8510), .A(n7110), .ZN(n7112) );
  OAI21_X1 U8986 ( .B1(n10034), .B2(n7526), .A(n7112), .ZN(n10035) );
  INV_X1 U8987 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7113) );
  OAI22_X1 U8988 ( .A1(n9703), .A2(n7113), .B1(n8049), .B2(n9705), .ZN(n7114)
         );
  NOR2_X1 U8989 ( .A1(n10035), .A2(n7114), .ZN(n7115) );
  MUX2_X1 U8990 ( .A(n7116), .B(n7115), .S(n9716), .Z(n7117) );
  OAI21_X1 U8991 ( .B1(n10034), .B2(n8386), .A(n7117), .ZN(P2_U3231) );
  NAND2_X1 U8992 ( .A1(n7155), .A2(n7262), .ZN(n8193) );
  XNOR2_X1 U8993 ( .A(n7118), .B(n8193), .ZN(n10048) );
  INV_X1 U8994 ( .A(n10048), .ZN(n7129) );
  INV_X1 U8995 ( .A(n8193), .ZN(n7120) );
  XNOR2_X1 U8996 ( .A(n7119), .B(n7120), .ZN(n7123) );
  INV_X1 U8997 ( .A(n7526), .ZN(n7444) );
  NAND2_X1 U8998 ( .A1(n10048), .A2(n7444), .ZN(n7122) );
  AOI22_X1 U8999 ( .A1(n6453), .A2(n8513), .B1(n8512), .B2(n8344), .ZN(n7121)
         );
  OAI211_X1 U9000 ( .C1(n7123), .C2(n10024), .A(n7122), .B(n7121), .ZN(n10051)
         );
  MUX2_X1 U9001 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10051), .S(n9716), .Z(n7124)
         );
  INV_X1 U9002 ( .A(n7124), .ZN(n7128) );
  INV_X1 U9003 ( .A(n8523), .ZN(n8425) );
  INV_X1 U9004 ( .A(n9703), .ZN(n8521) );
  AOI22_X1 U9005 ( .A1(n8425), .A2(n7126), .B1(n8521), .B2(n7125), .ZN(n7127)
         );
  OAI211_X1 U9006 ( .C1(n7129), .C2(n8386), .A(n7128), .B(n7127), .ZN(P2_U3228) );
  INV_X1 U9007 ( .A(n7148), .ZN(n7132) );
  NAND2_X1 U9008 ( .A1(n7130), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8229) );
  NAND2_X1 U9009 ( .A1(n8775), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7131) );
  OAI211_X1 U9010 ( .C1(n7132), .C2(n8777), .A(n8229), .B(n7131), .ZN(P2_U3272) );
  INV_X1 U9011 ( .A(n7138), .ZN(n10069) );
  NAND2_X1 U9012 ( .A1(n7135), .A2(n7442), .ZN(n7136) );
  XNOR2_X1 U9013 ( .A(n7138), .B(n7974), .ZN(n7302) );
  XNOR2_X1 U9014 ( .A(n7302), .B(n7278), .ZN(n7140) );
  AOI21_X1 U9015 ( .B1(n7139), .B2(n7140), .A(n8328), .ZN(n7141) );
  NAND2_X1 U9016 ( .A1(n7141), .A2(n7305), .ZN(n7146) );
  INV_X1 U9017 ( .A(n8299), .ZN(n8320) );
  AOI21_X1 U9018 ( .B1(n8320), .B2(n8339), .A(n7142), .ZN(n7143) );
  OAI21_X1 U9019 ( .B1(n8322), .B2(n7442), .A(n7143), .ZN(n7144) );
  AOI21_X1 U9020 ( .B1(n8291), .B2(n7447), .A(n7144), .ZN(n7145) );
  OAI211_X1 U9021 ( .C1(n10069), .C2(n8323), .A(n7146), .B(n7145), .ZN(
        P2_U3171) );
  NAND2_X1 U9022 ( .A1(n7148), .A2(n7147), .ZN(n7149) );
  OAI211_X1 U9023 ( .C1(n7150), .C2(n7993), .A(n7149), .B(n9186), .ZN(P1_U3332) );
  INV_X1 U9024 ( .A(n8062), .ZN(n8072) );
  NOR2_X1 U9025 ( .A1(n8194), .A2(n8072), .ZN(n7153) );
  INV_X1 U9026 ( .A(n7272), .ZN(n7151) );
  AOI21_X1 U9027 ( .B1(n7153), .B2(n7152), .A(n7151), .ZN(n10061) );
  INV_X1 U9028 ( .A(n10061), .ZN(n7169) );
  OAI22_X1 U9029 ( .A1(n7442), .A2(n9712), .B1(n7154), .B2(n9710), .ZN(n7164)
         );
  NAND2_X1 U9030 ( .A1(n7119), .A2(n7155), .ZN(n7263) );
  NAND2_X1 U9031 ( .A1(n7263), .A2(n7156), .ZN(n7275) );
  OR2_X1 U9032 ( .A1(n8194), .A2(n4852), .ZN(n7157) );
  AND2_X1 U9033 ( .A1(n7275), .A2(n7157), .ZN(n7162) );
  NAND2_X1 U9034 ( .A1(n7263), .A2(n7158), .ZN(n7159) );
  AND2_X1 U9035 ( .A1(n7159), .A2(n4852), .ZN(n7160) );
  NAND2_X1 U9036 ( .A1(n7160), .A2(n8194), .ZN(n7161) );
  AOI21_X1 U9037 ( .B1(n7162), .B2(n7161), .A(n10024), .ZN(n7163) );
  AOI211_X1 U9038 ( .C1(n10061), .C2(n7444), .A(n7164), .B(n7163), .ZN(n10058)
         );
  MUX2_X1 U9039 ( .A(n7924), .B(n10058), .S(n9716), .Z(n7168) );
  AOI22_X1 U9040 ( .A1(n8425), .A2(n7166), .B1(n8521), .B2(n7165), .ZN(n7167)
         );
  OAI211_X1 U9041 ( .C1(n7169), .C2(n8386), .A(n7168), .B(n7167), .ZN(P2_U3226) );
  NAND2_X1 U9042 ( .A1(n7438), .A2(n8084), .ZN(n7171) );
  XNOR2_X1 U9043 ( .A(n7336), .B(n8339), .ZN(n8200) );
  INV_X1 U9044 ( .A(n8200), .ZN(n7170) );
  XNOR2_X1 U9045 ( .A(n7171), .B(n7170), .ZN(n7177) );
  INV_X1 U9046 ( .A(n7177), .ZN(n10077) );
  XNOR2_X1 U9047 ( .A(n7172), .B(n8200), .ZN(n7173) );
  NAND2_X1 U9048 ( .A1(n7173), .A2(n8510), .ZN(n7179) );
  NAND2_X1 U9049 ( .A1(n8340), .A2(n8512), .ZN(n7175) );
  NAND2_X1 U9050 ( .A1(n8338), .A2(n8513), .ZN(n7174) );
  NAND2_X1 U9051 ( .A1(n7175), .A2(n7174), .ZN(n7176) );
  AOI21_X1 U9052 ( .B1(n7177), .B2(n7444), .A(n7176), .ZN(n7178) );
  NAND2_X1 U9053 ( .A1(n7179), .A2(n7178), .ZN(n10079) );
  NAND2_X1 U9054 ( .A1(n10079), .A2(n9716), .ZN(n7183) );
  INV_X1 U9055 ( .A(n7341), .ZN(n7180) );
  OAI22_X1 U9056 ( .A1(n9716), .A2(n5885), .B1(n7180), .B2(n9703), .ZN(n7181)
         );
  AOI21_X1 U9057 ( .B1(n8425), .B2(n7336), .A(n7181), .ZN(n7182) );
  OAI211_X1 U9058 ( .C1(n10077), .C2(n8386), .A(n7183), .B(n7182), .ZN(
        P2_U3223) );
  AND2_X1 U9059 ( .A1(n8060), .A2(n8069), .ZN(n8189) );
  NAND2_X1 U9060 ( .A1(n7198), .A2(n7184), .ZN(n7186) );
  NAND2_X1 U9061 ( .A1(n7186), .A2(n7185), .ZN(n7187) );
  XOR2_X1 U9062 ( .A(n8189), .B(n7187), .Z(n7188) );
  AOI222_X1 U9063 ( .A1(n8510), .A2(n7188), .B1(n8343), .B2(n8513), .C1(n8345), 
        .C2(n8512), .ZN(n10043) );
  XNOR2_X1 U9064 ( .A(n7189), .B(n8189), .ZN(n10046) );
  INV_X1 U9065 ( .A(n7190), .ZN(n7191) );
  NAND2_X1 U9066 ( .A1(n7526), .A2(n7191), .ZN(n9714) );
  AOI22_X1 U9067 ( .A1(n8425), .A2(n7193), .B1(n8521), .B2(n7192), .ZN(n7194)
         );
  OAI21_X1 U9068 ( .B1(n7195), .B2(n9716), .A(n7194), .ZN(n7196) );
  AOI21_X1 U9069 ( .B1(n10046), .B2(n8525), .A(n7196), .ZN(n7197) );
  OAI21_X1 U9070 ( .B1(n10043), .B2(n9719), .A(n7197), .ZN(P2_U3229) );
  XOR2_X1 U9071 ( .A(n8190), .B(n7198), .Z(n7199) );
  AOI222_X1 U9072 ( .A1(n8510), .A2(n7199), .B1(n8344), .B2(n8513), .C1(n8346), 
        .C2(n8512), .ZN(n10039) );
  XNOR2_X1 U9073 ( .A(n7200), .B(n8190), .ZN(n10042) );
  AOI22_X1 U9074 ( .A1(n8425), .A2(n7202), .B1(n8521), .B2(n7201), .ZN(n7203)
         );
  OAI21_X1 U9075 ( .B1(n7204), .B2(n9716), .A(n7203), .ZN(n7205) );
  AOI21_X1 U9076 ( .B1(n10042), .B2(n8525), .A(n7205), .ZN(n7206) );
  OAI21_X1 U9077 ( .B1(n10039), .B2(n9719), .A(n7206), .ZN(P2_U3230) );
  XNOR2_X1 U9078 ( .A(n4349), .B(n7354), .ZN(n7208) );
  NOR2_X1 U9079 ( .A1(n7208), .A2(n5148), .ZN(n7353) );
  AOI21_X1 U9080 ( .B1(n5148), .B2(n7208), .A(n7353), .ZN(n7213) );
  OAI22_X1 U9081 ( .A1(n7209), .A2(n9469), .B1(n7230), .B2(n9467), .ZN(n9866)
         );
  AOI22_X1 U9082 ( .A1(n9866), .A2(n8888), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n7210) );
  OAI21_X1 U9083 ( .B1(n8893), .B2(n9868), .A(n7210), .ZN(n7211) );
  AOI21_X1 U9084 ( .B1(n9870), .B2(n8887), .A(n7211), .ZN(n7212) );
  OAI21_X1 U9085 ( .B1(n7213), .B2(n5697), .A(n7212), .ZN(P1_U3227) );
  NAND2_X1 U9086 ( .A1(n8043), .A2(n8036), .ZN(n7214) );
  NAND2_X1 U9087 ( .A1(n7215), .A2(n7214), .ZN(n10032) );
  INV_X1 U9088 ( .A(n10032), .ZN(n7226) );
  NAND2_X1 U9089 ( .A1(n10032), .A2(n7444), .ZN(n7221) );
  OAI21_X1 U9090 ( .B1(n7217), .B2(n8043), .A(n7216), .ZN(n7218) );
  NAND2_X1 U9091 ( .A1(n7218), .A2(n8510), .ZN(n7220) );
  AOI22_X1 U9092 ( .A1(n8513), .A2(n8346), .B1(n8349), .B2(n8512), .ZN(n7219)
         );
  NAND3_X1 U9093 ( .A1(n7221), .A2(n7220), .A3(n7219), .ZN(n10030) );
  MUX2_X1 U9094 ( .A(n10030), .B(P2_REG2_REG_1__SCAN_IN), .S(n9719), .Z(n7222)
         );
  INV_X1 U9095 ( .A(n7222), .ZN(n7225) );
  AOI22_X1 U9096 ( .A1(n8425), .A2(n7223), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8521), .ZN(n7224) );
  OAI211_X1 U9097 ( .C1(n7226), .C2(n8386), .A(n7225), .B(n7224), .ZN(P2_U3232) );
  XOR2_X1 U9098 ( .A(n7228), .B(n7227), .Z(n7234) );
  NAND2_X1 U9099 ( .A1(n9204), .A2(n9431), .ZN(n7229) );
  OAI21_X1 U9100 ( .B1(n7230), .B2(n9469), .A(n7229), .ZN(n9853) );
  AOI22_X1 U9101 ( .A1(n9853), .A2(n8888), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7231) );
  OAI21_X1 U9102 ( .B1(n8862), .B2(n9855), .A(n7231), .ZN(n7232) );
  AOI21_X1 U9103 ( .B1(n9857), .B2(n8887), .A(n7232), .ZN(n7233) );
  OAI21_X1 U9104 ( .B1(n7234), .B2(n5697), .A(n7233), .ZN(P1_U3213) );
  XOR2_X1 U9105 ( .A(n7235), .B(n7237), .Z(n9951) );
  INV_X1 U9106 ( .A(n9862), .ZN(n7248) );
  INV_X1 U9107 ( .A(n8969), .ZN(n8972) );
  AOI21_X1 U9108 ( .B1(n8973), .B2(n8971), .A(n8972), .ZN(n9848) );
  OAI21_X1 U9109 ( .B1(n9848), .B2(n9847), .A(n7236), .ZN(n7238) );
  AOI21_X1 U9110 ( .B1(n7238), .B2(n7237), .A(n9465), .ZN(n7240) );
  OR2_X1 U9111 ( .A1(n7238), .A2(n7237), .ZN(n7326) );
  NAND2_X1 U9112 ( .A1(n9205), .A2(n9433), .ZN(n7239) );
  OAI21_X1 U9113 ( .B1(n7287), .B2(n9467), .A(n7239), .ZN(n7456) );
  AOI21_X1 U9114 ( .B1(n7240), .B2(n7326), .A(n7456), .ZN(n7241) );
  OAI21_X1 U9115 ( .B1(n9951), .B2(n9851), .A(n7241), .ZN(n9954) );
  NAND2_X1 U9116 ( .A1(n9954), .A2(n9346), .ZN(n7247) );
  OAI22_X1 U9117 ( .A1(n9528), .A2(n7242), .B1(n7460), .B2(n9501), .ZN(n7245)
         );
  INV_X1 U9118 ( .A(n9859), .ZN(n7243) );
  OAI211_X1 U9119 ( .C1(n7243), .C2(n9953), .A(n9892), .B(n7322), .ZN(n9952)
         );
  NOR2_X1 U9120 ( .A1(n9952), .A2(n9351), .ZN(n7244) );
  AOI211_X1 U9121 ( .C1(n9884), .C2(n7457), .A(n7245), .B(n7244), .ZN(n7246)
         );
  OAI211_X1 U9122 ( .C1(n9951), .C2(n7248), .A(n7247), .B(n7246), .ZN(P1_U3285) );
  INV_X1 U9123 ( .A(n8525), .ZN(n7436) );
  OR2_X1 U9124 ( .A1(n7250), .A2(n8203), .ZN(n7251) );
  NAND2_X1 U9125 ( .A1(n7249), .A2(n7251), .ZN(n10089) );
  XNOR2_X1 U9126 ( .A(n7252), .B(n8203), .ZN(n7253) );
  NAND2_X1 U9127 ( .A1(n7253), .A2(n8510), .ZN(n7255) );
  AOI22_X1 U9128 ( .A1(n8512), .A2(n8338), .B1(n8336), .B2(n8513), .ZN(n7254)
         );
  NAND2_X1 U9129 ( .A1(n7255), .A2(n7254), .ZN(n10091) );
  NAND2_X1 U9130 ( .A1(n10091), .A2(n9716), .ZN(n7259) );
  INV_X1 U9131 ( .A(n7318), .ZN(n7256) );
  OAI22_X1 U9132 ( .A1(n9716), .A2(n4585), .B1(n7256), .B2(n9703), .ZN(n7257)
         );
  AOI21_X1 U9133 ( .B1(n7315), .B2(n8425), .A(n7257), .ZN(n7258) );
  OAI211_X1 U9134 ( .C1(n7436), .C2(n10089), .A(n7259), .B(n7258), .ZN(
        P2_U3221) );
  AND2_X1 U9135 ( .A1(n8063), .A2(n8062), .ZN(n8195) );
  NAND2_X1 U9136 ( .A1(n7260), .A2(n8059), .ZN(n7261) );
  XOR2_X1 U9137 ( .A(n8195), .B(n7261), .Z(n10055) );
  INV_X1 U9138 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7266) );
  NAND2_X1 U9139 ( .A1(n7263), .A2(n7262), .ZN(n7264) );
  XNOR2_X1 U9140 ( .A(n7264), .B(n8195), .ZN(n7265) );
  AOI222_X1 U9141 ( .A1(n8510), .A2(n7265), .B1(n8342), .B2(n8513), .C1(n8343), 
        .C2(n8512), .ZN(n10054) );
  MUX2_X1 U9142 ( .A(n7266), .B(n10054), .S(n9716), .Z(n7270) );
  AOI22_X1 U9143 ( .A1(n8425), .A2(n7268), .B1(n8521), .B2(n7267), .ZN(n7269)
         );
  OAI211_X1 U9144 ( .C1(n7436), .C2(n10055), .A(n7270), .B(n7269), .ZN(
        P2_U3227) );
  NAND2_X1 U9145 ( .A1(n8085), .A2(n8083), .ZN(n8198) );
  NAND2_X1 U9146 ( .A1(n7272), .A2(n7271), .ZN(n7273) );
  XOR2_X1 U9147 ( .A(n8198), .B(n7273), .Z(n10064) );
  NAND2_X1 U9148 ( .A1(n7275), .A2(n7274), .ZN(n7276) );
  XOR2_X1 U9149 ( .A(n8198), .B(n7276), .Z(n7277) );
  OAI222_X1 U9150 ( .A1(n9712), .A2(n7278), .B1(n9710), .B2(n6222), .C1(n10024), .C2(n7277), .ZN(n10066) );
  NAND2_X1 U9151 ( .A1(n10066), .A2(n9716), .ZN(n7285) );
  INV_X1 U9152 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7281) );
  INV_X1 U9153 ( .A(n7279), .ZN(n7280) );
  OAI22_X1 U9154 ( .A1(n9716), .A2(n7281), .B1(n7280), .B2(n9703), .ZN(n7282)
         );
  AOI21_X1 U9155 ( .B1(n8425), .B2(n7283), .A(n7282), .ZN(n7284) );
  OAI211_X1 U9156 ( .C1(n10064), .C2(n7436), .A(n7285), .B(n7284), .ZN(
        P2_U3225) );
  XNOR2_X1 U9157 ( .A(n7286), .B(n8931), .ZN(n7290) );
  OR2_X1 U9158 ( .A1(n9201), .A2(n9467), .ZN(n7289) );
  OR2_X1 U9159 ( .A1(n7287), .A2(n9469), .ZN(n7288) );
  NAND2_X1 U9160 ( .A1(n7289), .A2(n7288), .ZN(n7575) );
  AOI21_X1 U9161 ( .B1(n7290), .B2(n9882), .A(n7575), .ZN(n9966) );
  XNOR2_X1 U9162 ( .A(n7291), .B(n8931), .ZN(n9970) );
  NAND2_X1 U9163 ( .A1(n9970), .A2(n9897), .ZN(n7298) );
  OAI22_X1 U9164 ( .A1(n9528), .A2(n7292), .B1(n7578), .B2(n9501), .ZN(n7296)
         );
  INV_X1 U9165 ( .A(n7574), .ZN(n9968) );
  INV_X1 U9166 ( .A(n7324), .ZN(n7294) );
  INV_X1 U9167 ( .A(n7293), .ZN(n7538) );
  OAI211_X1 U9168 ( .C1(n9968), .C2(n7294), .A(n7538), .B(n9892), .ZN(n9965)
         );
  NOR2_X1 U9169 ( .A1(n9965), .A2(n9351), .ZN(n7295) );
  AOI211_X1 U9170 ( .C1(n9884), .C2(n7574), .A(n7296), .B(n7295), .ZN(n7297)
         );
  OAI211_X1 U9171 ( .C1(n9523), .C2(n9966), .A(n7298), .B(n7297), .ZN(P1_U3283) );
  INV_X1 U9172 ( .A(n7299), .ZN(n7371) );
  OAI222_X1 U9173 ( .A1(n7301), .A2(P1_U3086), .B1(n9658), .B2(n7371), .C1(
        n7300), .C2(n7993), .ZN(P1_U3331) );
  INV_X1 U9174 ( .A(n7302), .ZN(n7303) );
  NAND2_X1 U9175 ( .A1(n7303), .A2(n8340), .ZN(n7304) );
  XNOR2_X1 U9176 ( .A(n7390), .B(n7974), .ZN(n7386) );
  XNOR2_X1 U9177 ( .A(n7336), .B(n7974), .ZN(n7335) );
  AOI22_X1 U9178 ( .A1(n7386), .A2(n7385), .B1(n7441), .B2(n7335), .ZN(n7306)
         );
  NAND2_X1 U9179 ( .A1(n7382), .A2(n7306), .ZN(n7311) );
  INV_X1 U9180 ( .A(n7386), .ZN(n7309) );
  OAI21_X1 U9181 ( .B1(n7335), .B2(n7441), .A(n7385), .ZN(n7308) );
  INV_X1 U9182 ( .A(n7335), .ZN(n7383) );
  AND2_X1 U9183 ( .A1(n8339), .A2(n8338), .ZN(n7307) );
  AOI22_X1 U9184 ( .A1(n7309), .A2(n7308), .B1(n7383), .B2(n7307), .ZN(n7310)
         );
  XNOR2_X1 U9185 ( .A(n7315), .B(n7961), .ZN(n7372) );
  XNOR2_X1 U9186 ( .A(n7372), .B(n9709), .ZN(n7312) );
  XNOR2_X1 U9187 ( .A(n7373), .B(n7312), .ZN(n7320) );
  INV_X1 U9188 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7313) );
  NOR2_X1 U9189 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7313), .ZN(n7849) );
  AOI21_X1 U9190 ( .B1(n8297), .B2(n8338), .A(n7849), .ZN(n7314) );
  OAI21_X1 U9191 ( .B1(n8112), .B2(n8299), .A(n7314), .ZN(n7317) );
  NAND2_X1 U9192 ( .A1(n7315), .A2(n10028), .ZN(n10087) );
  NOR2_X1 U9193 ( .A1(n10087), .A2(n8313), .ZN(n7316) );
  AOI211_X1 U9194 ( .C1(n7318), .C2(n8291), .A(n7317), .B(n7316), .ZN(n7319)
         );
  OAI21_X1 U9195 ( .B1(n7320), .B2(n8328), .A(n7319), .ZN(P2_U3164) );
  XOR2_X1 U9196 ( .A(n7327), .B(n7321), .Z(n9958) );
  AOI21_X1 U9197 ( .B1(n7322), .B2(n9959), .A(n9909), .ZN(n7325) );
  NOR2_X1 U9198 ( .A1(n7540), .A2(n9467), .ZN(n7323) );
  AOI21_X1 U9199 ( .B1(n7325), .B2(n7324), .A(n7323), .ZN(n9960) );
  NAND2_X1 U9200 ( .A1(n7326), .A2(n8977), .ZN(n7328) );
  XNOR2_X1 U9201 ( .A(n7328), .B(n7327), .ZN(n7329) );
  AOI22_X1 U9202 ( .A1(n7329), .A2(n9882), .B1(n9433), .B2(n9204), .ZN(n9961)
         );
  OAI21_X1 U9203 ( .B1(n9308), .B2(n9960), .A(n9961), .ZN(n7330) );
  NAND2_X1 U9204 ( .A1(n7330), .A2(n9346), .ZN(n7334) );
  OAI22_X1 U9205 ( .A1(n9528), .A2(n7331), .B1(n7557), .B2(n9501), .ZN(n7332)
         );
  AOI21_X1 U9206 ( .B1(n9884), .B2(n9959), .A(n7332), .ZN(n7333) );
  OAI211_X1 U9207 ( .C1(n9958), .C2(n9530), .A(n7334), .B(n7333), .ZN(P1_U3284) );
  XNOR2_X1 U9208 ( .A(n7382), .B(n8339), .ZN(n7384) );
  XNOR2_X1 U9209 ( .A(n7384), .B(n7335), .ZN(n7343) );
  NAND2_X1 U9210 ( .A1(n7336), .A2(n10028), .ZN(n10075) );
  NOR2_X1 U9211 ( .A1(n10075), .A2(n8313), .ZN(n7340) );
  INV_X1 U9212 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7337) );
  NOR2_X1 U9213 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7337), .ZN(n7886) );
  AOI21_X1 U9214 ( .B1(n8297), .B2(n8340), .A(n7886), .ZN(n7338) );
  OAI21_X1 U9215 ( .B1(n7385), .B2(n8299), .A(n7338), .ZN(n7339) );
  AOI211_X1 U9216 ( .C1(n8291), .C2(n7341), .A(n7340), .B(n7339), .ZN(n7342)
         );
  OAI21_X1 U9217 ( .B1(n7343), .B2(n8328), .A(n7342), .ZN(P2_U3157) );
  AND2_X1 U9218 ( .A1(n8101), .A2(n8099), .ZN(n8202) );
  XNOR2_X1 U9219 ( .A(n7344), .B(n8202), .ZN(n7345) );
  OAI222_X1 U9220 ( .A1(n9712), .A2(n9709), .B1(n9710), .B2(n7441), .C1(n10024), .C2(n7345), .ZN(n10082) );
  INV_X1 U9221 ( .A(n10082), .ZN(n7352) );
  NAND2_X1 U9222 ( .A1(n7346), .A2(n8090), .ZN(n7347) );
  XNOR2_X1 U9223 ( .A(n7347), .B(n8202), .ZN(n10085) );
  INV_X1 U9224 ( .A(n7390), .ZN(n7349) );
  AOI22_X1 U9225 ( .A1(n9719), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n8521), .B2(
        n7393), .ZN(n7348) );
  OAI21_X1 U9226 ( .B1(n7349), .B2(n8523), .A(n7348), .ZN(n7350) );
  AOI21_X1 U9227 ( .B1(n10085), .B2(n8525), .A(n7350), .ZN(n7351) );
  OAI21_X1 U9228 ( .B1(n7352), .B2(n9719), .A(n7351), .ZN(P2_U3222) );
  AOI21_X1 U9229 ( .B1(n7354), .B2(n4349), .A(n7353), .ZN(n7358) );
  XOR2_X1 U9230 ( .A(n7356), .B(n7355), .Z(n7357) );
  XNOR2_X1 U9231 ( .A(n7358), .B(n7357), .ZN(n7365) );
  AOI22_X1 U9232 ( .A1(n7359), .A2(n8888), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7360) );
  OAI21_X1 U9233 ( .B1(n8893), .B2(n7361), .A(n7360), .ZN(n7362) );
  AOI21_X1 U9234 ( .B1(n7363), .B2(n8887), .A(n7362), .ZN(n7364) );
  OAI21_X1 U9235 ( .B1(n7365), .B2(n5697), .A(n7364), .ZN(P1_U3239) );
  INV_X1 U9236 ( .A(n7366), .ZN(n7749) );
  OAI222_X1 U9237 ( .A1(P1_U3086), .A2(n7368), .B1(n9658), .B2(n7749), .C1(
        n7367), .C2(n7993), .ZN(P1_U3330) );
  OAI222_X1 U9238 ( .A1(n8777), .A2(n7371), .B1(P2_U3151), .B2(n7370), .C1(
        n7369), .C2(n7747), .ZN(P2_U3271) );
  OAI21_X1 U9239 ( .B1(n7373), .B2(n8337), .A(n7372), .ZN(n7375) );
  NAND2_X1 U9240 ( .A1(n7373), .A2(n8337), .ZN(n7374) );
  NAND2_X1 U9241 ( .A1(n7375), .A2(n7374), .ZN(n7497) );
  XNOR2_X1 U9242 ( .A(n8113), .B(n7961), .ZN(n7493) );
  XNOR2_X1 U9243 ( .A(n7493), .B(n8112), .ZN(n7376) );
  XNOR2_X1 U9244 ( .A(n7497), .B(n7376), .ZN(n7381) );
  AND2_X1 U9245 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n7830) );
  AOI21_X1 U9246 ( .B1(n8320), .B2(n8335), .A(n7830), .ZN(n7377) );
  OAI21_X1 U9247 ( .B1(n8322), .B2(n9709), .A(n7377), .ZN(n7379) );
  INV_X1 U9248 ( .A(n8113), .ZN(n9720) );
  NOR2_X1 U9249 ( .A1(n9720), .A2(n8323), .ZN(n7378) );
  AOI211_X1 U9250 ( .C1(n9702), .C2(n8291), .A(n7379), .B(n7378), .ZN(n7380)
         );
  OAI21_X1 U9251 ( .B1(n7381), .B2(n8328), .A(n7380), .ZN(P2_U3174) );
  OAI22_X1 U9252 ( .A1(n7384), .A2(n7383), .B1(n8339), .B2(n7382), .ZN(n7388)
         );
  XNOR2_X1 U9253 ( .A(n7386), .B(n7385), .ZN(n7387) );
  XNOR2_X1 U9254 ( .A(n7388), .B(n7387), .ZN(n7395) );
  AND2_X1 U9255 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7872) );
  AOI21_X1 U9256 ( .B1(n8297), .B2(n8339), .A(n7872), .ZN(n7389) );
  OAI21_X1 U9257 ( .B1(n9709), .B2(n8299), .A(n7389), .ZN(n7392) );
  NAND2_X1 U9258 ( .A1(n7390), .A2(n10028), .ZN(n10081) );
  NOR2_X1 U9259 ( .A1(n10081), .A2(n8313), .ZN(n7391) );
  AOI211_X1 U9260 ( .C1(n7393), .C2(n8291), .A(n7392), .B(n7391), .ZN(n7394)
         );
  OAI21_X1 U9261 ( .B1(n7395), .B2(n8328), .A(n7394), .ZN(P2_U3176) );
  INV_X1 U9262 ( .A(n7396), .ZN(n8934) );
  XNOR2_X1 U9263 ( .A(n7397), .B(n8934), .ZN(n7466) );
  INV_X1 U9264 ( .A(n7466), .ZN(n7409) );
  INV_X1 U9265 ( .A(n7417), .ZN(n7399) );
  AOI211_X1 U9266 ( .C1(n7523), .C2(n7398), .A(n9909), .B(n7399), .ZN(n7465)
         );
  INV_X1 U9267 ( .A(n7523), .ZN(n7400) );
  NOR2_X1 U9268 ( .A1(n7400), .A2(n9526), .ZN(n7403) );
  OAI22_X1 U9269 ( .A1(n9528), .A2(n7401), .B1(n7518), .B2(n9501), .ZN(n7402)
         );
  AOI211_X1 U9270 ( .C1(n7465), .C2(n9896), .A(n7403), .B(n7402), .ZN(n7408)
         );
  NAND2_X1 U9271 ( .A1(n7404), .A2(n8995), .ZN(n7405) );
  XNOR2_X1 U9272 ( .A(n7405), .B(n8934), .ZN(n7406) );
  OAI222_X1 U9273 ( .A1(n9469), .A2(n9201), .B1(n9467), .B2(n9004), .C1(n9465), 
        .C2(n7406), .ZN(n7464) );
  NAND2_X1 U9274 ( .A1(n7464), .A2(n9346), .ZN(n7407) );
  OAI211_X1 U9275 ( .C1(n7409), .C2(n9530), .A(n7408), .B(n7407), .ZN(P1_U3281) );
  XNOR2_X1 U9276 ( .A(n7410), .B(n8935), .ZN(n7411) );
  NAND2_X1 U9277 ( .A1(n7411), .A2(n9882), .ZN(n7415) );
  OR2_X1 U9278 ( .A1(n7539), .A2(n9469), .ZN(n7413) );
  NAND2_X1 U9279 ( .A1(n9198), .A2(n9431), .ZN(n7412) );
  NAND2_X1 U9280 ( .A1(n7413), .A2(n7412), .ZN(n7604) );
  INV_X1 U9281 ( .A(n7604), .ZN(n7414) );
  NAND2_X1 U9282 ( .A1(n7415), .A2(n7414), .ZN(n7477) );
  INV_X1 U9283 ( .A(n7477), .ZN(n7424) );
  XNOR2_X1 U9284 ( .A(n7416), .B(n8935), .ZN(n7479) );
  NAND2_X1 U9285 ( .A1(n7479), .A2(n9897), .ZN(n7423) );
  AOI211_X1 U9286 ( .C1(n9005), .C2(n7417), .A(n9909), .B(n7648), .ZN(n7478)
         );
  INV_X1 U9287 ( .A(n9005), .ZN(n7418) );
  NOR2_X1 U9288 ( .A1(n7418), .A2(n9526), .ZN(n7421) );
  OAI22_X1 U9289 ( .A1(n9528), .A2(n7419), .B1(n7606), .B2(n9501), .ZN(n7420)
         );
  AOI211_X1 U9290 ( .C1(n7478), .C2(n9896), .A(n7421), .B(n7420), .ZN(n7422)
         );
  OAI211_X1 U9291 ( .C1(n9900), .C2(n7424), .A(n7423), .B(n7422), .ZN(P1_U3280) );
  OR2_X1 U9292 ( .A1(n7425), .A2(n8121), .ZN(n7426) );
  NAND2_X1 U9293 ( .A1(n7427), .A2(n7426), .ZN(n7564) );
  OAI211_X1 U9294 ( .C1(n7428), .C2(n8207), .A(n7506), .B(n8510), .ZN(n7431)
         );
  OAI22_X1 U9295 ( .A1(n9711), .A2(n9710), .B1(n7731), .B2(n9712), .ZN(n7429)
         );
  INV_X1 U9296 ( .A(n7429), .ZN(n7430) );
  NAND2_X1 U9297 ( .A1(n7431), .A2(n7430), .ZN(n7566) );
  NAND2_X1 U9298 ( .A1(n7566), .A2(n9716), .ZN(n7435) );
  INV_X1 U9299 ( .A(n7596), .ZN(n7432) );
  OAI22_X1 U9300 ( .A1(n9716), .A2(n8363), .B1(n7432), .B2(n9703), .ZN(n7433)
         );
  AOI21_X1 U9301 ( .B1(n7589), .B2(n8425), .A(n7433), .ZN(n7434) );
  OAI211_X1 U9302 ( .C1(n7564), .C2(n7436), .A(n7435), .B(n7434), .ZN(P2_U3218) );
  XOR2_X1 U9303 ( .A(n7437), .B(n8197), .Z(n7446) );
  INV_X1 U9304 ( .A(n7438), .ZN(n7439) );
  AOI21_X1 U9305 ( .B1(n8197), .B2(n7440), .A(n7439), .ZN(n10073) );
  OAI22_X1 U9306 ( .A1(n7442), .A2(n9710), .B1(n7441), .B2(n9712), .ZN(n7443)
         );
  AOI21_X1 U9307 ( .B1(n10073), .B2(n7444), .A(n7443), .ZN(n7445) );
  OAI21_X1 U9308 ( .B1(n10024), .B2(n7446), .A(n7445), .ZN(n10070) );
  INV_X1 U9309 ( .A(n10070), .ZN(n7452) );
  INV_X1 U9310 ( .A(n8386), .ZN(n7450) );
  AOI22_X1 U9311 ( .A1(n9719), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n8521), .B2(
        n7447), .ZN(n7448) );
  OAI21_X1 U9312 ( .B1(n10069), .B2(n8523), .A(n7448), .ZN(n7449) );
  AOI21_X1 U9313 ( .B1(n10073), .B2(n7450), .A(n7449), .ZN(n7451) );
  OAI21_X1 U9314 ( .B1(n7452), .B2(n9719), .A(n7451), .ZN(P2_U3224) );
  XOR2_X1 U9315 ( .A(n7552), .B(n7551), .Z(n7455) );
  INV_X1 U9316 ( .A(n7453), .ZN(n7454) );
  NAND2_X1 U9317 ( .A1(n7455), .A2(n7454), .ZN(n7550) );
  OAI21_X1 U9318 ( .B1(n7455), .B2(n7454), .A(n7550), .ZN(n7462) );
  AOI22_X1 U9319 ( .A1(n7456), .A2(n8888), .B1(P1_REG3_REG_8__SCAN_IN), .B2(
        P1_U3086), .ZN(n7459) );
  NAND2_X1 U9320 ( .A1(n8887), .A2(n7457), .ZN(n7458) );
  OAI211_X1 U9321 ( .C1(n8893), .C2(n7460), .A(n7459), .B(n7458), .ZN(n7461)
         );
  AOI21_X1 U9322 ( .B1(n7462), .B2(n8895), .A(n7461), .ZN(n7463) );
  INV_X1 U9323 ( .A(n7463), .ZN(P1_U3221) );
  AOI211_X1 U9324 ( .C1(n7466), .C2(n9971), .A(n7465), .B(n7464), .ZN(n7470)
         );
  AOI22_X1 U9325 ( .A1(n7523), .A2(n6004), .B1(n9996), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7467) );
  OAI21_X1 U9326 ( .B1(n7470), .B2(n9996), .A(n7467), .ZN(P1_U3534) );
  INV_X1 U9327 ( .A(n9645), .ZN(n7481) );
  NOR2_X1 U9328 ( .A1(n9983), .A2(n5278), .ZN(n7468) );
  AOI21_X1 U9329 ( .B1(n7523), .B2(n7481), .A(n7468), .ZN(n7469) );
  OAI21_X1 U9330 ( .B1(n7470), .B2(n9982), .A(n7469), .ZN(P1_U3489) );
  INV_X1 U9331 ( .A(n7471), .ZN(n7475) );
  OAI222_X1 U9332 ( .A1(P1_U3086), .A2(n7473), .B1(n9658), .B2(n7475), .C1(
        n7472), .C2(n7993), .ZN(P1_U3329) );
  OAI222_X1 U9333 ( .A1(n7747), .A2(n7476), .B1(n7750), .B2(n7475), .C1(n7474), 
        .C2(P2_U3151), .ZN(P2_U3269) );
  AOI211_X1 U9334 ( .C1(n7479), .C2(n9971), .A(n7478), .B(n7477), .ZN(n7484)
         );
  NOR2_X1 U9335 ( .A1(n9983), .A2(n5300), .ZN(n7480) );
  AOI21_X1 U9336 ( .B1(n9005), .B2(n7481), .A(n7480), .ZN(n7482) );
  OAI21_X1 U9337 ( .B1(n7484), .B2(n9982), .A(n7482), .ZN(P1_U3492) );
  AOI22_X1 U9338 ( .A1(n9005), .A2(n6004), .B1(n9996), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n7483) );
  OAI21_X1 U9339 ( .B1(n7484), .B2(n9996), .A(n7483), .ZN(P1_U3535) );
  INV_X1 U9340 ( .A(n7498), .ZN(n7534) );
  NOR2_X1 U9341 ( .A1(n7534), .A2(n9705), .ZN(n7489) );
  INV_X1 U9342 ( .A(n7485), .ZN(n7486) );
  AOI21_X1 U9343 ( .B1(n8205), .B2(n7487), .A(n7486), .ZN(n7488) );
  OAI222_X1 U9344 ( .A1(n9712), .A2(n7693), .B1(n9710), .B2(n8112), .C1(n10024), .C2(n7488), .ZN(n7527) );
  AOI211_X1 U9345 ( .C1(n8521), .C2(n7502), .A(n7489), .B(n7527), .ZN(n7492)
         );
  XOR2_X1 U9346 ( .A(n7490), .B(n8205), .Z(n7528) );
  AOI22_X1 U9347 ( .A1(n7528), .A2(n8525), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9719), .ZN(n7491) );
  OAI21_X1 U9348 ( .B1(n7492), .B2(n9719), .A(n7491), .ZN(P2_U3219) );
  AND2_X1 U9349 ( .A1(n7493), .A2(n8336), .ZN(n7496) );
  INV_X1 U9350 ( .A(n7493), .ZN(n7494) );
  NAND2_X1 U9351 ( .A1(n7494), .A2(n8112), .ZN(n7495) );
  XNOR2_X1 U9352 ( .A(n7498), .B(n7974), .ZN(n7587) );
  XNOR2_X1 U9353 ( .A(n7587), .B(n8335), .ZN(n7585) );
  XOR2_X1 U9354 ( .A(n7586), .B(n7585), .Z(n7504) );
  NAND2_X1 U9355 ( .A1(n8297), .A2(n8336), .ZN(n7499) );
  NAND2_X1 U9356 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7817) );
  OAI211_X1 U9357 ( .C1(n7693), .C2(n8299), .A(n7499), .B(n7817), .ZN(n7501)
         );
  NOR2_X1 U9358 ( .A1(n7534), .A2(n8323), .ZN(n7500) );
  AOI211_X1 U9359 ( .C1(n7502), .C2(n8291), .A(n7501), .B(n7500), .ZN(n7503)
         );
  OAI21_X1 U9360 ( .B1(n7504), .B2(n8328), .A(n7503), .ZN(P2_U3155) );
  NAND2_X1 U9361 ( .A1(n7506), .A2(n7505), .ZN(n7507) );
  XNOR2_X1 U9362 ( .A(n7507), .B(n8208), .ZN(n7508) );
  OAI222_X1 U9363 ( .A1(n9712), .A2(n8311), .B1(n9710), .B2(n7693), .C1(n7508), 
        .C2(n10024), .ZN(n7669) );
  INV_X1 U9364 ( .A(n7669), .ZN(n7515) );
  OAI21_X1 U9365 ( .B1(n7510), .B2(n8126), .A(n7509), .ZN(n7511) );
  INV_X1 U9366 ( .A(n7511), .ZN(n7670) );
  INV_X1 U9367 ( .A(n7688), .ZN(n7698) );
  AOI22_X1 U9368 ( .A1(n9719), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8521), .B2(
        n7695), .ZN(n7512) );
  OAI21_X1 U9369 ( .B1(n7698), .B2(n8523), .A(n7512), .ZN(n7513) );
  AOI21_X1 U9370 ( .B1(n7670), .B2(n8525), .A(n7513), .ZN(n7514) );
  OAI21_X1 U9371 ( .B1(n7515), .B2(n9719), .A(n7514), .ZN(P2_U3217) );
  XOR2_X1 U9372 ( .A(n7517), .B(n7516), .Z(n7525) );
  INV_X1 U9373 ( .A(n7518), .ZN(n7519) );
  AOI22_X1 U9374 ( .A1(n8813), .A2(n9199), .B1(n8880), .B2(n7519), .ZN(n7521)
         );
  OAI211_X1 U9375 ( .C1(n9201), .C2(n8876), .A(n7521), .B(n7520), .ZN(n7522)
         );
  AOI21_X1 U9376 ( .B1(n7523), .B2(n8887), .A(n7522), .ZN(n7524) );
  OAI21_X1 U9377 ( .B1(n7525), .B2(n5697), .A(n7524), .ZN(P1_U3224) );
  INV_X1 U9378 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7529) );
  INV_X1 U9379 ( .A(n10072), .ZN(n10076) );
  NAND2_X1 U9380 ( .A1(n7526), .A2(n10076), .ZN(n10084) );
  AOI21_X1 U9381 ( .B1(n10084), .B2(n7528), .A(n7527), .ZN(n7531) );
  MUX2_X1 U9382 ( .A(n7529), .B(n7531), .S(n10094), .Z(n7530) );
  OAI21_X1 U9383 ( .B1(n7534), .B2(n8768), .A(n7530), .ZN(P2_U3432) );
  INV_X1 U9384 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7532) );
  MUX2_X1 U9385 ( .A(n7532), .B(n7531), .S(n10121), .Z(n7533) );
  OAI21_X1 U9386 ( .B1(n7534), .B2(n8576), .A(n7533), .ZN(P2_U3473) );
  INV_X1 U9387 ( .A(n9977), .ZN(n9957) );
  OAI21_X1 U9388 ( .B1(n7536), .B2(n8921), .A(n7535), .ZN(n9843) );
  INV_X1 U9389 ( .A(n7398), .ZN(n7537) );
  AOI211_X1 U9390 ( .C1(n9841), .C2(n7538), .A(n9909), .B(n7537), .ZN(n9842)
         );
  OAI22_X1 U9391 ( .A1(n7540), .A2(n9469), .B1(n7539), .B2(n9467), .ZN(n7628)
         );
  INV_X1 U9392 ( .A(n7404), .ZN(n7541) );
  AOI211_X1 U9393 ( .C1(n8921), .C2(n7542), .A(n9465), .B(n7541), .ZN(n7543)
         );
  AOI211_X1 U9394 ( .C1(n9981), .C2(n9843), .A(n7628), .B(n7543), .ZN(n9846)
         );
  INV_X1 U9395 ( .A(n9846), .ZN(n7544) );
  AOI211_X1 U9396 ( .C1(n9957), .C2(n9843), .A(n9842), .B(n7544), .ZN(n7549)
         );
  AOI22_X1 U9397 ( .A1(n9841), .A2(n6004), .B1(n9996), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7545) );
  OAI21_X1 U9398 ( .B1(n7549), .B2(n9996), .A(n7545), .ZN(P1_U3533) );
  OAI22_X1 U9399 ( .A1(n7546), .A2(n9645), .B1(n9983), .B2(n5238), .ZN(n7547)
         );
  INV_X1 U9400 ( .A(n7547), .ZN(n7548) );
  OAI21_X1 U9401 ( .B1(n7549), .B2(n9982), .A(n7548), .ZN(P1_U3486) );
  OAI21_X1 U9402 ( .B1(n7552), .B2(n7551), .A(n7550), .ZN(n7556) );
  XNOR2_X1 U9403 ( .A(n7554), .B(n7553), .ZN(n7555) );
  XNOR2_X1 U9404 ( .A(n7556), .B(n7555), .ZN(n7563) );
  OAI22_X1 U9405 ( .A1(n8876), .A2(n7558), .B1(n8893), .B2(n7557), .ZN(n7559)
         );
  AOI211_X1 U9406 ( .C1(n8813), .C2(n9202), .A(n7560), .B(n7559), .ZN(n7562)
         );
  NAND2_X1 U9407 ( .A1(n8887), .A2(n9959), .ZN(n7561) );
  OAI211_X1 U9408 ( .C1(n7563), .C2(n5697), .A(n7562), .B(n7561), .ZN(P1_U3231) );
  INV_X1 U9409 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7567) );
  INV_X1 U9410 ( .A(n10084), .ZN(n10088) );
  INV_X1 U9411 ( .A(n7589), .ZN(n7599) );
  OAI22_X1 U9412 ( .A1(n7564), .A2(n10088), .B1(n7599), .B2(n10068), .ZN(n7565) );
  NOR2_X1 U9413 ( .A1(n7566), .A2(n7565), .ZN(n7569) );
  MUX2_X1 U9414 ( .A(n7567), .B(n7569), .S(n10094), .Z(n7568) );
  INV_X1 U9415 ( .A(n7568), .ZN(P2_U3435) );
  MUX2_X1 U9416 ( .A(n8351), .B(n7569), .S(n10121), .Z(n7570) );
  INV_X1 U9417 ( .A(n7570), .ZN(P2_U3474) );
  XNOR2_X1 U9418 ( .A(n7622), .B(n7571), .ZN(n7572) );
  NAND2_X1 U9419 ( .A1(n7572), .A2(n7573), .ZN(n7621) );
  OAI21_X1 U9420 ( .B1(n7573), .B2(n7572), .A(n7621), .ZN(n7580) );
  NAND2_X1 U9421 ( .A1(n7574), .A2(n8887), .ZN(n7577) );
  AOI22_X1 U9422 ( .A1(n7575), .A2(n8888), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n7576) );
  OAI211_X1 U9423 ( .C1(n8893), .C2(n7578), .A(n7577), .B(n7576), .ZN(n7579)
         );
  AOI21_X1 U9424 ( .B1(n7580), .B2(n8895), .A(n7579), .ZN(n7581) );
  INV_X1 U9425 ( .A(n7581), .ZN(P1_U3217) );
  INV_X1 U9426 ( .A(n7582), .ZN(n7656) );
  OAI222_X1 U9427 ( .A1(n7747), .A2(n7584), .B1(n7750), .B2(n7656), .C1(
        P2_U3151), .C2(n7583), .ZN(P2_U3268) );
  NAND2_X1 U9428 ( .A1(n7587), .A2(n9711), .ZN(n7588) );
  XNOR2_X1 U9429 ( .A(n7589), .B(n7974), .ZN(n7684) );
  XNOR2_X1 U9430 ( .A(n7684), .B(n7693), .ZN(n7591) );
  AOI21_X1 U9431 ( .B1(n7590), .B2(n7591), .A(n8328), .ZN(n7593) );
  NAND2_X1 U9432 ( .A1(n7593), .A2(n7687), .ZN(n7598) );
  AND2_X1 U9433 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8353) );
  AOI21_X1 U9434 ( .B1(n8297), .B2(n8335), .A(n8353), .ZN(n7594) );
  OAI21_X1 U9435 ( .B1(n7731), .B2(n8299), .A(n7594), .ZN(n7595) );
  AOI21_X1 U9436 ( .B1(n8291), .B2(n7596), .A(n7595), .ZN(n7597) );
  OAI211_X1 U9437 ( .C1(n7599), .C2(n8323), .A(n7598), .B(n7597), .ZN(P2_U3181) );
  INV_X1 U9438 ( .A(n7600), .ZN(n7619) );
  OAI222_X1 U9439 ( .A1(n8777), .A2(n7619), .B1(n8223), .B2(P2_U3151), .C1(
        n7601), .C2(n7747), .ZN(P2_U3267) );
  XOR2_X1 U9440 ( .A(n7603), .B(n7602), .Z(n7609) );
  AOI22_X1 U9441 ( .A1(n7604), .A2(n8888), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n7605) );
  OAI21_X1 U9442 ( .B1(n8893), .B2(n7606), .A(n7605), .ZN(n7607) );
  AOI21_X1 U9443 ( .B1(n9005), .B2(n8887), .A(n7607), .ZN(n7608) );
  OAI21_X1 U9444 ( .B1(n7609), .B2(n5697), .A(n7608), .ZN(P1_U3234) );
  XNOR2_X1 U9445 ( .A(n7611), .B(n6459), .ZN(n7612) );
  AOI222_X1 U9446 ( .A1(n8510), .A2(n7612), .B1(n8511), .B2(n8513), .C1(n8333), 
        .C2(n8512), .ZN(n8585) );
  OAI21_X1 U9447 ( .B1(n7614), .B2(n6459), .A(n7613), .ZN(n8583) );
  INV_X1 U9448 ( .A(n8582), .ZN(n7732) );
  AOI22_X1 U9449 ( .A1(n9719), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8521), .B2(
        n7735), .ZN(n7615) );
  OAI21_X1 U9450 ( .B1(n7732), .B2(n8523), .A(n7615), .ZN(n7616) );
  AOI21_X1 U9451 ( .B1(n8583), .B2(n8525), .A(n7616), .ZN(n7617) );
  OAI21_X1 U9452 ( .B1(n8585), .B2(n9719), .A(n7617), .ZN(P2_U3216) );
  OAI222_X1 U9453 ( .A1(n7620), .A2(P1_U3086), .B1(n9658), .B2(n7619), .C1(
        n7618), .C2(n7993), .ZN(P1_U3327) );
  OAI21_X1 U9454 ( .B1(n7623), .B2(n7622), .A(n7621), .ZN(n7627) );
  XNOR2_X1 U9455 ( .A(n7625), .B(n7624), .ZN(n7626) );
  XNOR2_X1 U9456 ( .A(n7627), .B(n7626), .ZN(n7632) );
  AOI22_X1 U9457 ( .A1(n7628), .A2(n8888), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n7629) );
  OAI21_X1 U9458 ( .B1(n8862), .B2(n9839), .A(n7629), .ZN(n7630) );
  AOI21_X1 U9459 ( .B1(n9841), .B2(n8887), .A(n7630), .ZN(n7631) );
  OAI21_X1 U9460 ( .B1(n7632), .B2(n5697), .A(n7631), .ZN(P1_U3236) );
  XNOR2_X1 U9461 ( .A(n7634), .B(n7633), .ZN(n7635) );
  XNOR2_X1 U9462 ( .A(n7636), .B(n7635), .ZN(n7642) );
  NAND2_X1 U9463 ( .A1(n9197), .A2(n9431), .ZN(n7638) );
  NAND2_X1 U9464 ( .A1(n9199), .A2(n9433), .ZN(n7637) );
  NAND2_X1 U9465 ( .A1(n7638), .A2(n7637), .ZN(n7644) );
  AOI22_X1 U9466 ( .A1(n7644), .A2(n8888), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n7639) );
  OAI21_X1 U9467 ( .B1(n8893), .B2(n7651), .A(n7639), .ZN(n7640) );
  AOI21_X1 U9468 ( .B1(n9973), .B2(n8887), .A(n7640), .ZN(n7641) );
  OAI21_X1 U9469 ( .B1(n7642), .B2(n5697), .A(n7641), .ZN(P1_U3215) );
  AOI21_X1 U9470 ( .B1(n7643), .B2(n8938), .A(n9465), .ZN(n7646) );
  AOI21_X1 U9471 ( .B1(n7646), .B2(n7645), .A(n7644), .ZN(n9976) );
  XOR2_X1 U9472 ( .A(n7647), .B(n8938), .Z(n9978) );
  INV_X1 U9473 ( .A(n9978), .ZN(n9980) );
  NAND2_X1 U9474 ( .A1(n9980), .A2(n9897), .ZN(n7655) );
  INV_X1 U9475 ( .A(n7648), .ZN(n7649) );
  AOI211_X1 U9476 ( .C1(n9973), .C2(n7649), .A(n9909), .B(n7659), .ZN(n9972)
         );
  NOR2_X1 U9477 ( .A1(n7650), .A2(n9526), .ZN(n7653) );
  OAI22_X1 U9478 ( .A1(n9528), .A2(n9260), .B1(n7651), .B2(n9501), .ZN(n7652)
         );
  AOI211_X1 U9479 ( .C1(n9972), .C2(n9896), .A(n7653), .B(n7652), .ZN(n7654)
         );
  OAI211_X1 U9480 ( .C1(n9900), .C2(n9976), .A(n7655), .B(n7654), .ZN(P1_U3279) );
  OAI222_X1 U9481 ( .A1(P1_U3086), .A2(n9728), .B1(n9658), .B2(n7656), .C1(
        n8684), .C2(n7993), .ZN(P1_U3328) );
  INV_X1 U9482 ( .A(n7662), .ZN(n8941) );
  XNOR2_X1 U9483 ( .A(n7657), .B(n8941), .ZN(n7716) );
  OAI22_X1 U9484 ( .A1(n9528), .A2(n7658), .B1(n8892), .B2(n9501), .ZN(n7661)
         );
  OAI211_X1 U9485 ( .C1(n7659), .C2(n7721), .A(n9892), .B(n7707), .ZN(n7714)
         );
  NOR2_X1 U9486 ( .A1(n7714), .A2(n9351), .ZN(n7660) );
  AOI211_X1 U9487 ( .C1(n9884), .C2(n9011), .A(n7661), .B(n7660), .ZN(n7668)
         );
  XNOR2_X1 U9488 ( .A(n7663), .B(n7662), .ZN(n7666) );
  NAND2_X1 U9489 ( .A1(n9198), .A2(n9433), .ZN(n7664) );
  OAI21_X1 U9490 ( .B1(n7665), .B2(n9467), .A(n7664), .ZN(n8889) );
  AOI21_X1 U9491 ( .B1(n7666), .B2(n9882), .A(n8889), .ZN(n7715) );
  OR2_X1 U9492 ( .A1(n7715), .A2(n9900), .ZN(n7667) );
  OAI211_X1 U9493 ( .C1(n7716), .C2(n9530), .A(n7668), .B(n7667), .ZN(P1_U3278) );
  AOI21_X1 U9494 ( .B1(n7670), .B2(n10084), .A(n7669), .ZN(n7673) );
  MUX2_X1 U9495 ( .A(n7671), .B(n7673), .S(n10121), .Z(n7672) );
  OAI21_X1 U9496 ( .B1(n7698), .B2(n8576), .A(n7672), .ZN(P2_U3475) );
  INV_X1 U9497 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n7674) );
  MUX2_X1 U9498 ( .A(n7674), .B(n7673), .S(n10094), .Z(n7675) );
  OAI21_X1 U9499 ( .B1(n7698), .B2(n8768), .A(n7675), .ZN(P2_U3438) );
  OAI21_X1 U9500 ( .B1(n4277), .B2(n6335), .A(n7676), .ZN(n7677) );
  AOI222_X1 U9501 ( .A1(n8510), .A2(n7677), .B1(n8500), .B2(n8513), .C1(n8332), 
        .C2(n8512), .ZN(n8581) );
  INV_X1 U9502 ( .A(n8316), .ZN(n7678) );
  OAI22_X1 U9503 ( .A1(n9716), .A2(n7679), .B1(n7678), .B2(n9703), .ZN(n7680)
         );
  AOI21_X1 U9504 ( .B1(n8312), .B2(n8425), .A(n7680), .ZN(n7683) );
  NAND2_X1 U9505 ( .A1(n7681), .A2(n6335), .ZN(n8577) );
  NAND3_X1 U9506 ( .A1(n8578), .A2(n8525), .A3(n8577), .ZN(n7682) );
  OAI211_X1 U9507 ( .C1(n8581), .C2(n9719), .A(n7683), .B(n7682), .ZN(P2_U3215) );
  INV_X1 U9508 ( .A(n7684), .ZN(n7685) );
  NAND2_X1 U9509 ( .A1(n7685), .A2(n8334), .ZN(n7686) );
  NAND2_X1 U9510 ( .A1(n7687), .A2(n7686), .ZN(n7690) );
  XNOR2_X1 U9511 ( .A(n7688), .B(n7974), .ZN(n7725) );
  XNOR2_X1 U9512 ( .A(n7725), .B(n8333), .ZN(n7689) );
  OAI211_X1 U9513 ( .C1(n7690), .C2(n7689), .A(n7728), .B(n8283), .ZN(n7697)
         );
  NOR2_X1 U9514 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7691), .ZN(n7797) );
  AOI21_X1 U9515 ( .B1(n8320), .B2(n8332), .A(n7797), .ZN(n7692) );
  OAI21_X1 U9516 ( .B1(n8322), .B2(n7693), .A(n7692), .ZN(n7694) );
  AOI21_X1 U9517 ( .B1(n8291), .B2(n7695), .A(n7694), .ZN(n7696) );
  OAI211_X1 U9518 ( .C1(n7698), .C2(n8323), .A(n7697), .B(n7696), .ZN(P2_U3166) );
  XOR2_X1 U9519 ( .A(n7699), .B(n8940), .Z(n9599) );
  INV_X1 U9520 ( .A(n9599), .ZN(n7713) );
  INV_X1 U9521 ( .A(n8940), .ZN(n7700) );
  XNOR2_X1 U9522 ( .A(n7701), .B(n7700), .ZN(n7702) );
  NAND2_X1 U9523 ( .A1(n7702), .A2(n9882), .ZN(n7705) );
  NAND2_X1 U9524 ( .A1(n9195), .A2(n9431), .ZN(n7704) );
  NAND2_X1 U9525 ( .A1(n9197), .A2(n9433), .ZN(n7703) );
  AND2_X1 U9526 ( .A1(n7704), .A2(n7703), .ZN(n8822) );
  NAND2_X1 U9527 ( .A1(n7705), .A2(n8822), .ZN(n9597) );
  INV_X1 U9528 ( .A(n7739), .ZN(n7706) );
  AOI211_X1 U9529 ( .C1(n8825), .C2(n7707), .A(n9909), .B(n7706), .ZN(n9598)
         );
  NAND2_X1 U9530 ( .A1(n9598), .A2(n9896), .ZN(n7710) );
  INV_X1 U9531 ( .A(n8821), .ZN(n7708) );
  AOI22_X1 U9532 ( .A1(n9523), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n7708), .B2(
        n9886), .ZN(n7709) );
  OAI211_X1 U9533 ( .C1(n4461), .C2(n9526), .A(n7710), .B(n7709), .ZN(n7711)
         );
  AOI21_X1 U9534 ( .B1(n9597), .B2(n9528), .A(n7711), .ZN(n7712) );
  OAI21_X1 U9535 ( .B1(n7713), .B2(n9530), .A(n7712), .ZN(P1_U3277) );
  INV_X1 U9536 ( .A(n9971), .ZN(n9931) );
  OAI211_X1 U9537 ( .C1(n7716), .C2(n9931), .A(n7715), .B(n7714), .ZN(n7717)
         );
  INV_X1 U9538 ( .A(n7717), .ZN(n7719) );
  MUX2_X1 U9539 ( .A(n5348), .B(n7719), .S(n9998), .Z(n7718) );
  OAI21_X1 U9540 ( .B1(n7721), .B2(n9602), .A(n7718), .ZN(P1_U3537) );
  MUX2_X1 U9541 ( .A(n5343), .B(n7719), .S(n9983), .Z(n7720) );
  OAI21_X1 U9542 ( .B1(n7721), .B2(n9645), .A(n7720), .ZN(P1_U3498) );
  INV_X1 U9543 ( .A(n7722), .ZN(n7991) );
  OAI222_X1 U9544 ( .A1(n8777), .A2(n7991), .B1(n7724), .B2(P2_U3151), .C1(
        n7723), .C2(n7747), .ZN(P2_U3266) );
  INV_X1 U9545 ( .A(n7725), .ZN(n7726) );
  NAND2_X1 U9546 ( .A1(n7726), .A2(n8333), .ZN(n7727) );
  NAND2_X1 U9547 ( .A1(n7728), .A2(n7727), .ZN(n7941) );
  XNOR2_X1 U9548 ( .A(n8582), .B(n7961), .ZN(n7940) );
  XNOR2_X1 U9549 ( .A(n7940), .B(n8311), .ZN(n7729) );
  XNOR2_X1 U9550 ( .A(n7941), .B(n7729), .ZN(n7737) );
  AND2_X1 U9551 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7771) );
  AOI21_X1 U9552 ( .B1(n8320), .B2(n8511), .A(n7771), .ZN(n7730) );
  OAI21_X1 U9553 ( .B1(n8322), .B2(n7731), .A(n7730), .ZN(n7734) );
  NOR2_X1 U9554 ( .A1(n7732), .A2(n8323), .ZN(n7733) );
  AOI211_X1 U9555 ( .C1(n7735), .C2(n8291), .A(n7734), .B(n7733), .ZN(n7736)
         );
  OAI21_X1 U9556 ( .B1(n7737), .B2(n8328), .A(n7736), .ZN(P2_U3168) );
  XOR2_X1 U9557 ( .A(n7738), .B(n8943), .Z(n9596) );
  AOI211_X1 U9558 ( .C1(n9594), .C2(n7739), .A(n9909), .B(n9517), .ZN(n9593)
         );
  NOR2_X1 U9559 ( .A1(n4460), .A2(n9526), .ZN(n7741) );
  OAI22_X1 U9560 ( .A1(n9528), .A2(n9280), .B1(n8830), .B2(n9501), .ZN(n7740)
         );
  AOI211_X1 U9561 ( .C1(n9593), .C2(n9896), .A(n7741), .B(n7740), .ZN(n7746)
         );
  OAI211_X1 U9562 ( .C1(n8943), .C2(n7742), .A(n9511), .B(n9882), .ZN(n7744)
         );
  AOI22_X1 U9563 ( .A1(n9196), .A2(n9433), .B1(n9431), .B2(n9194), .ZN(n7743)
         );
  NAND2_X1 U9564 ( .A1(n7744), .A2(n7743), .ZN(n9592) );
  NAND2_X1 U9565 ( .A1(n9592), .A2(n9346), .ZN(n7745) );
  OAI211_X1 U9566 ( .C1(n9596), .C2(n9530), .A(n7746), .B(n7745), .ZN(P1_U3276) );
  INV_X1 U9567 ( .A(n7996), .ZN(n9657) );
  OAI222_X1 U9568 ( .A1(n7747), .A2(n7997), .B1(n8777), .B2(n9657), .C1(
        P2_U3151), .C2(n6117), .ZN(P2_U3265) );
  OAI222_X1 U9569 ( .A1(n7747), .A2(n7751), .B1(n7750), .B2(n7749), .C1(n7748), 
        .C2(P2_U3151), .ZN(P2_U3270) );
  AOI21_X1 U9570 ( .B1(n7753), .B2(n7752), .A(n4315), .ZN(n7767) );
  INV_X1 U9571 ( .A(n7754), .ZN(n7756) );
  NAND2_X1 U9572 ( .A1(n7756), .A2(n7755), .ZN(n7758) );
  OAI21_X1 U9573 ( .B1(n8348), .B2(n7758), .A(n5954), .ZN(n7764) );
  INV_X1 U9574 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10129) );
  NAND3_X1 U9575 ( .A1(n7758), .A2(n10006), .A3(n7757), .ZN(n7760) );
  AND2_X1 U9576 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8309) );
  INV_X1 U9577 ( .A(n8309), .ZN(n7759) );
  OAI211_X1 U9578 ( .C1(n10021), .C2(n10129), .A(n7760), .B(n7759), .ZN(n7763)
         );
  OAI21_X1 U9579 ( .B1(n7767), .B2(n9999), .A(n7766), .ZN(P2_U3200) );
  AOI21_X1 U9580 ( .B1(n7770), .B2(n7769), .A(n7768), .ZN(n7787) );
  INV_X1 U9581 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7773) );
  INV_X1 U9582 ( .A(n7771), .ZN(n7772) );
  OAI21_X1 U9583 ( .B1(n10021), .B2(n7773), .A(n7772), .ZN(n7779) );
  AOI21_X1 U9584 ( .B1(n7776), .B2(n7775), .A(n7774), .ZN(n7777) );
  NOR2_X1 U9585 ( .A1(n10014), .A2(n7777), .ZN(n7778) );
  AOI211_X1 U9586 ( .C1(n8369), .C2(n7780), .A(n7779), .B(n7778), .ZN(n7786)
         );
  OAI21_X1 U9587 ( .B1(n7783), .B2(n7782), .A(n7781), .ZN(n7784) );
  NAND2_X1 U9588 ( .A1(n7784), .A2(n10006), .ZN(n7785) );
  OAI211_X1 U9589 ( .C1(n7787), .C2(n9999), .A(n7786), .B(n7785), .ZN(P2_U3199) );
  AOI21_X1 U9590 ( .B1(n7790), .B2(n7789), .A(n7788), .ZN(n7808) );
  INV_X1 U9591 ( .A(n7791), .ZN(n7792) );
  NAND2_X1 U9592 ( .A1(n7793), .A2(n7792), .ZN(n7794) );
  XNOR2_X1 U9593 ( .A(n7795), .B(n7794), .ZN(n7806) );
  INV_X1 U9594 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U9595 ( .A1(n8369), .A2(n7796), .ZN(n7799) );
  INV_X1 U9596 ( .A(n7797), .ZN(n7798) );
  OAI211_X1 U9597 ( .C1(n7800), .C2(n10021), .A(n7799), .B(n7798), .ZN(n7805)
         );
  AOI21_X1 U9598 ( .B1(n4289), .B2(n7802), .A(n7801), .ZN(n7803) );
  NOR2_X1 U9599 ( .A1(n7803), .A2(n10014), .ZN(n7804) );
  AOI211_X1 U9600 ( .C1(n10006), .C2(n7806), .A(n7805), .B(n7804), .ZN(n7807)
         );
  OAI21_X1 U9601 ( .B1(n7808), .B2(n9999), .A(n7807), .ZN(P2_U3198) );
  AOI21_X1 U9602 ( .B1(n7811), .B2(n7810), .A(n7809), .ZN(n7827) );
  INV_X1 U9603 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7818) );
  AOI21_X1 U9604 ( .B1(n7814), .B2(n7813), .A(n7812), .ZN(n7815) );
  OR2_X1 U9605 ( .A1(n7815), .A2(n8357), .ZN(n7816) );
  OAI211_X1 U9606 ( .C1(n10021), .C2(n7818), .A(n7817), .B(n7816), .ZN(n7824)
         );
  AOI21_X1 U9607 ( .B1(n7821), .B2(n7820), .A(n7819), .ZN(n7822) );
  NOR2_X1 U9608 ( .A1(n7822), .A2(n10014), .ZN(n7823) );
  AOI211_X1 U9609 ( .C1(n8369), .C2(n7825), .A(n7824), .B(n7823), .ZN(n7826)
         );
  OAI21_X1 U9610 ( .B1(n7827), .B2(n9999), .A(n7826), .ZN(P2_U3196) );
  AOI21_X1 U9611 ( .B1(n9718), .B2(n7829), .A(n7828), .ZN(n7845) );
  INV_X1 U9612 ( .A(n7830), .ZN(n7836) );
  AOI21_X1 U9613 ( .B1(n7833), .B2(n7832), .A(n7831), .ZN(n7834) );
  OR2_X1 U9614 ( .A1(n7834), .A2(n8357), .ZN(n7835) );
  OAI211_X1 U9615 ( .C1(n10021), .C2(n7837), .A(n7836), .B(n7835), .ZN(n7842)
         );
  AOI21_X1 U9616 ( .B1(n9724), .B2(n7839), .A(n7838), .ZN(n7840) );
  NOR2_X1 U9617 ( .A1(n7840), .A2(n10014), .ZN(n7841) );
  AOI211_X1 U9618 ( .C1(n8369), .C2(n7843), .A(n7842), .B(n7841), .ZN(n7844)
         );
  OAI21_X1 U9619 ( .B1(n7845), .B2(n9999), .A(n7844), .ZN(P2_U3195) );
  AOI21_X1 U9620 ( .B1(n7848), .B2(n7847), .A(n7846), .ZN(n7864) );
  INV_X1 U9621 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7856) );
  INV_X1 U9622 ( .A(n7849), .ZN(n7855) );
  AOI21_X1 U9623 ( .B1(n7852), .B2(n7851), .A(n7850), .ZN(n7853) );
  OR2_X1 U9624 ( .A1(n7853), .A2(n8357), .ZN(n7854) );
  OAI211_X1 U9625 ( .C1(n10021), .C2(n7856), .A(n7855), .B(n7854), .ZN(n7861)
         );
  AOI21_X1 U9626 ( .B1(n4350), .B2(n7858), .A(n7857), .ZN(n7859) );
  NOR2_X1 U9627 ( .A1(n7859), .A2(n10014), .ZN(n7860) );
  AOI211_X1 U9628 ( .C1(n8369), .C2(n7862), .A(n7861), .B(n7860), .ZN(n7863)
         );
  OAI21_X1 U9629 ( .B1(n7864), .B2(n9999), .A(n7863), .ZN(P2_U3194) );
  AOI21_X1 U9630 ( .B1(n7867), .B2(n7866), .A(n7865), .ZN(n7883) );
  AOI21_X1 U9631 ( .B1(n7870), .B2(n7869), .A(n7868), .ZN(n7875) );
  INV_X1 U9632 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7871) );
  OR2_X1 U9633 ( .A1(n10021), .A2(n7871), .ZN(n7874) );
  INV_X1 U9634 ( .A(n7872), .ZN(n7873) );
  OAI211_X1 U9635 ( .C1(n7875), .C2(n8357), .A(n7874), .B(n7873), .ZN(n7880)
         );
  AOI21_X1 U9636 ( .B1(n10117), .B2(n7877), .A(n7876), .ZN(n7878) );
  NOR2_X1 U9637 ( .A1(n7878), .A2(n10014), .ZN(n7879) );
  AOI211_X1 U9638 ( .C1(n8369), .C2(n7881), .A(n7880), .B(n7879), .ZN(n7882)
         );
  OAI21_X1 U9639 ( .B1(n7883), .B2(n9999), .A(n7882), .ZN(P2_U3193) );
  AOI21_X1 U9640 ( .B1(n7885), .B2(n7884), .A(n4351), .ZN(n7902) );
  INV_X1 U9641 ( .A(n7886), .ZN(n7887) );
  OAI21_X1 U9642 ( .B1(n10021), .B2(n7888), .A(n7887), .ZN(n7894) );
  AOI21_X1 U9643 ( .B1(n7891), .B2(n7890), .A(n7889), .ZN(n7892) );
  NOR2_X1 U9644 ( .A1(n7892), .A2(n10014), .ZN(n7893) );
  AOI211_X1 U9645 ( .C1(n8369), .C2(n7895), .A(n7894), .B(n7893), .ZN(n7901)
         );
  AOI21_X1 U9646 ( .B1(n7898), .B2(n7897), .A(n7896), .ZN(n7899) );
  OR2_X1 U9647 ( .A1(n7899), .A2(n8357), .ZN(n7900) );
  OAI211_X1 U9648 ( .C1(n7902), .C2(n9999), .A(n7901), .B(n7900), .ZN(P2_U3192) );
  AOI21_X1 U9649 ( .B1(n7905), .B2(n7904), .A(n7903), .ZN(n7922) );
  OAI21_X1 U9650 ( .B1(n7908), .B2(n7907), .A(n7906), .ZN(n7909) );
  NAND2_X1 U9651 ( .A1(n7909), .A2(n10006), .ZN(n7921) );
  INV_X1 U9652 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7912) );
  INV_X1 U9653 ( .A(n7910), .ZN(n7911) );
  OAI21_X1 U9654 ( .B1(n10021), .B2(n7912), .A(n7911), .ZN(n7918) );
  AOI21_X1 U9655 ( .B1(n7915), .B2(n7914), .A(n7913), .ZN(n7916) );
  NOR2_X1 U9656 ( .A1(n7916), .A2(n10014), .ZN(n7917) );
  AOI211_X1 U9657 ( .C1(n8369), .C2(n7919), .A(n7918), .B(n7917), .ZN(n7920)
         );
  OAI211_X1 U9658 ( .C1(n7922), .C2(n9999), .A(n7921), .B(n7920), .ZN(P2_U3190) );
  AOI21_X1 U9659 ( .B1(n7925), .B2(n7924), .A(n7923), .ZN(n7939) );
  XNOR2_X1 U9660 ( .A(n7927), .B(n7926), .ZN(n7928) );
  NAND2_X1 U9661 ( .A1(n7928), .A2(n10006), .ZN(n7938) );
  INV_X1 U9662 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7930) );
  OAI21_X1 U9663 ( .B1(n10021), .B2(n7930), .A(n7929), .ZN(n7935) );
  AOI21_X1 U9664 ( .B1(n7932), .B2(n10109), .A(n7931), .ZN(n7933) );
  NOR2_X1 U9665 ( .A1(n7933), .A2(n10014), .ZN(n7934) );
  AOI211_X1 U9666 ( .C1(n8369), .C2(n7936), .A(n7935), .B(n7934), .ZN(n7937)
         );
  OAI211_X1 U9667 ( .C1(n7939), .C2(n9999), .A(n7938), .B(n7937), .ZN(P2_U3189) );
  XNOR2_X1 U9668 ( .A(n8312), .B(n7974), .ZN(n7943) );
  NAND2_X1 U9669 ( .A1(n7943), .A2(n7942), .ZN(n7946) );
  INV_X1 U9670 ( .A(n7943), .ZN(n7944) );
  NAND2_X1 U9671 ( .A1(n7944), .A2(n8511), .ZN(n7945) );
  NAND2_X1 U9672 ( .A1(n7946), .A2(n7945), .ZN(n8308) );
  NAND2_X1 U9673 ( .A1(n8305), .A2(n7946), .ZN(n7950) );
  INV_X1 U9674 ( .A(n7950), .ZN(n7948) );
  XNOR2_X1 U9675 ( .A(n8236), .B(n7974), .ZN(n7949) );
  INV_X1 U9676 ( .A(n7949), .ZN(n7947) );
  NAND2_X1 U9677 ( .A1(n7950), .A2(n7949), .ZN(n8279) );
  XNOR2_X1 U9678 ( .A(n8278), .B(n7974), .ZN(n7952) );
  NAND2_X1 U9679 ( .A1(n7952), .A2(n8488), .ZN(n8247) );
  INV_X1 U9680 ( .A(n7952), .ZN(n7953) );
  NAND2_X1 U9681 ( .A1(n7953), .A2(n8514), .ZN(n7954) );
  AND2_X1 U9682 ( .A1(n8247), .A2(n7954), .ZN(n8280) );
  NAND2_X1 U9683 ( .A1(n8246), .A2(n8247), .ZN(n7955) );
  XNOR2_X1 U9684 ( .A(n8245), .B(n7974), .ZN(n7956) );
  XNOR2_X1 U9685 ( .A(n7956), .B(n8501), .ZN(n8248) );
  NAND2_X1 U9686 ( .A1(n7955), .A2(n8248), .ZN(n8250) );
  NAND2_X1 U9687 ( .A1(n7956), .A2(n8288), .ZN(n7957) );
  XNOR2_X1 U9688 ( .A(n8029), .B(n7974), .ZN(n8294) );
  INV_X1 U9689 ( .A(n8294), .ZN(n7958) );
  NAND2_X1 U9690 ( .A1(n7958), .A2(n8253), .ZN(n7960) );
  AND2_X1 U9691 ( .A1(n8294), .A2(n8489), .ZN(n7959) );
  XNOR2_X1 U9692 ( .A(n8273), .B(n7974), .ZN(n8269) );
  XNOR2_X1 U9693 ( .A(n7962), .B(n7961), .ZN(n8266) );
  INV_X1 U9694 ( .A(n8266), .ZN(n7963) );
  OAI22_X1 U9695 ( .A1(n8269), .A2(n8464), .B1(n8300), .B2(n7963), .ZN(n7967)
         );
  OAI21_X1 U9696 ( .B1(n8266), .B2(n8475), .A(n8331), .ZN(n7965) );
  NOR2_X1 U9697 ( .A1(n8331), .A2(n8475), .ZN(n7964) );
  AOI22_X1 U9698 ( .A1(n8269), .A2(n7965), .B1(n7964), .B2(n7963), .ZN(n7966)
         );
  XNOR2_X1 U9699 ( .A(n8261), .B(n7974), .ZN(n7968) );
  XNOR2_X1 U9700 ( .A(n7968), .B(n8455), .ZN(n8259) );
  INV_X1 U9701 ( .A(n7968), .ZN(n7969) );
  XNOR2_X1 U9702 ( .A(n8743), .B(n7974), .ZN(n7970) );
  XNOR2_X1 U9703 ( .A(n7970), .B(n8405), .ZN(n8319) );
  XNOR2_X1 U9704 ( .A(n8414), .B(n7974), .ZN(n7971) );
  NAND2_X1 U9705 ( .A1(n7971), .A2(n8391), .ZN(n7972) );
  OAI21_X1 U9706 ( .B1(n7971), .B2(n8391), .A(n7972), .ZN(n7983) );
  INV_X1 U9707 ( .A(n7972), .ZN(n7973) );
  NOR2_X1 U9708 ( .A1(n7982), .A2(n7973), .ZN(n7976) );
  XNOR2_X1 U9709 ( .A(n8395), .B(n7974), .ZN(n7975) );
  XNOR2_X1 U9710 ( .A(n7976), .B(n7975), .ZN(n7981) );
  AOI22_X1 U9711 ( .A1(n8297), .A2(n8391), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7977) );
  OAI21_X1 U9712 ( .B1(n8015), .B2(n8299), .A(n7977), .ZN(n7979) );
  NOR2_X1 U9713 ( .A1(n8399), .A2(n8323), .ZN(n7978) );
  AOI211_X1 U9714 ( .C1(n8397), .C2(n8326), .A(n7979), .B(n7978), .ZN(n7980)
         );
  OAI21_X1 U9715 ( .B1(n7981), .B2(n8328), .A(n7980), .ZN(P2_U3160) );
  AOI22_X1 U9716 ( .A1(n8320), .A2(n8404), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7987) );
  OAI21_X1 U9717 ( .B1(n8438), .B2(n8322), .A(n7987), .ZN(n7988) );
  AOI21_X1 U9718 ( .B1(n8291), .B2(n8412), .A(n7988), .ZN(n7989) );
  OAI211_X1 U9719 ( .C1(n8414), .C2(n8323), .A(n7990), .B(n7989), .ZN(P2_U3154) );
  OAI222_X1 U9720 ( .A1(n7993), .A2(n7992), .B1(P1_U3086), .B2(n4281), .C1(
        n7991), .C2(n9658), .ZN(P1_U3326) );
  INV_X1 U9721 ( .A(n8017), .ZN(n7994) );
  AOI21_X1 U9722 ( .B1(n7995), .B2(n8177), .A(n7994), .ZN(n8006) );
  NAND2_X1 U9723 ( .A1(n7996), .A2(n6219), .ZN(n7999) );
  OR2_X1 U9724 ( .A1(n8001), .A2(n7997), .ZN(n7998) );
  NAND2_X1 U9725 ( .A1(n8591), .A2(n8004), .ZN(n8216) );
  INV_X1 U9726 ( .A(n8216), .ZN(n8005) );
  NAND2_X1 U9727 ( .A1(n8772), .A2(n6219), .ZN(n8003) );
  OR2_X1 U9728 ( .A1(n8001), .A2(n8000), .ZN(n8002) );
  OAI22_X1 U9729 ( .A1(n8006), .A2(n8005), .B1(n8376), .B2(n8217), .ZN(n8013)
         );
  NAND2_X1 U9730 ( .A1(n6170), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U9731 ( .A1(n6437), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8008) );
  NAND2_X1 U9732 ( .A1(n6159), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8007) );
  INV_X1 U9733 ( .A(n8373), .ZN(n8330) );
  OAI21_X1 U9734 ( .B1(n8330), .B2(n8591), .A(n8376), .ZN(n8012) );
  AOI21_X1 U9735 ( .B1(n8013), .B2(n8012), .A(n8011), .ZN(n8014) );
  NOR2_X1 U9736 ( .A1(n8015), .A2(n8137), .ZN(n8390) );
  NAND2_X1 U9737 ( .A1(n8179), .A2(n8176), .ZN(n8016) );
  NAND2_X1 U9738 ( .A1(n8017), .A2(n8016), .ZN(n8019) );
  INV_X1 U9739 ( .A(n8390), .ZN(n8018) );
  NAND2_X1 U9740 ( .A1(n8019), .A2(n8018), .ZN(n8175) );
  OR2_X1 U9741 ( .A1(n8414), .A2(n8391), .ZN(n8021) );
  MUX2_X1 U9742 ( .A(n8021), .B(n8020), .S(n8137), .Z(n8026) );
  MUX2_X1 U9743 ( .A(n8023), .B(n8022), .S(n8176), .Z(n8024) );
  NAND2_X1 U9744 ( .A1(n8024), .A2(n8410), .ZN(n8025) );
  NAND2_X1 U9745 ( .A1(n8026), .A2(n8025), .ZN(n8169) );
  INV_X1 U9746 ( .A(n8027), .ZN(n8028) );
  NOR2_X1 U9747 ( .A1(n8186), .A2(n8028), .ZN(n8032) );
  NAND2_X1 U9748 ( .A1(n8029), .A2(n8489), .ZN(n8030) );
  AND2_X1 U9749 ( .A1(n8184), .A2(n8030), .ZN(n8031) );
  MUX2_X1 U9750 ( .A(n8032), .B(n8031), .S(n8137), .Z(n8156) );
  INV_X1 U9751 ( .A(n8498), .ZN(n8504) );
  AOI22_X1 U9752 ( .A1(n8504), .A2(n8033), .B1(n8176), .B2(n8145), .ZN(n8150)
         );
  AOI21_X1 U9753 ( .B1(n8133), .B2(n8034), .A(n8137), .ZN(n8140) );
  NAND2_X1 U9754 ( .A1(n8045), .A2(n6804), .ZN(n8035) );
  NAND2_X1 U9755 ( .A1(n8036), .A2(n8035), .ZN(n8037) );
  NAND2_X1 U9756 ( .A1(n8037), .A2(n8137), .ZN(n8044) );
  INV_X1 U9757 ( .A(n8038), .ZN(n8039) );
  OAI21_X1 U9758 ( .B1(n8044), .B2(n8039), .A(n8137), .ZN(n8041) );
  MUX2_X1 U9759 ( .A(n8137), .B(n8041), .S(n8040), .Z(n8047) );
  NAND3_X1 U9760 ( .A1(n6449), .A2(n8045), .A3(n8044), .ZN(n8046) );
  NAND3_X1 U9761 ( .A1(n8047), .A2(n8042), .A3(n8046), .ZN(n8056) );
  NAND2_X1 U9762 ( .A1(n8345), .A2(n8048), .ZN(n8058) );
  NAND2_X1 U9763 ( .A1(n8346), .A2(n8049), .ZN(n8050) );
  NAND2_X1 U9764 ( .A1(n8058), .A2(n8050), .ZN(n8053) );
  NAND2_X1 U9765 ( .A1(n8067), .A2(n8051), .ZN(n8052) );
  MUX2_X1 U9766 ( .A(n8053), .B(n8052), .S(n8137), .Z(n8054) );
  INV_X1 U9767 ( .A(n8054), .ZN(n8055) );
  NAND2_X1 U9768 ( .A1(n8056), .A2(n8055), .ZN(n8057) );
  NAND2_X1 U9769 ( .A1(n8057), .A2(n8189), .ZN(n8071) );
  INV_X1 U9770 ( .A(n8058), .ZN(n8061) );
  OAI211_X1 U9771 ( .C1(n8071), .C2(n8061), .A(n8060), .B(n8059), .ZN(n8066)
         );
  AND2_X1 U9772 ( .A1(n8062), .A2(n8068), .ZN(n8065) );
  INV_X1 U9773 ( .A(n8063), .ZN(n8064) );
  AOI21_X1 U9774 ( .B1(n8066), .B2(n8065), .A(n8064), .ZN(n8076) );
  INV_X1 U9775 ( .A(n8067), .ZN(n8070) );
  OAI211_X1 U9776 ( .C1(n8071), .C2(n8070), .A(n8069), .B(n8068), .ZN(n8074)
         );
  AOI21_X1 U9777 ( .B1(n8074), .B2(n8073), .A(n8072), .ZN(n8075) );
  MUX2_X1 U9778 ( .A(n8076), .B(n8075), .S(n8176), .Z(n8077) );
  NAND2_X1 U9779 ( .A1(n8077), .A2(n8194), .ZN(n8082) );
  AND2_X1 U9780 ( .A1(n8085), .A2(n8078), .ZN(n8079) );
  MUX2_X1 U9781 ( .A(n8080), .B(n8079), .S(n8176), .Z(n8081) );
  NAND2_X1 U9782 ( .A1(n8082), .A2(n8081), .ZN(n8096) );
  NAND2_X1 U9783 ( .A1(n8084), .A2(n8083), .ZN(n8087) );
  NAND2_X1 U9784 ( .A1(n8089), .A2(n8085), .ZN(n8086) );
  MUX2_X1 U9785 ( .A(n8087), .B(n8086), .S(n8137), .Z(n8088) );
  INV_X1 U9786 ( .A(n8088), .ZN(n8095) );
  AND2_X1 U9787 ( .A1(n8090), .A2(n8089), .ZN(n8092) );
  MUX2_X1 U9788 ( .A(n8092), .B(n8091), .S(n8137), .Z(n8093) );
  NAND2_X1 U9789 ( .A1(n8202), .A2(n8093), .ZN(n8094) );
  AOI21_X1 U9790 ( .B1(n8096), .B2(n8095), .A(n8094), .ZN(n8107) );
  INV_X1 U9791 ( .A(n8097), .ZN(n8098) );
  NAND2_X1 U9792 ( .A1(n8099), .A2(n8098), .ZN(n8100) );
  NAND2_X1 U9793 ( .A1(n8100), .A2(n8101), .ZN(n8105) );
  INV_X1 U9794 ( .A(n8101), .ZN(n8102) );
  NOR2_X1 U9795 ( .A1(n8103), .A2(n8102), .ZN(n8104) );
  MUX2_X1 U9796 ( .A(n8105), .B(n8104), .S(n8137), .Z(n8106) );
  OAI21_X1 U9797 ( .B1(n8107), .B2(n8106), .A(n8203), .ZN(n8111) );
  MUX2_X1 U9798 ( .A(n8109), .B(n8108), .S(n8137), .Z(n8110) );
  NAND3_X1 U9799 ( .A1(n8111), .A2(n9707), .A3(n8110), .ZN(n8117) );
  NAND2_X1 U9800 ( .A1(n8113), .A2(n8112), .ZN(n8115) );
  MUX2_X1 U9801 ( .A(n8115), .B(n8114), .S(n8137), .Z(n8116) );
  NAND3_X1 U9802 ( .A1(n8117), .A2(n8205), .A3(n8116), .ZN(n8122) );
  MUX2_X1 U9803 ( .A(n8119), .B(n8118), .S(n8176), .Z(n8120) );
  NAND3_X1 U9804 ( .A1(n8122), .A2(n8121), .A3(n8120), .ZN(n8127) );
  MUX2_X1 U9805 ( .A(n8124), .B(n8123), .S(n8176), .Z(n8125) );
  NAND3_X1 U9806 ( .A1(n8127), .A2(n8126), .A3(n8125), .ZN(n8131) );
  MUX2_X1 U9807 ( .A(n8129), .B(n8128), .S(n8137), .Z(n8130) );
  NAND3_X1 U9808 ( .A1(n8131), .A2(n6459), .A3(n8130), .ZN(n8136) );
  OAI21_X1 U9809 ( .B1(n8311), .B2(n8582), .A(n8517), .ZN(n8132) );
  NAND2_X1 U9810 ( .A1(n8132), .A2(n8137), .ZN(n8135) );
  INV_X1 U9811 ( .A(n8133), .ZN(n8134) );
  AOI21_X1 U9812 ( .B1(n8136), .B2(n8135), .A(n8134), .ZN(n8139) );
  OAI22_X1 U9813 ( .A1(n8140), .A2(n8139), .B1(n8138), .B2(n8137), .ZN(n8142)
         );
  MUX2_X1 U9814 ( .A(n8137), .B(n8142), .S(n8141), .Z(n8143) );
  INV_X1 U9815 ( .A(n8143), .ZN(n8149) );
  AND2_X1 U9816 ( .A1(n8151), .A2(n8144), .ZN(n8147) );
  AND2_X1 U9817 ( .A1(n8152), .A2(n8145), .ZN(n8146) );
  MUX2_X1 U9818 ( .A(n8147), .B(n8146), .S(n8137), .Z(n8148) );
  OAI21_X1 U9819 ( .B1(n8150), .B2(n8149), .A(n8148), .ZN(n8154) );
  MUX2_X1 U9820 ( .A(n8152), .B(n8151), .S(n8137), .Z(n8153) );
  NAND3_X1 U9821 ( .A1(n8154), .A2(n8478), .A3(n8153), .ZN(n8155) );
  AND2_X1 U9822 ( .A1(n8156), .A2(n8155), .ZN(n8164) );
  INV_X1 U9823 ( .A(n8186), .ZN(n8157) );
  NAND2_X1 U9824 ( .A1(n8160), .A2(n8157), .ZN(n8159) );
  NAND2_X1 U9825 ( .A1(n8161), .A2(n8184), .ZN(n8158) );
  MUX2_X1 U9826 ( .A(n8159), .B(n8158), .S(n8176), .Z(n8163) );
  MUX2_X1 U9827 ( .A(n8161), .B(n8160), .S(n8176), .Z(n8162) );
  OAI211_X1 U9828 ( .C1(n8164), .C2(n8163), .A(n8447), .B(n8162), .ZN(n8167)
         );
  MUX2_X1 U9829 ( .A(n8427), .B(n8165), .S(n8176), .Z(n8166) );
  NAND4_X1 U9830 ( .A1(n8410), .A2(n8428), .A3(n8167), .A4(n8166), .ZN(n8168)
         );
  NAND2_X1 U9831 ( .A1(n8169), .A2(n8168), .ZN(n8170) );
  AND2_X1 U9832 ( .A1(n8175), .A2(n8170), .ZN(n8173) );
  INV_X1 U9833 ( .A(n8173), .ZN(n8172) );
  MUX2_X1 U9834 ( .A(n8404), .B(n8533), .S(n8137), .Z(n8174) );
  INV_X1 U9835 ( .A(n8174), .ZN(n8171) );
  INV_X1 U9836 ( .A(n8180), .ZN(n8181) );
  NAND2_X1 U9837 ( .A1(n8180), .A2(n8216), .ZN(n8182) );
  INV_X1 U9838 ( .A(n8184), .ZN(n8185) );
  NOR2_X1 U9839 ( .A1(n8186), .A2(n8185), .ZN(n8466) );
  INV_X1 U9840 ( .A(n8187), .ZN(n8491) );
  NAND4_X1 U9841 ( .A1(n6449), .A2(n8189), .A3(n10023), .A4(n8188), .ZN(n8192)
         );
  NAND2_X1 U9842 ( .A1(n8042), .A2(n8190), .ZN(n8191) );
  NOR2_X1 U9843 ( .A1(n8192), .A2(n8191), .ZN(n8196) );
  NAND4_X1 U9844 ( .A1(n8196), .A2(n8195), .A3(n8194), .A4(n8193), .ZN(n8199)
         );
  NOR3_X1 U9845 ( .A1(n8199), .A2(n8198), .A3(n8197), .ZN(n8201) );
  AND4_X1 U9846 ( .A1(n8203), .A2(n8202), .A3(n8201), .A4(n8200), .ZN(n8204)
         );
  NAND3_X1 U9847 ( .A1(n8205), .A2(n8204), .A3(n9707), .ZN(n8206) );
  NOR3_X1 U9848 ( .A1(n8208), .A2(n8207), .A3(n8206), .ZN(n8209) );
  NAND4_X1 U9849 ( .A1(n8519), .A2(n8210), .A3(n8209), .A4(n6459), .ZN(n8211)
         );
  NOR2_X1 U9850 ( .A1(n8498), .A2(n8211), .ZN(n8212) );
  NAND4_X1 U9851 ( .A1(n8466), .A2(n8491), .A3(n8212), .A4(n8478), .ZN(n8213)
         );
  NOR2_X1 U9852 ( .A1(n8436), .A2(n8213), .ZN(n8214) );
  NAND4_X1 U9853 ( .A1(n8410), .A2(n8428), .A3(n8458), .A4(n8214), .ZN(n8215)
         );
  NOR2_X1 U9854 ( .A1(n8395), .A2(n8215), .ZN(n8218) );
  NAND2_X1 U9855 ( .A1(n8220), .A2(n4849), .ZN(n8222) );
  XNOR2_X1 U9856 ( .A(n8222), .B(n8221), .ZN(n8230) );
  NOR3_X1 U9857 ( .A1(n8225), .A2(n8224), .A3(n8223), .ZN(n8228) );
  OAI21_X1 U9858 ( .B1(n8229), .B2(n8226), .A(P2_B_REG_SCAN_IN), .ZN(n8227) );
  OAI22_X1 U9859 ( .A1(n8230), .A2(n8229), .B1(n8228), .B2(n8227), .ZN(
        P2_U3296) );
  XNOR2_X1 U9860 ( .A(n8267), .B(n8266), .ZN(n8268) );
  XNOR2_X1 U9861 ( .A(n8268), .B(n8300), .ZN(n8235) );
  AOI22_X1 U9862 ( .A1(n8253), .A2(n8297), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8231) );
  OAI21_X1 U9863 ( .B1(n8464), .B2(n8299), .A(n8231), .ZN(n8233) );
  NOR2_X1 U9864 ( .A1(n8752), .A2(n8323), .ZN(n8232) );
  AOI211_X1 U9865 ( .C1(n8467), .C2(n8326), .A(n8233), .B(n8232), .ZN(n8234)
         );
  OAI21_X1 U9866 ( .B1(n8235), .B2(n8328), .A(n8234), .ZN(P2_U3156) );
  INV_X1 U9867 ( .A(n8236), .ZN(n8769) );
  OAI21_X1 U9868 ( .B1(n8286), .B2(n8238), .A(n8237), .ZN(n8239) );
  NAND2_X1 U9869 ( .A1(n8239), .A2(n8283), .ZN(n8244) );
  NAND2_X1 U9870 ( .A1(n8297), .A2(n8511), .ZN(n8241) );
  OAI211_X1 U9871 ( .C1(n8488), .C2(n8299), .A(n8241), .B(n8240), .ZN(n8242)
         );
  AOI21_X1 U9872 ( .B1(n8291), .B2(n8520), .A(n8242), .ZN(n8243) );
  OAI211_X1 U9873 ( .C1(n8769), .C2(n8323), .A(n8244), .B(n8243), .ZN(P2_U3159) );
  INV_X1 U9874 ( .A(n8245), .ZN(n8760) );
  INV_X1 U9875 ( .A(n8246), .ZN(n8284) );
  INV_X1 U9876 ( .A(n8247), .ZN(n8249) );
  NOR3_X1 U9877 ( .A1(n8284), .A2(n8249), .A3(n8248), .ZN(n8252) );
  INV_X1 U9878 ( .A(n8250), .ZN(n8251) );
  OAI21_X1 U9879 ( .B1(n8252), .B2(n8251), .A(n8283), .ZN(n8257) );
  AOI22_X1 U9880 ( .A1(n8253), .A2(n8320), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8254) );
  OAI21_X1 U9881 ( .B1(n8488), .B2(n8322), .A(n8254), .ZN(n8255) );
  AOI21_X1 U9882 ( .B1(n8492), .B2(n8326), .A(n8255), .ZN(n8256) );
  OAI211_X1 U9883 ( .C1(n8760), .C2(n8323), .A(n8257), .B(n8256), .ZN(P2_U3163) );
  XOR2_X1 U9884 ( .A(n8259), .B(n8258), .Z(n8265) );
  AOI22_X1 U9885 ( .A1(n8320), .A2(n8405), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8260) );
  OAI21_X1 U9886 ( .B1(n8464), .B2(n8322), .A(n8260), .ZN(n8263) );
  NOR2_X1 U9887 ( .A1(n8261), .A2(n8323), .ZN(n8262) );
  AOI211_X1 U9888 ( .C1(n8443), .C2(n8326), .A(n8263), .B(n8262), .ZN(n8264)
         );
  OAI21_X1 U9889 ( .B1(n8265), .B2(n8328), .A(n8264), .ZN(P2_U3165) );
  OAI22_X1 U9890 ( .A1(n8268), .A2(n8475), .B1(n8267), .B2(n8266), .ZN(n8271)
         );
  XNOR2_X1 U9891 ( .A(n8269), .B(n8464), .ZN(n8270) );
  XNOR2_X1 U9892 ( .A(n8271), .B(n8270), .ZN(n8277) );
  AOI22_X1 U9893 ( .A1(n8475), .A2(n8297), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8272) );
  OAI21_X1 U9894 ( .B1(n8455), .B2(n8299), .A(n8272), .ZN(n8275) );
  INV_X1 U9895 ( .A(n8273), .ZN(n8748) );
  NOR2_X1 U9896 ( .A1(n8748), .A2(n8323), .ZN(n8274) );
  AOI211_X1 U9897 ( .C1(n8457), .C2(n8326), .A(n8275), .B(n8274), .ZN(n8276)
         );
  OAI21_X1 U9898 ( .B1(n8277), .B2(n8328), .A(n8276), .ZN(P2_U3169) );
  INV_X1 U9899 ( .A(n8278), .ZN(n8764) );
  INV_X1 U9900 ( .A(n8237), .ZN(n8282) );
  INV_X1 U9901 ( .A(n8279), .ZN(n8281) );
  NOR3_X1 U9902 ( .A1(n8282), .A2(n8281), .A3(n8280), .ZN(n8285) );
  OAI21_X1 U9903 ( .B1(n8285), .B2(n8284), .A(n8283), .ZN(n8293) );
  NOR2_X1 U9904 ( .A1(n8322), .A2(n8286), .ZN(n8290) );
  OAI22_X1 U9905 ( .A1(n8288), .A2(n8299), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8287), .ZN(n8289) );
  AOI211_X1 U9906 ( .C1(n8291), .C2(n8505), .A(n8290), .B(n8289), .ZN(n8292)
         );
  OAI211_X1 U9907 ( .C1(n8764), .C2(n8323), .A(n8293), .B(n8292), .ZN(P2_U3173) );
  XNOR2_X1 U9908 ( .A(n8294), .B(n8489), .ZN(n8295) );
  XNOR2_X1 U9909 ( .A(n8296), .B(n8295), .ZN(n8304) );
  AOI22_X1 U9910 ( .A1(n8501), .A2(n8297), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8298) );
  OAI21_X1 U9911 ( .B1(n8300), .B2(n8299), .A(n8298), .ZN(n8302) );
  NOR2_X1 U9912 ( .A1(n8756), .A2(n8323), .ZN(n8301) );
  AOI211_X1 U9913 ( .C1(n8481), .C2(n8326), .A(n8302), .B(n8301), .ZN(n8303)
         );
  OAI21_X1 U9914 ( .B1(n8304), .B2(n8328), .A(n8303), .ZN(P2_U3175) );
  INV_X1 U9915 ( .A(n8305), .ZN(n8306) );
  AOI21_X1 U9916 ( .B1(n8308), .B2(n8307), .A(n8306), .ZN(n8318) );
  AOI21_X1 U9917 ( .B1(n8320), .B2(n8500), .A(n8309), .ZN(n8310) );
  OAI21_X1 U9918 ( .B1(n8322), .B2(n8311), .A(n8310), .ZN(n8315) );
  NAND2_X1 U9919 ( .A1(n8312), .A2(n10028), .ZN(n8580) );
  NOR2_X1 U9920 ( .A1(n8580), .A2(n8313), .ZN(n8314) );
  AOI211_X1 U9921 ( .C1(n8316), .C2(n8326), .A(n8315), .B(n8314), .ZN(n8317)
         );
  OAI21_X1 U9922 ( .B1(n8318), .B2(n8328), .A(n8317), .ZN(P2_U3178) );
  AOI22_X1 U9923 ( .A1(n8320), .A2(n8391), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8321) );
  OAI21_X1 U9924 ( .B1(n8455), .B2(n8322), .A(n8321), .ZN(n8325) );
  NOR2_X1 U9925 ( .A1(n8743), .A2(n8323), .ZN(n8324) );
  AOI211_X1 U9926 ( .C1(n8421), .C2(n8326), .A(n8325), .B(n8324), .ZN(n8327)
         );
  OAI21_X1 U9927 ( .B1(n8329), .B2(n8328), .A(n8327), .ZN(P2_U3180) );
  MUX2_X1 U9928 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8330), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9929 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8404), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9930 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8391), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9931 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8405), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9932 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8331), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9933 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8501), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9934 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8514), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9935 ( .A(n8500), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8348), .Z(
        P2_U3510) );
  MUX2_X1 U9936 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8511), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9937 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8332), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9938 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8333), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9939 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8334), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9940 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8335), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9941 ( .A(n8336), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8348), .Z(
        P2_U3504) );
  MUX2_X1 U9942 ( .A(n8337), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8348), .Z(
        P2_U3503) );
  MUX2_X1 U9943 ( .A(n8338), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8348), .Z(
        P2_U3502) );
  MUX2_X1 U9944 ( .A(n8339), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8348), .Z(
        P2_U3501) );
  MUX2_X1 U9945 ( .A(n8340), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8348), .Z(
        P2_U3500) );
  MUX2_X1 U9946 ( .A(n8341), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8348), .Z(
        P2_U3499) );
  MUX2_X1 U9947 ( .A(n8342), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8348), .Z(
        P2_U3498) );
  MUX2_X1 U9948 ( .A(n6453), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8348), .Z(
        P2_U3497) );
  MUX2_X1 U9949 ( .A(n8343), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8348), .Z(
        P2_U3496) );
  MUX2_X1 U9950 ( .A(n8344), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8348), .Z(
        P2_U3495) );
  MUX2_X1 U9951 ( .A(n8345), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8348), .Z(
        P2_U3494) );
  MUX2_X1 U9952 ( .A(n8346), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8348), .Z(
        P2_U3493) );
  MUX2_X1 U9953 ( .A(n8347), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8348), .Z(
        P2_U3492) );
  MUX2_X1 U9954 ( .A(n8349), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8348), .Z(
        P2_U3491) );
  AOI21_X1 U9955 ( .B1(n8352), .B2(n8351), .A(n8350), .ZN(n8371) );
  INV_X1 U9956 ( .A(n8353), .ZN(n8360) );
  AOI21_X1 U9957 ( .B1(n8356), .B2(n8355), .A(n8354), .ZN(n8358) );
  OR2_X1 U9958 ( .A1(n8358), .A2(n8357), .ZN(n8359) );
  OAI211_X1 U9959 ( .C1(n10021), .C2(n8361), .A(n8360), .B(n8359), .ZN(n8367)
         );
  AOI21_X1 U9960 ( .B1(n8364), .B2(n8363), .A(n8362), .ZN(n8365) );
  NOR2_X1 U9961 ( .A1(n8365), .A2(n9999), .ZN(n8366) );
  AOI211_X1 U9962 ( .C1(n8369), .C2(n8368), .A(n8367), .B(n8366), .ZN(n8370)
         );
  OAI21_X1 U9963 ( .B1(n8371), .B2(n10014), .A(n8370), .ZN(P2_U3197) );
  NOR2_X1 U9964 ( .A1(n8373), .A2(n8372), .ZN(n8587) );
  NOR2_X1 U9965 ( .A1(n9703), .A2(n8374), .ZN(n8383) );
  AOI21_X1 U9966 ( .B1(n9716), .B2(n8587), .A(n8383), .ZN(n8378) );
  NAND2_X1 U9967 ( .A1(n9719), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8375) );
  OAI211_X1 U9968 ( .C1(n8376), .C2(n8523), .A(n8378), .B(n8375), .ZN(P2_U3202) );
  INV_X1 U9969 ( .A(n8591), .ZN(n8379) );
  NAND2_X1 U9970 ( .A1(n9719), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8377) );
  OAI211_X1 U9971 ( .C1(n8379), .C2(n8523), .A(n8378), .B(n8377), .ZN(P2_U3203) );
  NAND2_X1 U9972 ( .A1(n8380), .A2(n9716), .ZN(n8385) );
  NOR2_X1 U9973 ( .A1(n8381), .A2(n8523), .ZN(n8382) );
  AOI211_X1 U9974 ( .C1(n9719), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8383), .B(
        n8382), .ZN(n8384) );
  OAI211_X1 U9975 ( .C1(n8387), .C2(n8386), .A(n8385), .B(n8384), .ZN(P2_U3204) );
  XNOR2_X1 U9976 ( .A(n8388), .B(n8395), .ZN(n8394) );
  AND2_X1 U9977 ( .A1(n8391), .A2(n8512), .ZN(n8392) );
  XNOR2_X1 U9978 ( .A(n8396), .B(n8395), .ZN(n8534) );
  AOI22_X1 U9979 ( .A1(n9719), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8521), .B2(
        n8397), .ZN(n8398) );
  OAI21_X1 U9980 ( .B1(n8399), .B2(n8523), .A(n8398), .ZN(n8400) );
  AOI21_X1 U9981 ( .B1(n8534), .B2(n8525), .A(n8400), .ZN(n8401) );
  OAI21_X1 U9982 ( .B1(n8536), .B2(n9719), .A(n8401), .ZN(P2_U3205) );
  INV_X1 U9983 ( .A(n8410), .ZN(n8402) );
  XNOR2_X1 U9984 ( .A(n8403), .B(n8402), .ZN(n8408) );
  OAI21_X1 U9985 ( .B1(n8411), .B2(n8410), .A(n8409), .ZN(n8540) );
  INV_X1 U9986 ( .A(n8540), .ZN(n8416) );
  AOI22_X1 U9987 ( .A1(n9719), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8521), .B2(
        n8412), .ZN(n8413) );
  OAI21_X1 U9988 ( .B1(n8414), .B2(n8523), .A(n8413), .ZN(n8415) );
  AOI21_X1 U9989 ( .B1(n8416), .B2(n8525), .A(n8415), .ZN(n8417) );
  OAI21_X1 U9990 ( .B1(n8539), .B2(n9719), .A(n8417), .ZN(P2_U3206) );
  XOR2_X1 U9991 ( .A(n8428), .B(n8418), .Z(n8419) );
  OAI222_X1 U9992 ( .A1(n9712), .A2(n8420), .B1(n9710), .B2(n8455), .C1(n8419), 
        .C2(n10024), .ZN(n8541) );
  INV_X1 U9993 ( .A(n8541), .ZN(n8434) );
  INV_X1 U9994 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8423) );
  INV_X1 U9995 ( .A(n8421), .ZN(n8422) );
  OAI22_X1 U9996 ( .A1(n9716), .A2(n8423), .B1(n8422), .B2(n9703), .ZN(n8424)
         );
  AOI21_X1 U9997 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8433) );
  NAND2_X1 U9998 ( .A1(n8448), .A2(n8447), .ZN(n8545) );
  NAND2_X1 U9999 ( .A1(n8545), .A2(n8427), .ZN(n8429) );
  NAND2_X1 U10000 ( .A1(n8429), .A2(n8428), .ZN(n8431) );
  OR2_X1 U10001 ( .A1(n8429), .A2(n8428), .ZN(n8430) );
  NAND2_X1 U10002 ( .A1(n8542), .A2(n8525), .ZN(n8432) );
  OAI211_X1 U10003 ( .C1(n8434), .C2(n9719), .A(n8433), .B(n8432), .ZN(
        P2_U3207) );
  INV_X1 U10004 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8451) );
  OAI211_X1 U10005 ( .C1(n8437), .C2(n8436), .A(n8435), .B(n8510), .ZN(n8441)
         );
  OAI22_X1 U10006 ( .A1(n8464), .A2(n9710), .B1(n8438), .B2(n9712), .ZN(n8439)
         );
  INV_X1 U10007 ( .A(n8439), .ZN(n8440) );
  NAND2_X1 U10008 ( .A1(n8441), .A2(n8440), .ZN(n8550) );
  NAND2_X1 U10009 ( .A1(n8442), .A2(n10028), .ZN(n8547) );
  INV_X1 U10010 ( .A(n8443), .ZN(n8444) );
  OAI22_X1 U10011 ( .A1(n8547), .A2(n8445), .B1(n8444), .B2(n9703), .ZN(n8446)
         );
  OAI21_X1 U10012 ( .B1(n8550), .B2(n8446), .A(n9716), .ZN(n8450) );
  OR2_X1 U10013 ( .A1(n8448), .A2(n8447), .ZN(n8546) );
  NAND3_X1 U10014 ( .A1(n8546), .A2(n8545), .A3(n8525), .ZN(n8449) );
  OAI211_X1 U10015 ( .C1(n9716), .C2(n8451), .A(n8450), .B(n8449), .ZN(
        P2_U3208) );
  NOR2_X1 U10016 ( .A1(n8748), .A2(n9705), .ZN(n8456) );
  OAI211_X1 U10017 ( .C1(n4318), .C2(n4722), .A(n8510), .B(n8452), .ZN(n8454)
         );
  NAND2_X1 U10018 ( .A1(n8475), .A2(n8512), .ZN(n8453) );
  OAI211_X1 U10019 ( .C1(n8455), .C2(n9712), .A(n8454), .B(n8453), .ZN(n8551)
         );
  AOI211_X1 U10020 ( .C1(n8521), .C2(n8457), .A(n8456), .B(n8551), .ZN(n8461)
         );
  XNOR2_X1 U10021 ( .A(n8459), .B(n8458), .ZN(n8552) );
  AOI22_X1 U10022 ( .A1(n8552), .A2(n8525), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9719), .ZN(n8460) );
  OAI21_X1 U10023 ( .B1(n8461), .B2(n9719), .A(n8460), .ZN(P2_U3209) );
  XNOR2_X1 U10024 ( .A(n8462), .B(n8466), .ZN(n8463) );
  OAI222_X1 U10025 ( .A1(n9712), .A2(n8464), .B1(n9710), .B2(n8489), .C1(
        n10024), .C2(n8463), .ZN(n8555) );
  INV_X1 U10026 ( .A(n8555), .ZN(n8471) );
  XOR2_X1 U10027 ( .A(n8466), .B(n8465), .Z(n8556) );
  AOI22_X1 U10028 ( .A1(n8521), .A2(n8467), .B1(n9719), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n8468) );
  OAI21_X1 U10029 ( .B1(n8752), .B2(n8523), .A(n8468), .ZN(n8469) );
  AOI21_X1 U10030 ( .B1(n8556), .B2(n8525), .A(n8469), .ZN(n8470) );
  OAI21_X1 U10031 ( .B1(n8471), .B2(n9719), .A(n8470), .ZN(P2_U3210) );
  OAI21_X1 U10032 ( .B1(n8474), .B2(n8473), .A(n8472), .ZN(n8476) );
  AOI222_X1 U10033 ( .A1(n8510), .A2(n8476), .B1(n8475), .B2(n8513), .C1(n8501), .C2(n8512), .ZN(n8477) );
  INV_X1 U10034 ( .A(n8477), .ZN(n8559) );
  NOR2_X1 U10035 ( .A1(n8479), .A2(n8478), .ZN(n8558) );
  INV_X1 U10036 ( .A(n8558), .ZN(n8480) );
  NAND3_X1 U10037 ( .A1(n8480), .A2(n8525), .A3(n8560), .ZN(n8483) );
  AOI22_X1 U10038 ( .A1(n9719), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8521), .B2(
        n8481), .ZN(n8482) );
  OAI211_X1 U10039 ( .C1(n8756), .C2(n8523), .A(n8483), .B(n8482), .ZN(n8484)
         );
  AOI21_X1 U10040 ( .B1(n8559), .B2(n9716), .A(n8484), .ZN(n8485) );
  INV_X1 U10041 ( .A(n8485), .ZN(P2_U3211) );
  XNOR2_X1 U10042 ( .A(n8486), .B(n8491), .ZN(n8487) );
  OAI222_X1 U10043 ( .A1(n9712), .A2(n8489), .B1(n9710), .B2(n8488), .C1(
        n10024), .C2(n8487), .ZN(n8563) );
  INV_X1 U10044 ( .A(n8563), .ZN(n8496) );
  XNOR2_X1 U10045 ( .A(n8490), .B(n8491), .ZN(n8564) );
  AOI22_X1 U10046 ( .A1(n9719), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8521), .B2(
        n8492), .ZN(n8493) );
  OAI21_X1 U10047 ( .B1(n8760), .B2(n8523), .A(n8493), .ZN(n8494) );
  AOI21_X1 U10048 ( .B1(n8564), .B2(n8525), .A(n8494), .ZN(n8495) );
  OAI21_X1 U10049 ( .B1(n8496), .B2(n9719), .A(n8495), .ZN(P2_U3212) );
  OAI21_X1 U10050 ( .B1(n8499), .B2(n8498), .A(n8497), .ZN(n8502) );
  AOI222_X1 U10051 ( .A1(n8510), .A2(n8502), .B1(n8501), .B2(n8513), .C1(n8500), .C2(n8512), .ZN(n8567) );
  XNOR2_X1 U10052 ( .A(n8503), .B(n8504), .ZN(n8569) );
  AOI22_X1 U10053 ( .A1(n9719), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8521), .B2(
        n8505), .ZN(n8506) );
  OAI21_X1 U10054 ( .B1(n8764), .B2(n8523), .A(n8506), .ZN(n8507) );
  AOI21_X1 U10055 ( .B1(n8569), .B2(n8525), .A(n8507), .ZN(n8508) );
  OAI21_X1 U10056 ( .B1(n8567), .B2(n9719), .A(n8508), .ZN(P2_U3213) );
  OAI211_X1 U10057 ( .C1(n4300), .C2(n6348), .A(n8510), .B(n8509), .ZN(n8516)
         );
  AOI22_X1 U10058 ( .A1(n8514), .A2(n8513), .B1(n8512), .B2(n8511), .ZN(n8515)
         );
  NAND2_X1 U10059 ( .A1(n8516), .A2(n8515), .ZN(n8572) );
  INV_X1 U10060 ( .A(n8572), .ZN(n8527) );
  NAND2_X1 U10061 ( .A1(n8578), .A2(n8517), .ZN(n8518) );
  XOR2_X1 U10062 ( .A(n8519), .B(n8518), .Z(n8573) );
  AOI22_X1 U10063 ( .A1(n9719), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8521), .B2(
        n8520), .ZN(n8522) );
  OAI21_X1 U10064 ( .B1(n8769), .B2(n8523), .A(n8522), .ZN(n8524) );
  AOI21_X1 U10065 ( .B1(n8573), .B2(n8525), .A(n8524), .ZN(n8526) );
  OAI21_X1 U10066 ( .B1(n8527), .B2(n9719), .A(n8526), .ZN(P2_U3214) );
  INV_X1 U10067 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8529) );
  INV_X1 U10068 ( .A(n8576), .ZN(n8530) );
  NAND2_X1 U10069 ( .A1(n8586), .A2(n8530), .ZN(n8528) );
  NAND2_X1 U10070 ( .A1(n8587), .A2(n10121), .ZN(n8531) );
  OAI211_X1 U10071 ( .C1(n10121), .C2(n8529), .A(n8528), .B(n8531), .ZN(
        P2_U3490) );
  INV_X1 U10072 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8628) );
  NAND2_X1 U10073 ( .A1(n8591), .A2(n8530), .ZN(n8532) );
  OAI211_X1 U10074 ( .C1(n10121), .C2(n8628), .A(n8532), .B(n8531), .ZN(
        P2_U3489) );
  AOI22_X1 U10075 ( .A1(n8534), .A2(n10084), .B1(n10028), .B2(n8533), .ZN(
        n8535) );
  NAND2_X1 U10076 ( .A1(n8536), .A2(n8535), .ZN(n8595) );
  MUX2_X1 U10077 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8595), .S(n10121), .Z(
        P2_U3487) );
  NAND2_X1 U10078 ( .A1(n8537), .A2(n10028), .ZN(n8538) );
  OAI211_X1 U10079 ( .C1(n10088), .C2(n8540), .A(n8539), .B(n8538), .ZN(n8596)
         );
  MUX2_X1 U10080 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8596), .S(n10121), .Z(
        P2_U3486) );
  INV_X1 U10081 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8543) );
  AOI21_X1 U10082 ( .B1(n8542), .B2(n10084), .A(n8541), .ZN(n8740) );
  MUX2_X1 U10083 ( .A(n8543), .B(n8740), .S(n10121), .Z(n8544) );
  OAI21_X1 U10084 ( .B1(n8743), .B2(n8576), .A(n8544), .ZN(P2_U3485) );
  NAND3_X1 U10085 ( .A1(n8546), .A2(n8545), .A3(n10084), .ZN(n8548) );
  NAND2_X1 U10086 ( .A1(n8548), .A2(n8547), .ZN(n8549) );
  MUX2_X1 U10087 ( .A(n8744), .B(P2_REG1_REG_25__SCAN_IN), .S(n10119), .Z(
        P2_U3484) );
  AOI21_X1 U10088 ( .B1(n8552), .B2(n10084), .A(n8551), .ZN(n8745) );
  MUX2_X1 U10089 ( .A(n8553), .B(n8745), .S(n10121), .Z(n8554) );
  OAI21_X1 U10090 ( .B1(n8748), .B2(n8576), .A(n8554), .ZN(P2_U3483) );
  AOI21_X1 U10091 ( .B1(n10084), .B2(n8556), .A(n8555), .ZN(n8749) );
  MUX2_X1 U10092 ( .A(n8685), .B(n8749), .S(n10121), .Z(n8557) );
  OAI21_X1 U10093 ( .B1(n8752), .B2(n8576), .A(n8557), .ZN(P2_U3482) );
  NOR2_X1 U10094 ( .A1(n8558), .A2(n10088), .ZN(n8561) );
  AOI21_X1 U10095 ( .B1(n8561), .B2(n8560), .A(n8559), .ZN(n8753) );
  MUX2_X1 U10096 ( .A(n8630), .B(n8753), .S(n10121), .Z(n8562) );
  OAI21_X1 U10097 ( .B1(n8756), .B2(n8576), .A(n8562), .ZN(P2_U3481) );
  INV_X1 U10098 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8565) );
  AOI21_X1 U10099 ( .B1(n8564), .B2(n10084), .A(n8563), .ZN(n8757) );
  MUX2_X1 U10100 ( .A(n8565), .B(n8757), .S(n10121), .Z(n8566) );
  OAI21_X1 U10101 ( .B1(n8760), .B2(n8576), .A(n8566), .ZN(P2_U3480) );
  INV_X1 U10102 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8570) );
  INV_X1 U10103 ( .A(n8567), .ZN(n8568) );
  AOI21_X1 U10104 ( .B1(n8569), .B2(n10084), .A(n8568), .ZN(n8761) );
  MUX2_X1 U10105 ( .A(n8570), .B(n8761), .S(n10121), .Z(n8571) );
  OAI21_X1 U10106 ( .B1(n8764), .B2(n8576), .A(n8571), .ZN(P2_U3479) );
  INV_X1 U10107 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8574) );
  AOI21_X1 U10108 ( .B1(n10084), .B2(n8573), .A(n8572), .ZN(n8765) );
  MUX2_X1 U10109 ( .A(n8574), .B(n8765), .S(n10121), .Z(n8575) );
  OAI21_X1 U10110 ( .B1(n8769), .B2(n8576), .A(n8575), .ZN(P2_U3478) );
  NAND3_X1 U10111 ( .A1(n8578), .A2(n10084), .A3(n8577), .ZN(n8579) );
  NAND3_X1 U10112 ( .A1(n8581), .A2(n8580), .A3(n8579), .ZN(n8770) );
  MUX2_X1 U10113 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8770), .S(n10121), .Z(
        P2_U3477) );
  AOI22_X1 U10114 ( .A1(n8583), .A2(n10084), .B1(n10028), .B2(n8582), .ZN(
        n8584) );
  NAND2_X1 U10115 ( .A1(n8585), .A2(n8584), .ZN(n8771) );
  MUX2_X1 U10116 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8771), .S(n10121), .Z(
        P2_U3476) );
  INV_X1 U10117 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8589) );
  INV_X1 U10118 ( .A(n8768), .ZN(n8590) );
  NAND2_X1 U10119 ( .A1(n8586), .A2(n8590), .ZN(n8588) );
  NAND2_X1 U10120 ( .A1(n10094), .A2(n8587), .ZN(n8592) );
  OAI211_X1 U10121 ( .C1(n8589), .C2(n10094), .A(n8588), .B(n8592), .ZN(
        P2_U3458) );
  INV_X1 U10122 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8594) );
  NAND2_X1 U10123 ( .A1(n8591), .A2(n8590), .ZN(n8593) );
  OAI211_X1 U10124 ( .C1(n8594), .C2(n10094), .A(n8593), .B(n8592), .ZN(
        P2_U3457) );
  MUX2_X1 U10125 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8595), .S(n10094), .Z(
        P2_U3455) );
  MUX2_X1 U10126 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8596), .S(n10094), .Z(
        n8739) );
  NAND3_X1 U10127 ( .A1(keyinput51), .A2(keyinput21), .A3(keyinput10), .ZN(
        n8610) );
  NAND2_X1 U10128 ( .A1(keyinput41), .A2(keyinput63), .ZN(n8597) );
  NOR3_X1 U10129 ( .A1(keyinput33), .A2(keyinput6), .A3(n8597), .ZN(n8601) );
  NAND2_X1 U10130 ( .A1(keyinput7), .A2(keyinput31), .ZN(n8598) );
  NOR3_X1 U10131 ( .A1(keyinput3), .A2(keyinput61), .A3(n8598), .ZN(n8600) );
  NOR3_X1 U10132 ( .A1(keyinput62), .A2(keyinput16), .A3(keyinput13), .ZN(
        n8599) );
  NAND4_X1 U10133 ( .A1(n8601), .A2(n8600), .A3(keyinput12), .A4(n8599), .ZN(
        n8609) );
  NOR3_X1 U10134 ( .A1(keyinput0), .A2(keyinput5), .A3(keyinput53), .ZN(n8607)
         );
  NAND2_X1 U10135 ( .A1(keyinput58), .A2(keyinput1), .ZN(n8602) );
  NOR3_X1 U10136 ( .A1(keyinput20), .A2(keyinput54), .A3(n8602), .ZN(n8606) );
  NAND3_X1 U10137 ( .A1(keyinput44), .A2(keyinput35), .A3(keyinput56), .ZN(
        n8604) );
  NAND3_X1 U10138 ( .A1(keyinput50), .A2(keyinput9), .A3(keyinput24), .ZN(
        n8603) );
  NOR4_X1 U10139 ( .A1(keyinput19), .A2(keyinput28), .A3(n8604), .A4(n8603), 
        .ZN(n8605) );
  NAND4_X1 U10140 ( .A1(keyinput27), .A2(n8607), .A3(n8606), .A4(n8605), .ZN(
        n8608) );
  NOR4_X1 U10141 ( .A1(keyinput15), .A2(n8610), .A3(n8609), .A4(n8608), .ZN(
        n8625) );
  NOR2_X1 U10142 ( .A1(keyinput60), .A2(keyinput32), .ZN(n8615) );
  NOR4_X1 U10143 ( .A1(keyinput8), .A2(keyinput37), .A3(keyinput29), .A4(
        keyinput55), .ZN(n8612) );
  NOR2_X1 U10144 ( .A1(keyinput23), .A2(keyinput52), .ZN(n8611) );
  NAND4_X1 U10145 ( .A1(n8612), .A2(keyinput49), .A3(keyinput45), .A4(n8611), 
        .ZN(n8613) );
  NOR4_X1 U10146 ( .A1(keyinput42), .A2(keyinput4), .A3(keyinput17), .A4(n8613), .ZN(n8614) );
  NAND4_X1 U10147 ( .A1(keyinput48), .A2(keyinput43), .A3(n8615), .A4(n8614), 
        .ZN(n8623) );
  NAND3_X1 U10148 ( .A1(keyinput38), .A2(keyinput18), .A3(keyinput59), .ZN(
        n8622) );
  NOR2_X1 U10149 ( .A1(keyinput39), .A2(keyinput34), .ZN(n8620) );
  NAND2_X1 U10150 ( .A1(keyinput36), .A2(keyinput26), .ZN(n8618) );
  NOR2_X1 U10151 ( .A1(keyinput30), .A2(keyinput22), .ZN(n8616) );
  NAND3_X1 U10152 ( .A1(keyinput25), .A2(keyinput2), .A3(n8616), .ZN(n8617) );
  NOR4_X1 U10153 ( .A1(keyinput57), .A2(keyinput47), .A3(n8618), .A4(n8617), 
        .ZN(n8619) );
  NAND4_X1 U10154 ( .A1(keyinput40), .A2(keyinput46), .A3(n8620), .A4(n8619), 
        .ZN(n8621) );
  NOR4_X1 U10155 ( .A1(keyinput14), .A2(n8623), .A3(n8622), .A4(n8621), .ZN(
        n8624) );
  AOI21_X1 U10156 ( .B1(n8625), .B2(n8624), .A(keyinput11), .ZN(n8737) );
  INV_X1 U10157 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8627) );
  OAI22_X1 U10158 ( .A1(n8628), .A2(keyinput24), .B1(n8627), .B2(keyinput20), 
        .ZN(n8626) );
  AOI221_X1 U10159 ( .B1(n8628), .B2(keyinput24), .C1(keyinput20), .C2(n8627), 
        .A(n8626), .ZN(n8633) );
  OAI22_X1 U10160 ( .A1(n8631), .A2(keyinput28), .B1(n8630), .B2(keyinput9), 
        .ZN(n8629) );
  AOI221_X1 U10161 ( .B1(n8631), .B2(keyinput28), .C1(keyinput9), .C2(n8630), 
        .A(n8629), .ZN(n8632) );
  AND2_X1 U10162 ( .A1(n8633), .A2(n8632), .ZN(n8642) );
  OAI22_X1 U10163 ( .A1(n9590), .A2(keyinput17), .B1(n4703), .B2(keyinput1), 
        .ZN(n8634) );
  AOI221_X1 U10164 ( .B1(n9590), .B2(keyinput17), .C1(keyinput1), .C2(n4703), 
        .A(n8634), .ZN(n8641) );
  INV_X1 U10165 ( .A(keyinput5), .ZN(n8636) );
  OAI22_X1 U10166 ( .A1(n6485), .A2(keyinput27), .B1(n8636), .B2(
        P2_REG3_REG_6__SCAN_IN), .ZN(n8635) );
  AOI221_X1 U10167 ( .B1(n6485), .B2(keyinput27), .C1(P2_REG3_REG_6__SCAN_IN), 
        .C2(n8636), .A(n8635), .ZN(n8640) );
  OAI22_X1 U10168 ( .A1(n8638), .A2(keyinput19), .B1(n10107), .B2(keyinput35), 
        .ZN(n8637) );
  AOI221_X1 U10169 ( .B1(n8638), .B2(keyinput19), .C1(keyinput35), .C2(n10107), 
        .A(n8637), .ZN(n8639) );
  NAND4_X1 U10170 ( .A1(n8642), .A2(n8641), .A3(n8640), .A4(n8639), .ZN(n8735)
         );
  INV_X1 U10171 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9903) );
  INV_X1 U10172 ( .A(keyinput44), .ZN(n8644) );
  OAI22_X1 U10173 ( .A1(n9903), .A2(keyinput53), .B1(n8644), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n8643) );
  AOI221_X1 U10174 ( .B1(n9903), .B2(keyinput53), .C1(P2_ADDR_REG_14__SCAN_IN), 
        .C2(n8644), .A(n8643), .ZN(n8648) );
  INV_X1 U10175 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n9902) );
  INV_X1 U10176 ( .A(keyinput56), .ZN(n8646) );
  OAI22_X1 U10177 ( .A1(n9902), .A2(keyinput50), .B1(n8646), .B2(
        P2_IR_REG_5__SCAN_IN), .ZN(n8645) );
  AOI221_X1 U10178 ( .B1(n9902), .B2(keyinput50), .C1(P2_IR_REG_5__SCAN_IN), 
        .C2(n8646), .A(n8645), .ZN(n8647) );
  NAND2_X1 U10179 ( .A1(n8648), .A2(n8647), .ZN(n8734) );
  INV_X1 U10180 ( .A(keyinput62), .ZN(n8650) );
  AOI22_X1 U10181 ( .A1(n8651), .A2(keyinput61), .B1(P2_REG2_REG_31__SCAN_IN), 
        .B2(n8650), .ZN(n8649) );
  OAI221_X1 U10182 ( .B1(n8651), .B2(keyinput61), .C1(n8650), .C2(
        P2_REG2_REG_31__SCAN_IN), .A(n8649), .ZN(n8656) );
  INV_X1 U10183 ( .A(SI_18_), .ZN(n8654) );
  INV_X1 U10184 ( .A(keyinput47), .ZN(n8653) );
  AOI22_X1 U10185 ( .A1(n8654), .A2(keyinput30), .B1(P1_ADDR_REG_10__SCAN_IN), 
        .B2(n8653), .ZN(n8652) );
  OAI221_X1 U10186 ( .B1(n8654), .B2(keyinput30), .C1(n8653), .C2(
        P1_ADDR_REG_10__SCAN_IN), .A(n8652), .ZN(n8655) );
  NOR2_X1 U10187 ( .A1(n8656), .A2(n8655), .ZN(n8678) );
  INV_X1 U10188 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n9901) );
  INV_X1 U10189 ( .A(keyinput59), .ZN(n8658) );
  AOI22_X1 U10190 ( .A1(n9901), .A2(keyinput18), .B1(P2_WR_REG_SCAN_IN), .B2(
        n8658), .ZN(n8657) );
  OAI221_X1 U10191 ( .B1(n9901), .B2(keyinput18), .C1(n8658), .C2(
        P2_WR_REG_SCAN_IN), .A(n8657), .ZN(n8663) );
  INV_X1 U10192 ( .A(keyinput52), .ZN(n8661) );
  INV_X1 U10193 ( .A(keyinput38), .ZN(n8660) );
  AOI22_X1 U10194 ( .A1(n8661), .A2(P2_ADDR_REG_6__SCAN_IN), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8660), .ZN(n8659) );
  OAI221_X1 U10195 ( .B1(n8661), .B2(P2_ADDR_REG_6__SCAN_IN), .C1(n8660), .C2(
        P1_ADDR_REG_15__SCAN_IN), .A(n8659), .ZN(n8662) );
  NOR2_X1 U10196 ( .A1(n8663), .A2(n8662), .ZN(n8677) );
  AOI22_X1 U10197 ( .A1(n8846), .A2(keyinput4), .B1(keyinput48), .B2(n6108), 
        .ZN(n8664) );
  OAI221_X1 U10198 ( .B1(n8846), .B2(keyinput4), .C1(n6108), .C2(keyinput48), 
        .A(n8664), .ZN(n8668) );
  INV_X1 U10199 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n9904) );
  INV_X1 U10200 ( .A(keyinput37), .ZN(n8666) );
  AOI22_X1 U10201 ( .A1(n9904), .A2(keyinput29), .B1(P1_ADDR_REG_13__SCAN_IN), 
        .B2(n8666), .ZN(n8665) );
  OAI221_X1 U10202 ( .B1(n9904), .B2(keyinput29), .C1(n8666), .C2(
        P1_ADDR_REG_13__SCAN_IN), .A(n8665), .ZN(n8667) );
  NOR2_X1 U10203 ( .A1(n8668), .A2(n8667), .ZN(n8676) );
  INV_X1 U10204 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9905) );
  AOI22_X1 U10205 ( .A1(n5081), .A2(keyinput55), .B1(n9905), .B2(keyinput49), 
        .ZN(n8669) );
  OAI221_X1 U10206 ( .B1(n5081), .B2(keyinput55), .C1(n9905), .C2(keyinput49), 
        .A(n8669), .ZN(n8674) );
  INV_X1 U10207 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n8671) );
  AOI22_X1 U10208 ( .A1(n8672), .A2(keyinput41), .B1(n8671), .B2(keyinput7), 
        .ZN(n8670) );
  OAI221_X1 U10209 ( .B1(n8672), .B2(keyinput41), .C1(n8671), .C2(keyinput7), 
        .A(n8670), .ZN(n8673) );
  NOR2_X1 U10210 ( .A1(n8674), .A2(n8673), .ZN(n8675) );
  NAND4_X1 U10211 ( .A1(n8678), .A2(n8677), .A3(n8676), .A4(n8675), .ZN(n8733)
         );
  AOI22_X1 U10212 ( .A1(n8680), .A2(keyinput25), .B1(keyinput2), .B2(n7658), 
        .ZN(n8679) );
  OAI221_X1 U10213 ( .B1(n8680), .B2(keyinput25), .C1(n7658), .C2(keyinput2), 
        .A(n8679), .ZN(n8688) );
  INV_X1 U10214 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8758) );
  AOI22_X1 U10215 ( .A1(n8682), .A2(keyinput60), .B1(keyinput43), .B2(n8758), 
        .ZN(n8681) );
  OAI221_X1 U10216 ( .B1(n8682), .B2(keyinput60), .C1(n8758), .C2(keyinput43), 
        .A(n8681), .ZN(n8687) );
  AOI22_X1 U10217 ( .A1(n8685), .A2(keyinput13), .B1(n8684), .B2(keyinput0), 
        .ZN(n8683) );
  OAI221_X1 U10218 ( .B1(n8685), .B2(keyinput13), .C1(n8684), .C2(keyinput0), 
        .A(n8683), .ZN(n8686) );
  OR3_X1 U10219 ( .A1(n8688), .A2(n8687), .A3(n8686), .ZN(n8731) );
  AOI22_X1 U10220 ( .A1(n8690), .A2(keyinput6), .B1(keyinput33), .B2(n6140), 
        .ZN(n8689) );
  OAI221_X1 U10221 ( .B1(n8690), .B2(keyinput6), .C1(n6140), .C2(keyinput33), 
        .A(n8689), .ZN(n8730) );
  AOI22_X1 U10222 ( .A1(n8693), .A2(keyinput39), .B1(keyinput34), .B2(n8692), 
        .ZN(n8691) );
  OAI221_X1 U10223 ( .B1(n8693), .B2(keyinput39), .C1(n8692), .C2(keyinput34), 
        .A(n8691), .ZN(n8729) );
  AOI22_X1 U10224 ( .A1(n9260), .A2(keyinput21), .B1(n8695), .B2(keyinput15), 
        .ZN(n8694) );
  OAI221_X1 U10225 ( .B1(n9260), .B2(keyinput21), .C1(n8695), .C2(keyinput15), 
        .A(n8694), .ZN(n8698) );
  AOI22_X1 U10226 ( .A1(n5097), .A2(keyinput46), .B1(keyinput36), .B2(n9985), 
        .ZN(n8696) );
  OAI221_X1 U10227 ( .B1(n5097), .B2(keyinput46), .C1(n9985), .C2(keyinput36), 
        .A(n8696), .ZN(n8697) );
  NOR2_X1 U10228 ( .A1(n8698), .A2(n8697), .ZN(n8727) );
  INV_X1 U10229 ( .A(keyinput57), .ZN(n8699) );
  XNOR2_X1 U10230 ( .A(n8699), .B(P1_REG2_REG_31__SCAN_IN), .ZN(n8703) );
  INV_X1 U10231 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10080) );
  XNOR2_X1 U10232 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput42), .ZN(n8701) );
  XNOR2_X1 U10233 ( .A(keyinput10), .B(P1_REG2_REG_28__SCAN_IN), .ZN(n8700) );
  OAI211_X1 U10234 ( .C1(keyinput11), .C2(n10080), .A(n8701), .B(n8700), .ZN(
        n8702) );
  NOR2_X1 U10235 ( .A1(n8703), .A2(n8702), .ZN(n8726) );
  XNOR2_X1 U10236 ( .A(P2_IR_REG_31__SCAN_IN), .B(keyinput63), .ZN(n8707) );
  XNOR2_X1 U10237 ( .A(SI_0_), .B(keyinput12), .ZN(n8706) );
  XNOR2_X1 U10238 ( .A(P2_REG1_REG_24__SCAN_IN), .B(keyinput3), .ZN(n8705) );
  XNOR2_X1 U10239 ( .A(P2_REG3_REG_21__SCAN_IN), .B(keyinput58), .ZN(n8704) );
  NAND4_X1 U10240 ( .A1(n8707), .A2(n8706), .A3(n8705), .A4(n8704), .ZN(n8713)
         );
  XNOR2_X1 U10241 ( .A(P2_REG2_REG_2__SCAN_IN), .B(keyinput31), .ZN(n8711) );
  XNOR2_X1 U10242 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput32), .ZN(n8710) );
  XNOR2_X1 U10243 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput54), .ZN(n8709) );
  XNOR2_X1 U10244 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput45), .ZN(n8708) );
  NAND4_X1 U10245 ( .A1(n8711), .A2(n8710), .A3(n8709), .A4(n8708), .ZN(n8712)
         );
  NOR2_X1 U10246 ( .A1(n8713), .A2(n8712), .ZN(n8725) );
  XNOR2_X1 U10247 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput40), .ZN(n8717) );
  XNOR2_X1 U10248 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(keyinput23), .ZN(n8716)
         );
  XNOR2_X1 U10249 ( .A(P2_IR_REG_13__SCAN_IN), .B(keyinput26), .ZN(n8715) );
  XNOR2_X1 U10250 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput22), .ZN(n8714) );
  NAND4_X1 U10251 ( .A1(n8717), .A2(n8716), .A3(n8715), .A4(n8714), .ZN(n8723)
         );
  XNOR2_X1 U10252 ( .A(keyinput8), .B(P1_IR_REG_29__SCAN_IN), .ZN(n8721) );
  XNOR2_X1 U10253 ( .A(SI_22_), .B(keyinput51), .ZN(n8720) );
  XNOR2_X1 U10254 ( .A(keyinput14), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n8719) );
  XNOR2_X1 U10255 ( .A(keyinput16), .B(P1_REG2_REG_29__SCAN_IN), .ZN(n8718) );
  NAND4_X1 U10256 ( .A1(n8721), .A2(n8720), .A3(n8719), .A4(n8718), .ZN(n8722)
         );
  NOR2_X1 U10257 ( .A1(n8723), .A2(n8722), .ZN(n8724) );
  NAND4_X1 U10258 ( .A1(n8727), .A2(n8726), .A3(n8725), .A4(n8724), .ZN(n8728)
         );
  OR4_X1 U10259 ( .A1(n8731), .A2(n8730), .A3(n8729), .A4(n8728), .ZN(n8732)
         );
  NOR4_X1 U10260 ( .A1(n8735), .A2(n8734), .A3(n8733), .A4(n8732), .ZN(n8736)
         );
  OAI21_X1 U10261 ( .B1(n8737), .B2(P2_REG0_REG_10__SCAN_IN), .A(n8736), .ZN(
        n8738) );
  XNOR2_X1 U10262 ( .A(n8739), .B(n8738), .ZN(P2_U3454) );
  INV_X1 U10263 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8741) );
  MUX2_X1 U10264 ( .A(n8741), .B(n8740), .S(n10094), .Z(n8742) );
  OAI21_X1 U10265 ( .B1(n8743), .B2(n8768), .A(n8742), .ZN(P2_U3453) );
  MUX2_X1 U10266 ( .A(n8744), .B(P2_REG0_REG_25__SCAN_IN), .S(n10092), .Z(
        P2_U3452) );
  INV_X1 U10267 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8746) );
  MUX2_X1 U10268 ( .A(n8746), .B(n8745), .S(n10094), .Z(n8747) );
  OAI21_X1 U10269 ( .B1(n8748), .B2(n8768), .A(n8747), .ZN(P2_U3451) );
  INV_X1 U10270 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8750) );
  MUX2_X1 U10271 ( .A(n8750), .B(n8749), .S(n10094), .Z(n8751) );
  OAI21_X1 U10272 ( .B1(n8752), .B2(n8768), .A(n8751), .ZN(P2_U3450) );
  INV_X1 U10273 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8754) );
  MUX2_X1 U10274 ( .A(n8754), .B(n8753), .S(n10094), .Z(n8755) );
  OAI21_X1 U10275 ( .B1(n8756), .B2(n8768), .A(n8755), .ZN(P2_U3449) );
  MUX2_X1 U10276 ( .A(n8758), .B(n8757), .S(n10094), .Z(n8759) );
  OAI21_X1 U10277 ( .B1(n8760), .B2(n8768), .A(n8759), .ZN(P2_U3448) );
  INV_X1 U10278 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8762) );
  MUX2_X1 U10279 ( .A(n8762), .B(n8761), .S(n10094), .Z(n8763) );
  OAI21_X1 U10280 ( .B1(n8764), .B2(n8768), .A(n8763), .ZN(P2_U3447) );
  INV_X1 U10281 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8766) );
  MUX2_X1 U10282 ( .A(n8766), .B(n8765), .S(n10094), .Z(n8767) );
  OAI21_X1 U10283 ( .B1(n8769), .B2(n8768), .A(n8767), .ZN(P2_U3446) );
  MUX2_X1 U10284 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8770), .S(n10094), .Z(
        P2_U3444) );
  MUX2_X1 U10285 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8771), .S(n10094), .Z(
        P2_U3441) );
  INV_X1 U10286 ( .A(n8772), .ZN(n9655) );
  NOR4_X1 U10287 ( .A1(n8773), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n6109), .ZN(n8774) );
  AOI21_X1 U10288 ( .B1(n8775), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8774), .ZN(
        n8776) );
  OAI21_X1 U10289 ( .B1(n9655), .B2(n8777), .A(n8776), .ZN(P2_U3264) );
  MUX2_X1 U10290 ( .A(n8778), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10291 ( .A1(n8781), .A2(n8780), .ZN(n8782) );
  XNOR2_X1 U10292 ( .A(n8779), .B(n8782), .ZN(n8789) );
  OAI22_X1 U10293 ( .A1(n8784), .A2(n8877), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8783), .ZN(n8787) );
  INV_X1 U10294 ( .A(n9424), .ZN(n8785) );
  OAI22_X1 U10295 ( .A1(n9466), .A2(n8876), .B1(n8785), .B2(n8862), .ZN(n8786)
         );
  AOI211_X1 U10296 ( .C1(n9563), .C2(n8887), .A(n8787), .B(n8786), .ZN(n8788)
         );
  OAI21_X1 U10297 ( .B1(n8789), .B2(n5697), .A(n8788), .ZN(P1_U3216) );
  INV_X1 U10298 ( .A(n8790), .ZN(n8791) );
  NAND2_X1 U10299 ( .A1(n8791), .A2(n8794), .ZN(n8792) );
  AOI22_X1 U10300 ( .A1(n4307), .A2(n8794), .B1(n8793), .B2(n8792), .ZN(n8799)
         );
  AOI22_X1 U10301 ( .A1(n9192), .A2(n9431), .B1(n9194), .B2(n9433), .ZN(n9493)
         );
  INV_X1 U10302 ( .A(n9493), .ZN(n8795) );
  AOI22_X1 U10303 ( .A1(n8795), .A2(n8888), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n8796) );
  OAI21_X1 U10304 ( .B1(n8893), .B2(n9502), .A(n8796), .ZN(n8797) );
  AOI21_X1 U10305 ( .B1(n9500), .B2(n8887), .A(n8797), .ZN(n8798) );
  OAI21_X1 U10306 ( .B1(n8799), .B2(n5697), .A(n8798), .ZN(P1_U3219) );
  NAND2_X1 U10307 ( .A1(n8800), .A2(n8844), .ZN(n8843) );
  NAND2_X1 U10308 ( .A1(n8843), .A2(n8801), .ZN(n8802) );
  XOR2_X1 U10309 ( .A(n8803), .B(n8802), .Z(n8808) );
  OAI22_X1 U10310 ( .A1(n8876), .A2(n9468), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8804), .ZN(n8806) );
  OAI22_X1 U10311 ( .A1(n9466), .A2(n8877), .B1(n8862), .B2(n9471), .ZN(n8805)
         );
  AOI211_X1 U10312 ( .C1(n9574), .C2(n8887), .A(n8806), .B(n8805), .ZN(n8807)
         );
  OAI21_X1 U10313 ( .B1(n8808), .B2(n5697), .A(n8807), .ZN(P1_U3223) );
  NAND2_X1 U10314 ( .A1(n8809), .A2(n8837), .ZN(n8836) );
  NAND2_X1 U10315 ( .A1(n8836), .A2(n8810), .ZN(n8811) );
  OAI21_X1 U10316 ( .B1(n8812), .B2(n8811), .A(n8871), .ZN(n8817) );
  AOI22_X1 U10317 ( .A1(n9432), .A2(n8832), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n8815) );
  AOI22_X1 U10318 ( .A1(n9394), .A2(n8813), .B1(n9398), .B2(n8880), .ZN(n8814)
         );
  OAI211_X1 U10319 ( .C1(n9401), .C2(n8883), .A(n8815), .B(n8814), .ZN(n8816)
         );
  AOI21_X1 U10320 ( .B1(n8817), .B2(n8895), .A(n8816), .ZN(n8818) );
  INV_X1 U10321 ( .A(n8818), .ZN(P1_U3225) );
  XOR2_X1 U10322 ( .A(n8820), .B(n8819), .Z(n8827) );
  NOR2_X1 U10323 ( .A1(n8893), .A2(n8821), .ZN(n8824) );
  NAND2_X1 U10324 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9271) );
  OAI21_X1 U10325 ( .B1(n8822), .B2(n8866), .A(n9271), .ZN(n8823) );
  AOI211_X1 U10326 ( .C1(n8825), .C2(n8887), .A(n8824), .B(n8823), .ZN(n8826)
         );
  OAI21_X1 U10327 ( .B1(n8827), .B2(n5697), .A(n8826), .ZN(P1_U3226) );
  XOR2_X1 U10328 ( .A(n8829), .B(n8828), .Z(n8835) );
  AND2_X1 U10329 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9289) );
  OAI22_X1 U10330 ( .A1(n8877), .A2(n9036), .B1(n8862), .B2(n8830), .ZN(n8831)
         );
  AOI211_X1 U10331 ( .C1(n8832), .C2(n9196), .A(n9289), .B(n8831), .ZN(n8834)
         );
  NAND2_X1 U10332 ( .A1(n9594), .A2(n8887), .ZN(n8833) );
  OAI211_X1 U10333 ( .C1(n8835), .C2(n5697), .A(n8834), .B(n8833), .ZN(
        P1_U3228) );
  INV_X1 U10334 ( .A(n9416), .ZN(n9623) );
  OAI21_X1 U10335 ( .B1(n8837), .B2(n8809), .A(n8836), .ZN(n8838) );
  NAND2_X1 U10336 ( .A1(n8838), .A2(n8895), .ZN(n8842) );
  OAI22_X1 U10337 ( .A1(n9447), .A2(n8876), .B1(n8893), .B2(n9414), .ZN(n8840)
         );
  NOR2_X1 U10338 ( .A1(n9409), .A2(n8877), .ZN(n8839) );
  AOI211_X1 U10339 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3086), .A(n8840), 
        .B(n8839), .ZN(n8841) );
  OAI211_X1 U10340 ( .C1(n9623), .C2(n8883), .A(n8842), .B(n8841), .ZN(
        P1_U3229) );
  OAI21_X1 U10341 ( .B1(n8844), .B2(n8800), .A(n8843), .ZN(n8845) );
  NAND2_X1 U10342 ( .A1(n8845), .A2(n8895), .ZN(n8849) );
  AOI22_X1 U10343 ( .A1(n9191), .A2(n9431), .B1(n9433), .B2(n9193), .ZN(n9480)
         );
  OAI22_X1 U10344 ( .A1(n9480), .A2(n8866), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8846), .ZN(n8847) );
  AOI21_X1 U10345 ( .B1(n9485), .B2(n8880), .A(n8847), .ZN(n8848) );
  OAI211_X1 U10346 ( .C1(n6085), .C2(n8883), .A(n8849), .B(n8848), .ZN(
        P1_U3233) );
  OAI21_X1 U10347 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8853) );
  NAND2_X1 U10348 ( .A1(n8853), .A2(n8895), .ZN(n8857) );
  OAI22_X1 U10349 ( .A1(n8876), .A2(n9448), .B1(n8862), .B2(n9451), .ZN(n8855)
         );
  NOR2_X1 U10350 ( .A1(n9447), .A2(n8877), .ZN(n8854) );
  AOI211_X1 U10351 ( .C1(P1_REG3_REG_22__SCAN_IN), .C2(P1_U3086), .A(n8855), 
        .B(n8854), .ZN(n8856) );
  OAI211_X1 U10352 ( .C1(n9628), .C2(n8883), .A(n8857), .B(n8856), .ZN(
        P1_U3235) );
  XOR2_X1 U10353 ( .A(n8859), .B(n8858), .Z(n8860) );
  XNOR2_X1 U10354 ( .A(n8861), .B(n8860), .ZN(n8870) );
  NOR2_X1 U10355 ( .A1(n8862), .A2(n9521), .ZN(n8868) );
  NAND2_X1 U10356 ( .A1(n9195), .A2(n9433), .ZN(n8864) );
  NAND2_X1 U10357 ( .A1(n9193), .A2(n9431), .ZN(n8863) );
  AND2_X1 U10358 ( .A1(n8864), .A2(n8863), .ZN(n9515) );
  OAI22_X1 U10359 ( .A1(n9515), .A2(n8866), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8865), .ZN(n8867) );
  AOI211_X1 U10360 ( .C1(n9520), .C2(n8887), .A(n8868), .B(n8867), .ZN(n8869)
         );
  OAI21_X1 U10361 ( .B1(n8870), .B2(n5697), .A(n8869), .ZN(P1_U3238) );
  OAI22_X1 U10362 ( .A1(n9409), .A2(n8876), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8875), .ZN(n8879) );
  NOR2_X1 U10363 ( .A1(n9377), .A2(n8877), .ZN(n8878) );
  AOI211_X1 U10364 ( .C1(n9384), .C2(n8880), .A(n8879), .B(n8878), .ZN(n8881)
         );
  OAI211_X1 U10365 ( .C1(n9618), .C2(n8883), .A(n8882), .B(n8881), .ZN(
        P1_U3240) );
  OAI21_X1 U10366 ( .B1(n8886), .B2(n8885), .A(n8884), .ZN(n8896) );
  NAND2_X1 U10367 ( .A1(n9011), .A2(n8887), .ZN(n8891) );
  AOI22_X1 U10368 ( .A1(n8889), .A2(n8888), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n8890) );
  OAI211_X1 U10369 ( .C1(n8893), .C2(n8892), .A(n8891), .B(n8890), .ZN(n8894)
         );
  AOI21_X1 U10370 ( .B1(n8896), .B2(n8895), .A(n8894), .ZN(n8897) );
  INV_X1 U10371 ( .A(n8897), .ZN(P1_U3241) );
  AND2_X1 U10372 ( .A1(n9097), .A2(n9091), .ZN(n9160) );
  NAND2_X1 U10373 ( .A1(n9628), .A2(n9434), .ZN(n8898) );
  NAND2_X1 U10374 ( .A1(n8899), .A2(n8898), .ZN(n9058) );
  NAND2_X1 U10375 ( .A1(n9058), .A2(n9059), .ZN(n8900) );
  NAND2_X1 U10376 ( .A1(n9068), .A2(n8900), .ZN(n8901) );
  NAND2_X1 U10377 ( .A1(n8901), .A2(n9067), .ZN(n8902) );
  NAND2_X1 U10378 ( .A1(n9073), .A2(n8902), .ZN(n8907) );
  INV_X1 U10379 ( .A(n8959), .ZN(n9459) );
  NAND2_X1 U10380 ( .A1(n9459), .A2(n9057), .ZN(n9047) );
  NOR2_X1 U10381 ( .A1(n8907), .A2(n9047), .ZN(n9153) );
  AOI21_X1 U10382 ( .B1(n9153), .B2(n8903), .A(n9159), .ZN(n8911) );
  INV_X1 U10383 ( .A(n9090), .ZN(n9083) );
  INV_X1 U10384 ( .A(n9077), .ZN(n8904) );
  NOR2_X1 U10385 ( .A1(n9083), .A2(n8904), .ZN(n9157) );
  INV_X1 U10386 ( .A(n9157), .ZN(n8910) );
  INV_X1 U10387 ( .A(n8960), .ZN(n8905) );
  NAND2_X1 U10388 ( .A1(n9048), .A2(n8905), .ZN(n9054) );
  NAND2_X1 U10389 ( .A1(n9059), .A2(n9428), .ZN(n9050) );
  INV_X1 U10390 ( .A(n9067), .ZN(n8906) );
  AOI211_X1 U10391 ( .C1(n9057), .C2(n9054), .A(n9050), .B(n8906), .ZN(n8908)
         );
  OAI21_X1 U10392 ( .B1(n8908), .B2(n8907), .A(n9074), .ZN(n8909) );
  NAND2_X1 U10393 ( .A1(n9095), .A2(n9085), .ZN(n9081) );
  AOI21_X1 U10394 ( .B1(n9157), .B2(n8909), .A(n9081), .ZN(n9163) );
  OAI21_X1 U10395 ( .B1(n8911), .B2(n8910), .A(n9163), .ZN(n8912) );
  INV_X1 U10396 ( .A(n9188), .ZN(n8951) );
  NAND2_X1 U10397 ( .A1(n9323), .A2(n8951), .ZN(n8952) );
  NAND2_X1 U10398 ( .A1(n8952), .A2(n9098), .ZN(n9166) );
  AOI21_X1 U10399 ( .B1(n9160), .B2(n8912), .A(n9166), .ZN(n8914) );
  NAND2_X1 U10400 ( .A1(n8916), .A2(n9188), .ZN(n9102) );
  NOR2_X1 U10401 ( .A1(n9323), .A2(n9102), .ZN(n8913) );
  OAI22_X1 U10402 ( .A1(n8914), .A2(n8913), .B1(n9610), .B2(n8916), .ZN(n8917)
         );
  INV_X1 U10403 ( .A(n8916), .ZN(n8915) );
  NAND2_X1 U10404 ( .A1(n9105), .A2(n8915), .ZN(n9165) );
  AOI21_X1 U10405 ( .B1(n8917), .B2(n9165), .A(n9101), .ZN(n8920) );
  INV_X1 U10406 ( .A(n8918), .ZN(n8919) );
  NOR2_X1 U10407 ( .A1(n8920), .A2(n8919), .ZN(n8956) );
  INV_X1 U10408 ( .A(n9165), .ZN(n9175) );
  INV_X1 U10409 ( .A(n9406), .ZN(n9411) );
  NAND4_X1 U10410 ( .A1(n8922), .A2(n4291), .A3(n4480), .A4(n9118), .ZN(n8925)
         );
  NAND2_X1 U10411 ( .A1(n8923), .A2(n6017), .ZN(n8924) );
  NOR3_X1 U10412 ( .A1(n8925), .A2(n8924), .A3(n8972), .ZN(n8930) );
  INV_X1 U10413 ( .A(n8926), .ZN(n8929) );
  INV_X1 U10414 ( .A(n9872), .ZN(n8927) );
  NAND4_X1 U10415 ( .A1(n8930), .A2(n8929), .A3(n8928), .A4(n8927), .ZN(n8932)
         );
  NOR2_X1 U10416 ( .A1(n8932), .A2(n8931), .ZN(n8933) );
  NAND3_X1 U10417 ( .A1(n8934), .A2(n4507), .A3(n8933), .ZN(n8937) );
  INV_X1 U10418 ( .A(n8935), .ZN(n8936) );
  OR3_X1 U10419 ( .A1(n8938), .A2(n8937), .A3(n8936), .ZN(n8939) );
  NOR2_X1 U10420 ( .A1(n8940), .A2(n8939), .ZN(n8942) );
  NAND3_X1 U10421 ( .A1(n8943), .A2(n8942), .A3(n8941), .ZN(n8944) );
  NOR2_X1 U10422 ( .A1(n9512), .A2(n8944), .ZN(n8945) );
  NAND2_X1 U10423 ( .A1(n9495), .A2(n8945), .ZN(n8946) );
  NOR2_X1 U10424 ( .A1(n9463), .A2(n8946), .ZN(n8947) );
  XNOR2_X1 U10425 ( .A(n9484), .B(n9192), .ZN(n9478) );
  AND4_X1 U10426 ( .A1(n9427), .A2(n8947), .A3(n9441), .A4(n9478), .ZN(n8948)
         );
  NAND4_X1 U10427 ( .A1(n9375), .A2(n9411), .A3(n9393), .A4(n8948), .ZN(n8949)
         );
  OR4_X1 U10428 ( .A1(n8950), .A2(n9335), .A3(n6055), .A4(n8949), .ZN(n8954)
         );
  OR2_X1 U10429 ( .A1(n9323), .A2(n8951), .ZN(n9164) );
  NAND2_X1 U10430 ( .A1(n9164), .A2(n8952), .ZN(n8953) );
  NOR4_X1 U10431 ( .A1(n9101), .A2(n9175), .A3(n8954), .A4(n8953), .ZN(n9110)
         );
  NOR4_X1 U10432 ( .A1(n8956), .A2(n9110), .A3(n9308), .A4(n8955), .ZN(n9174)
         );
  MUX2_X1 U10433 ( .A(n8957), .B(n9104), .S(n9193), .Z(n8961) );
  NAND2_X1 U10434 ( .A1(n9152), .A2(n9104), .ZN(n8958) );
  OAI22_X1 U10435 ( .A1(n8961), .A2(n8960), .B1(n8959), .B2(n8958), .ZN(n9046)
         );
  NAND2_X1 U10436 ( .A1(n9143), .A2(n8962), .ZN(n9016) );
  NOR2_X1 U10437 ( .A1(n9011), .A2(n9111), .ZN(n8963) );
  AOI21_X1 U10438 ( .B1(n9016), .B2(n9141), .A(n8963), .ZN(n9026) );
  AOI21_X1 U10439 ( .B1(n9143), .B2(n9197), .A(n9111), .ZN(n9025) );
  NAND2_X1 U10440 ( .A1(n8964), .A2(n9121), .ZN(n8967) );
  NAND3_X1 U10441 ( .A1(n8967), .A2(n8966), .A3(n8965), .ZN(n8968) );
  NAND3_X1 U10442 ( .A1(n8968), .A2(n8971), .A3(n4311), .ZN(n8970) );
  NAND2_X1 U10443 ( .A1(n8970), .A2(n8969), .ZN(n8975) );
  OAI21_X1 U10444 ( .B1(n8973), .B2(n8972), .A(n8971), .ZN(n8974) );
  INV_X1 U10445 ( .A(n9847), .ZN(n9850) );
  NAND2_X1 U10446 ( .A1(n8977), .A2(n8976), .ZN(n8978) );
  MUX2_X1 U10447 ( .A(n8979), .B(n8978), .S(n9104), .Z(n8980) );
  INV_X1 U10448 ( .A(n8980), .ZN(n8981) );
  MUX2_X1 U10449 ( .A(n8983), .B(n8982), .S(n9104), .Z(n8984) );
  NAND2_X1 U10450 ( .A1(n8992), .A2(n8985), .ZN(n8986) );
  NAND2_X1 U10451 ( .A1(n8986), .A2(n9124), .ZN(n8987) );
  AND2_X1 U10452 ( .A1(n8997), .A2(n8993), .ZN(n9129) );
  NAND2_X1 U10453 ( .A1(n8987), .A2(n9129), .ZN(n8989) );
  INV_X1 U10454 ( .A(n9134), .ZN(n8988) );
  AOI21_X1 U10455 ( .B1(n8989), .B2(n9131), .A(n8988), .ZN(n9003) );
  OAI21_X1 U10456 ( .B1(n8992), .B2(n8991), .A(n8990), .ZN(n8994) );
  NAND2_X1 U10457 ( .A1(n8994), .A2(n8993), .ZN(n8996) );
  NAND3_X1 U10458 ( .A1(n8996), .A2(n9124), .A3(n8995), .ZN(n9001) );
  AND2_X1 U10459 ( .A1(n9134), .A2(n8997), .ZN(n9000) );
  INV_X1 U10460 ( .A(n8998), .ZN(n8999) );
  AOI21_X1 U10461 ( .B1(n9001), .B2(n9000), .A(n8999), .ZN(n9002) );
  MUX2_X1 U10462 ( .A(n9003), .B(n9002), .S(n9104), .Z(n9008) );
  NAND2_X1 U10463 ( .A1(n9141), .A2(n9137), .ZN(n9017) );
  OR2_X1 U10464 ( .A1(n9005), .A2(n9004), .ZN(n9136) );
  NAND2_X1 U10465 ( .A1(n9136), .A2(n9104), .ZN(n9018) );
  INV_X1 U10466 ( .A(n9133), .ZN(n9006) );
  NAND2_X1 U10467 ( .A1(n9014), .A2(n9111), .ZN(n9009) );
  OAI22_X1 U10468 ( .A1(n9017), .A2(n9018), .B1(n9006), .B2(n9009), .ZN(n9007)
         );
  OAI22_X1 U10469 ( .A1(n9141), .A2(n9104), .B1(n9136), .B2(n9009), .ZN(n9013)
         );
  OR2_X1 U10470 ( .A1(n9011), .A2(n9010), .ZN(n9142) );
  OAI21_X1 U10471 ( .B1(n9104), .B2(n9137), .A(n9142), .ZN(n9012) );
  NOR2_X1 U10472 ( .A1(n9013), .A2(n9012), .ZN(n9023) );
  INV_X1 U10473 ( .A(n9014), .ZN(n9015) );
  OR2_X1 U10474 ( .A1(n9016), .A2(n9015), .ZN(n9115) );
  NAND3_X1 U10475 ( .A1(n9115), .A2(n9104), .A3(n9141), .ZN(n9022) );
  INV_X1 U10476 ( .A(n9017), .ZN(n9020) );
  NOR2_X1 U10477 ( .A1(n9018), .A2(n9133), .ZN(n9019) );
  NAND2_X1 U10478 ( .A1(n9020), .A2(n9019), .ZN(n9021) );
  OAI21_X1 U10479 ( .B1(n9026), .B2(n9025), .A(n9024), .ZN(n9032) );
  INV_X1 U10480 ( .A(n9027), .ZN(n9028) );
  OAI211_X1 U10481 ( .C1(n9029), .C2(n9028), .A(n9151), .B(n9148), .ZN(n9030)
         );
  INV_X1 U10482 ( .A(n9030), .ZN(n9031) );
  NAND4_X1 U10483 ( .A1(n9032), .A2(n9031), .A3(n9152), .A4(n9156), .ZN(n9044)
         );
  OR2_X1 U10484 ( .A1(n9147), .A2(n9194), .ZN(n9035) );
  OR2_X1 U10485 ( .A1(n9594), .A2(n9036), .ZN(n9039) );
  AOI21_X1 U10486 ( .B1(n9194), .B2(n9195), .A(n9104), .ZN(n9033) );
  NAND2_X1 U10487 ( .A1(n9039), .A2(n9033), .ZN(n9034) );
  AOI21_X1 U10488 ( .B1(n9640), .B2(n9035), .A(n9034), .ZN(n9042) );
  NAND2_X1 U10489 ( .A1(n9195), .A2(n9104), .ZN(n9038) );
  OAI22_X1 U10490 ( .A1(n9594), .A2(n9038), .B1(n9036), .B2(n9111), .ZN(n9037)
         );
  INV_X1 U10491 ( .A(n9037), .ZN(n9040) );
  OAI22_X1 U10492 ( .A1(n9040), .A2(n9520), .B1(n9039), .B2(n9038), .ZN(n9041)
         );
  AOI22_X1 U10493 ( .A1(n9042), .A2(n9152), .B1(n9156), .B2(n9041), .ZN(n9043)
         );
  INV_X1 U10494 ( .A(n9047), .ZN(n9049) );
  INV_X1 U10495 ( .A(n9048), .ZN(n9440) );
  AOI21_X1 U10496 ( .B1(n9056), .B2(n9049), .A(n9440), .ZN(n9053) );
  INV_X1 U10497 ( .A(n9441), .ZN(n9052) );
  INV_X1 U10498 ( .A(n9050), .ZN(n9051) );
  OAI21_X1 U10499 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(n9064) );
  INV_X1 U10500 ( .A(n9054), .ZN(n9055) );
  INV_X1 U10501 ( .A(n9058), .ZN(n9061) );
  INV_X1 U10502 ( .A(n9059), .ZN(n9060) );
  AOI21_X1 U10503 ( .B1(n9062), .B2(n9061), .A(n9060), .ZN(n9063) );
  NAND3_X1 U10504 ( .A1(n9426), .A2(n9111), .A3(n9065), .ZN(n9066) );
  MUX2_X1 U10505 ( .A(n9068), .B(n9067), .S(n9111), .Z(n9069) );
  NAND2_X1 U10506 ( .A1(n9070), .A2(n9069), .ZN(n9076) );
  INV_X1 U10507 ( .A(n9074), .ZN(n9071) );
  OAI211_X1 U10508 ( .C1(n9076), .C2(n9071), .A(n9077), .B(n9073), .ZN(n9072)
         );
  NAND2_X1 U10509 ( .A1(n9072), .A2(n9365), .ZN(n9080) );
  INV_X1 U10510 ( .A(n9073), .ZN(n9075) );
  OAI21_X1 U10511 ( .B1(n9076), .B2(n9075), .A(n9074), .ZN(n9078) );
  AOI21_X1 U10512 ( .B1(n9078), .B2(n9077), .A(n9159), .ZN(n9079) );
  INV_X1 U10513 ( .A(n9081), .ZN(n9082) );
  INV_X1 U10514 ( .A(n9085), .ZN(n9086) );
  NAND2_X1 U10515 ( .A1(n9086), .A2(n9111), .ZN(n9087) );
  AND2_X1 U10516 ( .A1(n9091), .A2(n9087), .ZN(n9088) );
  NAND2_X1 U10517 ( .A1(n9091), .A2(n9090), .ZN(n9092) );
  NAND2_X1 U10518 ( .A1(n9092), .A2(n9111), .ZN(n9093) );
  MUX2_X1 U10519 ( .A(n9098), .B(n9097), .S(n9111), .Z(n9099) );
  INV_X1 U10520 ( .A(n9099), .ZN(n9100) );
  NAND2_X1 U10521 ( .A1(n9176), .A2(n9102), .ZN(n9108) );
  NAND3_X1 U10522 ( .A1(n9106), .A2(n9105), .A3(n9188), .ZN(n9107) );
  NAND2_X1 U10523 ( .A1(n9308), .A2(n9114), .ZN(n9112) );
  INV_X1 U10524 ( .A(n9110), .ZN(n9113) );
  OAI22_X1 U10525 ( .A1(n9113), .A2(n9112), .B1(n9111), .B2(n9177), .ZN(n9173)
         );
  INV_X1 U10526 ( .A(n5695), .ZN(n9171) );
  NOR2_X1 U10527 ( .A1(n9410), .A2(n9114), .ZN(n9170) );
  INV_X1 U10528 ( .A(n9115), .ZN(n9140) );
  NOR2_X1 U10529 ( .A1(n9117), .A2(n9116), .ZN(n9123) );
  AND2_X1 U10530 ( .A1(n9120), .A2(n9119), .ZN(n9122) );
  AND4_X1 U10531 ( .A1(n9123), .A2(n9122), .A3(n9121), .A4(n4311), .ZN(n9127)
         );
  AND2_X1 U10532 ( .A1(n9125), .A2(n9124), .ZN(n9126) );
  OAI211_X1 U10533 ( .C1(n9128), .C2(n9127), .A(n9131), .B(n9126), .ZN(n9135)
         );
  INV_X1 U10534 ( .A(n9129), .ZN(n9130) );
  NAND2_X1 U10535 ( .A1(n9131), .A2(n9130), .ZN(n9132) );
  NAND4_X1 U10536 ( .A1(n9135), .A2(n9134), .A3(n9133), .A4(n9132), .ZN(n9138)
         );
  NAND3_X1 U10537 ( .A1(n9138), .A2(n9137), .A3(n9136), .ZN(n9139) );
  NAND2_X1 U10538 ( .A1(n9140), .A2(n9139), .ZN(n9146) );
  INV_X1 U10539 ( .A(n9142), .ZN(n9144) );
  OAI21_X1 U10540 ( .B1(n4756), .B2(n9144), .A(n9143), .ZN(n9145) );
  NAND3_X1 U10541 ( .A1(n9146), .A2(n9510), .A3(n9145), .ZN(n9149) );
  NAND3_X1 U10542 ( .A1(n9149), .A2(n9148), .A3(n9147), .ZN(n9150) );
  NAND3_X1 U10543 ( .A1(n9152), .A2(n9151), .A3(n9150), .ZN(n9155) );
  INV_X1 U10544 ( .A(n9153), .ZN(n9154) );
  AOI21_X1 U10545 ( .B1(n9156), .B2(n9155), .A(n9154), .ZN(n9158) );
  OAI21_X1 U10546 ( .B1(n9159), .B2(n9158), .A(n9157), .ZN(n9162) );
  INV_X1 U10547 ( .A(n9160), .ZN(n9161) );
  AOI21_X1 U10548 ( .B1(n9163), .B2(n9162), .A(n9161), .ZN(n9167) );
  OAI211_X1 U10549 ( .C1(n9167), .C2(n9166), .A(n9165), .B(n9164), .ZN(n9168)
         );
  NAND2_X1 U10550 ( .A1(n9168), .A2(n9176), .ZN(n9169) );
  MUX2_X1 U10551 ( .A(n9171), .B(n9170), .S(n9169), .Z(n9172) );
  NOR2_X1 U10552 ( .A1(n9176), .A2(n9410), .ZN(n9178) );
  NOR3_X1 U10553 ( .A1(n9180), .A2(n9728), .A3(n9179), .ZN(n9181) );
  NAND3_X1 U10554 ( .A1(n9182), .A2(n9181), .A3(n9647), .ZN(n9183) );
  OAI211_X1 U10555 ( .C1(n9184), .C2(n9186), .A(n9183), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9185) );
  OAI21_X1 U10556 ( .B1(n9187), .B2(n9186), .A(n9185), .ZN(P1_U3242) );
  MUX2_X1 U10557 ( .A(n9188), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9211), .Z(
        P1_U3584) );
  MUX2_X1 U10558 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9368), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10559 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9189), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10560 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9394), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10561 ( .A(n9190), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9211), .Z(
        P1_U3579) );
  MUX2_X1 U10562 ( .A(n9432), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9211), .Z(
        P1_U3578) );
  MUX2_X1 U10563 ( .A(n9434), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9211), .Z(
        P1_U3576) );
  MUX2_X1 U10564 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9191), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10565 ( .A(n9192), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9211), .Z(
        P1_U3574) );
  MUX2_X1 U10566 ( .A(n9193), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9211), .Z(
        P1_U3573) );
  MUX2_X1 U10567 ( .A(n9194), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9211), .Z(
        P1_U3572) );
  MUX2_X1 U10568 ( .A(n9195), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9211), .Z(
        P1_U3571) );
  MUX2_X1 U10569 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9196), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10570 ( .A(n9197), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9211), .Z(
        P1_U3569) );
  MUX2_X1 U10571 ( .A(n9198), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9211), .Z(
        P1_U3568) );
  MUX2_X1 U10572 ( .A(n9199), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9211), .Z(
        P1_U3567) );
  MUX2_X1 U10573 ( .A(n9200), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9211), .Z(
        P1_U3566) );
  MUX2_X1 U10574 ( .A(n4510), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9211), .Z(
        P1_U3565) );
  MUX2_X1 U10575 ( .A(n9202), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9211), .Z(
        P1_U3564) );
  MUX2_X1 U10576 ( .A(n9203), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9211), .Z(
        P1_U3563) );
  MUX2_X1 U10577 ( .A(n9204), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9211), .Z(
        P1_U3562) );
  MUX2_X1 U10578 ( .A(n9205), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9211), .Z(
        P1_U3561) );
  MUX2_X1 U10579 ( .A(n9206), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9211), .Z(
        P1_U3560) );
  MUX2_X1 U10580 ( .A(n9207), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9211), .Z(
        P1_U3559) );
  MUX2_X1 U10581 ( .A(n9208), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9211), .Z(
        P1_U3558) );
  MUX2_X1 U10582 ( .A(n9209), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9211), .Z(
        P1_U3557) );
  MUX2_X1 U10583 ( .A(n6010), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9211), .Z(
        P1_U3556) );
  MUX2_X1 U10584 ( .A(n9210), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9211), .Z(
        P1_U3555) );
  MUX2_X1 U10585 ( .A(n9212), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9211), .Z(
        P1_U3554) );
  OAI211_X1 U10586 ( .C1(n9215), .C2(n9214), .A(n9778), .B(n9213), .ZN(n9223)
         );
  OAI211_X1 U10587 ( .C1(n9218), .C2(n9217), .A(n9827), .B(n9216), .ZN(n9222)
         );
  AOI22_X1 U10588 ( .A1(n9735), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9221) );
  NAND2_X1 U10589 ( .A1(n9835), .A2(n9219), .ZN(n9220) );
  NAND4_X1 U10590 ( .A1(n9223), .A2(n9222), .A3(n9221), .A4(n9220), .ZN(
        P1_U3244) );
  INV_X1 U10591 ( .A(n9224), .ZN(n9228) );
  INV_X1 U10592 ( .A(n9735), .ZN(n9838) );
  INV_X1 U10593 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9226) );
  NAND2_X1 U10594 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9225) );
  OAI21_X1 U10595 ( .B1(n9838), .B2(n9226), .A(n9225), .ZN(n9227) );
  AOI21_X1 U10596 ( .B1(n9228), .B2(n9835), .A(n9227), .ZN(n9237) );
  OAI211_X1 U10597 ( .C1(n9231), .C2(n9230), .A(n9827), .B(n9229), .ZN(n9236)
         );
  OAI211_X1 U10598 ( .C1(n9234), .C2(n9233), .A(n9778), .B(n9232), .ZN(n9235)
         );
  NAND3_X1 U10599 ( .A1(n9237), .A2(n9236), .A3(n9235), .ZN(P1_U3246) );
  NAND2_X1 U10600 ( .A1(n9735), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n9238) );
  OAI211_X1 U10601 ( .C1(n9782), .C2(n9240), .A(n9239), .B(n9238), .ZN(n9241)
         );
  INV_X1 U10602 ( .A(n9241), .ZN(n9251) );
  OAI211_X1 U10603 ( .C1(n9244), .C2(n9243), .A(n9778), .B(n9242), .ZN(n9250)
         );
  INV_X1 U10604 ( .A(n9245), .ZN(n9246) );
  OAI211_X1 U10605 ( .C1(n9248), .C2(n9247), .A(n9827), .B(n9246), .ZN(n9249)
         );
  NAND4_X1 U10606 ( .A1(n9252), .A2(n9251), .A3(n9250), .A4(n9249), .ZN(
        P1_U3247) );
  XNOR2_X1 U10607 ( .A(n9281), .B(n9600), .ZN(n9278) );
  NOR2_X1 U10608 ( .A1(n9808), .A2(n9253), .ZN(n9254) );
  AOI21_X1 U10609 ( .B1(n9808), .B2(n9253), .A(n9254), .ZN(n9802) );
  NOR2_X1 U10610 ( .A1(n9256), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9255) );
  AOI21_X1 U10611 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n9256), .A(n9255), .ZN(
        n9789) );
  OAI21_X1 U10612 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n9264), .A(n9257), .ZN(
        n9790) );
  NOR2_X1 U10613 ( .A1(n9789), .A2(n9790), .ZN(n9788) );
  AOI21_X1 U10614 ( .B1(n9796), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9788), .ZN(
        n9801) );
  NOR2_X1 U10615 ( .A1(n9802), .A2(n9801), .ZN(n9800) );
  AOI21_X1 U10616 ( .B1(n9808), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9800), .ZN(
        n9258) );
  NOR2_X1 U10617 ( .A1(n9258), .A2(n9265), .ZN(n9259) );
  XNOR2_X1 U10618 ( .A(n9258), .B(n9265), .ZN(n9813) );
  NOR2_X1 U10619 ( .A1(n5348), .A2(n9813), .ZN(n9812) );
  NOR2_X1 U10620 ( .A1(n9259), .A2(n9812), .ZN(n9279) );
  XOR2_X1 U10621 ( .A(n9278), .B(n9279), .Z(n9276) );
  NOR2_X1 U10622 ( .A1(n9808), .A2(n9260), .ZN(n9261) );
  AOI21_X1 U10623 ( .B1(n9808), .B2(n9260), .A(n9261), .ZN(n9804) );
  NAND2_X1 U10624 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9796), .ZN(n9262) );
  OAI21_X1 U10625 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9796), .A(n9262), .ZN(
        n9792) );
  NOR2_X1 U10626 ( .A1(n9792), .A2(n9793), .ZN(n9791) );
  NOR2_X1 U10627 ( .A1(n9804), .A2(n9805), .ZN(n9803) );
  NOR2_X1 U10628 ( .A1(n9266), .A2(n9265), .ZN(n9267) );
  XOR2_X1 U10629 ( .A(n9819), .B(n9266), .Z(n9816) );
  NOR2_X1 U10630 ( .A1(n7658), .A2(n9816), .ZN(n9815) );
  XNOR2_X1 U10631 ( .A(n9281), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9268) );
  AOI21_X1 U10632 ( .B1(n9269), .B2(n9268), .A(n9814), .ZN(n9270) );
  NAND2_X1 U10633 ( .A1(n9270), .A2(n9283), .ZN(n9275) );
  INV_X1 U10634 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9272) );
  OAI21_X1 U10635 ( .B1(n9838), .B2(n9272), .A(n9271), .ZN(n9273) );
  AOI21_X1 U10636 ( .B1(n9281), .B2(n9835), .A(n9273), .ZN(n9274) );
  OAI211_X1 U10637 ( .C1(n9276), .C2(n9824), .A(n9275), .B(n9274), .ZN(
        P1_U3259) );
  XNOR2_X1 U10638 ( .A(n9298), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9299) );
  AOI22_X1 U10639 ( .A1(n9279), .A2(n9278), .B1(n9277), .B2(n9600), .ZN(n9300)
         );
  XOR2_X1 U10640 ( .A(n9299), .B(n9300), .Z(n9292) );
  XNOR2_X1 U10641 ( .A(n9298), .B(n9280), .ZN(n9285) );
  NAND2_X1 U10642 ( .A1(n9281), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9282) );
  NAND2_X1 U10643 ( .A1(n9284), .A2(n9285), .ZN(n9294) );
  OAI21_X1 U10644 ( .B1(n9285), .B2(n9284), .A(n9294), .ZN(n9286) );
  NAND2_X1 U10645 ( .A1(n9286), .A2(n9827), .ZN(n9291) );
  NOR2_X1 U10646 ( .A1(n9782), .A2(n9287), .ZN(n9288) );
  AOI211_X1 U10647 ( .C1(n9735), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9289), .B(
        n9288), .ZN(n9290) );
  OAI211_X1 U10648 ( .C1(n9824), .C2(n9292), .A(n9291), .B(n9290), .ZN(
        P1_U3260) );
  OR2_X1 U10649 ( .A1(n9298), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U10650 ( .A1(n9834), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9296) );
  OR2_X1 U10651 ( .A1(n9834), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9295) );
  AND2_X1 U10652 ( .A1(n9296), .A2(n9295), .ZN(n9829) );
  NAND2_X1 U10653 ( .A1(n9830), .A2(n9829), .ZN(n9828) );
  NAND2_X1 U10654 ( .A1(n9828), .A2(n9296), .ZN(n9297) );
  XNOR2_X1 U10655 ( .A(n9297), .B(n9503), .ZN(n9304) );
  OAI22_X1 U10656 ( .A1(n9300), .A2(n9299), .B1(n9298), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n9825) );
  NAND2_X1 U10657 ( .A1(n9834), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9301) );
  OAI21_X1 U10658 ( .B1(n9834), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9301), .ZN(
        n9826) );
  NOR2_X1 U10659 ( .A1(n9825), .A2(n9826), .ZN(n9823) );
  INV_X1 U10660 ( .A(n9301), .ZN(n9302) );
  NOR2_X1 U10661 ( .A1(n9823), .A2(n9302), .ZN(n9303) );
  XNOR2_X1 U10662 ( .A(n9303), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9305) );
  AOI22_X1 U10663 ( .A1(n9304), .A2(n9827), .B1(n9778), .B2(n9305), .ZN(n9310)
         );
  INV_X1 U10664 ( .A(n9304), .ZN(n9307) );
  OAI21_X1 U10665 ( .B1(n9305), .B2(n9824), .A(n9782), .ZN(n9306) );
  AOI21_X1 U10666 ( .B1(n9307), .B2(n9827), .A(n9306), .ZN(n9309) );
  NAND2_X1 U10667 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9311) );
  OAI211_X1 U10668 ( .C1(n9313), .C2(n9838), .A(n9312), .B(n9311), .ZN(
        P1_U3262) );
  NAND2_X1 U10669 ( .A1(n9314), .A2(n9896), .ZN(n9317) );
  INV_X1 U10670 ( .A(n9315), .ZN(n9532) );
  NOR2_X1 U10671 ( .A1(n9532), .A2(n9523), .ZN(n9321) );
  AOI21_X1 U10672 ( .B1(n9523), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9321), .ZN(
        n9316) );
  OAI211_X1 U10673 ( .C1(n9606), .C2(n9526), .A(n9317), .B(n9316), .ZN(
        P1_U3263) );
  OAI211_X1 U10674 ( .C1(n9610), .C2(n9319), .A(n9892), .B(n9318), .ZN(n9533)
         );
  NOR2_X1 U10675 ( .A1(n9528), .A2(n9320), .ZN(n9322) );
  AOI211_X1 U10676 ( .C1(n9323), .C2(n9884), .A(n9322), .B(n9321), .ZN(n9324)
         );
  OAI21_X1 U10677 ( .B1(n9533), .B2(n9351), .A(n9324), .ZN(P1_U3264) );
  INV_X1 U10678 ( .A(n9325), .ZN(n9334) );
  NOR2_X1 U10679 ( .A1(n4474), .A2(n9526), .ZN(n9329) );
  OAI22_X1 U10680 ( .A1(n9327), .A2(n9501), .B1(n9326), .B2(n9346), .ZN(n9328)
         );
  AOI211_X1 U10681 ( .C1(n9330), .C2(n9896), .A(n9329), .B(n9328), .ZN(n9333)
         );
  NAND2_X1 U10682 ( .A1(n9331), .A2(n9346), .ZN(n9332) );
  OAI211_X1 U10683 ( .C1(n9334), .C2(n9530), .A(n9333), .B(n9332), .ZN(
        P1_U3356) );
  NAND2_X1 U10684 ( .A1(n9336), .A2(n9335), .ZN(n9337) );
  NAND2_X1 U10685 ( .A1(n9338), .A2(n9337), .ZN(n9341) );
  OAI22_X1 U10686 ( .A1(n9377), .A2(n9469), .B1(n9339), .B2(n9467), .ZN(n9340)
         );
  NAND2_X1 U10687 ( .A1(n9539), .A2(n9897), .ZN(n9356) );
  OAI22_X1 U10688 ( .A1(n9348), .A2(n9501), .B1(n9347), .B2(n9346), .ZN(n9353)
         );
  AOI21_X1 U10689 ( .B1(n9354), .B2(n9358), .A(n9909), .ZN(n9350) );
  NAND2_X1 U10690 ( .A1(n9350), .A2(n9349), .ZN(n9536) );
  NOR2_X1 U10691 ( .A1(n9536), .A2(n9351), .ZN(n9352) );
  AOI211_X1 U10692 ( .C1(n9884), .C2(n9354), .A(n9353), .B(n9352), .ZN(n9355)
         );
  OAI211_X1 U10693 ( .C1(n9537), .C2(n9900), .A(n9356), .B(n9355), .ZN(
        P1_U3265) );
  XNOR2_X1 U10694 ( .A(n9357), .B(n6055), .ZN(n9546) );
  INV_X1 U10695 ( .A(n9381), .ZN(n9360) );
  INV_X1 U10696 ( .A(n9358), .ZN(n9359) );
  AOI211_X1 U10697 ( .C1(n9543), .C2(n9360), .A(n9909), .B(n9359), .ZN(n9542)
         );
  AOI22_X1 U10698 ( .A1(n9361), .A2(n9886), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9523), .ZN(n9362) );
  OAI21_X1 U10699 ( .B1(n9363), .B2(n9526), .A(n9362), .ZN(n9371) );
  NAND2_X1 U10700 ( .A1(n9364), .A2(n9365), .ZN(n9367) );
  XNOR2_X1 U10701 ( .A(n9367), .B(n9366), .ZN(n9369) );
  AOI222_X1 U10702 ( .A1(n9882), .A2(n9369), .B1(n9394), .B2(n9433), .C1(n9368), .C2(n9431), .ZN(n9545) );
  NOR2_X1 U10703 ( .A1(n9545), .A2(n9900), .ZN(n9370) );
  OAI21_X1 U10704 ( .B1(n9530), .B2(n9546), .A(n9372), .ZN(P1_U3266) );
  XNOR2_X1 U10705 ( .A(n9373), .B(n9375), .ZN(n9549) );
  INV_X1 U10706 ( .A(n9549), .ZN(n9389) );
  OAI21_X1 U10707 ( .B1(n9375), .B2(n9374), .A(n9364), .ZN(n9376) );
  NAND2_X1 U10708 ( .A1(n9376), .A2(n9882), .ZN(n9380) );
  OAI22_X1 U10709 ( .A1(n9377), .A2(n9467), .B1(n9409), .B2(n9469), .ZN(n9378)
         );
  INV_X1 U10710 ( .A(n9378), .ZN(n9379) );
  NAND2_X1 U10711 ( .A1(n9380), .A2(n9379), .ZN(n9547) );
  INV_X1 U10712 ( .A(n9396), .ZN(n9382) );
  AOI211_X1 U10713 ( .C1(n9383), .C2(n9382), .A(n9909), .B(n9381), .ZN(n9548)
         );
  NAND2_X1 U10714 ( .A1(n9548), .A2(n9896), .ZN(n9386) );
  AOI22_X1 U10715 ( .A1(n9384), .A2(n9886), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9523), .ZN(n9385) );
  OAI211_X1 U10716 ( .C1(n9618), .C2(n9526), .A(n9386), .B(n9385), .ZN(n9387)
         );
  AOI21_X1 U10717 ( .B1(n9547), .B2(n9528), .A(n9387), .ZN(n9388) );
  OAI21_X1 U10718 ( .B1(n9389), .B2(n9530), .A(n9388), .ZN(P1_U3267) );
  XNOR2_X1 U10719 ( .A(n9390), .B(n9393), .ZN(n9556) );
  OAI21_X1 U10720 ( .B1(n9393), .B2(n9392), .A(n9391), .ZN(n9395) );
  AOI222_X1 U10721 ( .A1(n9882), .A2(n9395), .B1(n9394), .B2(n9431), .C1(n9432), .C2(n9433), .ZN(n9555) );
  INV_X1 U10722 ( .A(n9555), .ZN(n9403) );
  INV_X1 U10723 ( .A(n9405), .ZN(n9397) );
  AOI211_X1 U10724 ( .C1(n9553), .C2(n9397), .A(n9909), .B(n9396), .ZN(n9552)
         );
  NAND2_X1 U10725 ( .A1(n9552), .A2(n9896), .ZN(n9400) );
  AOI22_X1 U10726 ( .A1(n9398), .A2(n9886), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9523), .ZN(n9399) );
  OAI211_X1 U10727 ( .C1(n9401), .C2(n9526), .A(n9400), .B(n9399), .ZN(n9402)
         );
  AOI21_X1 U10728 ( .B1(n9403), .B2(n9528), .A(n9402), .ZN(n9404) );
  OAI21_X1 U10729 ( .B1(n9556), .B2(n9530), .A(n9404), .ZN(P1_U3268) );
  AOI211_X1 U10730 ( .C1(n9416), .C2(n9421), .A(n9909), .B(n9405), .ZN(n9558)
         );
  XNOR2_X1 U10731 ( .A(n9407), .B(n9406), .ZN(n9408) );
  OAI222_X1 U10732 ( .A1(n9467), .A2(n9409), .B1(n9469), .B2(n9447), .C1(n9408), .C2(n9465), .ZN(n9557) );
  AOI21_X1 U10733 ( .B1(n9558), .B2(n9410), .A(n9557), .ZN(n9419) );
  XNOR2_X1 U10734 ( .A(n9412), .B(n9411), .ZN(n9559) );
  NAND2_X1 U10735 ( .A1(n9559), .A2(n9897), .ZN(n9418) );
  OAI22_X1 U10736 ( .A1(n9414), .A2(n9501), .B1(n9413), .B2(n9528), .ZN(n9415)
         );
  AOI21_X1 U10737 ( .B1(n9416), .B2(n9884), .A(n9415), .ZN(n9417) );
  OAI211_X1 U10738 ( .C1(n9419), .C2(n9900), .A(n9418), .B(n9417), .ZN(
        P1_U3269) );
  XNOR2_X1 U10739 ( .A(n9420), .B(n9427), .ZN(n9566) );
  INV_X1 U10740 ( .A(n9449), .ZN(n9423) );
  INV_X1 U10741 ( .A(n9421), .ZN(n9422) );
  AOI211_X1 U10742 ( .C1(n9563), .C2(n9423), .A(n9909), .B(n9422), .ZN(n9562)
         );
  AOI22_X1 U10743 ( .A1(n9424), .A2(n9886), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9523), .ZN(n9425) );
  OAI21_X1 U10744 ( .B1(n9426), .B2(n9526), .A(n9425), .ZN(n9437) );
  NAND3_X1 U10745 ( .A1(n9443), .A2(n9428), .A3(n4767), .ZN(n9429) );
  NAND2_X1 U10746 ( .A1(n9430), .A2(n9429), .ZN(n9435) );
  AOI222_X1 U10747 ( .A1(n9882), .A2(n9435), .B1(n9434), .B2(n9433), .C1(n9432), .C2(n9431), .ZN(n9565) );
  NOR2_X1 U10748 ( .A1(n9565), .A2(n9523), .ZN(n9436) );
  AOI211_X1 U10749 ( .C1(n9562), .C2(n9896), .A(n9437), .B(n9436), .ZN(n9438)
         );
  OAI21_X1 U10750 ( .B1(n9566), .B2(n9530), .A(n9438), .ZN(P1_U3270) );
  XNOR2_X1 U10751 ( .A(n9439), .B(n9441), .ZN(n9569) );
  INV_X1 U10752 ( .A(n9569), .ZN(n9457) );
  NOR2_X1 U10753 ( .A1(n9441), .A2(n9440), .ZN(n9445) );
  INV_X1 U10754 ( .A(n9443), .ZN(n9444) );
  AOI21_X1 U10755 ( .B1(n9445), .B2(n9442), .A(n9444), .ZN(n9446) );
  OAI222_X1 U10756 ( .A1(n9469), .A2(n9448), .B1(n9467), .B2(n9447), .C1(n9465), .C2(n9446), .ZN(n9567) );
  AOI211_X1 U10757 ( .C1(n9450), .C2(n4467), .A(n9909), .B(n9449), .ZN(n9568)
         );
  NAND2_X1 U10758 ( .A1(n9568), .A2(n9896), .ZN(n9454) );
  INV_X1 U10759 ( .A(n9451), .ZN(n9452) );
  AOI22_X1 U10760 ( .A1(n9452), .A2(n9886), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9523), .ZN(n9453) );
  OAI211_X1 U10761 ( .C1(n9628), .C2(n9526), .A(n9454), .B(n9453), .ZN(n9455)
         );
  AOI21_X1 U10762 ( .B1(n9567), .B2(n9528), .A(n9455), .ZN(n9456) );
  OAI21_X1 U10763 ( .B1(n9457), .B2(n9530), .A(n9456), .ZN(P1_U3271) );
  XOR2_X1 U10764 ( .A(n9463), .B(n9458), .Z(n9576) );
  NAND2_X1 U10765 ( .A1(n9460), .A2(n9459), .ZN(n9462) );
  INV_X1 U10766 ( .A(n9442), .ZN(n9461) );
  AOI21_X1 U10767 ( .B1(n9463), .B2(n9462), .A(n9461), .ZN(n9464) );
  OAI222_X1 U10768 ( .A1(n9469), .A2(n9468), .B1(n9467), .B2(n9466), .C1(n9465), .C2(n9464), .ZN(n9572) );
  AOI211_X1 U10769 ( .C1(n9574), .C2(n9482), .A(n9909), .B(n9470), .ZN(n9573)
         );
  NAND2_X1 U10770 ( .A1(n9573), .A2(n9896), .ZN(n9474) );
  INV_X1 U10771 ( .A(n9471), .ZN(n9472) );
  AOI22_X1 U10772 ( .A1(n9472), .A2(n9886), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9523), .ZN(n9473) );
  OAI211_X1 U10773 ( .C1(n4465), .C2(n9526), .A(n9474), .B(n9473), .ZN(n9475)
         );
  AOI21_X1 U10774 ( .B1(n9572), .B2(n9528), .A(n9475), .ZN(n9476) );
  OAI21_X1 U10775 ( .B1(n9576), .B2(n9530), .A(n9476), .ZN(P1_U3272) );
  XNOR2_X1 U10776 ( .A(n9477), .B(n9478), .ZN(n9579) );
  INV_X1 U10777 ( .A(n9579), .ZN(n9490) );
  XNOR2_X1 U10778 ( .A(n8903), .B(n9478), .ZN(n9479) );
  NAND2_X1 U10779 ( .A1(n9479), .A2(n9882), .ZN(n9481) );
  NAND2_X1 U10780 ( .A1(n9481), .A2(n9480), .ZN(n9577) );
  INV_X1 U10781 ( .A(n9482), .ZN(n9483) );
  AOI211_X1 U10782 ( .C1(n9484), .C2(n9497), .A(n9909), .B(n9483), .ZN(n9578)
         );
  NAND2_X1 U10783 ( .A1(n9578), .A2(n9896), .ZN(n9487) );
  AOI22_X1 U10784 ( .A1(n9523), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9485), .B2(
        n9886), .ZN(n9486) );
  OAI211_X1 U10785 ( .C1(n6085), .C2(n9526), .A(n9487), .B(n9486), .ZN(n9488)
         );
  AOI21_X1 U10786 ( .B1(n9577), .B2(n9528), .A(n9488), .ZN(n9489) );
  OAI21_X1 U10787 ( .B1(n9490), .B2(n9530), .A(n9489), .ZN(P1_U3273) );
  XNOR2_X1 U10788 ( .A(n9491), .B(n9495), .ZN(n9492) );
  NAND2_X1 U10789 ( .A1(n9492), .A2(n9882), .ZN(n9494) );
  NAND2_X1 U10790 ( .A1(n9494), .A2(n9493), .ZN(n9582) );
  INV_X1 U10791 ( .A(n9582), .ZN(n9508) );
  XNOR2_X1 U10792 ( .A(n9496), .B(n9495), .ZN(n9584) );
  NAND2_X1 U10793 ( .A1(n9584), .A2(n9897), .ZN(n9507) );
  INV_X1 U10794 ( .A(n9518), .ZN(n9499) );
  INV_X1 U10795 ( .A(n9497), .ZN(n9498) );
  AOI211_X1 U10796 ( .C1(n9500), .C2(n9499), .A(n9909), .B(n9498), .ZN(n9583)
         );
  NOR2_X1 U10797 ( .A1(n9636), .A2(n9526), .ZN(n9505) );
  OAI22_X1 U10798 ( .A1(n9528), .A2(n9503), .B1(n9502), .B2(n9501), .ZN(n9504)
         );
  AOI211_X1 U10799 ( .C1(n9583), .C2(n9896), .A(n9505), .B(n9504), .ZN(n9506)
         );
  OAI211_X1 U10800 ( .C1(n9523), .C2(n9508), .A(n9507), .B(n9506), .ZN(
        P1_U3274) );
  XNOR2_X1 U10801 ( .A(n9509), .B(n9512), .ZN(n9589) );
  INV_X1 U10802 ( .A(n9589), .ZN(n9531) );
  NAND2_X1 U10803 ( .A1(n9511), .A2(n9510), .ZN(n9513) );
  XNOR2_X1 U10804 ( .A(n9513), .B(n9512), .ZN(n9514) );
  NAND2_X1 U10805 ( .A1(n9514), .A2(n9882), .ZN(n9516) );
  NAND2_X1 U10806 ( .A1(n9516), .A2(n9515), .ZN(n9587) );
  INV_X1 U10807 ( .A(n9517), .ZN(n9519) );
  AOI211_X1 U10808 ( .C1(n9520), .C2(n9519), .A(n9909), .B(n9518), .ZN(n9588)
         );
  NAND2_X1 U10809 ( .A1(n9588), .A2(n9896), .ZN(n9525) );
  INV_X1 U10810 ( .A(n9521), .ZN(n9522) );
  AOI22_X1 U10811 ( .A1(n9523), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9522), .B2(
        n9886), .ZN(n9524) );
  OAI211_X1 U10812 ( .C1(n9640), .C2(n9526), .A(n9525), .B(n9524), .ZN(n9527)
         );
  AOI21_X1 U10813 ( .B1(n9587), .B2(n9528), .A(n9527), .ZN(n9529) );
  OAI21_X1 U10814 ( .B1(n9531), .B2(n9530), .A(n9529), .ZN(P1_U3275) );
  AND2_X1 U10815 ( .A1(n9533), .A2(n9532), .ZN(n9607) );
  MUX2_X1 U10816 ( .A(n9534), .B(n9607), .S(n9994), .Z(n9535) );
  OAI21_X1 U10817 ( .B1(n9610), .B2(n9602), .A(n9535), .ZN(P1_U3552) );
  NAND2_X1 U10818 ( .A1(n9537), .A2(n9536), .ZN(n9538) );
  MUX2_X1 U10819 ( .A(n9540), .B(n9611), .S(n9994), .Z(n9541) );
  OAI21_X1 U10820 ( .B1(n4473), .B2(n9602), .A(n9541), .ZN(P1_U3550) );
  AOI21_X1 U10821 ( .B1(n9974), .B2(n9543), .A(n9542), .ZN(n9544) );
  OAI211_X1 U10822 ( .C1(n9546), .C2(n9931), .A(n9545), .B(n9544), .ZN(n9614)
         );
  MUX2_X1 U10823 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9614), .S(n9994), .Z(
        P1_U3549) );
  MUX2_X1 U10824 ( .A(n9550), .B(n9615), .S(n9998), .Z(n9551) );
  OAI21_X1 U10825 ( .B1(n9618), .B2(n9602), .A(n9551), .ZN(P1_U3548) );
  AOI21_X1 U10826 ( .B1(n9974), .B2(n9553), .A(n9552), .ZN(n9554) );
  OAI211_X1 U10827 ( .C1(n9556), .C2(n9931), .A(n9555), .B(n9554), .ZN(n9619)
         );
  MUX2_X1 U10828 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9619), .S(n9998), .Z(
        P1_U3547) );
  AOI211_X1 U10829 ( .C1(n9559), .C2(n9971), .A(n9558), .B(n9557), .ZN(n9620)
         );
  MUX2_X1 U10830 ( .A(n9560), .B(n9620), .S(n9998), .Z(n9561) );
  OAI21_X1 U10831 ( .B1(n9623), .B2(n9602), .A(n9561), .ZN(P1_U3546) );
  AOI21_X1 U10832 ( .B1(n9974), .B2(n9563), .A(n9562), .ZN(n9564) );
  OAI211_X1 U10833 ( .C1(n9566), .C2(n9931), .A(n9565), .B(n9564), .ZN(n9624)
         );
  MUX2_X1 U10834 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9624), .S(n9998), .Z(
        P1_U3545) );
  INV_X1 U10835 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9570) );
  AOI211_X1 U10836 ( .C1(n9971), .C2(n9569), .A(n9568), .B(n9567), .ZN(n9625)
         );
  MUX2_X1 U10837 ( .A(n9570), .B(n9625), .S(n9998), .Z(n9571) );
  OAI21_X1 U10838 ( .B1(n9628), .B2(n9602), .A(n9571), .ZN(P1_U3544) );
  AOI211_X1 U10839 ( .C1(n9974), .C2(n9574), .A(n9573), .B(n9572), .ZN(n9575)
         );
  OAI21_X1 U10840 ( .B1(n9931), .B2(n9576), .A(n9575), .ZN(n9629) );
  MUX2_X1 U10841 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9629), .S(n9998), .Z(
        P1_U3543) );
  AOI211_X1 U10842 ( .C1(n9579), .C2(n9971), .A(n9578), .B(n9577), .ZN(n9630)
         );
  MUX2_X1 U10843 ( .A(n9580), .B(n9630), .S(n9998), .Z(n9581) );
  OAI21_X1 U10844 ( .B1(n6085), .B2(n9602), .A(n9581), .ZN(P1_U3542) );
  AOI211_X1 U10845 ( .C1(n9584), .C2(n9971), .A(n9583), .B(n9582), .ZN(n9633)
         );
  MUX2_X1 U10846 ( .A(n9585), .B(n9633), .S(n9998), .Z(n9586) );
  OAI21_X1 U10847 ( .B1(n9636), .B2(n9602), .A(n9586), .ZN(P1_U3541) );
  AOI211_X1 U10848 ( .C1(n9589), .C2(n9971), .A(n9588), .B(n9587), .ZN(n9637)
         );
  MUX2_X1 U10849 ( .A(n9590), .B(n9637), .S(n9998), .Z(n9591) );
  OAI21_X1 U10850 ( .B1(n9640), .B2(n9602), .A(n9591), .ZN(P1_U3540) );
  AOI211_X1 U10851 ( .C1(n9974), .C2(n9594), .A(n9593), .B(n9592), .ZN(n9595)
         );
  OAI21_X1 U10852 ( .B1(n9596), .B2(n9931), .A(n9595), .ZN(n9641) );
  MUX2_X1 U10853 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9641), .S(n9998), .Z(
        P1_U3539) );
  AOI211_X1 U10854 ( .C1(n9599), .C2(n9971), .A(n9598), .B(n9597), .ZN(n9642)
         );
  MUX2_X1 U10855 ( .A(n9600), .B(n9642), .S(n9998), .Z(n9601) );
  OAI21_X1 U10856 ( .B1(n4461), .B2(n9602), .A(n9601), .ZN(P1_U3538) );
  MUX2_X1 U10857 ( .A(n9604), .B(n9603), .S(n9983), .Z(n9605) );
  OAI21_X1 U10858 ( .B1(n9606), .B2(n9645), .A(n9605), .ZN(P1_U3521) );
  MUX2_X1 U10859 ( .A(n9608), .B(n9607), .S(n9983), .Z(n9609) );
  OAI21_X1 U10860 ( .B1(n9610), .B2(n9645), .A(n9609), .ZN(P1_U3520) );
  MUX2_X1 U10861 ( .A(n9612), .B(n9611), .S(n9983), .Z(n9613) );
  OAI21_X1 U10862 ( .B1(n4473), .B2(n9645), .A(n9613), .ZN(P1_U3518) );
  MUX2_X1 U10863 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9614), .S(n9983), .Z(
        P1_U3517) );
  MUX2_X1 U10864 ( .A(n9616), .B(n9615), .S(n9983), .Z(n9617) );
  OAI21_X1 U10865 ( .B1(n9618), .B2(n9645), .A(n9617), .ZN(P1_U3516) );
  MUX2_X1 U10866 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9619), .S(n9983), .Z(
        P1_U3515) );
  MUX2_X1 U10867 ( .A(n9621), .B(n9620), .S(n9983), .Z(n9622) );
  OAI21_X1 U10868 ( .B1(n9623), .B2(n9645), .A(n9622), .ZN(P1_U3514) );
  MUX2_X1 U10869 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9624), .S(n9983), .Z(
        P1_U3513) );
  MUX2_X1 U10870 ( .A(n9626), .B(n9625), .S(n9983), .Z(n9627) );
  OAI21_X1 U10871 ( .B1(n9628), .B2(n9645), .A(n9627), .ZN(P1_U3512) );
  MUX2_X1 U10872 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9629), .S(n9983), .Z(
        P1_U3511) );
  MUX2_X1 U10873 ( .A(n9631), .B(n9630), .S(n9983), .Z(n9632) );
  OAI21_X1 U10874 ( .B1(n6085), .B2(n9645), .A(n9632), .ZN(P1_U3510) );
  MUX2_X1 U10875 ( .A(n9634), .B(n9633), .S(n9983), .Z(n9635) );
  OAI21_X1 U10876 ( .B1(n9636), .B2(n9645), .A(n9635), .ZN(P1_U3509) );
  MUX2_X1 U10877 ( .A(n9638), .B(n9637), .S(n9983), .Z(n9639) );
  OAI21_X1 U10878 ( .B1(n9640), .B2(n9645), .A(n9639), .ZN(P1_U3507) );
  MUX2_X1 U10879 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9641), .S(n9983), .Z(
        P1_U3504) );
  MUX2_X1 U10880 ( .A(n9643), .B(n9642), .S(n9983), .Z(n9644) );
  OAI21_X1 U10881 ( .B1(n4461), .B2(n9645), .A(n9644), .ZN(P1_U3501) );
  AND2_X1 U10882 ( .A1(n9647), .A2(n9646), .ZN(n9906) );
  MUX2_X1 U10883 ( .A(P1_D_REG_1__SCAN_IN), .B(n9648), .S(n9906), .Z(P1_U3440)
         );
  MUX2_X1 U10884 ( .A(P1_D_REG_0__SCAN_IN), .B(n9649), .S(n9906), .Z(P1_U3439)
         );
  NAND2_X1 U10885 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), 
        .ZN(n9651) );
  OAI22_X1 U10886 ( .A1(n9652), .A2(n9651), .B1(n9650), .B2(n7993), .ZN(n9653)
         );
  INV_X1 U10887 ( .A(n9653), .ZN(n9654) );
  OAI21_X1 U10888 ( .B1(n9655), .B2(n9658), .A(n9654), .ZN(P1_U3324) );
  OAI222_X1 U10889 ( .A1(n9659), .A2(P1_U3086), .B1(n9658), .B2(n9657), .C1(
        n9656), .C2(n7993), .ZN(P1_U3325) );
  MUX2_X1 U10890 ( .A(n9660), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI211_X1 U10891 ( .C1(n9663), .C2(n9662), .A(n9661), .B(n9824), .ZN(n9668)
         );
  AOI211_X1 U10892 ( .C1(n9666), .C2(n9665), .A(n9664), .B(n9814), .ZN(n9667)
         );
  AOI211_X1 U10893 ( .C1(n9835), .C2(n9669), .A(n9668), .B(n9667), .ZN(n9671)
         );
  NAND2_X1 U10894 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9670) );
  OAI211_X1 U10895 ( .C1(n9672), .C2(n9838), .A(n9671), .B(n9670), .ZN(
        P1_U3253) );
  INV_X1 U10896 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9686) );
  INV_X1 U10897 ( .A(n9673), .ZN(n9677) );
  INV_X1 U10898 ( .A(n9674), .ZN(n9676) );
  AOI211_X1 U10899 ( .C1(n9677), .C2(n9676), .A(n9675), .B(n9824), .ZN(n9682)
         );
  AOI211_X1 U10900 ( .C1(n9680), .C2(n9679), .A(n9678), .B(n9814), .ZN(n9681)
         );
  AOI211_X1 U10901 ( .C1(n9835), .C2(n9683), .A(n9682), .B(n9681), .ZN(n9685)
         );
  NAND2_X1 U10902 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9684) );
  OAI211_X1 U10903 ( .C1(n9838), .C2(n9686), .A(n9685), .B(n9684), .ZN(
        P1_U3250) );
  INV_X1 U10904 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9699) );
  NOR2_X1 U10905 ( .A1(n9688), .A2(n9687), .ZN(n9689) );
  NOR3_X1 U10906 ( .A1(n9824), .A2(n9690), .A3(n9689), .ZN(n9695) );
  AOI211_X1 U10907 ( .C1(n9693), .C2(n9692), .A(n9691), .B(n9814), .ZN(n9694)
         );
  AOI211_X1 U10908 ( .C1(n9835), .C2(n9696), .A(n9695), .B(n9694), .ZN(n9698)
         );
  NAND2_X1 U10909 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9697) );
  OAI211_X1 U10910 ( .C1(n9838), .C2(n9699), .A(n9698), .B(n9697), .ZN(
        P1_U3251) );
  OAI21_X1 U10911 ( .B1(n9701), .B2(n9707), .A(n9700), .ZN(n9721) );
  INV_X1 U10912 ( .A(n9721), .ZN(n9715) );
  INV_X1 U10913 ( .A(n9702), .ZN(n9704) );
  OAI22_X1 U10914 ( .A1(n9720), .A2(n9705), .B1(n9704), .B2(n9703), .ZN(n9713)
         );
  XNOR2_X1 U10915 ( .A(n9706), .B(n9707), .ZN(n9708) );
  OAI222_X1 U10916 ( .A1(n9712), .A2(n9711), .B1(n9710), .B2(n9709), .C1(n9708), .C2(n10024), .ZN(n9723) );
  AOI211_X1 U10917 ( .C1(n9715), .C2(n9714), .A(n9713), .B(n9723), .ZN(n9717)
         );
  AOI22_X1 U10918 ( .A1(n9719), .A2(n9718), .B1(n9717), .B2(n9716), .ZN(
        P2_U3220) );
  OAI22_X1 U10919 ( .A1(n9721), .A2(n10088), .B1(n9720), .B2(n10068), .ZN(
        n9722) );
  NOR2_X1 U10920 ( .A1(n9723), .A2(n9722), .ZN(n9726) );
  AOI22_X1 U10921 ( .A1(n10121), .A2(n9726), .B1(n9724), .B2(n10119), .ZN(
        P2_U3472) );
  INV_X1 U10922 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9725) );
  AOI22_X1 U10923 ( .A1(n10094), .A2(n9726), .B1(n9725), .B2(n10092), .ZN(
        P2_U3429) );
  XNOR2_X1 U10924 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10925 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10926 ( .A(n9727), .ZN(n9729) );
  NAND2_X1 U10927 ( .A1(n9728), .A2(n5081), .ZN(n9731) );
  NAND2_X1 U10928 ( .A1(n9729), .A2(n9731), .ZN(n9732) );
  MUX2_X1 U10929 ( .A(n9732), .B(n9731), .S(n9730), .Z(n9734) );
  NAND2_X1 U10930 ( .A1(n9734), .A2(n9733), .ZN(n9737) );
  AOI22_X1 U10931 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n9735), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9736) );
  OAI21_X1 U10932 ( .B1(n9738), .B2(n9737), .A(n9736), .ZN(P1_U3243) );
  INV_X1 U10933 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9753) );
  AOI21_X1 U10934 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9742) );
  NAND2_X1 U10935 ( .A1(n9778), .A2(n9742), .ZN(n9748) );
  AOI21_X1 U10936 ( .B1(n9745), .B2(n9744), .A(n9743), .ZN(n9746) );
  NAND2_X1 U10937 ( .A1(n9827), .A2(n9746), .ZN(n9747) );
  OAI211_X1 U10938 ( .C1(n9782), .C2(n9749), .A(n9748), .B(n9747), .ZN(n9750)
         );
  INV_X1 U10939 ( .A(n9750), .ZN(n9752) );
  NAND2_X1 U10940 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9751) );
  OAI211_X1 U10941 ( .C1(n9838), .C2(n9753), .A(n9752), .B(n9751), .ZN(
        P1_U3248) );
  INV_X1 U10942 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9768) );
  AOI21_X1 U10943 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(n9757) );
  NAND2_X1 U10944 ( .A1(n9778), .A2(n9757), .ZN(n9763) );
  AOI21_X1 U10945 ( .B1(n9760), .B2(n9759), .A(n9758), .ZN(n9761) );
  NAND2_X1 U10946 ( .A1(n9827), .A2(n9761), .ZN(n9762) );
  OAI211_X1 U10947 ( .C1(n9782), .C2(n9764), .A(n9763), .B(n9762), .ZN(n9765)
         );
  INV_X1 U10948 ( .A(n9765), .ZN(n9767) );
  NAND2_X1 U10949 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9766) );
  OAI211_X1 U10950 ( .C1(n9838), .C2(n9768), .A(n9767), .B(n9766), .ZN(
        P1_U3249) );
  INV_X1 U10951 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9787) );
  INV_X1 U10952 ( .A(n9769), .ZN(n9781) );
  AOI21_X1 U10953 ( .B1(n9772), .B2(n9771), .A(n9770), .ZN(n9773) );
  NAND2_X1 U10954 ( .A1(n9827), .A2(n9773), .ZN(n9780) );
  AOI21_X1 U10955 ( .B1(n9776), .B2(n9775), .A(n9774), .ZN(n9777) );
  NAND2_X1 U10956 ( .A1(n9778), .A2(n9777), .ZN(n9779) );
  OAI211_X1 U10957 ( .C1(n9782), .C2(n9781), .A(n9780), .B(n9779), .ZN(n9783)
         );
  INV_X1 U10958 ( .A(n9783), .ZN(n9786) );
  NAND2_X1 U10959 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9785) );
  OAI211_X1 U10960 ( .C1(n9838), .C2(n9787), .A(n9786), .B(n9785), .ZN(
        P1_U3254) );
  AOI211_X1 U10961 ( .C1(n9790), .C2(n9789), .A(n9788), .B(n9824), .ZN(n9795)
         );
  AOI211_X1 U10962 ( .C1(n9793), .C2(n9792), .A(n9791), .B(n9814), .ZN(n9794)
         );
  AOI211_X1 U10963 ( .C1(n9835), .C2(n9796), .A(n9795), .B(n9794), .ZN(n9798)
         );
  NAND2_X1 U10964 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9797) );
  OAI211_X1 U10965 ( .C1(n9799), .C2(n9838), .A(n9798), .B(n9797), .ZN(
        P1_U3256) );
  INV_X1 U10966 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9811) );
  AOI211_X1 U10967 ( .C1(n9802), .C2(n9801), .A(n9800), .B(n9824), .ZN(n9807)
         );
  AOI211_X1 U10968 ( .C1(n9805), .C2(n9804), .A(n9803), .B(n9814), .ZN(n9806)
         );
  AOI211_X1 U10969 ( .C1(n9835), .C2(n9808), .A(n9807), .B(n9806), .ZN(n9810)
         );
  NAND2_X1 U10970 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9809) );
  OAI211_X1 U10971 ( .C1(n9838), .C2(n9811), .A(n9810), .B(n9809), .ZN(
        P1_U3257) );
  AOI211_X1 U10972 ( .C1(n5348), .C2(n9813), .A(n9812), .B(n9824), .ZN(n9818)
         );
  AOI211_X1 U10973 ( .C1(n9816), .C2(n7658), .A(n9815), .B(n9814), .ZN(n9817)
         );
  AOI211_X1 U10974 ( .C1(n9835), .C2(n9819), .A(n9818), .B(n9817), .ZN(n9821)
         );
  NAND2_X1 U10975 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9820) );
  OAI211_X1 U10976 ( .C1(n9822), .C2(n9838), .A(n9821), .B(n9820), .ZN(
        P1_U3258) );
  AOI211_X1 U10977 ( .C1(n9826), .C2(n9825), .A(n9824), .B(n9823), .ZN(n9833)
         );
  OAI211_X1 U10978 ( .C1(n9830), .C2(n9829), .A(n9828), .B(n9827), .ZN(n9831)
         );
  INV_X1 U10979 ( .A(n9831), .ZN(n9832) );
  AOI211_X1 U10980 ( .C1(n9835), .C2(n9834), .A(n9833), .B(n9832), .ZN(n9837)
         );
  NAND2_X1 U10981 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9836) );
  OAI211_X1 U10982 ( .C1(n9838), .C2(n10127), .A(n9837), .B(n9836), .ZN(
        P1_U3261) );
  INV_X1 U10983 ( .A(n9839), .ZN(n9840) );
  AOI222_X1 U10984 ( .A1(n9841), .A2(n9884), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n9523), .C1(n9886), .C2(n9840), .ZN(n9845) );
  AOI22_X1 U10985 ( .A1(n9843), .A2(n9862), .B1(n9896), .B2(n9842), .ZN(n9844)
         );
  OAI211_X1 U10986 ( .C1(n9900), .C2(n9846), .A(n9845), .B(n9844), .ZN(
        P1_U3282) );
  XNOR2_X1 U10987 ( .A(n9848), .B(n9847), .ZN(n9854) );
  XNOR2_X1 U10988 ( .A(n9849), .B(n9850), .ZN(n9858) );
  NOR2_X1 U10989 ( .A1(n9858), .A2(n9851), .ZN(n9852) );
  AOI211_X1 U10990 ( .C1(n9882), .C2(n9854), .A(n9853), .B(n9852), .ZN(n9947)
         );
  INV_X1 U10991 ( .A(n9855), .ZN(n9856) );
  AOI222_X1 U10992 ( .A1(n9857), .A2(n9884), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n9523), .C1(n9886), .C2(n9856), .ZN(n9864) );
  INV_X1 U10993 ( .A(n9858), .ZN(n9950) );
  OAI211_X1 U10994 ( .C1(n9860), .C2(n9946), .A(n9892), .B(n9859), .ZN(n9945)
         );
  INV_X1 U10995 ( .A(n9945), .ZN(n9861) );
  AOI22_X1 U10996 ( .A1(n9950), .A2(n9862), .B1(n9896), .B2(n9861), .ZN(n9863)
         );
  OAI211_X1 U10997 ( .C1(n9900), .C2(n9947), .A(n9864), .B(n9863), .ZN(
        P1_U3286) );
  XNOR2_X1 U10998 ( .A(n9865), .B(n9872), .ZN(n9867) );
  AOI21_X1 U10999 ( .B1(n9867), .B2(n9882), .A(n9866), .ZN(n9935) );
  INV_X1 U11000 ( .A(n9868), .ZN(n9869) );
  AOI222_X1 U11001 ( .A1(n9870), .A2(n9884), .B1(n9869), .B2(n9886), .C1(
        P1_REG2_REG_5__SCAN_IN), .C2(n9900), .ZN(n9878) );
  XNOR2_X1 U11002 ( .A(n9871), .B(n9872), .ZN(n9938) );
  INV_X1 U11003 ( .A(n9873), .ZN(n9874) );
  OAI211_X1 U11004 ( .C1(n9934), .C2(n9875), .A(n9874), .B(n9892), .ZN(n9933)
         );
  INV_X1 U11005 ( .A(n9933), .ZN(n9876) );
  AOI22_X1 U11006 ( .A1(n9938), .A2(n9897), .B1(n9896), .B2(n9876), .ZN(n9877)
         );
  OAI211_X1 U11007 ( .C1(n9900), .C2(n9935), .A(n9878), .B(n9877), .ZN(
        P1_U3288) );
  XNOR2_X1 U11008 ( .A(n9880), .B(n9890), .ZN(n9883) );
  AOI21_X1 U11009 ( .B1(n9883), .B2(n9882), .A(n9881), .ZN(n9922) );
  AOI222_X1 U11010 ( .A1(n9887), .A2(n9886), .B1(P1_REG2_REG_3__SCAN_IN), .B2(
        n9523), .C1(n9885), .C2(n9884), .ZN(n9899) );
  NAND2_X1 U11011 ( .A1(n9889), .A2(n9888), .ZN(n9891) );
  XNOR2_X1 U11012 ( .A(n9891), .B(n9890), .ZN(n9925) );
  OAI211_X1 U11013 ( .C1(n9894), .C2(n9921), .A(n9893), .B(n9892), .ZN(n9920)
         );
  INV_X1 U11014 ( .A(n9920), .ZN(n9895) );
  AOI22_X1 U11015 ( .A1(n9925), .A2(n9897), .B1(n9896), .B2(n9895), .ZN(n9898)
         );
  OAI211_X1 U11016 ( .C1(n9900), .C2(n9922), .A(n9899), .B(n9898), .ZN(
        P1_U3290) );
  AND2_X1 U11017 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9907), .ZN(P1_U3294) );
  NOR2_X1 U11018 ( .A1(n9906), .A2(n9901), .ZN(P1_U3295) );
  AND2_X1 U11019 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9907), .ZN(P1_U3296) );
  NOR2_X1 U11020 ( .A1(n9906), .A2(n9902), .ZN(P1_U3297) );
  AND2_X1 U11021 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9907), .ZN(P1_U3298) );
  AND2_X1 U11022 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9907), .ZN(P1_U3299) );
  AND2_X1 U11023 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9907), .ZN(P1_U3300) );
  AND2_X1 U11024 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9907), .ZN(P1_U3301) );
  AND2_X1 U11025 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9907), .ZN(P1_U3302) );
  AND2_X1 U11026 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9907), .ZN(P1_U3303) );
  AND2_X1 U11027 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9907), .ZN(P1_U3304) );
  AND2_X1 U11028 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9907), .ZN(P1_U3305) );
  NOR2_X1 U11029 ( .A1(n9906), .A2(n9903), .ZN(P1_U3306) );
  AND2_X1 U11030 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9907), .ZN(P1_U3307) );
  AND2_X1 U11031 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9907), .ZN(P1_U3308) );
  AND2_X1 U11032 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9907), .ZN(P1_U3309) );
  AND2_X1 U11033 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9907), .ZN(P1_U3310) );
  AND2_X1 U11034 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9907), .ZN(P1_U3311) );
  AND2_X1 U11035 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9907), .ZN(P1_U3312) );
  NOR2_X1 U11036 ( .A1(n9906), .A2(n9904), .ZN(P1_U3313) );
  AND2_X1 U11037 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9907), .ZN(P1_U3314) );
  AND2_X1 U11038 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9907), .ZN(P1_U3315) );
  AND2_X1 U11039 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9907), .ZN(P1_U3316) );
  AND2_X1 U11040 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9907), .ZN(P1_U3317) );
  AND2_X1 U11041 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9907), .ZN(P1_U3318) );
  AND2_X1 U11042 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9907), .ZN(P1_U3319) );
  AND2_X1 U11043 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9907), .ZN(P1_U3320) );
  NOR2_X1 U11044 ( .A1(n9906), .A2(n9905), .ZN(P1_U3321) );
  AND2_X1 U11045 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9907), .ZN(P1_U3322) );
  AND2_X1 U11046 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9907), .ZN(P1_U3323) );
  INV_X1 U11047 ( .A(n9908), .ZN(n9910) );
  INV_X1 U11048 ( .A(n9974), .ZN(n9967) );
  AOI211_X1 U11049 ( .C1(n9957), .C2(n9913), .A(n9912), .B(n9911), .ZN(n9984)
         );
  AOI22_X1 U11050 ( .A1(n9983), .A2(n9984), .B1(n5049), .B2(n9982), .ZN(
        P1_U3456) );
  NAND2_X1 U11051 ( .A1(n9914), .A2(n9957), .ZN(n9916) );
  OAI211_X1 U11052 ( .C1(n9917), .C2(n9967), .A(n9916), .B(n9915), .ZN(n9918)
         );
  NOR2_X1 U11053 ( .A1(n9919), .A2(n9918), .ZN(n9986) );
  AOI22_X1 U11054 ( .A1(n9983), .A2(n9986), .B1(n5036), .B2(n9982), .ZN(
        P1_U3459) );
  OAI21_X1 U11055 ( .B1(n9921), .B2(n9967), .A(n9920), .ZN(n9924) );
  INV_X1 U11056 ( .A(n9922), .ZN(n9923) );
  AOI211_X1 U11057 ( .C1(n9925), .C2(n9971), .A(n9924), .B(n9923), .ZN(n9987)
         );
  AOI22_X1 U11058 ( .A1(n9983), .A2(n9987), .B1(n5091), .B2(n9982), .ZN(
        P1_U3462) );
  AOI21_X1 U11059 ( .B1(n9974), .B2(n9927), .A(n9926), .ZN(n9928) );
  OAI211_X1 U11060 ( .C1(n9931), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9932)
         );
  INV_X1 U11061 ( .A(n9932), .ZN(n9988) );
  AOI22_X1 U11062 ( .A1(n9983), .A2(n9988), .B1(n5020), .B2(n9982), .ZN(
        P1_U3465) );
  OAI21_X1 U11063 ( .B1(n9934), .B2(n9967), .A(n9933), .ZN(n9937) );
  INV_X1 U11064 ( .A(n9935), .ZN(n9936) );
  AOI211_X1 U11065 ( .C1(n9938), .C2(n9971), .A(n9937), .B(n9936), .ZN(n9989)
         );
  AOI22_X1 U11066 ( .A1(n9983), .A2(n9989), .B1(n5132), .B2(n9982), .ZN(
        P1_U3468) );
  OAI21_X1 U11067 ( .B1(n9940), .B2(n9967), .A(n9939), .ZN(n9943) );
  INV_X1 U11068 ( .A(n9941), .ZN(n9942) );
  AOI211_X1 U11069 ( .C1(n9971), .C2(n9944), .A(n9943), .B(n9942), .ZN(n9990)
         );
  AOI22_X1 U11070 ( .A1(n9983), .A2(n9990), .B1(n5112), .B2(n9982), .ZN(
        P1_U3471) );
  OAI21_X1 U11071 ( .B1(n9946), .B2(n9967), .A(n9945), .ZN(n9949) );
  INV_X1 U11072 ( .A(n9947), .ZN(n9948) );
  AOI211_X1 U11073 ( .C1(n9957), .C2(n9950), .A(n9949), .B(n9948), .ZN(n9991)
         );
  AOI22_X1 U11074 ( .A1(n9983), .A2(n9991), .B1(n5161), .B2(n9982), .ZN(
        P1_U3474) );
  INV_X1 U11075 ( .A(n9951), .ZN(n9956) );
  OAI21_X1 U11076 ( .B1(n9953), .B2(n9967), .A(n9952), .ZN(n9955) );
  AOI211_X1 U11077 ( .C1(n9957), .C2(n9956), .A(n9955), .B(n9954), .ZN(n9992)
         );
  AOI22_X1 U11078 ( .A1(n9983), .A2(n9992), .B1(n5203), .B2(n9982), .ZN(
        P1_U3477) );
  INV_X1 U11079 ( .A(n9958), .ZN(n9964) );
  OAI21_X1 U11080 ( .B1(n4468), .B2(n9967), .A(n9960), .ZN(n9963) );
  INV_X1 U11081 ( .A(n9961), .ZN(n9962) );
  AOI211_X1 U11082 ( .C1(n9971), .C2(n9964), .A(n9963), .B(n9962), .ZN(n9993)
         );
  AOI22_X1 U11083 ( .A1(n9983), .A2(n9993), .B1(n5181), .B2(n9982), .ZN(
        P1_U3480) );
  OAI211_X1 U11084 ( .C1(n9968), .C2(n9967), .A(n9966), .B(n9965), .ZN(n9969)
         );
  AOI21_X1 U11085 ( .B1(n9971), .B2(n9970), .A(n9969), .ZN(n9995) );
  AOI22_X1 U11086 ( .A1(n9983), .A2(n9995), .B1(n5253), .B2(n9982), .ZN(
        P1_U3483) );
  AOI21_X1 U11087 ( .B1(n9974), .B2(n9973), .A(n9972), .ZN(n9975) );
  OAI211_X1 U11088 ( .C1(n9978), .C2(n9977), .A(n9976), .B(n9975), .ZN(n9979)
         );
  AOI21_X1 U11089 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(n9997) );
  AOI22_X1 U11090 ( .A1(n9983), .A2(n9997), .B1(n5328), .B2(n9982), .ZN(
        P1_U3495) );
  AOI22_X1 U11091 ( .A1(n9998), .A2(n9984), .B1(n5054), .B2(n9996), .ZN(
        P1_U3523) );
  AOI22_X1 U11092 ( .A1(n9994), .A2(n9986), .B1(n9985), .B2(n9996), .ZN(
        P1_U3524) );
  AOI22_X1 U11093 ( .A1(n9994), .A2(n9987), .B1(n6607), .B2(n9996), .ZN(
        P1_U3525) );
  AOI22_X1 U11094 ( .A1(n9994), .A2(n9988), .B1(n5019), .B2(n9996), .ZN(
        P1_U3526) );
  AOI22_X1 U11095 ( .A1(n9994), .A2(n9989), .B1(n5125), .B2(n9996), .ZN(
        P1_U3527) );
  AOI22_X1 U11096 ( .A1(n9994), .A2(n9990), .B1(n5113), .B2(n9996), .ZN(
        P1_U3528) );
  AOI22_X1 U11097 ( .A1(n9994), .A2(n9991), .B1(n6603), .B2(n9996), .ZN(
        P1_U3529) );
  AOI22_X1 U11098 ( .A1(n9998), .A2(n9992), .B1(n5209), .B2(n9996), .ZN(
        P1_U3530) );
  AOI22_X1 U11099 ( .A1(n9994), .A2(n9993), .B1(n5180), .B2(n9996), .ZN(
        P1_U3531) );
  AOI22_X1 U11100 ( .A1(n9998), .A2(n9995), .B1(n6868), .B2(n9996), .ZN(
        P1_U3532) );
  AOI22_X1 U11101 ( .A1(n9998), .A2(n9997), .B1(n9253), .B2(n9996), .ZN(
        P1_U3536) );
  INV_X1 U11102 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10022) );
  INV_X1 U11103 ( .A(n9999), .ZN(n10005) );
  OAI21_X1 U11104 ( .B1(n10002), .B2(n10001), .A(n10000), .ZN(n10004) );
  AOI22_X1 U11105 ( .A1(n10005), .A2(n10004), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(P2_U3151), .ZN(n10011) );
  OAI211_X1 U11106 ( .C1(n10009), .C2(n10008), .A(n10007), .B(n10006), .ZN(
        n10010) );
  OAI211_X1 U11107 ( .C1(n5954), .C2(n10012), .A(n10011), .B(n10010), .ZN(
        n10013) );
  INV_X1 U11108 ( .A(n10013), .ZN(n10020) );
  OAI21_X1 U11109 ( .B1(n10015), .B2(n10017), .A(n10016), .ZN(n10018) );
  NAND2_X1 U11110 ( .A1(n4658), .A2(n10018), .ZN(n10019) );
  OAI211_X1 U11111 ( .C1(n10022), .C2(n10021), .A(n10020), .B(n10019), .ZN(
        P2_U3184) );
  AOI21_X1 U11112 ( .B1(n10024), .B2(n10088), .A(n10023), .ZN(n10025) );
  AOI211_X1 U11113 ( .C1(n10028), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        n10096) );
  INV_X1 U11114 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10029) );
  AOI22_X1 U11115 ( .A1(n10094), .A2(n10096), .B1(n10029), .B2(n10092), .ZN(
        P2_U3390) );
  AOI211_X1 U11116 ( .C1(n10072), .C2(n10032), .A(n10031), .B(n10030), .ZN(
        n10098) );
  INV_X1 U11117 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10033) );
  AOI22_X1 U11118 ( .A1(n10094), .A2(n10098), .B1(n10033), .B2(n10092), .ZN(
        P2_U3393) );
  INV_X1 U11119 ( .A(n10034), .ZN(n10037) );
  AOI211_X1 U11120 ( .C1(n10072), .C2(n10037), .A(n10036), .B(n10035), .ZN(
        n10100) );
  INV_X1 U11121 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U11122 ( .A1(n10094), .A2(n10100), .B1(n10038), .B2(n10092), .ZN(
        P2_U3396) );
  INV_X1 U11123 ( .A(n10039), .ZN(n10040) );
  AOI211_X1 U11124 ( .C1(n10084), .C2(n10042), .A(n10041), .B(n10040), .ZN(
        n10102) );
  AOI22_X1 U11125 ( .A1(n10094), .A2(n10102), .B1(n6140), .B2(n10092), .ZN(
        P2_U3399) );
  INV_X1 U11126 ( .A(n10043), .ZN(n10044) );
  AOI211_X1 U11127 ( .C1(n10046), .C2(n10084), .A(n10045), .B(n10044), .ZN(
        n10104) );
  INV_X1 U11128 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10047) );
  AOI22_X1 U11129 ( .A1(n10094), .A2(n10104), .B1(n10047), .B2(n10092), .ZN(
        P2_U3402) );
  AND2_X1 U11130 ( .A1(n10048), .A2(n10072), .ZN(n10050) );
  NOR3_X1 U11131 ( .A1(n10051), .A2(n10050), .A3(n10049), .ZN(n10106) );
  INV_X1 U11132 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10052) );
  AOI22_X1 U11133 ( .A1(n10094), .A2(n10106), .B1(n10052), .B2(n10092), .ZN(
        P2_U3405) );
  OAI211_X1 U11134 ( .C1(n10088), .C2(n10055), .A(n10054), .B(n10053), .ZN(
        n10056) );
  INV_X1 U11135 ( .A(n10056), .ZN(n10108) );
  INV_X1 U11136 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10057) );
  AOI22_X1 U11137 ( .A1(n10094), .A2(n10108), .B1(n10057), .B2(n10092), .ZN(
        P2_U3408) );
  INV_X1 U11138 ( .A(n10058), .ZN(n10059) );
  AOI211_X1 U11139 ( .C1(n10072), .C2(n10061), .A(n10060), .B(n10059), .ZN(
        n10110) );
  INV_X1 U11140 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10062) );
  AOI22_X1 U11141 ( .A1(n10094), .A2(n10110), .B1(n10062), .B2(n10092), .ZN(
        P2_U3411) );
  OAI22_X1 U11142 ( .A1(n10064), .A2(n10088), .B1(n10063), .B2(n10068), .ZN(
        n10065) );
  NOR2_X1 U11143 ( .A1(n10066), .A2(n10065), .ZN(n10112) );
  INV_X1 U11144 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U11145 ( .A1(n10094), .A2(n10112), .B1(n10067), .B2(n10092), .ZN(
        P2_U3414) );
  NOR2_X1 U11146 ( .A1(n10069), .A2(n10068), .ZN(n10071) );
  AOI211_X1 U11147 ( .C1(n10073), .C2(n10072), .A(n10071), .B(n10070), .ZN(
        n10114) );
  INV_X1 U11148 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10074) );
  AOI22_X1 U11149 ( .A1(n10094), .A2(n10114), .B1(n10074), .B2(n10092), .ZN(
        P2_U3417) );
  OAI21_X1 U11150 ( .B1(n10077), .B2(n10076), .A(n10075), .ZN(n10078) );
  NOR2_X1 U11151 ( .A1(n10079), .A2(n10078), .ZN(n10116) );
  AOI22_X1 U11152 ( .A1(n10094), .A2(n10116), .B1(n10080), .B2(n10092), .ZN(
        P2_U3420) );
  INV_X1 U11153 ( .A(n10081), .ZN(n10083) );
  AOI211_X1 U11154 ( .C1(n10085), .C2(n10084), .A(n10083), .B(n10082), .ZN(
        n10118) );
  INV_X1 U11155 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10086) );
  AOI22_X1 U11156 ( .A1(n10094), .A2(n10118), .B1(n10086), .B2(n10092), .ZN(
        P2_U3423) );
  OAI21_X1 U11157 ( .B1(n10089), .B2(n10088), .A(n10087), .ZN(n10090) );
  NOR2_X1 U11158 ( .A1(n10091), .A2(n10090), .ZN(n10120) );
  INV_X1 U11159 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10093) );
  AOI22_X1 U11160 ( .A1(n10094), .A2(n10120), .B1(n10093), .B2(n10092), .ZN(
        P2_U3426) );
  AOI22_X1 U11161 ( .A1(n10121), .A2(n10096), .B1(n10095), .B2(n10119), .ZN(
        P2_U3459) );
  AOI22_X1 U11162 ( .A1(n10121), .A2(n10098), .B1(n10097), .B2(n10119), .ZN(
        P2_U3460) );
  INV_X1 U11163 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U11164 ( .A1(n10121), .A2(n10100), .B1(n10099), .B2(n10119), .ZN(
        P2_U3461) );
  AOI22_X1 U11165 ( .A1(n10121), .A2(n10102), .B1(n10101), .B2(n10119), .ZN(
        P2_U3462) );
  AOI22_X1 U11166 ( .A1(n10121), .A2(n10104), .B1(n10103), .B2(n10119), .ZN(
        P2_U3463) );
  AOI22_X1 U11167 ( .A1(n10121), .A2(n10106), .B1(n10105), .B2(n10119), .ZN(
        P2_U3464) );
  AOI22_X1 U11168 ( .A1(n10121), .A2(n10108), .B1(n10107), .B2(n10119), .ZN(
        P2_U3465) );
  AOI22_X1 U11169 ( .A1(n10121), .A2(n10110), .B1(n10109), .B2(n10119), .ZN(
        P2_U3466) );
  INV_X1 U11170 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U11171 ( .A1(n10121), .A2(n10112), .B1(n10111), .B2(n10119), .ZN(
        P2_U3467) );
  AOI22_X1 U11172 ( .A1(n10121), .A2(n10114), .B1(n10113), .B2(n10119), .ZN(
        P2_U3468) );
  AOI22_X1 U11173 ( .A1(n10121), .A2(n10116), .B1(n10115), .B2(n10119), .ZN(
        P2_U3469) );
  AOI22_X1 U11174 ( .A1(n10121), .A2(n10118), .B1(n10117), .B2(n10119), .ZN(
        P2_U3470) );
  AOI22_X1 U11175 ( .A1(n10121), .A2(n10120), .B1(n4372), .B2(n10119), .ZN(
        P2_U3471) );
  OAI222_X1 U11176 ( .A1(n6686), .A2(n10125), .B1(n6686), .B2(n10124), .C1(
        n10123), .C2(n10122), .ZN(ADD_1068_U5) );
  XOR2_X1 U11177 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11178 ( .B1(n10128), .B2(n10127), .A(n10126), .ZN(n10130) );
  XNOR2_X1 U11179 ( .A(n10130), .B(n10129), .ZN(ADD_1068_U55) );
  OAI21_X1 U11180 ( .B1(n10133), .B2(n10132), .A(n10131), .ZN(ADD_1068_U56) );
  OAI21_X1 U11181 ( .B1(n10136), .B2(n10135), .A(n10134), .ZN(ADD_1068_U57) );
  OAI21_X1 U11182 ( .B1(n10139), .B2(n10138), .A(n10137), .ZN(ADD_1068_U58) );
  OAI21_X1 U11183 ( .B1(n10142), .B2(n10141), .A(n10140), .ZN(ADD_1068_U59) );
  OAI21_X1 U11184 ( .B1(n10145), .B2(n10144), .A(n10143), .ZN(ADD_1068_U60) );
  OAI21_X1 U11185 ( .B1(n10148), .B2(n10147), .A(n10146), .ZN(ADD_1068_U61) );
  OAI21_X1 U11186 ( .B1(n10151), .B2(n10150), .A(n10149), .ZN(ADD_1068_U62) );
  OAI21_X1 U11187 ( .B1(n10154), .B2(n10153), .A(n10152), .ZN(ADD_1068_U63) );
  OAI21_X1 U11188 ( .B1(n10157), .B2(n10156), .A(n10155), .ZN(ADD_1068_U50) );
  OAI21_X1 U11189 ( .B1(n10160), .B2(n10159), .A(n10158), .ZN(ADD_1068_U51) );
  OAI21_X1 U11190 ( .B1(n10163), .B2(n10162), .A(n10161), .ZN(ADD_1068_U47) );
  OAI21_X1 U11191 ( .B1(n10166), .B2(n10165), .A(n10164), .ZN(ADD_1068_U49) );
  OAI21_X1 U11192 ( .B1(n10169), .B2(n10168), .A(n10167), .ZN(ADD_1068_U48) );
  AOI21_X1 U11193 ( .B1(n10172), .B2(n10171), .A(n10170), .ZN(ADD_1068_U54) );
  AOI21_X1 U11194 ( .B1(n10175), .B2(n10174), .A(n10173), .ZN(ADD_1068_U53) );
  OAI21_X1 U11195 ( .B1(n10178), .B2(n10177), .A(n10176), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4980 ( .A(n5096), .Z(n5987) );
  CLKBUF_X1 U4981 ( .A(n6155), .Z(n6443) );
  CLKBUF_X1 U5249 ( .A(n5199), .Z(n5986) );
endmodule

