

module b22_C_SARLock_k_64_10 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15191;

  INV_X4 U7182 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NAND2_X1 U7183 ( .A1(n6939), .A2(n6938), .ZN(n13801) );
  AND2_X1 U7184 ( .A1(n13994), .A2(n11612), .ZN(n13793) );
  NOR2_X1 U7185 ( .A1(n11384), .A2(n11096), .ZN(n12008) );
  NAND2_X1 U7186 ( .A1(n7903), .A2(n7902), .ZN(n10933) );
  NAND3_X1 U7187 ( .A1(n10469), .A2(n7008), .A3(n14692), .ZN(n10748) );
  AND2_X1 U7188 ( .A1(n14684), .A2(n14676), .ZN(n7008) );
  INV_X1 U7189 ( .A(n13367), .ZN(n7444) );
  INV_X2 U7190 ( .A(n13264), .ZN(n6443) );
  INV_X1 U7191 ( .A(n7762), .ZN(n9305) );
  BUF_X2 U7192 ( .A(n7769), .Z(n9306) );
  CLKBUF_X3 U7193 ( .A(n9213), .Z(n6445) );
  XNOR2_X1 U7194 ( .A(n7675), .B(n7674), .ZN(n11429) );
  NAND2_X1 U7195 ( .A1(n8382), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8386) );
  OR2_X1 U7196 ( .A1(n8411), .A2(n9629), .ZN(n8390) );
  BUF_X2 U7197 ( .A(n8405), .Z(n6449) );
  OAI21_X1 U7198 ( .B1(n8318), .B2(n8314), .A(n8319), .ZN(n8969) );
  NOR2_X1 U7199 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7652) );
  OR2_X1 U7200 ( .A1(n13016), .A2(n13142), .ZN(n12993) );
  NOR2_X2 U7201 ( .A1(n13067), .A2(n13157), .ZN(n13041) );
  OR2_X2 U7202 ( .A1(n11393), .A2(n11394), .ZN(n8179) );
  AND2_X1 U7203 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n14775), .ZN(n6433) );
  NOR2_X1 U7204 ( .A1(n6433), .A2(n14768), .ZN(n10897) );
  NAND2_X1 U7205 ( .A1(n6437), .A2(n8969), .ZN(n6447) );
  NAND2_X1 U7206 ( .A1(n7218), .A2(SI_3_), .ZN(n7591) );
  XNOR2_X1 U7207 ( .A(n8349), .B(P3_IR_REG_30__SCAN_IN), .ZN(n8351) );
  INV_X1 U7208 ( .A(n12604), .ZN(n12576) );
  CLKBUF_X2 U7210 ( .A(n8781), .Z(n6436) );
  XNOR2_X1 U7211 ( .A(n8322), .B(n8321), .ZN(n8968) );
  INV_X1 U7212 ( .A(n10731), .ZN(n14692) );
  INV_X1 U7213 ( .A(n13484), .ZN(n6749) );
  INV_X2 U7214 ( .A(n15191), .ZN(n11731) );
  INV_X2 U7215 ( .A(n11044), .ZN(n11726) );
  OR2_X1 U7216 ( .A1(n13890), .A2(n13699), .ZN(n13673) );
  INV_X1 U7217 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n13973) );
  INV_X1 U7218 ( .A(n10892), .ZN(n10839) );
  XNOR2_X1 U7219 ( .A(n10904), .B(n10905), .ZN(n14858) );
  INV_X1 U7220 ( .A(n12954), .ZN(n13124) );
  NAND2_X1 U7221 ( .A1(n7983), .A2(n7982), .ZN(n13134) );
  INV_X1 U7222 ( .A(n12923), .ZN(n13113) );
  INV_X1 U7223 ( .A(n12909), .ZN(n13108) );
  INV_X2 U7224 ( .A(n10022), .ZN(n6438) );
  INV_X1 U7225 ( .A(n13700), .ZN(n13898) );
  NAND2_X1 U7226 ( .A1(n10559), .A2(n7184), .ZN(n10994) );
  NAND2_X1 U7227 ( .A1(n7073), .A2(n14063), .ZN(n14065) );
  NAND2_X1 U7228 ( .A1(n7771), .A2(n7772), .ZN(n12744) );
  XNOR2_X1 U7229 ( .A(n14065), .B(n6818), .ZN(n15147) );
  OR2_X1 U7230 ( .A1(n6929), .A2(n6928), .ZN(n6434) );
  NAND2_X2 U7231 ( .A1(n9061), .A2(n9062), .ZN(n6452) );
  XNOR2_X2 U7232 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14044) );
  OAI21_X2 U7233 ( .B1(n6484), .B2(P3_IR_REG_23__SCAN_IN), .A(n6780), .ZN(
        n8959) );
  NAND2_X2 U7234 ( .A1(n12962), .A2(n8189), .ZN(n12945) );
  OAI21_X2 U7235 ( .B1(n12992), .B2(n7529), .A(n7528), .ZN(n12962) );
  NAND2_X2 U7236 ( .A1(n12349), .A2(n12348), .ZN(n12347) );
  NAND2_X2 U7237 ( .A1(n7372), .A2(n7370), .ZN(n12349) );
  OAI21_X2 U7238 ( .B1(n11969), .B2(n9107), .A(n9106), .ZN(n11886) );
  NAND2_X2 U7239 ( .A1(n9105), .A2(n9104), .ZN(n11969) );
  OAI22_X2 U7240 ( .A1(n7699), .A2(n7004), .B1(n7697), .B2(n9938), .ZN(n7629)
         );
  NAND2_X2 U7241 ( .A1(n7627), .A2(n7626), .ZN(n7699) );
  OAI211_X2 U7242 ( .C1(n12973), .C2(n6670), .A(n7157), .B(n6669), .ZN(n12916)
         );
  BUF_X4 U7243 ( .A(n6452), .Z(n6435) );
  OR2_X2 U7245 ( .A1(n14327), .A2(n14328), .ZN(n7072) );
  OAI21_X2 U7246 ( .B1(n14082), .B2(n14081), .A(n14322), .ZN(n14327) );
  NAND2_X1 U7247 ( .A1(n8351), .A2(n12524), .ZN(n8781) );
  XNOR2_X2 U7248 ( .A(n8131), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8193) );
  XNOR2_X2 U7249 ( .A(n9412), .B(P1_IR_REG_24__SCAN_IN), .ZN(n11240) );
  OAI211_X2 U7250 ( .C1(n14746), .C2(n6448), .A(n8390), .B(n8389), .ZN(n10124)
         );
  XNOR2_X2 U7251 ( .A(n8349), .B(n12518), .ZN(n11825) );
  XOR2_X2 U7252 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(n14040), .Z(n14041) );
  XNOR2_X2 U7253 ( .A(n14004), .B(n7077), .ZN(n14040) );
  AND2_X2 U7254 ( .A1(n11434), .A2(n9610), .ZN(n11446) );
  XNOR2_X1 U7256 ( .A(n8322), .B(n8321), .ZN(n6437) );
  INV_X8 U7257 ( .A(n12168), .ZN(n14738) );
  NOR2_X2 U7258 ( .A1(n11094), .A2(n6763), .ZN(n12006) );
  NOR2_X2 U7259 ( .A1(n14324), .A2(n14323), .ZN(n14082) );
  OAI21_X2 U7260 ( .B1(n14078), .B2(n14077), .A(n14318), .ZN(n14324) );
  AOI22_X2 U7261 ( .A1(P3_REG2_REG_2__SCAN_IN), .A2(n10839), .B1(n10892), .B2(
        n10317), .ZN(n10305) );
  OR2_X2 U7262 ( .A1(n8376), .A2(n7027), .ZN(n8378) );
  NAND2_X1 U7263 ( .A1(n7244), .A2(n7238), .ZN(n7242) );
  AND2_X1 U7264 ( .A1(n7006), .A2(n11690), .ZN(n13719) );
  NAND2_X1 U7265 ( .A1(n11676), .A2(n11675), .ZN(n13648) );
  AND2_X1 U7266 ( .A1(n8012), .A2(n8011), .ZN(n12954) );
  NAND2_X1 U7267 ( .A1(n11039), .A2(n11038), .ZN(n11175) );
  OAI21_X1 U7268 ( .B1(n14222), .B2(n6645), .A(n6643), .ZN(n14195) );
  AND2_X1 U7269 ( .A1(n10601), .A2(n10545), .ZN(n10559) );
  NAND2_X1 U7270 ( .A1(n10670), .A2(n10671), .ZN(n10768) );
  AOI21_X1 U7271 ( .B1(n10323), .B2(n10322), .A(n10321), .ZN(n14760) );
  NAND2_X1 U7272 ( .A1(n6749), .A2(n6748), .ZN(n14405) );
  INV_X2 U7273 ( .A(n10707), .ZN(n11994) );
  AND4_X1 U7274 ( .A1(n8427), .A2(n8426), .A3(n8425), .A4(n8424), .ZN(n10707)
         );
  INV_X1 U7275 ( .A(n13482), .ZN(n14383) );
  INV_X4 U7276 ( .A(n13364), .ZN(n13331) );
  INV_X2 U7277 ( .A(n13485), .ZN(n10215) );
  INV_X2 U7278 ( .A(n8968), .ZN(n12168) );
  BUF_X2 U7279 ( .A(n10107), .Z(n11744) );
  AND2_X1 U7280 ( .A1(n11446), .A2(n10095), .ZN(n13206) );
  BUF_X2 U7281 ( .A(n7778), .Z(n9338) );
  INV_X1 U7282 ( .A(n13822), .ZN(n14414) );
  INV_X2 U7283 ( .A(n9454), .ZN(n7942) );
  NOR2_X1 U7284 ( .A1(n7731), .A2(n7642), .ZN(n7653) );
  INV_X2 U7285 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7027) );
  OR2_X1 U7286 ( .A1(n9183), .A2(n14987), .ZN(n9057) );
  NAND2_X1 U7287 ( .A1(n9141), .A2(n11874), .ZN(n11876) );
  AOI21_X1 U7288 ( .B1(n6717), .B2(n9359), .A(n9358), .ZN(n9387) );
  NAND2_X1 U7289 ( .A1(n13894), .A2(n14429), .ZN(n7231) );
  AND2_X1 U7290 ( .A1(n13696), .A2(n13695), .ZN(n13904) );
  AOI21_X1 U7291 ( .B1(n13711), .B2(n13710), .A(n14540), .ZN(n13713) );
  XNOR2_X1 U7292 ( .A(n6744), .B(n13672), .ZN(n13894) );
  AND2_X1 U7293 ( .A1(n11833), .A2(n12282), .ZN(n11902) );
  AND2_X1 U7294 ( .A1(n6845), .A2(n11899), .ZN(n11833) );
  OR3_X2 U7295 ( .A1(n13727), .A2(n13721), .A3(n13709), .ZN(n13710) );
  AOI211_X1 U7296 ( .C1(n14538), .C2(n13919), .A(n13918), .B(n13917), .ZN(
        n13923) );
  OR2_X1 U7297 ( .A1(n12862), .A2(n14655), .ZN(n6795) );
  NAND2_X1 U7298 ( .A1(n13459), .A2(n13460), .ZN(n13458) );
  OAI21_X1 U7299 ( .B1(n6844), .B2(n13736), .A(n14429), .ZN(n6843) );
  AOI21_X1 U7300 ( .B1(n13771), .B2(n13757), .A(n13756), .ZN(n13760) );
  NAND2_X1 U7301 ( .A1(n13399), .A2(n13327), .ZN(n13459) );
  NOR2_X1 U7302 ( .A1(n13673), .A2(n13626), .ZN(n13621) );
  OAI21_X1 U7303 ( .B1(n12655), .B2(n6702), .A(n6699), .ZN(n6703) );
  NAND2_X1 U7304 ( .A1(n11746), .A2(n11745), .ZN(n13881) );
  NAND2_X1 U7305 ( .A1(n13326), .A2(n13397), .ZN(n13399) );
  INV_X1 U7306 ( .A(n13094), .ZN(n12856) );
  AOI21_X1 U7307 ( .B1(n6862), .B2(n14874), .A(n6859), .ZN(n6858) );
  AND2_X1 U7308 ( .A1(n9340), .A2(n9339), .ZN(n13094) );
  NAND2_X1 U7309 ( .A1(n13752), .A2(n7212), .ZN(n13921) );
  NAND2_X1 U7310 ( .A1(n7242), .A2(n7246), .ZN(n13773) );
  INV_X1 U7311 ( .A(n9132), .ZN(n6591) );
  INV_X1 U7312 ( .A(n7242), .ZN(n6439) );
  XNOR2_X1 U7313 ( .A(n9302), .B(n9301), .ZN(n13187) );
  NAND2_X1 U7314 ( .A1(n9336), .A2(n9299), .ZN(n9302) );
  NAND2_X1 U7315 ( .A1(n9336), .A2(n9335), .ZN(n13981) );
  OAI21_X1 U7316 ( .B1(n13346), .B2(n6633), .A(n6630), .ZN(n6634) );
  NAND2_X1 U7317 ( .A1(n11842), .A2(n11841), .ZN(n11910) );
  OR2_X1 U7318 ( .A1(n9334), .A2(n9333), .ZN(n9336) );
  INV_X1 U7319 ( .A(n6989), .ZN(n6986) );
  AND2_X1 U7320 ( .A1(n7058), .A2(n7057), .ZN(n14135) );
  NAND2_X1 U7321 ( .A1(n8287), .A2(n6592), .ZN(n8715) );
  OAI21_X1 U7322 ( .B1(n13010), .B2(n8186), .A(n8187), .ZN(n12992) );
  OR2_X1 U7323 ( .A1(n6593), .A2(n15122), .ZN(n8287) );
  OR2_X1 U7324 ( .A1(n14339), .A2(n14340), .ZN(n7057) );
  OAI21_X1 U7325 ( .B1(n8096), .B2(n8095), .A(n8098), .ZN(n8118) );
  NAND2_X1 U7326 ( .A1(n12082), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12109) );
  NAND2_X1 U7327 ( .A1(n8675), .A2(n8674), .ZN(n12432) );
  NAND2_X1 U7328 ( .A1(n7195), .A2(n7198), .ZN(n13828) );
  NAND2_X1 U7329 ( .A1(n11663), .A2(n11662), .ZN(n13919) );
  XNOR2_X1 U7330 ( .A(n12108), .B(n12087), .ZN(n12082) );
  AND2_X1 U7331 ( .A1(n8055), .A2(n8054), .ZN(n12923) );
  OAI21_X1 U7332 ( .B1(n8673), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n6595), .ZN(
        n8685) );
  NAND2_X1 U7333 ( .A1(n11629), .A2(n11628), .ZN(n13780) );
  OAI21_X1 U7334 ( .B1(n14231), .B2(n6642), .A(n6639), .ZN(n13258) );
  NAND2_X1 U7335 ( .A1(n6973), .A2(n6804), .ZN(n14242) );
  NAND2_X1 U7336 ( .A1(n6595), .A2(n6594), .ZN(n8673) );
  XNOR2_X1 U7337 ( .A(n8063), .B(n8062), .ZN(n11661) );
  AND3_X1 U7338 ( .A1(n7140), .A2(n7138), .A3(n7137), .ZN(n12103) );
  OR2_X1 U7339 ( .A1(n6596), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6594) );
  XNOR2_X1 U7340 ( .A(n13249), .B(n13247), .ZN(n14231) );
  AND2_X1 U7341 ( .A1(n7999), .A2(n7998), .ZN(n13129) );
  XNOR2_X1 U7342 ( .A(n7981), .B(n7980), .ZN(n11597) );
  INV_X1 U7343 ( .A(n12079), .ZN(n6440) );
  NAND2_X1 U7344 ( .A1(n7967), .A2(n7966), .ZN(n13142) );
  NAND2_X1 U7345 ( .A1(n7979), .A2(n7978), .ZN(n7981) );
  INV_X1 U7346 ( .A(n13069), .ZN(n6441) );
  OAI21_X2 U7347 ( .B1(n7993), .B2(n7005), .A(n7997), .ZN(n8027) );
  INV_X1 U7348 ( .A(n11233), .ZN(n6442) );
  NAND2_X1 U7349 ( .A1(n11080), .A2(n6776), .ZN(n11283) );
  AND2_X2 U7350 ( .A1(n7658), .A2(n7657), .ZN(n13022) );
  OR2_X1 U7351 ( .A1(n14237), .A2(n14208), .ZN(n13655) );
  NAND2_X1 U7352 ( .A1(n14219), .A2(n13217), .ZN(n14222) );
  NAND2_X1 U7353 ( .A1(n11221), .A2(n11220), .ZN(n14237) );
  NAND2_X1 U7354 ( .A1(n7735), .A2(n7734), .ZN(n13167) );
  NAND2_X1 U7355 ( .A1(n8616), .A2(n8270), .ZN(n8633) );
  NAND2_X1 U7356 ( .A1(n6914), .A2(n6912), .ZN(n7965) );
  NAND2_X1 U7357 ( .A1(n10768), .A2(n6672), .ZN(n10771) );
  XNOR2_X1 U7358 ( .A(n6740), .B(n7729), .ZN(n11219) );
  NAND2_X1 U7359 ( .A1(n8614), .A2(n8613), .ZN(n8616) );
  NAND2_X1 U7360 ( .A1(n10970), .A2(n11314), .ZN(n11211) );
  NAND2_X1 U7361 ( .A1(n11179), .A2(n11178), .ZN(n14285) );
  OR2_X1 U7362 ( .A1(n7681), .A2(n7237), .ZN(n6914) );
  XNOR2_X1 U7363 ( .A(n7746), .B(n7745), .ZN(n11176) );
  NAND2_X1 U7364 ( .A1(n8452), .A2(n8798), .ZN(n10946) );
  AOI21_X1 U7365 ( .B1(n6455), .B2(n7449), .A(n7448), .ZN(n7447) );
  OAI21_X1 U7366 ( .B1(n7165), .B2(n14858), .A(n7164), .ZN(n11094) );
  NAND2_X1 U7367 ( .A1(n8585), .A2(n8584), .ZN(n8587) );
  NAND2_X1 U7368 ( .A1(n6803), .A2(n6802), .ZN(n10750) );
  NAND2_X1 U7369 ( .A1(n14850), .A2(n6849), .ZN(n10846) );
  INV_X1 U7370 ( .A(n11091), .ZN(n14716) );
  NOR2_X1 U7371 ( .A1(n14841), .A2(n14840), .ZN(n14839) );
  NOR2_X1 U7372 ( .A1(n14819), .A2(n10902), .ZN(n14841) );
  OR2_X1 U7373 ( .A1(n10269), .A2(n9337), .ZN(n7852) );
  NAND2_X1 U7374 ( .A1(n8561), .A2(n8560), .ZN(n8563) );
  NAND2_X1 U7375 ( .A1(n7882), .A2(n7608), .ZN(n7610) );
  NAND2_X2 U7376 ( .A1(n10371), .A2(n12998), .ZN(n13038) );
  XNOR2_X1 U7377 ( .A(n10901), .B(n14829), .ZN(n14820) );
  NAND2_X1 U7378 ( .A1(n7013), .A2(n10383), .ZN(n10429) );
  AND3_X1 U7379 ( .A1(n7152), .A2(n7151), .A3(n6561), .ZN(n10901) );
  NAND2_X1 U7380 ( .A1(n8544), .A2(n8543), .ZN(n8546) );
  NAND2_X1 U7381 ( .A1(n7810), .A2(n7148), .ZN(n14659) );
  INV_X1 U7382 ( .A(n10947), .ZN(n14888) );
  OR2_X1 U7383 ( .A1(n14786), .A2(n7153), .ZN(n7152) );
  AND4_X1 U7384 ( .A1(n8410), .A2(n8409), .A3(n8408), .A4(n8407), .ZN(n14902)
         );
  AND2_X2 U7385 ( .A1(n13679), .A2(n14416), .ZN(n14439) );
  NAND2_X1 U7386 ( .A1(n7143), .A2(n7142), .ZN(n14768) );
  CLKBUF_X3 U7387 ( .A(n8421), .Z(n8756) );
  BUF_X2 U7388 ( .A(n8400), .Z(n8617) );
  BUF_X2 U7389 ( .A(n8411), .Z(n6787) );
  NAND2_X1 U7390 ( .A1(n6447), .A2(n9657), .ZN(n8411) );
  NAND4_X1 U7391 ( .A1(n10239), .A2(n10238), .A3(n10237), .A4(n10236), .ZN(
        n13482) );
  NAND2_X1 U7392 ( .A1(n9028), .A2(n9027), .ZN(n9147) );
  OR2_X1 U7393 ( .A1(n14752), .A2(n7144), .ZN(n7143) );
  NAND2_X1 U7394 ( .A1(n7020), .A2(n14054), .ZN(n14057) );
  XNOR2_X1 U7395 ( .A(n10893), .B(n14765), .ZN(n14752) );
  AND4_X1 U7396 ( .A1(n9710), .A2(n9709), .A3(n9708), .A4(n9707), .ZN(n10221)
         );
  CLKBUF_X1 U7397 ( .A(n8969), .Z(n12531) );
  NAND3_X1 U7398 ( .A1(n7788), .A2(n7789), .A3(n6489), .ZN(n12743) );
  AND2_X1 U7399 ( .A1(n9060), .A2(n9059), .ZN(n9061) );
  NAND2_X2 U7400 ( .A1(n8347), .A2(n12517), .ZN(n12524) );
  XNOR2_X1 U7401 ( .A(n10804), .B(P3_B_REG_SCAN_IN), .ZN(n9025) );
  INV_X1 U7402 ( .A(n13367), .ZN(n6444) );
  NOR2_X1 U7403 ( .A1(n10306), .A2(n10305), .ZN(n10891) );
  NAND4_X1 U7404 ( .A1(n7767), .A2(n7766), .A3(n7764), .A4(n7765), .ZN(n12746)
         );
  OR2_X2 U7405 ( .A1(n11446), .A2(n9586), .ZN(n13365) );
  NAND2_X1 U7406 ( .A1(n12177), .A2(n10169), .ZN(n9060) );
  MUX2_X1 U7407 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8345), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8347) );
  NOR2_X1 U7408 ( .A1(n8316), .A2(n8315), .ZN(n8319) );
  OR2_X1 U7409 ( .A1(n8317), .A2(n7027), .ZN(n8318) );
  NAND2_X1 U7410 ( .A1(n8959), .A2(n8958), .ZN(n10804) );
  NAND2_X1 U7411 ( .A1(n8320), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8322) );
  AND2_X1 U7412 ( .A1(n8313), .A2(n7438), .ZN(n8317) );
  NAND2_X1 U7413 ( .A1(n7078), .A2(n14003), .ZN(n14004) );
  NAND2_X1 U7414 ( .A1(n8415), .A2(n8244), .ZN(n8429) );
  NOR2_X1 U7415 ( .A1(n10138), .A2(n14932), .ZN(n10303) );
  NAND2_X1 U7416 ( .A1(n9575), .A2(n7296), .ZN(n13822) );
  MUX2_X1 U7417 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9536), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n9538) );
  XNOR2_X1 U7418 ( .A(n9553), .B(n6902), .ZN(n13979) );
  INV_X2 U7419 ( .A(n12515), .ZN(n12528) );
  NAND2_X1 U7420 ( .A1(n9575), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9568) );
  OAI21_X1 U7421 ( .B1(n7218), .B2(SI_3_), .A(n7591), .ZN(n7217) );
  NAND2_X1 U7422 ( .A1(n8135), .A2(n8134), .ZN(n10942) );
  AND2_X2 U7423 ( .A1(n8311), .A2(n8310), .ZN(n8313) );
  NAND2_X2 U7424 ( .A1(n7012), .A2(P1_U3086), .ZN(n13986) );
  NAND2_X1 U7425 ( .A1(n8413), .A2(n8412), .ZN(n8415) );
  NAND2_X1 U7426 ( .A1(n13974), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9553) );
  NOR2_X1 U7427 ( .A1(n8618), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n8621) );
  XNOR2_X1 U7428 ( .A(n8140), .B(n8139), .ZN(n8194) );
  XNOR2_X1 U7429 ( .A(n9572), .B(n15080), .ZN(n11433) );
  NAND2_X1 U7430 ( .A1(n9554), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9556) );
  INV_X1 U7431 ( .A(n8956), .ZN(n8311) );
  MUX2_X1 U7432 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8133), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n8135) );
  INV_X1 U7433 ( .A(n6627), .ZN(n9412) );
  NAND2_X2 U7434 ( .A1(n9657), .A2(P1_U3086), .ZN(n13988) );
  MUX2_X1 U7435 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9540), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n9541) );
  NAND2_X1 U7436 ( .A1(n9574), .A2(n9573), .ZN(n9575) );
  NAND2_X2 U7437 ( .A1(n9657), .A2(P2_U3088), .ZN(n13199) );
  NAND2_X1 U7438 ( .A1(n8134), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8131) );
  NAND2_X1 U7439 ( .A1(n6724), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7673) );
  NAND2_X1 U7440 ( .A1(n9571), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9574) );
  OR2_X1 U7441 ( .A1(n6624), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n8618) );
  OAI21_X1 U7442 ( .B1(n9571), .B2(n9570), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9572) );
  NOR2_X1 U7443 ( .A1(n9576), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U7444 ( .A1(n7655), .A2(n7297), .ZN(n8134) );
  AND3_X1 U7445 ( .A1(n7200), .A2(n7199), .A3(n6560), .ZN(n9552) );
  AND2_X1 U7446 ( .A1(n7567), .A2(n7653), .ZN(n7655) );
  AND2_X1 U7447 ( .A1(n7730), .A2(n7653), .ZN(n6725) );
  AND3_X1 U7448 ( .A1(n7573), .A2(n6930), .A3(n9415), .ZN(n7199) );
  AND3_X1 U7449 ( .A1(n9408), .A2(n9407), .A3(n7294), .ZN(n10174) );
  INV_X1 U7450 ( .A(n9414), .ZN(n9415) );
  NAND2_X1 U7451 ( .A1(n7649), .A2(n7539), .ZN(n7808) );
  AND4_X1 U7452 ( .A1(n8301), .A2(n8300), .A3(n8492), .A4(n8478), .ZN(n8302)
         );
  AND4_X1 U7453 ( .A1(n9406), .A2(n9404), .A3(n9405), .A4(n9653), .ZN(n9407)
         );
  AND4_X1 U7454 ( .A1(n6947), .A2(n6948), .A3(n6949), .A4(n9577), .ZN(n7573)
         );
  AND2_X1 U7455 ( .A1(n7352), .A2(n7351), .ZN(n6620) );
  INV_X4 U7456 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7457 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8310) );
  INV_X1 U7458 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7732) );
  INV_X1 U7459 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8208) );
  INV_X1 U7460 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7578) );
  NOR2_X1 U7461 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n7293) );
  INV_X1 U7462 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8222) );
  INV_X1 U7463 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6902) );
  NOR2_X1 U7464 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n6948) );
  NOR2_X1 U7465 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n6949) );
  INV_X4 U7466 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X2 U7467 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7649) );
  NOR2_X1 U7468 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9815) );
  INV_X1 U7469 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8478) );
  NOR2_X1 U7470 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8301) );
  NOR2_X1 U7471 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n8300) );
  NOR2_X1 U7472 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n9405) );
  NOR2_X1 U7473 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7636) );
  NOR2_X1 U7474 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n9404) );
  NOR2_X1 U7475 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7637) );
  NAND2_X1 U7476 ( .A1(n11825), .A2(n12524), .ZN(n6446) );
  NAND2_X2 U7477 ( .A1(n11825), .A2(n12524), .ZN(n8653) );
  NAND2_X1 U7478 ( .A1(n12205), .A2(n8774), .ZN(n8975) );
  NAND4_X4 U7479 ( .A1(n8386), .A2(n8385), .A3(n8384), .A4(n8383), .ZN(n14918)
         );
  AND2_X2 U7480 ( .A1(n10942), .A2(n8193), .ZN(n9186) );
  NOR2_X2 U7481 ( .A1(n14070), .A2(n14071), .ZN(n14074) );
  NAND2_X1 U7482 ( .A1(n6437), .A2(n8969), .ZN(n6448) );
  NAND2_X1 U7483 ( .A1(n14738), .A2(n8969), .ZN(n10134) );
  BUF_X4 U7484 ( .A(n8405), .Z(n6450) );
  AND2_X2 U7485 ( .A1(n11825), .A2(n8350), .ZN(n8405) );
  OAI222_X1 U7486 ( .A1(P3_U3151), .A2(n11825), .B1(n12521), .B2(n11824), .C1(
        n12528), .C2(n11823), .ZN(P3_U3265) );
  NOR2_X2 U7487 ( .A1(n11106), .A2(n11105), .ZN(n12001) );
  NOR2_X2 U7488 ( .A1(n12934), .A2(n13113), .ZN(n12920) );
  AND2_X1 U7489 ( .A1(n11612), .A2(n11609), .ZN(n10107) );
  NAND2_X2 U7490 ( .A1(n12253), .A2(n8897), .ZN(n12240) );
  OAI22_X2 U7491 ( .A1(n14242), .A2(n14249), .B1(n13657), .B2(n13866), .ZN(
        n13869) );
  OR2_X1 U7493 ( .A1(n11446), .A2(n9858), .ZN(n13367) );
  AOI21_X2 U7494 ( .B1(n9025), .B2(n11016), .A(n11201), .ZN(n11424) );
  NAND2_X1 U7495 ( .A1(n9192), .A2(n9191), .ZN(n6704) );
  INV_X1 U7496 ( .A(n9237), .ZN(n6731) );
  OAI22_X1 U7497 ( .A1(n14716), .A2(n9342), .B1(n11288), .B2(n9213), .ZN(n9237) );
  INV_X1 U7498 ( .A(n12524), .ZN(n8350) );
  AND2_X1 U7499 ( .A1(n8997), .A2(n7368), .ZN(n7367) );
  OR2_X1 U7500 ( .A1(n11353), .A2(n7369), .ZN(n7368) );
  OAI21_X1 U7501 ( .B1(n12900), .B2(n8078), .A(n9360), .ZN(n12885) );
  NAND2_X1 U7502 ( .A1(n8081), .A2(n8082), .ZN(n8096) );
  NAND2_X1 U7503 ( .A1(n8080), .A2(n11200), .ZN(n8081) );
  NAND2_X1 U7504 ( .A1(n11298), .A2(n9089), .ZN(n11364) );
  INV_X1 U7505 ( .A(n8617), .ZN(n8778) );
  AND4_X1 U7506 ( .A1(n11706), .A2(n11705), .A3(n11704), .A4(n11703), .ZN(
        n13675) );
  NAND2_X1 U7507 ( .A1(n7170), .A2(n6921), .ZN(n13703) );
  NAND2_X1 U7508 ( .A1(n7174), .A2(n7171), .ZN(n7170) );
  NAND2_X1 U7509 ( .A1(n13726), .A2(n6922), .ZN(n6921) );
  INV_X1 U7510 ( .A(n7175), .ZN(n7171) );
  INV_X1 U7511 ( .A(n13626), .ZN(n13887) );
  NAND2_X1 U7512 ( .A1(n6736), .A2(n6762), .ZN(n6735) );
  OAI22_X1 U7513 ( .A1(n10431), .A2(n6445), .B1(n10090), .B2(n9342), .ZN(n9212) );
  AND2_X1 U7514 ( .A1(n7485), .A2(n9214), .ZN(n6779) );
  NAND2_X1 U7515 ( .A1(n7484), .A2(n7483), .ZN(n7487) );
  AOI21_X1 U7516 ( .B1(n7523), .B2(n9244), .A(n7522), .ZN(n7521) );
  INV_X1 U7517 ( .A(n9242), .ZN(n7522) );
  NAND2_X1 U7518 ( .A1(n9235), .A2(n6730), .ZN(n6728) );
  INV_X1 U7519 ( .A(n9236), .ZN(n6729) );
  NAND2_X1 U7520 ( .A1(n6731), .A2(n9238), .ZN(n6730) );
  INV_X1 U7521 ( .A(n9287), .ZN(n6720) );
  INV_X1 U7522 ( .A(n9288), .ZN(n6716) );
  AOI21_X1 U7523 ( .B1(n6476), .B2(n11720), .A(n6882), .ZN(n6881) );
  INV_X1 U7524 ( .A(n11722), .ZN(n6882) );
  OAI21_X1 U7525 ( .B1(n6990), .B2(n13772), .A(n13669), .ZN(n6989) );
  NAND2_X1 U7526 ( .A1(n7965), .A2(n7964), .ZN(n7993) );
  NAND2_X1 U7527 ( .A1(n14050), .A2(n14051), .ZN(n7078) );
  NOR2_X1 U7528 ( .A1(n8908), .A2(n8909), .ZN(n9015) );
  OR2_X1 U7529 ( .A1(n8678), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8688) );
  INV_X1 U7530 ( .A(n10198), .ZN(n9047) );
  AND2_X1 U7531 ( .A1(n9381), .A2(n9316), .ZN(n9349) );
  OR2_X1 U7532 ( .A1(n13096), .A2(n12602), .ZN(n8116) );
  OR2_X1 U7533 ( .A1(n13108), .A2(n12629), .ZN(n9361) );
  NAND2_X1 U7534 ( .A1(n13124), .A2(n12675), .ZN(n7162) );
  OR2_X1 U7535 ( .A1(n7984), .A2(n12620), .ZN(n8001) );
  INV_X1 U7536 ( .A(n12736), .ZN(n10787) );
  AND2_X1 U7537 ( .A1(n10718), .A2(n8164), .ZN(n7514) );
  NAND2_X1 U7538 ( .A1(n10436), .A2(n10437), .ZN(n7843) );
  OAI21_X1 U7539 ( .B1(n10422), .B2(n7544), .A(n8159), .ZN(n7543) );
  AND2_X1 U7540 ( .A1(n8194), .A2(n10418), .ZN(n9343) );
  NAND2_X1 U7541 ( .A1(n6798), .A2(n6796), .ZN(n9393) );
  NOR2_X1 U7542 ( .A1(n7671), .A2(n6797), .ZN(n6796) );
  NAND2_X1 U7543 ( .A1(n7648), .A2(n6470), .ZN(n6798) );
  NOR2_X1 U7544 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n6797) );
  OR2_X1 U7545 ( .A1(n7868), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7884) );
  INV_X1 U7546 ( .A(n9558), .ZN(n9557) );
  NAND2_X1 U7547 ( .A1(n13719), .A2(n13651), .ZN(n7174) );
  INV_X1 U7548 ( .A(n7248), .ZN(n7243) );
  OR2_X1 U7549 ( .A1(n14285), .A2(n13236), .ZN(n11508) );
  INV_X1 U7550 ( .A(n11431), .ZN(n9586) );
  NAND2_X1 U7551 ( .A1(n6998), .A2(n8064), .ZN(n8080) );
  INV_X1 U7552 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9577) );
  AND2_X1 U7553 ( .A1(n6906), .A2(n7254), .ZN(n6905) );
  AOI21_X1 U7554 ( .B1(n7257), .B2(n7259), .A(n7255), .ZN(n7254) );
  XNOR2_X1 U7555 ( .A(n7726), .B(SI_14_), .ZN(n7746) );
  OAI21_X1 U7556 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14017), .A(n14016), .ZN(
        n14072) );
  AOI22_X1 U7557 ( .A1(n7048), .A2(n9144), .B1(n7047), .B2(n7045), .ZN(n7044)
         );
  INV_X1 U7558 ( .A(n11962), .ZN(n7045) );
  AOI21_X1 U7559 ( .B1(n7051), .B2(n7054), .A(n6612), .ZN(n6611) );
  INV_X1 U7560 ( .A(n11951), .ZN(n6612) );
  AOI21_X1 U7561 ( .B1(n11910), .B2(n9123), .A(n7569), .ZN(n11851) );
  NAND2_X1 U7562 ( .A1(n11165), .A2(n6510), .ZN(n11298) );
  NAND2_X1 U7563 ( .A1(n7062), .A2(n12294), .ZN(n7061) );
  NAND2_X1 U7564 ( .A1(n11365), .A2(n9092), .ZN(n11861) );
  NAND2_X1 U7565 ( .A1(n7066), .A2(n9067), .ZN(n7065) );
  NOR2_X1 U7566 ( .A1(n8927), .A2(n8788), .ZN(n7399) );
  OR2_X1 U7567 ( .A1(n8925), .A2(n6556), .ZN(n7398) );
  NAND2_X1 U7568 ( .A1(n8975), .A2(n8919), .ZN(n7400) );
  AND4_X1 U7569 ( .A1(n8559), .A2(n8558), .A3(n8557), .A4(n8556), .ZN(n11937)
         );
  INV_X1 U7570 ( .A(n6436), .ZN(n8769) );
  AND2_X1 U7571 ( .A1(n8351), .A2(n8350), .ZN(n8421) );
  NAND2_X1 U7572 ( .A1(n14852), .A2(n14851), .ZN(n14850) );
  XNOR2_X1 U7573 ( .A(n10846), .B(n10905), .ZN(n14873) );
  OR2_X1 U7574 ( .A1(n11883), .A2(n12249), .ZN(n7568) );
  NAND2_X1 U7575 ( .A1(n8903), .A2(n8736), .ZN(n12239) );
  NAND2_X1 U7576 ( .A1(n7419), .A2(n7427), .ZN(n7418) );
  AND2_X1 U7577 ( .A1(n7427), .A2(n7425), .ZN(n7420) );
  NAND2_X1 U7578 ( .A1(n12286), .A2(n12294), .ZN(n8888) );
  NAND2_X1 U7579 ( .A1(n7382), .A2(n6516), .ZN(n12308) );
  XNOR2_X1 U7580 ( .A(n12432), .B(n12295), .ZN(n12311) );
  AOI21_X1 U7581 ( .B1(n7367), .B2(n7369), .A(n6567), .ZN(n7365) );
  AOI21_X1 U7582 ( .B1(n7362), .B2(n7364), .A(n7360), .ZN(n7359) );
  INV_X1 U7583 ( .A(n8852), .ZN(n7360) );
  OAI21_X1 U7584 ( .B1(n10949), .B2(n7402), .A(n7401), .ZN(n11248) );
  AOI21_X1 U7585 ( .B1(n7403), .B2(n7408), .A(n6465), .ZN(n7401) );
  INV_X1 U7586 ( .A(n7403), .ZN(n7402) );
  NAND2_X1 U7587 ( .A1(n7405), .A2(n7406), .ZN(n11154) );
  AOI21_X1 U7588 ( .B1(n7379), .B2(n7381), .A(n7377), .ZN(n7376) );
  INV_X1 U7589 ( .A(n8827), .ZN(n7377) );
  AND2_X1 U7590 ( .A1(n9020), .A2(n9019), .ZN(n14891) );
  AND2_X1 U7591 ( .A1(n9162), .A2(n10132), .ZN(n14919) );
  NAND2_X1 U7592 ( .A1(n8740), .A2(n8739), .ZN(n11959) );
  OR2_X1 U7593 ( .A1(n6787), .A2(n11200), .ZN(n8739) );
  INV_X1 U7594 ( .A(n6787), .ZN(n8663) );
  INV_X1 U7595 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8312) );
  OR2_X1 U7596 ( .A1(n8474), .A2(n8473), .ZN(n8476) );
  INV_X1 U7597 ( .A(n7340), .ZN(n7339) );
  OAI21_X1 U7598 ( .B1(n7343), .B2(n7344), .A(n7341), .ZN(n7340) );
  NAND2_X1 U7599 ( .A1(n7346), .A2(n7342), .ZN(n7341) );
  INV_X1 U7600 ( .A(n12599), .ZN(n7342) );
  NAND2_X1 U7601 ( .A1(n10084), .A2(n7303), .ZN(n7302) );
  INV_X1 U7602 ( .A(n7763), .ZN(n8122) );
  AND4_X1 U7604 ( .A1(n7878), .A2(n7877), .A3(n7876), .A4(n7875), .ZN(n10741)
         );
  AND2_X1 U7605 ( .A1(n6815), .A2(n11426), .ZN(n8056) );
  AND2_X1 U7606 ( .A1(n11426), .A2(n11429), .ZN(n7769) );
  NAND2_X1 U7607 ( .A1(n7495), .A2(n7503), .ZN(n7494) );
  AOI21_X1 U7608 ( .B1(n7495), .B2(n7493), .A(n6535), .ZN(n7492) );
  XNOR2_X1 U7609 ( .A(n13103), .B(n12727), .ZN(n12884) );
  AOI21_X1 U7610 ( .B1(n12916), .B2(n12915), .A(n6531), .ZN(n12900) );
  AOI21_X1 U7611 ( .B1(n7532), .B2(n7531), .A(n9374), .ZN(n7528) );
  INV_X1 U7612 ( .A(n13002), .ZN(n13055) );
  AND2_X1 U7613 ( .A1(n9454), .A2(n7012), .ZN(n7778) );
  NAND2_X1 U7614 ( .A1(n8142), .A2(n8141), .ZN(n13065) );
  NAND2_X2 U7615 ( .A1(n6739), .A2(n10583), .ZN(n14689) );
  XNOR2_X1 U7616 ( .A(n9186), .B(n8194), .ZN(n6739) );
  OR2_X1 U7617 ( .A1(n7671), .A2(n13189), .ZN(n7647) );
  INV_X1 U7618 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8215) );
  INV_X1 U7619 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8212) );
  INV_X1 U7620 ( .A(n7474), .ZN(n7473) );
  OAI21_X1 U7621 ( .B1(n7476), .B2(n7475), .A(n13442), .ZN(n7474) );
  AND2_X1 U7622 ( .A1(n13416), .A2(n13306), .ZN(n13345) );
  NOR2_X1 U7623 ( .A1(n13335), .A2(n13334), .ZN(n13336) );
  AND2_X1 U7624 ( .A1(n13337), .A2(n7457), .ZN(n7456) );
  OR2_X1 U7625 ( .A1(n13460), .A2(n13336), .ZN(n7457) );
  NAND2_X1 U7626 ( .A1(n13321), .A2(n13322), .ZN(n13327) );
  NAND2_X2 U7627 ( .A1(n6444), .A2(n14468), .ZN(n13364) );
  NAND2_X1 U7628 ( .A1(n7446), .A2(n6513), .ZN(n7445) );
  NAND2_X1 U7629 ( .A1(n11743), .A2(n9543), .ZN(n7446) );
  NAND3_X1 U7630 ( .A1(n7459), .A2(n7461), .A3(n7460), .ZN(n10488) );
  NAND2_X1 U7631 ( .A1(n6480), .A2(n10120), .ZN(n7460) );
  NAND2_X1 U7632 ( .A1(n10116), .A2(n6480), .ZN(n7461) );
  NAND2_X1 U7633 ( .A1(n7468), .A2(n13263), .ZN(n7466) );
  NAND2_X1 U7634 ( .A1(n14199), .A2(n13243), .ZN(n13249) );
  NAND2_X1 U7635 ( .A1(n9557), .A2(n13979), .ZN(n11730) );
  AND2_X1 U7636 ( .A1(n13652), .A2(n11754), .ZN(n13704) );
  AND2_X1 U7637 ( .A1(n11708), .A2(n11707), .ZN(n13700) );
  AND2_X1 U7638 ( .A1(n13728), .A2(n13719), .ZN(n13714) );
  NAND2_X1 U7639 ( .A1(n13921), .A2(n13647), .ZN(n13726) );
  INV_X1 U7640 ( .A(n13644), .ZN(n13756) );
  OR2_X1 U7641 ( .A1(n13945), .A2(n13817), .ZN(n7248) );
  AOI21_X1 U7642 ( .B1(n7210), .B2(n13663), .A(n6526), .ZN(n7208) );
  AND2_X1 U7643 ( .A1(n7204), .A2(n13631), .ZN(n7201) );
  NAND2_X1 U7644 ( .A1(n7203), .A2(n14249), .ZN(n7205) );
  AND2_X1 U7645 ( .A1(n6977), .A2(n6485), .ZN(n6976) );
  INV_X1 U7646 ( .A(n6981), .ZN(n6978) );
  INV_X1 U7647 ( .A(n6980), .ZN(n6979) );
  AOI21_X1 U7648 ( .B1(n11036), .B2(n6959), .A(n6525), .ZN(n6958) );
  INV_X1 U7649 ( .A(n10993), .ZN(n6959) );
  AOI21_X1 U7650 ( .B1(n7186), .B2(n11767), .A(n6523), .ZN(n7185) );
  INV_X1 U7651 ( .A(n14380), .ZN(n13835) );
  INV_X1 U7652 ( .A(n14382), .ZN(n13865) );
  INV_X1 U7653 ( .A(n13719), .ZN(n13906) );
  INV_X1 U7654 ( .A(n14528), .ZN(n14538) );
  OR2_X1 U7655 ( .A1(n14468), .A2(n13822), .ZN(n9915) );
  XNOR2_X1 U7656 ( .A(n8096), .B(n8084), .ZN(n13195) );
  XNOR2_X1 U7657 ( .A(n7909), .B(n7908), .ZN(n10995) );
  OAI21_X1 U7658 ( .B1(n7610), .B2(n7612), .A(n7251), .ZN(n7909) );
  NAND2_X1 U7659 ( .A1(n7830), .A2(n7600), .ZN(n7845) );
  NAND2_X1 U7660 ( .A1(n7845), .A2(n7844), .ZN(n7846) );
  INV_X1 U7661 ( .A(n9657), .ZN(n7012) );
  NAND2_X1 U7662 ( .A1(n8766), .A2(n8765), .ZN(n11819) );
  INV_X1 U7663 ( .A(n10931), .ZN(n6696) );
  NAND2_X1 U7664 ( .A1(n11725), .A2(n11724), .ZN(n13626) );
  OR2_X1 U7665 ( .A1(n13981), .A2(n11723), .ZN(n11725) );
  NAND2_X1 U7666 ( .A1(n13703), .A2(n13704), .ZN(n13896) );
  AOI22_X1 U7667 ( .A1(n12746), .A2(n9342), .B1(n10515), .B2(n6445), .ZN(n9188) );
  NAND2_X1 U7668 ( .A1(n6734), .A2(n6733), .ZN(n6732) );
  INV_X1 U7669 ( .A(n9196), .ZN(n6733) );
  INV_X1 U7670 ( .A(n6704), .ZN(n6734) );
  OAI22_X1 U7671 ( .A1(n11467), .A2(n6900), .B1(n11466), .B2(n6899), .ZN(
        n11470) );
  INV_X1 U7672 ( .A(n11465), .ZN(n6899) );
  NOR2_X1 U7673 ( .A1(n6901), .A2(n11465), .ZN(n6900) );
  NAND2_X1 U7674 ( .A1(n7285), .A2(n11476), .ZN(n7284) );
  NOR2_X1 U7675 ( .A1(n7486), .A2(n7483), .ZN(n7482) );
  AND2_X1 U7676 ( .A1(n6711), .A2(n6708), .ZN(n9229) );
  INV_X1 U7677 ( .A(n9228), .ZN(n6707) );
  NOR2_X1 U7678 ( .A1(n9225), .A2(n9228), .ZN(n6710) );
  AOI21_X1 U7679 ( .B1(n6897), .B2(n6896), .A(n6894), .ZN(n6893) );
  OR4_X1 U7680 ( .A1(n13636), .A2(n13864), .A3(n13860), .A4(n11719), .ZN(
        n11572) );
  AOI22_X1 U7681 ( .A1(n7520), .A2(n7525), .B1(n7524), .B2(n7521), .ZN(n7516)
         );
  OR2_X1 U7682 ( .A1(n7525), .A2(n9243), .ZN(n7524) );
  INV_X1 U7683 ( .A(n9255), .ZN(n7552) );
  AOI21_X1 U7684 ( .B1(n9253), .B2(n9252), .A(n6536), .ZN(n6723) );
  NAND2_X1 U7685 ( .A1(n6887), .A2(n11600), .ZN(n6886) );
  OR2_X1 U7686 ( .A1(n11614), .A2(n11613), .ZN(n11618) );
  NAND2_X1 U7687 ( .A1(n7286), .A2(n11631), .ZN(n7290) );
  NAND2_X1 U7688 ( .A1(n9271), .A2(n7555), .ZN(n7554) );
  AND2_X1 U7689 ( .A1(n9270), .A2(n9269), .ZN(n7556) );
  NOR2_X1 U7690 ( .A1(n6892), .A2(n11665), .ZN(n6890) );
  NAND2_X1 U7691 ( .A1(n11665), .A2(n6892), .ZN(n6891) );
  NAND2_X1 U7692 ( .A1(n7620), .A2(SI_15_), .ZN(n7622) );
  INV_X1 U7693 ( .A(n7908), .ZN(n7250) );
  NAND2_X1 U7694 ( .A1(n7553), .A2(n6679), .ZN(n6678) );
  INV_X1 U7695 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6679) );
  INV_X1 U7696 ( .A(n6881), .ZN(n6878) );
  INV_X1 U7697 ( .A(n13709), .ZN(n6813) );
  AND2_X1 U7698 ( .A1(n13756), .A2(n13757), .ZN(n7245) );
  NAND2_X1 U7699 ( .A1(n7247), .A2(n13772), .ZN(n7240) );
  NAND2_X1 U7700 ( .A1(n13995), .A2(n13822), .ZN(n11431) );
  NAND2_X1 U7701 ( .A1(n13485), .A2(n9925), .ZN(n10228) );
  NAND2_X1 U7702 ( .A1(n8034), .A2(n8033), .ZN(n8048) );
  NAND2_X1 U7703 ( .A1(n8027), .A2(n8026), .ZN(n8034) );
  NOR2_X1 U7704 ( .A1(n6913), .A2(n7962), .ZN(n6912) );
  INV_X1 U7705 ( .A(n7630), .ZN(n6913) );
  NAND2_X1 U7706 ( .A1(n7631), .A2(n10018), .ZN(n7964) );
  NOR2_X1 U7707 ( .A1(n7628), .A2(SI_17_), .ZN(n7004) );
  NOR3_X1 U7708 ( .A1(n11803), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n10307) );
  NOR2_X1 U7709 ( .A1(n10891), .A2(n6490), .ZN(n10893) );
  NAND2_X1 U7710 ( .A1(n14778), .A2(n6850), .ZN(n10842) );
  NAND2_X1 U7711 ( .A1(n14775), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n6850) );
  OR2_X1 U7712 ( .A1(n8767), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12184) );
  OR2_X1 U7713 ( .A1(n11819), .A2(n12214), .ZN(n8914) );
  AND2_X1 U7714 ( .A1(n11959), .A2(n12215), .ZN(n8909) );
  NOR2_X1 U7715 ( .A1(n11959), .A2(n12215), .ZN(n8908) );
  OR2_X1 U7716 ( .A1(n8741), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8754) );
  NOR2_X1 U7717 ( .A1(n9014), .A2(n7426), .ZN(n7425) );
  INV_X1 U7718 ( .A(n7566), .ZN(n7426) );
  NAND2_X1 U7719 ( .A1(n8338), .A2(n15079), .ZN(n8697) );
  INV_X1 U7720 ( .A(n8688), .ZN(n8338) );
  NOR2_X1 U7721 ( .A1(n12356), .A2(n7374), .ZN(n7373) );
  NOR2_X1 U7722 ( .A1(n12372), .A2(n7375), .ZN(n7374) );
  INV_X1 U7723 ( .A(n8861), .ZN(n7375) );
  OR2_X1 U7724 ( .A1(n8626), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8637) );
  NAND2_X1 U7725 ( .A1(n8333), .A2(n11973), .ZN(n8626) );
  INV_X1 U7726 ( .A(n8606), .ZN(n8333) );
  NAND2_X1 U7727 ( .A1(n8332), .A2(n11925), .ZN(n8591) );
  INV_X1 U7728 ( .A(n8577), .ZN(n8332) );
  INV_X1 U7729 ( .A(n8837), .ZN(n7411) );
  INV_X1 U7730 ( .A(n8841), .ZN(n7410) );
  NAND2_X1 U7731 ( .A1(n6537), .A2(n6453), .ZN(n7406) );
  NAND2_X1 U7732 ( .A1(n14921), .A2(n14910), .ZN(n8807) );
  NAND2_X1 U7733 ( .A1(n11246), .A2(n8994), .ZN(n11378) );
  NAND2_X1 U7734 ( .A1(n8312), .A2(n8321), .ZN(n7440) );
  AOI21_X1 U7735 ( .B1(n7099), .B2(n7097), .A(n6585), .ZN(n7096) );
  INV_X1 U7736 ( .A(n7099), .ZN(n7098) );
  NAND2_X1 U7737 ( .A1(n8563), .A2(n8263), .ZN(n8264) );
  NAND2_X1 U7738 ( .A1(n7084), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U7739 ( .A1(n9646), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8241) );
  NOR2_X1 U7740 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n8375) );
  XNOR2_X1 U7741 ( .A(n13022), .B(n12576), .ZN(n12547) );
  NOR2_X1 U7742 ( .A1(n9290), .A2(n9291), .ZN(n7479) );
  NAND2_X1 U7743 ( .A1(n7548), .A2(n7547), .ZN(n7546) );
  AND2_X1 U7744 ( .A1(n6563), .A2(n6714), .ZN(n6713) );
  NAND2_X1 U7745 ( .A1(n6720), .A2(n6716), .ZN(n6714) );
  NOR2_X1 U7746 ( .A1(n6720), .A2(n6716), .ZN(n6715) );
  AND2_X1 U7747 ( .A1(n9349), .A2(n9320), .ZN(n9328) );
  NAND2_X1 U7748 ( .A1(n9347), .A2(n9381), .ZN(n6789) );
  NAND2_X1 U7749 ( .A1(n8129), .A2(n7129), .ZN(n7128) );
  OR2_X1 U7750 ( .A1(n13124), .A2(n12931), .ZN(n9363) );
  NAND2_X1 U7751 ( .A1(n10452), .A2(n7115), .ZN(n6684) );
  NOR2_X1 U7752 ( .A1(n7880), .A2(n7116), .ZN(n7115) );
  INV_X1 U7753 ( .A(n7859), .ZN(n7116) );
  NAND2_X1 U7754 ( .A1(n7860), .A2(n7859), .ZN(n7119) );
  INV_X1 U7755 ( .A(n8158), .ZN(n7544) );
  NAND2_X2 U7756 ( .A1(n14689), .A2(n10020), .ZN(n12604) );
  INV_X1 U7757 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7641) );
  INV_X1 U7758 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7640) );
  INV_X1 U7759 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n7639) );
  INV_X1 U7760 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8136) );
  NOR2_X1 U7761 ( .A1(n11061), .A2(n7453), .ZN(n7449) );
  INV_X1 U7762 ( .A(n13365), .ZN(n13318) );
  INV_X1 U7763 ( .A(n13979), .ZN(n6968) );
  INV_X1 U7764 ( .A(n7261), .ZN(n6991) );
  AND2_X1 U7765 ( .A1(n6991), .A2(n6989), .ZN(n6987) );
  OAI21_X1 U7766 ( .B1(n7261), .B2(n7267), .A(n13721), .ZN(n7260) );
  INV_X1 U7767 ( .A(n13634), .ZN(n7197) );
  NOR2_X1 U7768 ( .A1(n6983), .A2(n6982), .ZN(n6981) );
  INV_X1 U7769 ( .A(n11502), .ZN(n6983) );
  AND2_X1 U7770 ( .A1(n11762), .A2(n10408), .ZN(n7190) );
  INV_X1 U7771 ( .A(n10410), .ZN(n7193) );
  OR2_X1 U7772 ( .A1(n10243), .A2(n10221), .ZN(n11447) );
  NAND2_X1 U7773 ( .A1(n14405), .A2(n10218), .ZN(n10232) );
  NAND2_X1 U7774 ( .A1(n10215), .A2(n7445), .ZN(n10230) );
  NAND2_X1 U7775 ( .A1(n10228), .A2(n10230), .ZN(n11444) );
  OAI21_X1 U7776 ( .B1(n8118), .B2(n8117), .A(n8119), .ZN(n9294) );
  INV_X1 U7777 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U7778 ( .A1(n8048), .A2(SI_24_), .ZN(n8049) );
  OR2_X1 U7779 ( .A1(n8046), .A2(n6784), .ZN(n8050) );
  INV_X1 U7780 ( .A(n8047), .ZN(n6784) );
  XNOR2_X1 U7781 ( .A(n8048), .B(SI_24_), .ZN(n8046) );
  NAND2_X1 U7782 ( .A1(n10174), .A2(n9410), .ZN(n9576) );
  NOR2_X1 U7783 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n9413) );
  OAI211_X1 U7784 ( .C1(n7965), .C2(n10167), .A(n7221), .B(n7219), .ZN(n7977)
         );
  NAND2_X1 U7785 ( .A1(n7220), .A2(SI_20_), .ZN(n7219) );
  NAND2_X1 U7786 ( .A1(n7965), .A2(n6564), .ZN(n7221) );
  INV_X1 U7787 ( .A(n7964), .ZN(n7220) );
  NAND2_X1 U7788 ( .A1(n7256), .A2(n7619), .ZN(n7726) );
  OAI21_X1 U7789 ( .B1(n7607), .B2(SI_9_), .A(n7609), .ZN(n7881) );
  NAND2_X1 U7790 ( .A1(n6903), .A2(n6993), .ZN(n7882) );
  AOI21_X1 U7791 ( .B1(n6995), .B2(n6997), .A(n6994), .ZN(n6993) );
  NAND2_X1 U7792 ( .A1(n7845), .A2(n6995), .ZN(n6903) );
  INV_X1 U7793 ( .A(n7606), .ZN(n6994) );
  INV_X1 U7794 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U7795 ( .A1(n14001), .A2(n6765), .ZN(n14002) );
  NAND2_X1 U7796 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6766), .ZN(n6765) );
  INV_X1 U7797 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6766) );
  XNOR2_X1 U7798 ( .A(n6452), .B(n10703), .ZN(n9075) );
  AND2_X1 U7799 ( .A1(n9142), .A2(n9140), .ZN(n11874) );
  NAND2_X1 U7800 ( .A1(n11851), .A2(n6509), .ZN(n7062) );
  NAND2_X1 U7801 ( .A1(n11851), .A2(n9124), .ZN(n9125) );
  AND2_X1 U7802 ( .A1(n7052), .A2(n9112), .ZN(n7051) );
  NAND2_X1 U7803 ( .A1(n11892), .A2(n7053), .ZN(n7052) );
  NAND2_X1 U7804 ( .A1(n11892), .A2(n7055), .ZN(n7054) );
  INV_X1 U7805 ( .A(n9109), .ZN(n7055) );
  AND4_X1 U7806 ( .A1(n8657), .A2(n8656), .A3(n8655), .A4(n8654), .ZN(n9007)
         );
  NAND2_X1 U7807 ( .A1(n7168), .A2(n7167), .ZN(n10138) );
  INV_X1 U7808 ( .A(n10304), .ZN(n7167) );
  NAND2_X1 U7809 ( .A1(n10142), .A2(n7169), .ZN(n7168) );
  NAND2_X1 U7810 ( .A1(P3_REG2_REG_0__SCAN_IN), .A2(n14746), .ZN(n7169) );
  INV_X1 U7811 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10692) );
  INV_X1 U7812 ( .A(n14769), .ZN(n7147) );
  NOR2_X1 U7813 ( .A1(n14765), .A2(n10893), .ZN(n10894) );
  XNOR2_X1 U7814 ( .A(n10842), .B(n10898), .ZN(n14797) );
  NAND2_X1 U7815 ( .A1(n14797), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n14796) );
  NAND2_X1 U7816 ( .A1(n7166), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7165) );
  NAND2_X1 U7817 ( .A1(n10906), .A2(n7166), .ZN(n7164) );
  INV_X1 U7818 ( .A(n10908), .ZN(n7166) );
  NAND2_X1 U7819 ( .A1(n14847), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U7820 ( .A1(n12032), .A2(n6851), .ZN(n12054) );
  OR2_X1 U7821 ( .A1(n12033), .A2(n12021), .ZN(n6851) );
  NAND2_X1 U7822 ( .A1(n12081), .A2(n12083), .ZN(n12108) );
  NAND2_X1 U7823 ( .A1(n7389), .A2(n7393), .ZN(n7386) );
  NAND2_X1 U7824 ( .A1(n7393), .A2(n7394), .ZN(n7387) );
  NAND2_X1 U7825 ( .A1(n8774), .A2(n8914), .ZN(n12199) );
  AND2_X1 U7826 ( .A1(n8761), .A2(n8760), .ZN(n12226) );
  INV_X1 U7827 ( .A(n9015), .ZN(n12227) );
  AND2_X1 U7828 ( .A1(n8735), .A2(n8734), .ZN(n12249) );
  NOR2_X1 U7829 ( .A1(n12247), .A2(n7424), .ZN(n7421) );
  NAND2_X1 U7830 ( .A1(n9013), .A2(n7425), .ZN(n7422) );
  INV_X1 U7831 ( .A(n12250), .ZN(n12247) );
  NAND2_X1 U7832 ( .A1(n8897), .A2(n8898), .ZN(n12250) );
  INV_X1 U7833 ( .A(n12306), .ZN(n12283) );
  NAND2_X1 U7834 ( .A1(n8672), .A2(n8928), .ZN(n7382) );
  OR2_X1 U7835 ( .A1(n12496), .A2(n12305), .ZN(n8929) );
  OAI21_X1 U7836 ( .B1(n9006), .B2(n7415), .A(n7414), .ZN(n12304) );
  AOI21_X1 U7837 ( .B1(n7416), .B2(n12334), .A(n6527), .ZN(n7414) );
  INV_X1 U7838 ( .A(n7416), .ZN(n7415) );
  AND2_X1 U7839 ( .A1(n7564), .A2(n9008), .ZN(n7416) );
  AOI21_X1 U7840 ( .B1(n7356), .B2(n7358), .A(n6569), .ZN(n7354) );
  NAND2_X1 U7841 ( .A1(n9006), .A2(n9005), .ZN(n12328) );
  NAND2_X1 U7842 ( .A1(n12373), .A2(n12372), .ZN(n12375) );
  INV_X1 U7843 ( .A(n11920), .ZN(n12384) );
  NAND2_X1 U7844 ( .A1(n11357), .A2(n11356), .ZN(n11359) );
  NAND2_X1 U7845 ( .A1(n11352), .A2(n11353), .ZN(n11351) );
  AND2_X1 U7846 ( .A1(n7406), .A2(n7404), .ZN(n7403) );
  NAND2_X1 U7847 ( .A1(n10949), .A2(n7407), .ZN(n7405) );
  INV_X1 U7848 ( .A(n11992), .ZN(n11155) );
  AND4_X1 U7849 ( .A1(n8524), .A2(n8523), .A3(n8522), .A4(n8521), .ZN(n11303)
         );
  INV_X1 U7850 ( .A(n14881), .ZN(n10918) );
  AND4_X1 U7851 ( .A1(n8472), .A2(n8471), .A3(n8470), .A4(n8469), .ZN(n10947)
         );
  OR2_X1 U7852 ( .A1(n8453), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8466) );
  NAND2_X1 U7853 ( .A1(n10946), .A2(n10945), .ZN(n10944) );
  AND3_X1 U7854 ( .A1(n8451), .A2(n8450), .A3(n8449), .ZN(n10630) );
  AND4_X1 U7855 ( .A1(n8459), .A2(n8458), .A3(n8457), .A4(n8456), .ZN(n10920)
         );
  NAND2_X1 U7856 ( .A1(n8753), .A2(n8752), .ZN(n9063) );
  OR2_X1 U7857 ( .A1(n6787), .A2(n11259), .ZN(n8752) );
  NAND2_X1 U7858 ( .A1(n8727), .A2(n8726), .ZN(n12413) );
  NAND2_X1 U7859 ( .A1(n9047), .A2(n10196), .ZN(n14915) );
  OR2_X1 U7860 ( .A1(n8653), .A2(n8391), .ZN(n8393) );
  NOR2_X1 U7861 ( .A1(n7440), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n7439) );
  OAI21_X1 U7862 ( .B1(n8776), .B2(n8299), .A(n8298), .ZN(n8358) );
  NAND2_X1 U7863 ( .A1(n8292), .A2(n8291), .ZN(n8751) );
  OR2_X1 U7864 ( .A1(n8738), .A2(n8290), .ZN(n8292) );
  NOR2_X1 U7865 ( .A1(n7430), .A2(n7435), .ZN(n7429) );
  NOR2_X1 U7866 ( .A1(n8955), .A2(n7027), .ZN(n6780) );
  INV_X1 U7867 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n8955) );
  NOR2_X1 U7868 ( .A1(n7435), .A2(n7433), .ZN(n7431) );
  NAND2_X1 U7869 ( .A1(n8599), .A2(n8598), .ZN(n8601) );
  NAND2_X1 U7870 ( .A1(n8264), .A2(n9991), .ZN(n7086) );
  INV_X1 U7871 ( .A(n7083), .ZN(n7082) );
  NAND2_X1 U7872 ( .A1(n8526), .A2(n8525), .ZN(n8528) );
  NAND2_X1 U7873 ( .A1(n9698), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8253) );
  AND2_X1 U7874 ( .A1(n8255), .A2(n8254), .ZN(n8496) );
  NAND2_X1 U7875 ( .A1(n8476), .A2(n8253), .ZN(n8497) );
  AND2_X1 U7876 ( .A1(n7107), .A2(n8496), .ZN(n7106) );
  NAND2_X1 U7877 ( .A1(n8473), .A2(n8253), .ZN(n7107) );
  NAND2_X1 U7878 ( .A1(n8251), .A2(n8250), .ZN(n8474) );
  OR2_X1 U7879 ( .A1(n8430), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n8432) );
  AND2_X1 U7880 ( .A1(n8248), .A2(n8247), .ZN(n8446) );
  NAND2_X1 U7881 ( .A1(n9648), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8246) );
  CLKBUF_X1 U7882 ( .A(n8375), .Z(n8376) );
  NAND2_X1 U7883 ( .A1(n7027), .A2(n6856), .ZN(n6855) );
  INV_X1 U7884 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6856) );
  AOI21_X1 U7885 ( .B1(n11283), .B2(n6499), .A(n7329), .ZN(n11414) );
  OAI21_X1 U7886 ( .B1(n7331), .B2(n7330), .A(n6533), .ZN(n7329) );
  NAND2_X1 U7887 ( .A1(n11414), .A2(n11415), .ZN(n12534) );
  AND2_X1 U7888 ( .A1(n12696), .A2(n12543), .ZN(n7309) );
  AND2_X1 U7889 ( .A1(n12589), .A2(n6500), .ZN(n7307) );
  NAND2_X1 U7890 ( .A1(n12606), .A2(n12599), .ZN(n7343) );
  INV_X1 U7891 ( .A(n12535), .ZN(n7324) );
  NAND2_X1 U7892 ( .A1(n8037), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8070) );
  INV_X1 U7893 ( .A(n8038), .ZN(n8037) );
  INV_X1 U7894 ( .A(n10032), .ZN(n7298) );
  INV_X1 U7895 ( .A(n10033), .ZN(n7299) );
  NAND2_X1 U7896 ( .A1(n10589), .A2(n10586), .ZN(n7315) );
  INV_X1 U7897 ( .A(n10533), .ZN(n7312) );
  NAND2_X1 U7898 ( .A1(n10788), .A2(n7317), .ZN(n7316) );
  INV_X1 U7899 ( .A(n7315), .ZN(n7314) );
  OAI21_X1 U7900 ( .B1(n12611), .B2(n12688), .A(n12687), .ZN(n12686) );
  XNOR2_X1 U7901 ( .A(n10029), .B(n10028), .ZN(n12687) );
  NAND2_X1 U7902 ( .A1(n7833), .A2(n7832), .ZN(n7841) );
  NAND2_X1 U7903 ( .A1(n10205), .A2(n6693), .ZN(n6695) );
  NOR2_X1 U7904 ( .A1(n10207), .A2(n6694), .ZN(n6693) );
  INV_X1 U7905 ( .A(n7560), .ZN(n6694) );
  XNOR2_X1 U7906 ( .A(n13167), .B(n6816), .ZN(n12535) );
  NAND2_X1 U7907 ( .A1(n12534), .A2(n12533), .ZN(n7327) );
  AND2_X1 U7908 ( .A1(n9381), .A2(n9380), .ZN(n9388) );
  AND4_X1 U7909 ( .A1(n7840), .A2(n7839), .A3(n7838), .A4(n7837), .ZN(n10453)
         );
  OR2_X1 U7910 ( .A1(n7763), .A2(n9965), .ZN(n7766) );
  NAND2_X1 U7911 ( .A1(n7128), .A2(n9377), .ZN(n7126) );
  INV_X1 U7912 ( .A(n12887), .ZN(n12602) );
  NAND2_X1 U7913 ( .A1(n12886), .A2(n6508), .ZN(n12866) );
  AND2_X1 U7914 ( .A1(n8104), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12859) );
  AOI21_X1 U7915 ( .B1(n12886), .B2(n12868), .A(n12867), .ZN(n6667) );
  NAND2_X1 U7916 ( .A1(n12866), .A2(n13065), .ZN(n6682) );
  NAND2_X1 U7917 ( .A1(n12885), .A2(n12884), .ZN(n12886) );
  INV_X1 U7918 ( .A(n7496), .ZN(n7495) );
  OAI21_X1 U7919 ( .B1(n12929), .B2(n7497), .A(n7504), .ZN(n7496) );
  NAND2_X1 U7920 ( .A1(n12923), .A2(n12657), .ZN(n7504) );
  XNOR2_X1 U7921 ( .A(n13113), .B(n12657), .ZN(n12924) );
  INV_X1 U7922 ( .A(n12941), .ZN(n7500) );
  AOI21_X1 U7923 ( .B1(n7158), .B2(n7161), .A(n6538), .ZN(n7157) );
  OR2_X1 U7924 ( .A1(n6670), .A2(n7563), .ZN(n6669) );
  INV_X1 U7925 ( .A(n12924), .ZN(n12915) );
  NAND2_X1 U7926 ( .A1(n6542), .A2(n7162), .ZN(n7160) );
  NAND2_X1 U7927 ( .A1(n9374), .A2(n7162), .ZN(n7161) );
  OR2_X1 U7928 ( .A1(n12959), .A2(n12963), .ZN(n7163) );
  NAND2_X1 U7929 ( .A1(n12973), .A2(n7563), .ZN(n12959) );
  INV_X1 U7930 ( .A(n7537), .ZN(n7534) );
  OR2_X1 U7931 ( .A1(n13142), .A2(n12976), .ZN(n7537) );
  NAND2_X1 U7932 ( .A1(n7536), .A2(n7538), .ZN(n7535) );
  INV_X1 U7933 ( .A(n12992), .ZN(n7536) );
  XNOR2_X1 U7934 ( .A(n13134), .B(n13005), .ZN(n12986) );
  NAND2_X1 U7935 ( .A1(n12974), .A2(n12986), .ZN(n12973) );
  AND2_X1 U7936 ( .A1(n6673), .A2(n6562), .ZN(n13000) );
  OR2_X1 U7937 ( .A1(n13012), .A2(n6554), .ZN(n6673) );
  INV_X1 U7938 ( .A(n7970), .ZN(n7968) );
  NAND2_X1 U7939 ( .A1(n13031), .A2(n13022), .ZN(n13016) );
  INV_X1 U7940 ( .A(n7721), .ZN(n7665) );
  AOI21_X1 U7941 ( .B1(n6685), .B2(n6662), .A(n6568), .ZN(n13027) );
  NOR2_X1 U7942 ( .A1(n7132), .A2(n7134), .ZN(n6662) );
  AND2_X1 U7943 ( .A1(n13157), .A2(n13058), .ZN(n7132) );
  NOR2_X1 U7944 ( .A1(n8181), .A2(n7558), .ZN(n7557) );
  NAND2_X1 U7945 ( .A1(n8179), .A2(n7559), .ZN(n13062) );
  AND2_X1 U7946 ( .A1(n9371), .A2(n8178), .ZN(n7559) );
  AOI21_X1 U7947 ( .B1(n6824), .B2(n6823), .A(n6822), .ZN(n13054) );
  NAND2_X1 U7948 ( .A1(n13167), .A2(n13056), .ZN(n6823) );
  NOR2_X1 U7949 ( .A1(n13056), .A2(n13167), .ZN(n6822) );
  NAND2_X2 U7950 ( .A1(n7750), .A2(n7749), .ZN(n11406) );
  OAI21_X1 U7951 ( .B1(n11114), .B2(n8173), .A(n8174), .ZN(n11209) );
  NAND2_X1 U7952 ( .A1(n6671), .A2(n7937), .ZN(n11116) );
  NAND2_X1 U7953 ( .A1(n10771), .A2(n7149), .ZN(n6671) );
  INV_X1 U7954 ( .A(n7915), .ZN(n7662) );
  NAND2_X1 U7955 ( .A1(n10771), .A2(n7922), .ZN(n10965) );
  AND2_X1 U7956 ( .A1(n8169), .A2(n7921), .ZN(n10776) );
  OAI211_X1 U7957 ( .C1(n8165), .C2(n7513), .A(n7511), .B(n10744), .ZN(n10747)
         );
  INV_X1 U7958 ( .A(n8166), .ZN(n7513) );
  NAND2_X1 U7959 ( .A1(n8165), .A2(n7514), .ZN(n10726) );
  OAI21_X1 U7960 ( .B1(n10389), .B2(n9337), .A(n7870), .ZN(n10731) );
  AND4_X1 U7961 ( .A1(n7858), .A2(n7857), .A3(n7856), .A4(n7855), .ZN(n10591)
         );
  NAND2_X1 U7962 ( .A1(n10422), .A2(n10417), .ZN(n10416) );
  INV_X1 U7963 ( .A(n13004), .ZN(n13057) );
  INV_X1 U7964 ( .A(n10663), .ZN(n7013) );
  XNOR2_X1 U7965 ( .A(n12743), .B(n10383), .ZN(n10377) );
  AND2_X1 U7966 ( .A1(n8143), .A2(n9958), .ZN(n13004) );
  AND2_X1 U7967 ( .A1(n8144), .A2(n9958), .ZN(n13002) );
  INV_X1 U7968 ( .A(n13022), .ZN(n13148) );
  INV_X1 U7969 ( .A(n13045), .ZN(n13157) );
  NAND2_X1 U7970 ( .A1(n10224), .A2(n7682), .ZN(n7148) );
  INV_X1 U7971 ( .A(n10383), .ZN(n14651) );
  OR3_X1 U7972 ( .A1(n13203), .A2(n11239), .A3(n11295), .ZN(n9946) );
  NAND2_X1 U7973 ( .A1(n8209), .A2(n8208), .ZN(n8214) );
  INV_X1 U7974 ( .A(n8207), .ZN(n8209) );
  AND2_X1 U7975 ( .A1(n7656), .A2(n8132), .ZN(n10418) );
  OR2_X1 U7976 ( .A1(n7655), .A2(n13189), .ZN(n7654) );
  NOR2_X1 U7977 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7539) );
  AND2_X1 U7978 ( .A1(n7456), .A2(n6647), .ZN(n6646) );
  INV_X1 U7979 ( .A(n13397), .ZN(n6648) );
  NAND2_X1 U7980 ( .A1(n11069), .A2(n11068), .ZN(n6760) );
  AND2_X1 U7981 ( .A1(n6455), .A2(n7454), .ZN(n7451) );
  AND2_X1 U7982 ( .A1(n11223), .A2(n11222), .ZN(n11514) );
  NAND2_X1 U7983 ( .A1(n6634), .A2(n13417), .ZN(n13395) );
  AOI21_X1 U7984 ( .B1(n13345), .B2(n6632), .A(n6631), .ZN(n6630) );
  INV_X1 U7985 ( .A(n13345), .ZN(n6633) );
  XNOR2_X1 U7986 ( .A(n10488), .B(n10486), .ZN(n10502) );
  NOR2_X1 U7987 ( .A1(n10502), .A2(n10503), .ZN(n10501) );
  OAI21_X1 U7988 ( .B1(n9861), .B2(n13364), .A(n9860), .ZN(n9862) );
  INV_X1 U7989 ( .A(n10221), .ZN(n10240) );
  XNOR2_X1 U7990 ( .A(n9926), .B(n13365), .ZN(n10002) );
  NAND2_X1 U7991 ( .A1(n7445), .A2(n6444), .ZN(n7443) );
  INV_X1 U7992 ( .A(n13262), .ZN(n7469) );
  NAND2_X1 U7993 ( .A1(n7277), .A2(n7276), .ZN(n7275) );
  NAND2_X1 U7994 ( .A1(n11786), .A2(n11788), .ZN(n7276) );
  NAND2_X1 U7995 ( .A1(n11787), .A2(n7278), .ZN(n7277) );
  AND2_X1 U7996 ( .A1(n7272), .A2(n6880), .ZN(n6879) );
  NAND2_X1 U7997 ( .A1(n6659), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6658) );
  INV_X1 U7998 ( .A(n11634), .ZN(n6659) );
  OAI21_X1 U7999 ( .B1(n6971), .B2(n6968), .A(n6969), .ZN(n6967) );
  NAND2_X1 U8000 ( .A1(n9557), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U8001 ( .A1(n9557), .A2(n6970), .ZN(n6969) );
  AND2_X1 U8002 ( .A1(n6968), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6970) );
  AND2_X1 U8003 ( .A1(n13737), .A2(n13738), .ZN(n6844) );
  NOR2_X1 U8004 ( .A1(n13737), .A2(n13738), .ZN(n13736) );
  OR2_X1 U8005 ( .A1(n13740), .A2(n14380), .ZN(n6842) );
  NAND2_X1 U8006 ( .A1(n13770), .A2(n7214), .ZN(n13752) );
  NOR2_X1 U8007 ( .A1(n13756), .A2(n7215), .ZN(n7214) );
  INV_X1 U8008 ( .A(n13643), .ZN(n7215) );
  NAND2_X1 U8009 ( .A1(n13773), .A2(n13772), .ZN(n13771) );
  NAND2_X1 U8010 ( .A1(n13784), .A2(n13785), .ZN(n6920) );
  NAND2_X1 U8011 ( .A1(n6920), .A2(n6918), .ZN(n13770) );
  NOR2_X1 U8012 ( .A1(n6919), .A2(n13772), .ZN(n6918) );
  INV_X1 U8013 ( .A(n13642), .ZN(n6919) );
  NOR2_X1 U8014 ( .A1(n13807), .A2(n7211), .ZN(n7210) );
  INV_X1 U8015 ( .A(n13640), .ZN(n7211) );
  NAND2_X1 U8016 ( .A1(n13829), .A2(n13662), .ZN(n13815) );
  OR2_X1 U8017 ( .A1(n13811), .A2(n13663), .ZN(n13812) );
  OR2_X1 U8018 ( .A1(n13873), .A2(n13633), .ZN(n13635) );
  NAND2_X1 U8019 ( .A1(n6539), .A2(n11502), .ZN(n6980) );
  NAND2_X1 U8020 ( .A1(n11175), .A2(n6981), .ZN(n6975) );
  NAND2_X1 U8021 ( .A1(n7207), .A2(n7206), .ZN(n13630) );
  INV_X1 U8022 ( .A(n6485), .ZN(n7206) );
  OR2_X1 U8023 ( .A1(n10994), .A2(n11767), .ZN(n6955) );
  INV_X1 U8024 ( .A(n11761), .ZN(n7181) );
  OR2_X1 U8025 ( .A1(n11747), .A2(n13505), .ZN(n14380) );
  INV_X1 U8026 ( .A(n13652), .ZN(n7234) );
  NAND2_X1 U8027 ( .A1(n10392), .A2(n10391), .ZN(n14515) );
  XNOR2_X1 U8028 ( .A(n8080), .B(n8065), .ZN(n13200) );
  NOR2_X1 U8029 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6947) );
  INV_X1 U8030 ( .A(n7200), .ZN(n7441) );
  XNOR2_X1 U8031 ( .A(n8010), .B(n8009), .ZN(n11627) );
  NAND2_X1 U8032 ( .A1(n10476), .A2(n9566), .ZN(n9571) );
  XNOR2_X1 U8033 ( .A(n7977), .B(n7994), .ZN(n11579) );
  XNOR2_X1 U8034 ( .A(n7963), .B(n7962), .ZN(n11533) );
  NAND2_X1 U8035 ( .A1(n6914), .A2(n7630), .ZN(n7963) );
  NAND2_X1 U8036 ( .A1(n7607), .A2(SI_9_), .ZN(n7609) );
  NAND2_X1 U8037 ( .A1(n9746), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9817) );
  INV_X1 U8038 ( .A(n6996), .ZN(n6995) );
  OAI21_X1 U8039 ( .B1(n7844), .B2(n6997), .A(n7861), .ZN(n6996) );
  NAND2_X1 U8040 ( .A1(n7807), .A2(n7594), .ZN(n7815) );
  NAND2_X1 U8041 ( .A1(n6917), .A2(n6916), .ZN(n6915) );
  AND2_X1 U8042 ( .A1(n7019), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14045) );
  INV_X1 U8043 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7019) );
  NOR2_X1 U8044 ( .A1(n14058), .A2(n14059), .ZN(n14060) );
  NAND2_X1 U8045 ( .A1(n14010), .A2(n14009), .ZN(n14061) );
  NAND2_X1 U8046 ( .A1(n14055), .A2(n15109), .ZN(n14009) );
  AOI21_X1 U8047 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n15066), .A(n14018), .ZN(
        n14037) );
  OAI22_X1 U8048 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14026), .B1(n14033), 
        .B2(n14025), .ZN(n14083) );
  NAND2_X1 U8049 ( .A1(n7056), .A2(n14134), .ZN(n14143) );
  OAI21_X1 U8050 ( .B1(n14135), .B2(n14136), .A(P2_ADDR_REG_17__SCAN_IN), .ZN(
        n7056) );
  INV_X1 U8051 ( .A(n7048), .ZN(n7042) );
  NAND2_X1 U8052 ( .A1(n7044), .A2(n7046), .ZN(n7043) );
  INV_X1 U8053 ( .A(n7047), .ZN(n7046) );
  AND3_X1 U8054 ( .A1(n8682), .A2(n8681), .A3(n8680), .ZN(n12295) );
  NAND2_X1 U8055 ( .A1(n11167), .A2(n11166), .ZN(n11165) );
  AND4_X1 U8056 ( .A1(n8612), .A2(n8611), .A3(n8610), .A4(n8609), .ZN(n12385)
         );
  NAND2_X1 U8057 ( .A1(n8625), .A2(n8624), .ZN(n12361) );
  OR2_X1 U8058 ( .A1(n9845), .A2(n8617), .ZN(n8625) );
  NAND2_X1 U8059 ( .A1(n10689), .A2(n6774), .ZN(n10805) );
  NAND2_X1 U8060 ( .A1(n9077), .A2(n10707), .ZN(n6774) );
  AND4_X1 U8061 ( .A1(n8596), .A2(n8595), .A3(n8594), .A4(n8593), .ZN(n12369)
         );
  OAI21_X1 U8062 ( .B1(n11861), .B2(n9093), .A(n9099), .ZN(n11923) );
  AND2_X1 U8063 ( .A1(n8713), .A2(n8712), .ZN(n12282) );
  NAND2_X1 U8064 ( .A1(n6601), .A2(n8926), .ZN(n7110) );
  NAND2_X1 U8065 ( .A1(n6604), .A2(n6602), .ZN(n6601) );
  INV_X1 U8066 ( .A(n12295), .ZN(n12319) );
  INV_X1 U8067 ( .A(n9007), .ZN(n12344) );
  INV_X1 U8068 ( .A(n12369), .ZN(n11989) );
  INV_X1 U8069 ( .A(n11937), .ZN(n11990) );
  NAND4_X1 U8070 ( .A1(n8509), .A2(n8508), .A3(n8507), .A4(n8506), .ZN(n14887)
         );
  INV_X1 U8071 ( .A(n10854), .ZN(n14765) );
  NOR2_X1 U8072 ( .A1(n10848), .A2(n10849), .ZN(n11097) );
  OR2_X1 U8073 ( .A1(n12029), .A2(n12061), .ZN(n7131) );
  INV_X1 U8074 ( .A(n12178), .ZN(n6860) );
  AOI21_X1 U8075 ( .B1(n12522), .B2(n8778), .A(n8777), .ZN(n12193) );
  OAI21_X1 U8076 ( .B1(n9024), .B2(n14891), .A(n9023), .ZN(n7350) );
  NAND2_X1 U8077 ( .A1(n7388), .A2(n7394), .ZN(n12212) );
  NAND2_X1 U8078 ( .A1(n7395), .A2(n8888), .ZN(n12260) );
  NAND2_X1 U8079 ( .A1(n8706), .A2(n8705), .ZN(n12276) );
  NAND2_X1 U8080 ( .A1(n8576), .A2(n8575), .ZN(n14162) );
  INV_X1 U8081 ( .A(n12193), .ZN(n8787) );
  INV_X1 U8082 ( .A(n9063), .ZN(n12475) );
  AND2_X1 U8083 ( .A1(n9031), .A2(n9030), .ZN(n12512) );
  XNOR2_X1 U8084 ( .A(n8797), .B(P3_IR_REG_22__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U8085 ( .A1(n10534), .A2(n10533), .ZN(n10588) );
  AND2_X1 U8086 ( .A1(n8077), .A2(n8076), .ZN(n12629) );
  NOR2_X1 U8087 ( .A1(n6469), .A2(n12724), .ZN(n7336) );
  NAND2_X1 U8088 ( .A1(n7339), .A2(n7343), .ZN(n7338) );
  NAND2_X1 U8089 ( .A1(n8103), .A2(n8102), .ZN(n13096) );
  NAND2_X1 U8090 ( .A1(n7334), .A2(n7332), .ZN(n11313) );
  AND2_X1 U8091 ( .A1(n7334), .A2(n7333), .ZN(n11284) );
  NAND2_X1 U8092 ( .A1(n11283), .A2(n11282), .ZN(n7334) );
  AND2_X1 U8093 ( .A1(n8022), .A2(n8021), .ZN(n12675) );
  INV_X1 U8094 ( .A(n12939), .ZN(n13118) );
  NAND2_X1 U8095 ( .A1(n10791), .A2(n10792), .ZN(n10932) );
  NAND2_X1 U8096 ( .A1(n7328), .A2(n7331), .ZN(n11413) );
  NAND2_X1 U8097 ( .A1(n11283), .A2(n6457), .ZN(n7328) );
  NAND2_X1 U8098 ( .A1(n6703), .A2(n12572), .ZN(n12707) );
  NAND2_X1 U8099 ( .A1(n8094), .A2(n8093), .ZN(n12727) );
  INV_X1 U8100 ( .A(n12629), .ZN(n12918) );
  INV_X1 U8101 ( .A(n12675), .ZN(n12931) );
  NAND4_X1 U8102 ( .A1(n7825), .A2(n7824), .A3(n7823), .A4(n7822), .ZN(n12741)
         );
  OR2_X1 U8103 ( .A1(n7762), .A2(n13080), .ZN(n6775) );
  AND3_X1 U8104 ( .A1(n7751), .A2(n6518), .A3(n7752), .ZN(n6769) );
  NAND2_X1 U8105 ( .A1(n9954), .A2(n14637), .ZN(n12998) );
  NAND2_X1 U8106 ( .A1(n7010), .A2(n9454), .ZN(n7009) );
  OR2_X1 U8107 ( .A1(n9454), .A2(n12749), .ZN(n7760) );
  NAND2_X1 U8108 ( .A1(n8229), .A2(n8228), .ZN(n14636) );
  NAND2_X1 U8109 ( .A1(n10272), .A2(n10271), .ZN(n14506) );
  OAI21_X1 U8110 ( .B1(n13459), .B2(n13336), .A(n7456), .ZN(n13363) );
  NAND2_X1 U8111 ( .A1(n13458), .A2(n6786), .ZN(n6785) );
  NOR2_X1 U8112 ( .A1(n13337), .A2(n13336), .ZN(n6786) );
  NAND2_X1 U8113 ( .A1(n14195), .A2(n13240), .ZN(n14199) );
  AND4_X1 U8114 ( .A1(n11183), .A2(n11182), .A3(n11181), .A4(n11180), .ZN(
        n14208) );
  NAND2_X1 U8115 ( .A1(n6637), .A2(n6636), .ZN(n6635) );
  INV_X1 U8116 ( .A(n11340), .ZN(n6636) );
  NAND2_X1 U8117 ( .A1(n10549), .A2(n10548), .ZN(n14537) );
  NAND2_X1 U8118 ( .A1(n11599), .A2(n11598), .ZN(n13945) );
  INV_X1 U8119 ( .A(n14265), .ZN(n13659) );
  NAND2_X1 U8120 ( .A1(n14231), .A2(n14232), .ZN(n14230) );
  AND2_X1 U8121 ( .A1(n10099), .A2(n11795), .ZN(n14241) );
  NAND2_X1 U8122 ( .A1(n14416), .A2(n9870), .ZN(n14238) );
  INV_X1 U8123 ( .A(n14221), .ZN(n14233) );
  OR2_X1 U8124 ( .A1(n11747), .A2(n13984), .ZN(n14382) );
  NAND4_X1 U8125 ( .A1(n10104), .A2(n10103), .A3(n10102), .A4(n10101), .ZN(
        n13483) );
  NAND2_X1 U8126 ( .A1(n6927), .A2(n6926), .ZN(n13886) );
  OR2_X1 U8127 ( .A1(n13622), .A2(n13887), .ZN(n6927) );
  NOR2_X1 U8128 ( .A1(n13621), .A2(n14468), .ZN(n6926) );
  NAND2_X1 U8129 ( .A1(n13691), .A2(n6514), .ZN(n6744) );
  NAND2_X1 U8130 ( .A1(n13692), .A2(n14429), .ZN(n13696) );
  NAND2_X1 U8131 ( .A1(n13725), .A2(n13649), .ZN(n13720) );
  NAND2_X1 U8132 ( .A1(n13195), .A2(n11743), .ZN(n7006) );
  NAND2_X1 U8133 ( .A1(n11513), .A2(n11512), .ZN(n14271) );
  NAND2_X1 U8134 ( .A1(n10997), .A2(n10996), .ZN(n14226) );
  NAND2_X1 U8135 ( .A1(n9611), .A2(n9866), .ZN(n14416) );
  NAND2_X1 U8136 ( .A1(n13653), .A2(n7234), .ZN(n7233) );
  NOR2_X1 U8137 ( .A1(n14489), .A2(n7230), .ZN(n7229) );
  OR2_X1 U8138 ( .A1(n7236), .A2(n7230), .ZN(n7227) );
  NAND2_X1 U8139 ( .A1(n7230), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7235) );
  NAND2_X1 U8140 ( .A1(n13896), .A2(n7232), .ZN(n7225) );
  NOR2_X1 U8141 ( .A1(n13653), .A2(n7234), .ZN(n7232) );
  INV_X1 U8142 ( .A(n13896), .ZN(n7223) );
  NAND2_X1 U8143 ( .A1(n6755), .A2(n14544), .ZN(n6754) );
  INV_X1 U8144 ( .A(n13916), .ZN(n6755) );
  NAND2_X1 U8145 ( .A1(n6759), .A2(n14544), .ZN(n6758) );
  INV_X1 U8146 ( .A(n13928), .ZN(n6759) );
  XNOR2_X1 U8147 ( .A(n14074), .B(n7076), .ZN(n14108) );
  INV_X1 U8148 ( .A(n14075), .ZN(n7076) );
  AND2_X1 U8149 ( .A1(n7072), .A2(n7070), .ZN(n14332) );
  NOR2_X1 U8150 ( .A1(n14332), .A2(n14333), .ZN(n14331) );
  OAI21_X1 U8151 ( .B1(n14088), .B2(n14087), .A(n14335), .ZN(n14339) );
  INV_X1 U8152 ( .A(n10228), .ZN(n11439) );
  INV_X1 U8153 ( .A(n10230), .ZN(n11440) );
  INV_X1 U8154 ( .A(n11466), .ZN(n6901) );
  OAI22_X1 U8155 ( .A1(n6712), .A2(n9201), .B1(n9200), .B2(n9199), .ZN(n9208)
         );
  NAND2_X1 U8156 ( .A1(n6735), .A2(n6732), .ZN(n9201) );
  INV_X1 U8157 ( .A(n11470), .ZN(n11473) );
  NAND2_X1 U8158 ( .A1(n11477), .A2(n7283), .ZN(n7282) );
  INV_X1 U8159 ( .A(n11476), .ZN(n7283) );
  NOR2_X1 U8160 ( .A1(n7488), .A2(n9210), .ZN(n7486) );
  NAND2_X1 U8161 ( .A1(n9216), .A2(n9218), .ZN(n6727) );
  NAND2_X1 U8162 ( .A1(n6867), .A2(n6866), .ZN(n6865) );
  OAI22_X1 U8163 ( .A1(n11489), .A2(n7270), .B1(n11490), .B2(n7269), .ZN(
        n11494) );
  INV_X1 U8164 ( .A(n11488), .ZN(n7269) );
  NOR2_X1 U8165 ( .A1(n11491), .A2(n11488), .ZN(n7270) );
  NOR2_X1 U8166 ( .A1(n6898), .A2(n11492), .ZN(n6897) );
  NAND2_X1 U8167 ( .A1(n6898), .A2(n11492), .ZN(n6896) );
  NAND2_X1 U8168 ( .A1(n9229), .A2(n9228), .ZN(n6741) );
  NAND2_X1 U8169 ( .A1(n6875), .A2(n6468), .ZN(n6872) );
  AOI21_X1 U8170 ( .B1(n6874), .B2(n6873), .A(n6870), .ZN(n6869) );
  INV_X1 U8171 ( .A(n11504), .ZN(n6873) );
  NAND2_X1 U8172 ( .A1(n6472), .A2(n6529), .ZN(n6870) );
  NOR2_X1 U8173 ( .A1(n7523), .A2(n9244), .ZN(n7520) );
  INV_X1 U8174 ( .A(n9240), .ZN(n7526) );
  NAND2_X1 U8175 ( .A1(n7519), .A2(n7518), .ZN(n7517) );
  INV_X1 U8176 ( .A(n7520), .ZN(n7519) );
  INV_X1 U8177 ( .A(n7521), .ZN(n7518) );
  NOR2_X1 U8178 ( .A1(n11566), .A2(n13846), .ZN(n11573) );
  NAND2_X1 U8179 ( .A1(n11601), .A2(n6885), .ZN(n6884) );
  INV_X1 U8180 ( .A(n11600), .ZN(n6885) );
  INV_X1 U8181 ( .A(n6723), .ZN(n6722) );
  AOI21_X1 U8182 ( .B1(n6471), .B2(n6723), .A(n6572), .ZN(n6721) );
  NAND2_X1 U8183 ( .A1(n11630), .A2(n7288), .ZN(n7287) );
  INV_X1 U8184 ( .A(n11631), .ZN(n7288) );
  AND2_X1 U8185 ( .A1(n9265), .A2(n6772), .ZN(n9266) );
  INV_X1 U8186 ( .A(n9269), .ZN(n7555) );
  NAND2_X1 U8187 ( .A1(n8900), .A2(n10132), .ZN(n6806) );
  NAND2_X1 U8188 ( .A1(n6808), .A2(n9044), .ZN(n6807) );
  NAND2_X1 U8189 ( .A1(n11677), .A2(n11679), .ZN(n7292) );
  NOR2_X1 U8190 ( .A1(n6491), .A2(n6890), .ZN(n6889) );
  INV_X1 U8191 ( .A(n8703), .ZN(n7100) );
  INV_X1 U8192 ( .A(n8285), .ZN(n7097) );
  INV_X1 U8193 ( .A(n9291), .ZN(n7480) );
  NAND2_X1 U8194 ( .A1(n7646), .A2(n6725), .ZN(n7648) );
  OR2_X1 U8195 ( .A1(n7831), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n7864) );
  OR2_X1 U8196 ( .A1(n11568), .A2(n13848), .ZN(n11567) );
  NAND2_X1 U8197 ( .A1(n8064), .A2(SI_26_), .ZN(n7001) );
  OAI21_X1 U8198 ( .B1(n7002), .B2(n7001), .A(n8079), .ZN(n7000) );
  INV_X1 U8199 ( .A(n7258), .ZN(n7257) );
  OAI21_X1 U8200 ( .B1(n7938), .B2(n7259), .A(n7576), .ZN(n7258) );
  INV_X1 U8201 ( .A(n7624), .ZN(n7255) );
  INV_X1 U8202 ( .A(n7619), .ZN(n7259) );
  AND2_X1 U8203 ( .A1(n7257), .A2(n6909), .ZN(n6908) );
  NAND2_X1 U8204 ( .A1(n6910), .A2(n7617), .ZN(n6909) );
  INV_X1 U8205 ( .A(n7923), .ZN(n6910) );
  NAND2_X1 U8206 ( .A1(n6908), .A2(n6911), .ZN(n6906) );
  INV_X1 U8207 ( .A(n7617), .ZN(n6911) );
  NAND2_X1 U8208 ( .A1(n7611), .A2(SI_10_), .ZN(n7613) );
  OAI21_X1 U8209 ( .B1(n9657), .B2(n9658), .A(n6840), .ZN(n7592) );
  NOR3_X1 U8210 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .A3(
        n14739), .ZN(n10304) );
  OR2_X1 U8211 ( .A1(n11097), .A2(n6857), .ZN(n12017) );
  NOR2_X1 U8212 ( .A1(n11098), .A2(n14988), .ZN(n6857) );
  NAND2_X1 U8213 ( .A1(n14151), .A2(n6812), .ZN(n12163) );
  OR2_X1 U8214 ( .A1(n12150), .A2(n12151), .ZN(n6812) );
  NAND2_X1 U8215 ( .A1(n8342), .A2(n8341), .ZN(n8767) );
  XNOR2_X1 U8216 ( .A(n9063), .B(n12226), .ZN(n9016) );
  OR2_X1 U8217 ( .A1(n12413), .A2(n12249), .ZN(n8903) );
  INV_X1 U8218 ( .A(n7421), .ZN(n7419) );
  NAND2_X1 U8219 ( .A1(n6591), .A2(n12266), .ZN(n7427) );
  OR2_X1 U8220 ( .A1(n12276), .A2(n12282), .ZN(n8899) );
  NAND2_X1 U8221 ( .A1(n6591), .A2(n6590), .ZN(n8898) );
  OR2_X1 U8222 ( .A1(n8697), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8707) );
  INV_X1 U8223 ( .A(n8888), .ZN(n8894) );
  INV_X1 U8224 ( .A(n7357), .ZN(n7356) );
  OAI21_X1 U8225 ( .B1(n12356), .B2(n7358), .A(n9004), .ZN(n7357) );
  INV_X1 U8226 ( .A(n9003), .ZN(n7358) );
  OR2_X1 U8227 ( .A1(n11954), .A2(n9007), .ZN(n8872) );
  OR2_X1 U8228 ( .A1(n8591), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8606) );
  INV_X1 U8229 ( .A(n8996), .ZN(n7369) );
  INV_X1 U8230 ( .A(n8851), .ZN(n7364) );
  INV_X1 U8231 ( .A(n7363), .ZN(n7362) );
  OAI21_X1 U8232 ( .B1(n11356), .B2(n7364), .A(n8853), .ZN(n7363) );
  INV_X1 U8233 ( .A(n7380), .ZN(n7379) );
  OAI21_X1 U8234 ( .B1(n10945), .B2(n7381), .A(n10918), .ZN(n7380) );
  INV_X1 U8235 ( .A(n8826), .ZN(n7381) );
  NAND2_X1 U8236 ( .A1(n10949), .A2(n8990), .ZN(n14882) );
  NAND2_X1 U8237 ( .A1(n10647), .A2(n10646), .ZN(n7397) );
  AND3_X1 U8238 ( .A1(n8381), .A2(n8380), .A3(n8379), .ZN(n9072) );
  NAND2_X1 U8239 ( .A1(n8403), .A2(n14916), .ZN(n8802) );
  INV_X1 U8240 ( .A(n8295), .ZN(n7114) );
  NOR2_X1 U8241 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), .ZN(
        n8315) );
  INV_X1 U8242 ( .A(n7440), .ZN(n7438) );
  INV_X1 U8243 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n8308) );
  INV_X1 U8244 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7434) );
  NAND2_X1 U8245 ( .A1(n6596), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6595) );
  INV_X1 U8246 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8303) );
  INV_X1 U8247 ( .A(n8253), .ZN(n7104) );
  OAI21_X1 U8248 ( .B1(n8428), .B2(n7092), .A(n8446), .ZN(n7091) );
  INV_X1 U8249 ( .A(n7091), .ZN(n7089) );
  INV_X1 U8250 ( .A(n11412), .ZN(n7330) );
  OR2_X1 U8251 ( .A1(n12598), .A2(n12597), .ZN(n12599) );
  INV_X1 U8252 ( .A(n12534), .ZN(n6691) );
  XNOR2_X1 U8253 ( .A(n12604), .B(n10021), .ZN(n10026) );
  NOR2_X1 U8254 ( .A1(n7502), .A2(n7498), .ZN(n7493) );
  AND2_X1 U8255 ( .A1(n7160), .A2(n12940), .ZN(n7158) );
  INV_X1 U8256 ( .A(n8180), .ZN(n7558) );
  NOR2_X1 U8257 ( .A1(n11211), .A2(n11406), .ZN(n7015) );
  INV_X1 U8258 ( .A(n7922), .ZN(n7150) );
  INV_X1 U8259 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U8260 ( .A1(n12744), .A2(n14645), .ZN(n7785) );
  NAND2_X1 U8261 ( .A1(n9887), .A2(n9886), .ZN(n10655) );
  AND2_X1 U8262 ( .A1(n13036), .A2(n13041), .ZN(n13031) );
  INV_X1 U8263 ( .A(n7808), .ZN(n6680) );
  NOR2_X1 U8264 ( .A1(n7642), .A2(n6678), .ZN(n6677) );
  NOR2_X1 U8265 ( .A1(n7189), .A2(n13490), .ZN(n7188) );
  AOI21_X1 U8266 ( .B1(n13250), .B2(n6641), .A(n6640), .ZN(n6639) );
  INV_X1 U8267 ( .A(n14207), .ZN(n6640) );
  INV_X1 U8268 ( .A(n14232), .ZN(n6641) );
  NAND2_X1 U8269 ( .A1(n11742), .A2(n7273), .ZN(n7272) );
  NAND2_X1 U8270 ( .A1(n6881), .A2(n11721), .ZN(n6880) );
  NAND2_X1 U8271 ( .A1(n6541), .A2(n6878), .ZN(n6877) );
  NOR2_X1 U8272 ( .A1(n7172), .A2(n7173), .ZN(n6922) );
  INV_X1 U8273 ( .A(n7174), .ZN(n7173) );
  NOR2_X1 U8274 ( .A1(n6481), .A2(n7265), .ZN(n7263) );
  INV_X1 U8275 ( .A(n7268), .ZN(n7265) );
  NAND2_X1 U8276 ( .A1(n11567), .A2(n13662), .ZN(n13636) );
  NAND2_X1 U8277 ( .A1(n11514), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11559) );
  NAND2_X1 U8278 ( .A1(n6485), .A2(n13629), .ZN(n7203) );
  OR2_X1 U8279 ( .A1(n13629), .A2(n7202), .ZN(n7204) );
  INV_X1 U8280 ( .A(n14249), .ZN(n7202) );
  NOR2_X1 U8281 ( .A1(n7184), .A2(n11036), .ZN(n7183) );
  INV_X1 U8282 ( .A(n11000), .ZN(n7186) );
  NOR2_X1 U8283 ( .A1(n6962), .A2(n6963), .ZN(n6961) );
  INV_X1 U8284 ( .A(n10282), .ZN(n6963) );
  INV_X1 U8285 ( .A(n14385), .ZN(n6962) );
  NAND2_X1 U8286 ( .A1(n10281), .A2(n11757), .ZN(n10283) );
  NAND2_X1 U8287 ( .A1(n10245), .A2(n10244), .ZN(n10297) );
  NOR2_X1 U8288 ( .A1(n14411), .A2(n10243), .ZN(n10244) );
  NAND2_X1 U8289 ( .A1(n6923), .A2(n11450), .ZN(n14411) );
  INV_X1 U8290 ( .A(n14433), .ZN(n6923) );
  INV_X1 U8291 ( .A(n14404), .ZN(n14401) );
  INV_X1 U8292 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7580) );
  INV_X1 U8293 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7581) );
  NAND2_X1 U8294 ( .A1(n6573), .A2(n6477), .ZN(n7005) );
  INV_X1 U8295 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9566) );
  INV_X1 U8296 ( .A(n7994), .ZN(n7992) );
  NAND2_X1 U8297 ( .A1(n7629), .A2(SI_18_), .ZN(n7630) );
  INV_X1 U8298 ( .A(n7680), .ZN(n7237) );
  NOR2_X1 U8299 ( .A1(n7295), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n10476) );
  XNOR2_X1 U8300 ( .A(n7625), .B(SI_16_), .ZN(n7713) );
  XNOR2_X1 U8301 ( .A(n7616), .B(SI_12_), .ZN(n7923) );
  AOI21_X1 U8302 ( .B1(n6459), .B2(n7251), .A(n6571), .ZN(n7249) );
  AOI21_X1 U8303 ( .B1(n7897), .B2(n7253), .A(n7252), .ZN(n7251) );
  INV_X1 U8304 ( .A(n7613), .ZN(n7252) );
  INV_X1 U8305 ( .A(n7609), .ZN(n7253) );
  AND2_X1 U8306 ( .A1(n9669), .A2(n9668), .ZN(n9696) );
  INV_X1 U8307 ( .A(n7217), .ZN(n7792) );
  NAND2_X1 U8308 ( .A1(n14006), .A2(n14007), .ZN(n14008) );
  XNOR2_X1 U8309 ( .A(n14008), .B(n6819), .ZN(n14055) );
  INV_X1 U8310 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6819) );
  AOI22_X1 U8311 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14012), .B1(n14061), .B2(
        n14011), .ZN(n14013) );
  NOR2_X1 U8312 ( .A1(n9144), .A2(n9145), .ZN(n7047) );
  NAND2_X1 U8313 ( .A1(n7040), .A2(n7039), .ZN(n7035) );
  NAND2_X1 U8314 ( .A1(n8337), .A2(n8336), .ZN(n8678) );
  INV_X1 U8315 ( .A(n8666), .ZN(n8337) );
  OR2_X1 U8316 ( .A1(n9122), .A2(n11911), .ZN(n11849) );
  NOR2_X1 U8317 ( .A1(n9108), .A2(n12368), .ZN(n7053) );
  NAND2_X1 U8318 ( .A1(n9128), .A2(n9129), .ZN(n11899) );
  AND2_X1 U8319 ( .A1(n11873), .A2(n9135), .ZN(n11900) );
  OR2_X1 U8320 ( .A1(n8707), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8718) );
  NAND2_X1 U8321 ( .A1(n6622), .A2(n10690), .ZN(n10689) );
  NAND2_X1 U8322 ( .A1(n8329), .A2(n11302), .ZN(n8518) );
  INV_X1 U8323 ( .A(n8504), .ZN(n8329) );
  NAND2_X1 U8324 ( .A1(n8335), .A2(n8334), .ZN(n8651) );
  INV_X1 U8325 ( .A(n8637), .ZN(n8335) );
  OR2_X1 U8326 ( .A1(n8651), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8666) );
  NOR2_X1 U8327 ( .A1(n9177), .A2(n9166), .ZN(n11974) );
  INV_X1 U8328 ( .A(n12177), .ZN(n9048) );
  AOI21_X1 U8329 ( .B1(n6605), .B2(n6502), .A(n8925), .ZN(n6604) );
  AND2_X1 U8330 ( .A1(n8784), .A2(n8367), .ZN(n8785) );
  AOI21_X1 U8331 ( .B1(n10142), .B2(n10141), .A(n10307), .ZN(n10143) );
  OR2_X1 U8332 ( .A1(n14752), .A2(n10852), .ZN(n7146) );
  AOI21_X1 U8333 ( .B1(n14772), .B2(n14771), .A(n14770), .ZN(n14789) );
  NAND2_X1 U8334 ( .A1(n14796), .A2(n10843), .ZN(n14814) );
  NAND2_X1 U8335 ( .A1(n10899), .A2(n7154), .ZN(n7151) );
  NAND2_X1 U8336 ( .A1(n7154), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7153) );
  OR2_X1 U8337 ( .A1(n14786), .A2(n10862), .ZN(n7156) );
  NAND2_X1 U8338 ( .A1(n14826), .A2(n10845), .ZN(n14852) );
  AOI21_X1 U8339 ( .B1(n14844), .B2(n14843), .A(n14842), .ZN(n14862) );
  NOR2_X1 U8340 ( .A1(n11098), .A2(n10907), .ZN(n6763) );
  XNOR2_X1 U8341 ( .A(n12017), .B(n12007), .ZN(n11099) );
  NAND2_X1 U8342 ( .A1(n11099), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n12019) );
  NAND2_X1 U8343 ( .A1(n12057), .A2(n12056), .ZN(n12059) );
  XNOR2_X1 U8344 ( .A(n12163), .B(n6811), .ZN(n12153) );
  NAND2_X1 U8345 ( .A1(n7385), .A2(n7383), .ZN(n12198) );
  AOI21_X1 U8346 ( .B1(n7386), .B2(n7387), .A(n7384), .ZN(n7383) );
  AND2_X1 U8347 ( .A1(n8748), .A2(n8747), .ZN(n12215) );
  NOR2_X1 U8348 ( .A1(n9015), .A2(n7392), .ZN(n7391) );
  INV_X1 U8349 ( .A(n7568), .ZN(n7392) );
  AOI21_X1 U8350 ( .B1(n12207), .B2(n8756), .A(n8773), .ZN(n12214) );
  INV_X1 U8351 ( .A(n9016), .ZN(n12217) );
  NAND2_X1 U8352 ( .A1(n8339), .A2(n11904), .ZN(n8728) );
  INV_X1 U8353 ( .A(n8718), .ZN(n8339) );
  NAND2_X1 U8354 ( .A1(n8340), .A2(n15102), .ZN(n8741) );
  INV_X1 U8355 ( .A(n8728), .ZN(n8340) );
  AOI21_X1 U8356 ( .B1(n9013), .B2(n7566), .A(n7565), .ZN(n12264) );
  NAND2_X1 U8357 ( .A1(n9010), .A2(n9009), .ZN(n12292) );
  AOI21_X1 U8358 ( .B1(n7373), .B2(n7375), .A(n7371), .ZN(n7370) );
  INV_X1 U8359 ( .A(n8865), .ZN(n7371) );
  AND4_X1 U8360 ( .A1(n8644), .A2(n8643), .A3(n8642), .A4(n8641), .ZN(n12358)
         );
  NAND2_X1 U8361 ( .A1(n8331), .A2(n8330), .ZN(n8577) );
  INV_X1 U8362 ( .A(n8553), .ZN(n8331) );
  AND3_X1 U8363 ( .A1(n8552), .A2(n8551), .A3(n8550), .ZN(n11381) );
  OR2_X1 U8364 ( .A1(n8518), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8536) );
  OR2_X1 U8365 ( .A1(n8536), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8553) );
  INV_X1 U8366 ( .A(n7413), .ZN(n7412) );
  AOI21_X1 U8367 ( .B1(n7413), .B2(n7411), .A(n7410), .ZN(n7409) );
  NOR2_X1 U8368 ( .A1(n11247), .A2(n6461), .ZN(n7413) );
  NAND2_X1 U8369 ( .A1(n11248), .A2(n11247), .ZN(n11246) );
  OR2_X1 U8370 ( .A1(n8483), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8504) );
  NAND2_X1 U8371 ( .A1(n8328), .A2(n8327), .ZN(n8483) );
  INV_X1 U8372 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n8327) );
  INV_X1 U8373 ( .A(n8466), .ZN(n8328) );
  NAND2_X1 U8374 ( .A1(n7397), .A2(n7396), .ZN(n10952) );
  AND2_X1 U8375 ( .A1(n8988), .A2(n8987), .ZN(n7396) );
  AND4_X1 U8376 ( .A1(n8445), .A2(n8444), .A3(n8443), .A4(n8442), .ZN(n10948)
         );
  NAND2_X1 U8377 ( .A1(n8326), .A2(n8325), .ZN(n8453) );
  INV_X1 U8378 ( .A(n8439), .ZN(n8326) );
  NAND2_X1 U8379 ( .A1(n10642), .A2(n10692), .ZN(n8439) );
  INV_X1 U8380 ( .A(n10646), .ZN(n10644) );
  OR2_X1 U8381 ( .A1(n8411), .A2(SI_3_), .ZN(n8420) );
  INV_X1 U8382 ( .A(n9072), .ZN(n14910) );
  NAND2_X1 U8383 ( .A1(n8802), .A2(n9067), .ZN(n8982) );
  AND2_X1 U8384 ( .A1(n9517), .A2(n12513), .ZN(n9175) );
  OR2_X1 U8385 ( .A1(n6787), .A2(n10802), .ZN(n8716) );
  NAND2_X1 U8386 ( .A1(n7111), .A2(n7112), .ZN(n8776) );
  AOI21_X1 U8387 ( .B1(n7113), .B2(n8294), .A(n6584), .ZN(n7112) );
  NAND2_X1 U8388 ( .A1(n8288), .A2(n15035), .ZN(n7095) );
  XNOR2_X1 U8389 ( .A(n8794), .B(P3_IR_REG_21__SCAN_IN), .ZN(n10628) );
  INV_X1 U8390 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7026) );
  NAND2_X1 U8391 ( .A1(n8661), .A2(n7026), .ZN(n7025) );
  XNOR2_X1 U8392 ( .A(n8661), .B(n7027), .ZN(n7023) );
  AND2_X1 U8393 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7024) );
  NAND2_X1 U8394 ( .A1(n6608), .A2(n8273), .ZN(n8646) );
  NAND2_X1 U8395 ( .A1(n8633), .A2(n8272), .ZN(n6608) );
  NAND2_X1 U8396 ( .A1(n8601), .A2(n8268), .ZN(n8614) );
  NAND2_X1 U8397 ( .A1(n8587), .A2(n8266), .ZN(n8599) );
  NAND2_X1 U8398 ( .A1(n7083), .A2(n7086), .ZN(n8585) );
  AND2_X1 U8399 ( .A1(n8266), .A2(n8265), .ZN(n8584) );
  NAND2_X1 U8400 ( .A1(n8546), .A2(n8261), .ZN(n8561) );
  AND2_X1 U8401 ( .A1(n8263), .A2(n8262), .ZN(n8560) );
  NAND2_X1 U8402 ( .A1(n8528), .A2(n8259), .ZN(n8544) );
  AND2_X1 U8403 ( .A1(n8261), .A2(n8260), .ZN(n8543) );
  AND2_X1 U8404 ( .A1(n8259), .A2(n8258), .ZN(n8525) );
  OAI21_X1 U8405 ( .B1(n8474), .B2(n7105), .A(n7102), .ZN(n8511) );
  AOI21_X1 U8406 ( .B1(n7106), .B2(n7104), .A(n7103), .ZN(n7102) );
  INV_X1 U8407 ( .A(n7106), .ZN(n7105) );
  INV_X1 U8408 ( .A(n8255), .ZN(n7103) );
  AND2_X1 U8409 ( .A1(n8257), .A2(n8256), .ZN(n8510) );
  OR2_X1 U8410 ( .A1(n8490), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n8491) );
  NOR2_X1 U8411 ( .A1(n8491), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8530) );
  INV_X1 U8412 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8477) );
  NAND2_X1 U8413 ( .A1(n6597), .A2(n7087), .ZN(n8463) );
  INV_X1 U8414 ( .A(n7088), .ZN(n7087) );
  NAND2_X1 U8415 ( .A1(n8429), .A2(n7089), .ZN(n6597) );
  OAI21_X1 U8416 ( .B1(n7091), .B2(n8246), .A(n8248), .ZN(n7088) );
  AND2_X1 U8417 ( .A1(n8244), .A2(n8243), .ZN(n8412) );
  NAND2_X1 U8418 ( .A1(n6610), .A2(n8399), .ZN(n6609) );
  AND2_X1 U8419 ( .A1(n8241), .A2(n8240), .ZN(n8373) );
  OR2_X1 U8420 ( .A1(n7853), .A2(n10525), .ZN(n7873) );
  NOR2_X1 U8421 ( .A1(n12600), .A2(n7345), .ZN(n7344) );
  INV_X1 U8422 ( .A(n12575), .ZN(n7345) );
  INV_X1 U8423 ( .A(n11281), .ZN(n7333) );
  AND2_X1 U8424 ( .A1(n11285), .A2(n7333), .ZN(n7332) );
  INV_X1 U8425 ( .A(n8015), .ZN(n8013) );
  AOI21_X1 U8426 ( .B1(n12673), .B2(n12672), .A(n12560), .ZN(n12564) );
  OR2_X1 U8427 ( .A1(n7873), .A2(n7872), .ZN(n7889) );
  INV_X1 U8428 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7888) );
  OAI21_X1 U8429 ( .B1(n12644), .B2(n7306), .A(n7304), .ZN(n12664) );
  AOI21_X1 U8430 ( .B1(n7307), .B2(n7305), .A(n12549), .ZN(n7304) );
  INV_X1 U8431 ( .A(n7309), .ZN(n7305) );
  OR2_X1 U8432 ( .A1(n7332), .A2(n11311), .ZN(n7331) );
  OR2_X1 U8433 ( .A1(n7889), .A2(n7888), .ZN(n7915) );
  AND2_X1 U8434 ( .A1(n12627), .A2(n6700), .ZN(n6699) );
  NAND2_X1 U8435 ( .A1(n6701), .A2(n12568), .ZN(n6700) );
  INV_X1 U8436 ( .A(n12654), .ZN(n6701) );
  INV_X1 U8437 ( .A(n12568), .ZN(n6702) );
  NAND2_X1 U8438 ( .A1(n7664), .A2(n7663), .ZN(n7954) );
  AND2_X1 U8439 ( .A1(n8193), .A2(n9952), .ZN(n9958) );
  NOR2_X1 U8440 ( .A1(n14633), .A2(n9951), .ZN(n9961) );
  NAND2_X1 U8441 ( .A1(n6830), .A2(n6719), .ZN(n6718) );
  AND2_X1 U8442 ( .A1(n9328), .A2(n6553), .ZN(n6830) );
  NAND2_X1 U8443 ( .A1(n6789), .A2(n6788), .ZN(n9350) );
  NAND2_X1 U8444 ( .A1(n9349), .A2(n9348), .ZN(n6788) );
  INV_X1 U8445 ( .A(n9186), .ZN(n10020) );
  AND3_X1 U8446 ( .A1(n7679), .A2(n7678), .A3(n7677), .ZN(n12697) );
  AND2_X1 U8447 ( .A1(n7770), .A2(n6771), .ZN(n7771) );
  OR2_X1 U8448 ( .A1(n7762), .A2(n9422), .ZN(n7770) );
  AND2_X1 U8449 ( .A1(n7769), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6737) );
  OR2_X1 U8450 ( .A1(n7763), .A2(n12760), .ZN(n7772) );
  OR2_X1 U8451 ( .A1(n9969), .A2(n9970), .ZN(n9967) );
  INV_X1 U8452 ( .A(n8116), .ZN(n7129) );
  INV_X1 U8453 ( .A(n7128), .ZN(n7125) );
  AND2_X1 U8454 ( .A1(n8108), .A2(n8107), .ZN(n12875) );
  NAND2_X1 U8455 ( .A1(n8116), .A2(n8115), .ZN(n12879) );
  AND2_X1 U8456 ( .A1(n8071), .A2(n8087), .ZN(n12907) );
  NAND2_X1 U8457 ( .A1(n7007), .A2(n12939), .ZN(n12934) );
  NAND2_X1 U8458 ( .A1(n13000), .A2(n13001), .ZN(n12999) );
  OR2_X1 U8459 ( .A1(n7709), .A2(n7668), .ZN(n7970) );
  NAND2_X1 U8460 ( .A1(n6833), .A2(n6506), .ZN(n13012) );
  NAND2_X1 U8461 ( .A1(n13027), .A2(n6834), .ZN(n6833) );
  NAND2_X1 U8462 ( .A1(n13036), .A2(n12728), .ZN(n6834) );
  NAND2_X1 U8463 ( .A1(n13054), .A2(n7135), .ZN(n6685) );
  NAND2_X1 U8464 ( .A1(n13074), .A2(n7136), .ZN(n7135) );
  NAND2_X1 U8465 ( .A1(n6441), .A2(n13074), .ZN(n13067) );
  AND3_X1 U8466 ( .A1(n7712), .A2(n7711), .A3(n7710), .ZN(n13058) );
  NAND2_X1 U8467 ( .A1(n7015), .A2(n7014), .ZN(n13069) );
  OAI21_X1 U8468 ( .B1(n7960), .B2(n11406), .A(n11315), .ZN(n7961) );
  INV_X1 U8469 ( .A(n7015), .ZN(n11390) );
  AND4_X1 U8470 ( .A1(n7935), .A2(n7934), .A3(n7933), .A4(n7932), .ZN(n11317)
         );
  AND2_X1 U8471 ( .A1(n7944), .A2(n7943), .ZN(n11314) );
  OR2_X1 U8472 ( .A1(n7930), .A2(n9971), .ZN(n7952) );
  NOR2_X1 U8473 ( .A1(n10776), .A2(n10769), .ZN(n6672) );
  INV_X1 U8474 ( .A(n10748), .ZN(n6803) );
  NAND2_X1 U8475 ( .A1(n6684), .A2(n7117), .ZN(n10737) );
  NAND2_X1 U8476 ( .A1(n6683), .A2(n6684), .ZN(n10739) );
  AND2_X1 U8477 ( .A1(n7895), .A2(n7117), .ZN(n6683) );
  AND2_X1 U8478 ( .A1(n10469), .A2(n14676), .ZN(n10456) );
  AND2_X1 U8479 ( .A1(n7008), .A2(n10469), .ZN(n10727) );
  CLKBUF_X1 U8480 ( .A(n10452), .Z(n6783) );
  NAND2_X1 U8481 ( .A1(n7541), .A2(n7540), .ZN(n10435) );
  INV_X1 U8482 ( .A(n7543), .ZN(n7542) );
  AOI21_X1 U8483 ( .B1(n7826), .B2(n6675), .A(n6498), .ZN(n6674) );
  INV_X1 U8484 ( .A(n7826), .ZN(n6676) );
  INV_X1 U8485 ( .A(n7813), .ZN(n6675) );
  XNOR2_X1 U8486 ( .A(n7841), .B(n12740), .ZN(n10437) );
  NAND2_X1 U8487 ( .A1(n7659), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7835) );
  NAND2_X1 U8488 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7820) );
  NAND2_X1 U8489 ( .A1(n14645), .A2(n10664), .ZN(n10663) );
  NOR2_X1 U8490 ( .A1(n10021), .A2(n10515), .ZN(n10664) );
  NAND2_X1 U8491 ( .A1(n7012), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7011) );
  NAND2_X1 U8492 ( .A1(n8121), .A2(n8120), .ZN(n12858) );
  AND2_X1 U8493 ( .A1(n7163), .A2(n6483), .ZN(n12947) );
  AND2_X1 U8494 ( .A1(n14689), .A2(n14688), .ZN(n14655) );
  OR2_X1 U8495 ( .A1(n8221), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8207) );
  NOR2_X1 U8496 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n7297) );
  OR2_X1 U8497 ( .A1(n7884), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n7910) );
  AND2_X1 U8498 ( .A1(n7869), .A2(n7884), .ZN(n12824) );
  INV_X1 U8499 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7634) );
  INV_X1 U8500 ( .A(n11341), .ZN(n6637) );
  INV_X1 U8501 ( .A(n13478), .ZN(n11346) );
  NOR2_X1 U8502 ( .A1(n13378), .A2(n7477), .ZN(n7476) );
  INV_X1 U8503 ( .A(n13281), .ZN(n7477) );
  AND2_X1 U8504 ( .A1(n13327), .A2(n13325), .ZN(n13397) );
  OR2_X1 U8505 ( .A1(n10399), .A2(n10398), .ZN(n10551) );
  OAI21_X1 U8506 ( .B1(n11062), .B2(n7450), .A(n7447), .ZN(n11339) );
  INV_X1 U8507 ( .A(n6761), .ZN(n7448) );
  NOR2_X1 U8508 ( .A1(n10563), .A2(n10562), .ZN(n10986) );
  OR2_X1 U8509 ( .A1(n10551), .A2(n10550), .ZN(n10563) );
  NAND2_X1 U8510 ( .A1(n7472), .A2(n7471), .ZN(n7470) );
  INV_X1 U8511 ( .A(n13409), .ZN(n7472) );
  NOR2_X1 U8512 ( .A1(n11041), .A2(n11040), .ZN(n11223) );
  AND4_X1 U8513 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n13651) );
  AND4_X1 U8514 ( .A1(n11048), .A2(n11047), .A3(n11046), .A4(n11045), .ZN(
        n13236) );
  CLKBUF_X1 U8515 ( .A(n10100), .Z(n11044) );
  NOR2_X1 U8516 ( .A1(n6944), .A2(n13648), .ZN(n6942) );
  NOR2_X1 U8517 ( .A1(n13721), .A2(n7176), .ZN(n7175) );
  INV_X1 U8518 ( .A(n13649), .ZN(n7176) );
  NOR2_X1 U8519 ( .A1(n7260), .A2(n6987), .ZN(n6985) );
  INV_X1 U8520 ( .A(n6481), .ZN(n7172) );
  OAI21_X1 U8521 ( .B1(n7242), .B2(n7241), .A(n7239), .ZN(n13755) );
  NAND2_X1 U8522 ( .A1(n13787), .A2(n6456), .ZN(n13762) );
  NAND2_X1 U8523 ( .A1(n13787), .A2(n13931), .ZN(n13774) );
  INV_X1 U8524 ( .A(n6939), .ZN(n13820) );
  NOR2_X1 U8525 ( .A1(n11575), .A2(n13428), .ZN(n11590) );
  NAND2_X1 U8526 ( .A1(n6941), .A2(n6940), .ZN(n13832) );
  INV_X1 U8527 ( .A(n6941), .ZN(n13856) );
  NOR2_X1 U8528 ( .A1(n13860), .A2(n13864), .ZN(n6746) );
  NAND2_X1 U8529 ( .A1(n14257), .A2(n13864), .ZN(n7198) );
  NAND2_X1 U8530 ( .A1(n13635), .A2(n7196), .ZN(n7195) );
  OAI21_X1 U8531 ( .B1(n13860), .B2(n7197), .A(n6534), .ZN(n7196) );
  INV_X1 U8532 ( .A(n13636), .ZN(n13830) );
  NOR2_X1 U8533 ( .A1(n14251), .A2(n14271), .ZN(n14250) );
  NAND2_X1 U8534 ( .A1(n6442), .A2(n6931), .ZN(n14251) );
  NAND2_X1 U8535 ( .A1(n6933), .A2(n6932), .ZN(n11233) );
  INV_X1 U8536 ( .A(n11187), .ZN(n6933) );
  NAND2_X1 U8537 ( .A1(n11175), .A2(n11769), .ZN(n6984) );
  NAND2_X1 U8538 ( .A1(n6935), .A2(n6934), .ZN(n11187) );
  INV_X1 U8539 ( .A(n14123), .ZN(n6935) );
  NAND2_X1 U8540 ( .A1(n6937), .A2(n6936), .ZN(n14123) );
  AND2_X1 U8541 ( .A1(n6965), .A2(n10539), .ZN(n6964) );
  AOI21_X1 U8542 ( .B1(n11762), .B2(n7193), .A(n6522), .ZN(n7192) );
  NAND2_X1 U8543 ( .A1(n10286), .A2(n11763), .ZN(n10388) );
  AOI21_X1 U8544 ( .B1(n11761), .B2(n7180), .A(n6524), .ZN(n7179) );
  INV_X1 U8545 ( .A(n10251), .ZN(n7180) );
  NAND2_X1 U8546 ( .A1(n10283), .A2(n10282), .ZN(n10337) );
  NAND2_X1 U8547 ( .A1(n10337), .A2(n7181), .ZN(n14386) );
  NAND2_X1 U8548 ( .A1(n11448), .A2(n11447), .ZN(n14404) );
  NAND2_X1 U8549 ( .A1(n14423), .A2(n11441), .ZN(n14422) );
  NAND2_X1 U8550 ( .A1(n10231), .A2(n10230), .ZN(n14423) );
  NAND2_X1 U8551 ( .A1(n9925), .A2(n10329), .ZN(n14433) );
  NAND2_X1 U8552 ( .A1(n9861), .A2(n6972), .ZN(n11437) );
  NAND2_X1 U8553 ( .A1(n11718), .A2(n11717), .ZN(n13890) );
  NAND2_X1 U8554 ( .A1(n13630), .A2(n13629), .ZN(n14248) );
  AND2_X1 U8555 ( .A1(n9726), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9678) );
  XNOR2_X1 U8556 ( .A(n9294), .B(n9293), .ZN(n11716) );
  XNOR2_X1 U8557 ( .A(n8118), .B(n8117), .ZN(n13192) );
  NAND2_X1 U8558 ( .A1(n7200), .A2(n7199), .ZN(n6655) );
  NAND2_X1 U8559 ( .A1(n8050), .A2(n8049), .ZN(n8063) );
  XNOR2_X1 U8560 ( .A(n8027), .B(SI_22_), .ZN(n11610) );
  NOR2_X1 U8561 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n9569) );
  INV_X1 U8562 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n15080) );
  NAND2_X1 U8563 ( .A1(n6794), .A2(n6792), .ZN(n6740) );
  NAND2_X1 U8564 ( .A1(n7726), .A2(n6793), .ZN(n6792) );
  AND2_X1 U8565 ( .A1(n10077), .A2(n9990), .ZN(n11025) );
  OR2_X1 U8566 ( .A1(n9700), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9702) );
  OR2_X1 U8567 ( .A1(n9702), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9746) );
  NOR2_X1 U8568 ( .A1(n9690), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9669) );
  OR2_X1 U8569 ( .A1(n9688), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9690) );
  NAND2_X1 U8570 ( .A1(n7018), .A2(n7016), .ZN(n14043) );
  NAND2_X1 U8571 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7017), .ZN(n7016) );
  INV_X1 U8572 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7017) );
  XNOR2_X1 U8573 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n14042) );
  XNOR2_X1 U8574 ( .A(n14002), .B(n7079), .ZN(n14050) );
  INV_X1 U8575 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14051) );
  NAND2_X1 U8576 ( .A1(n14106), .A2(n14105), .ZN(n7073) );
  OAI21_X1 U8577 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14020), .A(n14019), .ZN(
        n14035) );
  AOI21_X1 U8578 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14024), .A(n14023), .ZN(
        n14033) );
  NOR2_X1 U8579 ( .A1(n14080), .A2(n14079), .ZN(n14023) );
  AND3_X1 U8580 ( .A1(n8482), .A2(n8481), .A3(n8480), .ZN(n14961) );
  INV_X1 U8581 ( .A(n11363), .ZN(n6846) );
  AND3_X1 U8582 ( .A1(n8534), .A2(n8533), .A3(n8532), .ZN(n11370) );
  AND2_X1 U8583 ( .A1(n7035), .A2(n7034), .ZN(n10637) );
  INV_X1 U8584 ( .A(n7031), .ZN(n7034) );
  NAND2_X1 U8585 ( .A1(n7035), .A2(n7038), .ZN(n10638) );
  INV_X1 U8586 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10642) );
  NAND2_X1 U8587 ( .A1(n6614), .A2(n9115), .ZN(n11842) );
  NAND2_X1 U8588 ( .A1(n6619), .A2(n7048), .ZN(n6618) );
  NOR2_X1 U8589 ( .A1(n9144), .A2(n6616), .ZN(n6615) );
  INV_X1 U8590 ( .A(n9142), .ZN(n6616) );
  AND2_X1 U8591 ( .A1(n11816), .A2(n6832), .ZN(n6831) );
  AND2_X1 U8592 ( .A1(n11812), .A2(n11963), .ZN(n6832) );
  NAND2_X1 U8593 ( .A1(n10978), .A2(n9083), .ZN(n11167) );
  NAND2_X1 U8594 ( .A1(n7064), .A2(n11996), .ZN(n7067) );
  INV_X1 U8595 ( .A(n7068), .ZN(n7064) );
  NAND2_X1 U8596 ( .A1(n8687), .A2(n8686), .ZN(n12298) );
  OR2_X1 U8597 ( .A1(n6787), .A2(n10194), .ZN(n8686) );
  OAI21_X1 U8598 ( .B1(n11886), .B2(n9109), .A(n7050), .ZN(n11893) );
  INV_X1 U8599 ( .A(n7053), .ZN(n7050) );
  AND3_X1 U8600 ( .A1(n8436), .A2(n8435), .A3(n8434), .ZN(n10695) );
  NAND2_X1 U8601 ( .A1(n11165), .A2(n9085), .ZN(n11300) );
  INV_X1 U8602 ( .A(n7063), .ZN(n7060) );
  NAND2_X1 U8603 ( .A1(n7062), .A2(n7063), .ZN(n11931) );
  NAND2_X1 U8604 ( .A1(n6607), .A2(n8696), .ZN(n12286) );
  AND4_X1 U8605 ( .A1(n8542), .A2(n8541), .A3(n8540), .A4(n8539), .ZN(n11945)
         );
  XNOR2_X1 U8606 ( .A(n9073), .B(n10708), .ZN(n10358) );
  NAND2_X1 U8607 ( .A1(n9161), .A2(n9160), .ZN(n11972) );
  AOI21_X1 U8608 ( .B1(n10805), .B2(n10806), .A(n6773), .ZN(n10830) );
  AND2_X1 U8609 ( .A1(n9078), .A2(n10948), .ZN(n6773) );
  INV_X1 U8610 ( .A(n11968), .ZN(n11979) );
  INV_X1 U8611 ( .A(n11963), .ZN(n11981) );
  INV_X1 U8612 ( .A(n12226), .ZN(n12201) );
  INV_X1 U8613 ( .A(n12215), .ZN(n12236) );
  OAI211_X1 U8614 ( .C1(n8772), .C2(n12430), .A(n8691), .B(n8690), .ZN(n12306)
         );
  INV_X1 U8615 ( .A(n12358), .ZN(n11952) );
  NAND4_X1 U8616 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8580), .ZN(n11920)
         );
  INV_X1 U8617 ( .A(n11945), .ZN(n11866) );
  INV_X1 U8618 ( .A(n11303), .ZN(n11991) );
  INV_X1 U8619 ( .A(n10920), .ZN(n11993) );
  INV_X1 U8620 ( .A(n10948), .ZN(n10832) );
  OR2_X1 U8621 ( .A1(n9517), .A2(n11423), .ZN(n11997) );
  INV_X1 U8622 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14750) );
  NOR2_X1 U8623 ( .A1(n10135), .A2(n14746), .ZN(n14744) );
  INV_X1 U8624 ( .A(n7146), .ZN(n14751) );
  NAND2_X1 U8625 ( .A1(n10894), .A2(n7147), .ZN(n7142) );
  NAND2_X1 U8626 ( .A1(n7147), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7144) );
  INV_X1 U8627 ( .A(n10894), .ZN(n7145) );
  NAND2_X1 U8628 ( .A1(n7152), .A2(n7151), .ZN(n14802) );
  NOR2_X1 U8629 ( .A1(n14858), .A2(n11272), .ZN(n14857) );
  AND2_X1 U8630 ( .A1(n10847), .A2(n14872), .ZN(n10848) );
  XNOR2_X1 U8631 ( .A(n12054), .B(n12061), .ZN(n12034) );
  NAND2_X1 U8632 ( .A1(n12034), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n12056) );
  AND2_X1 U8633 ( .A1(n12030), .A2(n12029), .ZN(n12048) );
  NOR2_X1 U8634 ( .A1(n7139), .A2(n12089), .ZN(n7138) );
  INV_X1 U8635 ( .A(n7141), .ZN(n7139) );
  NAND2_X1 U8636 ( .A1(n12109), .A2(n12110), .ZN(n12138) );
  NOR2_X1 U8637 ( .A1(n14147), .A2(n6520), .ZN(n12133) );
  NAND2_X1 U8638 ( .A1(n8362), .A2(n8361), .ZN(n12181) );
  NAND2_X1 U8639 ( .A1(n12234), .A2(n7568), .ZN(n12224) );
  NAND2_X1 U8640 ( .A1(n7422), .A2(n7423), .ZN(n12246) );
  NAND2_X1 U8641 ( .A1(n7382), .A2(n8929), .ZN(n12310) );
  NAND2_X1 U8642 ( .A1(n12328), .A2(n7416), .ZN(n12318) );
  NAND2_X1 U8643 ( .A1(n8636), .A2(n8635), .ZN(n12444) );
  NAND2_X1 U8644 ( .A1(n7355), .A2(n9003), .ZN(n12343) );
  NAND2_X1 U8645 ( .A1(n12355), .A2(n12356), .ZN(n7355) );
  NAND2_X1 U8646 ( .A1(n12375), .A2(n8861), .ZN(n12360) );
  NAND2_X1 U8647 ( .A1(n8605), .A2(n8604), .ZN(n12452) );
  NAND2_X1 U8648 ( .A1(n11359), .A2(n8851), .ZN(n11401) );
  NAND2_X1 U8649 ( .A1(n11351), .A2(n8996), .ZN(n11398) );
  NAND2_X1 U8650 ( .A1(n11244), .A2(n11243), .ZN(n12393) );
  NAND2_X1 U8651 ( .A1(n7405), .A2(n7403), .ZN(n11157) );
  AND3_X1 U8652 ( .A1(n8517), .A2(n8516), .A3(n8515), .ZN(n11276) );
  NAND2_X1 U8653 ( .A1(n10944), .A2(n8826), .ZN(n10917) );
  INV_X1 U8654 ( .A(n14929), .ZN(n12271) );
  NAND2_X1 U8655 ( .A1(n14896), .A2(n14960), .ZN(n12391) );
  INV_X2 U8656 ( .A(n14933), .ZN(n14935) );
  INV_X1 U8657 ( .A(n12181), .ZN(n12462) );
  NAND2_X1 U8658 ( .A1(n8324), .A2(n8323), .ZN(n12463) );
  INV_X1 U8659 ( .A(n11819), .ZN(n12471) );
  OR2_X1 U8660 ( .A1(n12424), .A2(n12423), .ZN(n12484) );
  NAND2_X1 U8661 ( .A1(n8665), .A2(n8664), .ZN(n12496) );
  INV_X1 U8662 ( .A(n11276), .ZN(n11306) );
  INV_X1 U8663 ( .A(n9147), .ZN(n12514) );
  AND2_X1 U8664 ( .A1(n7439), .A2(n7437), .ZN(n7436) );
  INV_X1 U8665 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7437) );
  OAI21_X1 U8666 ( .B1(n8751), .B2(n8294), .A(n8295), .ZN(n8764) );
  XNOR2_X1 U8667 ( .A(n8961), .B(n8312), .ZN(n11201) );
  OAI21_X1 U8668 ( .B1(n8715), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n8287), .ZN(
        n8725) );
  XNOR2_X1 U8669 ( .A(n8715), .B(n15035), .ZN(n10801) );
  NOR2_X1 U8670 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), .ZN(
        n8957) );
  NAND2_X1 U8671 ( .A1(n8792), .A2(n8793), .ZN(n10169) );
  NAND2_X1 U8672 ( .A1(n7082), .A2(n7086), .ZN(n8573) );
  NAND2_X1 U8673 ( .A1(n7084), .A2(n7086), .ZN(n8571) );
  NAND2_X1 U8674 ( .A1(n7101), .A2(n7106), .ZN(n8499) );
  NAND2_X1 U8675 ( .A1(n8474), .A2(n8253), .ZN(n7101) );
  NAND2_X1 U8676 ( .A1(n7090), .A2(n8246), .ZN(n8447) );
  NAND2_X1 U8677 ( .A1(n8429), .A2(n8428), .ZN(n7090) );
  OAI21_X1 U8678 ( .B1(n8396), .B2(n6856), .A(n6855), .ZN(n6854) );
  AND2_X1 U8679 ( .A1(n9945), .A2(n9401), .ZN(n9452) );
  NAND2_X1 U8680 ( .A1(n8086), .A2(n8085), .ZN(n13103) );
  NAND2_X1 U8681 ( .A1(n13195), .A2(n7682), .ZN(n8086) );
  XNOR2_X1 U8682 ( .A(n12564), .B(n12561), .ZN(n12583) );
  NAND2_X1 U8683 ( .A1(n10932), .A2(n10931), .ZN(n10934) );
  NAND2_X1 U8684 ( .A1(n10028), .A2(n6689), .ZN(n6688) );
  INV_X1 U8685 ( .A(n10029), .ZN(n6689) );
  INV_X1 U8686 ( .A(n7301), .ZN(n10042) );
  INV_X1 U8687 ( .A(n12744), .ZN(n10037) );
  NAND2_X1 U8688 ( .A1(n7308), .A2(n7307), .ZN(n12588) );
  AND2_X1 U8689 ( .A1(n7308), .A2(n6500), .ZN(n12590) );
  NAND2_X1 U8690 ( .A1(n12644), .A2(n7309), .ZN(n7308) );
  OR2_X1 U8691 ( .A1(n10588), .A2(n7315), .ZN(n10789) );
  NOR2_X1 U8692 ( .A1(n10588), .A2(n10587), .ZN(n10590) );
  AND4_X1 U8693 ( .A1(n7920), .A2(n7919), .A3(n7918), .A4(n7917), .ZN(n11288)
         );
  NAND2_X1 U8694 ( .A1(n6698), .A2(n12568), .ZN(n12626) );
  NAND2_X1 U8695 ( .A1(n12655), .A2(n12654), .ZN(n6698) );
  AND2_X1 U8696 ( .A1(n7325), .A2(n7326), .ZN(n12637) );
  OR2_X1 U8697 ( .A1(n7327), .A2(n7324), .ZN(n7326) );
  NAND2_X1 U8698 ( .A1(n12715), .A2(n12714), .ZN(n7325) );
  AND2_X1 U8699 ( .A1(n10040), .A2(n10043), .ZN(n7300) );
  NAND2_X1 U8700 ( .A1(n10534), .A2(n7314), .ZN(n7313) );
  OAI21_X1 U8701 ( .B1(n7315), .B2(n7312), .A(n7316), .ZN(n7311) );
  INV_X1 U8702 ( .A(n11314), .ZN(n11324) );
  INV_X1 U8703 ( .A(n13129), .ZN(n12679) );
  NAND2_X1 U8704 ( .A1(n11079), .A2(n6777), .ZN(n6776) );
  INV_X1 U8705 ( .A(n11081), .ZN(n6777) );
  NAND2_X1 U8706 ( .A1(n6668), .A2(n7912), .ZN(n11091) );
  NAND2_X1 U8707 ( .A1(n10995), .A2(n7682), .ZN(n6668) );
  AND2_X1 U8708 ( .A1(n12717), .A2(n13004), .ZN(n12685) );
  AND2_X1 U8709 ( .A1(n12644), .A2(n12543), .ZN(n12695) );
  INV_X1 U8710 ( .A(n12741), .ZN(n10438) );
  INV_X1 U8711 ( .A(n12683), .ZN(n12658) );
  NAND2_X1 U8712 ( .A1(n10205), .A2(n7560), .ZN(n10206) );
  INV_X1 U8713 ( .A(n12708), .ZN(n12720) );
  XNOR2_X1 U8714 ( .A(n7327), .B(n12535), .ZN(n12715) );
  INV_X1 U8715 ( .A(n12631), .ZN(n12917) );
  NAND2_X1 U8716 ( .A1(n8056), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7764) );
  OR2_X1 U8717 ( .A1(n7762), .A2(n7761), .ZN(n7767) );
  NAND2_X1 U8718 ( .A1(n6836), .A2(n6438), .ZN(n13091) );
  XNOR2_X1 U8719 ( .A(n12851), .B(n6837), .ZN(n6836) );
  INV_X1 U8720 ( .A(n12862), .ZN(n7550) );
  AOI21_X1 U8721 ( .B1(n7121), .B2(n6458), .A(n8151), .ZN(n7120) );
  INV_X1 U8722 ( .A(n12866), .ZN(n7121) );
  NAND2_X1 U8723 ( .A1(n12866), .A2(n7123), .ZN(n7122) );
  NOR2_X1 U8724 ( .A1(n7124), .A2(n13029), .ZN(n7123) );
  NOR2_X1 U8725 ( .A1(n7125), .A2(n7127), .ZN(n7124) );
  NOR2_X1 U8726 ( .A1(n8129), .A2(n7129), .ZN(n7127) );
  AND2_X1 U8727 ( .A1(n12874), .A2(n12873), .ZN(n13095) );
  NOR2_X1 U8728 ( .A1(n6682), .A2(n6667), .ZN(n6666) );
  AOI21_X1 U8729 ( .B1(n12891), .B2(n13065), .A(n12890), .ZN(n13105) );
  NAND2_X1 U8730 ( .A1(n12889), .A2(n12888), .ZN(n12890) );
  NAND2_X1 U8731 ( .A1(n12886), .A2(n7577), .ZN(n12891) );
  NAND2_X1 U8732 ( .A1(n7491), .A2(n7495), .ZN(n12910) );
  NAND2_X1 U8733 ( .A1(n12941), .A2(n7498), .ZN(n7491) );
  AND2_X1 U8734 ( .A1(n8067), .A2(n8066), .ZN(n12909) );
  AOI21_X1 U8735 ( .B1(n12903), .B2(n13065), .A(n12902), .ZN(n13110) );
  NAND2_X1 U8736 ( .A1(n7499), .A2(n7505), .ZN(n12925) );
  NAND2_X1 U8737 ( .A1(n7500), .A2(n12929), .ZN(n7499) );
  NAND2_X1 U8738 ( .A1(n7159), .A2(n7160), .ZN(n12930) );
  OR2_X1 U8739 ( .A1(n12959), .A2(n7161), .ZN(n7159) );
  NAND2_X1 U8740 ( .A1(n7530), .A2(n7531), .ZN(n12964) );
  NAND2_X1 U8741 ( .A1(n12992), .A2(n7533), .ZN(n7530) );
  INV_X1 U8742 ( .A(n12967), .ZN(n12979) );
  NAND2_X1 U8743 ( .A1(n7535), .A2(n7533), .ZN(n13136) );
  NAND2_X1 U8744 ( .A1(n7535), .A2(n7537), .ZN(n12987) );
  NAND2_X1 U8745 ( .A1(n11533), .A2(n7682), .ZN(n7658) );
  AND2_X1 U8746 ( .A1(n7702), .A2(n7701), .ZN(n13045) );
  NAND2_X1 U8747 ( .A1(n13062), .A2(n8180), .ZN(n13040) );
  NAND2_X1 U8748 ( .A1(n8179), .A2(n8178), .ZN(n13060) );
  INV_X1 U8749 ( .A(n7960), .ZN(n11207) );
  NAND2_X1 U8750 ( .A1(n10726), .A2(n8166), .ZN(n10745) );
  NAND2_X1 U8751 ( .A1(n8165), .A2(n8164), .ZN(n10724) );
  NAND2_X1 U8752 ( .A1(n10416), .A2(n8158), .ZN(n10462) );
  NAND2_X1 U8753 ( .A1(n10424), .A2(n7813), .ZN(n10464) );
  NAND2_X1 U8754 ( .A1(n10108), .A2(n7682), .ZN(n7796) );
  NAND2_X1 U8755 ( .A1(n13038), .A2(n10382), .ZN(n13073) );
  INV_X1 U8756 ( .A(n13073), .ZN(n13082) );
  INV_X1 U8757 ( .A(n13085), .ZN(n12984) );
  NAND2_X1 U8758 ( .A1(n13091), .A2(n6800), .ZN(n13171) );
  INV_X1 U8759 ( .A(n6801), .ZN(n6800) );
  OAI21_X1 U8760 ( .B1(n6837), .B2(n14715), .A(n13092), .ZN(n6801) );
  AND3_X2 U8761 ( .A1(n8230), .A2(n10368), .A3(n14636), .ZN(n14723) );
  AND2_X1 U8762 ( .A1(n9945), .A2(n8224), .ZN(n14637) );
  NAND2_X1 U8763 ( .A1(n6692), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U8764 ( .A1(n7646), .A2(n6460), .ZN(n6692) );
  XNOR2_X1 U8765 ( .A(n8216), .B(n8215), .ZN(n13203) );
  XNOR2_X1 U8766 ( .A(n8213), .B(n8212), .ZN(n11295) );
  NAND2_X1 U8767 ( .A1(n8138), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8140) );
  INV_X1 U8768 ( .A(n8193), .ZN(n11010) );
  INV_X1 U8769 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10585) );
  INV_X1 U8770 ( .A(n10418), .ZN(n10583) );
  INV_X1 U8771 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10178) );
  INV_X1 U8772 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10083) );
  INV_X1 U8773 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9924) );
  INV_X1 U8774 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9821) );
  INV_X1 U8775 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9757) );
  INV_X1 U8776 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9751) );
  INV_X1 U8777 ( .A(n9484), .ZN(n9749) );
  INV_X1 U8778 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9705) );
  INV_X1 U8779 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9683) );
  INV_X1 U8780 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9672) );
  INV_X1 U8781 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9663) );
  INV_X1 U8782 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9648) );
  INV_X1 U8783 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9646) );
  INV_X1 U8784 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9682) );
  NAND2_X1 U8785 ( .A1(n13346), .A2(n13344), .ZN(n6629) );
  CLKBUF_X1 U8786 ( .A(n13346), .Z(n13347) );
  INV_X1 U8787 ( .A(n10120), .ZN(n7458) );
  NAND2_X1 U8788 ( .A1(n10118), .A2(n10117), .ZN(n10119) );
  NAND2_X1 U8789 ( .A1(n7462), .A2(n7464), .ZN(n13356) );
  NAND2_X1 U8790 ( .A1(n13409), .A2(n7468), .ZN(n7462) );
  AOI21_X1 U8791 ( .B1(n7456), .B2(n13336), .A(n13362), .ZN(n7455) );
  XNOR2_X1 U8792 ( .A(n13369), .B(n13368), .ZN(n13370) );
  NAND2_X1 U8793 ( .A1(n7452), .A2(n7451), .ZN(n11261) );
  NAND2_X1 U8794 ( .A1(n11062), .A2(n11061), .ZN(n7452) );
  XNOR2_X1 U8795 ( .A(n10002), .B(n9927), .ZN(n9931) );
  NAND2_X1 U8796 ( .A1(n13282), .A2(n13281), .ZN(n13379) );
  NAND2_X1 U8797 ( .A1(n14222), .A2(n13221), .ZN(n13387) );
  NAND2_X1 U8798 ( .A1(n14222), .A2(n6492), .ZN(n13388) );
  NOR2_X1 U8799 ( .A1(n10501), .A2(n10491), .ZN(n10759) );
  AND2_X1 U8800 ( .A1(n10490), .A2(n10489), .ZN(n10491) );
  XNOR2_X1 U8801 ( .A(n11339), .B(n11340), .ZN(n6638) );
  NAND2_X1 U8802 ( .A1(n10544), .A2(n10543), .ZN(n14525) );
  AOI21_X1 U8803 ( .B1(n7464), .B2(n7467), .A(n6528), .ZN(n7463) );
  INV_X1 U8804 ( .A(n6644), .ZN(n6643) );
  OAI21_X1 U8805 ( .B1(n6492), .B2(n6645), .A(n13435), .ZN(n6644) );
  INV_X1 U8806 ( .A(n13230), .ZN(n6645) );
  NAND2_X1 U8807 ( .A1(n13388), .A2(n13230), .ZN(n13434) );
  NAND2_X1 U8808 ( .A1(n10001), .A2(n6828), .ZN(n10004) );
  NAND2_X1 U8809 ( .A1(n6829), .A2(n9927), .ZN(n6828) );
  INV_X1 U8810 ( .A(n10002), .ZN(n6829) );
  NAND2_X1 U8811 ( .A1(n7470), .A2(n13262), .ZN(n13451) );
  NAND2_X1 U8812 ( .A1(n6652), .A2(n6651), .ZN(n10818) );
  NAND2_X1 U8813 ( .A1(n10757), .A2(n10758), .ZN(n6651) );
  NAND2_X1 U8814 ( .A1(n10759), .A2(n6653), .ZN(n6652) );
  NAND2_X1 U8815 ( .A1(n6810), .A2(n6654), .ZN(n6653) );
  NOR2_X1 U8816 ( .A1(n11789), .A2(n7275), .ZN(n7274) );
  INV_X1 U8817 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n9711) );
  OR2_X1 U8818 ( .A1(n11730), .A2(n9733), .ZN(n9708) );
  OR2_X1 U8819 ( .A1(n11730), .A2(n9731), .ZN(n9583) );
  OR2_X1 U8820 ( .A1(n10100), .A2(n9559), .ZN(n6657) );
  OR2_X1 U8821 ( .A1(n11730), .A2(n9732), .ZN(n6656) );
  NAND2_X1 U8822 ( .A1(n15191), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6660) );
  INV_X1 U8823 ( .A(n6967), .ZN(n6966) );
  NAND2_X1 U8824 ( .A1(n7262), .A2(n6750), .ZN(n13914) );
  OR2_X1 U8825 ( .A1(n13736), .A2(n6751), .ZN(n6750) );
  OR2_X1 U8826 ( .A1(n7172), .A2(n7268), .ZN(n6751) );
  OR2_X1 U8827 ( .A1(n13739), .A2(n14382), .ZN(n6841) );
  NOR2_X1 U8828 ( .A1(n13747), .A2(n7213), .ZN(n7212) );
  INV_X1 U8829 ( .A(n13646), .ZN(n7213) );
  NAND2_X1 U8830 ( .A1(n13752), .A2(n13646), .ZN(n13748) );
  NAND2_X1 U8831 ( .A1(n13770), .A2(n13643), .ZN(n13754) );
  NAND2_X1 U8832 ( .A1(n11627), .A2(n11743), .ZN(n11629) );
  NAND2_X1 U8833 ( .A1(n7244), .A2(n7248), .ZN(n13786) );
  NAND2_X1 U8834 ( .A1(n13812), .A2(n13640), .ZN(n13806) );
  INV_X1 U8835 ( .A(n6805), .ZN(n13814) );
  NAND2_X1 U8836 ( .A1(n11581), .A2(n11580), .ZN(n13950) );
  NAND2_X1 U8837 ( .A1(n11579), .A2(n11743), .ZN(n11581) );
  NAND2_X1 U8838 ( .A1(n13635), .A2(n13634), .ZN(n13845) );
  AND2_X1 U8839 ( .A1(n11522), .A2(n11521), .ZN(n14265) );
  OAI21_X1 U8840 ( .B1(n11175), .B2(n6979), .A(n6976), .ZN(n13656) );
  NAND2_X1 U8841 ( .A1(n6955), .A2(n6958), .ZN(n14115) );
  NAND2_X1 U8842 ( .A1(n10994), .A2(n10993), .ZN(n11037) );
  NAND2_X1 U8843 ( .A1(n7187), .A2(n11000), .ZN(n11017) );
  NAND2_X1 U8844 ( .A1(n10999), .A2(n11768), .ZN(n7187) );
  NAND2_X1 U8845 ( .A1(n7194), .A2(n10410), .ZN(n10576) );
  NAND2_X1 U8846 ( .A1(n10409), .A2(n10408), .ZN(n7194) );
  OR2_X1 U8847 ( .A1(n13679), .A2(n14414), .ZN(n13875) );
  NAND2_X1 U8848 ( .A1(n10252), .A2(n10251), .ZN(n10336) );
  NAND2_X1 U8849 ( .A1(n14420), .A2(n9617), .ZN(n13876) );
  INV_X1 U8850 ( .A(n13876), .ZN(n14430) );
  NAND2_X1 U8851 ( .A1(n13886), .A2(n6924), .ZN(n13961) );
  INV_X1 U8852 ( .A(n6925), .ZN(n6924) );
  OAI21_X1 U8853 ( .B1(n13887), .B2(n14528), .A(n13885), .ZN(n6925) );
  AND2_X1 U8854 ( .A1(n13902), .A2(n13901), .ZN(n13903) );
  AND2_X1 U8855 ( .A1(n13900), .A2(n13899), .ZN(n13901) );
  AND2_X1 U8856 ( .A1(n6809), .A2(n13907), .ZN(n6745) );
  NAND2_X1 U8857 ( .A1(n7573), .A2(n9415), .ZN(n9416) );
  AOI21_X1 U8858 ( .B1(n6628), .B2(n9411), .A(n13973), .ZN(n6627) );
  INV_X1 U8859 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11007) );
  INV_X1 U8860 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10582) );
  OR2_X1 U8861 ( .A1(n9574), .A2(n9573), .ZN(n7296) );
  INV_X1 U8862 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10076) );
  INV_X1 U8863 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10176) );
  INV_X1 U8864 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10079) );
  INV_X1 U8865 ( .A(n11177), .ZN(n11137) );
  INV_X1 U8866 ( .A(n11025), .ZN(n10186) );
  INV_X1 U8867 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9819) );
  INV_X1 U8868 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9755) );
  NAND2_X1 U8869 ( .A1(n7898), .A2(n7897), .ZN(n7900) );
  INV_X1 U8870 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9748) );
  INV_X1 U8871 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9704) );
  OAI21_X1 U8872 ( .B1(n7845), .B2(n6997), .A(n6995), .ZN(n7863) );
  NAND2_X1 U8873 ( .A1(n7846), .A2(n6817), .ZN(n7862) );
  NOR2_X1 U8874 ( .A1(n7861), .A2(n6997), .ZN(n6817) );
  OAI21_X1 U8875 ( .B1(n7844), .B2(n7845), .A(n7846), .ZN(n10269) );
  INV_X1 U8876 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9698) );
  INV_X1 U8877 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9671) );
  OR2_X1 U8878 ( .A1(n7828), .A2(n7827), .ZN(n7829) );
  INV_X1 U8879 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9667) );
  INV_X1 U8880 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9692) );
  INV_X1 U8881 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9687) );
  INV_X1 U8882 ( .A(n7773), .ZN(n7775) );
  NAND2_X1 U8883 ( .A1(n6915), .A2(n7587), .ZN(n7755) );
  INV_X1 U8884 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7021) );
  XNOR2_X1 U8885 ( .A(n14060), .B(n7074), .ZN(n14106) );
  INV_X1 U8886 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7074) );
  INV_X1 U8887 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6818) );
  NAND2_X1 U8888 ( .A1(n7075), .A2(n14076), .ZN(n14111) );
  NAND2_X1 U8889 ( .A1(n14108), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7075) );
  NAND2_X1 U8890 ( .A1(n6764), .A2(n14109), .ZN(n14320) );
  OAI21_X1 U8891 ( .B1(n14111), .B2(n14110), .A(P2_ADDR_REG_10__SCAN_IN), .ZN(
        n6764) );
  INV_X1 U8892 ( .A(n14331), .ZN(n6768) );
  INV_X1 U8893 ( .A(n7069), .ZN(n6767) );
  NAND2_X1 U8894 ( .A1(n14135), .A2(n14136), .ZN(n14134) );
  OAI21_X1 U8895 ( .B1(n12475), .B2(n11968), .A(n9169), .ZN(n9170) );
  INV_X1 U8896 ( .A(n6826), .ZN(n6825) );
  OAI21_X1 U8897 ( .B1(n12479), .B2(n11968), .A(n11967), .ZN(n6826) );
  OAI21_X1 U8898 ( .B1(n8951), .B2(n6599), .A(n8970), .ZN(n6606) );
  XNOR2_X1 U8899 ( .A(n12173), .B(n12174), .ZN(n6862) );
  MUX2_X1 U8900 ( .A(n12406), .B(n12472), .S(n14990), .Z(n12407) );
  OAI21_X1 U8901 ( .B1(n9183), .B2(n14973), .A(n6570), .ZN(P3_U3456) );
  NAND2_X1 U8902 ( .A1(n14973), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n6820) );
  MUX2_X1 U8903 ( .A(n12473), .B(n12472), .S(n14974), .Z(n12474) );
  NAND2_X1 U8904 ( .A1(n7338), .A2(n12689), .ZN(n7337) );
  AND2_X1 U8905 ( .A1(n9397), .A2(n9396), .ZN(n9398) );
  OAI211_X1 U8906 ( .C1(n12865), .C2(n13078), .A(n7551), .B(n7549), .ZN(
        P2_U3236) );
  AOI21_X1 U8907 ( .B1(n12864), .B2(n13085), .A(n12863), .ZN(n7551) );
  AND2_X1 U8908 ( .A1(n7120), .A2(n7122), .ZN(n12865) );
  NAND2_X1 U8909 ( .A1(n7550), .A2(n12988), .ZN(n7549) );
  INV_X1 U8910 ( .A(n13342), .ZN(n6790) );
  NAND2_X1 U8911 ( .A1(n14230), .A2(n13250), .ZN(n14206) );
  INV_X1 U8912 ( .A(n6782), .ZN(n6781) );
  OAI21_X1 U8913 ( .B1(n13895), .B2(n14489), .A(n7236), .ZN(n6782) );
  AND2_X1 U8914 ( .A1(n7227), .A2(n7235), .ZN(n7226) );
  AND2_X1 U8915 ( .A1(n7233), .A2(n7229), .ZN(n7224) );
  NAND2_X1 U8916 ( .A1(n6753), .A2(n6752), .ZN(P1_U3522) );
  NAND2_X1 U8917 ( .A1(n7230), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6752) );
  NAND2_X1 U8918 ( .A1(n6757), .A2(n6756), .ZN(P1_U3520) );
  NAND2_X1 U8919 ( .A1(n7230), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6756) );
  INV_X1 U8920 ( .A(n7057), .ZN(n14338) );
  XNOR2_X1 U8921 ( .A(n14146), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n7080) );
  AOI21_X1 U8922 ( .B1(n7533), .B2(n8188), .A(n6462), .ZN(n7531) );
  CLKBUF_X3 U8923 ( .A(n11449), .Z(n11719) );
  NOR2_X1 U8924 ( .A1(n12986), .A2(n7534), .ZN(n7533) );
  OR2_X1 U8925 ( .A1(n8993), .A2(n8992), .ZN(n6453) );
  INV_X1 U8926 ( .A(n14114), .ZN(n6957) );
  NAND2_X2 U8927 ( .A1(n11010), .A2(n8195), .ZN(n10022) );
  AND2_X1 U8928 ( .A1(n13282), .A2(n7476), .ZN(n6454) );
  AND2_X1 U8929 ( .A1(n6761), .A2(n6760), .ZN(n6455) );
  NAND3_X1 U8930 ( .A1(n6966), .A2(n9562), .A3(n9563), .ZN(n13486) );
  INV_X1 U8931 ( .A(n13486), .ZN(n9861) );
  OAI22_X1 U8932 ( .A1(n14676), .A2(n9342), .B1(n10453), .B2(n6445), .ZN(n9217) );
  AND2_X1 U8933 ( .A1(n13931), .A2(n6946), .ZN(n6456) );
  NAND2_X1 U8934 ( .A1(n11558), .A2(n11557), .ZN(n13860) );
  INV_X1 U8935 ( .A(n13648), .ZN(n13911) );
  AND2_X1 U8936 ( .A1(n11312), .A2(n11282), .ZN(n6457) );
  AND2_X1 U8937 ( .A1(n7126), .A2(n13065), .ZN(n6458) );
  AND2_X1 U8938 ( .A1(n7612), .A2(n7250), .ZN(n6459) );
  AND3_X1 U8939 ( .A1(n7730), .A2(n7653), .A3(n6551), .ZN(n6460) );
  INV_X1 U8940 ( .A(n14803), .ZN(n7154) );
  XNOR2_X1 U8941 ( .A(n10090), .B(n14659), .ZN(n10422) );
  AND2_X1 U8942 ( .A1(n8835), .A2(n8837), .ZN(n6461) );
  AND2_X1 U8943 ( .A1(n13134), .A2(n13005), .ZN(n6462) );
  NAND2_X1 U8944 ( .A1(n6623), .A2(n6501), .ZN(n6463) );
  AND2_X1 U8945 ( .A1(n8872), .A2(n8876), .ZN(n12334) );
  AND2_X1 U8946 ( .A1(n9014), .A2(n8888), .ZN(n6464) );
  AND2_X1 U8947 ( .A1(n14887), .A2(n11276), .ZN(n6465) );
  OR2_X1 U8948 ( .A1(n11503), .A2(n11738), .ZN(n6466) );
  NOR2_X1 U8949 ( .A1(n7061), .A2(n7060), .ZN(n6467) );
  NOR2_X1 U8950 ( .A1(n7527), .A2(n9240), .ZN(n7523) );
  NAND2_X1 U8951 ( .A1(n6548), .A2(n13655), .ZN(n6468) );
  AND2_X1 U8952 ( .A1(n7339), .A2(n6530), .ZN(n6469) );
  AND2_X1 U8953 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n6470) );
  NAND2_X1 U8954 ( .A1(n8717), .A2(n8716), .ZN(n9132) );
  INV_X1 U8955 ( .A(n8246), .ZN(n7092) );
  INV_X1 U8956 ( .A(n13036), .ZN(n13153) );
  AND2_X1 U8957 ( .A1(n7689), .A2(n7688), .ZN(n13036) );
  NOR2_X1 U8958 ( .A1(n9253), .A2(n9252), .ZN(n6471) );
  OR2_X1 U8959 ( .A1(n6466), .A2(n6974), .ZN(n6472) );
  AND2_X1 U8960 ( .A1(n6551), .A2(n7674), .ZN(n6473) );
  AND3_X1 U8961 ( .A1(n6681), .A2(n6680), .A3(n6677), .ZN(n6474) );
  OR2_X1 U8962 ( .A1(n7181), .A2(n6962), .ZN(n6475) );
  AND2_X1 U8963 ( .A1(n11710), .A2(n11709), .ZN(n6476) );
  INV_X1 U8964 ( .A(n8188), .ZN(n7538) );
  INV_X1 U8965 ( .A(n13344), .ZN(n6632) );
  OR2_X1 U8966 ( .A1(n7995), .A2(SI_21_), .ZN(n6477) );
  INV_X1 U8967 ( .A(n12724), .ZN(n12689) );
  NAND2_X1 U8968 ( .A1(n11021), .A2(n11020), .ZN(n14120) );
  INV_X1 U8969 ( .A(n14120), .ZN(n6936) );
  INV_X1 U8970 ( .A(n11766), .ZN(n6965) );
  INV_X2 U8971 ( .A(n14973), .ZN(n14974) );
  OAI21_X1 U8972 ( .B1(n6783), .B2(n7860), .A(n7859), .ZN(n10717) );
  AND3_X1 U8973 ( .A1(n10117), .A2(n7458), .A3(n10118), .ZN(n6478) );
  AND2_X1 U8974 ( .A1(n8289), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6479) );
  INV_X1 U8975 ( .A(n6435), .ZN(n10347) );
  INV_X2 U8976 ( .A(n8056), .ZN(n7786) );
  NAND2_X1 U8977 ( .A1(n10483), .A2(n10482), .ZN(n6480) );
  XOR2_X2 U8978 ( .A(n13648), .B(n13671), .Z(n6481) );
  NAND2_X2 U8979 ( .A1(n9538), .A2(n9554), .ZN(n13984) );
  INV_X1 U8980 ( .A(n11769), .ZN(n6982) );
  AND2_X1 U8981 ( .A1(n6768), .A2(n6767), .ZN(n6482) );
  NAND2_X1 U8982 ( .A1(n13129), .A2(n12975), .ZN(n6483) );
  OR2_X1 U8983 ( .A1(n8952), .A2(P3_IR_REG_22__SCAN_IN), .ZN(n6484) );
  INV_X1 U8984 ( .A(n6852), .ZN(n10142) );
  NAND2_X1 U8985 ( .A1(n8397), .A2(n6853), .ZN(n6852) );
  AND2_X1 U8986 ( .A1(n13655), .A2(n11510), .ZN(n6485) );
  AND2_X1 U8987 ( .A1(n13787), .A2(n6943), .ZN(n6486) );
  AND2_X1 U8988 ( .A1(n6629), .A2(n13345), .ZN(n6487) );
  NAND2_X1 U8989 ( .A1(n7649), .A2(n7634), .ZN(n7781) );
  AND2_X1 U8990 ( .A1(n7470), .A2(n7468), .ZN(n6488) );
  AND2_X1 U8991 ( .A1(n7787), .A2(n7790), .ZN(n6489) );
  AND2_X1 U8992 ( .A1(n10892), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n6490) );
  INV_X1 U8993 ( .A(n7498), .ZN(n7497) );
  NOR2_X1 U8994 ( .A1(n8191), .A2(n7506), .ZN(n7498) );
  NOR2_X1 U8995 ( .A1(n11679), .A2(n11677), .ZN(n6491) );
  AND2_X1 U8996 ( .A1(n13226), .A2(n13221), .ZN(n6492) );
  INV_X1 U8997 ( .A(n11741), .ZN(n7273) );
  OR3_X1 U8998 ( .A1(n8647), .A2(n7025), .A3(P3_IR_REG_18__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U8999 ( .A1(n7676), .A2(n11429), .ZN(n7762) );
  INV_X1 U9000 ( .A(n10329), .ZN(n6972) );
  OR2_X1 U9001 ( .A1(n13433), .A2(n14194), .ZN(n6494) );
  INV_X1 U9002 ( .A(n11433), .ZN(n9610) );
  INV_X1 U9003 ( .A(n7454), .ZN(n7453) );
  NAND2_X1 U9004 ( .A1(n13664), .A2(n13836), .ZN(n6495) );
  INV_X1 U9005 ( .A(n10243), .ZN(n14480) );
  NAND2_X1 U9006 ( .A1(n10110), .A2(n10109), .ZN(n10243) );
  INV_X1 U9007 ( .A(n11768), .ZN(n7184) );
  INV_X1 U9008 ( .A(n13167), .ZN(n7014) );
  NOR4_X1 U9009 ( .A1(n12991), .A2(n13026), .A3(n13011), .A4(n9373), .ZN(n6496) );
  NAND2_X1 U9010 ( .A1(n7887), .A2(n7886), .ZN(n10793) );
  INV_X1 U9011 ( .A(n10793), .ZN(n6802) );
  INV_X1 U9012 ( .A(n12848), .ZN(n6837) );
  INV_X1 U9013 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9555) );
  AND2_X1 U9014 ( .A1(n11341), .A2(n11340), .ZN(n6497) );
  AND2_X1 U9015 ( .A1(n10471), .A2(n10438), .ZN(n6498) );
  XNOR2_X1 U9016 ( .A(n13118), .B(n12631), .ZN(n12929) );
  INV_X1 U9017 ( .A(n11786), .ZN(n7278) );
  AND2_X1 U9018 ( .A1(n6457), .A2(n11412), .ZN(n6499) );
  INV_X1 U9019 ( .A(n7603), .ZN(n6997) );
  NAND2_X1 U9020 ( .A1(n12546), .A2(n12545), .ZN(n6500) );
  AND2_X1 U9021 ( .A1(n8036), .A2(n8035), .ZN(n12939) );
  INV_X1 U9022 ( .A(n11493), .ZN(n6898) );
  OR2_X1 U9023 ( .A1(n11899), .A2(n9136), .ZN(n6501) );
  AND2_X1 U9024 ( .A1(n8923), .A2(n9044), .ZN(n6502) );
  AND3_X1 U9025 ( .A1(n9997), .A2(n9996), .A3(n9995), .ZN(n11450) );
  INV_X1 U9026 ( .A(n11450), .ZN(n6748) );
  INV_X1 U9027 ( .A(n9290), .ZN(n7481) );
  INV_X1 U9028 ( .A(n12199), .ZN(n7384) );
  OAI22_X1 U9029 ( .A1(n14716), .A2(n9213), .B1(n11288), .B2(n9342), .ZN(n9238) );
  AND2_X1 U9030 ( .A1(n7177), .A2(n14384), .ZN(n6503) );
  OR3_X1 U9031 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6504) );
  INV_X1 U9032 ( .A(n7007), .ZN(n12952) );
  NOR2_X1 U9033 ( .A1(n7526), .A2(n9241), .ZN(n7525) );
  AND2_X1 U9034 ( .A1(n6920), .A2(n13642), .ZN(n6505) );
  OR2_X1 U9035 ( .A1(n13036), .A2(n12728), .ZN(n6506) );
  AND2_X1 U9036 ( .A1(n13725), .A2(n7175), .ZN(n6507) );
  INV_X1 U9037 ( .A(n9374), .ZN(n12963) );
  AND2_X1 U9038 ( .A1(n12867), .A2(n12868), .ZN(n6508) );
  AND2_X1 U9039 ( .A1(n9127), .A2(n9124), .ZN(n6509) );
  AND2_X1 U9040 ( .A1(n9086), .A2(n9085), .ZN(n6510) );
  INV_X1 U9041 ( .A(n7394), .ZN(n7390) );
  AND2_X1 U9042 ( .A1(n9225), .A2(n9223), .ZN(n6511) );
  AND2_X1 U9043 ( .A1(n9225), .A2(n9221), .ZN(n6512) );
  AND2_X1 U9044 ( .A1(n9548), .A2(n9549), .ZN(n6513) );
  INV_X1 U9045 ( .A(n7408), .ZN(n7407) );
  NAND2_X1 U9046 ( .A1(n6453), .A2(n8990), .ZN(n7408) );
  INV_X1 U9047 ( .A(n7424), .ZN(n7423) );
  OAI22_X1 U9048 ( .A1(n9014), .A2(n7428), .B1(n12282), .B2(n12420), .ZN(n7424) );
  NAND2_X1 U9049 ( .A1(n13898), .A2(n13675), .ZN(n6514) );
  AND2_X1 U9050 ( .A1(n13812), .A2(n7210), .ZN(n6515) );
  AND2_X1 U9051 ( .A1(n8683), .A2(n8929), .ZN(n6516) );
  AND2_X1 U9052 ( .A1(n7422), .A2(n7421), .ZN(n6517) );
  OR2_X1 U9053 ( .A1(n7763), .A2(n12747), .ZN(n6518) );
  AND2_X1 U9054 ( .A1(n7324), .A2(n7322), .ZN(n6519) );
  INV_X1 U9055 ( .A(n7533), .ZN(n7532) );
  AND2_X1 U9056 ( .A1(n12129), .A2(n14157), .ZN(n6520) );
  OR2_X1 U9057 ( .A1(n7481), .A2(n7480), .ZN(n6521) );
  NOR2_X1 U9058 ( .A1(n14515), .A2(n13479), .ZN(n6522) );
  NOR2_X1 U9059 ( .A1(n14226), .A2(n13476), .ZN(n6523) );
  NOR2_X1 U9060 ( .A1(n11464), .A2(n13482), .ZN(n6524) );
  NOR2_X1 U9061 ( .A1(n14226), .A2(n11344), .ZN(n6525) );
  NOR2_X1 U9062 ( .A1(n13945), .A2(n13641), .ZN(n6526) );
  NOR2_X1 U9063 ( .A1(n12496), .A2(n12332), .ZN(n6527) );
  NOR2_X1 U9064 ( .A1(n13274), .A2(n13273), .ZN(n6528) );
  NAND2_X1 U9065 ( .A1(n11509), .A2(n11738), .ZN(n6529) );
  INV_X1 U9066 ( .A(n7503), .ZN(n7502) );
  NAND2_X1 U9067 ( .A1(n12909), .A2(n12629), .ZN(n7503) );
  INV_X1 U9068 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13189) );
  INV_X1 U9069 ( .A(n6944), .ZN(n6943) );
  NAND2_X1 U9070 ( .A1(n6456), .A2(n6945), .ZN(n6944) );
  AND2_X1 U9071 ( .A1(n7646), .A2(n6474), .ZN(n7671) );
  NAND2_X1 U9072 ( .A1(n7344), .A2(n7346), .ZN(n6530) );
  INV_X1 U9073 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8137) );
  INV_X1 U9074 ( .A(n7506), .ZN(n7505) );
  NOR2_X1 U9075 ( .A1(n12939), .A2(n12631), .ZN(n7506) );
  INV_X1 U9076 ( .A(n7565), .ZN(n7428) );
  INV_X1 U9077 ( .A(n7433), .ZN(n7432) );
  NAND2_X1 U9078 ( .A1(n8303), .A2(n7434), .ZN(n7433) );
  INV_X1 U9079 ( .A(n7267), .ZN(n7266) );
  NOR2_X1 U9080 ( .A1(n6481), .A2(n13738), .ZN(n7267) );
  INV_X1 U9081 ( .A(n6990), .ZN(n7239) );
  NAND2_X1 U9082 ( .A1(n7240), .A2(n7245), .ZN(n6990) );
  INV_X1 U9083 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8314) );
  INV_X1 U9084 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9658) );
  AND2_X1 U9085 ( .A1(n13113), .A2(n12657), .ZN(n6531) );
  INV_X1 U9086 ( .A(n7465), .ZN(n7464) );
  NAND2_X1 U9087 ( .A1(n13272), .A2(n7466), .ZN(n7465) );
  OR2_X1 U9088 ( .A1(n7441), .A2(n9416), .ZN(n6532) );
  INV_X1 U9089 ( .A(n11477), .ZN(n7285) );
  NAND2_X1 U9090 ( .A1(n11410), .A2(n11411), .ZN(n6533) );
  NAND2_X1 U9091 ( .A1(n13634), .A2(n13864), .ZN(n6534) );
  NAND2_X1 U9092 ( .A1(n9663), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8248) );
  XNOR2_X1 U9093 ( .A(n14692), .B(n6816), .ZN(n10788) );
  INV_X1 U9094 ( .A(n9014), .ZN(n12263) );
  AND2_X1 U9095 ( .A1(n8899), .A2(n8714), .ZN(n9014) );
  AND2_X1 U9096 ( .A1(n13108), .A2(n12918), .ZN(n6535) );
  NOR2_X1 U9097 ( .A1(n9255), .A2(n9257), .ZN(n6536) );
  NAND2_X1 U9098 ( .A1(n14881), .A2(n8991), .ZN(n6537) );
  INV_X1 U9099 ( .A(n11630), .ZN(n7286) );
  NOR2_X1 U9100 ( .A1(n12939), .A2(n12917), .ZN(n6538) );
  OAI21_X1 U9101 ( .B1(n7391), .B2(n7390), .A(n9016), .ZN(n7389) );
  NAND2_X1 U9102 ( .A1(n11508), .A2(n6494), .ZN(n6539) );
  OR2_X1 U9103 ( .A1(n11069), .A2(n11068), .ZN(n6761) );
  INV_X1 U9104 ( .A(n6875), .ZN(n6874) );
  INV_X1 U9105 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7553) );
  INV_X1 U9106 ( .A(n11601), .ZN(n6887) );
  NAND2_X1 U9107 ( .A1(n9292), .A2(n7479), .ZN(n6540) );
  OR2_X1 U9108 ( .A1(n11720), .A2(n6476), .ZN(n6541) );
  NAND2_X1 U9109 ( .A1(n8023), .A2(n6483), .ZN(n6542) );
  OR2_X1 U9110 ( .A1(n9218), .A2(n9216), .ZN(n6543) );
  AND2_X1 U9111 ( .A1(n7251), .A2(n7250), .ZN(n6544) );
  INV_X1 U9112 ( .A(n13655), .ZN(n6974) );
  INV_X1 U9113 ( .A(n9371), .ZN(n13059) );
  OR2_X1 U9114 ( .A1(n14144), .A2(n14143), .ZN(n6545) );
  AND3_X1 U9115 ( .A1(n8945), .A2(n8921), .A3(n8923), .ZN(n6546) );
  AND2_X1 U9116 ( .A1(n7044), .A2(n7042), .ZN(n6547) );
  NAND2_X1 U9117 ( .A1(n9125), .A2(n9126), .ZN(n7063) );
  NOR2_X1 U9118 ( .A1(n11771), .A2(n11504), .ZN(n6548) );
  AND2_X1 U9119 ( .A1(n8196), .A2(n7122), .ZN(n6549) );
  NOR2_X1 U9120 ( .A1(n10471), .A2(n12741), .ZN(n6550) );
  AND2_X1 U9121 ( .A1(n7670), .A2(n7553), .ZN(n6551) );
  AND2_X1 U9122 ( .A1(n7319), .A2(n12638), .ZN(n6552) );
  AND2_X1 U9123 ( .A1(n6540), .A2(n9323), .ZN(n6553) );
  AND2_X1 U9124 ( .A1(n8798), .A2(n8822), .ZN(n10616) );
  INV_X1 U9125 ( .A(n10616), .ZN(n8988) );
  AND2_X1 U9126 ( .A1(n13148), .A2(n12697), .ZN(n6554) );
  AND2_X1 U9127 ( .A1(n12190), .A2(n11983), .ZN(n8924) );
  AND2_X1 U9128 ( .A1(n9535), .A2(n7478), .ZN(n6555) );
  AND2_X1 U9129 ( .A1(n8924), .A2(n12181), .ZN(n6556) );
  NOR2_X1 U9130 ( .A1(n8205), .A2(n7645), .ZN(n7646) );
  OR2_X1 U9131 ( .A1(n11742), .A2(n7273), .ZN(n6557) );
  OR2_X1 U9132 ( .A1(n11709), .A2(n11710), .ZN(n6558) );
  AND2_X1 U9133 ( .A1(n7278), .A2(n11753), .ZN(n6559) );
  AND2_X1 U9134 ( .A1(n6555), .A2(n9537), .ZN(n6560) );
  NOR2_X1 U9135 ( .A1(n9211), .A2(n9212), .ZN(n7489) );
  INV_X1 U9136 ( .A(n14405), .ZN(n6953) );
  INV_X1 U9137 ( .A(n13672), .ZN(n13653) );
  XNOR2_X1 U9138 ( .A(n13890), .B(n13693), .ZN(n13672) );
  NAND2_X1 U9139 ( .A1(n14809), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U9140 ( .A1(n13022), .A2(n13003), .ZN(n6562) );
  INV_X1 U9141 ( .A(n7037), .ZN(n7036) );
  NAND2_X1 U9142 ( .A1(n9076), .A2(n11995), .ZN(n7037) );
  AND2_X1 U9143 ( .A1(n12535), .A2(n12714), .ZN(n7321) );
  INV_X1 U9144 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7352) );
  AND2_X1 U9145 ( .A1(n9292), .A2(n6521), .ZN(n6563) );
  INV_X1 U9146 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7478) );
  NAND2_X1 U9147 ( .A1(n11535), .A2(n11534), .ZN(n11568) );
  INV_X1 U9148 ( .A(n11568), .ZN(n6940) );
  AOI21_X1 U9149 ( .B1(n12255), .B2(n8756), .A(n8722), .ZN(n12266) );
  INV_X1 U9150 ( .A(n12266), .ZN(n6590) );
  INV_X1 U9151 ( .A(n11153), .ZN(n7404) );
  XNOR2_X1 U9152 ( .A(n13780), .B(n13667), .ZN(n13772) );
  INV_X1 U9153 ( .A(n13772), .ZN(n7241) );
  INV_X1 U9154 ( .A(n13919), .ZN(n6945) );
  INV_X1 U9155 ( .A(n14237), .ZN(n6931) );
  NAND2_X1 U9156 ( .A1(n11642), .A2(n11641), .ZN(n13926) );
  INV_X1 U9157 ( .A(n13926), .ZN(n6946) );
  NAND2_X1 U9158 ( .A1(n8564), .A2(n8303), .ZN(n8566) );
  OAI211_X1 U9159 ( .C1(n8772), .C2(n15025), .A(n8700), .B(n8699), .ZN(n11987)
         );
  INV_X1 U9160 ( .A(n11987), .ZN(n12294) );
  INV_X1 U9161 ( .A(n9264), .ZN(n6772) );
  INV_X1 U9162 ( .A(n12657), .ZN(n12932) );
  AND2_X1 U9163 ( .A1(n8061), .A2(n8060), .ZN(n12657) );
  INV_X1 U9164 ( .A(SI_1_), .ZN(n6916) );
  NAND2_X1 U9165 ( .A1(n7366), .A2(n7365), .ZN(n12381) );
  INV_X1 U9166 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7351) );
  INV_X1 U9167 ( .A(n13945), .ZN(n6938) );
  AND2_X1 U9168 ( .A1(n11565), .A2(n11564), .ZN(n13864) );
  INV_X1 U9169 ( .A(n13416), .ZN(n6631) );
  INV_X1 U9170 ( .A(n13441), .ZN(n7475) );
  INV_X1 U9171 ( .A(n7731), .ZN(n6681) );
  INV_X1 U9172 ( .A(n11498), .ZN(n6894) );
  AND2_X1 U9173 ( .A1(n7696), .A2(n7695), .ZN(n13014) );
  AND4_X1 U9174 ( .A1(n7725), .A2(n7724), .A3(n7723), .A4(n7722), .ZN(n12648)
         );
  INV_X1 U9175 ( .A(n12648), .ZN(n7136) );
  AOI22_X1 U9176 ( .A1(n11464), .A2(n6443), .B1(n13331), .B2(n13482), .ZN(
        n10758) );
  INV_X1 U9177 ( .A(n10758), .ZN(n6654) );
  INV_X1 U9178 ( .A(n7468), .ZN(n7467) );
  NOR2_X1 U9179 ( .A1(n13452), .A2(n7469), .ZN(n7468) );
  INV_X1 U9180 ( .A(n13263), .ZN(n7471) );
  AND2_X1 U9181 ( .A1(n7964), .A2(n10167), .ZN(n6564) );
  INV_X1 U9182 ( .A(n11232), .ZN(n7207) );
  OR2_X1 U9183 ( .A1(n8647), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6565) );
  AND2_X1 U9184 ( .A1(n6975), .A2(n6980), .ZN(n6566) );
  AND2_X1 U9185 ( .A1(n14162), .A2(n11920), .ZN(n6567) );
  AND2_X1 U9186 ( .A1(n13045), .A2(n12729), .ZN(n6568) );
  AND2_X1 U9187 ( .A1(n12444), .A2(n11952), .ZN(n6569) );
  INV_X1 U9188 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10012) );
  INV_X1 U9189 ( .A(n13074), .ZN(n13162) );
  AND2_X1 U9190 ( .A1(n7717), .A2(n7716), .ZN(n13074) );
  AND2_X1 U9191 ( .A1(n9185), .A2(n6820), .ZN(n6570) );
  AND2_X1 U9192 ( .A1(n7615), .A2(n9660), .ZN(n6571) );
  NOR2_X1 U9193 ( .A1(n7552), .A2(n9256), .ZN(n6572) );
  INV_X1 U9194 ( .A(n9285), .ZN(n7548) );
  OR2_X1 U9195 ( .A1(n7992), .A2(SI_20_), .ZN(n6573) );
  AND2_X1 U9196 ( .A1(n6984), .A2(n6494), .ZN(n6574) );
  INV_X1 U9197 ( .A(n7745), .ZN(n7727) );
  AND2_X1 U9198 ( .A1(n12328), .A2(n9008), .ZN(n6575) );
  AND2_X1 U9199 ( .A1(n6842), .A2(n6841), .ZN(n6576) );
  OR2_X1 U9200 ( .A1(n7548), .A2(n7547), .ZN(n6577) );
  INV_X1 U9201 ( .A(n7134), .ZN(n7133) );
  NOR2_X1 U9202 ( .A1(n13074), .A2(n7136), .ZN(n7134) );
  INV_X1 U9203 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9991) );
  INV_X1 U9204 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7028) );
  INV_X1 U9205 ( .A(n10132), .ZN(n9044) );
  NAND2_X1 U9206 ( .A1(n11027), .A2(n11026), .ZN(n13433) );
  INV_X1 U9207 ( .A(n13433), .ZN(n6934) );
  OAI22_X1 U9208 ( .A1(n10818), .A2(n10817), .B1(n10815), .B2(n10816), .ZN(
        n11062) );
  AOI21_X1 U9209 ( .B1(n11339), .B2(n6635), .A(n6497), .ZN(n13212) );
  AND2_X1 U9210 ( .A1(n6695), .A2(n10529), .ZN(n10534) );
  OAI21_X1 U9211 ( .B1(n10424), .B2(n6676), .A(n6674), .ZN(n10436) );
  INV_X1 U9212 ( .A(n14285), .ZN(n6932) );
  AND2_X1 U9213 ( .A1(n12029), .A2(n12061), .ZN(n6578) );
  INV_X1 U9214 ( .A(n14122), .ZN(n6937) );
  NAND2_X1 U9215 ( .A1(n7397), .A2(n8987), .ZN(n10615) );
  AND2_X1 U9216 ( .A1(n10540), .A2(n10539), .ZN(n6579) );
  NOR2_X1 U9217 ( .A1(n14857), .A2(n10906), .ZN(n6580) );
  NAND3_X1 U9218 ( .A1(n9408), .A2(n9407), .A3(n7293), .ZN(n7295) );
  OR2_X1 U9219 ( .A1(n6628), .A2(n13973), .ZN(n6581) );
  AND2_X1 U9220 ( .A1(n7452), .A2(n7454), .ZN(n6582) );
  INV_X1 U9221 ( .A(n14546), .ZN(n7230) );
  INV_X1 U9222 ( .A(n12165), .ZN(n6811) );
  NOR2_X1 U9223 ( .A1(n12177), .A2(n9150), .ZN(n6583) );
  AND2_X1 U9224 ( .A1(n10198), .A2(n10628), .ZN(n10132) );
  AND2_X1 U9225 ( .A1(n12612), .A2(n12613), .ZN(n12611) );
  NAND2_X1 U9226 ( .A1(n9365), .A2(n6686), .ZN(n10375) );
  INV_X1 U9227 ( .A(n14468), .ZN(n14412) );
  INV_X1 U9228 ( .A(n13065), .ZN(n13029) );
  AND2_X1 U9229 ( .A1(n8762), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6584) );
  AND2_X1 U9230 ( .A1(n8286), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6585) );
  INV_X1 U9231 ( .A(n14911), .ZN(n7109) );
  AND2_X1 U9232 ( .A1(n12087), .A2(n12084), .ZN(n6586) );
  NOR2_X1 U9233 ( .A1(n8296), .A2(n7114), .ZN(n7113) );
  AND2_X1 U9234 ( .A1(n7156), .A2(n7155), .ZN(n6587) );
  INV_X1 U9235 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n7077) );
  INV_X1 U9236 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n7294) );
  NAND3_X1 U9237 ( .A1(n6725), .A2(n6473), .A3(n7646), .ZN(n6724) );
  AND2_X1 U9238 ( .A1(n7146), .A2(n7145), .ZN(n6588) );
  AND2_X1 U9239 ( .A1(n8313), .A2(n7436), .ZN(n8346) );
  AND3_X1 U9240 ( .A1(n9386), .A2(n9390), .A3(n11202), .ZN(n6589) );
  INV_X1 U9241 ( .A(SI_14_), .ZN(n6793) );
  INV_X1 U9242 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7079) );
  INV_X1 U9243 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6839) );
  NAND2_X1 U9244 ( .A1(n6593), .A2(n15122), .ZN(n6592) );
  OAI21_X1 U9245 ( .B1(n8694), .B2(n7098), .A(n7096), .ZN(n6593) );
  NAND2_X1 U9246 ( .A1(n8280), .A2(n8279), .ZN(n6596) );
  NAND2_X1 U9247 ( .A1(n8513), .A2(n8257), .ZN(n8526) );
  NAND2_X1 U9248 ( .A1(n7085), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7084) );
  NAND2_X1 U9249 ( .A1(n6598), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U9250 ( .A1(n11609), .A2(n6598), .ZN(n6848) );
  OAI22_X1 U9251 ( .A1(n6600), .A2(n9019), .B1(n8950), .B2(n8949), .ZN(n6599)
         );
  XNOR2_X1 U9252 ( .A(n8789), .B(n9048), .ZN(n6600) );
  NAND2_X1 U9253 ( .A1(n6603), .A2(n10132), .ZN(n6602) );
  NAND2_X1 U9254 ( .A1(n6605), .A2(n8945), .ZN(n6603) );
  NAND2_X1 U9255 ( .A1(n8922), .A2(n6546), .ZN(n6605) );
  NAND2_X1 U9256 ( .A1(n8242), .A2(n8241), .ZN(n8413) );
  NAND2_X1 U9257 ( .A1(n6606), .A2(n8973), .ZN(P3_U3296) );
  NAND2_X1 U9258 ( .A1(n10197), .A2(n8778), .ZN(n6607) );
  INV_X1 U9259 ( .A(n8398), .ZN(n6610) );
  NAND2_X1 U9260 ( .A1(n6609), .A2(n8239), .ZN(n8374) );
  XNOR2_X1 U9261 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8399) );
  NAND2_X1 U9262 ( .A1(n8511), .A2(n8510), .ZN(n8513) );
  NAND2_X1 U9263 ( .A1(n8685), .A2(n8282), .ZN(n8284) );
  OAI21_X1 U9264 ( .B1(n11886), .B2(n7054), .A(n7051), .ZN(n11950) );
  NAND2_X1 U9265 ( .A1(n6613), .A2(n6611), .ZN(n6614) );
  NAND2_X1 U9266 ( .A1(n11886), .A2(n7051), .ZN(n6613) );
  NAND2_X2 U9267 ( .A1(n11876), .A2(n9142), .ZN(n11961) );
  NAND2_X1 U9268 ( .A1(n11876), .A2(n6615), .ZN(n6619) );
  OAI211_X1 U9269 ( .C1(n6618), .C2(n11821), .A(n11820), .B(n6617), .ZN(
        P3_U3160) );
  NAND2_X1 U9270 ( .A1(n6618), .A2(n6831), .ZN(n6617) );
  AND3_X2 U9271 ( .A1(n6620), .A2(n8375), .A3(n6621), .ZN(n8460) );
  NAND2_X1 U9272 ( .A1(n8376), .A2(n6621), .ZN(n8430) );
  NOR2_X2 U9273 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n6621) );
  OAI21_X1 U9274 ( .B1(n10690), .B2(n6622), .A(n10689), .ZN(n10691) );
  NAND2_X1 U9275 ( .A1(n7030), .A2(n7032), .ZN(n6622) );
  NAND2_X1 U9276 ( .A1(n11833), .A2(n9137), .ZN(n6623) );
  NAND3_X1 U9277 ( .A1(n6623), .A2(n6501), .A3(n11873), .ZN(n9141) );
  NAND2_X1 U9278 ( .A1(n6624), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U9279 ( .A1(n8564), .A2(n7432), .ZN(n6624) );
  NAND2_X2 U9280 ( .A1(n6493), .A2(n6625), .ZN(n12177) );
  AOI22_X1 U9281 ( .A1(n8647), .A2(n7024), .B1(n7022), .B2(n7023), .ZN(n6625)
         );
  NAND3_X1 U9282 ( .A1(n10004), .A2(n6480), .A3(n6626), .ZN(n7459) );
  OAI21_X1 U9283 ( .B1(n10004), .B2(n6626), .A(n10118), .ZN(n10005) );
  NAND2_X1 U9284 ( .A1(n10004), .A2(n6626), .ZN(n10118) );
  XNOR2_X1 U9285 ( .A(n10114), .B(n10113), .ZN(n6626) );
  XNOR2_X1 U9286 ( .A(n6638), .B(n11341), .ZN(n11270) );
  INV_X1 U9287 ( .A(n13250), .ZN(n6642) );
  OAI21_X1 U9288 ( .B1(n13326), .B2(n6649), .A(n6646), .ZN(n6650) );
  NAND2_X1 U9289 ( .A1(n6648), .A2(n13327), .ZN(n6647) );
  INV_X1 U9290 ( .A(n13327), .ZN(n6649) );
  NAND2_X1 U9291 ( .A1(n6650), .A2(n7455), .ZN(n13371) );
  NAND2_X1 U9292 ( .A1(n6655), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9417) );
  NAND4_X1 U9293 ( .A1(n6660), .A2(n6658), .A3(n6657), .A4(n6656), .ZN(n13485)
         );
  NAND2_X1 U9294 ( .A1(n13979), .A2(n9558), .ZN(n10100) );
  OR2_X4 U9295 ( .A1(n13979), .A2(n9558), .ZN(n11634) );
  NAND2_X1 U9298 ( .A1(n6685), .A2(n7133), .ZN(n13047) );
  NAND2_X1 U9299 ( .A1(n7814), .A2(n7597), .ZN(n6663) );
  OAI211_X2 U9300 ( .C1(n7815), .C2(n6665), .A(n7827), .B(n6663), .ZN(n7830)
         );
  NAND2_X1 U9301 ( .A1(n6664), .A2(n7597), .ZN(n7828) );
  NAND2_X1 U9302 ( .A1(n7815), .A2(n7596), .ZN(n6664) );
  INV_X1 U9303 ( .A(n7597), .ZN(n6665) );
  NOR2_X2 U9304 ( .A1(n6666), .A2(n12872), .ZN(n13101) );
  INV_X1 U9305 ( .A(n7158), .ZN(n6670) );
  NOR2_X2 U9306 ( .A1(n7808), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n7730) );
  AOI21_X2 U9307 ( .B1(n11116), .B2(n11115), .A(n7950), .ZN(n7960) );
  NAND2_X1 U9308 ( .A1(n10654), .A2(n10655), .ZN(n6686) );
  XNOR2_X2 U9309 ( .A(n10021), .B(n12745), .ZN(n9886) );
  NAND3_X1 U9310 ( .A1(n7771), .A2(n12684), .A3(n7772), .ZN(n10376) );
  NAND3_X2 U9311 ( .A1(n7783), .A2(n6687), .A3(n7784), .ZN(n12684) );
  AND2_X1 U9312 ( .A1(n7785), .A2(n10376), .ZN(n9365) );
  OR2_X1 U9313 ( .A1(n9337), .A2(n9992), .ZN(n6687) );
  NAND2_X1 U9314 ( .A1(n12686), .A2(n6688), .ZN(n10033) );
  NAND3_X1 U9315 ( .A1(n7318), .A2(n6552), .A3(n6690), .ZN(n12636) );
  NAND2_X1 U9316 ( .A1(n6691), .A2(n7321), .ZN(n6690) );
  INV_X1 U9317 ( .A(n6725), .ZN(n7683) );
  INV_X1 U9318 ( .A(n6695), .ZN(n10530) );
  NOR2_X1 U9319 ( .A1(n10935), .A2(n6696), .ZN(n6697) );
  NAND2_X1 U9320 ( .A1(n10932), .A2(n6697), .ZN(n11080) );
  NAND2_X1 U9321 ( .A1(n6704), .A2(n9196), .ZN(n6736) );
  NAND3_X1 U9322 ( .A1(n7510), .A2(n7509), .A3(n9227), .ZN(n6711) );
  AND2_X1 U9323 ( .A1(n6741), .A2(n6705), .ZN(n9234) );
  NAND3_X1 U9324 ( .A1(n6709), .A2(n9230), .A3(n6706), .ZN(n6705) );
  NAND4_X1 U9325 ( .A1(n7510), .A2(n7509), .A3(n9227), .A4(n6707), .ZN(n6706)
         );
  NAND3_X1 U9326 ( .A1(n7508), .A2(n7507), .A3(n9226), .ZN(n6708) );
  NAND3_X1 U9327 ( .A1(n7508), .A2(n7507), .A3(n6710), .ZN(n6709) );
  NOR2_X1 U9328 ( .A1(n9202), .A2(n6742), .ZN(n6712) );
  INV_X1 U9329 ( .A(n9208), .ZN(n9205) );
  OAI21_X1 U9330 ( .B1(n9289), .B2(n6715), .A(n6713), .ZN(n6719) );
  NAND2_X1 U9331 ( .A1(n9351), .A2(n6718), .ZN(n6717) );
  OAI21_X1 U9332 ( .B1(n9254), .B2(n6722), .A(n6721), .ZN(n9258) );
  INV_X1 U9333 ( .A(n9258), .ZN(n9261) );
  NAND3_X1 U9334 ( .A1(n6778), .A2(n7490), .A3(n6543), .ZN(n6726) );
  NAND2_X1 U9335 ( .A1(n6726), .A2(n6727), .ZN(n9220) );
  OAI22_X1 U9336 ( .A1(n6729), .A2(n6728), .B1(n6731), .B2(n9238), .ZN(n9239)
         );
  AOI22_X1 U9337 ( .A1(n9263), .A2(n9262), .B1(n9261), .B2(n9260), .ZN(n9265)
         );
  OAI21_X1 U9338 ( .B1(n9205), .B2(n9204), .A(n9203), .ZN(n9206) );
  OAI21_X1 U9339 ( .B1(n9272), .B2(n7556), .A(n7554), .ZN(n9275) );
  NAND2_X1 U9340 ( .A1(n7515), .A2(n7516), .ZN(n9246) );
  INV_X1 U9341 ( .A(n9199), .ZN(n6742) );
  OR2_X4 U9342 ( .A1(n11426), .A2(n11429), .ZN(n7763) );
  NAND2_X1 U9343 ( .A1(n7545), .A2(n7546), .ZN(n9289) );
  AOI21_X1 U9344 ( .B1(n9278), .B2(n9277), .A(n9276), .ZN(n9282) );
  AOI22_X1 U9345 ( .A1(n9250), .A2(n9249), .B1(n9248), .B2(n9247), .ZN(n9254)
         );
  INV_X1 U9346 ( .A(n9215), .ZN(n7483) );
  OAI21_X1 U9347 ( .B1(n9282), .B2(n9281), .A(n9280), .ZN(n9284) );
  NOR2_X1 U9348 ( .A1(n7936), .A2(n7150), .ZN(n7149) );
  NAND2_X1 U9349 ( .A1(n10739), .A2(n7896), .ZN(n10670) );
  NAND2_X1 U9350 ( .A1(n7442), .A2(n7443), .ZN(n9926) );
  OAI22_X1 U9351 ( .A1(n12619), .A2(n12618), .B1(n12556), .B2(n12555), .ZN(
        n12557) );
  NAND2_X1 U9352 ( .A1(n7299), .A2(n7298), .ZN(n7301) );
  NAND2_X1 U9353 ( .A1(n10087), .A2(n10088), .ZN(n10205) );
  AOI21_X1 U9354 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n8056), .A(n6737), .ZN(
        n6771) );
  INV_X2 U9355 ( .A(n9337), .ZN(n7682) );
  NAND2_X2 U9356 ( .A1(n9454), .A2(n9657), .ZN(n9337) );
  OAI21_X1 U9357 ( .B1(n9208), .B2(n9207), .A(n9206), .ZN(n9209) );
  INV_X1 U9358 ( .A(n9195), .ZN(n6762) );
  OAI21_X1 U9359 ( .B1(n9234), .B2(n9233), .A(n9232), .ZN(n9236) );
  NAND2_X1 U9360 ( .A1(n7960), .A2(n11406), .ZN(n6738) );
  NAND2_X1 U9361 ( .A1(n7961), .A2(n6738), .ZN(n11387) );
  NAND2_X1 U9362 ( .A1(n7843), .A2(n7842), .ZN(n10452) );
  OAI21_X1 U9363 ( .B1(n11609), .B2(n6839), .A(n6838), .ZN(n7585) );
  NAND2_X1 U9364 ( .A1(n7655), .A2(n7562), .ZN(n8138) );
  NAND2_X1 U9365 ( .A1(n11609), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6838) );
  INV_X1 U9366 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7216) );
  NAND2_X1 U9367 ( .A1(n9657), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6840) );
  NAND2_X1 U9368 ( .A1(n12645), .A2(n12646), .ZN(n12644) );
  XNOR2_X2 U9369 ( .A(n7673), .B(n7672), .ZN(n11426) );
  NAND2_X1 U9370 ( .A1(n10085), .A2(n7302), .ZN(n10087) );
  AOI21_X1 U9371 ( .B1(n9268), .B2(n9267), .A(n9266), .ZN(n9272) );
  OR2_X1 U9372 ( .A1(n9275), .A2(n9274), .ZN(n9278) );
  INV_X1 U9373 ( .A(n7311), .ZN(n7310) );
  NAND2_X1 U9374 ( .A1(n12663), .A2(n12553), .ZN(n12619) );
  NAND2_X1 U9375 ( .A1(n7209), .A2(n7208), .ZN(n13784) );
  OR2_X1 U9376 ( .A1(n13909), .A2(n14489), .ZN(n6809) );
  NAND2_X1 U9377 ( .A1(n7191), .A2(n7192), .ZN(n10600) );
  NAND2_X1 U9378 ( .A1(n7182), .A2(n7185), .ZN(n14113) );
  NAND2_X1 U9379 ( .A1(n9304), .A2(n9303), .ZN(n12848) );
  NAND2_X1 U9380 ( .A1(n11195), .A2(n11771), .ZN(n14284) );
  AND2_X2 U9381 ( .A1(n9408), .A2(n9407), .ZN(n7200) );
  BUF_X1 U9382 ( .A(n11730), .Z(n6743) );
  NAND2_X1 U9383 ( .A1(n11995), .A2(n10636), .ZN(n8812) );
  NAND2_X2 U9384 ( .A1(n7395), .A2(n6464), .ZN(n12262) );
  NAND2_X2 U9385 ( .A1(n8597), .A2(n8857), .ZN(n12373) );
  OAI21_X2 U9386 ( .B1(n11375), .B2(n11377), .A(n8843), .ZN(n11357) );
  AOI21_X2 U9387 ( .B1(n12228), .B2(n8749), .A(n8908), .ZN(n12218) );
  INV_X1 U9388 ( .A(n8313), .ZN(n8960) );
  INV_X1 U9389 ( .A(n7307), .ZN(n7306) );
  AOI21_X2 U9390 ( .B1(n12240), .B2(n8942), .A(n8905), .ZN(n12228) );
  OAI21_X2 U9391 ( .B1(n11152), .B2(n7412), .A(n7409), .ZN(n11375) );
  NAND2_X1 U9392 ( .A1(n6807), .A2(n6806), .ZN(n8901) );
  NAND2_X1 U9393 ( .A1(n7110), .A2(n8979), .ZN(n7108) );
  OAI21_X1 U9394 ( .B1(n8900), .B2(n8899), .A(n8898), .ZN(n6808) );
  NAND2_X1 U9395 ( .A1(n6814), .A2(n6813), .ZN(n7261) );
  NAND2_X1 U9396 ( .A1(n7231), .A2(n6781), .ZN(n13962) );
  AOI21_X1 U9397 ( .B1(n6976), .B2(n6979), .A(n6974), .ZN(n6973) );
  NAND2_X1 U9398 ( .A1(n6821), .A2(n13807), .ZN(n7244) );
  NAND2_X1 U9399 ( .A1(n7321), .A2(n12532), .ZN(n7319) );
  NAND2_X1 U9400 ( .A1(n6747), .A2(n13663), .ZN(n6805) );
  AOI21_X1 U9401 ( .B1(n13847), .B2(n13661), .A(n6746), .ZN(n13831) );
  NAND2_X1 U9402 ( .A1(n7746), .A2(n7745), .ZN(n6794) );
  NOR2_X1 U9403 ( .A1(n13737), .A2(n7266), .ZN(n7264) );
  INV_X1 U9404 ( .A(n13815), .ZN(n6747) );
  NAND2_X1 U9405 ( .A1(n13908), .A2(n6745), .ZN(n13964) );
  NAND2_X1 U9406 ( .A1(n10397), .A2(n10396), .ZN(n10540) );
  NAND4_X2 U9407 ( .A1(n9583), .A2(n9584), .A3(n9582), .A4(n9585), .ZN(n13484)
         );
  NAND2_X1 U9408 ( .A1(n13258), .A2(n13257), .ZN(n13409) );
  OAI21_X2 U9409 ( .B1(n13282), .B2(n7475), .A(n7473), .ZN(n13346) );
  NAND2_X1 U9410 ( .A1(n9931), .A2(n9930), .ZN(n10001) );
  NAND2_X1 U9411 ( .A1(n6978), .A2(n6980), .ZN(n6977) );
  NAND2_X1 U9412 ( .A1(n13965), .A2(n14546), .ZN(n6753) );
  NAND2_X1 U9413 ( .A1(n13915), .A2(n6754), .ZN(n13965) );
  NAND2_X1 U9414 ( .A1(n13967), .A2(n14546), .ZN(n6757) );
  NAND2_X1 U9415 ( .A1(n13927), .A2(n6758), .ZN(n13967) );
  INV_X1 U9416 ( .A(n7451), .ZN(n7450) );
  NOR2_X2 U9417 ( .A1(n12031), .A2(n8579), .ZN(n12049) );
  NOR2_X1 U9418 ( .A1(n12103), .A2(n12104), .ZN(n12106) );
  INV_X1 U9419 ( .A(n6854), .ZN(n6853) );
  NOR2_X1 U9420 ( .A1(n12133), .A2(n12132), .ZN(n12160) );
  AOI21_X2 U9421 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n14847), .A(n14839), .ZN(
        n10904) );
  NAND2_X1 U9422 ( .A1(n15147), .A2(n15148), .ZN(n14066) );
  NAND2_X1 U9423 ( .A1(n12745), .A2(n9213), .ZN(n9194) );
  NAND2_X2 U9424 ( .A1(n6769), .A2(n6775), .ZN(n12745) );
  NAND2_X1 U9425 ( .A1(n7059), .A2(n14602), .ZN(n7058) );
  NAND2_X1 U9426 ( .A1(n6440), .A2(n6586), .ZN(n7140) );
  OAI21_X1 U9427 ( .B1(n14145), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6545), .ZN(
        n7081) );
  INV_X1 U9428 ( .A(n11426), .ZN(n7676) );
  OR2_X1 U9429 ( .A1(n9265), .A2(n6772), .ZN(n9268) );
  NAND2_X1 U9430 ( .A1(n7033), .A2(n7040), .ZN(n7032) );
  NAND2_X1 U9431 ( .A1(n9387), .A2(n6589), .ZN(n9399) );
  INV_X1 U9432 ( .A(n11748), .ZN(n6835) );
  OAI21_X1 U9433 ( .B1(n9209), .B2(n7487), .A(n6779), .ZN(n6778) );
  NAND2_X1 U9434 ( .A1(n7029), .A2(n7038), .ZN(n7031) );
  NAND2_X1 U9435 ( .A1(n7031), .A2(n7037), .ZN(n7030) );
  OAI22_X1 U9436 ( .A1(n11923), .A2(n9101), .B1(n12384), .B2(n9100), .ZN(
        n11827) );
  NAND2_X1 U9437 ( .A1(n6992), .A2(n7249), .ZN(n7924) );
  OAI21_X1 U9438 ( .B1(n6439), .B2(n6988), .A(n6985), .ZN(n13711) );
  INV_X1 U9439 ( .A(n7263), .ZN(n6814) );
  INV_X2 U9440 ( .A(n7841), .ZN(n14676) );
  NAND2_X2 U9441 ( .A1(n8503), .A2(n8502), .ZN(n11152) );
  OR2_X1 U9442 ( .A1(n8781), .A2(n10317), .ZN(n8369) );
  NAND2_X1 U9443 ( .A1(n10702), .A2(n8811), .ZN(n10645) );
  NAND2_X1 U9444 ( .A1(n12347), .A2(n8658), .ZN(n12333) );
  INV_X1 U9445 ( .A(n10757), .ZN(n6810) );
  NAND2_X1 U9446 ( .A1(n13363), .A2(n6785), .ZN(n13343) );
  NAND2_X1 U9447 ( .A1(n12206), .A2(n7384), .ZN(n12205) );
  AOI21_X1 U9448 ( .B1(n7094), .B2(n8288), .A(n6479), .ZN(n7093) );
  OAI21_X1 U9449 ( .B1(n7110), .B2(n7109), .A(n7108), .ZN(n8951) );
  OAI21_X1 U9450 ( .B1(n8918), .B2(n8917), .A(n8974), .ZN(n8922) );
  OR2_X1 U9451 ( .A1(n11209), .A2(n8175), .ZN(n8177) );
  AOI21_X1 U9452 ( .B1(n7542), .B2(n7544), .A(n6550), .ZN(n7540) );
  NAND2_X1 U9453 ( .A1(n8172), .A2(n8171), .ZN(n11114) );
  XNOR2_X1 U9454 ( .A(n8192), .B(n9377), .ZN(n12862) );
  NAND3_X1 U9455 ( .A1(n6795), .A2(n7120), .A3(n6549), .ZN(n8236) );
  NAND2_X1 U9456 ( .A1(n6805), .A2(n6495), .ZN(n6821) );
  XNOR2_X1 U9457 ( .A(n14485), .B(n13483), .ZN(n11757) );
  INV_X1 U9458 ( .A(n8049), .ZN(n7003) );
  NAND2_X1 U9459 ( .A1(n6791), .A2(n6790), .ZN(P1_U3214) );
  NAND2_X1 U9460 ( .A1(n13343), .A2(n14233), .ZN(n6791) );
  NAND2_X1 U9461 ( .A1(n7812), .A2(n7811), .ZN(n10424) );
  INV_X1 U9462 ( .A(n12746), .ZN(n9187) );
  INV_X1 U9463 ( .A(n11429), .ZN(n6815) );
  OAI21_X1 U9464 ( .B1(n9209), .B2(n7489), .A(n7482), .ZN(n7490) );
  AND2_X2 U9465 ( .A1(n10971), .A2(n14186), .ZN(n10970) );
  INV_X1 U9466 ( .A(n6799), .ZN(n12892) );
  NOR2_X2 U9467 ( .A1(n12904), .A2(n13103), .ZN(n6799) );
  NOR2_X4 U9468 ( .A1(n12993), .A2(n13134), .ZN(n12967) );
  NOR2_X2 U9469 ( .A1(n10750), .A2(n10933), .ZN(n10779) );
  AOI21_X1 U9470 ( .B1(n10024), .B2(n10022), .A(n10023), .ZN(n12613) );
  NAND2_X1 U9471 ( .A1(n6976), .A2(n11175), .ZN(n6804) );
  OAI21_X2 U9472 ( .B1(n7588), .B2(SI_2_), .A(n7590), .ZN(n7774) );
  INV_X1 U9473 ( .A(n6821), .ZN(n13798) );
  INV_X1 U9474 ( .A(n7262), .ZN(n13727) );
  NAND2_X1 U9475 ( .A1(n7429), .A2(n8564), .ZN(n8956) );
  NAND2_X1 U9476 ( .A1(n12179), .A2(n14863), .ZN(n6861) );
  NAND2_X1 U9477 ( .A1(n6861), .A2(n6860), .ZN(n6859) );
  NAND2_X1 U9478 ( .A1(n7561), .A2(n7432), .ZN(n7430) );
  NAND2_X1 U9479 ( .A1(n6991), .A2(n7239), .ZN(n6988) );
  NAND2_X1 U9480 ( .A1(n7065), .A2(n7068), .ZN(n9070) );
  NAND2_X1 U9481 ( .A1(n7061), .A2(n7063), .ZN(n9128) );
  NAND2_X1 U9482 ( .A1(n6847), .A2(n6846), .ZN(n11365) );
  NAND4_X1 U9483 ( .A1(n8305), .A2(n8306), .A3(n8304), .A4(n7028), .ZN(n7435)
         );
  NAND2_X1 U9484 ( .A1(n9224), .A2(n6511), .ZN(n7509) );
  INV_X1 U9485 ( .A(n10639), .ZN(n7029) );
  NAND2_X1 U9486 ( .A1(n8564), .A2(n7431), .ZN(n8791) );
  CLKBUF_X3 U9487 ( .A(n12604), .Z(n6816) );
  INV_X1 U9488 ( .A(n7514), .ZN(n7512) );
  INV_X1 U9489 ( .A(n7501), .ZN(n12883) );
  NAND2_X1 U9490 ( .A1(n14043), .A2(n14042), .ZN(n14001) );
  XNOR2_X1 U9491 ( .A(n14057), .B(n14056), .ZN(n15144) );
  XNOR2_X1 U9492 ( .A(n7081), .B(n7080), .ZN(SUB_1596_U4) );
  NAND2_X1 U9493 ( .A1(n14339), .A2(n14340), .ZN(n7059) );
  NAND2_X1 U9494 ( .A1(n14044), .A2(n14045), .ZN(n7018) );
  XNOR2_X1 U9495 ( .A(n14041), .B(n7021), .ZN(n15143) );
  NAND2_X1 U9496 ( .A1(n15143), .A2(n15142), .ZN(n7020) );
  NOR2_X1 U9497 ( .A1(n7003), .A2(n8062), .ZN(n7002) );
  INV_X1 U9498 ( .A(n7000), .ZN(n6999) );
  NAND2_X1 U9499 ( .A1(n8702), .A2(n8701), .ZN(n7395) );
  NAND2_X1 U9500 ( .A1(n6843), .A2(n6576), .ZN(n13917) );
  AND2_X1 U9501 ( .A1(n12195), .A2(n14972), .ZN(n7349) );
  NAND2_X1 U9502 ( .A1(n7378), .A2(n7376), .ZN(n14880) );
  NAND2_X1 U9503 ( .A1(n7361), .A2(n7359), .ZN(n12386) );
  INV_X1 U9504 ( .A(n11387), .ZN(n6824) );
  NOR2_X1 U9505 ( .A1(n12559), .A2(n12558), .ZN(n12560) );
  NAND2_X1 U9506 ( .A1(n7301), .A2(n7300), .ZN(n10085) );
  NAND2_X1 U9507 ( .A1(n11240), .A2(n9419), .ZN(n10095) );
  NAND2_X1 U9508 ( .A1(n6827), .A2(n6825), .ZN(P3_U3180) );
  NAND2_X1 U9509 ( .A1(n11964), .A2(n11963), .ZN(n6827) );
  XNOR2_X1 U9510 ( .A(n6452), .B(n9072), .ZN(n9073) );
  NAND2_X1 U9511 ( .A1(n9222), .A2(n6512), .ZN(n7510) );
  NAND2_X1 U9512 ( .A1(n7483), .A2(n7486), .ZN(n7485) );
  NAND2_X1 U9513 ( .A1(n7313), .A2(n7310), .ZN(n10791) );
  INV_X1 U9514 ( .A(n9212), .ZN(n7488) );
  NOR2_X1 U9515 ( .A1(n12049), .A2(n12050), .ZN(n12053) );
  NOR2_X1 U9516 ( .A1(n12009), .A2(n12008), .ZN(n12012) );
  OAI21_X1 U9517 ( .B1(n12180), .B2(n14878), .A(n6858), .ZN(P3_U3201) );
  NAND2_X1 U9518 ( .A1(n13426), .A2(n13427), .ZN(n13282) );
  INV_X1 U9519 ( .A(n7489), .ZN(n7484) );
  INV_X1 U9520 ( .A(n7118), .ZN(n7117) );
  NAND2_X1 U9521 ( .A1(n7067), .A2(n9070), .ZN(n10351) );
  INV_X1 U9522 ( .A(n11364), .ZN(n6847) );
  OR2_X1 U9523 ( .A1(n10349), .A2(n9071), .ZN(n7040) );
  NAND2_X2 U9524 ( .A1(n8143), .A2(n9393), .ZN(n9454) );
  INV_X1 U9525 ( .A(n12743), .ZN(n10420) );
  NAND2_X2 U9526 ( .A1(n6835), .A2(n11433), .ZN(n14468) );
  AOI22_X1 U9527 ( .A1(n13331), .A2(n13484), .B1(n6748), .B2(n13206), .ZN(
        n10113) );
  INV_X2 U9528 ( .A(n11609), .ZN(n9542) );
  INV_X8 U9529 ( .A(n9542), .ZN(n9657) );
  OAI21_X1 U9530 ( .B1(n7119), .B2(n7880), .A(n7879), .ZN(n7118) );
  NAND2_X1 U9531 ( .A1(n12920), .A2(n12909), .ZN(n12904) );
  AND2_X4 U9532 ( .A1(n7852), .A2(n7851), .ZN(n14684) );
  NAND2_X2 U9533 ( .A1(n12967), .A2(n13129), .ZN(n12966) );
  NAND2_X1 U9534 ( .A1(n6907), .A2(n7617), .ZN(n7939) );
  NAND2_X1 U9535 ( .A1(n9131), .A2(n9130), .ZN(n6845) );
  NOR2_X1 U9536 ( .A1(n10358), .A2(n7036), .ZN(n7033) );
  NOR2_X2 U9537 ( .A1(n8791), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n8796) );
  OAI21_X2 U9538 ( .B1(n13409), .B2(n7465), .A(n7463), .ZN(n13426) );
  NAND2_X1 U9539 ( .A1(n7773), .A2(n7589), .ZN(n7776) );
  NAND2_X1 U9540 ( .A1(n7863), .A2(n7862), .ZN(n10389) );
  OAI21_X1 U9541 ( .B1(n11609), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6848), .ZN(
        n7586) );
  NAND2_X1 U9542 ( .A1(n6865), .A2(n6863), .ZN(n11482) );
  NAND2_X1 U9543 ( .A1(n6864), .A2(n11478), .ZN(n6863) );
  NAND2_X1 U9544 ( .A1(n6868), .A2(n11479), .ZN(n6864) );
  INV_X1 U9545 ( .A(n11479), .ZN(n6866) );
  INV_X1 U9546 ( .A(n6868), .ZN(n6867) );
  NAND2_X1 U9547 ( .A1(n7281), .A2(n7284), .ZN(n6868) );
  AND4_X2 U9548 ( .A1(n9545), .A2(n9403), .A3(n9402), .A4(n9815), .ZN(n9408)
         );
  NAND2_X1 U9549 ( .A1(n6871), .A2(n6869), .ZN(n11531) );
  NAND3_X1 U9550 ( .A1(n11501), .A2(n11500), .A3(n6872), .ZN(n6871) );
  NAND2_X1 U9551 ( .A1(n11506), .A2(n11507), .ZN(n6875) );
  NAND2_X1 U9552 ( .A1(n6876), .A2(n6879), .ZN(n7271) );
  NAND2_X1 U9553 ( .A1(n7280), .A2(n6877), .ZN(n6876) );
  NAND2_X1 U9554 ( .A1(n6883), .A2(n6886), .ZN(n11614) );
  NAND3_X1 U9555 ( .A1(n11589), .A2(n6884), .A3(n11588), .ZN(n6883) );
  NAND2_X1 U9556 ( .A1(n6888), .A2(n6889), .ZN(n7291) );
  NAND3_X1 U9557 ( .A1(n11650), .A2(n6891), .A3(n11649), .ZN(n6888) );
  INV_X1 U9558 ( .A(n11664), .ZN(n6892) );
  OAI21_X1 U9559 ( .B1(n11494), .B2(n6897), .A(n6896), .ZN(n11497) );
  NAND2_X1 U9560 ( .A1(n6895), .A2(n6893), .ZN(n11496) );
  NAND2_X1 U9561 ( .A1(n11494), .A2(n6896), .ZN(n6895) );
  NAND2_X1 U9562 ( .A1(n7924), .A2(n6908), .ZN(n6904) );
  NAND2_X1 U9563 ( .A1(n6904), .A2(n6905), .ZN(n7714) );
  NAND2_X1 U9564 ( .A1(n7924), .A2(n7923), .ZN(n6907) );
  XNOR2_X1 U9565 ( .A(n7629), .B(SI_18_), .ZN(n7681) );
  NAND2_X1 U9566 ( .A1(n7757), .A2(n7587), .ZN(n7773) );
  NAND3_X1 U9567 ( .A1(n6915), .A2(n7587), .A3(n7753), .ZN(n7757) );
  INV_X1 U9568 ( .A(n7585), .ZN(n6917) );
  NAND2_X2 U9569 ( .A1(n13984), .A2(n14344), .ZN(n11612) );
  NAND2_X1 U9570 ( .A1(n7188), .A2(n13984), .ZN(n9548) );
  NAND4_X1 U9571 ( .A1(n9408), .A2(n9415), .A3(n6930), .A4(n6555), .ZN(n6929)
         );
  NAND2_X1 U9572 ( .A1(n9407), .A2(n7573), .ZN(n6928) );
  NOR2_X2 U9573 ( .A1(n13832), .A2(n13950), .ZN(n6939) );
  NOR2_X2 U9574 ( .A1(n13874), .A2(n13860), .ZN(n6941) );
  AND2_X2 U9575 ( .A1(n13787), .A2(n6942), .ZN(n13728) );
  NAND2_X1 U9576 ( .A1(n6952), .A2(n6950), .ZN(n14403) );
  INV_X1 U9577 ( .A(n6951), .ZN(n6950) );
  OAI21_X1 U9578 ( .B1(n6953), .B2(n11441), .A(n14401), .ZN(n6951) );
  NAND3_X1 U9579 ( .A1(n10231), .A2(n10230), .A3(n14405), .ZN(n6952) );
  NAND2_X1 U9580 ( .A1(n6954), .A2(n6956), .ZN(n11039) );
  NAND2_X1 U9581 ( .A1(n10994), .A2(n6958), .ZN(n6954) );
  AOI21_X1 U9582 ( .B1(n6958), .B2(n11767), .A(n6957), .ZN(n6956) );
  INV_X1 U9583 ( .A(n9552), .ZN(n9554) );
  NAND2_X1 U9584 ( .A1(n10283), .A2(n6961), .ZN(n6960) );
  NAND3_X1 U9585 ( .A1(n10284), .A2(n6960), .A3(n6475), .ZN(n14388) );
  NAND2_X1 U9586 ( .A1(n10540), .A2(n6964), .ZN(n10601) );
  OAI21_X2 U9587 ( .B1(n6439), .B2(n6990), .A(n6986), .ZN(n13737) );
  NAND2_X1 U9588 ( .A1(n7610), .A2(n6544), .ZN(n6992) );
  NAND2_X1 U9589 ( .A1(n8050), .A2(n7002), .ZN(n6998) );
  OAI21_X1 U9590 ( .B1(n8050), .B2(n7001), .A(n6999), .ZN(n8082) );
  NOR2_X2 U9591 ( .A1(n12966), .A2(n13124), .ZN(n7007) );
  XNOR2_X2 U9592 ( .A(n7647), .B(n7670), .ZN(n8143) );
  OAI21_X1 U9593 ( .B1(n9699), .B2(n7012), .A(n7011), .ZN(n7010) );
  NAND2_X2 U9594 ( .A1(n7760), .A2(n7009), .ZN(n10021) );
  NOR2_X1 U9595 ( .A1(n10429), .A2(n14659), .ZN(n10468) );
  AND2_X2 U9596 ( .A1(n7797), .A2(n7796), .ZN(n10383) );
  NAND3_X1 U9597 ( .A1(n7028), .A2(P3_IR_REG_19__SCAN_IN), .A3(n7026), .ZN(
        n7022) );
  INV_X1 U9598 ( .A(n10358), .ZN(n7039) );
  INV_X1 U9599 ( .A(n7040), .ZN(n10357) );
  OR2_X1 U9600 ( .A1(n9074), .A2(n14921), .ZN(n7038) );
  NAND2_X1 U9601 ( .A1(n11961), .A2(n6547), .ZN(n7041) );
  OAI211_X1 U9602 ( .C1(n11961), .C2(n7043), .A(n11963), .B(n7041), .ZN(n9172)
         );
  NAND2_X1 U9603 ( .A1(n11961), .A2(n11962), .ZN(n11960) );
  AND2_X1 U9604 ( .A1(n9145), .A2(n7049), .ZN(n7048) );
  OR2_X1 U9605 ( .A1(n11962), .A2(n9144), .ZN(n7049) );
  NAND3_X1 U9606 ( .A1(n9061), .A2(n9068), .A3(n9062), .ZN(n7068) );
  NAND3_X1 U9607 ( .A1(n9066), .A2(n9062), .A3(n9061), .ZN(n7066) );
  INV_X1 U9608 ( .A(n7072), .ZN(n14326) );
  AOI21_X1 U9609 ( .B1(n14332), .B2(n14333), .A(P2_ADDR_REG_14__SCAN_IN), .ZN(
        n7069) );
  NAND2_X1 U9610 ( .A1(n7071), .A2(n14329), .ZN(n7070) );
  NAND2_X1 U9611 ( .A1(n14327), .A2(n14328), .ZN(n7071) );
  INV_X1 U9612 ( .A(n8264), .ZN(n7085) );
  INV_X1 U9613 ( .A(n8287), .ZN(n7094) );
  OAI21_X1 U9614 ( .B1(n8715), .B2(n7095), .A(n7093), .ZN(n8738) );
  OAI21_X1 U9615 ( .B1(n8694), .B2(n8693), .A(n8285), .ZN(n8704) );
  AOI21_X1 U9616 ( .B1(n8693), .B2(n8285), .A(n7100), .ZN(n7099) );
  NAND2_X1 U9617 ( .A1(n8751), .A2(n7113), .ZN(n7111) );
  NOR2_X2 U9618 ( .A1(n14148), .A2(n8639), .ZN(n14147) );
  XNOR2_X2 U9619 ( .A(n12129), .B(n14157), .ZN(n14148) );
  NAND2_X1 U9620 ( .A1(n12030), .A2(n6578), .ZN(n7130) );
  OAI211_X1 U9621 ( .C1(n12030), .C2(n12061), .A(n7131), .B(n7130), .ZN(n12031) );
  NAND2_X1 U9622 ( .A1(n12079), .A2(n12112), .ZN(n7137) );
  NAND3_X1 U9623 ( .A1(n7140), .A2(n7141), .A3(n7137), .ZN(n12080) );
  NAND2_X1 U9624 ( .A1(n6440), .A2(n12084), .ZN(n12102) );
  OR2_X1 U9625 ( .A1(n12084), .A2(n12087), .ZN(n7141) );
  INV_X1 U9626 ( .A(n14659), .ZN(n10431) );
  INV_X1 U9627 ( .A(n7156), .ZN(n14785) );
  INV_X1 U9628 ( .A(n10899), .ZN(n7155) );
  INV_X1 U9629 ( .A(n7163), .ZN(n12958) );
  NAND2_X1 U9630 ( .A1(n13726), .A2(n6481), .ZN(n13725) );
  OAI21_X1 U9631 ( .B1(n10252), .B2(n7181), .A(n7179), .ZN(n14379) );
  NAND2_X1 U9632 ( .A1(n7178), .A2(n6503), .ZN(n10268) );
  NAND2_X1 U9633 ( .A1(n7179), .A2(n7181), .ZN(n7177) );
  NAND2_X1 U9634 ( .A1(n10252), .A2(n7179), .ZN(n7178) );
  NAND2_X1 U9635 ( .A1(n10999), .A2(n7183), .ZN(n7182) );
  INV_X1 U9636 ( .A(n14344), .ZN(n7189) );
  INV_X2 U9637 ( .A(n11612), .ZN(n11556) );
  NAND2_X2 U9638 ( .A1(n9541), .A2(n6434), .ZN(n14344) );
  NAND2_X1 U9639 ( .A1(n10409), .A2(n7190), .ZN(n7191) );
  NAND3_X1 U9640 ( .A1(n7200), .A2(n7199), .A3(n7478), .ZN(n9539) );
  OAI21_X1 U9641 ( .B1(n11232), .B2(n7205), .A(n7201), .ZN(n13873) );
  INV_X2 U9642 ( .A(n7445), .ZN(n9925) );
  NAND2_X1 U9643 ( .A1(n13811), .A2(n7210), .ZN(n7209) );
  NAND2_X2 U9644 ( .A1(n12128), .A2(n12127), .ZN(n12129) );
  NAND2_X1 U9645 ( .A1(n8284), .A2(n8283), .ZN(n8694) );
  NAND2_X1 U9646 ( .A1(n8277), .A2(n8276), .ZN(n8660) );
  NAND2_X1 U9647 ( .A1(n8660), .A2(n8659), .ZN(n8280) );
  NAND2_X1 U9648 ( .A1(n8646), .A2(n8275), .ZN(n8277) );
  NOR2_X2 U9649 ( .A1(n14537), .A2(n10607), .ZN(n11001) );
  NOR2_X2 U9650 ( .A1(n14394), .A2(n14393), .ZN(n14395) );
  NOR2_X4 U9651 ( .A1(n13801), .A2(n13793), .ZN(n13787) );
  NAND2_X1 U9652 ( .A1(n7223), .A2(n13653), .ZN(n7222) );
  NAND3_X1 U9653 ( .A1(n14140), .A2(P3_ADDR_REG_19__SCAN_IN), .A3(n7216), .ZN(
        n7579) );
  INV_X2 U9654 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n14140) );
  MUX2_X1 U9655 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n9542), .Z(n7218) );
  NAND3_X1 U9656 ( .A1(n7225), .A2(n7233), .A3(n7222), .ZN(n13895) );
  NAND3_X1 U9657 ( .A1(n7225), .A2(n7224), .A3(n7222), .ZN(n7228) );
  OAI211_X1 U9658 ( .C1(n7231), .C2(n7230), .A(n7228), .B(n7226), .ZN(P1_U3525) );
  INV_X1 U9659 ( .A(n13893), .ZN(n7236) );
  NOR2_X1 U9660 ( .A1(n13785), .A2(n7243), .ZN(n7238) );
  INV_X1 U9661 ( .A(n7247), .ZN(n7246) );
  NOR2_X1 U9662 ( .A1(n13939), .A2(n13666), .ZN(n7247) );
  NAND2_X1 U9663 ( .A1(n7610), .A2(n7609), .ZN(n7898) );
  NAND2_X1 U9664 ( .A1(n7939), .A2(n7938), .ZN(n7256) );
  NOR2_X1 U9665 ( .A1(n7264), .A2(n7263), .ZN(n7262) );
  AND2_X1 U9666 ( .A1(n13919), .A2(n13670), .ZN(n7268) );
  NAND2_X1 U9667 ( .A1(n7271), .A2(n6557), .ZN(n11750) );
  NAND2_X1 U9668 ( .A1(n11750), .A2(n6559), .ZN(n7279) );
  NAND2_X1 U9669 ( .A1(n7279), .A2(n7274), .ZN(n11790) );
  NAND3_X1 U9670 ( .A1(n11698), .A2(n6558), .A3(n11697), .ZN(n7280) );
  NAND3_X1 U9671 ( .A1(n11475), .A2(n7282), .A3(n11474), .ZN(n7281) );
  NAND2_X1 U9672 ( .A1(n7289), .A2(n7287), .ZN(n11645) );
  NAND3_X1 U9673 ( .A1(n7290), .A2(n11618), .A3(n11617), .ZN(n7289) );
  NAND2_X1 U9674 ( .A1(n7291), .A2(n7292), .ZN(n11693) );
  INV_X1 U9675 ( .A(n7295), .ZN(n10127) );
  NAND2_X1 U9676 ( .A1(n7655), .A2(n8137), .ZN(n8132) );
  NOR2_X1 U9677 ( .A1(n10042), .A2(n10041), .ZN(n10044) );
  INV_X1 U9678 ( .A(n10086), .ZN(n7303) );
  INV_X1 U9679 ( .A(n10790), .ZN(n7317) );
  NAND2_X1 U9680 ( .A1(n12534), .A2(n7320), .ZN(n7318) );
  NOR2_X1 U9681 ( .A1(n6519), .A2(n12532), .ZN(n7320) );
  OR2_X1 U9682 ( .A1(n12535), .A2(n7323), .ZN(n7322) );
  INV_X1 U9683 ( .A(n12714), .ZN(n7323) );
  NAND2_X1 U9684 ( .A1(n12704), .A2(n7336), .ZN(n7335) );
  OAI211_X1 U9685 ( .C1(n12704), .C2(n7337), .A(n12610), .B(n7335), .ZN(
        P2_U3192) );
  NAND2_X1 U9686 ( .A1(n12704), .A2(n12575), .ZN(n12601) );
  INV_X1 U9687 ( .A(n12606), .ZN(n7346) );
  NAND2_X1 U9688 ( .A1(n7347), .A2(n14904), .ZN(n8404) );
  INV_X1 U9689 ( .A(n14905), .ZN(n7347) );
  NAND3_X1 U9690 ( .A1(n10644), .A2(n10918), .A3(n7348), .ZN(n8931) );
  NOR2_X1 U9691 ( .A1(n8988), .A2(n14905), .ZN(n7348) );
  INV_X1 U9692 ( .A(n7350), .ZN(n12197) );
  NOR2_X1 U9693 ( .A1(n7350), .A2(n7349), .ZN(n9183) );
  NAND2_X1 U9694 ( .A1(n12355), .A2(n7356), .ZN(n7353) );
  NAND2_X1 U9695 ( .A1(n7353), .A2(n7354), .ZN(n12330) );
  NAND2_X1 U9696 ( .A1(n11357), .A2(n7362), .ZN(n7361) );
  NAND2_X1 U9697 ( .A1(n11352), .A2(n7367), .ZN(n7366) );
  NAND2_X1 U9698 ( .A1(n12373), .A2(n7373), .ZN(n7372) );
  NAND2_X1 U9699 ( .A1(n10946), .A2(n7379), .ZN(n7378) );
  NAND2_X1 U9700 ( .A1(n12234), .A2(n7386), .ZN(n7385) );
  NAND2_X1 U9701 ( .A1(n12234), .A2(n7391), .ZN(n7388) );
  OAI21_X1 U9702 ( .B1(n12234), .B2(n7387), .A(n7386), .ZN(n12200) );
  NAND2_X1 U9703 ( .A1(n12475), .A2(n12226), .ZN(n7393) );
  OR2_X1 U9704 ( .A1(n11959), .A2(n12236), .ZN(n7394) );
  AOI21_X2 U9705 ( .B1(n7400), .B2(n7399), .A(n7398), .ZN(n8789) );
  OAI21_X1 U9706 ( .B1(n11152), .B2(n8835), .A(n8837), .ZN(n11245) );
  NAND2_X1 U9707 ( .A1(n7417), .A2(n7418), .ZN(n12235) );
  NAND2_X1 U9708 ( .A1(n9013), .A2(n7420), .ZN(n7417) );
  NAND2_X1 U9709 ( .A1(n8313), .A2(n7439), .ZN(n8344) );
  NAND2_X1 U9710 ( .A1(n8313), .A2(n8312), .ZN(n8320) );
  NAND2_X1 U9711 ( .A1(n7441), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U9712 ( .A1(n13485), .A2(n13206), .ZN(n7442) );
  NAND2_X1 U9713 ( .A1(n11059), .A2(n11060), .ZN(n7454) );
  NAND2_X1 U9714 ( .A1(n6434), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9536) );
  OAI21_X1 U9715 ( .B1(n12941), .B2(n7494), .A(n7492), .ZN(n7501) );
  NAND2_X1 U9716 ( .A1(n9224), .A2(n9223), .ZN(n7507) );
  NAND2_X1 U9717 ( .A1(n9222), .A2(n9221), .ZN(n7508) );
  NAND2_X1 U9718 ( .A1(n7512), .A2(n8166), .ZN(n7511) );
  NAND2_X1 U9719 ( .A1(n9239), .A2(n7517), .ZN(n7515) );
  INV_X1 U9720 ( .A(n9241), .ZN(n7527) );
  INV_X1 U9721 ( .A(n7531), .ZN(n7529) );
  NAND2_X1 U9722 ( .A1(n10417), .A2(n7542), .ZN(n7541) );
  NAND3_X1 U9723 ( .A1(n9284), .A2(n9283), .A3(n6577), .ZN(n7545) );
  INV_X1 U9724 ( .A(n9286), .ZN(n7547) );
  AND2_X1 U9725 ( .A1(n9275), .A2(n9274), .ZN(n9276) );
  NAND2_X1 U9726 ( .A1(n13062), .A2(n7557), .ZN(n8183) );
  NAND3_X1 U9727 ( .A1(n7581), .A2(n7580), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7582) );
  NAND2_X1 U9728 ( .A1(n13101), .A2(n13100), .ZN(n13173) );
  INV_X1 U9729 ( .A(n13099), .ZN(n13100) );
  INV_X1 U9730 ( .A(n11833), .ZN(n11834) );
  OAI21_X1 U9731 ( .B1(n13098), .B2(n14655), .A(n13097), .ZN(n13099) );
  XNOR2_X1 U9732 ( .A(n8046), .B(n8047), .ZN(n11640) );
  INV_X1 U9733 ( .A(n11730), .ZN(n11711) );
  NAND2_X1 U9734 ( .A1(n6447), .A2(n7012), .ZN(n8400) );
  INV_X1 U9735 ( .A(n8344), .ZN(n8316) );
  OAI22_X2 U9736 ( .A1(n13869), .A2(n13660), .B1(n14209), .B2(n13659), .ZN(
        n13847) );
  OR2_X1 U9737 ( .A1(n7683), .A2(n8205), .ZN(n8221) );
  NAND2_X1 U9738 ( .A1(n14905), .A2(n14900), .ZN(n14899) );
  INV_X1 U9739 ( .A(n12557), .ZN(n12559) );
  INV_X4 U9740 ( .A(n9213), .ZN(n9342) );
  AND2_X2 U9741 ( .A1(n9186), .A2(n9343), .ZN(n9213) );
  INV_X1 U9742 ( .A(n12334), .ZN(n9005) );
  NAND2_X1 U9743 ( .A1(n14990), .A2(n14960), .ZN(n12459) );
  INV_X1 U9744 ( .A(n12459), .ZN(n9055) );
  AND2_X2 U9745 ( .A1(n10627), .A2(n9052), .ZN(n14990) );
  OR2_X1 U9746 ( .A1(n10204), .A2(n10203), .ZN(n7560) );
  OR2_X1 U9747 ( .A1(n14633), .A2(n8235), .ZN(n14735) );
  AND4_X1 U9748 ( .A1(n8309), .A2(n8795), .A3(n8308), .A4(n8307), .ZN(n7561)
         );
  AND3_X1 U9749 ( .A1(n8130), .A2(n8137), .A3(n8136), .ZN(n7562) );
  OR2_X1 U9750 ( .A1(n9279), .A2(n13005), .ZN(n7563) );
  NAND2_X1 U9751 ( .A1(n8929), .A2(n8928), .ZN(n7564) );
  INV_X1 U9752 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8343) );
  AND2_X1 U9753 ( .A1(n12286), .A2(n11987), .ZN(n7565) );
  OR2_X1 U9754 ( .A1(n12286), .A2(n11987), .ZN(n7566) );
  OR2_X1 U9755 ( .A1(n14973), .A2(n14915), .ZN(n12510) );
  INV_X1 U9756 ( .A(n12510), .ZN(n9184) );
  AND4_X1 U9757 ( .A1(n7649), .A2(n7652), .A3(n7651), .A4(n7650), .ZN(n7567)
         );
  NOR2_X1 U9758 ( .A1(n11854), .A2(n11849), .ZN(n7569) );
  AND3_X1 U9759 ( .A1(n9384), .A2(n11202), .A3(n10418), .ZN(n7570) );
  AND3_X1 U9760 ( .A1(n9328), .A2(n9327), .A3(n9326), .ZN(n7571) );
  NAND4_X1 U9761 ( .A1(n11572), .A2(n11571), .A3(n11570), .A4(n11569), .ZN(
        n7572) );
  NOR3_X1 U9762 ( .A1(n11529), .A2(n11528), .A3(n11547), .ZN(n7574) );
  NAND2_X1 U9763 ( .A1(n11992), .A2(n11171), .ZN(n7575) );
  AND2_X1 U9764 ( .A1(n7621), .A2(n7622), .ZN(n7576) );
  OR2_X1 U9765 ( .A1(n12885), .A2(n12884), .ZN(n7577) );
  INV_X2 U9766 ( .A(n14439), .ZN(n14420) );
  INV_X1 U9767 ( .A(n9862), .ZN(n9929) );
  MUX2_X1 U9768 ( .A(n14485), .B(n13483), .S(n11738), .Z(n11458) );
  OAI22_X1 U9769 ( .A1(n14676), .A2(n6445), .B1(n10453), .B2(n9342), .ZN(n9216) );
  INV_X1 U9770 ( .A(n9220), .ZN(n9224) );
  AOI21_X1 U9771 ( .B1(n11574), .B2(n11573), .A(n7572), .ZN(n11585) );
  AOI22_X1 U9772 ( .A1(n11406), .A2(n9213), .B1(n12731), .B2(n9342), .ZN(n9247) );
  NOR2_X1 U9773 ( .A1(n14404), .A2(n11444), .ZN(n11759) );
  INV_X1 U9774 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8307) );
  INV_X1 U9775 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n8304) );
  INV_X1 U9776 ( .A(n9066), .ZN(n8403) );
  INV_X1 U9777 ( .A(n10744), .ZN(n7895) );
  INV_X1 U9778 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n7635) );
  AND2_X1 U9779 ( .A1(n9858), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n9859) );
  AOI21_X1 U9780 ( .B1(n13206), .B2(n6972), .A(n9859), .ZN(n9860) );
  INV_X1 U9781 ( .A(n8754), .ZN(n8342) );
  INV_X1 U9782 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U9783 ( .A1(n8463), .A2(n8249), .ZN(n8251) );
  INV_X1 U9784 ( .A(n7952), .ZN(n7664) );
  OR2_X1 U9785 ( .A1(n8070), .A2(n8069), .ZN(n8087) );
  NOR2_X1 U9786 ( .A1(n10115), .A2(n10114), .ZN(n10116) );
  INV_X1 U9787 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10398) );
  INV_X1 U9788 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10273) );
  INV_X1 U9789 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9653) );
  INV_X1 U9790 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8325) );
  CLKBUF_X1 U9791 ( .A(n11974), .Z(n11940) );
  INV_X1 U9792 ( .A(n12239), .ZN(n8942) );
  NAND2_X1 U9793 ( .A1(n11378), .A2(n11377), .ZN(n11376) );
  NAND2_X1 U9794 ( .A1(n9704), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8255) );
  NAND2_X1 U9795 ( .A1(n9711), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8244) );
  OR2_X1 U9796 ( .A1(n10930), .A2(n10929), .ZN(n10931) );
  OR2_X1 U9797 ( .A1(n7739), .A2(n7719), .ZN(n7721) );
  NAND2_X1 U9798 ( .A1(n7665), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n7709) );
  NAND2_X1 U9799 ( .A1(n7662), .A2(n7661), .ZN(n7930) );
  NOR2_X1 U9800 ( .A1(n7571), .A2(n9350), .ZN(n9351) );
  NOR2_X1 U9801 ( .A1(n8087), .A2(n12577), .ZN(n8104) );
  OR2_X1 U9802 ( .A1(n8001), .A2(n8000), .ZN(n8015) );
  OR2_X1 U9803 ( .A1(n7954), .A2(n7737), .ZN(n7739) );
  XNOR2_X1 U9804 ( .A(n12858), .B(n12869), .ZN(n9377) );
  NAND2_X1 U9805 ( .A1(n8013), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n8038) );
  NAND2_X1 U9806 ( .A1(n7968), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7984) );
  INV_X1 U9807 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7670) );
  INV_X1 U9808 ( .A(n10116), .ZN(n10117) );
  OR2_X1 U9809 ( .A1(n13220), .A2(n13219), .ZN(n13221) );
  INV_X1 U9810 ( .A(n10489), .ZN(n10486) );
  AND2_X1 U9811 ( .A1(n14217), .A2(n14218), .ZN(n13217) );
  OAI22_X1 U9812 ( .A1(n10215), .A2(n13364), .B1(n9925), .B2(n13264), .ZN(
        n10003) );
  OR2_X1 U9813 ( .A1(n11559), .A2(n11538), .ZN(n11575) );
  NOR2_X1 U9814 ( .A1(n10274), .A2(n10273), .ZN(n10287) );
  INV_X1 U9815 ( .A(n11762), .ZN(n10396) );
  NAND2_X1 U9816 ( .A1(n7714), .A2(n7713), .ZN(n7627) );
  NAND2_X1 U9817 ( .A1(n7604), .A2(SI_8_), .ZN(n7606) );
  NOR2_X2 U9818 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n9545) );
  NOR2_X1 U9819 ( .A1(n14073), .A2(n14072), .ZN(n14018) );
  OR2_X1 U9820 ( .A1(n6787), .A2(n11015), .ZN(n8726) );
  INV_X1 U9821 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n11302) );
  NAND2_X1 U9822 ( .A1(n12308), .A2(n8883), .ZN(n12297) );
  INV_X1 U9823 ( .A(n9004), .ZN(n12348) );
  INV_X1 U9824 ( .A(n14919), .ZN(n14903) );
  INV_X1 U9825 ( .A(n10134), .ZN(n8662) );
  NAND2_X1 U9826 ( .A1(n9165), .A2(n10132), .ZN(n14901) );
  AND2_X1 U9827 ( .A1(n8268), .A2(n8267), .ZN(n8598) );
  INV_X1 U9828 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n8492) );
  AND2_X1 U9829 ( .A1(n8246), .A2(n8245), .ZN(n8428) );
  AND2_X1 U9830 ( .A1(n10942), .A2(n10583), .ZN(n9956) );
  NAND2_X1 U9831 ( .A1(n7660), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7853) );
  INV_X1 U9832 ( .A(n8194), .ZN(n9952) );
  OR2_X1 U9833 ( .A1(n12936), .A2(n7763), .ZN(n8045) );
  INV_X1 U9834 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10525) );
  OR2_X1 U9835 ( .A1(n9902), .A2(n9901), .ZN(n9900) );
  INV_X1 U9836 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9971) );
  OR2_X1 U9837 ( .A1(n10370), .A2(n14636), .ZN(n10371) );
  INV_X1 U9838 ( .A(n14715), .ZN(n14660) );
  INV_X1 U9839 ( .A(n9943), .ZN(n9954) );
  AND2_X1 U9840 ( .A1(n13396), .A2(n13315), .ZN(n13417) );
  AND2_X1 U9841 ( .A1(n13344), .A2(n13297), .ZN(n13442) );
  OR2_X1 U9842 ( .A1(n11029), .A2(n11028), .ZN(n11041) );
  AND2_X1 U9843 ( .A1(n11602), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11619) );
  AND2_X1 U9844 ( .A1(n11590), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11602) );
  AND2_X1 U9845 ( .A1(n9677), .A2(n11293), .ZN(n9419) );
  INV_X1 U9846 ( .A(n13650), .ZN(n13721) );
  INV_X1 U9847 ( .A(n13860), .ZN(n14257) );
  OR2_X1 U9848 ( .A1(n10212), .A2(n14414), .ZN(n14509) );
  INV_X1 U9849 ( .A(n14429), .ZN(n14540) );
  NAND2_X1 U9850 ( .A1(n8008), .A2(n8007), .ZN(n8010) );
  XNOR2_X1 U9851 ( .A(n7618), .B(SI_13_), .ZN(n7938) );
  XNOR2_X1 U9852 ( .A(n7614), .B(SI_11_), .ZN(n7908) );
  OAI21_X1 U9853 ( .B1(P3_ADDR_REG_11__SCAN_IN), .B2(n14022), .A(n14021), .ZN(
        n14079) );
  NAND2_X1 U9854 ( .A1(n9152), .A2(n9151), .ZN(n11963) );
  INV_X1 U9855 ( .A(n6449), .ZN(n8772) );
  AND4_X1 U9856 ( .A1(n8631), .A2(n8630), .A3(n8629), .A4(n8628), .ZN(n12368)
         );
  INV_X1 U9857 ( .A(n14741), .ZN(n14874) );
  INV_X1 U9858 ( .A(n14901), .ZN(n14920) );
  INV_X1 U9859 ( .A(n14891), .ZN(n14923) );
  NOR2_X1 U9860 ( .A1(n14990), .A2(n9053), .ZN(n9054) );
  AND2_X1 U9861 ( .A1(n9043), .A2(n9042), .ZN(n10627) );
  INV_X1 U9862 ( .A(n14915), .ZN(n14960) );
  OR2_X1 U9863 ( .A1(n14906), .A2(n14968), .ZN(n14972) );
  AND2_X1 U9864 ( .A1(n14911), .A2(n9047), .ZN(n14968) );
  XNOR2_X1 U9865 ( .A(n8954), .B(n8953), .ZN(n10131) );
  NOR2_X1 U9866 ( .A1(n8311), .A2(n8957), .ZN(n8958) );
  INV_X1 U9867 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n8377) );
  AND2_X1 U9868 ( .A1(n9961), .A2(n9956), .ZN(n12717) );
  NAND2_X1 U9869 ( .A1(n9955), .A2(n12998), .ZN(n12722) );
  AND2_X1 U9870 ( .A1(n8045), .A2(n8044), .ZN(n12631) );
  AND4_X1 U9871 ( .A1(n7949), .A2(n7948), .A3(n7947), .A4(n7946), .ZN(n11418)
         );
  AND2_X1 U9872 ( .A1(n9978), .A2(n9439), .ZN(n10071) );
  AND2_X1 U9873 ( .A1(n9507), .A2(n9506), .ZN(n14579) );
  AND2_X1 U9874 ( .A1(n13038), .A2(n10583), .ZN(n13085) );
  NAND2_X1 U9875 ( .A1(n9343), .A2(n10942), .ZN(n14688) );
  OR2_X1 U9876 ( .A1(n10774), .A2(n11086), .ZN(n14717) );
  AOI21_X1 U9877 ( .B1(n8217), .B2(n11295), .A(n13203), .ZN(n14630) );
  AND2_X1 U9878 ( .A1(n7885), .A2(n7910), .ZN(n9484) );
  AND3_X1 U9879 ( .A1(n11542), .A2(n11541), .A3(n11540), .ZN(n13848) );
  AND2_X1 U9880 ( .A1(n9737), .A2(n9736), .ZN(n9760) );
  INV_X1 U9881 ( .A(n14354), .ZN(n14367) );
  INV_X1 U9882 ( .A(n14375), .ZN(n14357) );
  INV_X1 U9883 ( .A(n14360), .ZN(n14370) );
  INV_X1 U9884 ( .A(n13663), .ZN(n13816) );
  INV_X1 U9885 ( .A(n13875), .ZN(n14436) );
  INV_X1 U9886 ( .A(n13844), .ZN(n14252) );
  AND2_X1 U9887 ( .A1(n14509), .A2(n14523), .ZN(n14489) );
  NAND2_X1 U9888 ( .A1(n11739), .A2(n9579), .ZN(n14429) );
  INV_X1 U9889 ( .A(n14489), .ZN(n14544) );
  INV_X1 U9890 ( .A(n9880), .ZN(n9918) );
  AND2_X1 U9891 ( .A1(n10095), .A2(n9678), .ZN(n9866) );
  AND2_X1 U9892 ( .A1(n10147), .A2(n10146), .ZN(n14871) );
  INV_X1 U9893 ( .A(n11972), .ZN(n11373) );
  INV_X1 U9894 ( .A(n8785), .ZN(n12183) );
  INV_X1 U9895 ( .A(n12368), .ZN(n12345) );
  INV_X1 U9896 ( .A(n9066), .ZN(n11996) );
  INV_X1 U9897 ( .A(n14871), .ZN(n14837) );
  OR2_X1 U9898 ( .A1(n10140), .A2(n10139), .ZN(n14878) );
  INV_X1 U9899 ( .A(n12463), .ZN(n12190) );
  AND2_X1 U9900 ( .A1(n11355), .A2(n11354), .ZN(n14169) );
  NAND2_X1 U9901 ( .A1(n10629), .A2(n12271), .ZN(n14933) );
  AOI21_X1 U9902 ( .B1(n8787), .B2(n9055), .A(n9054), .ZN(n9056) );
  INV_X1 U9903 ( .A(n14990), .ZN(n14987) );
  AND2_X1 U9904 ( .A1(n14170), .A2(n14169), .ZN(n14177) );
  AND2_X1 U9905 ( .A1(n9182), .A2(n9181), .ZN(n14973) );
  OR2_X1 U9906 ( .A1(n11424), .A2(n11423), .ZN(n11425) );
  AND2_X1 U9907 ( .A1(n10131), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12513) );
  INV_X1 U9908 ( .A(n10628), .ZN(n10196) );
  OR2_X1 U9909 ( .A1(n8568), .A2(n8567), .ZN(n12036) );
  NAND2_X1 U9910 ( .A1(n9961), .A2(n9960), .ZN(n12724) );
  NAND2_X1 U9911 ( .A1(n8114), .A2(n8113), .ZN(n12887) );
  INV_X1 U9912 ( .A(n11288), .ZN(n12734) );
  INV_X1 U9913 ( .A(n10591), .ZN(n12739) );
  INV_X1 U9914 ( .A(n14579), .ZN(n14620) );
  INV_X1 U9915 ( .A(n14577), .ZN(n14628) );
  NAND2_X1 U9916 ( .A1(n13038), .A2(n10373), .ZN(n13053) );
  INV_X1 U9917 ( .A(n14723), .ZN(n14721) );
  INV_X1 U9918 ( .A(n14631), .ZN(n14632) );
  OR2_X1 U9919 ( .A1(n10368), .A2(n14635), .ZN(n14633) );
  INV_X1 U9920 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10081) );
  OR2_X1 U9921 ( .A1(n13463), .A2(n14380), .ZN(n14215) );
  INV_X1 U9922 ( .A(n13793), .ZN(n13939) );
  OR2_X1 U9923 ( .A1(n9869), .A2(n9868), .ZN(n14221) );
  INV_X1 U9924 ( .A(n13675), .ZN(n13472) );
  OR2_X1 U9925 ( .A1(n11227), .A2(n11226), .ZN(n13866) );
  OR2_X1 U9926 ( .A1(n14348), .A2(n9729), .ZN(n14360) );
  OR2_X1 U9927 ( .A1(n14348), .A2(n13505), .ZN(n14375) );
  NAND2_X1 U9928 ( .A1(n14420), .A2(n10213), .ZN(n13844) );
  NAND2_X1 U9929 ( .A1(n13904), .A2(n13903), .ZN(n13963) );
  AND2_X1 U9930 ( .A1(n14290), .A2(n14289), .ZN(n14313) );
  AND2_X2 U9931 ( .A1(n9919), .A2(n9918), .ZN(n14546) );
  INV_X1 U9932 ( .A(n11430), .ZN(n13995) );
  INV_X1 U9933 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10129) );
  INV_X1 U9934 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9914) );
  INV_X2 U9935 ( .A(n11997), .ZN(P3_U3897) );
  AND2_X1 U9936 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9452), .ZN(P2_U3947) );
  OR3_X1 U9937 ( .A1(n9516), .A2(n12594), .A3(n9515), .ZN(P2_U3233) );
  INV_X1 U9938 ( .A(n14991), .ZN(P1_U4016) );
  NAND2_X1 U9939 ( .A1(n7579), .A2(n7578), .ZN(n7584) );
  NAND2_X1 U9940 ( .A1(n7582), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n7583) );
  NAND2_X4 U9941 ( .A1(n7584), .A2(n7583), .ZN(n11609) );
  NAND2_X1 U9942 ( .A1(n7585), .A2(SI_1_), .ZN(n7587) );
  INV_X1 U9943 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8387) );
  INV_X1 U9944 ( .A(SI_0_), .ZN(n9629) );
  NOR2_X1 U9945 ( .A1(n7586), .A2(n9629), .ZN(n7753) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n11609), .Z(n7588) );
  NAND2_X1 U9947 ( .A1(n7588), .A2(SI_2_), .ZN(n7590) );
  INV_X1 U9948 ( .A(n7774), .ZN(n7589) );
  NAND2_X1 U9949 ( .A1(n7776), .A2(n7590), .ZN(n7793) );
  NAND2_X1 U9950 ( .A1(n7793), .A2(n7792), .ZN(n7795) );
  NAND2_X1 U9951 ( .A1(n7795), .A2(n7591), .ZN(n7805) );
  NAND2_X1 U9952 ( .A1(n7592), .A2(SI_4_), .ZN(n7594) );
  OAI21_X1 U9953 ( .B1(n7592), .B2(SI_4_), .A(n7594), .ZN(n7593) );
  INV_X1 U9954 ( .A(n7593), .ZN(n7804) );
  NAND2_X1 U9955 ( .A1(n7805), .A2(n7804), .ZN(n7807) );
  MUX2_X1 U9956 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9657), .Z(n7595) );
  NAND2_X1 U9957 ( .A1(n7595), .A2(SI_5_), .ZN(n7597) );
  OAI21_X1 U9958 ( .B1(SI_5_), .B2(n7595), .A(n7597), .ZN(n7814) );
  INV_X1 U9959 ( .A(n7814), .ZN(n7596) );
  MUX2_X1 U9960 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9657), .Z(n7598) );
  NAND2_X1 U9961 ( .A1(n7598), .A2(SI_6_), .ZN(n7600) );
  OAI21_X1 U9962 ( .B1(SI_6_), .B2(n7598), .A(n7600), .ZN(n7599) );
  INV_X1 U9963 ( .A(n7599), .ZN(n7827) );
  MUX2_X1 U9964 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n11609), .Z(n7601) );
  NAND2_X1 U9965 ( .A1(n7601), .A2(SI_7_), .ZN(n7603) );
  OAI21_X1 U9966 ( .B1(n7601), .B2(SI_7_), .A(n7603), .ZN(n7602) );
  INV_X1 U9967 ( .A(n7602), .ZN(n7844) );
  MUX2_X1 U9968 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n11609), .Z(n7604) );
  OAI21_X1 U9969 ( .B1(SI_8_), .B2(n7604), .A(n7606), .ZN(n7605) );
  INV_X1 U9970 ( .A(n7605), .ZN(n7861) );
  MUX2_X1 U9971 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n11609), .Z(n7607) );
  INV_X1 U9972 ( .A(n7881), .ZN(n7608) );
  MUX2_X1 U9973 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n11609), .Z(n7611) );
  OAI21_X1 U9974 ( .B1(n7611), .B2(SI_10_), .A(n7613), .ZN(n7612) );
  INV_X1 U9975 ( .A(n7612), .ZN(n7897) );
  MUX2_X1 U9976 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n11609), .Z(n7614) );
  INV_X1 U9977 ( .A(n7614), .ZN(n7615) );
  INV_X1 U9978 ( .A(SI_11_), .ZN(n9660) );
  MUX2_X1 U9979 ( .A(n9914), .B(n9924), .S(n11609), .Z(n7616) );
  INV_X1 U9980 ( .A(SI_12_), .ZN(n9673) );
  NAND2_X1 U9981 ( .A1(n7616), .A2(n9673), .ZN(n7617) );
  MUX2_X1 U9982 ( .A(n9991), .B(n10012), .S(n11609), .Z(n7618) );
  INV_X1 U9983 ( .A(SI_13_), .ZN(n9713) );
  NAND2_X1 U9984 ( .A1(n7618), .A2(n9713), .ZN(n7619) );
  MUX2_X1 U9985 ( .A(n10079), .B(n10083), .S(n11609), .Z(n7745) );
  NAND2_X1 U9986 ( .A1(n7727), .A2(SI_14_), .ZN(n7621) );
  MUX2_X1 U9987 ( .A(n10176), .B(n10178), .S(n11609), .Z(n7728) );
  INV_X1 U9988 ( .A(n7728), .ZN(n7620) );
  NOR2_X1 U9989 ( .A1(n7727), .A2(SI_14_), .ZN(n7623) );
  INV_X1 U9990 ( .A(SI_15_), .ZN(n9813) );
  AOI22_X1 U9991 ( .A1(n7623), .A2(n7622), .B1(n9813), .B2(n7728), .ZN(n7624)
         );
  MUX2_X1 U9992 ( .A(n10076), .B(n10081), .S(n11609), .Z(n7625) );
  INV_X1 U9993 ( .A(SI_16_), .ZN(n9844) );
  NAND2_X1 U9994 ( .A1(n7625), .A2(n9844), .ZN(n7626) );
  INV_X1 U9995 ( .A(SI_17_), .ZN(n9938) );
  INV_X1 U9996 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10171) );
  MUX2_X1 U9997 ( .A(n10129), .B(n10171), .S(n9657), .Z(n7697) );
  INV_X1 U9998 ( .A(n7697), .ZN(n7628) );
  MUX2_X1 U9999 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9657), .Z(n7680) );
  MUX2_X1 U10000 ( .A(n10582), .B(n10585), .S(n9657), .Z(n7631) );
  INV_X1 U10001 ( .A(SI_19_), .ZN(n10018) );
  INV_X1 U10002 ( .A(n7631), .ZN(n7632) );
  NAND2_X1 U10003 ( .A1(n7632), .A2(SI_19_), .ZN(n7633) );
  NAND2_X1 U10004 ( .A1(n7964), .A2(n7633), .ZN(n7962) );
  NOR2_X1 U10005 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7638) );
  NAND4_X1 U10006 ( .A1(n7638), .A2(n7637), .A3(n7636), .A4(n7635), .ZN(n7731)
         );
  NAND4_X1 U10007 ( .A1(n7641), .A2(n7732), .A3(n7640), .A4(n7639), .ZN(n7642)
         );
  NOR2_X1 U10008 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n7644) );
  NOR2_X1 U10009 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .ZN(n7643) );
  NAND4_X1 U10010 ( .A1(n7652), .A2(n7644), .A3(n7643), .A4(n8136), .ZN(n8205)
         );
  NAND4_X1 U10011 ( .A1(n8212), .A2(n8208), .A3(n8222), .A4(n8215), .ZN(n7645)
         );
  NOR2_X1 U10012 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n7651) );
  NOR2_X1 U10013 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7650) );
  MUX2_X1 U10014 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7654), .S(
        P2_IR_REG_19__SCAN_IN), .Z(n7656) );
  AOI22_X1 U10015 ( .A1(n9338), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7942), 
        .B2(n10418), .ZN(n7657) );
  INV_X1 U10016 ( .A(n7820), .ZN(n7659) );
  INV_X1 U10017 ( .A(n7835), .ZN(n7660) );
  AND2_X1 U10018 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n7661) );
  AND2_X1 U10019 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n7663) );
  INV_X1 U10020 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n7737) );
  INV_X1 U10021 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7719) );
  INV_X1 U10022 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7667) );
  INV_X1 U10023 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7666) );
  OAI21_X1 U10024 ( .B1(n7709), .B2(n7667), .A(n7666), .ZN(n7669) );
  NAND2_X1 U10025 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .ZN(n7668) );
  AND2_X1 U10026 ( .A1(n7669), .A2(n7970), .ZN(n13019) );
  INV_X1 U10027 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7672) );
  INV_X1 U10028 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7674) );
  NAND2_X1 U10029 ( .A1(n13019), .A2(n8122), .ZN(n7679) );
  AOI22_X1 U10030 ( .A1(n9306), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n9305), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n7678) );
  NAND2_X1 U10031 ( .A1(n8056), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7677) );
  INV_X1 U10032 ( .A(n12697), .ZN(n13003) );
  XNOR2_X1 U10033 ( .A(n7681), .B(n7680), .ZN(n11555) );
  NAND2_X1 U10034 ( .A1(n11555), .A2(n7682), .ZN(n7689) );
  OR2_X1 U10035 ( .A1(n7683), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n7684) );
  NAND2_X1 U10036 ( .A1(n7684), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7700) );
  INV_X1 U10037 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7685) );
  NAND2_X1 U10038 ( .A1(n7700), .A2(n7685), .ZN(n7686) );
  NAND2_X1 U10039 ( .A1(n7686), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7687) );
  XNOR2_X1 U10040 ( .A(n7687), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9502) );
  AOI22_X1 U10041 ( .A1(n9338), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7942), 
        .B2(n9502), .ZN(n7688) );
  XNOR2_X1 U10042 ( .A(n7709), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n13033) );
  NAND2_X1 U10043 ( .A1(n13033), .A2(n8122), .ZN(n7696) );
  INV_X1 U10044 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7693) );
  NAND2_X1 U10045 ( .A1(n9306), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7692) );
  INV_X1 U10046 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n7690) );
  OR2_X1 U10047 ( .A1(n6770), .A2(n7690), .ZN(n7691) );
  OAI211_X1 U10048 ( .C1(n7693), .C2(n7786), .A(n7692), .B(n7691), .ZN(n7694)
         );
  INV_X1 U10049 ( .A(n7694), .ZN(n7695) );
  INV_X1 U10050 ( .A(n13014), .ZN(n12728) );
  XNOR2_X1 U10051 ( .A(n7697), .B(SI_17_), .ZN(n7698) );
  XNOR2_X1 U10052 ( .A(n7699), .B(n7698), .ZN(n11520) );
  NAND2_X1 U10053 ( .A1(n11520), .A2(n7682), .ZN(n7702) );
  XNOR2_X1 U10054 ( .A(n7700), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9457) );
  AOI22_X1 U10055 ( .A1(n9338), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7942), 
        .B2(n9457), .ZN(n7701) );
  INV_X1 U10056 ( .A(n9306), .ZN(n8147) );
  INV_X1 U10057 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n7703) );
  OR2_X1 U10058 ( .A1(n8147), .A2(n7703), .ZN(n7706) );
  INV_X1 U10059 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7704) );
  OR2_X1 U10060 ( .A1(n6770), .A2(n7704), .ZN(n7705) );
  AND2_X1 U10061 ( .A1(n7706), .A2(n7705), .ZN(n7712) );
  INV_X1 U10062 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U10063 ( .A1(n7721), .A2(n7707), .ZN(n7708) );
  NAND2_X1 U10064 ( .A1(n7709), .A2(n7708), .ZN(n13042) );
  OR2_X1 U10065 ( .A1(n13042), .A2(n7763), .ZN(n7711) );
  INV_X1 U10066 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9500) );
  OR2_X1 U10067 ( .A1(n7786), .A2(n9500), .ZN(n7710) );
  INV_X1 U10068 ( .A(n13058), .ZN(n12729) );
  XNOR2_X1 U10069 ( .A(n7714), .B(n7713), .ZN(n11511) );
  NAND2_X1 U10070 ( .A1(n11511), .A2(n7682), .ZN(n7717) );
  NAND2_X1 U10071 ( .A1(n7683), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7715) );
  XNOR2_X1 U10072 ( .A(n7715), .B(P2_IR_REG_16__SCAN_IN), .ZN(n9458) );
  AOI22_X1 U10073 ( .A1(n9338), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7942), 
        .B2(n9458), .ZN(n7716) );
  NAND2_X1 U10074 ( .A1(n9306), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7725) );
  INV_X1 U10075 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7718) );
  OR2_X1 U10076 ( .A1(n6770), .A2(n7718), .ZN(n7724) );
  NAND2_X1 U10077 ( .A1(n7739), .A2(n7719), .ZN(n7720) );
  NAND2_X1 U10078 ( .A1(n7721), .A2(n7720), .ZN(n13070) );
  OR2_X1 U10079 ( .A1(n7763), .A2(n13070), .ZN(n7723) );
  INV_X1 U10080 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9499) );
  OR2_X1 U10081 ( .A1(n7786), .A2(n9499), .ZN(n7722) );
  XNOR2_X1 U10082 ( .A(n7728), .B(SI_15_), .ZN(n7729) );
  NAND2_X1 U10083 ( .A1(n11219), .A2(n7682), .ZN(n7735) );
  AND2_X1 U10084 ( .A1(n7730), .A2(n6681), .ZN(n7925) );
  NAND2_X1 U10085 ( .A1(n7925), .A2(n7732), .ZN(n7940) );
  OR2_X1 U10086 ( .A1(n7940), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n7747) );
  OAI21_X1 U10087 ( .B1(n7747), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7733) );
  XNOR2_X1 U10088 ( .A(n7733), .B(P2_IR_REG_15__SCAN_IN), .ZN(n14584) );
  AOI22_X1 U10089 ( .A1(n9338), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7942), 
        .B2(n14584), .ZN(n7734) );
  INV_X1 U10090 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7736) );
  OR2_X1 U10091 ( .A1(n6770), .A2(n7736), .ZN(n7744) );
  NAND2_X1 U10092 ( .A1(n9306), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n7743) );
  NAND2_X1 U10093 ( .A1(n7954), .A2(n7737), .ZN(n7738) );
  NAND2_X1 U10094 ( .A1(n7739), .A2(n7738), .ZN(n12719) );
  OR2_X1 U10095 ( .A1(n7763), .A2(n12719), .ZN(n7742) );
  INV_X1 U10096 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7740) );
  OR2_X1 U10097 ( .A1(n7786), .A2(n7740), .ZN(n7741) );
  NAND4_X1 U10098 ( .A1(n7744), .A2(n7743), .A3(n7742), .A4(n7741), .ZN(n12730) );
  INV_X1 U10099 ( .A(n12730), .ZN(n13056) );
  NAND2_X1 U10100 ( .A1(n11176), .A2(n7682), .ZN(n7750) );
  NAND2_X1 U10101 ( .A1(n7747), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7748) );
  XNOR2_X1 U10102 ( .A(n7748), .B(P2_IR_REG_14__SCAN_IN), .ZN(n9496) );
  AOI22_X1 U10103 ( .A1(n9338), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7942), 
        .B2(n9496), .ZN(n7749) );
  INV_X1 U10104 ( .A(n11406), .ZN(n14180) );
  NAND2_X1 U10105 ( .A1(n7769), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7752) );
  NAND2_X1 U10106 ( .A1(n8056), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7751) );
  INV_X1 U10107 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n12747) );
  INV_X1 U10108 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n13080) );
  INV_X1 U10109 ( .A(n7753), .ZN(n7754) );
  NAND2_X1 U10110 ( .A1(n7755), .A2(n7754), .ZN(n7756) );
  NAND2_X1 U10111 ( .A1(n7757), .A2(n7756), .ZN(n9699) );
  INV_X1 U10112 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n12751) );
  NAND2_X1 U10113 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n7758) );
  MUX2_X1 U10114 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7758), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n7759) );
  INV_X1 U10115 ( .A(n7649), .ZN(n7779) );
  NAND2_X1 U10116 ( .A1(n7759), .A2(n7779), .ZN(n12749) );
  INV_X1 U10117 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7761) );
  INV_X1 U10118 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U10119 ( .A1(n7769), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7765) );
  NAND2_X1 U10120 ( .A1(n9657), .A2(SI_0_), .ZN(n7768) );
  XNOR2_X1 U10121 ( .A(n7768), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13204) );
  MUX2_X2 U10122 ( .A(P2_IR_REG_0__SCAN_IN), .B(n13204), .S(n9454), .Z(n10515)
         );
  INV_X1 U10123 ( .A(n10515), .ZN(n9957) );
  NOR2_X1 U10124 ( .A1(n12746), .A2(n9957), .ZN(n9887) );
  INV_X1 U10125 ( .A(n12745), .ZN(n8154) );
  NAND2_X1 U10126 ( .A1(n8154), .A2(n10021), .ZN(n10654) );
  INV_X1 U10127 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n12760) );
  INV_X1 U10128 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U10129 ( .A1(n7775), .A2(n7774), .ZN(n7777) );
  NAND2_X1 U10130 ( .A1(n7777), .A2(n7776), .ZN(n9992) );
  NAND2_X1 U10131 ( .A1(n7778), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7784) );
  NAND2_X1 U10132 ( .A1(n7779), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7780) );
  MUX2_X1 U10133 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7780), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n7782) );
  NAND2_X1 U10134 ( .A1(n7782), .A2(n7781), .ZN(n12761) );
  INV_X1 U10135 ( .A(n12761), .ZN(n9465) );
  NAND2_X1 U10136 ( .A1(n7942), .A2(n9465), .ZN(n7783) );
  INV_X2 U10137 ( .A(n12684), .ZN(n14645) );
  NAND2_X1 U10138 ( .A1(n10375), .A2(n10376), .ZN(n7799) );
  NAND2_X1 U10139 ( .A1(n7769), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7790) );
  OR2_X1 U10140 ( .A1(n7763), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7789) );
  INV_X1 U10141 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9466) );
  OR2_X1 U10142 ( .A1(n7786), .A2(n9466), .ZN(n7788) );
  INV_X1 U10143 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10380) );
  OR2_X1 U10144 ( .A1(n7762), .A2(n10380), .ZN(n7787) );
  NAND2_X1 U10145 ( .A1(n7781), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7791) );
  XNOR2_X1 U10146 ( .A(n7791), .B(P2_IR_REG_3__SCAN_IN), .ZN(n9806) );
  AOI22_X1 U10147 ( .A1(n7778), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n7942), .B2(
        n9806), .ZN(n7797) );
  OR2_X1 U10148 ( .A1(n7793), .A2(n7792), .ZN(n7794) );
  AND2_X1 U10149 ( .A1(n7795), .A2(n7794), .ZN(n10108) );
  INV_X1 U10150 ( .A(n10377), .ZN(n7798) );
  NAND2_X1 U10151 ( .A1(n7799), .A2(n7798), .ZN(n10374) );
  NAND2_X1 U10152 ( .A1(n10420), .A2(n14651), .ZN(n10421) );
  NAND2_X1 U10153 ( .A1(n10374), .A2(n10421), .ZN(n7812) );
  NAND2_X1 U10154 ( .A1(n9306), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7803) );
  INV_X1 U10155 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10428) );
  OR2_X1 U10156 ( .A1(n6770), .A2(n10428), .ZN(n7802) );
  OAI21_X1 U10157 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n7820), .ZN(n10430) );
  OR2_X1 U10158 ( .A1(n7763), .A2(n10430), .ZN(n7801) );
  INV_X1 U10159 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9469) );
  OR2_X1 U10160 ( .A1(n7786), .A2(n9469), .ZN(n7800) );
  AND4_X2 U10161 ( .A1(n7803), .A2(n7802), .A3(n7801), .A4(n7800), .ZN(n10090)
         );
  OR2_X1 U10162 ( .A1(n7805), .A2(n7804), .ZN(n7806) );
  AND2_X1 U10163 ( .A1(n7807), .A2(n7806), .ZN(n10224) );
  NAND2_X1 U10164 ( .A1(n7808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7809) );
  XNOR2_X1 U10165 ( .A(n7809), .B(P2_IR_REG_4__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U10166 ( .A1(n7778), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7942), .B2(
        n12777), .ZN(n7810) );
  INV_X1 U10167 ( .A(n10422), .ZN(n7811) );
  NAND2_X1 U10168 ( .A1(n14659), .A2(n10090), .ZN(n7813) );
  XNOR2_X1 U10169 ( .A(n7815), .B(n7814), .ZN(n10253) );
  NAND2_X1 U10170 ( .A1(n10253), .A2(n7682), .ZN(n7818) );
  INV_X1 U10171 ( .A(n7730), .ZN(n7831) );
  NAND2_X1 U10172 ( .A1(n7831), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7816) );
  XNOR2_X1 U10173 ( .A(n7816), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9850) );
  AOI22_X1 U10174 ( .A1(n9338), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7942), .B2(
        n9850), .ZN(n7817) );
  NAND2_X1 U10175 ( .A1(n7818), .A2(n7817), .ZN(n10471) );
  NAND2_X1 U10176 ( .A1(n9305), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7825) );
  NAND2_X1 U10177 ( .A1(n9306), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7824) );
  INV_X1 U10178 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U10179 ( .A1(n7820), .A2(n7819), .ZN(n7821) );
  NAND2_X1 U10180 ( .A1(n7835), .A2(n7821), .ZN(n10472) );
  OR2_X1 U10181 ( .A1(n7763), .A2(n10472), .ZN(n7823) );
  INV_X1 U10182 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n9472) );
  OR2_X1 U10183 ( .A1(n7786), .A2(n9472), .ZN(n7822) );
  OR2_X1 U10184 ( .A1(n10471), .A2(n10438), .ZN(n7826) );
  NAND2_X1 U10185 ( .A1(n7830), .A2(n7829), .ZN(n10257) );
  OR2_X1 U10186 ( .A1(n10257), .A2(n9337), .ZN(n7833) );
  NAND2_X1 U10187 ( .A1(n7864), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7848) );
  XNOR2_X1 U10188 ( .A(n7848), .B(P2_IR_REG_6__SCAN_IN), .ZN(n12793) );
  AOI22_X1 U10189 ( .A1(n9338), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7942), .B2(
        n12793), .ZN(n7832) );
  NAND2_X1 U10190 ( .A1(n9306), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7840) );
  INV_X1 U10191 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10443) );
  OR2_X1 U10192 ( .A1(n6770), .A2(n10443), .ZN(n7839) );
  INV_X1 U10193 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U10194 ( .A1(n7835), .A2(n7834), .ZN(n7836) );
  NAND2_X1 U10195 ( .A1(n7853), .A2(n7836), .ZN(n10445) );
  OR2_X1 U10196 ( .A1(n7763), .A2(n10445), .ZN(n7838) );
  OR2_X1 U10197 ( .A1(n7786), .A2(n14729), .ZN(n7837) );
  INV_X1 U10198 ( .A(n10453), .ZN(n12740) );
  NAND2_X1 U10199 ( .A1(n7841), .A2(n10453), .ZN(n7842) );
  INV_X1 U10200 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7847) );
  NAND2_X1 U10201 ( .A1(n7848), .A2(n7847), .ZN(n7849) );
  NAND2_X1 U10202 ( .A1(n7849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7850) );
  XNOR2_X1 U10203 ( .A(n7850), .B(P2_IR_REG_7__SCAN_IN), .ZN(n12808) );
  AOI22_X1 U10204 ( .A1(n9338), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7942), .B2(
        n12808), .ZN(n7851) );
  NAND2_X1 U10205 ( .A1(n9306), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7858) );
  INV_X1 U10206 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10455) );
  OR2_X1 U10207 ( .A1(n6770), .A2(n10455), .ZN(n7857) );
  NAND2_X1 U10208 ( .A1(n7853), .A2(n10525), .ZN(n7854) );
  NAND2_X1 U10209 ( .A1(n7873), .A2(n7854), .ZN(n10528) );
  OR2_X1 U10210 ( .A1(n7763), .A2(n10528), .ZN(n7856) );
  INV_X1 U10211 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9477) );
  OR2_X1 U10212 ( .A1(n7786), .A2(n9477), .ZN(n7855) );
  NOR2_X1 U10213 ( .A1(n14684), .A2(n12739), .ZN(n7860) );
  NAND2_X1 U10214 ( .A1(n14684), .A2(n12739), .ZN(n7859) );
  INV_X1 U10215 ( .A(n7864), .ZN(n7866) );
  NOR2_X1 U10216 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n7865) );
  NAND2_X1 U10217 ( .A1(n7866), .A2(n7865), .ZN(n7868) );
  NAND2_X1 U10218 ( .A1(n7868), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7867) );
  MUX2_X1 U10219 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7867), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n7869) );
  AOI22_X1 U10220 ( .A1(n9338), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7942), .B2(
        n12824), .ZN(n7870) );
  NAND2_X1 U10221 ( .A1(n9305), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7878) );
  INV_X1 U10222 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n7871) );
  OR2_X1 U10223 ( .A1(n8147), .A2(n7871), .ZN(n7877) );
  NAND2_X1 U10224 ( .A1(n7873), .A2(n7872), .ZN(n7874) );
  NAND2_X1 U10225 ( .A1(n7889), .A2(n7874), .ZN(n10728) );
  OR2_X1 U10226 ( .A1(n7763), .A2(n10728), .ZN(n7876) );
  INV_X1 U10227 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9480) );
  OR2_X1 U10228 ( .A1(n7786), .A2(n9480), .ZN(n7875) );
  INV_X1 U10229 ( .A(n10741), .ZN(n12738) );
  AND2_X1 U10230 ( .A1(n14692), .A2(n12738), .ZN(n7880) );
  OR2_X1 U10231 ( .A1(n14692), .A2(n12738), .ZN(n7879) );
  XNOR2_X1 U10232 ( .A(n7882), .B(n7881), .ZN(n10541) );
  NAND2_X1 U10233 ( .A1(n10541), .A2(n7682), .ZN(n7887) );
  NAND2_X1 U10234 ( .A1(n7884), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7883) );
  MUX2_X1 U10235 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7883), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n7885) );
  AOI22_X1 U10236 ( .A1(n9338), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7942), .B2(
        n9484), .ZN(n7886) );
  NAND2_X1 U10237 ( .A1(n9305), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7894) );
  NAND2_X1 U10238 ( .A1(n9306), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7893) );
  NAND2_X1 U10239 ( .A1(n7889), .A2(n7888), .ZN(n7890) );
  NAND2_X1 U10240 ( .A1(n7915), .A2(n7890), .ZN(n10797) );
  OR2_X1 U10241 ( .A1(n7763), .A2(n10797), .ZN(n7892) );
  INV_X1 U10242 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9518) );
  OR2_X1 U10243 ( .A1(n7786), .A2(n9518), .ZN(n7891) );
  NAND4_X1 U10244 ( .A1(n7894), .A2(n7893), .A3(n7892), .A4(n7891), .ZN(n12736) );
  XNOR2_X1 U10245 ( .A(n10793), .B(n10787), .ZN(n10744) );
  OR2_X1 U10246 ( .A1(n10793), .A2(n10787), .ZN(n7896) );
  OR2_X1 U10247 ( .A1(n7898), .A2(n7897), .ZN(n7899) );
  NAND2_X1 U10248 ( .A1(n7900), .A2(n7899), .ZN(n10546) );
  OR2_X1 U10249 ( .A1(n10546), .A2(n9337), .ZN(n7903) );
  NAND2_X1 U10250 ( .A1(n7910), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7901) );
  XNOR2_X1 U10251 ( .A(n7901), .B(P2_IR_REG_10__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U10252 ( .A1(n9338), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7942), 
        .B2(n12840), .ZN(n7902) );
  NAND2_X1 U10253 ( .A1(n9305), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7907) );
  NAND2_X1 U10254 ( .A1(n9306), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7906) );
  INV_X1 U10255 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7914) );
  XNOR2_X1 U10256 ( .A(n7915), .B(n7914), .ZN(n10937) );
  OR2_X1 U10257 ( .A1(n7763), .A2(n10937), .ZN(n7905) );
  INV_X1 U10258 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9487) );
  OR2_X1 U10259 ( .A1(n7786), .A2(n9487), .ZN(n7904) );
  NAND4_X1 U10260 ( .A1(n7907), .A2(n7906), .A3(n7905), .A4(n7904), .ZN(n12735) );
  INV_X1 U10261 ( .A(n12735), .ZN(n10773) );
  XNOR2_X1 U10262 ( .A(n10933), .B(n10773), .ZN(n10676) );
  INV_X1 U10263 ( .A(n10676), .ZN(n10671) );
  OAI21_X1 U10264 ( .B1(n7910), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7911) );
  XNOR2_X1 U10265 ( .A(n7911), .B(P2_IR_REG_11__SCAN_IN), .ZN(n9905) );
  AOI22_X1 U10266 ( .A1(n9338), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n9905), 
        .B2(n7942), .ZN(n7912) );
  NAND2_X1 U10267 ( .A1(n9306), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7920) );
  INV_X1 U10268 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10781) );
  OR2_X1 U10269 ( .A1(n6770), .A2(n10781), .ZN(n7919) );
  INV_X1 U10270 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7913) );
  OAI21_X1 U10271 ( .B1(n7915), .B2(n7914), .A(n7913), .ZN(n7916) );
  NAND2_X1 U10272 ( .A1(n7916), .A2(n7930), .ZN(n11089) );
  OR2_X1 U10273 ( .A1(n7763), .A2(n11089), .ZN(n7918) );
  INV_X1 U10274 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9488) );
  OR2_X1 U10275 ( .A1(n7786), .A2(n9488), .ZN(n7917) );
  NAND2_X1 U10276 ( .A1(n11091), .A2(n12734), .ZN(n8169) );
  OR2_X1 U10277 ( .A1(n11091), .A2(n12734), .ZN(n7921) );
  NOR2_X1 U10278 ( .A1(n10933), .A2(n10773), .ZN(n10769) );
  OR2_X1 U10279 ( .A1(n14716), .A2(n12734), .ZN(n7922) );
  XNOR2_X1 U10280 ( .A(n7924), .B(n7923), .ZN(n11018) );
  NAND2_X1 U10281 ( .A1(n11018), .A2(n7682), .ZN(n7929) );
  INV_X1 U10282 ( .A(n7925), .ZN(n7926) );
  NAND2_X1 U10283 ( .A1(n7926), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7927) );
  XNOR2_X1 U10284 ( .A(n7927), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9922) );
  AOI22_X1 U10285 ( .A1(n9338), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7942), 
        .B2(n9922), .ZN(n7928) );
  AND2_X2 U10286 ( .A1(n7929), .A2(n7928), .ZN(n14186) );
  NAND2_X1 U10287 ( .A1(n9306), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7935) );
  INV_X1 U10288 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10969) );
  OR2_X1 U10289 ( .A1(n6770), .A2(n10969), .ZN(n7934) );
  NAND2_X1 U10290 ( .A1(n7930), .A2(n9971), .ZN(n7931) );
  NAND2_X1 U10291 ( .A1(n7952), .A2(n7931), .ZN(n11287) );
  OR2_X1 U10292 ( .A1(n7763), .A2(n11287), .ZN(n7933) );
  INV_X1 U10293 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9492) );
  OR2_X1 U10294 ( .A1(n7786), .A2(n9492), .ZN(n7932) );
  INV_X1 U10295 ( .A(n11317), .ZN(n12733) );
  NOR2_X1 U10296 ( .A1(n14186), .A2(n12733), .ZN(n7936) );
  NAND2_X1 U10297 ( .A1(n14186), .A2(n12733), .ZN(n7937) );
  XNOR2_X1 U10298 ( .A(n7939), .B(n7938), .ZN(n11024) );
  NAND2_X1 U10299 ( .A1(n11024), .A2(n7682), .ZN(n7944) );
  NAND2_X1 U10300 ( .A1(n7940), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7941) );
  XNOR2_X1 U10301 ( .A(n7941), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10011) );
  AOI22_X1 U10302 ( .A1(n9338), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7942), 
        .B2(n10011), .ZN(n7943) );
  NAND2_X1 U10303 ( .A1(n9306), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7949) );
  INV_X1 U10304 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10063) );
  XNOR2_X1 U10305 ( .A(n7952), .B(n10063), .ZN(n11316) );
  OR2_X1 U10306 ( .A1(n7763), .A2(n11316), .ZN(n7948) );
  INV_X1 U10307 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7945) );
  OR2_X1 U10308 ( .A1(n7786), .A2(n7945), .ZN(n7947) );
  INV_X1 U10309 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n11120) );
  OR2_X1 U10310 ( .A1(n6770), .A2(n11120), .ZN(n7946) );
  XNOR2_X1 U10311 ( .A(n11324), .B(n11418), .ZN(n11113) );
  INV_X1 U10312 ( .A(n11113), .ZN(n11115) );
  INV_X1 U10313 ( .A(n11418), .ZN(n12732) );
  AND2_X1 U10314 ( .A1(n11314), .A2(n12732), .ZN(n7950) );
  NAND2_X1 U10315 ( .A1(n9305), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7959) );
  NAND2_X1 U10316 ( .A1(n9306), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n7958) );
  INV_X1 U10317 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7951) );
  OAI21_X1 U10318 ( .B1(n7952), .B2(n10063), .A(n7951), .ZN(n7953) );
  NAND2_X1 U10319 ( .A1(n7954), .A2(n7953), .ZN(n11417) );
  OR2_X1 U10320 ( .A1(n7763), .A2(n11417), .ZN(n7957) );
  INV_X1 U10321 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7955) );
  OR2_X1 U10322 ( .A1(n7786), .A2(n7955), .ZN(n7956) );
  NAND4_X1 U10323 ( .A1(n7959), .A2(n7958), .A3(n7957), .A4(n7956), .ZN(n12731) );
  INV_X1 U10324 ( .A(n12731), .ZN(n11315) );
  INV_X1 U10325 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10943) );
  MUX2_X1 U10326 ( .A(n11007), .B(n10943), .S(n9657), .Z(n7994) );
  NAND2_X1 U10327 ( .A1(n11579), .A2(n7682), .ZN(n7967) );
  NAND2_X1 U10328 ( .A1(n9338), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7966) );
  INV_X1 U10329 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n7974) );
  INV_X1 U10330 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7969) );
  NAND2_X1 U10331 ( .A1(n7970), .A2(n7969), .ZN(n7971) );
  NAND2_X1 U10332 ( .A1(n7984), .A2(n7971), .ZN(n12997) );
  OR2_X1 U10333 ( .A1(n12997), .A2(n7763), .ZN(n7973) );
  AOI22_X1 U10334 ( .A1(n9306), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n9305), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n7972) );
  OAI211_X1 U10335 ( .C1(n7786), .C2(n7974), .A(n7973), .B(n7972), .ZN(n12976)
         );
  INV_X1 U10336 ( .A(n12976), .ZN(n13015) );
  NAND2_X1 U10337 ( .A1(n13142), .A2(n13015), .ZN(n7976) );
  OR2_X1 U10338 ( .A1(n13142), .A2(n13015), .ZN(n7975) );
  NAND2_X1 U10339 ( .A1(n7976), .A2(n7975), .ZN(n12991) );
  INV_X1 U10340 ( .A(n12991), .ZN(n13001) );
  NAND2_X1 U10341 ( .A1(n12999), .A2(n7976), .ZN(n12974) );
  NAND2_X1 U10342 ( .A1(n7977), .A2(n7992), .ZN(n7979) );
  INV_X1 U10343 ( .A(SI_20_), .ZN(n10167) );
  OR2_X1 U10344 ( .A1(n7993), .A2(n10167), .ZN(n7978) );
  MUX2_X1 U10345 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9657), .Z(n7995) );
  XNOR2_X1 U10346 ( .A(n7995), .B(SI_21_), .ZN(n7980) );
  NAND2_X1 U10347 ( .A1(n11597), .A2(n7682), .ZN(n7983) );
  NAND2_X1 U10348 ( .A1(n9338), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n7982) );
  INV_X1 U10349 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12620) );
  NAND2_X1 U10350 ( .A1(n7984), .A2(n12620), .ZN(n7985) );
  NAND2_X1 U10351 ( .A1(n8001), .A2(n7985), .ZN(n12980) );
  OR2_X1 U10352 ( .A1(n12980), .A2(n7763), .ZN(n7991) );
  INV_X1 U10353 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U10354 ( .A1(n9305), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n7987) );
  NAND2_X1 U10355 ( .A1(n9306), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7986) );
  OAI211_X1 U10356 ( .C1(n7988), .C2(n7786), .A(n7987), .B(n7986), .ZN(n7989)
         );
  INV_X1 U10357 ( .A(n7989), .ZN(n7990) );
  NAND2_X1 U10358 ( .A1(n7991), .A2(n7990), .ZN(n13005) );
  INV_X1 U10359 ( .A(n13134), .ZN(n9279) );
  NOR2_X1 U10360 ( .A1(n7994), .A2(n10167), .ZN(n7996) );
  AOI22_X1 U10361 ( .A1(n7996), .A2(n6477), .B1(n7995), .B2(SI_21_), .ZN(n7997) );
  MUX2_X1 U10362 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9657), .Z(n8028) );
  XNOR2_X1 U10363 ( .A(n11610), .B(n8028), .ZN(n11149) );
  NAND2_X1 U10364 ( .A1(n11149), .A2(n7682), .ZN(n7999) );
  NAND2_X1 U10365 ( .A1(n9338), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n7998) );
  INV_X1 U10366 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10367 ( .A1(n8001), .A2(n8000), .ZN(n8002) );
  AND2_X1 U10368 ( .A1(n8015), .A2(n8002), .ZN(n12968) );
  INV_X1 U10369 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n15052) );
  NAND2_X1 U10370 ( .A1(n9305), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8004) );
  NAND2_X1 U10371 ( .A1(n9306), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8003) );
  OAI211_X1 U10372 ( .C1(n15052), .C2(n7786), .A(n8004), .B(n8003), .ZN(n8005)
         );
  AOI21_X1 U10373 ( .B1(n12968), .B2(n8122), .A(n8005), .ZN(n12621) );
  INV_X1 U10374 ( .A(n12621), .ZN(n12975) );
  XNOR2_X1 U10375 ( .A(n12679), .B(n12975), .ZN(n9374) );
  INV_X1 U10376 ( .A(n11610), .ZN(n8006) );
  NAND2_X1 U10377 ( .A1(n8006), .A2(n8028), .ZN(n8008) );
  NAND2_X1 U10378 ( .A1(n8027), .A2(SI_22_), .ZN(n8007) );
  MUX2_X1 U10379 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9657), .Z(n8030) );
  XNOR2_X1 U10380 ( .A(n8030), .B(SI_23_), .ZN(n8009) );
  NAND2_X1 U10381 ( .A1(n11627), .A2(n7682), .ZN(n8012) );
  NAND2_X1 U10382 ( .A1(n9338), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8011) );
  INV_X1 U10383 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10384 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  NAND2_X1 U10385 ( .A1(n8038), .A2(n8016), .ZN(n12950) );
  OR2_X1 U10386 ( .A1(n12950), .A2(n7763), .ZN(n8022) );
  INV_X1 U10387 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8019) );
  NAND2_X1 U10388 ( .A1(n9305), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8018) );
  NAND2_X1 U10389 ( .A1(n9306), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8017) );
  OAI211_X1 U10390 ( .C1(n8019), .C2(n7786), .A(n8018), .B(n8017), .ZN(n8020)
         );
  INV_X1 U10391 ( .A(n8020), .ZN(n8021) );
  NAND2_X1 U10392 ( .A1(n12954), .A2(n12931), .ZN(n8023) );
  INV_X1 U10393 ( .A(n8030), .ZN(n8024) );
  INV_X1 U10394 ( .A(SI_23_), .ZN(n10513) );
  NAND2_X1 U10395 ( .A1(n8024), .A2(n10513), .ZN(n8031) );
  OAI21_X1 U10396 ( .B1(SI_22_), .B2(n8028), .A(n8031), .ZN(n8025) );
  INV_X1 U10397 ( .A(n8025), .ZN(n8026) );
  INV_X1 U10398 ( .A(n8028), .ZN(n8029) );
  INV_X1 U10399 ( .A(SI_22_), .ZN(n8695) );
  NOR2_X1 U10400 ( .A1(n8029), .A2(n8695), .ZN(n8032) );
  AOI22_X1 U10401 ( .A1(n8032), .A2(n8031), .B1(n8030), .B2(SI_23_), .ZN(n8033) );
  MUX2_X1 U10402 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9657), .Z(n8047) );
  NAND2_X1 U10403 ( .A1(n11640), .A2(n7682), .ZN(n8036) );
  NAND2_X1 U10404 ( .A1(n9338), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8035) );
  INV_X1 U10405 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n15051) );
  NAND2_X1 U10406 ( .A1(n8038), .A2(n15051), .ZN(n8039) );
  NAND2_X1 U10407 ( .A1(n8070), .A2(n8039), .ZN(n12936) );
  INV_X1 U10408 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8042) );
  NAND2_X1 U10409 ( .A1(n9305), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8041) );
  NAND2_X1 U10410 ( .A1(n9306), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8040) );
  OAI211_X1 U10411 ( .C1(n8042), .C2(n7786), .A(n8041), .B(n8040), .ZN(n8043)
         );
  INV_X1 U10412 ( .A(n8043), .ZN(n8044) );
  INV_X1 U10413 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8289) );
  INV_X1 U10414 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11297) );
  MUX2_X1 U10415 ( .A(n8289), .B(n11297), .S(n9657), .Z(n8051) );
  INV_X1 U10416 ( .A(SI_25_), .ZN(n11015) );
  NAND2_X1 U10417 ( .A1(n8051), .A2(n11015), .ZN(n8064) );
  INV_X1 U10418 ( .A(n8051), .ZN(n8052) );
  NAND2_X1 U10419 ( .A1(n8052), .A2(SI_25_), .ZN(n8053) );
  NAND2_X1 U10420 ( .A1(n8064), .A2(n8053), .ZN(n8062) );
  NAND2_X1 U10421 ( .A1(n11661), .A2(n7682), .ZN(n8055) );
  NAND2_X1 U10422 ( .A1(n9338), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8054) );
  XNOR2_X1 U10423 ( .A(n8070), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n12921) );
  NAND2_X1 U10424 ( .A1(n12921), .A2(n8122), .ZN(n8061) );
  INV_X1 U10425 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n15124) );
  NAND2_X1 U10426 ( .A1(n9305), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8058) );
  NAND2_X1 U10427 ( .A1(n8056), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8057) );
  OAI211_X1 U10428 ( .C1(n8147), .C2(n15124), .A(n8058), .B(n8057), .ZN(n8059)
         );
  INV_X1 U10429 ( .A(n8059), .ZN(n8060) );
  INV_X1 U10430 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n13991) );
  INV_X1 U10431 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13202) );
  MUX2_X1 U10432 ( .A(n13991), .B(n13202), .S(n9657), .Z(n8079) );
  XNOR2_X1 U10433 ( .A(n8079), .B(SI_26_), .ZN(n8065) );
  NAND2_X1 U10434 ( .A1(n13200), .A2(n7682), .ZN(n8067) );
  NAND2_X1 U10435 ( .A1(n9338), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8066) );
  INV_X1 U10436 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12628) );
  INV_X1 U10437 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8068) );
  OAI21_X1 U10438 ( .B1(n8070), .B2(n12628), .A(n8068), .ZN(n8071) );
  NAND2_X1 U10439 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .ZN(n8069) );
  NAND2_X1 U10440 ( .A1(n12907), .A2(n8122), .ZN(n8077) );
  INV_X1 U10441 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10442 ( .A1(n9305), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8073) );
  NAND2_X1 U10443 ( .A1(n9306), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8072) );
  OAI211_X1 U10444 ( .C1(n8074), .C2(n7786), .A(n8073), .B(n8072), .ZN(n8075)
         );
  INV_X1 U10445 ( .A(n8075), .ZN(n8076) );
  INV_X1 U10446 ( .A(n9361), .ZN(n8078) );
  NAND2_X1 U10447 ( .A1(n13108), .A2(n12629), .ZN(n9360) );
  INV_X1 U10448 ( .A(SI_26_), .ZN(n11200) );
  MUX2_X1 U10449 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9657), .Z(n8097) );
  INV_X1 U10450 ( .A(n8097), .ZN(n8083) );
  XNOR2_X1 U10451 ( .A(n8083), .B(SI_27_), .ZN(n8084) );
  NAND2_X1 U10452 ( .A1(n9338), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8085) );
  INV_X1 U10453 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12577) );
  INV_X1 U10454 ( .A(n8104), .ZN(n8106) );
  NAND2_X1 U10455 ( .A1(n8087), .A2(n12577), .ZN(n8088) );
  NAND2_X1 U10456 ( .A1(n8106), .A2(n8088), .ZN(n12893) );
  OR2_X1 U10457 ( .A1(n12893), .A2(n7763), .ZN(n8094) );
  INV_X1 U10458 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8091) );
  NAND2_X1 U10459 ( .A1(n9306), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8090) );
  NAND2_X1 U10460 ( .A1(n9305), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8089) );
  OAI211_X1 U10461 ( .C1(n8091), .C2(n7786), .A(n8090), .B(n8089), .ZN(n8092)
         );
  INV_X1 U10462 ( .A(n8092), .ZN(n8093) );
  NOR2_X1 U10463 ( .A1(n8097), .A2(SI_27_), .ZN(n8095) );
  NAND2_X1 U10464 ( .A1(n8097), .A2(SI_27_), .ZN(n8098) );
  INV_X1 U10465 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13987) );
  INV_X1 U10466 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8762) );
  MUX2_X1 U10467 ( .A(n13987), .B(n8762), .S(n9657), .Z(n8099) );
  INV_X1 U10468 ( .A(SI_28_), .ZN(n12529) );
  NAND2_X1 U10469 ( .A1(n8099), .A2(n12529), .ZN(n8119) );
  INV_X1 U10470 ( .A(n8099), .ZN(n8100) );
  NAND2_X1 U10471 ( .A1(n8100), .A2(SI_28_), .ZN(n8101) );
  NAND2_X1 U10472 ( .A1(n8119), .A2(n8101), .ZN(n8117) );
  NAND2_X1 U10473 ( .A1(n13192), .A2(n7682), .ZN(n8103) );
  NAND2_X1 U10474 ( .A1(n9338), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8102) );
  INV_X1 U10475 ( .A(n12859), .ZN(n8108) );
  INV_X1 U10476 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8105) );
  NAND2_X1 U10477 ( .A1(n8106), .A2(n8105), .ZN(n8107) );
  NAND2_X1 U10478 ( .A1(n12875), .A2(n8122), .ZN(n8114) );
  INV_X1 U10479 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8111) );
  NAND2_X1 U10480 ( .A1(n9305), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8110) );
  NAND2_X1 U10481 ( .A1(n9306), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8109) );
  OAI211_X1 U10482 ( .C1(n8111), .C2(n7786), .A(n8110), .B(n8109), .ZN(n8112)
         );
  INV_X1 U10483 ( .A(n8112), .ZN(n8113) );
  NAND2_X1 U10484 ( .A1(n13096), .A2(n12602), .ZN(n8115) );
  INV_X1 U10485 ( .A(n12879), .ZN(n12867) );
  INV_X1 U10486 ( .A(n12727), .ZN(n12870) );
  NAND2_X1 U10487 ( .A1(n13103), .A2(n12870), .ZN(n12868) );
  INV_X1 U10488 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13982) );
  INV_X1 U10489 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11428) );
  MUX2_X1 U10490 ( .A(n13982), .B(n11428), .S(n9657), .Z(n9295) );
  XNOR2_X1 U10491 ( .A(n9295), .B(SI_29_), .ZN(n9293) );
  NAND2_X1 U10492 ( .A1(n11716), .A2(n7682), .ZN(n8121) );
  NAND2_X1 U10493 ( .A1(n9338), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U10494 ( .A1(n12859), .A2(n8122), .ZN(n8128) );
  INV_X1 U10495 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8125) );
  NAND2_X1 U10496 ( .A1(n9306), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8124) );
  NAND2_X1 U10497 ( .A1(n9305), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8123) );
  OAI211_X1 U10498 ( .C1(n8125), .C2(n7786), .A(n8124), .B(n8123), .ZN(n8126)
         );
  INV_X1 U10499 ( .A(n8126), .ZN(n8127) );
  NAND2_X1 U10500 ( .A1(n8128), .A2(n8127), .ZN(n12869) );
  INV_X1 U10501 ( .A(n9377), .ZN(n8129) );
  INV_X1 U10502 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8130) );
  NAND2_X1 U10503 ( .A1(n8132), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8133) );
  INV_X1 U10504 ( .A(n10942), .ZN(n10519) );
  NAND2_X1 U10505 ( .A1(n8193), .A2(n10519), .ZN(n8142) );
  INV_X1 U10506 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8139) );
  NAND2_X1 U10507 ( .A1(n9952), .A2(n10418), .ZN(n8141) );
  INV_X1 U10508 ( .A(n8143), .ZN(n8144) );
  INV_X1 U10509 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8145) );
  OR2_X1 U10510 ( .A1(n7786), .A2(n8145), .ZN(n8150) );
  INV_X1 U10511 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n12853) );
  OR2_X1 U10512 ( .A1(n6770), .A2(n12853), .ZN(n8149) );
  INV_X1 U10513 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8146) );
  OR2_X1 U10514 ( .A1(n8147), .A2(n8146), .ZN(n8148) );
  AND3_X1 U10515 ( .A1(n8150), .A2(n8149), .A3(n8148), .ZN(n9341) );
  INV_X1 U10516 ( .A(P2_B_REG_SCAN_IN), .ZN(n8211) );
  OAI21_X1 U10517 ( .B1(n9393), .B2(n8211), .A(n13004), .ZN(n12845) );
  OAI22_X1 U10518 ( .A1(n12602), .A2(n13055), .B1(n9341), .B2(n12845), .ZN(
        n8151) );
  INV_X1 U10519 ( .A(n9886), .ZN(n8152) );
  NAND2_X1 U10520 ( .A1(n12746), .A2(n10515), .ZN(n9883) );
  NAND2_X1 U10521 ( .A1(n8152), .A2(n9883), .ZN(n9885) );
  INV_X1 U10522 ( .A(n10021), .ZN(n8153) );
  NAND2_X1 U10523 ( .A1(n8154), .A2(n8153), .ZN(n8155) );
  NAND2_X1 U10524 ( .A1(n9885), .A2(n8155), .ZN(n10662) );
  INV_X1 U10525 ( .A(n9365), .ZN(n10661) );
  NAND2_X1 U10526 ( .A1(n10662), .A2(n10661), .ZN(n10660) );
  NAND2_X1 U10527 ( .A1(n10037), .A2(n14645), .ZN(n8156) );
  NAND2_X1 U10528 ( .A1(n10660), .A2(n8156), .ZN(n10365) );
  NAND2_X1 U10529 ( .A1(n10365), .A2(n10377), .ZN(n10364) );
  NAND2_X1 U10530 ( .A1(n10420), .A2(n10383), .ZN(n8157) );
  NAND2_X1 U10531 ( .A1(n10364), .A2(n8157), .ZN(n10417) );
  NAND2_X1 U10532 ( .A1(n10431), .A2(n10090), .ZN(n8158) );
  NAND2_X1 U10533 ( .A1(n10471), .A2(n12741), .ZN(n8159) );
  INV_X1 U10534 ( .A(n10437), .ZN(n8160) );
  NAND2_X1 U10535 ( .A1(n10435), .A2(n8160), .ZN(n8162) );
  NAND2_X1 U10536 ( .A1(n14676), .A2(n10453), .ZN(n8161) );
  NAND2_X1 U10537 ( .A1(n8162), .A2(n8161), .ZN(n10450) );
  INV_X1 U10538 ( .A(n14684), .ZN(n10537) );
  XNOR2_X1 U10539 ( .A(n10537), .B(n12739), .ZN(n10451) );
  INV_X1 U10540 ( .A(n10451), .ZN(n8163) );
  NAND2_X1 U10541 ( .A1(n10450), .A2(n8163), .ZN(n8165) );
  NAND2_X1 U10542 ( .A1(n14684), .A2(n10591), .ZN(n8164) );
  XNOR2_X1 U10543 ( .A(n10731), .B(n10741), .ZN(n10718) );
  INV_X1 U10544 ( .A(n10718), .ZN(n10723) );
  OR2_X1 U10545 ( .A1(n14692), .A2(n10741), .ZN(n8166) );
  NAND2_X1 U10546 ( .A1(n10793), .A2(n12736), .ZN(n8167) );
  NAND2_X1 U10547 ( .A1(n10747), .A2(n8167), .ZN(n10677) );
  NAND2_X1 U10548 ( .A1(n10677), .A2(n10676), .ZN(n10679) );
  NAND2_X1 U10549 ( .A1(n10933), .A2(n12735), .ZN(n8168) );
  NAND2_X1 U10550 ( .A1(n10679), .A2(n8168), .ZN(n10777) );
  NAND2_X1 U10551 ( .A1(n10777), .A2(n10776), .ZN(n10775) );
  NAND2_X1 U10552 ( .A1(n10775), .A2(n8169), .ZN(n10963) );
  NAND2_X1 U10553 ( .A1(n14186), .A2(n11317), .ZN(n8170) );
  NAND2_X1 U10554 ( .A1(n10963), .A2(n8170), .ZN(n8172) );
  OR2_X1 U10555 ( .A1(n14186), .A2(n11317), .ZN(n8171) );
  NOR2_X1 U10556 ( .A1(n11314), .A2(n11418), .ZN(n8173) );
  NAND2_X1 U10557 ( .A1(n11314), .A2(n11418), .ZN(n8174) );
  NOR2_X1 U10558 ( .A1(n11406), .A2(n12731), .ZN(n8175) );
  NAND2_X1 U10559 ( .A1(n11406), .A2(n12731), .ZN(n8176) );
  NAND2_X1 U10560 ( .A1(n8177), .A2(n8176), .ZN(n11393) );
  XNOR2_X1 U10561 ( .A(n13167), .B(n12730), .ZN(n11394) );
  OR2_X1 U10562 ( .A1(n13167), .A2(n12730), .ZN(n8178) );
  XNOR2_X1 U10563 ( .A(n13162), .B(n12648), .ZN(n9371) );
  OR2_X1 U10564 ( .A1(n13074), .A2(n12648), .ZN(n8180) );
  NOR2_X1 U10565 ( .A1(n13045), .A2(n13058), .ZN(n8181) );
  NAND2_X1 U10566 ( .A1(n13045), .A2(n13058), .ZN(n8182) );
  NAND2_X1 U10567 ( .A1(n8183), .A2(n8182), .ZN(n13025) );
  XNOR2_X1 U10568 ( .A(n13153), .B(n13014), .ZN(n13026) );
  NAND2_X1 U10569 ( .A1(n13025), .A2(n13026), .ZN(n8185) );
  NAND2_X1 U10570 ( .A1(n13036), .A2(n13014), .ZN(n8184) );
  NAND2_X1 U10571 ( .A1(n8185), .A2(n8184), .ZN(n13010) );
  AND2_X1 U10572 ( .A1(n13022), .A2(n12697), .ZN(n8186) );
  OR2_X1 U10573 ( .A1(n13022), .A2(n12697), .ZN(n8187) );
  AND2_X1 U10574 ( .A1(n13142), .A2(n12976), .ZN(n8188) );
  OR2_X1 U10575 ( .A1(n13129), .A2(n12621), .ZN(n8189) );
  NAND2_X1 U10576 ( .A1(n13124), .A2(n12931), .ZN(n9362) );
  INV_X1 U10577 ( .A(n9362), .ZN(n8190) );
  AOI21_X2 U10578 ( .B1(n12945), .B2(n9363), .A(n8190), .ZN(n12941) );
  INV_X1 U10579 ( .A(n12929), .ZN(n12940) );
  NOR2_X1 U10580 ( .A1(n12923), .A2(n12657), .ZN(n8191) );
  INV_X1 U10581 ( .A(n13103), .ZN(n12896) );
  OAI22_X1 U10582 ( .A1(n12883), .A2(n12884), .B1(n12896), .B2(n12870), .ZN(
        n12880) );
  AOI22_X1 U10583 ( .A1(n12880), .A2(n12879), .B1(n13096), .B2(n12887), .ZN(
        n8192) );
  NOR2_X1 U10584 ( .A1(n8193), .A2(n9952), .ZN(n10514) );
  INV_X1 U10585 ( .A(n9956), .ZN(n8220) );
  NAND2_X1 U10586 ( .A1(n10514), .A2(n8220), .ZN(n14715) );
  INV_X1 U10587 ( .A(n10471), .ZN(n14670) );
  AND2_X1 U10588 ( .A1(n10468), .A2(n14670), .ZN(n10469) );
  AND2_X2 U10589 ( .A1(n14716), .A2(n10779), .ZN(n10971) );
  OR2_X2 U10590 ( .A1(n12892), .A2(n13096), .ZN(n12873) );
  AND2_X1 U10591 ( .A1(n10942), .A2(n8194), .ZN(n8195) );
  NOR2_X2 U10592 ( .A1(n12873), .A2(n12858), .ZN(n12852) );
  AOI211_X1 U10593 ( .C1(n12858), .C2(n12873), .A(n10022), .B(n12852), .ZN(
        n12864) );
  AOI21_X1 U10594 ( .B1(n14660), .B2(n12858), .A(n12864), .ZN(n8196) );
  NOR4_X1 U10595 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n8200) );
  NOR4_X1 U10596 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n8199) );
  NOR4_X1 U10597 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8198) );
  NOR4_X1 U10598 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n8197) );
  NAND4_X1 U10599 ( .A1(n8200), .A2(n8199), .A3(n8198), .A4(n8197), .ZN(n8219)
         );
  NOR2_X1 U10600 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .ZN(
        n8204) );
  NOR4_X1 U10601 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n8203) );
  NOR4_X1 U10602 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n8202) );
  NOR4_X1 U10603 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8201) );
  NAND4_X1 U10604 ( .A1(n8204), .A2(n8203), .A3(n8202), .A4(n8201), .ZN(n8218)
         );
  NAND2_X1 U10605 ( .A1(n8207), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8206) );
  MUX2_X1 U10606 ( .A(n8206), .B(P2_IR_REG_31__SCAN_IN), .S(n8208), .Z(n8210)
         );
  NAND2_X1 U10607 ( .A1(n8210), .A2(n8214), .ZN(n11239) );
  XOR2_X1 U10608 ( .A(n11239), .B(n8211), .Z(n8217) );
  NAND2_X1 U10609 ( .A1(n8214), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8213) );
  OAI21_X1 U10610 ( .B1(n8214), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8216) );
  OAI21_X1 U10611 ( .B1(n8219), .B2(n8218), .A(n14630), .ZN(n9942) );
  NAND2_X1 U10612 ( .A1(n8220), .A2(n9958), .ZN(n9947) );
  NAND2_X1 U10613 ( .A1(n8221), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8223) );
  XNOR2_X1 U10614 ( .A(n8223), .B(n8222), .ZN(n9945) );
  AND2_X1 U10615 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9946), .ZN(n8224) );
  AND2_X1 U10616 ( .A1(n9947), .A2(n14637), .ZN(n8225) );
  NAND2_X1 U10617 ( .A1(n9942), .A2(n8225), .ZN(n10367) );
  OR2_X1 U10618 ( .A1(n14688), .A2(n8193), .ZN(n9943) );
  NOR2_X1 U10619 ( .A1(n10367), .A2(n9954), .ZN(n8230) );
  INV_X1 U10620 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14634) );
  NAND2_X1 U10621 ( .A1(n14630), .A2(n14634), .ZN(n8227) );
  NAND2_X1 U10622 ( .A1(n13203), .A2(n11239), .ZN(n8226) );
  NAND2_X1 U10623 ( .A1(n8227), .A2(n8226), .ZN(n10368) );
  INV_X1 U10624 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15046) );
  NAND2_X1 U10625 ( .A1(n14630), .A2(n15046), .ZN(n8229) );
  NAND2_X1 U10626 ( .A1(n13203), .A2(n11295), .ZN(n8228) );
  NAND2_X1 U10627 ( .A1(n8236), .A2(n14723), .ZN(n8233) );
  INV_X1 U10628 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8231) );
  OR2_X1 U10629 ( .A1(n14723), .A2(n8231), .ZN(n8232) );
  NAND2_X1 U10630 ( .A1(n8233), .A2(n8232), .ZN(P2_U3496) );
  INV_X1 U10631 ( .A(n14637), .ZN(n14635) );
  AND3_X1 U10632 ( .A1(n9942), .A2(n9943), .A3(n9947), .ZN(n8234) );
  NAND2_X1 U10633 ( .A1(n14636), .A2(n8234), .ZN(n8235) );
  INV_X2 U10634 ( .A(n14735), .ZN(n14737) );
  NAND2_X1 U10635 ( .A1(n8236), .A2(n14737), .ZN(n8238) );
  NAND2_X1 U10636 ( .A1(n14735), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8237) );
  NAND2_X1 U10637 ( .A1(n8238), .A2(n8237), .ZN(P2_U3528) );
  NAND2_X1 U10638 ( .A1(n9682), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U10639 ( .A1(n9687), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8240) );
  NAND2_X1 U10640 ( .A1(n8374), .A2(n8373), .ZN(n8242) );
  NAND2_X1 U10641 ( .A1(n9692), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8243) );
  NAND2_X1 U10642 ( .A1(n9658), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U10643 ( .A1(n9667), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8247) );
  NAND2_X1 U10644 ( .A1(n9671), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8249) );
  NAND2_X1 U10645 ( .A1(n9672), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8250) );
  NAND2_X1 U10646 ( .A1(n9683), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8252) );
  NAND2_X1 U10647 ( .A1(n8253), .A2(n8252), .ZN(n8473) );
  NAND2_X1 U10648 ( .A1(n9705), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8254) );
  NAND2_X1 U10649 ( .A1(n9748), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8257) );
  NAND2_X1 U10650 ( .A1(n9751), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8256) );
  NAND2_X1 U10651 ( .A1(n9755), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U10652 ( .A1(n9757), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8258) );
  NAND2_X1 U10653 ( .A1(n9819), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8261) );
  NAND2_X1 U10654 ( .A1(n9821), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8260) );
  NAND2_X1 U10655 ( .A1(n9914), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10656 ( .A1(n9924), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8262) );
  NAND2_X1 U10657 ( .A1(n10079), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8266) );
  NAND2_X1 U10658 ( .A1(n10083), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8265) );
  NAND2_X1 U10659 ( .A1(n10176), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8268) );
  NAND2_X1 U10660 ( .A1(n10178), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8267) );
  NAND2_X1 U10661 ( .A1(n10076), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U10662 ( .A1(n10081), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8269) );
  AND2_X1 U10663 ( .A1(n8270), .A2(n8269), .ZN(n8613) );
  NAND2_X1 U10664 ( .A1(n10129), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8273) );
  NAND2_X1 U10665 ( .A1(n10171), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8271) );
  NAND2_X1 U10666 ( .A1(n8273), .A2(n8271), .ZN(n8632) );
  INV_X1 U10667 ( .A(n8632), .ZN(n8272) );
  INV_X1 U10668 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10479) );
  NAND2_X1 U10669 ( .A1(n10479), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8276) );
  INV_X1 U10670 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10481) );
  NAND2_X1 U10671 ( .A1(n10481), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8274) );
  NAND2_X1 U10672 ( .A1(n8276), .A2(n8274), .ZN(n8645) );
  INV_X1 U10673 ( .A(n8645), .ZN(n8275) );
  NAND2_X1 U10674 ( .A1(n10582), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8279) );
  NAND2_X1 U10675 ( .A1(n10585), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8278) );
  AND2_X1 U10676 ( .A1(n8279), .A2(n8278), .ZN(n8659) );
  INV_X1 U10677 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11009) );
  NAND2_X1 U10678 ( .A1(n11009), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8283) );
  INV_X1 U10679 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11012) );
  NAND2_X1 U10680 ( .A1(n11012), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U10681 ( .A1(n8283), .A2(n8281), .ZN(n8684) );
  INV_X1 U10682 ( .A(n8684), .ZN(n8282) );
  INV_X1 U10683 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11151) );
  XNOR2_X1 U10684 ( .A(n11151), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U10685 ( .A1(n11151), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8285) );
  XNOR2_X1 U10686 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8703) );
  INV_X1 U10687 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8286) );
  INV_X1 U10688 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n15122) );
  NAND2_X1 U10689 ( .A1(n11297), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8288) );
  AND2_X1 U10690 ( .A1(n13991), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8290) );
  NAND2_X1 U10691 ( .A1(n13202), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8291) );
  INV_X1 U10692 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8293) );
  AND2_X1 U10693 ( .A1(n8293), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8294) );
  INV_X1 U10694 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n13989) );
  NAND2_X1 U10695 ( .A1(n13989), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8295) );
  AND2_X1 U10696 ( .A1(n13987), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U10697 ( .A1(n13982), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8298) );
  NAND2_X1 U10698 ( .A1(n11428), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8297) );
  AND2_X1 U10699 ( .A1(n8298), .A2(n8297), .ZN(n8775) );
  INV_X1 U10700 ( .A(n8775), .ZN(n8299) );
  INV_X1 U10701 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11427) );
  XNOR2_X1 U10702 ( .A(n11427), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n8357) );
  XNOR2_X1 U10703 ( .A(n8358), .B(n8357), .ZN(n11822) );
  AND2_X2 U10704 ( .A1(n8460), .A2(n8302), .ZN(n8564) );
  NOR2_X1 U10705 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_15__SCAN_IN), 
        .ZN(n8306) );
  NOR2_X1 U10706 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), 
        .ZN(n8305) );
  NOR2_X1 U10707 ( .A1(P3_IR_REG_23__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n8309) );
  INV_X1 U10708 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8321) );
  NAND2_X1 U10709 ( .A1(n11822), .A2(n8778), .ZN(n8324) );
  INV_X1 U10710 ( .A(SI_30_), .ZN(n11824) );
  OR2_X1 U10711 ( .A1(n6787), .A2(n11824), .ZN(n8323) );
  INV_X1 U10712 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8330) );
  INV_X1 U10713 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n11925) );
  INV_X1 U10714 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n11973) );
  INV_X1 U10715 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8334) );
  INV_X1 U10716 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n8336) );
  INV_X1 U10717 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15079) );
  INV_X1 U10718 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n11904) );
  INV_X1 U10719 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15102) );
  INV_X1 U10720 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8341) );
  INV_X1 U10721 ( .A(n12184), .ZN(n8348) );
  OR2_X2 U10722 ( .A1(n8346), .A2(n8343), .ZN(n8349) );
  INV_X1 U10723 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12518) );
  NAND2_X1 U10724 ( .A1(n8344), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8345) );
  INV_X1 U10725 ( .A(n8346), .ZN(n12517) );
  NAND2_X1 U10726 ( .A1(n8348), .A2(n8756), .ZN(n8784) );
  INV_X1 U10727 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n8354) );
  INV_X4 U10728 ( .A(n8653), .ZN(n8382) );
  NAND2_X1 U10729 ( .A1(n8382), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10730 ( .A1(n8769), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8352) );
  OAI211_X1 U10731 ( .C1(n8354), .C2(n8772), .A(n8353), .B(n8352), .ZN(n8355)
         );
  INV_X1 U10732 ( .A(n8355), .ZN(n8356) );
  NAND2_X1 U10733 ( .A1(n8784), .A2(n8356), .ZN(n11983) );
  INV_X1 U10734 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13980) );
  OAI22_X1 U10735 ( .A1(n8358), .A2(n8357), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n13980), .ZN(n8360) );
  XNOR2_X1 U10736 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n8359) );
  XNOR2_X1 U10737 ( .A(n8360), .B(n8359), .ZN(n12516) );
  NAND2_X1 U10738 ( .A1(n12516), .A2(n8778), .ZN(n8362) );
  OR2_X1 U10739 ( .A1(n6787), .A2(n15060), .ZN(n8361) );
  INV_X1 U10740 ( .A(P3_REG2_REG_31__SCAN_IN), .ZN(n12187) );
  NAND2_X1 U10741 ( .A1(n6449), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8365) );
  INV_X1 U10742 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n8363) );
  OR2_X1 U10743 ( .A1(n8653), .A2(n8363), .ZN(n8364) );
  OAI211_X1 U10744 ( .C1(n6436), .C2(n12187), .A(n8365), .B(n8364), .ZN(n8366)
         );
  INV_X1 U10745 ( .A(n8366), .ZN(n8367) );
  NOR2_X1 U10746 ( .A1(n12462), .A2(n12183), .ZN(n8925) );
  NAND2_X1 U10747 ( .A1(n8421), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U10748 ( .A1(n8405), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8371) );
  INV_X1 U10749 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8368) );
  OR2_X1 U10750 ( .A1(n6446), .A2(n8368), .ZN(n8370) );
  INV_X1 U10751 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10317) );
  AND4_X2 U10752 ( .A1(n8372), .A2(n8371), .A3(n8370), .A4(n8369), .ZN(n10708)
         );
  INV_X1 U10753 ( .A(n10708), .ZN(n14921) );
  OR2_X1 U10754 ( .A1(n8411), .A2(SI_2_), .ZN(n8381) );
  XNOR2_X1 U10755 ( .A(n8374), .B(n8373), .ZN(n9635) );
  OR2_X1 U10756 ( .A1(n8400), .A2(n9635), .ZN(n8380) );
  XNOR2_X2 U10757 ( .A(n8378), .B(n8377), .ZN(n10892) );
  OR2_X1 U10758 ( .A1(n6448), .A2(n10839), .ZN(n8379) );
  NAND2_X1 U10759 ( .A1(n10708), .A2(n9072), .ZN(n8808) );
  NAND2_X2 U10760 ( .A1(n8807), .A2(n8808), .ZN(n14905) );
  NAND2_X1 U10761 ( .A1(n6449), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U10762 ( .A1(n8421), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8384) );
  INV_X1 U10763 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n14739) );
  OR2_X1 U10764 ( .A1(n8781), .A2(n14739), .ZN(n8383) );
  INV_X1 U10765 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n14746) );
  NAND2_X1 U10766 ( .A1(n8387), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8388) );
  AND2_X1 U10767 ( .A1(n8398), .A2(n8388), .ZN(n9630) );
  OR2_X1 U10768 ( .A1(n8400), .A2(n9630), .ZN(n8389) );
  INV_X2 U10769 ( .A(n10124), .ZN(n11809) );
  NOR2_X4 U10770 ( .A1(n14918), .A2(n11809), .ZN(n14917) );
  NAND2_X1 U10771 ( .A1(n6450), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8395) );
  NAND2_X1 U10772 ( .A1(n8421), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8394) );
  INV_X1 U10773 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8391) );
  INV_X1 U10774 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n14932) );
  OR2_X1 U10775 ( .A1(n8781), .A2(n14932), .ZN(n8392) );
  AND4_X2 U10776 ( .A1(n8395), .A2(n8394), .A3(n8393), .A4(n8392), .ZN(n9066)
         );
  NAND2_X1 U10777 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8396) );
  INV_X1 U10778 ( .A(n8376), .ZN(n8397) );
  OR2_X1 U10779 ( .A1(n8411), .A2(n6916), .ZN(n8402) );
  XNOR2_X1 U10780 ( .A(n8399), .B(n8398), .ZN(n9634) );
  OR2_X1 U10781 ( .A1(n8400), .A2(n9634), .ZN(n8401) );
  OAI211_X1 U10782 ( .C1(n6448), .C2(n6852), .A(n8402), .B(n8401), .ZN(n9068)
         );
  INV_X1 U10783 ( .A(n9068), .ZN(n14916) );
  NAND2_X1 U10784 ( .A1(n14917), .A2(n8802), .ZN(n9064) );
  NAND2_X1 U10785 ( .A1(n9066), .A2(n9068), .ZN(n9067) );
  NAND2_X1 U10786 ( .A1(n9064), .A2(n9067), .ZN(n14904) );
  NAND2_X1 U10787 ( .A1(n8404), .A2(n8808), .ZN(n10700) );
  NAND2_X1 U10788 ( .A1(n6449), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10789 ( .A1(n8421), .A2(n10642), .ZN(n8409) );
  INV_X1 U10790 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8406) );
  OR2_X1 U10791 ( .A1(n8653), .A2(n8406), .ZN(n8408) );
  INV_X1 U10792 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n10852) );
  OR2_X1 U10793 ( .A1(n8781), .A2(n10852), .ZN(n8407) );
  OR2_X1 U10794 ( .A1(n8413), .A2(n8412), .ZN(n8414) );
  NAND2_X1 U10795 ( .A1(n8415), .A2(n8414), .ZN(n9624) );
  OR2_X1 U10796 ( .A1(n8617), .A2(n9624), .ZN(n8419) );
  INV_X1 U10797 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8417) );
  NAND2_X1 U10798 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6504), .ZN(n8416) );
  XNOR2_X1 U10799 ( .A(n8417), .B(n8416), .ZN(n10854) );
  OR2_X1 U10800 ( .A1(n6448), .A2(n14765), .ZN(n8418) );
  AND3_X2 U10801 ( .A1(n8420), .A2(n8419), .A3(n8418), .ZN(n10703) );
  NAND2_X1 U10802 ( .A1(n14902), .A2(n10703), .ZN(n8811) );
  INV_X2 U10803 ( .A(n14902), .ZN(n11995) );
  INV_X1 U10804 ( .A(n10703), .ZN(n10636) );
  NAND2_X1 U10805 ( .A1(n8811), .A2(n8812), .ZN(n10705) );
  INV_X1 U10806 ( .A(n10705), .ZN(n10699) );
  NAND2_X1 U10807 ( .A1(n10700), .A2(n10699), .ZN(n10702) );
  NAND2_X1 U10808 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8422) );
  NAND2_X1 U10809 ( .A1(n8439), .A2(n8422), .ZN(n10688) );
  NAND2_X1 U10810 ( .A1(n8756), .A2(n10688), .ZN(n8427) );
  NAND2_X1 U10811 ( .A1(n6450), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8426) );
  INV_X1 U10812 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8423) );
  OR2_X1 U10813 ( .A1(n8653), .A2(n8423), .ZN(n8425) );
  INV_X1 U10814 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10896) );
  OR2_X1 U10815 ( .A1(n6436), .A2(n10896), .ZN(n8424) );
  OR2_X1 U10816 ( .A1(n8411), .A2(SI_4_), .ZN(n8436) );
  XNOR2_X1 U10817 ( .A(n8429), .B(n8428), .ZN(n9641) );
  OR2_X1 U10818 ( .A1(n8617), .A2(n9641), .ZN(n8435) );
  NAND2_X1 U10819 ( .A1(n8430), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8431) );
  MUX2_X1 U10820 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8431), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n8433) );
  AND2_X1 U10821 ( .A1(n8433), .A2(n8432), .ZN(n10895) );
  OR2_X1 U10822 ( .A1(n6448), .A2(n10895), .ZN(n8434) );
  NAND2_X1 U10823 ( .A1(n10707), .A2(n10695), .ZN(n8816) );
  INV_X1 U10824 ( .A(n10695), .ZN(n8437) );
  NAND2_X1 U10825 ( .A1(n11994), .A2(n8437), .ZN(n8817) );
  NAND2_X1 U10826 ( .A1(n8816), .A2(n8817), .ZN(n10646) );
  NAND2_X1 U10827 ( .A1(n10645), .A2(n10644), .ZN(n8438) );
  NAND2_X1 U10828 ( .A1(n8438), .A2(n8816), .ZN(n10614) );
  NAND2_X1 U10829 ( .A1(n6450), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8445) );
  NAND2_X1 U10830 ( .A1(n8439), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n8440) );
  NAND2_X1 U10831 ( .A1(n8453), .A2(n8440), .ZN(n10811) );
  NAND2_X1 U10832 ( .A1(n8756), .A2(n10811), .ZN(n8444) );
  INV_X1 U10833 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8441) );
  OR2_X1 U10834 ( .A1(n8653), .A2(n8441), .ZN(n8443) );
  INV_X1 U10835 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10862) );
  OR2_X1 U10836 ( .A1(n6436), .A2(n10862), .ZN(n8442) );
  OR2_X1 U10837 ( .A1(n6787), .A2(SI_5_), .ZN(n8451) );
  XNOR2_X1 U10838 ( .A(n8447), .B(n8446), .ZN(n9644) );
  OR2_X1 U10839 ( .A1(n8617), .A2(n9644), .ZN(n8450) );
  NAND2_X1 U10840 ( .A1(n8432), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8448) );
  XNOR2_X1 U10841 ( .A(n8448), .B(n7351), .ZN(n14793) );
  INV_X1 U10842 ( .A(n14793), .ZN(n10898) );
  OR2_X1 U10843 ( .A1(n10134), .A2(n10898), .ZN(n8449) );
  NAND2_X1 U10844 ( .A1(n10948), .A2(n10630), .ZN(n8798) );
  INV_X1 U10845 ( .A(n10630), .ZN(n10809) );
  NAND2_X1 U10846 ( .A1(n10832), .A2(n10809), .ZN(n8822) );
  NAND2_X1 U10847 ( .A1(n10614), .A2(n10616), .ZN(n8452) );
  NAND2_X1 U10848 ( .A1(n8453), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8454) );
  NAND2_X1 U10849 ( .A1(n8466), .A2(n8454), .ZN(n10959) );
  NAND2_X1 U10850 ( .A1(n8756), .A2(n10959), .ZN(n8459) );
  NAND2_X1 U10851 ( .A1(n6449), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8458) );
  INV_X1 U10852 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8455) );
  OR2_X1 U10853 ( .A1(n8653), .A2(n8455), .ZN(n8457) );
  INV_X1 U10854 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10957) );
  OR2_X1 U10855 ( .A1(n6436), .A2(n10957), .ZN(n8456) );
  OR2_X1 U10856 ( .A1(n8460), .A2(n7027), .ZN(n8461) );
  XNOR2_X1 U10857 ( .A(n8461), .B(n8477), .ZN(n14809) );
  INV_X1 U10858 ( .A(SI_6_), .ZN(n9622) );
  OR2_X1 U10859 ( .A1(n8411), .A2(n9622), .ZN(n8465) );
  XNOR2_X1 U10860 ( .A(n9672), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8462) );
  XNOR2_X1 U10861 ( .A(n8463), .B(n8462), .ZN(n9623) );
  OR2_X1 U10862 ( .A1(n8617), .A2(n9623), .ZN(n8464) );
  OAI211_X1 U10863 ( .C1(n10134), .C2(n14809), .A(n8465), .B(n8464), .ZN(
        n10958) );
  NAND2_X1 U10864 ( .A1(n10920), .A2(n10958), .ZN(n8826) );
  INV_X1 U10865 ( .A(n10958), .ZN(n9079) );
  NAND2_X1 U10866 ( .A1(n11993), .A2(n9079), .ZN(n8824) );
  NAND2_X1 U10867 ( .A1(n8826), .A2(n8824), .ZN(n10950) );
  INV_X1 U10868 ( .A(n10950), .ZN(n10945) );
  NAND2_X1 U10869 ( .A1(n8466), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8467) );
  NAND2_X1 U10870 ( .A1(n8483), .A2(n8467), .ZN(n10977) );
  NAND2_X1 U10871 ( .A1(n8756), .A2(n10977), .ZN(n8472) );
  NAND2_X1 U10872 ( .A1(n6449), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8471) );
  INV_X1 U10873 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10872) );
  OR2_X1 U10874 ( .A1(n6436), .A2(n10872), .ZN(n8470) );
  INV_X1 U10875 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8468) );
  OR2_X1 U10876 ( .A1(n6446), .A2(n8468), .ZN(n8469) );
  OR2_X1 U10877 ( .A1(n6787), .A2(SI_7_), .ZN(n8482) );
  NAND2_X1 U10878 ( .A1(n8474), .A2(n8473), .ZN(n8475) );
  AND2_X1 U10879 ( .A1(n8476), .A2(n8475), .ZN(n9638) );
  OR2_X1 U10880 ( .A1(n8617), .A2(n9638), .ZN(n8481) );
  NAND2_X1 U10881 ( .A1(n8460), .A2(n8477), .ZN(n8490) );
  NAND2_X1 U10882 ( .A1(n8490), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8479) );
  XNOR2_X1 U10883 ( .A(n8479), .B(n8478), .ZN(n10900) );
  INV_X1 U10884 ( .A(n10900), .ZN(n14829) );
  OR2_X1 U10885 ( .A1(n6448), .A2(n14829), .ZN(n8480) );
  NAND2_X1 U10886 ( .A1(n10947), .A2(n14961), .ZN(n8827) );
  INV_X1 U10887 ( .A(n14961), .ZN(n10925) );
  NAND2_X1 U10888 ( .A1(n14888), .A2(n10925), .ZN(n8828) );
  NAND2_X1 U10889 ( .A1(n8827), .A2(n8828), .ZN(n14881) );
  NAND2_X1 U10890 ( .A1(n8769), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8489) );
  NAND2_X1 U10891 ( .A1(n8483), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U10892 ( .A1(n8504), .A2(n8484), .ZN(n14895) );
  NAND2_X1 U10893 ( .A1(n8756), .A2(n14895), .ZN(n8488) );
  NAND2_X1 U10894 ( .A1(n6450), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8487) );
  INV_X1 U10895 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8485) );
  OR2_X1 U10896 ( .A1(n6446), .A2(n8485), .ZN(n8486) );
  NAND4_X1 U10897 ( .A1(n8489), .A2(n8488), .A3(n8487), .A4(n8486), .ZN(n11992) );
  INV_X1 U10898 ( .A(n8530), .ZN(n8495) );
  NAND2_X1 U10899 ( .A1(n8491), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8493) );
  MUX2_X1 U10900 ( .A(n8493), .B(P3_IR_REG_31__SCAN_IN), .S(n8492), .Z(n8494)
         );
  NAND2_X1 U10901 ( .A1(n8495), .A2(n8494), .ZN(n14847) );
  INV_X1 U10902 ( .A(SI_8_), .ZN(n9628) );
  OR2_X1 U10903 ( .A1(n6787), .A2(n9628), .ZN(n8501) );
  OR2_X1 U10904 ( .A1(n8497), .A2(n8496), .ZN(n8498) );
  NAND2_X1 U10905 ( .A1(n8499), .A2(n8498), .ZN(n9627) );
  OR2_X1 U10906 ( .A1(n8617), .A2(n9627), .ZN(n8500) );
  OAI211_X1 U10907 ( .C1(n10134), .C2(n14847), .A(n8501), .B(n8500), .ZN(
        n11171) );
  XNOR2_X1 U10908 ( .A(n11992), .B(n11171), .ZN(n14886) );
  NAND2_X1 U10909 ( .A1(n14880), .A2(n14886), .ZN(n8503) );
  NAND2_X1 U10910 ( .A1(n11155), .A2(n11171), .ZN(n8502) );
  NAND2_X1 U10911 ( .A1(n8382), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U10912 ( .A1(n6450), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8508) );
  NAND2_X1 U10913 ( .A1(n8504), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U10914 ( .A1(n8518), .A2(n8505), .ZN(n11308) );
  NAND2_X1 U10915 ( .A1(n8756), .A2(n11308), .ZN(n8507) );
  INV_X1 U10916 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11272) );
  OR2_X1 U10917 ( .A1(n6436), .A2(n11272), .ZN(n8506) );
  OR2_X1 U10918 ( .A1(n8511), .A2(n8510), .ZN(n8512) );
  AND2_X1 U10919 ( .A1(n8513), .A2(n8512), .ZN(n9631) );
  OR2_X1 U10920 ( .A1(n8617), .A2(n9631), .ZN(n8517) );
  OR2_X1 U10921 ( .A1(n6787), .A2(SI_9_), .ZN(n8516) );
  OR2_X1 U10922 ( .A1(n8530), .A2(n8343), .ZN(n8514) );
  INV_X1 U10923 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n8529) );
  XNOR2_X1 U10924 ( .A(n8514), .B(n8529), .ZN(n14867) );
  INV_X1 U10925 ( .A(n14867), .ZN(n10905) );
  OR2_X1 U10926 ( .A1(n10134), .A2(n10905), .ZN(n8515) );
  NOR2_X1 U10927 ( .A1(n14887), .A2(n11306), .ZN(n8835) );
  NAND2_X1 U10928 ( .A1(n14887), .A2(n11306), .ZN(n8837) );
  NAND2_X1 U10929 ( .A1(n8518), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U10930 ( .A1(n8536), .A2(n8519), .ZN(n11251) );
  NAND2_X1 U10931 ( .A1(n8756), .A2(n11251), .ZN(n8524) );
  NAND2_X1 U10932 ( .A1(n6449), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8523) );
  INV_X1 U10933 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8520) );
  OR2_X1 U10934 ( .A1(n8653), .A2(n8520), .ZN(n8522) );
  INV_X1 U10935 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n10907) );
  OR2_X1 U10936 ( .A1(n6436), .A2(n10907), .ZN(n8521) );
  OR2_X1 U10937 ( .A1(n8526), .A2(n8525), .ZN(n8527) );
  AND2_X1 U10938 ( .A1(n8528), .A2(n8527), .ZN(n9650) );
  OR2_X1 U10939 ( .A1(n8617), .A2(n9650), .ZN(n8534) );
  OR2_X1 U10940 ( .A1(n6787), .A2(SI_10_), .ZN(n8533) );
  NAND2_X1 U10941 ( .A1(n8530), .A2(n8529), .ZN(n8547) );
  NAND2_X1 U10942 ( .A1(n8547), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8531) );
  XNOR2_X1 U10943 ( .A(n8531), .B(P3_IR_REG_10__SCAN_IN), .ZN(n11098) );
  OR2_X1 U10944 ( .A1(n10134), .A2(n11098), .ZN(n8532) );
  NAND2_X1 U10945 ( .A1(n11303), .A2(n11370), .ZN(n8840) );
  INV_X1 U10946 ( .A(n11370), .ZN(n8535) );
  NAND2_X1 U10947 ( .A1(n11991), .A2(n8535), .ZN(n8841) );
  NAND2_X1 U10948 ( .A1(n8840), .A2(n8841), .ZN(n11247) );
  NAND2_X1 U10949 ( .A1(n8536), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U10950 ( .A1(n8553), .A2(n8537), .ZN(n11948) );
  NAND2_X1 U10951 ( .A1(n8756), .A2(n11948), .ZN(n8542) );
  NAND2_X1 U10952 ( .A1(n6450), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8541) );
  INV_X1 U10953 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n8538) );
  OR2_X1 U10954 ( .A1(n8653), .A2(n8538), .ZN(n8540) );
  INV_X1 U10955 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11384) );
  OR2_X1 U10956 ( .A1(n6436), .A2(n11384), .ZN(n8539) );
  OR2_X1 U10957 ( .A1(n8544), .A2(n8543), .ZN(n8545) );
  NAND2_X1 U10958 ( .A1(n8546), .A2(n8545), .ZN(n9661) );
  NAND2_X1 U10959 ( .A1(n8778), .A2(n9661), .ZN(n8552) );
  OR2_X1 U10960 ( .A1(n6787), .A2(SI_11_), .ZN(n8551) );
  OAI21_X1 U10961 ( .B1(n8547), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8549) );
  INV_X1 U10962 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8548) );
  XNOR2_X1 U10963 ( .A(n8549), .B(n8548), .ZN(n12018) );
  INV_X1 U10964 ( .A(n12018), .ZN(n12007) );
  OR2_X1 U10965 ( .A1(n10134), .A2(n12007), .ZN(n8550) );
  NAND2_X1 U10966 ( .A1(n11945), .A2(n11381), .ZN(n8843) );
  INV_X1 U10967 ( .A(n11381), .ZN(n11942) );
  NAND2_X1 U10968 ( .A1(n11866), .A2(n11942), .ZN(n8847) );
  NAND2_X1 U10969 ( .A1(n8843), .A2(n8847), .ZN(n11377) );
  NAND2_X1 U10970 ( .A1(n8553), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8554) );
  NAND2_X1 U10971 ( .A1(n8577), .A2(n8554), .ZN(n11870) );
  NAND2_X1 U10972 ( .A1(n8756), .A2(n11870), .ZN(n8559) );
  NAND2_X1 U10973 ( .A1(n6450), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8558) );
  INV_X1 U10974 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8555) );
  OR2_X1 U10975 ( .A1(n6446), .A2(n8555), .ZN(n8557) );
  INV_X1 U10976 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n12010) );
  OR2_X1 U10977 ( .A1(n6436), .A2(n12010), .ZN(n8556) );
  OR2_X1 U10978 ( .A1(n8561), .A2(n8560), .ZN(n8562) );
  NAND2_X1 U10979 ( .A1(n8563), .A2(n8562), .ZN(n9674) );
  OR2_X1 U10980 ( .A1(n9674), .A2(n8617), .ZN(n8570) );
  NOR2_X1 U10981 ( .A1(n8564), .A2(n8343), .ZN(n8565) );
  MUX2_X1 U10982 ( .A(n7027), .B(n8565), .S(P3_IR_REG_12__SCAN_IN), .Z(n8568)
         );
  INV_X1 U10983 ( .A(n8566), .ZN(n8567) );
  INV_X1 U10984 ( .A(n12036), .ZN(n12033) );
  AOI22_X1 U10985 ( .A1(n8663), .A2(SI_12_), .B1(n8662), .B2(n12033), .ZN(
        n8569) );
  NAND2_X1 U10986 ( .A1(n8570), .A2(n8569), .ZN(n14167) );
  NAND2_X1 U10987 ( .A1(n11937), .A2(n14167), .ZN(n8851) );
  INV_X1 U10988 ( .A(n14167), .ZN(n11868) );
  NAND2_X1 U10989 ( .A1(n11868), .A2(n11990), .ZN(n8849) );
  NAND2_X1 U10990 ( .A1(n8851), .A2(n8849), .ZN(n11353) );
  INV_X1 U10991 ( .A(n11353), .ZN(n11356) );
  NAND2_X1 U10992 ( .A1(n8571), .A2(n10012), .ZN(n8572) );
  NAND2_X1 U10993 ( .A1(n8573), .A2(n8572), .ZN(n9714) );
  OR2_X1 U10994 ( .A1(n9714), .A2(n8617), .ZN(n8576) );
  NAND2_X1 U10995 ( .A1(n8566), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8574) );
  XNOR2_X1 U10996 ( .A(n8574), .B(P3_IR_REG_13__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U10997 ( .A1(n8663), .A2(SI_13_), .B1(n8662), .B2(n12061), .ZN(
        n8575) );
  NAND2_X1 U10998 ( .A1(n8382), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U10999 ( .A1(n8577), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U11000 ( .A1(n8591), .A2(n8578), .ZN(n11924) );
  NAND2_X1 U11001 ( .A1(n8756), .A2(n11924), .ZN(n8582) );
  NAND2_X1 U11002 ( .A1(n6449), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8581) );
  INV_X1 U11003 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n8579) );
  OR2_X1 U11004 ( .A1(n6436), .A2(n8579), .ZN(n8580) );
  OR2_X1 U11005 ( .A1(n14162), .A2(n12384), .ZN(n8853) );
  NAND2_X1 U11006 ( .A1(n14162), .A2(n12384), .ZN(n8852) );
  OR2_X1 U11007 ( .A1(n8585), .A2(n8584), .ZN(n8586) );
  NAND2_X1 U11008 ( .A1(n8587), .A2(n8586), .ZN(n9775) );
  OR2_X1 U11009 ( .A1(n9775), .A2(n8617), .ZN(n8590) );
  XNOR2_X1 U11010 ( .A(n8588), .B(P3_IR_REG_14__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U11011 ( .A1(n8663), .A2(SI_14_), .B1(n8662), .B2(n12071), .ZN(
        n8589) );
  NAND2_X1 U11012 ( .A1(n8590), .A2(n8589), .ZN(n12388) );
  NAND2_X1 U11013 ( .A1(n8591), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U11014 ( .A1(n8606), .A2(n8592), .ZN(n12389) );
  NAND2_X1 U11015 ( .A1(n8756), .A2(n12389), .ZN(n8596) );
  NAND2_X1 U11016 ( .A1(n6449), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8595) );
  INV_X1 U11017 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12051) );
  OR2_X1 U11018 ( .A1(n6436), .A2(n12051), .ZN(n8594) );
  INV_X1 U11019 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12508) );
  OR2_X1 U11020 ( .A1(n6446), .A2(n12508), .ZN(n8593) );
  OR2_X1 U11021 ( .A1(n12388), .A2(n12369), .ZN(n8858) );
  NAND2_X1 U11022 ( .A1(n12386), .A2(n8858), .ZN(n8597) );
  NAND2_X1 U11023 ( .A1(n12388), .A2(n12369), .ZN(n8857) );
  OR2_X1 U11024 ( .A1(n8599), .A2(n8598), .ZN(n8600) );
  NAND2_X1 U11025 ( .A1(n8601), .A2(n8600), .ZN(n9814) );
  OR2_X1 U11026 ( .A1(n9814), .A2(n8617), .ZN(n8605) );
  NAND2_X1 U11027 ( .A1(n8618), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8603) );
  INV_X1 U11028 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8602) );
  XNOR2_X1 U11029 ( .A(n8603), .B(n8602), .ZN(n12112) );
  INV_X1 U11030 ( .A(n12112), .ZN(n12087) );
  AOI22_X1 U11031 ( .A1(n8663), .A2(SI_15_), .B1(n8662), .B2(n12087), .ZN(
        n8604) );
  NAND2_X1 U11032 ( .A1(n6449), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8612) );
  NAND2_X1 U11033 ( .A1(n8606), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8607) );
  NAND2_X1 U11034 ( .A1(n8626), .A2(n8607), .ZN(n12376) );
  NAND2_X1 U11035 ( .A1(n8756), .A2(n12376), .ZN(n8611) );
  INV_X1 U11036 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n8608) );
  OR2_X1 U11037 ( .A1(n8653), .A2(n8608), .ZN(n8610) );
  INV_X1 U11038 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12089) );
  OR2_X1 U11039 ( .A1(n6436), .A2(n12089), .ZN(n8609) );
  OR2_X1 U11040 ( .A1(n12452), .A2(n12385), .ZN(n8862) );
  NAND2_X1 U11041 ( .A1(n12452), .A2(n12385), .ZN(n8861) );
  NAND2_X1 U11042 ( .A1(n8862), .A2(n8861), .ZN(n9000) );
  INV_X1 U11043 ( .A(n9000), .ZN(n12372) );
  OR2_X1 U11044 ( .A1(n8614), .A2(n8613), .ZN(n8615) );
  NAND2_X1 U11045 ( .A1(n8616), .A2(n8615), .ZN(n9845) );
  NOR2_X1 U11046 ( .A1(n8621), .A2(n8343), .ZN(n8619) );
  MUX2_X1 U11047 ( .A(n7027), .B(n8619), .S(P3_IR_REG_16__SCAN_IN), .Z(n8623)
         );
  INV_X1 U11048 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8620) );
  NAND2_X1 U11049 ( .A1(n8621), .A2(n8620), .ZN(n8647) );
  INV_X1 U11050 ( .A(n8647), .ZN(n8622) );
  NOR2_X1 U11051 ( .A1(n8623), .A2(n8622), .ZN(n12126) );
  AOI22_X1 U11052 ( .A1(n8663), .A2(SI_16_), .B1(n8662), .B2(n12126), .ZN(
        n8624) );
  NAND2_X1 U11053 ( .A1(n8626), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11054 ( .A1(n8637), .A2(n8627), .ZN(n12362) );
  NAND2_X1 U11055 ( .A1(n8756), .A2(n12362), .ZN(n8631) );
  NAND2_X1 U11056 ( .A1(n6450), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8630) );
  INV_X1 U11057 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12125) );
  OR2_X1 U11058 ( .A1(n6436), .A2(n12125), .ZN(n8629) );
  INV_X1 U11059 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12503) );
  OR2_X1 U11060 ( .A1(n8653), .A2(n12503), .ZN(n8628) );
  OR2_X1 U11061 ( .A1(n12361), .A2(n12368), .ZN(n8866) );
  NAND2_X1 U11062 ( .A1(n12361), .A2(n12368), .ZN(n8865) );
  NAND2_X1 U11063 ( .A1(n8866), .A2(n8865), .ZN(n12356) );
  INV_X1 U11064 ( .A(n12356), .ZN(n12359) );
  XNOR2_X1 U11065 ( .A(n8633), .B(n8632), .ZN(n9937) );
  NAND2_X1 U11066 ( .A1(n9937), .A2(n8778), .ZN(n8636) );
  NAND2_X1 U11067 ( .A1(n8647), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8634) );
  XNOR2_X1 U11068 ( .A(n8634), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U11069 ( .A1(n8663), .A2(SI_17_), .B1(n8662), .B2(n12151), .ZN(
        n8635) );
  NAND2_X1 U11070 ( .A1(n8637), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U11071 ( .A1(n8651), .A2(n8638), .ZN(n12350) );
  NAND2_X1 U11072 ( .A1(n8756), .A2(n12350), .ZN(n8644) );
  NAND2_X1 U11073 ( .A1(n6450), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8643) );
  INV_X1 U11074 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n8639) );
  OR2_X1 U11075 ( .A1(n6436), .A2(n8639), .ZN(n8642) );
  INV_X1 U11076 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n8640) );
  OR2_X1 U11077 ( .A1(n6446), .A2(n8640), .ZN(n8641) );
  OR2_X1 U11078 ( .A1(n12444), .A2(n12358), .ZN(n8871) );
  NAND2_X1 U11079 ( .A1(n12444), .A2(n12358), .ZN(n12335) );
  NAND2_X1 U11080 ( .A1(n8871), .A2(n12335), .ZN(n9004) );
  XNOR2_X1 U11081 ( .A(n8646), .B(n8645), .ZN(n10014) );
  NAND2_X1 U11082 ( .A1(n10014), .A2(n8778), .ZN(n8650) );
  NAND2_X1 U11083 ( .A1(n6565), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8648) );
  XNOR2_X1 U11084 ( .A(n8648), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U11085 ( .A1(n8663), .A2(SI_18_), .B1(n8662), .B2(n12165), .ZN(
        n8649) );
  NAND2_X1 U11086 ( .A1(n8650), .A2(n8649), .ZN(n11954) );
  NAND2_X1 U11087 ( .A1(n8651), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U11088 ( .A1(n8666), .A2(n8652), .ZN(n12338) );
  NAND2_X1 U11089 ( .A1(n8756), .A2(n12338), .ZN(n8657) );
  NAND2_X1 U11090 ( .A1(n6450), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8656) );
  INV_X1 U11091 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12130) );
  OR2_X1 U11092 ( .A1(n6436), .A2(n12130), .ZN(n8655) );
  INV_X1 U11093 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12498) );
  OR2_X1 U11094 ( .A1(n8653), .A2(n12498), .ZN(n8654) );
  NAND2_X1 U11095 ( .A1(n11954), .A2(n9007), .ZN(n8876) );
  INV_X1 U11096 ( .A(n12335), .ZN(n8875) );
  NOR2_X1 U11097 ( .A1(n9005), .A2(n8875), .ZN(n8658) );
  NAND2_X1 U11098 ( .A1(n12333), .A2(n8872), .ZN(n12317) );
  INV_X1 U11099 ( .A(n12317), .ZN(n8672) );
  XNOR2_X1 U11100 ( .A(n8660), .B(n8659), .ZN(n10019) );
  NAND2_X1 U11101 ( .A1(n10019), .A2(n8778), .ZN(n8665) );
  INV_X1 U11102 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8661) );
  AOI22_X1 U11103 ( .A1(n8663), .A2(n10018), .B1(n8662), .B2(n12177), .ZN(
        n8664) );
  NAND2_X1 U11104 ( .A1(n8382), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U11105 ( .A1(n8666), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11106 ( .A1(n8678), .A2(n8667), .ZN(n12322) );
  NAND2_X1 U11107 ( .A1(n8756), .A2(n12322), .ZN(n8670) );
  NAND2_X1 U11108 ( .A1(n6450), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8669) );
  INV_X1 U11109 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12161) );
  OR2_X1 U11110 ( .A1(n6436), .A2(n12161), .ZN(n8668) );
  NAND4_X1 U11111 ( .A1(n8671), .A2(n8670), .A3(n8669), .A4(n8668), .ZN(n12305) );
  NAND2_X1 U11112 ( .A1(n12496), .A2(n12305), .ZN(n8928) );
  XNOR2_X1 U11113 ( .A(n8673), .B(n11007), .ZN(n10166) );
  NAND2_X1 U11114 ( .A1(n10166), .A2(n8778), .ZN(n8675) );
  OR2_X1 U11115 ( .A1(n6787), .A2(n10167), .ZN(n8674) );
  NAND2_X1 U11116 ( .A1(n8769), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8677) );
  NAND2_X1 U11117 ( .A1(n8382), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n8676) );
  AND2_X1 U11118 ( .A1(n8677), .A2(n8676), .ZN(n8682) );
  NAND2_X1 U11119 ( .A1(n8678), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U11120 ( .A1(n8688), .A2(n8679), .ZN(n12312) );
  NAND2_X1 U11121 ( .A1(n12312), .A2(n8756), .ZN(n8681) );
  NAND2_X1 U11122 ( .A1(n6449), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8680) );
  INV_X1 U11123 ( .A(n12311), .ZN(n8683) );
  OR2_X1 U11124 ( .A1(n12432), .A2(n12295), .ZN(n8883) );
  XNOR2_X1 U11125 ( .A(n8685), .B(n8684), .ZN(n10193) );
  NAND2_X1 U11126 ( .A1(n10193), .A2(n8778), .ZN(n8687) );
  INV_X1 U11127 ( .A(SI_21_), .ZN(n10194) );
  INV_X1 U11128 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12430) );
  NAND2_X1 U11129 ( .A1(n8688), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8689) );
  NAND2_X1 U11130 ( .A1(n8697), .A2(n8689), .ZN(n12299) );
  NAND2_X1 U11131 ( .A1(n12299), .A2(n8756), .ZN(n8691) );
  AOI22_X1 U11132 ( .A1(n8769), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n8382), .B2(
        P3_REG0_REG_21__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U11133 ( .A1(n12298), .A2(n12283), .ZN(n8890) );
  NAND2_X1 U11134 ( .A1(n12297), .A2(n8890), .ZN(n8692) );
  OR2_X1 U11135 ( .A1(n12298), .A2(n12283), .ZN(n8889) );
  NAND2_X1 U11136 ( .A1(n8692), .A2(n8889), .ZN(n12285) );
  INV_X1 U11137 ( .A(n12285), .ZN(n8702) );
  XNOR2_X1 U11138 ( .A(n8694), .B(n8693), .ZN(n10197) );
  OR2_X1 U11139 ( .A1(n6787), .A2(n8695), .ZN(n8696) );
  INV_X1 U11140 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n15025) );
  NAND2_X1 U11141 ( .A1(n8697), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8698) );
  NAND2_X1 U11142 ( .A1(n8707), .A2(n8698), .ZN(n12287) );
  NAND2_X1 U11143 ( .A1(n12287), .A2(n8756), .ZN(n8700) );
  AOI22_X1 U11144 ( .A1(n8769), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n8382), .B2(
        P3_REG0_REG_22__SCAN_IN), .ZN(n8699) );
  NOR2_X1 U11145 ( .A1(n12286), .A2(n12294), .ZN(n8893) );
  INV_X1 U11146 ( .A(n8893), .ZN(n8701) );
  XNOR2_X1 U11147 ( .A(n8704), .B(n8703), .ZN(n10510) );
  NAND2_X1 U11148 ( .A1(n10510), .A2(n8778), .ZN(n8706) );
  OR2_X1 U11149 ( .A1(n6787), .A2(n10513), .ZN(n8705) );
  NAND2_X1 U11150 ( .A1(n8707), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8708) );
  NAND2_X1 U11151 ( .A1(n8718), .A2(n8708), .ZN(n12270) );
  NAND2_X1 U11152 ( .A1(n12270), .A2(n8756), .ZN(n8713) );
  INV_X1 U11153 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12273) );
  NAND2_X1 U11154 ( .A1(n6450), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U11155 ( .A1(n8382), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8709) );
  OAI211_X1 U11156 ( .C1(n6436), .C2(n12273), .A(n8710), .B(n8709), .ZN(n8711)
         );
  INV_X1 U11157 ( .A(n8711), .ZN(n8712) );
  NAND2_X1 U11158 ( .A1(n12276), .A2(n12282), .ZN(n8714) );
  INV_X1 U11159 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n15035) );
  NAND2_X1 U11160 ( .A1(n10801), .A2(n8778), .ZN(n8717) );
  INV_X1 U11161 ( .A(SI_24_), .ZN(n10802) );
  NAND2_X1 U11162 ( .A1(n8718), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U11163 ( .A1(n8728), .A2(n8719), .ZN(n12255) );
  INV_X1 U11164 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12418) );
  NAND2_X1 U11165 ( .A1(n8769), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U11166 ( .A1(n8382), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8720) );
  OAI211_X1 U11167 ( .C1(n12418), .C2(n8772), .A(n8721), .B(n8720), .ZN(n8722)
         );
  NAND2_X1 U11168 ( .A1(n9132), .A2(n12266), .ZN(n8897) );
  INV_X1 U11169 ( .A(n8899), .ZN(n12251) );
  NOR2_X1 U11170 ( .A1(n12250), .A2(n12251), .ZN(n8723) );
  NAND2_X1 U11171 ( .A1(n12262), .A2(n8723), .ZN(n12253) );
  XNOR2_X1 U11172 ( .A(n11297), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8724) );
  XNOR2_X1 U11173 ( .A(n8725), .B(n8724), .ZN(n11013) );
  NAND2_X1 U11174 ( .A1(n11013), .A2(n8778), .ZN(n8727) );
  NAND2_X1 U11175 ( .A1(n8728), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8729) );
  NAND2_X1 U11176 ( .A1(n8741), .A2(n8729), .ZN(n12241) );
  NAND2_X1 U11177 ( .A1(n12241), .A2(n8756), .ZN(n8735) );
  INV_X1 U11178 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n8732) );
  NAND2_X1 U11179 ( .A1(n8769), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8731) );
  NAND2_X1 U11180 ( .A1(n8382), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8730) );
  OAI211_X1 U11181 ( .C1(n8732), .C2(n8772), .A(n8731), .B(n8730), .ZN(n8733)
         );
  INV_X1 U11182 ( .A(n8733), .ZN(n8734) );
  NAND2_X1 U11183 ( .A1(n12413), .A2(n12249), .ZN(n8736) );
  INV_X1 U11184 ( .A(n8736), .ZN(n8905) );
  XNOR2_X1 U11185 ( .A(n13202), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8737) );
  XNOR2_X1 U11186 ( .A(n8738), .B(n8737), .ZN(n11198) );
  NAND2_X1 U11187 ( .A1(n11198), .A2(n8778), .ZN(n8740) );
  NAND2_X1 U11188 ( .A1(n8741), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8742) );
  NAND2_X1 U11189 ( .A1(n8754), .A2(n8742), .ZN(n12229) );
  NAND2_X1 U11190 ( .A1(n12229), .A2(n8756), .ZN(n8748) );
  INV_X1 U11191 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n8745) );
  NAND2_X1 U11192 ( .A1(n6449), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U11193 ( .A1(n8382), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8743) );
  OAI211_X1 U11194 ( .C1(n6436), .C2(n8745), .A(n8744), .B(n8743), .ZN(n8746)
         );
  INV_X1 U11195 ( .A(n8746), .ZN(n8747) );
  INV_X1 U11196 ( .A(n8909), .ZN(n8749) );
  XNOR2_X1 U11197 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8750) );
  XNOR2_X1 U11198 ( .A(n8751), .B(n8750), .ZN(n11258) );
  NAND2_X1 U11199 ( .A1(n11258), .A2(n8778), .ZN(n8753) );
  INV_X1 U11200 ( .A(SI_27_), .ZN(n11259) );
  NAND2_X1 U11201 ( .A1(n8754), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11202 ( .A1(n8767), .A2(n8755), .ZN(n12219) );
  NAND2_X1 U11203 ( .A1(n12219), .A2(n8756), .ZN(n8761) );
  INV_X1 U11204 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U11205 ( .A1(n8382), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U11206 ( .A1(n8769), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8757) );
  OAI211_X1 U11207 ( .C1(n8772), .C2(n12406), .A(n8758), .B(n8757), .ZN(n8759)
         );
  INV_X1 U11208 ( .A(n8759), .ZN(n8760) );
  NAND2_X1 U11209 ( .A1(n12218), .A2(n12217), .ZN(n12216) );
  NAND2_X1 U11210 ( .A1(n9063), .A2(n12226), .ZN(n8916) );
  NAND2_X1 U11211 ( .A1(n12216), .A2(n8916), .ZN(n12206) );
  XNOR2_X1 U11212 ( .A(n8762), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8763) );
  XNOR2_X1 U11213 ( .A(n8764), .B(n8763), .ZN(n12526) );
  NAND2_X1 U11214 ( .A1(n12526), .A2(n8778), .ZN(n8766) );
  OR2_X1 U11215 ( .A1(n6787), .A2(n12529), .ZN(n8765) );
  NAND2_X1 U11216 ( .A1(n8767), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U11217 ( .A1(n12184), .A2(n8768), .ZN(n12207) );
  INV_X1 U11218 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12402) );
  NAND2_X1 U11219 ( .A1(n8382), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U11220 ( .A1(n8769), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8770) );
  OAI211_X1 U11221 ( .C1(n12402), .C2(n8772), .A(n8771), .B(n8770), .ZN(n8773)
         );
  NAND2_X1 U11222 ( .A1(n11819), .A2(n12214), .ZN(n8774) );
  XNOR2_X1 U11223 ( .A(n8776), .B(n8775), .ZN(n12522) );
  INV_X1 U11224 ( .A(SI_29_), .ZN(n12523) );
  NOR2_X1 U11225 ( .A1(n6787), .A2(n12523), .ZN(n8777) );
  INV_X1 U11226 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n15048) );
  NAND2_X1 U11227 ( .A1(n8382), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U11228 ( .A1(n6450), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8779) );
  OAI211_X1 U11229 ( .C1(n15048), .C2(n6436), .A(n8780), .B(n8779), .ZN(n8782)
         );
  INV_X1 U11230 ( .A(n8782), .ZN(n8783) );
  NAND2_X1 U11231 ( .A1(n8784), .A2(n8783), .ZN(n11984) );
  NAND2_X1 U11232 ( .A1(n12193), .A2(n11984), .ZN(n8919) );
  OR2_X1 U11233 ( .A1(n12181), .A2(n8785), .ZN(n8926) );
  INV_X1 U11234 ( .A(n11983), .ZN(n8786) );
  NAND2_X1 U11235 ( .A1(n12463), .A2(n8786), .ZN(n8923) );
  NAND2_X1 U11236 ( .A1(n8926), .A2(n8923), .ZN(n8927) );
  INV_X1 U11237 ( .A(n11984), .ZN(n12204) );
  NAND2_X1 U11238 ( .A1(n8787), .A2(n12204), .ZN(n8920) );
  OAI21_X1 U11239 ( .B1(n12190), .B2(n12183), .A(n8920), .ZN(n8788) );
  NAND2_X1 U11240 ( .A1(n8791), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8790) );
  MUX2_X1 U11241 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8790), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8792) );
  INV_X1 U11242 ( .A(n8796), .ZN(n8793) );
  INV_X1 U11243 ( .A(n10169), .ZN(n9046) );
  NAND2_X1 U11244 ( .A1(n8793), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8794) );
  NAND2_X1 U11245 ( .A1(n9046), .A2(n10628), .ZN(n9019) );
  INV_X1 U11246 ( .A(n9060), .ZN(n8979) );
  AND2_X1 U11247 ( .A1(n9048), .A2(n10169), .ZN(n14911) );
  NAND2_X1 U11248 ( .A1(n8796), .A2(n8795), .ZN(n8952) );
  NAND2_X1 U11249 ( .A1(n8952), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8797) );
  INV_X1 U11250 ( .A(n12276), .ZN(n12420) );
  INV_X1 U11251 ( .A(n12282), .ZN(n11835) );
  AND2_X1 U11252 ( .A1(n8826), .A2(n8798), .ZN(n8821) );
  INV_X1 U11253 ( .A(n8982), .ZN(n10348) );
  AND2_X1 U11254 ( .A1(n14918), .A2(n11809), .ZN(n8930) );
  INV_X1 U11255 ( .A(n8930), .ZN(n8799) );
  NAND3_X1 U11256 ( .A1(n10348), .A2(n10198), .A3(n8799), .ZN(n8801) );
  OAI211_X1 U11257 ( .C1(n8930), .C2(n10196), .A(n9044), .B(n9067), .ZN(n8800)
         );
  AOI22_X1 U11258 ( .A1(n8801), .A2(n8800), .B1(n14917), .B2(n10196), .ZN(
        n8806) );
  INV_X1 U11259 ( .A(n8802), .ZN(n8804) );
  INV_X1 U11260 ( .A(n9067), .ZN(n8803) );
  MUX2_X1 U11261 ( .A(n8804), .B(n8803), .S(n10132), .Z(n8805) );
  NOR3_X1 U11262 ( .A1(n8806), .A2(n8805), .A3(n14905), .ZN(n8815) );
  NAND2_X1 U11263 ( .A1(n8812), .A2(n8807), .ZN(n8810) );
  NAND2_X1 U11264 ( .A1(n8811), .A2(n8808), .ZN(n8809) );
  MUX2_X1 U11265 ( .A(n8810), .B(n8809), .S(n9044), .Z(n8814) );
  MUX2_X1 U11266 ( .A(n8812), .B(n8811), .S(n10132), .Z(n8813) );
  OAI211_X1 U11267 ( .C1(n8815), .C2(n8814), .A(n10644), .B(n8813), .ZN(n8819)
         );
  MUX2_X1 U11268 ( .A(n8817), .B(n8816), .S(n9044), .Z(n8818) );
  NAND3_X1 U11269 ( .A1(n8819), .A2(n10616), .A3(n8818), .ZN(n8820) );
  OAI21_X1 U11270 ( .B1(n8821), .B2(n9044), .A(n8820), .ZN(n8825) );
  AOI21_X1 U11271 ( .B1(n8824), .B2(n8822), .A(n10132), .ZN(n8823) );
  AOI21_X1 U11272 ( .B1(n8825), .B2(n8824), .A(n8823), .ZN(n8831) );
  OAI21_X1 U11273 ( .B1(n10132), .B2(n8826), .A(n10918), .ZN(n8830) );
  MUX2_X1 U11274 ( .A(n8828), .B(n8827), .S(n10132), .Z(n8829) );
  OAI211_X1 U11275 ( .C1(n8831), .C2(n8830), .A(n14886), .B(n8829), .ZN(n8834)
         );
  XNOR2_X1 U11276 ( .A(n14887), .B(n11276), .ZN(n11153) );
  MUX2_X1 U11277 ( .A(n10132), .B(n11155), .S(n11171), .Z(n8832) );
  OAI21_X1 U11278 ( .B1(n9044), .B2(n11992), .A(n8832), .ZN(n8833) );
  NAND3_X1 U11279 ( .A1(n8834), .A2(n11153), .A3(n8833), .ZN(n8839) );
  INV_X1 U11280 ( .A(n8835), .ZN(n8836) );
  MUX2_X1 U11281 ( .A(n8837), .B(n8836), .S(n10132), .Z(n8838) );
  AOI21_X1 U11282 ( .B1(n8839), .B2(n8838), .A(n11247), .ZN(n8846) );
  INV_X1 U11283 ( .A(n11377), .ZN(n8934) );
  MUX2_X1 U11284 ( .A(n8841), .B(n8840), .S(n10132), .Z(n8842) );
  NAND2_X1 U11285 ( .A1(n8934), .A2(n8842), .ZN(n8845) );
  AND2_X1 U11286 ( .A1(n8851), .A2(n8843), .ZN(n8844) );
  OAI22_X1 U11287 ( .A1(n8846), .A2(n8845), .B1(n10132), .B2(n8844), .ZN(n8850) );
  AOI21_X1 U11288 ( .B1(n8849), .B2(n8847), .A(n9044), .ZN(n8848) );
  AOI21_X1 U11289 ( .B1(n8850), .B2(n8849), .A(n8848), .ZN(n8856) );
  AND2_X1 U11290 ( .A1(n8853), .A2(n8852), .ZN(n11400) );
  OAI21_X1 U11291 ( .B1(n9044), .B2(n8851), .A(n11400), .ZN(n8855) );
  NAND2_X1 U11292 ( .A1(n8858), .A2(n8857), .ZN(n12382) );
  INV_X1 U11293 ( .A(n12382), .ZN(n12387) );
  MUX2_X1 U11294 ( .A(n8853), .B(n8852), .S(n9044), .Z(n8854) );
  OAI211_X1 U11295 ( .C1(n8856), .C2(n8855), .A(n12387), .B(n8854), .ZN(n8860)
         );
  MUX2_X1 U11296 ( .A(n8858), .B(n8857), .S(n10132), .Z(n8859) );
  AOI21_X1 U11297 ( .B1(n8860), .B2(n8859), .A(n9000), .ZN(n8869) );
  NAND2_X1 U11298 ( .A1(n8865), .A2(n8861), .ZN(n8864) );
  NAND2_X1 U11299 ( .A1(n8866), .A2(n8862), .ZN(n8863) );
  MUX2_X1 U11300 ( .A(n8864), .B(n8863), .S(n9044), .Z(n8868) );
  MUX2_X1 U11301 ( .A(n8866), .B(n8865), .S(n9044), .Z(n8867) );
  OAI21_X1 U11302 ( .B1(n8869), .B2(n8868), .A(n8867), .ZN(n8870) );
  AND3_X1 U11303 ( .A1(n8870), .A2(n12334), .A3(n12348), .ZN(n8882) );
  NAND2_X1 U11304 ( .A1(n8872), .A2(n8871), .ZN(n8873) );
  NAND2_X1 U11305 ( .A1(n8873), .A2(n8876), .ZN(n8874) );
  NAND2_X1 U11306 ( .A1(n8928), .A2(n8874), .ZN(n8879) );
  NAND2_X1 U11307 ( .A1(n12334), .A2(n8875), .ZN(n8877) );
  NAND3_X1 U11308 ( .A1(n8877), .A2(n8929), .A3(n8876), .ZN(n8878) );
  MUX2_X1 U11309 ( .A(n8879), .B(n8878), .S(n9044), .Z(n8881) );
  MUX2_X1 U11310 ( .A(n8928), .B(n8929), .S(n10132), .Z(n8880) );
  OAI21_X1 U11311 ( .B1(n8882), .B2(n8881), .A(n8880), .ZN(n8887) );
  NAND2_X1 U11312 ( .A1(n8889), .A2(n8890), .ZN(n12296) );
  INV_X1 U11313 ( .A(n12296), .ZN(n8886) );
  NAND2_X1 U11314 ( .A1(n12432), .A2(n12295), .ZN(n8884) );
  MUX2_X1 U11315 ( .A(n8884), .B(n8883), .S(n10132), .Z(n8885) );
  OAI211_X1 U11316 ( .C1(n8887), .C2(n12311), .A(n8886), .B(n8885), .ZN(n8892)
         );
  OR2_X1 U11317 ( .A1(n8893), .A2(n8894), .ZN(n12284) );
  INV_X1 U11318 ( .A(n12284), .ZN(n12279) );
  MUX2_X1 U11319 ( .A(n8890), .B(n8889), .S(n9044), .Z(n8891) );
  AND3_X1 U11320 ( .A1(n8892), .A2(n12279), .A3(n8891), .ZN(n8896) );
  MUX2_X1 U11321 ( .A(n8894), .B(n8893), .S(n10132), .Z(n8895) );
  OAI33_X1 U11322 ( .A1(n9044), .A2(n12420), .A3(n11835), .B1(n12263), .B2(
        n8896), .B3(n8895), .ZN(n8902) );
  INV_X1 U11323 ( .A(n8897), .ZN(n8900) );
  AOI211_X1 U11324 ( .C1(n8902), .C2(n12247), .A(n8901), .B(n12239), .ZN(n8907) );
  INV_X1 U11325 ( .A(n8903), .ZN(n8904) );
  MUX2_X1 U11326 ( .A(n8905), .B(n8904), .S(n10132), .Z(n8906) );
  NOR3_X1 U11327 ( .A1(n8907), .A2(n8906), .A3(n12227), .ZN(n8911) );
  MUX2_X1 U11328 ( .A(n8909), .B(n8908), .S(n9044), .Z(n8910) );
  OAI21_X1 U11329 ( .B1(n8911), .B2(n8910), .A(n12217), .ZN(n8913) );
  NAND3_X1 U11330 ( .A1(n12475), .A2(n12201), .A3(n9044), .ZN(n8912) );
  AOI21_X1 U11331 ( .B1(n8913), .B2(n8912), .A(n12199), .ZN(n8918) );
  XNOR2_X1 U11332 ( .A(n8914), .B(n9044), .ZN(n8915) );
  AOI21_X1 U11333 ( .B1(n7384), .B2(n8916), .A(n8915), .ZN(n8917) );
  NAND2_X1 U11334 ( .A1(n8919), .A2(n8920), .ZN(n9017) );
  INV_X1 U11335 ( .A(n9017), .ZN(n8974) );
  INV_X1 U11336 ( .A(n8924), .ZN(n8945) );
  MUX2_X1 U11337 ( .A(n8920), .B(n8919), .S(n9044), .Z(n8921) );
  INV_X1 U11338 ( .A(n8925), .ZN(n8944) );
  INV_X1 U11339 ( .A(n8927), .ZN(n8947) );
  NOR2_X1 U11340 ( .A1(n14917), .A2(n8930), .ZN(n11798) );
  NAND4_X1 U11341 ( .A1(n11798), .A2(n10699), .A3(n10945), .A4(n10348), .ZN(
        n8932) );
  NOR2_X1 U11342 ( .A1(n8932), .A2(n8931), .ZN(n8935) );
  NOR2_X1 U11343 ( .A1(n7404), .A2(n11247), .ZN(n8933) );
  AND4_X1 U11344 ( .A1(n8935), .A2(n8934), .A3(n8933), .A4(n14886), .ZN(n8936)
         );
  NAND4_X1 U11345 ( .A1(n12387), .A2(n11356), .A3(n11400), .A4(n8936), .ZN(
        n8937) );
  NOR2_X1 U11346 ( .A1(n8937), .A2(n9000), .ZN(n8938) );
  NAND4_X1 U11347 ( .A1(n12334), .A2(n12348), .A3(n12359), .A4(n8938), .ZN(
        n8939) );
  OR4_X1 U11348 ( .A1(n12296), .A2(n12311), .A3(n7564), .A4(n8939), .ZN(n8940)
         );
  NOR4_X1 U11349 ( .A1(n12250), .A2(n12263), .A3(n12284), .A4(n8940), .ZN(
        n8941) );
  NAND4_X1 U11350 ( .A1(n7384), .A2(n8942), .A3(n9015), .A4(n8941), .ZN(n8943)
         );
  NOR3_X1 U11351 ( .A1(n9017), .A2(n8943), .A3(n9016), .ZN(n8946) );
  NAND4_X1 U11352 ( .A1(n8947), .A2(n8946), .A3(n8945), .A4(n8944), .ZN(n8948)
         );
  XNOR2_X1 U11353 ( .A(n8948), .B(n12177), .ZN(n8950) );
  NOR2_X1 U11354 ( .A1(n10628), .A2(n10169), .ZN(n9149) );
  INV_X1 U11355 ( .A(n9149), .ZN(n8949) );
  NAND2_X1 U11356 ( .A1(n6484), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8954) );
  INV_X1 U11357 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8953) );
  NOR2_X1 U11358 ( .A1(n10131), .A2(P3_U3151), .ZN(n8970) );
  INV_X1 U11359 ( .A(n10804), .ZN(n8967) );
  NAND2_X1 U11360 ( .A1(n8960), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8961) );
  INV_X1 U11361 ( .A(n11201), .ZN(n8965) );
  NAND2_X1 U11362 ( .A1(n8956), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8962) );
  MUX2_X1 U11363 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8962), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n8963) );
  NAND2_X1 U11364 ( .A1(n8963), .A2(n8960), .ZN(n11016) );
  INV_X1 U11365 ( .A(n11016), .ZN(n8964) );
  AND2_X1 U11366 ( .A1(n8965), .A2(n8964), .ZN(n8966) );
  NAND2_X1 U11367 ( .A1(n8967), .A2(n8966), .ZN(n9517) );
  NOR2_X1 U11368 ( .A1(n9060), .A2(n9044), .ZN(n11797) );
  NAND2_X1 U11369 ( .A1(n9175), .A2(n11797), .ZN(n9178) );
  NOR3_X1 U11370 ( .A1(n9178), .A2(n12168), .A3(n12531), .ZN(n8972) );
  INV_X1 U11371 ( .A(n8970), .ZN(n10511) );
  OAI21_X1 U11372 ( .B1(n10511), .B2(n10198), .A(P3_B_REG_SCAN_IN), .ZN(n8971)
         );
  OR2_X1 U11373 ( .A1(n8972), .A2(n8971), .ZN(n8973) );
  XNOR2_X1 U11374 ( .A(n8975), .B(n8974), .ZN(n12195) );
  NAND2_X1 U11375 ( .A1(n12177), .A2(n10196), .ZN(n8978) );
  NAND2_X1 U11376 ( .A1(n10196), .A2(n10169), .ZN(n8976) );
  XNOR2_X1 U11377 ( .A(n10198), .B(n8976), .ZN(n8977) );
  NAND2_X1 U11378 ( .A1(n8978), .A2(n8977), .ZN(n9174) );
  NAND3_X1 U11379 ( .A1(n9174), .A2(n8979), .A3(n14915), .ZN(n8981) );
  AND2_X1 U11380 ( .A1(n10198), .A2(n9046), .ZN(n8980) );
  NAND2_X1 U11381 ( .A1(n12177), .A2(n8980), .ZN(n9045) );
  NAND2_X1 U11382 ( .A1(n8981), .A2(n9045), .ZN(n14906) );
  NAND2_X1 U11383 ( .A1(n14918), .A2(n10124), .ZN(n14922) );
  NAND2_X1 U11384 ( .A1(n8982), .A2(n14922), .ZN(n8984) );
  NAND2_X1 U11385 ( .A1(n9066), .A2(n14916), .ZN(n8983) );
  NAND2_X1 U11386 ( .A1(n8984), .A2(n8983), .ZN(n14900) );
  NAND2_X1 U11387 ( .A1(n10708), .A2(n14910), .ZN(n10706) );
  AND2_X1 U11388 ( .A1(n10705), .A2(n10706), .ZN(n8985) );
  NAND2_X1 U11389 ( .A1(n14899), .A2(n8985), .ZN(n10704) );
  NAND2_X1 U11390 ( .A1(n11995), .A2(n10703), .ZN(n8986) );
  NAND2_X1 U11391 ( .A1(n10704), .A2(n8986), .ZN(n10647) );
  NAND2_X1 U11392 ( .A1(n11994), .A2(n10695), .ZN(n8987) );
  NAND2_X1 U11393 ( .A1(n10948), .A2(n10809), .ZN(n10951) );
  AND2_X1 U11394 ( .A1(n10950), .A2(n10951), .ZN(n8989) );
  NAND2_X1 U11395 ( .A1(n10952), .A2(n8989), .ZN(n10949) );
  NAND2_X1 U11396 ( .A1(n11993), .A2(n10958), .ZN(n8990) );
  INV_X1 U11397 ( .A(n11171), .ZN(n14894) );
  NAND2_X1 U11398 ( .A1(n11155), .A2(n14894), .ZN(n8991) );
  INV_X1 U11399 ( .A(n8991), .ZN(n8993) );
  NAND2_X1 U11400 ( .A1(n14888), .A2(n14961), .ZN(n14883) );
  AND2_X1 U11401 ( .A1(n7575), .A2(n14883), .ZN(n8992) );
  NAND2_X1 U11402 ( .A1(n11991), .A2(n11370), .ZN(n8994) );
  NAND2_X1 U11403 ( .A1(n11866), .A2(n11381), .ZN(n8995) );
  NAND2_X1 U11404 ( .A1(n11376), .A2(n8995), .ZN(n11352) );
  NAND2_X1 U11405 ( .A1(n11990), .A2(n14167), .ZN(n8996) );
  OR2_X1 U11406 ( .A1(n14162), .A2(n11920), .ZN(n8997) );
  NAND2_X1 U11407 ( .A1(n12381), .A2(n12382), .ZN(n8999) );
  NAND2_X1 U11408 ( .A1(n12388), .A2(n11989), .ZN(n8998) );
  NAND2_X1 U11409 ( .A1(n8999), .A2(n8998), .ZN(n12367) );
  NAND2_X1 U11410 ( .A1(n12367), .A2(n9000), .ZN(n9002) );
  INV_X1 U11411 ( .A(n12385), .ZN(n11988) );
  NAND2_X1 U11412 ( .A1(n12452), .A2(n11988), .ZN(n9001) );
  NAND2_X1 U11413 ( .A1(n9002), .A2(n9001), .ZN(n12355) );
  NAND2_X1 U11414 ( .A1(n12361), .A2(n12345), .ZN(n9003) );
  INV_X1 U11415 ( .A(n12330), .ZN(n9006) );
  OR2_X1 U11416 ( .A1(n11954), .A2(n12344), .ZN(n9008) );
  INV_X1 U11417 ( .A(n12305), .ZN(n12332) );
  NAND2_X1 U11418 ( .A1(n12304), .A2(n12311), .ZN(n9010) );
  NAND2_X1 U11419 ( .A1(n12432), .A2(n12319), .ZN(n9009) );
  AND2_X1 U11420 ( .A1(n12298), .A2(n12306), .ZN(n9012) );
  OR2_X1 U11421 ( .A1(n12298), .A2(n12306), .ZN(n9011) );
  OAI21_X1 U11422 ( .B1(n12292), .B2(n9012), .A(n9011), .ZN(n12280) );
  INV_X1 U11423 ( .A(n12280), .ZN(n9013) );
  NAND2_X1 U11424 ( .A1(n12235), .A2(n12239), .ZN(n12234) );
  INV_X1 U11425 ( .A(n12413), .ZN(n11883) );
  OAI21_X1 U11426 ( .B1(n12214), .B2(n12471), .A(n12198), .ZN(n9018) );
  XNOR2_X1 U11427 ( .A(n9018), .B(n9017), .ZN(n9024) );
  NAND2_X1 U11428 ( .A1(n9048), .A2(n10198), .ZN(n9020) );
  OR2_X1 U11429 ( .A1(n12531), .A2(n14738), .ZN(n10139) );
  NAND2_X1 U11430 ( .A1(n10139), .A2(n10134), .ZN(n9165) );
  INV_X1 U11431 ( .A(n9165), .ZN(n9162) );
  INV_X1 U11432 ( .A(n12214), .ZN(n11985) );
  INV_X1 U11433 ( .A(P3_B_REG_SCAN_IN), .ZN(n9021) );
  NOR2_X1 U11434 ( .A1(n12531), .A2(n9021), .ZN(n9022) );
  NOR2_X1 U11435 ( .A1(n14901), .A2(n9022), .ZN(n12182) );
  AOI22_X1 U11436 ( .A1(n14919), .A2(n11985), .B1(n11983), .B2(n12182), .ZN(
        n9023) );
  INV_X1 U11437 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n9026) );
  NAND2_X1 U11438 ( .A1(n11424), .A2(n9026), .ZN(n9028) );
  NAND2_X1 U11439 ( .A1(n10804), .A2(n11201), .ZN(n9027) );
  INV_X1 U11440 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U11441 ( .A1(n11424), .A2(n9029), .ZN(n9031) );
  NAND2_X1 U11442 ( .A1(n11201), .A2(n11016), .ZN(n9030) );
  XNOR2_X1 U11443 ( .A(n9147), .B(n12512), .ZN(n9043) );
  NOR2_X1 U11444 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n9035) );
  NOR4_X1 U11445 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9034) );
  NOR4_X1 U11446 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n9033) );
  NOR4_X1 U11447 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n9032) );
  NAND4_X1 U11448 ( .A1(n9035), .A2(n9034), .A3(n9033), .A4(n9032), .ZN(n9041)
         );
  NOR4_X1 U11449 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9039) );
  NOR4_X1 U11450 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9038) );
  NOR4_X1 U11451 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9037) );
  NOR4_X1 U11452 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9036) );
  NAND4_X1 U11453 ( .A1(n9039), .A2(n9038), .A3(n9037), .A4(n9036), .ZN(n9040)
         );
  OAI21_X1 U11454 ( .B1(n9041), .B2(n9040), .A(n11424), .ZN(n9146) );
  AND2_X1 U11455 ( .A1(n9146), .A2(n9175), .ZN(n9042) );
  NAND2_X1 U11456 ( .A1(n9060), .A2(n10132), .ZN(n9154) );
  NAND2_X1 U11457 ( .A1(n9045), .A2(n9044), .ZN(n10622) );
  AND2_X1 U11458 ( .A1(n9154), .A2(n10622), .ZN(n10624) );
  OAI22_X1 U11459 ( .A1(n9048), .A2(n9047), .B1(n9046), .B2(n14915), .ZN(n9049) );
  AOI21_X1 U11460 ( .B1(n9049), .B2(n9060), .A(n10132), .ZN(n9051) );
  INV_X1 U11461 ( .A(n12512), .ZN(n9050) );
  MUX2_X1 U11462 ( .A(n10624), .B(n9051), .S(n9050), .Z(n9052) );
  INV_X1 U11463 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U11464 ( .A1(n9057), .A2(n9056), .ZN(P3_U3488) );
  NAND2_X2 U11465 ( .A1(n12514), .A2(n9149), .ZN(n9062) );
  NAND2_X1 U11466 ( .A1(n10628), .A2(n10169), .ZN(n9059) );
  XNOR2_X1 U11467 ( .A(n9063), .B(n10347), .ZN(n11815) );
  NOR2_X1 U11468 ( .A1(n11815), .A2(n12201), .ZN(n11811) );
  AOI21_X1 U11469 ( .B1(n11815), .B2(n12201), .A(n11811), .ZN(n9145) );
  XNOR2_X1 U11470 ( .A(n6435), .B(n10695), .ZN(n9077) );
  INV_X1 U11471 ( .A(n9075), .ZN(n9076) );
  NAND2_X1 U11472 ( .A1(n9064), .A2(n6452), .ZN(n9065) );
  NAND2_X1 U11473 ( .A1(n14922), .A2(n9065), .ZN(n9069) );
  NOR2_X1 U11474 ( .A1(n9069), .A2(n10351), .ZN(n10349) );
  INV_X1 U11475 ( .A(n9070), .ZN(n9071) );
  INV_X1 U11476 ( .A(n9073), .ZN(n9074) );
  XNOR2_X1 U11477 ( .A(n9075), .B(n14902), .ZN(n10639) );
  XNOR2_X1 U11478 ( .A(n9077), .B(n11994), .ZN(n10690) );
  XNOR2_X1 U11479 ( .A(n6435), .B(n10630), .ZN(n9078) );
  XNOR2_X1 U11480 ( .A(n9078), .B(n10832), .ZN(n10806) );
  XNOR2_X1 U11481 ( .A(n6435), .B(n9079), .ZN(n9080) );
  XNOR2_X1 U11482 ( .A(n9080), .B(n10920), .ZN(n10829) );
  NAND2_X1 U11483 ( .A1(n10830), .A2(n10829), .ZN(n10828) );
  NAND2_X1 U11484 ( .A1(n9080), .A2(n11993), .ZN(n9081) );
  NAND2_X1 U11485 ( .A1(n10828), .A2(n9081), .ZN(n10980) );
  XNOR2_X1 U11486 ( .A(n14881), .B(n10347), .ZN(n10979) );
  NAND2_X1 U11487 ( .A1(n10980), .A2(n10979), .ZN(n10978) );
  INV_X1 U11488 ( .A(n10979), .ZN(n9082) );
  NAND2_X1 U11489 ( .A1(n9082), .A2(n14888), .ZN(n9083) );
  XNOR2_X1 U11490 ( .A(n6435), .B(n14894), .ZN(n9084) );
  XNOR2_X1 U11491 ( .A(n9084), .B(n11155), .ZN(n11166) );
  NAND2_X1 U11492 ( .A1(n9084), .A2(n11992), .ZN(n9085) );
  XNOR2_X1 U11493 ( .A(n6435), .B(n11306), .ZN(n9087) );
  XNOR2_X1 U11494 ( .A(n9087), .B(n14887), .ZN(n11301) );
  INV_X1 U11495 ( .A(n11301), .ZN(n9086) );
  INV_X1 U11496 ( .A(n9087), .ZN(n9088) );
  INV_X1 U11497 ( .A(n14887), .ZN(n11169) );
  NAND2_X1 U11498 ( .A1(n9088), .A2(n11169), .ZN(n9089) );
  XNOR2_X1 U11499 ( .A(n6435), .B(n11370), .ZN(n9090) );
  XNOR2_X1 U11500 ( .A(n9090), .B(n11303), .ZN(n11363) );
  INV_X1 U11501 ( .A(n9090), .ZN(n9091) );
  NAND2_X1 U11502 ( .A1(n9091), .A2(n11991), .ZN(n9092) );
  XNOR2_X1 U11503 ( .A(n6435), .B(n11381), .ZN(n9095) );
  XNOR2_X1 U11504 ( .A(n11868), .B(n6435), .ZN(n11862) );
  NAND2_X1 U11505 ( .A1(n11862), .A2(n11990), .ZN(n9094) );
  OAI21_X1 U11506 ( .B1(n11945), .B2(n9095), .A(n9094), .ZN(n9093) );
  INV_X1 U11507 ( .A(n11862), .ZN(n9098) );
  INV_X1 U11508 ( .A(n9094), .ZN(n9096) );
  INV_X1 U11509 ( .A(n9095), .ZN(n11860) );
  NOR3_X1 U11510 ( .A1(n9096), .A2(n11860), .A3(n11866), .ZN(n9097) );
  AOI21_X1 U11511 ( .B1(n11937), .B2(n9098), .A(n9097), .ZN(n9099) );
  XNOR2_X1 U11512 ( .A(n14162), .B(n10347), .ZN(n11921) );
  NOR2_X1 U11513 ( .A1(n11921), .A2(n11920), .ZN(n9101) );
  INV_X1 U11514 ( .A(n11921), .ZN(n9100) );
  XNOR2_X1 U11515 ( .A(n12388), .B(n6435), .ZN(n9102) );
  XNOR2_X1 U11516 ( .A(n9102), .B(n11989), .ZN(n11826) );
  NAND2_X1 U11517 ( .A1(n11827), .A2(n11826), .ZN(n9105) );
  INV_X1 U11518 ( .A(n9102), .ZN(n9103) );
  NAND2_X1 U11519 ( .A1(n9103), .A2(n11989), .ZN(n9104) );
  XNOR2_X1 U11520 ( .A(n12452), .B(n6435), .ZN(n11970) );
  NOR2_X1 U11521 ( .A1(n11970), .A2(n12385), .ZN(n9107) );
  NAND2_X1 U11522 ( .A1(n11970), .A2(n12385), .ZN(n9106) );
  XNOR2_X1 U11523 ( .A(n12361), .B(n10347), .ZN(n11884) );
  NOR2_X1 U11524 ( .A1(n11884), .A2(n12345), .ZN(n9109) );
  INV_X1 U11525 ( .A(n11884), .ZN(n9108) );
  XNOR2_X1 U11526 ( .A(n12444), .B(n6435), .ZN(n9110) );
  XNOR2_X1 U11527 ( .A(n9110), .B(n11952), .ZN(n11892) );
  INV_X1 U11528 ( .A(n9110), .ZN(n9111) );
  NAND2_X1 U11529 ( .A1(n9111), .A2(n11952), .ZN(n9112) );
  XNOR2_X1 U11530 ( .A(n11954), .B(n6435), .ZN(n9113) );
  XNOR2_X1 U11531 ( .A(n9113), .B(n12344), .ZN(n11951) );
  INV_X1 U11532 ( .A(n9113), .ZN(n9114) );
  NAND2_X1 U11533 ( .A1(n9114), .A2(n12344), .ZN(n9115) );
  XNOR2_X1 U11534 ( .A(n12496), .B(n6435), .ZN(n9116) );
  XNOR2_X1 U11535 ( .A(n9116), .B(n12332), .ZN(n11841) );
  NAND2_X1 U11536 ( .A1(n9116), .A2(n12305), .ZN(n11909) );
  XNOR2_X1 U11537 ( .A(n12432), .B(n6435), .ZN(n9121) );
  INV_X1 U11538 ( .A(n9121), .ZN(n9117) );
  NAND2_X1 U11539 ( .A1(n9117), .A2(n12319), .ZN(n9120) );
  AND2_X1 U11540 ( .A1(n11909), .A2(n9120), .ZN(n11848) );
  XNOR2_X1 U11541 ( .A(n12298), .B(n6435), .ZN(n9118) );
  NAND2_X1 U11542 ( .A1(n9118), .A2(n12283), .ZN(n9124) );
  OAI21_X1 U11543 ( .B1(n9118), .B2(n12283), .A(n9124), .ZN(n11854) );
  INV_X1 U11544 ( .A(n11854), .ZN(n9119) );
  AND2_X1 U11545 ( .A1(n11848), .A2(n9119), .ZN(n9123) );
  INV_X1 U11546 ( .A(n9120), .ZN(n9122) );
  XNOR2_X1 U11547 ( .A(n9121), .B(n12319), .ZN(n11911) );
  XNOR2_X1 U11548 ( .A(n12286), .B(n6435), .ZN(n9126) );
  INV_X1 U11549 ( .A(n9126), .ZN(n9127) );
  XNOR2_X1 U11550 ( .A(n12276), .B(n6435), .ZN(n9129) );
  INV_X1 U11551 ( .A(n9128), .ZN(n9131) );
  INV_X1 U11552 ( .A(n9129), .ZN(n9130) );
  XNOR2_X1 U11553 ( .A(n9132), .B(n6435), .ZN(n9133) );
  NAND2_X1 U11554 ( .A1(n9133), .A2(n12266), .ZN(n11873) );
  INV_X1 U11555 ( .A(n9133), .ZN(n9134) );
  NAND2_X1 U11556 ( .A1(n9134), .A2(n6590), .ZN(n9135) );
  AND2_X1 U11557 ( .A1(n12282), .A2(n11900), .ZN(n9137) );
  INV_X1 U11558 ( .A(n11900), .ZN(n9136) );
  XNOR2_X1 U11559 ( .A(n12413), .B(n6452), .ZN(n9138) );
  NAND2_X1 U11560 ( .A1(n9138), .A2(n12249), .ZN(n9142) );
  INV_X1 U11561 ( .A(n9138), .ZN(n9139) );
  INV_X1 U11562 ( .A(n12249), .ZN(n11986) );
  NAND2_X1 U11563 ( .A1(n9139), .A2(n11986), .ZN(n9140) );
  XNOR2_X1 U11564 ( .A(n11959), .B(n10347), .ZN(n9143) );
  NOR2_X1 U11565 ( .A1(n9143), .A2(n12236), .ZN(n9144) );
  AOI21_X1 U11566 ( .B1(n9143), .B2(n12236), .A(n9144), .ZN(n11962) );
  NAND3_X1 U11567 ( .A1(n12514), .A2(n12512), .A3(n9146), .ZN(n9179) );
  INV_X1 U11568 ( .A(n9175), .ZN(n10130) );
  NOR2_X1 U11569 ( .A1(n9179), .A2(n10130), .ZN(n9173) );
  NAND3_X1 U11570 ( .A1(n9173), .A2(n9174), .A3(n14915), .ZN(n9152) );
  NAND2_X1 U11571 ( .A1(n9147), .A2(n9146), .ZN(n9148) );
  OR2_X1 U11572 ( .A1(n12512), .A2(n9148), .ZN(n9177) );
  INV_X1 U11573 ( .A(n9177), .ZN(n9164) );
  NAND2_X1 U11574 ( .A1(n9149), .A2(n10198), .ZN(n9150) );
  NAND3_X1 U11575 ( .A1(n9164), .A2(n9175), .A3(n6583), .ZN(n9151) );
  AND2_X1 U11576 ( .A1(n14911), .A2(n14960), .ZN(n9153) );
  AND2_X2 U11577 ( .A1(n9175), .A2(n9153), .ZN(n14929) );
  AOI21_X2 U11578 ( .B1(n9173), .B2(n14960), .A(n14929), .ZN(n11968) );
  NAND2_X1 U11579 ( .A1(n9179), .A2(n9174), .ZN(n9157) );
  AND2_X1 U11580 ( .A1(n9517), .A2(n10131), .ZN(n9156) );
  NAND2_X1 U11581 ( .A1(n9177), .A2(n6583), .ZN(n9155) );
  NAND4_X1 U11582 ( .A1(n9157), .A2(n9156), .A3(n9155), .A4(n9154), .ZN(n9158)
         );
  NAND2_X1 U11583 ( .A1(n9158), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9161) );
  INV_X1 U11584 ( .A(n9178), .ZN(n9159) );
  NAND2_X1 U11585 ( .A1(n9177), .A2(n9159), .ZN(n9160) );
  NOR2_X1 U11586 ( .A1(n9178), .A2(n9162), .ZN(n9163) );
  NAND2_X1 U11587 ( .A1(n9164), .A2(n9163), .ZN(n11977) );
  OR2_X1 U11588 ( .A1(n9178), .A2(n9165), .ZN(n9166) );
  AOI22_X1 U11589 ( .A1(n12236), .A2(n11940), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n9167) );
  OAI21_X1 U11590 ( .B1(n12214), .B2(n11977), .A(n9167), .ZN(n9168) );
  AOI21_X1 U11591 ( .B1(n12219), .B2(n11972), .A(n9168), .ZN(n9169) );
  INV_X1 U11592 ( .A(n9170), .ZN(n9171) );
  NAND2_X1 U11593 ( .A1(n9172), .A2(n9171), .ZN(P3_U3154) );
  NAND2_X1 U11594 ( .A1(n9173), .A2(n6583), .ZN(n9182) );
  NAND2_X1 U11595 ( .A1(n9175), .A2(n9174), .ZN(n9176) );
  OAI22_X1 U11596 ( .A1(n9179), .A2(n9178), .B1(n9177), .B2(n9176), .ZN(n9180)
         );
  INV_X1 U11597 ( .A(n9180), .ZN(n9181) );
  NAND2_X1 U11598 ( .A1(n8787), .A2(n9184), .ZN(n9185) );
  NAND2_X1 U11599 ( .A1(n9187), .A2(n9957), .ZN(n9364) );
  NAND2_X1 U11600 ( .A1(n9188), .A2(n9364), .ZN(n9192) );
  NAND2_X1 U11601 ( .A1(n12746), .A2(n9957), .ZN(n9190) );
  INV_X1 U11602 ( .A(n9343), .ZN(n9189) );
  NAND3_X1 U11603 ( .A1(n9190), .A2(n9186), .A3(n9189), .ZN(n9191) );
  NAND2_X1 U11604 ( .A1(n10021), .A2(n9342), .ZN(n9193) );
  NAND2_X1 U11605 ( .A1(n9194), .A2(n9193), .ZN(n9196) );
  AOI22_X1 U11606 ( .A1(n12745), .A2(n9342), .B1(n6445), .B2(n10021), .ZN(
        n9195) );
  NAND2_X1 U11607 ( .A1(n12744), .A2(n9342), .ZN(n9198) );
  NAND2_X1 U11608 ( .A1(n12684), .A2(n6445), .ZN(n9197) );
  NAND2_X1 U11609 ( .A1(n9198), .A2(n9197), .ZN(n9200) );
  INV_X1 U11610 ( .A(n9200), .ZN(n9202) );
  AOI22_X1 U11611 ( .A1(n12744), .A2(n6445), .B1(n12684), .B2(n9342), .ZN(
        n9199) );
  AOI22_X1 U11612 ( .A1(n12743), .A2(n6445), .B1(n14651), .B2(n9342), .ZN(
        n9204) );
  INV_X1 U11613 ( .A(n9204), .ZN(n9207) );
  OAI22_X1 U11614 ( .A1(n10420), .A2(n6445), .B1(n10383), .B2(n9342), .ZN(
        n9203) );
  OAI22_X1 U11615 ( .A1(n10431), .A2(n9342), .B1(n10090), .B2(n6445), .ZN(
        n9210) );
  INV_X1 U11616 ( .A(n9210), .ZN(n9211) );
  AOI22_X1 U11617 ( .A1(n10471), .A2(n9342), .B1(n9213), .B2(n12741), .ZN(
        n9215) );
  OAI22_X1 U11618 ( .A1(n14670), .A2(n9342), .B1(n10438), .B2(n6445), .ZN(
        n9214) );
  INV_X1 U11619 ( .A(n9217), .ZN(n9218) );
  OAI22_X1 U11620 ( .A1(n14684), .A2(n9213), .B1(n10591), .B2(n9342), .ZN(
        n9219) );
  INV_X1 U11621 ( .A(n9219), .ZN(n9223) );
  NAND2_X1 U11622 ( .A1(n9220), .A2(n9219), .ZN(n9222) );
  OAI22_X1 U11623 ( .A1(n14684), .A2(n9342), .B1(n10591), .B2(n9213), .ZN(
        n9221) );
  OAI22_X1 U11624 ( .A1(n14692), .A2(n9342), .B1(n10741), .B2(n6445), .ZN(
        n9225) );
  OAI22_X1 U11625 ( .A1(n14692), .A2(n9213), .B1(n10741), .B2(n9342), .ZN(
        n9227) );
  INV_X1 U11626 ( .A(n9225), .ZN(n9226) );
  AOI22_X1 U11627 ( .A1(n10793), .A2(n9342), .B1(n9213), .B2(n12736), .ZN(
        n9228) );
  OAI22_X1 U11628 ( .A1(n6802), .A2(n9342), .B1(n10787), .B2(n9213), .ZN(n9230) );
  AOI22_X1 U11629 ( .A1(n10933), .A2(n9213), .B1(n12735), .B2(n9342), .ZN(
        n9233) );
  AOI22_X1 U11630 ( .A1(n10933), .A2(n9342), .B1(n9213), .B2(n12735), .ZN(
        n9231) );
  INV_X1 U11631 ( .A(n9231), .ZN(n9232) );
  NAND2_X1 U11632 ( .A1(n9234), .A2(n9233), .ZN(n9235) );
  OAI22_X1 U11633 ( .A1(n14186), .A2(n9342), .B1(n11317), .B2(n9213), .ZN(
        n9240) );
  OAI22_X1 U11634 ( .A1(n14186), .A2(n6445), .B1(n11317), .B2(n9342), .ZN(
        n9241) );
  OAI22_X1 U11635 ( .A1(n11314), .A2(n6445), .B1(n11418), .B2(n9342), .ZN(
        n9244) );
  INV_X1 U11636 ( .A(n9244), .ZN(n9243) );
  OAI22_X1 U11637 ( .A1(n11314), .A2(n9342), .B1(n11418), .B2(n9213), .ZN(
        n9242) );
  INV_X1 U11638 ( .A(n9247), .ZN(n9245) );
  NAND2_X1 U11639 ( .A1(n9246), .A2(n9245), .ZN(n9250) );
  OAI22_X1 U11640 ( .A1(n14180), .A2(n6445), .B1(n11315), .B2(n9342), .ZN(
        n9249) );
  INV_X1 U11641 ( .A(n9246), .ZN(n9248) );
  AOI22_X1 U11642 ( .A1(n13167), .A2(n9342), .B1(n6445), .B2(n12730), .ZN(
        n9253) );
  AOI22_X1 U11643 ( .A1(n13167), .A2(n6445), .B1(n12730), .B2(n9342), .ZN(
        n9251) );
  INV_X1 U11644 ( .A(n9251), .ZN(n9252) );
  OAI22_X1 U11645 ( .A1(n13074), .A2(n9342), .B1(n12648), .B2(n9213), .ZN(
        n9256) );
  OAI22_X1 U11646 ( .A1(n13074), .A2(n6445), .B1(n12648), .B2(n9342), .ZN(
        n9255) );
  INV_X1 U11647 ( .A(n9256), .ZN(n9257) );
  OAI22_X1 U11648 ( .A1(n13045), .A2(n6445), .B1(n13058), .B2(n9342), .ZN(
        n9259) );
  NAND2_X1 U11649 ( .A1(n9258), .A2(n9259), .ZN(n9263) );
  OAI22_X1 U11650 ( .A1(n13045), .A2(n9342), .B1(n13058), .B2(n6445), .ZN(
        n9262) );
  INV_X1 U11651 ( .A(n9259), .ZN(n9260) );
  OAI22_X1 U11652 ( .A1(n13036), .A2(n9342), .B1(n13014), .B2(n6445), .ZN(
        n9264) );
  OAI22_X1 U11653 ( .A1(n13036), .A2(n6445), .B1(n13014), .B2(n9342), .ZN(
        n9267) );
  OAI22_X1 U11654 ( .A1(n13022), .A2(n6445), .B1(n12697), .B2(n9342), .ZN(
        n9271) );
  INV_X1 U11655 ( .A(n9271), .ZN(n9270) );
  OAI22_X1 U11656 ( .A1(n13022), .A2(n9342), .B1(n12697), .B2(n6445), .ZN(
        n9269) );
  AOI22_X1 U11657 ( .A1(n13142), .A2(n9213), .B1(n12976), .B2(n9342), .ZN(
        n9274) );
  INV_X1 U11658 ( .A(n13142), .ZN(n9273) );
  OAI22_X1 U11659 ( .A1(n9273), .A2(n6445), .B1(n13015), .B2(n9342), .ZN(n9277) );
  AOI22_X1 U11660 ( .A1(n13134), .A2(n9342), .B1(n6445), .B2(n13005), .ZN(
        n9281) );
  INV_X1 U11661 ( .A(n13005), .ZN(n12674) );
  OAI22_X1 U11662 ( .A1(n9279), .A2(n9342), .B1(n12674), .B2(n6445), .ZN(n9280) );
  NAND2_X1 U11663 ( .A1(n9282), .A2(n9281), .ZN(n9283) );
  OAI22_X1 U11664 ( .A1(n13129), .A2(n9342), .B1(n12621), .B2(n6445), .ZN(
        n9286) );
  AOI22_X1 U11665 ( .A1(n12679), .A2(n9342), .B1(n6445), .B2(n12975), .ZN(
        n9285) );
  OAI22_X1 U11666 ( .A1(n12954), .A2(n6445), .B1(n12675), .B2(n9342), .ZN(
        n9288) );
  AOI22_X1 U11667 ( .A1(n13124), .A2(n6445), .B1(n12931), .B2(n9342), .ZN(
        n9287) );
  OAI22_X1 U11668 ( .A1(n12939), .A2(n9342), .B1(n12631), .B2(n6445), .ZN(
        n9291) );
  AOI22_X1 U11669 ( .A1(n13118), .A2(n9342), .B1(n6445), .B2(n12917), .ZN(
        n9290) );
  AOI22_X1 U11670 ( .A1(n13113), .A2(n6445), .B1(n12932), .B2(n9342), .ZN(
        n9322) );
  OAI22_X1 U11671 ( .A1(n12923), .A2(n6445), .B1(n12657), .B2(n9342), .ZN(
        n9321) );
  OR2_X1 U11672 ( .A1(n9322), .A2(n9321), .ZN(n9292) );
  NAND2_X1 U11673 ( .A1(n9294), .A2(n9293), .ZN(n9297) );
  NAND2_X1 U11674 ( .A1(n9295), .A2(n12523), .ZN(n9296) );
  NAND2_X1 U11675 ( .A1(n9297), .A2(n9296), .ZN(n9334) );
  MUX2_X1 U11676 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9657), .Z(n9298) );
  NAND2_X1 U11677 ( .A1(n9298), .A2(SI_30_), .ZN(n9299) );
  OAI21_X1 U11678 ( .B1(n9298), .B2(SI_30_), .A(n9299), .ZN(n9333) );
  MUX2_X1 U11679 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9657), .Z(n9300) );
  XNOR2_X1 U11680 ( .A(n9300), .B(SI_31_), .ZN(n9301) );
  NAND2_X1 U11681 ( .A1(n13187), .A2(n7682), .ZN(n9304) );
  NAND2_X1 U11682 ( .A1(n9338), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9303) );
  INV_X1 U11683 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9309) );
  NAND2_X1 U11684 ( .A1(n9305), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9308) );
  NAND2_X1 U11685 ( .A1(n9306), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9307) );
  OAI211_X1 U11686 ( .C1(n7786), .C2(n9309), .A(n9308), .B(n9307), .ZN(n12847)
         );
  XNOR2_X1 U11687 ( .A(n12848), .B(n12847), .ZN(n9381) );
  AND2_X1 U11688 ( .A1(n12869), .A2(n9342), .ZN(n9310) );
  AOI21_X1 U11689 ( .B1(n12858), .B2(n6445), .A(n9310), .ZN(n9346) );
  NAND2_X1 U11690 ( .A1(n12858), .A2(n9342), .ZN(n9312) );
  NAND2_X1 U11691 ( .A1(n12869), .A2(n6445), .ZN(n9311) );
  NAND2_X1 U11692 ( .A1(n9312), .A2(n9311), .ZN(n9345) );
  AND2_X1 U11693 ( .A1(n12887), .A2(n9342), .ZN(n9313) );
  AOI21_X1 U11694 ( .B1(n13096), .B2(n6445), .A(n9313), .ZN(n9332) );
  NAND2_X1 U11695 ( .A1(n13096), .A2(n9342), .ZN(n9315) );
  NAND2_X1 U11696 ( .A1(n12887), .A2(n9213), .ZN(n9314) );
  NAND2_X1 U11697 ( .A1(n9315), .A2(n9314), .ZN(n9331) );
  AOI22_X1 U11698 ( .A1(n9346), .A2(n9345), .B1(n9332), .B2(n9331), .ZN(n9316)
         );
  AND2_X1 U11699 ( .A1(n12727), .A2(n9342), .ZN(n9317) );
  AOI21_X1 U11700 ( .B1(n13103), .B2(n9213), .A(n9317), .ZN(n9330) );
  NAND2_X1 U11701 ( .A1(n13103), .A2(n9342), .ZN(n9319) );
  NAND2_X1 U11702 ( .A1(n12727), .A2(n9213), .ZN(n9318) );
  NAND2_X1 U11703 ( .A1(n9319), .A2(n9318), .ZN(n9329) );
  NAND2_X1 U11704 ( .A1(n9330), .A2(n9329), .ZN(n9320) );
  OAI22_X1 U11705 ( .A1(n12909), .A2(n6445), .B1(n12629), .B2(n9342), .ZN(
        n9324) );
  AOI22_X1 U11706 ( .A1(n13108), .A2(n6445), .B1(n12918), .B2(n9342), .ZN(
        n9325) );
  AOI22_X1 U11707 ( .A1(n9324), .A2(n9325), .B1(n9322), .B2(n9321), .ZN(n9323)
         );
  INV_X1 U11708 ( .A(n9324), .ZN(n9327) );
  INV_X1 U11709 ( .A(n9325), .ZN(n9326) );
  OAI22_X1 U11710 ( .A1(n9332), .A2(n9331), .B1(n9330), .B2(n9329), .ZN(n9348)
         );
  NAND2_X1 U11711 ( .A1(n9334), .A2(n9333), .ZN(n9335) );
  OR2_X1 U11712 ( .A1(n13981), .A2(n9337), .ZN(n9340) );
  NAND2_X1 U11713 ( .A1(n9338), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9339) );
  OAI22_X1 U11714 ( .A1(n13094), .A2(n6445), .B1(n9341), .B2(n9342), .ZN(n9353) );
  INV_X1 U11715 ( .A(n9341), .ZN(n12726) );
  NAND2_X1 U11716 ( .A1(n12847), .A2(n9342), .ZN(n9354) );
  OAI211_X1 U11717 ( .C1(n10519), .C2(n9343), .A(n9354), .B(n8193), .ZN(n9344)
         );
  AOI22_X1 U11718 ( .A1(n12856), .A2(n9213), .B1(n12726), .B2(n9344), .ZN(
        n9352) );
  OAI22_X1 U11719 ( .A1(n9353), .A2(n9352), .B1(n9346), .B2(n9345), .ZN(n9347)
         );
  NAND2_X1 U11720 ( .A1(n9353), .A2(n9352), .ZN(n9359) );
  AND2_X1 U11721 ( .A1(n12847), .A2(n6445), .ZN(n9357) );
  INV_X1 U11722 ( .A(n9354), .ZN(n9355) );
  NOR2_X1 U11723 ( .A1(n9355), .A2(n6445), .ZN(n9356) );
  MUX2_X1 U11724 ( .A(n9357), .B(n9356), .S(n12848), .Z(n9358) );
  INV_X1 U11725 ( .A(n9387), .ZN(n9385) );
  XNOR2_X1 U11726 ( .A(n12856), .B(n12726), .ZN(n9379) );
  NAND2_X1 U11727 ( .A1(n9361), .A2(n9360), .ZN(n12911) );
  NAND2_X1 U11728 ( .A1(n9363), .A2(n9362), .ZN(n12946) );
  XNOR2_X1 U11729 ( .A(n13148), .B(n12697), .ZN(n13011) );
  NAND2_X1 U11730 ( .A1(n9364), .A2(n9883), .ZN(n14638) );
  NAND4_X1 U11731 ( .A1(n9365), .A2(n10519), .A3(n9886), .A4(n14638), .ZN(
        n9366) );
  NOR3_X1 U11732 ( .A1(n9366), .A2(n10422), .A3(n10377), .ZN(n9367) );
  XNOR2_X1 U11733 ( .A(n10471), .B(n12741), .ZN(n10463) );
  NAND4_X1 U11734 ( .A1(n10451), .A2(n9367), .A3(n10437), .A4(n10463), .ZN(
        n9368) );
  OR4_X1 U11735 ( .A1(n10676), .A2(n10744), .A3(n10718), .A4(n9368), .ZN(n9369) );
  INV_X1 U11736 ( .A(n14186), .ZN(n10974) );
  XNOR2_X1 U11737 ( .A(n10974), .B(n11317), .ZN(n10964) );
  OR4_X1 U11738 ( .A1(n11113), .A2(n9369), .A3(n10776), .A4(n10964), .ZN(n9370) );
  NOR2_X1 U11739 ( .A1(n9371), .A2(n9370), .ZN(n9372) );
  XNOR2_X1 U11740 ( .A(n11406), .B(n12731), .ZN(n11210) );
  XNOR2_X1 U11741 ( .A(n13157), .B(n12729), .ZN(n13046) );
  NAND4_X1 U11742 ( .A1(n11394), .A2(n9372), .A3(n11210), .A4(n13046), .ZN(
        n9373) );
  NAND4_X1 U11743 ( .A1(n12946), .A2(n6496), .A3(n9374), .A4(n12986), .ZN(
        n9375) );
  OR4_X1 U11744 ( .A1(n12911), .A2(n12929), .A3(n12924), .A4(n9375), .ZN(n9376) );
  NOR2_X1 U11745 ( .A1(n12879), .A2(n9376), .ZN(n9378) );
  AND4_X1 U11746 ( .A1(n9379), .A2(n9378), .A3(n9377), .A4(n12884), .ZN(n9380)
         );
  MUX2_X1 U11747 ( .A(n9388), .B(n10942), .S(n8193), .Z(n9382) );
  OAI21_X1 U11748 ( .B1(n10519), .B2(n8194), .A(n9382), .ZN(n9384) );
  INV_X1 U11749 ( .A(n9945), .ZN(n9383) );
  AND2_X1 U11750 ( .A1(n9383), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11202) );
  NAND2_X1 U11751 ( .A1(n9385), .A2(n7570), .ZN(n9400) );
  OAI21_X1 U11752 ( .B1(n10020), .B2(n9952), .A(n10418), .ZN(n9386) );
  NAND2_X1 U11753 ( .A1(n11010), .A2(n10519), .ZN(n9390) );
  INV_X1 U11754 ( .A(n9388), .ZN(n9389) );
  XOR2_X1 U11755 ( .A(n10583), .B(n9389), .Z(n9392) );
  INV_X1 U11756 ( .A(n9390), .ZN(n9391) );
  NAND3_X1 U11757 ( .A1(n9392), .A2(n11202), .A3(n9391), .ZN(n9397) );
  INV_X1 U11758 ( .A(n11202), .ZN(n9395) );
  INV_X1 U11759 ( .A(n9393), .ZN(n9505) );
  NAND4_X1 U11760 ( .A1(n13002), .A2(n9505), .A3(n14637), .A4(n9956), .ZN(
        n9394) );
  OAI211_X1 U11761 ( .C1(n9952), .C2(n9395), .A(n9394), .B(P2_B_REG_SCAN_IN), 
        .ZN(n9396) );
  NAND3_X1 U11762 ( .A1(n9400), .A2(n9399), .A3(n9398), .ZN(P2_U3328) );
  INV_X1 U11763 ( .A(n9946), .ZN(n9401) );
  NOR2_X1 U11764 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n9403) );
  NOR2_X1 U11765 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), 
        .ZN(n9402) );
  NOR2_X1 U11766 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n9406) );
  NAND2_X1 U11767 ( .A1(n9569), .A2(n15080), .ZN(n9414) );
  NAND2_X1 U11768 ( .A1(n9413), .A2(n9566), .ZN(n9409) );
  NOR2_X1 U11769 ( .A1(n9414), .A2(n9409), .ZN(n9410) );
  INV_X1 U11770 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9411) );
  XNOR2_X1 U11771 ( .A(n6581), .B(n9411), .ZN(n9726) );
  INV_X1 U11772 ( .A(n9678), .ZN(n9420) );
  XNOR2_X1 U11773 ( .A(n9417), .B(P1_IR_REG_26__SCAN_IN), .ZN(n9677) );
  NAND2_X1 U11774 ( .A1(n6532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9418) );
  XNOR2_X1 U11775 ( .A(n9418), .B(P1_IR_REG_25__SCAN_IN), .ZN(n11293) );
  OR2_X2 U11776 ( .A1(n9420), .A2(n10095), .ZN(n14991) );
  NAND2_X1 U11777 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n9457), .ZN(n9448) );
  INV_X1 U11778 ( .A(n9457), .ZN(n14611) );
  AOI22_X1 U11779 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n9457), .B1(n14611), 
        .B2(n7704), .ZN(n14605) );
  NAND2_X1 U11780 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n9458), .ZN(n9447) );
  INV_X1 U11781 ( .A(n9458), .ZN(n14598) );
  AOI22_X1 U11782 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n9458), .B1(n14598), 
        .B2(n7718), .ZN(n14592) );
  MUX2_X1 U11783 ( .A(n13080), .B(P2_REG2_REG_1__SCAN_IN), .S(n12749), .Z(
        n12755) );
  AND2_X1 U11784 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n12756) );
  NAND2_X1 U11785 ( .A1(n12755), .A2(n12756), .ZN(n12754) );
  INV_X1 U11786 ( .A(n12749), .ZN(n9462) );
  NAND2_X1 U11787 ( .A1(n9462), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9421) );
  NAND2_X1 U11788 ( .A1(n12754), .A2(n9421), .ZN(n12767) );
  MUX2_X1 U11789 ( .A(n9422), .B(P2_REG2_REG_2__SCAN_IN), .S(n12761), .Z(
        n12768) );
  NAND2_X1 U11790 ( .A1(n12767), .A2(n12768), .ZN(n12766) );
  NAND2_X1 U11791 ( .A1(n9465), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9801) );
  NAND2_X1 U11792 ( .A1(n12766), .A2(n9801), .ZN(n9424) );
  MUX2_X1 U11793 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10380), .S(n9806), .Z(n9423) );
  NAND2_X1 U11794 ( .A1(n9424), .A2(n9423), .ZN(n9803) );
  NAND2_X1 U11795 ( .A1(n9806), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9425) );
  NAND2_X1 U11796 ( .A1(n9803), .A2(n9425), .ZN(n12774) );
  MUX2_X1 U11797 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10428), .S(n12777), .Z(
        n12773) );
  NAND2_X1 U11798 ( .A1(n12774), .A2(n12773), .ZN(n12772) );
  NAND2_X1 U11799 ( .A1(n12777), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9847) );
  NAND2_X1 U11800 ( .A1(n12772), .A2(n9847), .ZN(n9427) );
  INV_X1 U11801 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10467) );
  MUX2_X1 U11802 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n10467), .S(n9850), .Z(n9426) );
  NAND2_X1 U11803 ( .A1(n9427), .A2(n9426), .ZN(n12791) );
  NAND2_X1 U11804 ( .A1(n9850), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n12790) );
  NAND2_X1 U11805 ( .A1(n12791), .A2(n12790), .ZN(n9429) );
  MUX2_X1 U11806 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10443), .S(n12793), .Z(
        n9428) );
  NAND2_X1 U11807 ( .A1(n9429), .A2(n9428), .ZN(n12806) );
  NAND2_X1 U11808 ( .A1(n12793), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n12805) );
  NAND2_X1 U11809 ( .A1(n12806), .A2(n12805), .ZN(n9431) );
  MUX2_X1 U11810 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10455), .S(n12808), .Z(
        n9430) );
  NAND2_X1 U11811 ( .A1(n9431), .A2(n9430), .ZN(n12821) );
  NAND2_X1 U11812 ( .A1(n12808), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n12820) );
  NAND2_X1 U11813 ( .A1(n12821), .A2(n12820), .ZN(n9433) );
  INV_X1 U11814 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10729) );
  MUX2_X1 U11815 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10729), .S(n12824), .Z(
        n9432) );
  NAND2_X1 U11816 ( .A1(n9433), .A2(n9432), .ZN(n12823) );
  NAND2_X1 U11817 ( .A1(n12824), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U11818 ( .A1(n12823), .A2(n9434), .ZN(n9526) );
  INV_X1 U11819 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10751) );
  MUX2_X1 U11820 ( .A(n10751), .B(P2_REG2_REG_9__SCAN_IN), .S(n9484), .Z(n9435) );
  OR2_X1 U11821 ( .A1(n9526), .A2(n9435), .ZN(n9522) );
  NAND2_X1 U11822 ( .A1(n9749), .A2(n10751), .ZN(n9436) );
  AND2_X1 U11823 ( .A1(n9522), .A2(n9436), .ZN(n12835) );
  INV_X1 U11824 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10682) );
  MUX2_X1 U11825 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n10682), .S(n12840), .Z(
        n12834) );
  NAND2_X1 U11826 ( .A1(n12835), .A2(n12834), .ZN(n12833) );
  NAND2_X1 U11827 ( .A1(n12840), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9437) );
  NAND2_X1 U11828 ( .A1(n12833), .A2(n9437), .ZN(n9902) );
  MUX2_X1 U11829 ( .A(n10781), .B(P2_REG2_REG_11__SCAN_IN), .S(n9905), .Z(
        n9901) );
  OR2_X1 U11830 ( .A1(n9905), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U11831 ( .A1(n9900), .A2(n9974), .ZN(n9438) );
  MUX2_X1 U11832 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n10969), .S(n9922), .Z(
        n9976) );
  NAND2_X1 U11833 ( .A1(n9438), .A2(n9976), .ZN(n9978) );
  OR2_X1 U11834 ( .A1(n9922), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9439) );
  MUX2_X1 U11835 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n11120), .S(n10011), .Z(
        n10070) );
  NAND2_X1 U11836 ( .A1(n10071), .A2(n10070), .ZN(n10069) );
  NAND2_X1 U11837 ( .A1(n10011), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9440) );
  NAND2_X1 U11838 ( .A1(n10069), .A2(n9440), .ZN(n9441) );
  NAND2_X1 U11839 ( .A1(n9496), .A2(n9441), .ZN(n9444) );
  XNOR2_X1 U11840 ( .A(n9441), .B(n9496), .ZN(n14564) );
  INV_X1 U11841 ( .A(n14564), .ZN(n9442) );
  NAND2_X1 U11842 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n9442), .ZN(n9443) );
  NAND2_X1 U11843 ( .A1(n9444), .A2(n9443), .ZN(n9445) );
  NAND2_X1 U11844 ( .A1(n14584), .A2(n9445), .ZN(n9446) );
  INV_X1 U11845 ( .A(n14584), .ZN(n10180) );
  XNOR2_X1 U11846 ( .A(n10180), .B(n9445), .ZN(n14583) );
  NAND2_X1 U11847 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n14583), .ZN(n14581) );
  NAND2_X1 U11848 ( .A1(n9446), .A2(n14581), .ZN(n14591) );
  NAND2_X1 U11849 ( .A1(n14592), .A2(n14591), .ZN(n14590) );
  NAND2_X1 U11850 ( .A1(n9447), .A2(n14590), .ZN(n14604) );
  NAND2_X1 U11851 ( .A1(n14605), .A2(n14604), .ZN(n14603) );
  NAND2_X1 U11852 ( .A1(n9448), .A2(n14603), .ZN(n9449) );
  NOR2_X1 U11853 ( .A1(n9502), .A2(n9449), .ZN(n9450) );
  INV_X1 U11854 ( .A(n9502), .ZN(n14623) );
  XOR2_X1 U11855 ( .A(n14623), .B(n9449), .Z(n14616) );
  NOR2_X1 U11856 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n14616), .ZN(n14615) );
  NOR2_X1 U11857 ( .A1(n9450), .A2(n14615), .ZN(n9451) );
  XNOR2_X1 U11858 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n9451), .ZN(n9511) );
  INV_X1 U11859 ( .A(n9511), .ZN(n9509) );
  NAND2_X1 U11860 ( .A1(n9958), .A2(n9945), .ZN(n9453) );
  AOI21_X1 U11861 ( .B1(n9454), .B2(n9453), .A(n9452), .ZN(n9514) );
  INV_X1 U11862 ( .A(n9514), .ZN(n9507) );
  NAND2_X1 U11863 ( .A1(n9505), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13197) );
  NOR2_X1 U11864 ( .A1(n13197), .A2(n8143), .ZN(n9455) );
  NAND2_X1 U11865 ( .A1(n9507), .A2(n9455), .ZN(n14622) );
  AND2_X1 U11866 ( .A1(n8143), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9456) );
  NAND2_X1 U11867 ( .A1(n9507), .A2(n9456), .ZN(n14624) );
  AOI22_X1 U11868 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n9457), .B1(n14611), 
        .B2(n9500), .ZN(n14608) );
  AOI22_X1 U11869 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n9458), .B1(n14598), 
        .B2(n9499), .ZN(n14595) );
  INV_X1 U11870 ( .A(n9496), .ZN(n14571) );
  INV_X1 U11871 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9459) );
  MUX2_X1 U11872 ( .A(n9459), .B(P2_REG1_REG_1__SCAN_IN), .S(n12749), .Z(n9461) );
  AND2_X1 U11873 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9460) );
  NAND2_X1 U11874 ( .A1(n9461), .A2(n9460), .ZN(n12753) );
  NAND2_X1 U11875 ( .A1(n9462), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U11876 ( .A1(n12753), .A2(n9463), .ZN(n12764) );
  INV_X1 U11877 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9464) );
  MUX2_X1 U11878 ( .A(n9464), .B(P2_REG1_REG_2__SCAN_IN), .S(n12761), .Z(
        n12765) );
  NAND2_X1 U11879 ( .A1(n12764), .A2(n12765), .ZN(n12763) );
  NAND2_X1 U11880 ( .A1(n9465), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9808) );
  NAND2_X1 U11881 ( .A1(n12763), .A2(n9808), .ZN(n9468) );
  MUX2_X1 U11882 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9466), .S(n9806), .Z(n9467)
         );
  NAND2_X1 U11883 ( .A1(n9468), .A2(n9467), .ZN(n12780) );
  NAND2_X1 U11884 ( .A1(n9806), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n12779) );
  NAND2_X1 U11885 ( .A1(n12780), .A2(n12779), .ZN(n9471) );
  MUX2_X1 U11886 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n9469), .S(n12777), .Z(n9470) );
  NAND2_X1 U11887 ( .A1(n9471), .A2(n9470), .ZN(n12782) );
  NAND2_X1 U11888 ( .A1(n12777), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9852) );
  NAND2_X1 U11889 ( .A1(n12782), .A2(n9852), .ZN(n9474) );
  MUX2_X1 U11890 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n9472), .S(n9850), .Z(n9473)
         );
  NAND2_X1 U11891 ( .A1(n9474), .A2(n9473), .ZN(n12796) );
  NAND2_X1 U11892 ( .A1(n9850), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n12795) );
  NAND2_X1 U11893 ( .A1(n12796), .A2(n12795), .ZN(n9476) );
  MUX2_X1 U11894 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n14729), .S(n12793), .Z(
        n9475) );
  NAND2_X1 U11895 ( .A1(n9476), .A2(n9475), .ZN(n12811) );
  NAND2_X1 U11896 ( .A1(n12793), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n12810) );
  NAND2_X1 U11897 ( .A1(n12811), .A2(n12810), .ZN(n9479) );
  MUX2_X1 U11898 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9477), .S(n12808), .Z(n9478) );
  NAND2_X1 U11899 ( .A1(n9479), .A2(n9478), .ZN(n12827) );
  NAND2_X1 U11900 ( .A1(n12808), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U11901 ( .A1(n12827), .A2(n12826), .ZN(n9482) );
  MUX2_X1 U11902 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n9480), .S(n12824), .Z(n9481) );
  NAND2_X1 U11903 ( .A1(n9482), .A2(n9481), .ZN(n12829) );
  NAND2_X1 U11904 ( .A1(n12824), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9483) );
  NAND2_X1 U11905 ( .A1(n12829), .A2(n9483), .ZN(n9523) );
  MUX2_X1 U11906 ( .A(n9518), .B(P2_REG1_REG_9__SCAN_IN), .S(n9484), .Z(n9485)
         );
  OR2_X1 U11907 ( .A1(n9523), .A2(n9485), .ZN(n9520) );
  NAND2_X1 U11908 ( .A1(n9749), .A2(n9518), .ZN(n9486) );
  AND2_X1 U11909 ( .A1(n9520), .A2(n9486), .ZN(n12838) );
  MUX2_X1 U11910 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9487), .S(n12840), .Z(
        n12837) );
  NAND2_X1 U11911 ( .A1(n12838), .A2(n12837), .ZN(n12836) );
  NAND2_X1 U11912 ( .A1(n12840), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9907) );
  NAND2_X1 U11913 ( .A1(n12836), .A2(n9907), .ZN(n9490) );
  MUX2_X1 U11914 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9488), .S(n9905), .Z(n9489) );
  NAND2_X1 U11915 ( .A1(n9490), .A2(n9489), .ZN(n9909) );
  NAND2_X1 U11916 ( .A1(n9905), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9491) );
  NAND2_X1 U11917 ( .A1(n9909), .A2(n9491), .ZN(n9969) );
  MUX2_X1 U11918 ( .A(n9492), .B(P2_REG1_REG_12__SCAN_IN), .S(n9922), .Z(n9970) );
  OR2_X1 U11919 ( .A1(n9922), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U11920 ( .A1(n9967), .A2(n9493), .ZN(n10065) );
  MUX2_X1 U11921 ( .A(n7945), .B(P2_REG1_REG_13__SCAN_IN), .S(n10011), .Z(
        n10066) );
  NOR2_X1 U11922 ( .A1(n10065), .A2(n10066), .ZN(n14569) );
  AND2_X1 U11923 ( .A1(n10011), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n14565) );
  OR2_X1 U11924 ( .A1(n14569), .A2(n14565), .ZN(n9495) );
  NAND2_X1 U11925 ( .A1(n9496), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9494) );
  OAI211_X1 U11926 ( .C1(n9496), .C2(P2_REG1_REG_14__SCAN_IN), .A(n9495), .B(
        n9494), .ZN(n14567) );
  OAI21_X1 U11927 ( .B1(n7955), .B2(n14571), .A(n14567), .ZN(n9497) );
  NAND2_X1 U11928 ( .A1(n14584), .A2(n9497), .ZN(n9498) );
  XNOR2_X1 U11929 ( .A(n9497), .B(n10180), .ZN(n14580) );
  NAND2_X1 U11930 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n14580), .ZN(n14578) );
  NAND2_X1 U11931 ( .A1(n9498), .A2(n14578), .ZN(n14594) );
  NAND2_X1 U11932 ( .A1(n14595), .A2(n14594), .ZN(n14593) );
  OAI21_X1 U11933 ( .B1(n14598), .B2(n9499), .A(n14593), .ZN(n14607) );
  NAND2_X1 U11934 ( .A1(n14608), .A2(n14607), .ZN(n14606) );
  OAI21_X1 U11935 ( .B1(n14611), .B2(n9500), .A(n14606), .ZN(n9501) );
  XNOR2_X1 U11936 ( .A(n14623), .B(n9501), .ZN(n14618) );
  NAND2_X1 U11937 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n14618), .ZN(n14617) );
  NAND2_X1 U11938 ( .A1(n9502), .A2(n9501), .ZN(n9503) );
  NAND2_X1 U11939 ( .A1(n14617), .A2(n9503), .ZN(n9504) );
  XNOR2_X1 U11940 ( .A(n9504), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9510) );
  OR2_X1 U11941 ( .A1(n8143), .A2(P2_U3088), .ZN(n13194) );
  NOR2_X1 U11942 ( .A1(n13194), .A2(n9505), .ZN(n9506) );
  NAND2_X1 U11943 ( .A1(n9510), .A2(n14579), .ZN(n9508) );
  OAI211_X1 U11944 ( .C1(n9509), .C2(n14622), .A(n14624), .B(n9508), .ZN(n9513) );
  OAI22_X1 U11945 ( .A1(n9511), .A2(n14622), .B1(n9510), .B2(n14620), .ZN(
        n9512) );
  MUX2_X1 U11946 ( .A(n9513), .B(n9512), .S(n10583), .Z(n9516) );
  AND2_X1 U11947 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12594) );
  AND2_X1 U11948 ( .A1(n9514), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14577) );
  NOR2_X1 U11949 ( .A1(n14628), .A2(n14140), .ZN(n9515) );
  INV_X1 U11950 ( .A(n12513), .ZN(n11423) );
  NAND3_X1 U11951 ( .A1(n9523), .A2(n9749), .A3(n9518), .ZN(n9519) );
  AOI21_X1 U11952 ( .B1(n9520), .B2(n9519), .A(n14620), .ZN(n9534) );
  NAND3_X1 U11953 ( .A1(n9526), .A2(n9749), .A3(n10751), .ZN(n9521) );
  AOI21_X1 U11954 ( .B1(n9522), .B2(n9521), .A(n14622), .ZN(n9533) );
  NOR2_X1 U11955 ( .A1(n14622), .A2(n10751), .ZN(n9527) );
  INV_X1 U11956 ( .A(n14624), .ZN(n14585) );
  INV_X1 U11957 ( .A(n9523), .ZN(n9524) );
  NOR3_X1 U11958 ( .A1(n9524), .A2(n9518), .A3(n14620), .ZN(n9525) );
  AOI211_X1 U11959 ( .C1(n9527), .C2(n9526), .A(n14585), .B(n9525), .ZN(n9528)
         );
  NOR2_X1 U11960 ( .A1(n9528), .A2(n9749), .ZN(n9532) );
  INV_X1 U11961 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9530) );
  NAND2_X1 U11962 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n9529) );
  OAI21_X1 U11963 ( .B1(n14628), .B2(n9530), .A(n9529), .ZN(n9531) );
  OR4_X1 U11964 ( .A1(n9534), .A2(n9533), .A3(n9532), .A4(n9531), .ZN(P2_U3223) );
  INV_X1 U11965 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9535) );
  INV_X1 U11966 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9537) );
  NAND2_X1 U11967 ( .A1(n9539), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9540) );
  NAND2_X1 U11968 ( .A1(n10107), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9549) );
  AND2_X4 U11969 ( .A1(n11612), .A2(n7012), .ZN(n11743) );
  INV_X1 U11970 ( .A(n9699), .ZN(n9543) );
  NAND2_X1 U11971 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9544) );
  MUX2_X1 U11972 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9544), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n9547) );
  INV_X1 U11973 ( .A(n9545), .ZN(n9546) );
  NAND2_X1 U11974 ( .A1(n9547), .A2(n9546), .ZN(n13490) );
  INV_X1 U11975 ( .A(n13490), .ZN(n13496) );
  INV_X1 U11976 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13506) );
  NOR2_X1 U11977 ( .A1(n9657), .A2(n9629), .ZN(n9550) );
  XNOR2_X1 U11978 ( .A(n9550), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n13996) );
  MUX2_X1 U11979 ( .A(n13506), .B(n13996), .S(n11612), .Z(n10329) );
  OR2_X1 U11980 ( .A1(n10329), .A2(n9925), .ZN(n9551) );
  NAND2_X1 U11981 ( .A1(n14433), .A2(n9551), .ZN(n14469) );
  NAND2_X1 U11982 ( .A1(n9552), .A2(n9555), .ZN(n13974) );
  INV_X1 U11983 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9732) );
  INV_X1 U11984 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9612) );
  INV_X1 U11985 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9559) );
  XNOR2_X1 U11986 ( .A(n14469), .B(n10215), .ZN(n9565) );
  INV_X1 U11987 ( .A(n11444), .ZN(n9564) );
  NAND2_X1 U11988 ( .A1(n15191), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9563) );
  INV_X1 U11989 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9560) );
  INV_X1 U11990 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14343) );
  INV_X1 U11991 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9561) );
  OR2_X1 U11992 ( .A1(n10100), .A2(n9561), .ZN(n9562) );
  MUX2_X1 U11993 ( .A(n9565), .B(n9564), .S(n13486), .Z(n9590) );
  INV_X1 U11994 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9573) );
  INV_X1 U11995 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9567) );
  INV_X1 U11996 ( .A(n11434), .ZN(n9616) );
  INV_X1 U11997 ( .A(n9569), .ZN(n9570) );
  NAND2_X1 U11998 ( .A1(n9616), .A2(n9610), .ZN(n11739) );
  NAND2_X1 U11999 ( .A1(n9576), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9578) );
  XNOR2_X1 U12000 ( .A(n9578), .B(n9577), .ZN(n11430) );
  NAND2_X1 U12001 ( .A1(n14414), .A2(n13995), .ZN(n9579) );
  NAND2_X1 U12002 ( .A1(n9610), .A2(n13995), .ZN(n11747) );
  NAND2_X1 U12003 ( .A1(n15191), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9585) );
  INV_X1 U12004 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9580) );
  OR2_X1 U12005 ( .A1(n11634), .A2(n9580), .ZN(n9584) );
  INV_X1 U12006 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9731) );
  INV_X1 U12007 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9581) );
  OR2_X1 U12008 ( .A1(n10100), .A2(n9581), .ZN(n9582) );
  INV_X1 U12009 ( .A(n13984), .ZN(n13505) );
  AOI22_X1 U12010 ( .A1(n13865), .A2(n13486), .B1(n13484), .B2(n13835), .ZN(
        n9589) );
  NAND2_X1 U12011 ( .A1(n13486), .A2(n6972), .ZN(n10214) );
  XNOR2_X1 U12012 ( .A(n11444), .B(n10214), .ZN(n14472) );
  NAND2_X1 U12013 ( .A1(n11446), .A2(n9586), .ZN(n9587) );
  NAND2_X1 U12014 ( .A1(n13365), .A2(n9587), .ZN(n10212) );
  INV_X1 U12015 ( .A(n14509), .ZN(n14532) );
  NAND2_X1 U12016 ( .A1(n14472), .A2(n14532), .ZN(n9588) );
  OAI211_X1 U12017 ( .C1(n9590), .C2(n14540), .A(n9589), .B(n9588), .ZN(n14470) );
  NAND2_X1 U12018 ( .A1(n11434), .A2(n13822), .ZN(n9867) );
  INV_X1 U12019 ( .A(n11747), .ZN(n9591) );
  NAND2_X1 U12020 ( .A1(n9867), .A2(n9591), .ZN(n10096) );
  NAND2_X1 U12021 ( .A1(n10096), .A2(n9866), .ZN(n11792) );
  INV_X1 U12022 ( .A(P1_B_REG_SCAN_IN), .ZN(n13616) );
  OR2_X1 U12023 ( .A1(n11293), .A2(n13616), .ZN(n9592) );
  OR2_X1 U12024 ( .A1(n11240), .A2(n9592), .ZN(n9594) );
  NAND2_X1 U12025 ( .A1(n11240), .A2(n13616), .ZN(n9593) );
  AND3_X1 U12026 ( .A1(n9594), .A2(n9593), .A3(n9677), .ZN(n9675) );
  NOR4_X1 U12027 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9603) );
  NOR4_X1 U12028 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n9602) );
  INV_X1 U12029 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n15086) );
  INV_X1 U12030 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n15125) );
  INV_X1 U12031 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n15108) );
  INV_X1 U12032 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14466) );
  NAND4_X1 U12033 ( .A1(n15086), .A2(n15125), .A3(n15108), .A4(n14466), .ZN(
        n9600) );
  NOR4_X1 U12034 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9598) );
  NOR4_X1 U12035 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n9597) );
  NOR4_X1 U12036 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9596) );
  NOR4_X1 U12037 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9595) );
  NAND4_X1 U12038 ( .A1(n9598), .A2(n9597), .A3(n9596), .A4(n9595), .ZN(n9599)
         );
  NOR4_X1 U12039 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n9600), .A4(n9599), .ZN(n9601) );
  NAND3_X1 U12040 ( .A1(n9603), .A2(n9602), .A3(n9601), .ZN(n9604) );
  NAND2_X1 U12041 ( .A1(n9675), .A2(n9604), .ZN(n9871) );
  INV_X1 U12042 ( .A(n9871), .ZN(n9605) );
  OR2_X1 U12043 ( .A1(n11792), .A2(n9605), .ZN(n9880) );
  INV_X1 U12044 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n9607) );
  NOR2_X1 U12045 ( .A1(n9677), .A2(n11293), .ZN(n9606) );
  AOI21_X1 U12046 ( .B1(n9675), .B2(n9607), .A(n9606), .ZN(n9872) );
  INV_X1 U12047 ( .A(n9872), .ZN(n9917) );
  NOR2_X1 U12048 ( .A1(n9880), .A2(n9917), .ZN(n9857) );
  INV_X1 U12049 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9609) );
  NOR2_X1 U12050 ( .A1(n11240), .A2(n9677), .ZN(n9608) );
  AOI21_X1 U12051 ( .B1(n9675), .B2(n9609), .A(n9608), .ZN(n9879) );
  INV_X1 U12052 ( .A(n9879), .ZN(n9916) );
  NAND2_X1 U12053 ( .A1(n9857), .A2(n9916), .ZN(n13679) );
  NAND2_X1 U12054 ( .A1(n11434), .A2(n11430), .ZN(n11748) );
  INV_X1 U12055 ( .A(n9915), .ZN(n9611) );
  MUX2_X1 U12056 ( .A(n14470), .B(P1_REG2_REG_1__SCAN_IN), .S(n14439), .Z(
        n9621) );
  OR2_X1 U12057 ( .A1(n13875), .A2(n14468), .ZN(n13857) );
  OAI22_X1 U12058 ( .A1(n13857), .A2(n14469), .B1(n9612), .B2(n14416), .ZN(
        n9620) );
  INV_X1 U12059 ( .A(n11446), .ZN(n9613) );
  OR2_X1 U12060 ( .A1(n9613), .A2(n13822), .ZN(n14410) );
  INV_X1 U12061 ( .A(n14410), .ZN(n9614) );
  NAND2_X1 U12062 ( .A1(n14420), .A2(n9614), .ZN(n14121) );
  INV_X1 U12063 ( .A(n14472), .ZN(n9615) );
  NOR2_X1 U12064 ( .A1(n14121), .A2(n9615), .ZN(n9619) );
  NAND2_X1 U12065 ( .A1(n9616), .A2(n11433), .ZN(n11781) );
  OR2_X1 U12066 ( .A1(n11781), .A2(n13995), .ZN(n14415) );
  INV_X1 U12067 ( .A(n14415), .ZN(n9617) );
  NOR2_X1 U12068 ( .A1(n13876), .A2(n9925), .ZN(n9618) );
  OR4_X1 U12069 ( .A1(n9621), .A2(n9620), .A3(n9619), .A4(n9618), .ZN(P1_U3292) );
  NOR2_X1 U12070 ( .A1(n9657), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12515) );
  NAND2_X1 U12071 ( .A1(n9657), .A2(P3_U3151), .ZN(n12530) );
  OAI222_X1 U12072 ( .A1(n14809), .A2(P3_U3151), .B1(n12528), .B2(n9623), .C1(
        n9622), .C2(n12530), .ZN(P3_U3289) );
  INV_X1 U12073 ( .A(n9624), .ZN(n9626) );
  INV_X1 U12074 ( .A(SI_3_), .ZN(n9625) );
  OAI222_X1 U12075 ( .A1(n10854), .A2(P3_U3151), .B1(n12528), .B2(n9626), .C1(
        n9625), .C2(n12530), .ZN(P3_U3292) );
  OAI222_X1 U12076 ( .A1(P3_U3151), .A2(n14847), .B1(n12530), .B2(n9628), .C1(
        n12528), .C2(n9627), .ZN(P3_U3287) );
  OAI222_X1 U12077 ( .A1(n14746), .A2(P3_U3151), .B1(n12528), .B2(n9630), .C1(
        n9629), .C2(n12530), .ZN(P3_U3295) );
  INV_X1 U12078 ( .A(n9631), .ZN(n9633) );
  CLKBUF_X1 U12079 ( .A(n12530), .Z(n12521) );
  INV_X1 U12080 ( .A(SI_9_), .ZN(n9632) );
  OAI222_X1 U12081 ( .A1(n12528), .A2(n9633), .B1(n12521), .B2(n9632), .C1(
        n14867), .C2(P3_U3151), .ZN(P3_U3286) );
  OAI222_X1 U12082 ( .A1(P3_U3151), .A2(n6852), .B1(n12521), .B2(n6916), .C1(
        n12528), .C2(n9634), .ZN(P3_U3294) );
  INV_X1 U12083 ( .A(n9635), .ZN(n9637) );
  INV_X1 U12084 ( .A(SI_2_), .ZN(n9636) );
  OAI222_X1 U12085 ( .A1(n12528), .A2(n9637), .B1(n12521), .B2(n9636), .C1(
        n10892), .C2(P3_U3151), .ZN(P3_U3293) );
  INV_X1 U12086 ( .A(n9638), .ZN(n9640) );
  INV_X1 U12087 ( .A(SI_7_), .ZN(n9639) );
  OAI222_X1 U12088 ( .A1(n12528), .A2(n9640), .B1(n12521), .B2(n9639), .C1(
        n10900), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U12089 ( .A(n9641), .ZN(n9643) );
  INV_X1 U12090 ( .A(SI_4_), .ZN(n9642) );
  INV_X1 U12091 ( .A(n10895), .ZN(n14775) );
  OAI222_X1 U12092 ( .A1(n12528), .A2(n9643), .B1(n12521), .B2(n9642), .C1(
        n14775), .C2(P3_U3151), .ZN(P3_U3291) );
  INV_X1 U12093 ( .A(n9644), .ZN(n9645) );
  INV_X1 U12094 ( .A(SI_5_), .ZN(n15097) );
  OAI222_X1 U12095 ( .A1(n12528), .A2(n9645), .B1(n12521), .B2(n15097), .C1(
        n14793), .C2(P3_U3151), .ZN(P3_U3290) );
  NOR2_X1 U12096 ( .A1(n9657), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13196) );
  INV_X2 U12097 ( .A(n13196), .ZN(n13201) );
  OAI222_X1 U12098 ( .A1(n13201), .A2(n9646), .B1(n13199), .B2(n9992), .C1(
        n12761), .C2(P2_U3088), .ZN(P2_U3325) );
  INV_X1 U12099 ( .A(n10224), .ZN(n9659) );
  INV_X1 U12100 ( .A(n12777), .ZN(n9647) );
  OAI222_X1 U12101 ( .A1(n13201), .A2(n9648), .B1(n13199), .B2(n9659), .C1(
        n9647), .C2(P2_U3088), .ZN(P2_U3323) );
  INV_X1 U12102 ( .A(n10108), .ZN(n9694) );
  INV_X1 U12103 ( .A(n9806), .ZN(n9649) );
  OAI222_X1 U12104 ( .A1(n13201), .A2(n9711), .B1(n13199), .B2(n9694), .C1(
        n9649), .C2(P2_U3088), .ZN(P2_U3324) );
  INV_X1 U12105 ( .A(n9650), .ZN(n9652) );
  INV_X1 U12106 ( .A(SI_10_), .ZN(n9651) );
  INV_X1 U12107 ( .A(n11098), .ZN(n11095) );
  OAI222_X1 U12108 ( .A1(n12528), .A2(n9652), .B1(n12521), .B2(n9651), .C1(
        n11095), .C2(P3_U3151), .ZN(P3_U3285) );
  NAND2_X1 U12109 ( .A1(n9545), .A2(n9653), .ZN(n9688) );
  NAND2_X1 U12110 ( .A1(n9690), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9654) );
  MUX2_X1 U12111 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9654), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n9656) );
  INV_X1 U12112 ( .A(n9669), .ZN(n9655) );
  AND2_X1 U12113 ( .A1(n9656), .A2(n9655), .ZN(n10225) );
  INV_X1 U12114 ( .A(n10225), .ZN(n13534) );
  OAI222_X1 U12115 ( .A1(n13986), .A2(n9659), .B1(n13534), .B2(P1_U3086), .C1(
        n9658), .C2(n13988), .ZN(P1_U3351) );
  OAI222_X1 U12116 ( .A1(n12528), .A2(n9661), .B1(n12521), .B2(n9660), .C1(
        n12018), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U12117 ( .A(n10253), .ZN(n9666) );
  INV_X1 U12118 ( .A(n9850), .ZN(n9662) );
  OAI222_X1 U12119 ( .A1(n13201), .A2(n9663), .B1(n13199), .B2(n9666), .C1(
        P2_U3088), .C2(n9662), .ZN(P2_U3322) );
  OR2_X1 U12120 ( .A1(n9669), .A2(n13973), .ZN(n9664) );
  XNOR2_X1 U12121 ( .A(n9664), .B(P1_IR_REG_5__SCAN_IN), .ZN(n13558) );
  INV_X1 U12122 ( .A(n13558), .ZN(n9665) );
  OAI222_X1 U12123 ( .A1(n13988), .A2(n9667), .B1(n13986), .B2(n9666), .C1(
        P1_U3086), .C2(n9665), .ZN(P1_U3350) );
  INV_X1 U12124 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9668) );
  OR2_X1 U12125 ( .A1(n9696), .A2(n13973), .ZN(n9670) );
  XNOR2_X1 U12126 ( .A(n9670), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10258) );
  INV_X1 U12127 ( .A(n10258), .ZN(n9723) );
  OAI222_X1 U12128 ( .A1(n13986), .A2(n10257), .B1(n9723), .B2(P1_U3086), .C1(
        n9671), .C2(n13988), .ZN(P1_U3349) );
  INV_X1 U12129 ( .A(n12793), .ZN(n12787) );
  OAI222_X1 U12130 ( .A1(n13201), .A2(n9672), .B1(n13199), .B2(n10257), .C1(
        n12787), .C2(P2_U3088), .ZN(P2_U3321) );
  OAI222_X1 U12131 ( .A1(n12528), .A2(n9674), .B1(n12036), .B2(P3_U3151), .C1(
        n9673), .C2(n12521), .ZN(P3_U3283) );
  INV_X1 U12132 ( .A(n9675), .ZN(n9676) );
  AND2_X2 U12133 ( .A1(n9676), .A2(n9866), .ZN(n14467) );
  INV_X1 U12134 ( .A(n9677), .ZN(n13992) );
  NAND2_X1 U12135 ( .A1(n9678), .A2(n13992), .ZN(n9680) );
  OAI22_X1 U12136 ( .A1(n14467), .A2(P1_D_REG_1__SCAN_IN), .B1(n11293), .B2(
        n9680), .ZN(n9679) );
  INV_X1 U12137 ( .A(n9679), .ZN(P1_U3446) );
  OAI22_X1 U12138 ( .A1(n14467), .A2(P1_D_REG_0__SCAN_IN), .B1(n11240), .B2(
        n9680), .ZN(n9681) );
  INV_X1 U12139 ( .A(n9681), .ZN(P1_U3445) );
  OAI222_X1 U12140 ( .A1(P2_U3088), .A2(n12749), .B1(n13199), .B2(n9699), .C1(
        n9682), .C2(n13201), .ZN(P2_U3326) );
  INV_X1 U12141 ( .A(n12808), .ZN(n12801) );
  OAI222_X1 U12142 ( .A1(n13201), .A2(n9683), .B1(n13199), .B2(n10269), .C1(
        n12801), .C2(P2_U3088), .ZN(P2_U3320) );
  NOR2_X1 U12143 ( .A1(n9545), .A2(n13973), .ZN(n9684) );
  MUX2_X1 U12144 ( .A(n13973), .B(n9684), .S(P1_IR_REG_2__SCAN_IN), .Z(n9686)
         );
  INV_X1 U12145 ( .A(n9688), .ZN(n9685) );
  NOR2_X1 U12146 ( .A1(n9686), .A2(n9685), .ZN(n9994) );
  INV_X1 U12147 ( .A(n9994), .ZN(n13512) );
  OAI222_X1 U12148 ( .A1(n13986), .A2(n9992), .B1(n13512), .B2(P1_U3086), .C1(
        n9687), .C2(n13988), .ZN(P1_U3353) );
  NAND2_X1 U12149 ( .A1(n9688), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9689) );
  MUX2_X1 U12150 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9689), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n9691) );
  AND2_X1 U12151 ( .A1(n9691), .A2(n9690), .ZN(n13524) );
  INV_X1 U12152 ( .A(n13524), .ZN(n9693) );
  OAI222_X1 U12153 ( .A1(n13986), .A2(n9694), .B1(n9693), .B2(P1_U3086), .C1(
        n9692), .C2(n13988), .ZN(P1_U3352) );
  INV_X1 U12154 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9695) );
  NAND2_X1 U12155 ( .A1(n9696), .A2(n9695), .ZN(n9700) );
  NAND2_X1 U12156 ( .A1(n9700), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9697) );
  XNOR2_X1 U12157 ( .A(n9697), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10270) );
  INV_X1 U12158 ( .A(n10270), .ZN(n9799) );
  OAI222_X1 U12159 ( .A1(n13986), .A2(n10269), .B1(n9799), .B2(P1_U3086), .C1(
        n9698), .C2(n13988), .ZN(P1_U3348) );
  OAI222_X1 U12160 ( .A1(n13988), .A2(n6839), .B1(n13490), .B2(P1_U3086), .C1(
        n13986), .C2(n9699), .ZN(P1_U3354) );
  NAND2_X1 U12161 ( .A1(n9702), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9701) );
  MUX2_X1 U12162 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9701), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n9703) );
  NAND2_X1 U12163 ( .A1(n9703), .A2(n9746), .ZN(n9764) );
  OAI222_X1 U12164 ( .A1(n13986), .A2(n10389), .B1(n9764), .B2(P1_U3086), .C1(
        n9704), .C2(n13988), .ZN(P1_U3347) );
  INV_X1 U12165 ( .A(n12824), .ZN(n12816) );
  OAI222_X1 U12166 ( .A1(n13201), .A2(n9705), .B1(n13199), .B2(n10389), .C1(
        n12816), .C2(P2_U3088), .ZN(P2_U3319) );
  NAND2_X1 U12167 ( .A1(n15191), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9710) );
  OR2_X1 U12168 ( .A1(n11634), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9709) );
  INV_X1 U12169 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9733) );
  INV_X1 U12170 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9706) );
  OR2_X1 U12171 ( .A1(n10100), .A2(n9706), .ZN(n9707) );
  MUX2_X1 U12172 ( .A(n9711), .B(n10221), .S(P1_U4016), .Z(n9712) );
  INV_X1 U12173 ( .A(n9712), .ZN(P1_U3563) );
  INV_X1 U12174 ( .A(n12061), .ZN(n12055) );
  OAI222_X1 U12175 ( .A1(n12528), .A2(n9714), .B1(n12055), .B2(P3_U3151), .C1(
        n9713), .C2(n12530), .ZN(P3_U3282) );
  INV_X1 U12176 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9715) );
  MUX2_X1 U12177 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n9715), .S(n9994), .Z(n13515) );
  INV_X1 U12178 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n13491) );
  MUX2_X1 U12179 ( .A(n13491), .B(P1_REG2_REG_1__SCAN_IN), .S(n13490), .Z(
        n9716) );
  AND2_X1 U12180 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13492) );
  NAND2_X1 U12181 ( .A1(n9716), .A2(n13492), .ZN(n13495) );
  OAI21_X1 U12182 ( .B1(n13491), .B2(n13490), .A(n13495), .ZN(n13514) );
  NAND2_X1 U12183 ( .A1(n13515), .A2(n13514), .ZN(n13527) );
  NAND2_X1 U12184 ( .A1(n9994), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13526) );
  NAND2_X1 U12185 ( .A1(n13527), .A2(n13526), .ZN(n9719) );
  INV_X1 U12186 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9717) );
  MUX2_X1 U12187 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9717), .S(n13524), .Z(n9718) );
  NAND2_X1 U12188 ( .A1(n9719), .A2(n9718), .ZN(n13538) );
  NAND2_X1 U12189 ( .A1(n13524), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13537) );
  INV_X1 U12190 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9720) );
  MUX2_X1 U12191 ( .A(n9720), .B(P1_REG2_REG_4__SCAN_IN), .S(n10225), .Z(
        n13539) );
  AOI21_X1 U12192 ( .B1(n13538), .B2(n13537), .A(n13539), .ZN(n13536) );
  NOR2_X1 U12193 ( .A1(n13534), .A2(n9720), .ZN(n13557) );
  INV_X1 U12194 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10234) );
  MUX2_X1 U12195 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10234), .S(n13558), .Z(
        n9721) );
  OAI21_X1 U12196 ( .B1(n13536), .B2(n13557), .A(n9721), .ZN(n13563) );
  NAND2_X1 U12197 ( .A1(n13558), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9780) );
  INV_X1 U12198 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9722) );
  MUX2_X1 U12199 ( .A(n9722), .B(P1_REG2_REG_6__SCAN_IN), .S(n10258), .Z(n9779) );
  AOI21_X1 U12200 ( .B1(n13563), .B2(n9780), .A(n9779), .ZN(n9788) );
  NOR2_X1 U12201 ( .A1(n9723), .A2(n9722), .ZN(n9787) );
  INV_X1 U12202 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10296) );
  MUX2_X1 U12203 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10296), .S(n10270), .Z(
        n9786) );
  OAI21_X1 U12204 ( .B1(n9788), .B2(n9787), .A(n9786), .ZN(n9790) );
  NAND2_X1 U12205 ( .A1(n10270), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9725) );
  INV_X1 U12206 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9763) );
  MUX2_X1 U12207 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n9763), .S(n9764), .Z(n9724)
         );
  AOI21_X1 U12208 ( .B1(n9790), .B2(n9725), .A(n9724), .ZN(n9767) );
  NAND3_X1 U12209 ( .A1(n9790), .A2(n9725), .A3(n9724), .ZN(n9730) );
  INV_X1 U12210 ( .A(n9726), .ZN(n9728) );
  OR2_X1 U12211 ( .A1(n11747), .A2(n9728), .ZN(n9727) );
  NAND2_X1 U12212 ( .A1(n9727), .A2(n11612), .ZN(n9740) );
  NAND2_X1 U12213 ( .A1(n9728), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11795) );
  INV_X1 U12214 ( .A(n11795), .ZN(n11204) );
  NOR2_X1 U12215 ( .A1(n9866), .A2(n11204), .ZN(n9739) );
  OR2_X1 U12216 ( .A1(n9740), .A2(n9739), .ZN(n14348) );
  NAND2_X1 U12217 ( .A1(n13505), .A2(n7189), .ZN(n9729) );
  NAND2_X1 U12218 ( .A1(n9730), .A2(n14370), .ZN(n9745) );
  MUX2_X1 U12219 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9731), .S(n9994), .Z(n13510) );
  MUX2_X1 U12220 ( .A(n9732), .B(P1_REG1_REG_1__SCAN_IN), .S(n13490), .Z(
        n13488) );
  AND2_X1 U12221 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13489) );
  NAND2_X1 U12222 ( .A1(n13488), .A2(n13489), .ZN(n13487) );
  OAI21_X1 U12223 ( .B1(n9732), .B2(n13490), .A(n13487), .ZN(n13509) );
  NAND2_X1 U12224 ( .A1(n13510), .A2(n13509), .ZN(n13522) );
  NAND2_X1 U12225 ( .A1(n9994), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13521) );
  NAND2_X1 U12226 ( .A1(n13522), .A2(n13521), .ZN(n9735) );
  MUX2_X1 U12227 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9733), .S(n13524), .Z(n9734) );
  NAND2_X1 U12228 ( .A1(n9735), .A2(n9734), .ZN(n13543) );
  NAND2_X1 U12229 ( .A1(n13524), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n13542) );
  INV_X1 U12230 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n15068) );
  MUX2_X1 U12231 ( .A(n15068), .B(P1_REG1_REG_4__SCAN_IN), .S(n10225), .Z(
        n13544) );
  AOI21_X1 U12232 ( .B1(n13543), .B2(n13542), .A(n13544), .ZN(n13541) );
  AOI21_X1 U12233 ( .B1(n10225), .B2(P1_REG1_REG_4__SCAN_IN), .A(n13541), .ZN(
        n13554) );
  INV_X1 U12234 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14551) );
  MUX2_X1 U12235 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n14551), .S(n13558), .Z(
        n13555) );
  NAND2_X1 U12236 ( .A1(n13554), .A2(n13555), .ZN(n13553) );
  OAI21_X1 U12237 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n13558), .A(n13553), .ZN(
        n9778) );
  INV_X1 U12238 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14553) );
  MUX2_X1 U12239 ( .A(n14553), .B(P1_REG1_REG_6__SCAN_IN), .S(n10258), .Z(
        n9777) );
  NOR2_X1 U12240 ( .A1(n9778), .A2(n9777), .ZN(n9776) );
  AOI21_X1 U12241 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n10258), .A(n9776), .ZN(
        n9793) );
  INV_X1 U12242 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14555) );
  MUX2_X1 U12243 ( .A(n14555), .B(P1_REG1_REG_7__SCAN_IN), .S(n10270), .Z(
        n9792) );
  NOR2_X1 U12244 ( .A1(n9793), .A2(n9792), .ZN(n9791) );
  AOI21_X1 U12245 ( .B1(n10270), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9791), .ZN(
        n9737) );
  INV_X1 U12246 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n14557) );
  MUX2_X1 U12247 ( .A(n14557), .B(P1_REG1_REG_8__SCAN_IN), .S(n9764), .Z(n9736) );
  NOR2_X1 U12248 ( .A1(n9737), .A2(n9736), .ZN(n9738) );
  OR2_X1 U12249 ( .A1(n14348), .A2(n7189), .ZN(n14354) );
  OAI21_X1 U12250 ( .B1(n9738), .B2(n9760), .A(n14367), .ZN(n9744) );
  INV_X1 U12251 ( .A(n9764), .ZN(n10390) );
  INV_X1 U12252 ( .A(n9739), .ZN(n9741) );
  AND2_X1 U12253 ( .A1(n9741), .A2(n9740), .ZN(n14346) );
  INV_X1 U12254 ( .A(n14346), .ZN(n14992) );
  INV_X1 U12255 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14017) );
  NAND2_X1 U12256 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11071) );
  OAI21_X1 U12257 ( .B1(n14992), .B2(n14017), .A(n11071), .ZN(n9742) );
  AOI21_X1 U12258 ( .B1(n10390), .B2(n14357), .A(n9742), .ZN(n9743) );
  OAI211_X1 U12259 ( .C1(n9767), .C2(n9745), .A(n9744), .B(n9743), .ZN(
        P1_U3251) );
  INV_X1 U12260 ( .A(n10541), .ZN(n9750) );
  XNOR2_X1 U12261 ( .A(n9817), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10542) );
  INV_X1 U12262 ( .A(n10542), .ZN(n9747) );
  OAI222_X1 U12263 ( .A1(n13988), .A2(n9748), .B1(n13986), .B2(n9750), .C1(
        P1_U3086), .C2(n9747), .ZN(P1_U3346) );
  OAI222_X1 U12264 ( .A1(n13201), .A2(n9751), .B1(n13199), .B2(n9750), .C1(
        P2_U3088), .C2(n9749), .ZN(P2_U3318) );
  INV_X1 U12265 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9752) );
  NAND2_X1 U12266 ( .A1(n9817), .A2(n9752), .ZN(n9753) );
  NAND2_X1 U12267 ( .A1(n9753), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9754) );
  XNOR2_X1 U12268 ( .A(n9754), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10547) );
  INV_X1 U12269 ( .A(n10547), .ZN(n10050) );
  OAI222_X1 U12270 ( .A1(n13986), .A2(n10546), .B1(n10050), .B2(P1_U3086), 
        .C1(n9755), .C2(n13988), .ZN(P1_U3345) );
  INV_X1 U12271 ( .A(n12840), .ZN(n9756) );
  OAI222_X1 U12272 ( .A1(n13201), .A2(n9757), .B1(n13199), .B2(n10546), .C1(
        n9756), .C2(P2_U3088), .ZN(P2_U3317) );
  NOR2_X1 U12273 ( .A1(n10390), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9758) );
  INV_X1 U12274 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n14559) );
  MUX2_X1 U12275 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n14559), .S(n10542), .Z(
        n9759) );
  OAI21_X1 U12276 ( .B1(n9760), .B2(n9758), .A(n9759), .ZN(n9822) );
  INV_X1 U12277 ( .A(n9822), .ZN(n9762) );
  NOR3_X1 U12278 ( .A1(n9760), .A2(n9759), .A3(n9758), .ZN(n9761) );
  OAI21_X1 U12279 ( .B1(n9762), .B2(n9761), .A(n14367), .ZN(n9773) );
  INV_X1 U12280 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n15066) );
  NAND2_X1 U12281 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n11265) );
  OAI21_X1 U12282 ( .B1(n14992), .B2(n15066), .A(n11265), .ZN(n9771) );
  NOR2_X1 U12283 ( .A1(n9764), .A2(n9763), .ZN(n9766) );
  INV_X1 U12284 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10608) );
  MUX2_X1 U12285 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10608), .S(n10542), .Z(
        n9765) );
  OAI21_X1 U12286 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(n9830) );
  INV_X1 U12287 ( .A(n9830), .ZN(n9769) );
  NOR3_X1 U12288 ( .A1(n9767), .A2(n9766), .A3(n9765), .ZN(n9768) );
  NOR3_X1 U12289 ( .A1(n9769), .A2(n9768), .A3(n14360), .ZN(n9770) );
  AOI211_X1 U12290 ( .C1(n14357), .C2(n10542), .A(n9771), .B(n9770), .ZN(n9772) );
  NAND2_X1 U12291 ( .A1(n9773), .A2(n9772), .ZN(P1_U3252) );
  INV_X1 U12292 ( .A(n12071), .ZN(n9774) );
  OAI222_X1 U12293 ( .A1(n12528), .A2(n9775), .B1(n12521), .B2(n6793), .C1(
        n9774), .C2(P3_U3151), .ZN(P3_U3281) );
  AOI211_X1 U12294 ( .C1(n9778), .C2(n9777), .A(n14354), .B(n9776), .ZN(n9785)
         );
  AND3_X1 U12295 ( .A1(n13563), .A2(n9780), .A3(n9779), .ZN(n9781) );
  NOR3_X1 U12296 ( .A1(n14360), .A2(n9788), .A3(n9781), .ZN(n9784) );
  INV_X1 U12297 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14012) );
  NAND2_X1 U12298 ( .A1(n14357), .A2(n10258), .ZN(n9782) );
  NAND2_X1 U12299 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10763) );
  OAI211_X1 U12300 ( .C1(n14992), .C2(n14012), .A(n9782), .B(n10763), .ZN(
        n9783) );
  OR3_X1 U12301 ( .A1(n9785), .A2(n9784), .A3(n9783), .ZN(P1_U3249) );
  OR3_X1 U12302 ( .A1(n9788), .A2(n9787), .A3(n9786), .ZN(n9789) );
  NAND3_X1 U12303 ( .A1(n9790), .A2(n14370), .A3(n9789), .ZN(n9798) );
  NAND2_X1 U12304 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n10822) );
  AOI211_X1 U12305 ( .C1(n9793), .C2(n9792), .A(n9791), .B(n14354), .ZN(n9794)
         );
  INV_X1 U12306 ( .A(n9794), .ZN(n9795) );
  NAND2_X1 U12307 ( .A1(n10822), .A2(n9795), .ZN(n9796) );
  AOI21_X1 U12308 ( .B1(n14346), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n9796), .ZN(
        n9797) );
  OAI211_X1 U12309 ( .C1(n14375), .C2(n9799), .A(n9798), .B(n9797), .ZN(
        P1_U3250) );
  MUX2_X1 U12310 ( .A(n10380), .B(P2_REG2_REG_3__SCAN_IN), .S(n9806), .Z(n9800) );
  NAND3_X1 U12311 ( .A1(n12766), .A2(n9801), .A3(n9800), .ZN(n9802) );
  NAND2_X1 U12312 ( .A1(n9803), .A2(n9802), .ZN(n9812) );
  INV_X1 U12313 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14052) );
  AOI22_X1 U12314 ( .A1(n14585), .A2(n9806), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        P2_U3088), .ZN(n9804) );
  OAI21_X1 U12315 ( .B1(n14628), .B2(n14052), .A(n9804), .ZN(n9805) );
  INV_X1 U12316 ( .A(n9805), .ZN(n9811) );
  MUX2_X1 U12317 ( .A(n9466), .B(P2_REG1_REG_3__SCAN_IN), .S(n9806), .Z(n9807)
         );
  NAND3_X1 U12318 ( .A1(n12763), .A2(n9808), .A3(n9807), .ZN(n9809) );
  NAND3_X1 U12319 ( .A1(n14579), .A2(n12780), .A3(n9809), .ZN(n9810) );
  OAI211_X1 U12320 ( .C1(n14622), .C2(n9812), .A(n9811), .B(n9810), .ZN(
        P2_U3217) );
  OAI222_X1 U12321 ( .A1(n12528), .A2(n9814), .B1(n12530), .B2(n9813), .C1(
        n12112), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12322 ( .A(n10995), .ZN(n9820) );
  OR2_X1 U12323 ( .A1(n9815), .A2(n13973), .ZN(n9816) );
  NAND2_X1 U12324 ( .A1(n9817), .A2(n9816), .ZN(n9913) );
  INV_X1 U12325 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9818) );
  XNOR2_X1 U12326 ( .A(n9913), .B(n9818), .ZN(n13572) );
  INV_X1 U12327 ( .A(n13572), .ZN(n10054) );
  OAI222_X1 U12328 ( .A1(n13988), .A2(n9819), .B1(n13986), .B2(n9820), .C1(
        P1_U3086), .C2(n10054), .ZN(P1_U3344) );
  INV_X1 U12329 ( .A(n9905), .ZN(n9903) );
  OAI222_X1 U12330 ( .A1(n13201), .A2(n9821), .B1(n13199), .B2(n9820), .C1(
        P2_U3088), .C2(n9903), .ZN(P2_U3316) );
  OAI21_X1 U12331 ( .B1(n10542), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9822), .ZN(
        n9826) );
  INV_X1 U12332 ( .A(n9826), .ZN(n9824) );
  INV_X1 U12333 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10553) );
  MUX2_X1 U12334 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10553), .S(n10547), .Z(
        n9823) );
  OAI21_X1 U12335 ( .B1(n9824), .B2(n9823), .A(n14367), .ZN(n9835) );
  MUX2_X1 U12336 ( .A(n10553), .B(P1_REG1_REG_10__SCAN_IN), .S(n10547), .Z(
        n9825) );
  NOR2_X1 U12337 ( .A1(n9826), .A2(n9825), .ZN(n10053) );
  INV_X1 U12338 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14020) );
  NAND2_X1 U12339 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n11343)
         );
  OAI21_X1 U12340 ( .B1(n14992), .B2(n14020), .A(n11343), .ZN(n9827) );
  AOI21_X1 U12341 ( .B1(n10547), .B2(n14357), .A(n9827), .ZN(n9834) );
  NAND2_X1 U12342 ( .A1(n10542), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9829) );
  INV_X1 U12343 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10571) );
  MUX2_X1 U12344 ( .A(n10571), .B(P1_REG2_REG_10__SCAN_IN), .S(n10547), .Z(
        n9828) );
  AOI21_X1 U12345 ( .B1(n9830), .B2(n9829), .A(n9828), .ZN(n13575) );
  INV_X1 U12346 ( .A(n13575), .ZN(n9832) );
  NAND3_X1 U12347 ( .A1(n9830), .A2(n9829), .A3(n9828), .ZN(n9831) );
  NAND3_X1 U12348 ( .A1(n9832), .A2(n14370), .A3(n9831), .ZN(n9833) );
  OAI211_X1 U12349 ( .C1(n9835), .C2(n10053), .A(n9834), .B(n9833), .ZN(
        P1_U3253) );
  INV_X1 U12350 ( .A(n14622), .ZN(n14582) );
  AOI22_X1 U12351 ( .A1(n14582), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n14579), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n9840) );
  INV_X1 U12352 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9836) );
  NAND2_X1 U12353 ( .A1(n14579), .A2(n9836), .ZN(n9837) );
  OAI211_X1 U12354 ( .C1(P2_REG2_REG_0__SCAN_IN), .C2(n14622), .A(n9837), .B(
        n14624), .ZN(n9838) );
  INV_X1 U12355 ( .A(n9838), .ZN(n9839) );
  MUX2_X1 U12356 ( .A(n9840), .B(n9839), .S(P2_IR_REG_0__SCAN_IN), .Z(n9843)
         );
  NOR2_X1 U12357 ( .A1(n9965), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9841) );
  AOI21_X1 U12358 ( .B1(n14577), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n9841), .ZN(
        n9842) );
  NAND2_X1 U12359 ( .A1(n9843), .A2(n9842), .ZN(P2_U3214) );
  INV_X1 U12360 ( .A(n12126), .ZN(n12136) );
  OAI222_X1 U12361 ( .A1(n12528), .A2(n9845), .B1(n12136), .B2(P3_U3151), .C1(
        n9844), .C2(n12530), .ZN(P3_U3279) );
  INV_X1 U12362 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9856) );
  AND2_X1 U12363 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10092) );
  MUX2_X1 U12364 ( .A(n10467), .B(P2_REG2_REG_5__SCAN_IN), .S(n9850), .Z(n9846) );
  NAND3_X1 U12365 ( .A1(n12772), .A2(n9847), .A3(n9846), .ZN(n9848) );
  AND3_X1 U12366 ( .A1(n14582), .A2(n12791), .A3(n9848), .ZN(n9849) );
  AOI211_X1 U12367 ( .C1(n14585), .C2(n9850), .A(n10092), .B(n9849), .ZN(n9855) );
  MUX2_X1 U12368 ( .A(n9472), .B(P2_REG1_REG_5__SCAN_IN), .S(n9850), .Z(n9851)
         );
  NAND3_X1 U12369 ( .A1(n12782), .A2(n9852), .A3(n9851), .ZN(n9853) );
  NAND3_X1 U12370 ( .A1(n14579), .A2(n12796), .A3(n9853), .ZN(n9854) );
  OAI211_X1 U12371 ( .C1(n9856), .C2(n14628), .A(n9855), .B(n9854), .ZN(
        P2_U3219) );
  NAND2_X1 U12372 ( .A1(n9857), .A2(n9879), .ZN(n13463) );
  INV_X1 U12373 ( .A(n10095), .ZN(n9858) );
  NAND2_X1 U12374 ( .A1(n13486), .A2(n13206), .ZN(n9865) );
  OAI22_X1 U12375 ( .A1(n13367), .A2(n10329), .B1(n10095), .B2(n14343), .ZN(
        n9863) );
  INV_X1 U12376 ( .A(n9863), .ZN(n9864) );
  NAND2_X1 U12377 ( .A1(n9865), .A2(n9864), .ZN(n9928) );
  XNOR2_X1 U12378 ( .A(n9929), .B(n9928), .ZN(n13501) );
  NAND4_X1 U12379 ( .A1(n9872), .A2(n9879), .A3(n9866), .A4(n9871), .ZN(n9869)
         );
  AND2_X1 U12380 ( .A1(n11433), .A2(n11430), .ZN(n9878) );
  NAND2_X1 U12381 ( .A1(n9867), .A2(n9878), .ZN(n14528) );
  NAND2_X1 U12382 ( .A1(n14528), .A2(n11747), .ZN(n9868) );
  NAND2_X1 U12383 ( .A1(n13501), .A2(n14233), .ZN(n9876) );
  OR2_X1 U12384 ( .A1(n9869), .A2(n14415), .ZN(n9870) );
  NAND3_X1 U12385 ( .A1(n9879), .A2(n9872), .A3(n9871), .ZN(n9873) );
  NAND2_X1 U12386 ( .A1(n9873), .A2(n9915), .ZN(n10097) );
  INV_X1 U12387 ( .A(n11792), .ZN(n9874) );
  NAND2_X1 U12388 ( .A1(n10097), .A2(n9874), .ZN(n10006) );
  AOI22_X1 U12389 ( .A1(n14238), .A2(n6972), .B1(n10006), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n9875) );
  OAI211_X1 U12390 ( .C1(n10215), .C2(n14215), .A(n9876), .B(n9875), .ZN(
        P1_U3232) );
  NOR2_X1 U12391 ( .A1(n10215), .A2(n14380), .ZN(n10332) );
  OR2_X1 U12392 ( .A1(n11748), .A2(n13822), .ZN(n14523) );
  NAND2_X1 U12393 ( .A1(n13486), .A2(n10329), .ZN(n11445) );
  NAND2_X1 U12394 ( .A1(n11437), .A2(n11445), .ZN(n10333) );
  INV_X1 U12395 ( .A(n10333), .ZN(n11758) );
  AOI21_X1 U12396 ( .B1(n14489), .B2(n14540), .A(n11758), .ZN(n9877) );
  AOI211_X1 U12397 ( .C1(n9878), .C2(n6972), .A(n10332), .B(n9877), .ZN(n9920)
         );
  AND3_X1 U12398 ( .A1(n9917), .A2(n9915), .A3(n9879), .ZN(n9881) );
  AND2_X2 U12399 ( .A1(n9881), .A2(n9918), .ZN(n14563) );
  INV_X1 U12400 ( .A(n14563), .ZN(n14561) );
  NAND2_X1 U12401 ( .A1(n14561), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9882) );
  OAI21_X1 U12402 ( .B1(n9920), .B2(n14561), .A(n9882), .ZN(P1_U3528) );
  INV_X1 U12403 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9899) );
  INV_X1 U12404 ( .A(n9883), .ZN(n10024) );
  NAND2_X1 U12405 ( .A1(n9886), .A2(n10024), .ZN(n9884) );
  NAND2_X1 U12406 ( .A1(n9885), .A2(n9884), .ZN(n13086) );
  INV_X1 U12407 ( .A(n13086), .ZN(n9897) );
  INV_X1 U12408 ( .A(n14689), .ZN(n14709) );
  NAND2_X1 U12409 ( .A1(n13086), .A2(n14709), .ZN(n9893) );
  OAI21_X1 U12410 ( .B1(n9887), .B2(n9886), .A(n10655), .ZN(n9891) );
  NAND2_X1 U12411 ( .A1(n12746), .A2(n13002), .ZN(n9889) );
  NAND2_X1 U12412 ( .A1(n12744), .A2(n13004), .ZN(n9888) );
  NAND2_X1 U12413 ( .A1(n9889), .A2(n9888), .ZN(n9890) );
  AOI21_X1 U12414 ( .B1(n9891), .B2(n13065), .A(n9890), .ZN(n9892) );
  AND2_X1 U12415 ( .A1(n9893), .A2(n9892), .ZN(n13079) );
  NAND2_X1 U12416 ( .A1(n10021), .A2(n10515), .ZN(n9894) );
  NAND2_X1 U12417 ( .A1(n9894), .A2(n6438), .ZN(n9895) );
  NOR2_X1 U12418 ( .A1(n10664), .A2(n9895), .ZN(n13084) );
  AOI21_X1 U12419 ( .B1(n14660), .B2(n10021), .A(n13084), .ZN(n9896) );
  OAI211_X1 U12420 ( .C1(n9897), .C2(n14688), .A(n13079), .B(n9896), .ZN(n9940) );
  NAND2_X1 U12421 ( .A1(n9940), .A2(n14723), .ZN(n9898) );
  OAI21_X1 U12422 ( .B1(n14723), .B2(n9899), .A(n9898), .ZN(P2_U3433) );
  INV_X1 U12423 ( .A(n9900), .ZN(n9977) );
  AOI21_X1 U12424 ( .B1(n9902), .B2(n9901), .A(n9977), .ZN(n9912) );
  NAND2_X1 U12425 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n11088)
         );
  OAI21_X1 U12426 ( .B1(n14624), .B2(n9903), .A(n11088), .ZN(n9904) );
  AOI21_X1 U12427 ( .B1(n14577), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9904), .ZN(
        n9911) );
  MUX2_X1 U12428 ( .A(n9488), .B(P2_REG1_REG_11__SCAN_IN), .S(n9905), .Z(n9906) );
  NAND3_X1 U12429 ( .A1(n12836), .A2(n9907), .A3(n9906), .ZN(n9908) );
  NAND3_X1 U12430 ( .A1(n9909), .A2(n14579), .A3(n9908), .ZN(n9910) );
  OAI211_X1 U12431 ( .C1(n9912), .C2(n14622), .A(n9911), .B(n9910), .ZN(
        P2_U3225) );
  INV_X1 U12432 ( .A(n11018), .ZN(n9923) );
  OAI21_X1 U12433 ( .B1(n9913), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9986) );
  XNOR2_X1 U12434 ( .A(n9986), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11019) );
  INV_X1 U12435 ( .A(n11019), .ZN(n10159) );
  OAI222_X1 U12436 ( .A1(n13986), .A2(n9923), .B1(n10159), .B2(P1_U3086), .C1(
        n9914), .C2(n13988), .ZN(P1_U3343) );
  AND3_X1 U12437 ( .A1(n9917), .A2(n9916), .A3(n9915), .ZN(n9919) );
  OR2_X1 U12438 ( .A1(n9920), .A2(n7230), .ZN(n9921) );
  OAI21_X1 U12439 ( .B1(n14546), .B2(n9561), .A(n9921), .ZN(P1_U3459) );
  INV_X1 U12440 ( .A(n9922), .ZN(n9972) );
  OAI222_X1 U12441 ( .A1(n13201), .A2(n9924), .B1(n13199), .B2(n9923), .C1(
        n9972), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U12442 ( .A(n10003), .ZN(n9927) );
  MUX2_X1 U12443 ( .A(n13365), .B(n9929), .S(n9928), .Z(n9930) );
  OAI21_X1 U12444 ( .B1(n9931), .B2(n9930), .A(n10001), .ZN(n9935) );
  OR2_X1 U12445 ( .A1(n13463), .A2(n14382), .ZN(n14214) );
  INV_X1 U12446 ( .A(n14214), .ZN(n13453) );
  NAND2_X1 U12447 ( .A1(n13453), .A2(n13486), .ZN(n9933) );
  AOI22_X1 U12448 ( .A1(n14238), .A2(n7445), .B1(n10006), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n9932) );
  OAI211_X1 U12449 ( .C1(n6749), .C2(n14215), .A(n9933), .B(n9932), .ZN(n9934)
         );
  AOI21_X1 U12450 ( .B1(n9935), .B2(n14233), .A(n9934), .ZN(n9936) );
  INV_X1 U12451 ( .A(n9936), .ZN(P1_U3222) );
  INV_X1 U12452 ( .A(n12151), .ZN(n14157) );
  INV_X1 U12453 ( .A(n9937), .ZN(n9939) );
  OAI222_X1 U12454 ( .A1(n14157), .A2(P3_U3151), .B1(n12528), .B2(n9939), .C1(
        n9938), .C2(n12530), .ZN(P3_U3278) );
  NAND2_X1 U12455 ( .A1(n9940), .A2(n14737), .ZN(n9941) );
  OAI21_X1 U12456 ( .B1(n14737), .B2(n9459), .A(n9941), .ZN(P2_U3500) );
  INV_X1 U12457 ( .A(n9942), .ZN(n9950) );
  OR2_X1 U12458 ( .A1(n10368), .A2(n9950), .ZN(n9944) );
  OAI21_X1 U12459 ( .B1(n9944), .B2(n14636), .A(n9943), .ZN(n9949) );
  AND3_X1 U12460 ( .A1(n9947), .A2(n9946), .A3(n9945), .ZN(n9948) );
  NAND2_X1 U12461 ( .A1(n9949), .A2(n9948), .ZN(n10034) );
  OR2_X1 U12462 ( .A1(n10034), .A2(P2_U3088), .ZN(n12682) );
  INV_X1 U12463 ( .A(n12682), .ZN(n9966) );
  OR2_X1 U12464 ( .A1(n14636), .A2(n9950), .ZN(n9951) );
  NOR2_X1 U12465 ( .A1(n9952), .A2(n10942), .ZN(n9953) );
  AND2_X1 U12466 ( .A1(n11010), .A2(n9953), .ZN(n10382) );
  NAND2_X1 U12467 ( .A1(n9961), .A2(n10382), .ZN(n9955) );
  INV_X1 U12468 ( .A(n12717), .ZN(n12710) );
  NAND2_X1 U12469 ( .A1(n12745), .A2(n13004), .ZN(n10516) );
  MUX2_X1 U12470 ( .A(n14638), .B(n9957), .S(n6438), .Z(n9962) );
  INV_X1 U12471 ( .A(n9958), .ZN(n9959) );
  AND2_X1 U12472 ( .A1(n14715), .A2(n9959), .ZN(n9960) );
  OAI22_X1 U12473 ( .A1(n12710), .A2(n10516), .B1(n9962), .B2(n12724), .ZN(
        n9963) );
  AOI21_X1 U12474 ( .B1(n10515), .B2(n12722), .A(n9963), .ZN(n9964) );
  OAI21_X1 U12475 ( .B1(n9966), .B2(n9965), .A(n9964), .ZN(P2_U3204) );
  INV_X1 U12476 ( .A(n9967), .ZN(n9968) );
  AOI21_X1 U12477 ( .B1(n9970), .B2(n9969), .A(n9968), .ZN(n9983) );
  NOR2_X1 U12478 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9971), .ZN(n11290) );
  NOR2_X1 U12479 ( .A1(n14624), .A2(n9972), .ZN(n9973) );
  AOI211_X1 U12480 ( .C1(n14577), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n11290), 
        .B(n9973), .ZN(n9982) );
  INV_X1 U12481 ( .A(n9974), .ZN(n9975) );
  NOR3_X1 U12482 ( .A1(n9977), .A2(n9976), .A3(n9975), .ZN(n9980) );
  INV_X1 U12483 ( .A(n9978), .ZN(n9979) );
  OAI21_X1 U12484 ( .B1(n9980), .B2(n9979), .A(n14582), .ZN(n9981) );
  OAI211_X1 U12485 ( .C1(n9983), .C2(n14620), .A(n9982), .B(n9981), .ZN(
        P2_U3226) );
  INV_X1 U12486 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n15027) );
  NAND2_X1 U12487 ( .A1(n11920), .A2(P3_U3897), .ZN(n9984) );
  OAI21_X1 U12488 ( .B1(P3_U3897), .B2(n15027), .A(n9984), .ZN(P3_U3504) );
  INV_X1 U12489 ( .A(n11024), .ZN(n10013) );
  INV_X1 U12490 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U12491 ( .A1(n9986), .A2(n9985), .ZN(n9987) );
  NAND2_X1 U12492 ( .A1(n9987), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9989) );
  INV_X1 U12493 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9988) );
  NAND2_X1 U12494 ( .A1(n9989), .A2(n9988), .ZN(n10077) );
  OR2_X1 U12495 ( .A1(n9989), .A2(n9988), .ZN(n9990) );
  OAI222_X1 U12496 ( .A1(n13986), .A2(n10013), .B1(n10186), .B2(P1_U3086), 
        .C1(n9991), .C2(n13988), .ZN(P1_U3342) );
  AOI22_X1 U12497 ( .A1(n10240), .A2(n13835), .B1(n13865), .B2(n13485), .ZN(
        n14424) );
  NAND2_X1 U12498 ( .A1(n13484), .A2(n13206), .ZN(n9999) );
  INV_X1 U12499 ( .A(n9992), .ZN(n9993) );
  NAND2_X1 U12500 ( .A1(n11743), .A2(n9993), .ZN(n9997) );
  NAND2_X1 U12501 ( .A1(n10107), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U12502 ( .A1(n11556), .A2(n9994), .ZN(n9995) );
  OR2_X1 U12503 ( .A1(n11450), .A2(n13367), .ZN(n9998) );
  NAND2_X1 U12504 ( .A1(n9999), .A2(n9998), .ZN(n10000) );
  XNOR2_X1 U12505 ( .A(n10000), .B(n13365), .ZN(n10114) );
  NAND2_X1 U12506 ( .A1(n10005), .A2(n14233), .ZN(n10008) );
  AOI22_X1 U12507 ( .A1(n14238), .A2(n6748), .B1(n10006), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n10007) );
  OAI211_X1 U12508 ( .C1(n14424), .C2(n13463), .A(n10008), .B(n10007), .ZN(
        P1_U3237) );
  INV_X1 U12509 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n15127) );
  NAND2_X1 U12510 ( .A1(n11952), .A2(P3_U3897), .ZN(n10009) );
  OAI21_X1 U12511 ( .B1(P3_U3897), .B2(n15127), .A(n10009), .ZN(P3_U3508) );
  INV_X1 U12512 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n15037) );
  NAND2_X1 U12513 ( .A1(n10832), .A2(P3_U3897), .ZN(n10010) );
  OAI21_X1 U12514 ( .B1(P3_U3897), .B2(n15037), .A(n10010), .ZN(P3_U3496) );
  INV_X1 U12515 ( .A(n10011), .ZN(n10064) );
  OAI222_X1 U12516 ( .A1(P2_U3088), .A2(n10064), .B1(n13199), .B2(n10013), 
        .C1(n10012), .C2(n13201), .ZN(P2_U3314) );
  INV_X1 U12517 ( .A(n10014), .ZN(n10016) );
  INV_X1 U12518 ( .A(SI_18_), .ZN(n10015) );
  OAI222_X1 U12519 ( .A1(n6811), .A2(P3_U3151), .B1(n12528), .B2(n10016), .C1(
        n10015), .C2(n12530), .ZN(P3_U3277) );
  INV_X1 U12520 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n15040) );
  NAND2_X1 U12521 ( .A1(n11866), .A2(P3_U3897), .ZN(n10017) );
  OAI21_X1 U12522 ( .B1(P3_U3897), .B2(n15040), .A(n10017), .ZN(P3_U3502) );
  OAI222_X1 U12523 ( .A1(n12177), .A2(P3_U3151), .B1(n12528), .B2(n10019), 
        .C1(n10018), .C2(n12521), .ZN(P3_U3276) );
  NAND2_X1 U12524 ( .A1(n12744), .A2(n10022), .ZN(n10028) );
  XNOR2_X1 U12525 ( .A(n12684), .B(n12604), .ZN(n10029) );
  NAND2_X1 U12526 ( .A1(n12745), .A2(n10022), .ZN(n10025) );
  XNOR2_X1 U12527 ( .A(n10026), .B(n10025), .ZN(n12612) );
  NOR2_X1 U12528 ( .A1(n10515), .A2(n12604), .ZN(n10023) );
  INV_X1 U12529 ( .A(n10025), .ZN(n10027) );
  NOR2_X1 U12530 ( .A1(n10027), .A2(n10026), .ZN(n12688) );
  NOR2_X1 U12531 ( .A1(n10420), .A2(n6438), .ZN(n10031) );
  XNOR2_X1 U12532 ( .A(n10383), .B(n12576), .ZN(n10030) );
  NAND2_X1 U12533 ( .A1(n10031), .A2(n10030), .ZN(n10040) );
  OAI21_X1 U12534 ( .B1(n10031), .B2(n10030), .A(n10040), .ZN(n10032) );
  AOI211_X1 U12535 ( .C1(n10033), .C2(n10032), .A(n12724), .B(n10042), .ZN(
        n10039) );
  NOR2_X1 U12536 ( .A1(n12710), .A2(n13055), .ZN(n12683) );
  INV_X1 U12537 ( .A(n10090), .ZN(n12742) );
  AOI22_X1 U12538 ( .A1(n12685), .A2(n12742), .B1(n14651), .B2(n12722), .ZN(
        n10036) );
  AND2_X1 U12539 ( .A1(n10034), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12708) );
  MUX2_X1 U12540 ( .A(n12720), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n10035) );
  OAI211_X1 U12541 ( .C1(n12658), .C2(n10037), .A(n10036), .B(n10035), .ZN(
        n10038) );
  OR2_X1 U12542 ( .A1(n10039), .A2(n10038), .ZN(P2_U3190) );
  INV_X1 U12543 ( .A(n10040), .ZN(n10041) );
  XNOR2_X1 U12544 ( .A(n10431), .B(n6816), .ZN(n10084) );
  NOR2_X1 U12545 ( .A1(n10090), .A2(n6438), .ZN(n10086) );
  XNOR2_X1 U12546 ( .A(n10084), .B(n10086), .ZN(n10043) );
  OAI21_X1 U12547 ( .B1(n10044), .B2(n10043), .A(n10085), .ZN(n10048) );
  INV_X1 U12548 ( .A(n12685), .ZN(n12656) );
  OAI22_X1 U12549 ( .A1(n10420), .A2(n12658), .B1(n12656), .B2(n10438), .ZN(
        n10047) );
  NAND2_X1 U12550 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n12776) );
  NAND2_X1 U12551 ( .A1(n12722), .A2(n14659), .ZN(n10045) );
  OAI211_X1 U12552 ( .C1(n12720), .C2(n10430), .A(n12776), .B(n10045), .ZN(
        n10046) );
  AOI211_X1 U12553 ( .C1(n10048), .C2(n12689), .A(n10047), .B(n10046), .ZN(
        n10049) );
  INV_X1 U12554 ( .A(n10049), .ZN(P2_U3202) );
  INV_X1 U12555 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n11002) );
  NOR2_X1 U12556 ( .A1(n10050), .A2(n10571), .ZN(n13574) );
  MUX2_X1 U12557 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n11002), .S(n13572), .Z(
        n13573) );
  OAI21_X1 U12558 ( .B1(n13575), .B2(n13574), .A(n13573), .ZN(n13577) );
  OAI21_X1 U12559 ( .B1(n10054), .B2(n11002), .A(n13577), .ZN(n10052) );
  INV_X1 U12560 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U12561 ( .A1(n11019), .A2(n10155), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n10159), .ZN(n10051) );
  NOR2_X1 U12562 ( .A1(n10051), .A2(n10052), .ZN(n10154) );
  AOI21_X1 U12563 ( .B1(n10052), .B2(n10051), .A(n10154), .ZN(n10062) );
  AOI21_X1 U12564 ( .B1(n10547), .B2(P1_REG1_REG_10__SCAN_IN), .A(n10053), 
        .ZN(n13568) );
  INV_X1 U12565 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14304) );
  MUX2_X1 U12566 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14304), .S(n13572), .Z(
        n13569) );
  NAND2_X1 U12567 ( .A1(n13568), .A2(n13569), .ZN(n13567) );
  NAND2_X1 U12568 ( .A1(n10054), .A2(n14304), .ZN(n10055) );
  INV_X1 U12569 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10988) );
  MUX2_X1 U12570 ( .A(n10988), .B(P1_REG1_REG_12__SCAN_IN), .S(n11019), .Z(
        n10056) );
  AOI21_X1 U12571 ( .B1(n13567), .B2(n10055), .A(n10056), .ZN(n10158) );
  AND3_X1 U12572 ( .A1(n13567), .A2(n10056), .A3(n10055), .ZN(n10057) );
  OAI21_X1 U12573 ( .B1(n10158), .B2(n10057), .A(n14367), .ZN(n10061) );
  INV_X1 U12574 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n13391) );
  NOR2_X1 U12575 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13391), .ZN(n10059) );
  NOR2_X1 U12576 ( .A1(n14375), .A2(n10159), .ZN(n10058) );
  AOI211_X1 U12577 ( .C1(n14346), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n10059), 
        .B(n10058), .ZN(n10060) );
  OAI211_X1 U12578 ( .C1(n10062), .C2(n14360), .A(n10061), .B(n10060), .ZN(
        P1_U3255) );
  OAI22_X1 U12579 ( .A1(n14624), .A2(n10064), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10063), .ZN(n10068) );
  AOI211_X1 U12580 ( .C1(n10066), .C2(n10065), .A(n14620), .B(n14569), .ZN(
        n10067) );
  AOI211_X1 U12581 ( .C1(n14577), .C2(P2_ADDR_REG_13__SCAN_IN), .A(n10068), 
        .B(n10067), .ZN(n10073) );
  OAI211_X1 U12582 ( .C1(n10071), .C2(n10070), .A(n10069), .B(n14582), .ZN(
        n10072) );
  NAND2_X1 U12583 ( .A1(n10073), .A2(n10072), .ZN(P2_U3227) );
  INV_X1 U12584 ( .A(n11511), .ZN(n10080) );
  NOR2_X1 U12585 ( .A1(n10174), .A2(n13973), .ZN(n10074) );
  MUX2_X1 U12586 ( .A(n13973), .B(n10074), .S(P1_IR_REG_16__SCAN_IN), .Z(
        n10075) );
  NOR2_X1 U12587 ( .A1(n10075), .A2(n10127), .ZN(n13585) );
  INV_X1 U12588 ( .A(n13585), .ZN(n11142) );
  OAI222_X1 U12589 ( .A1(n13986), .A2(n10080), .B1(n11142), .B2(P1_U3086), 
        .C1(n10076), .C2(n13988), .ZN(P1_U3339) );
  INV_X1 U12590 ( .A(n11176), .ZN(n10082) );
  NAND2_X1 U12591 ( .A1(n10077), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10078) );
  XNOR2_X1 U12592 ( .A(n10078), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11177) );
  OAI222_X1 U12593 ( .A1(n13986), .A2(n10082), .B1(n11137), .B2(P1_U3086), 
        .C1(n10079), .C2(n13988), .ZN(P1_U3341) );
  OAI222_X1 U12594 ( .A1(n13201), .A2(n10081), .B1(n13199), .B2(n10080), .C1(
        n14598), .C2(P2_U3088), .ZN(P2_U3311) );
  OAI222_X1 U12595 ( .A1(n13201), .A2(n10083), .B1(n13199), .B2(n10082), .C1(
        n14571), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U12596 ( .A(n12722), .ZN(n12653) );
  NOR2_X1 U12597 ( .A1(n10438), .A2(n6438), .ZN(n10204) );
  XNOR2_X1 U12598 ( .A(n10471), .B(n6816), .ZN(n10203) );
  XOR2_X1 U12599 ( .A(n10204), .B(n10203), .Z(n10088) );
  OAI21_X1 U12600 ( .B1(n10088), .B2(n10087), .A(n10205), .ZN(n10089) );
  NAND2_X1 U12601 ( .A1(n10089), .A2(n12689), .ZN(n10094) );
  OAI22_X1 U12602 ( .A1(n10090), .A2(n13055), .B1(n10453), .B2(n13057), .ZN(
        n10465) );
  NOR2_X1 U12603 ( .A1(n12720), .A2(n10472), .ZN(n10091) );
  AOI211_X1 U12604 ( .C1(n12717), .C2(n10465), .A(n10092), .B(n10091), .ZN(
        n10093) );
  OAI211_X1 U12605 ( .C1(n14670), .C2(n12653), .A(n10094), .B(n10093), .ZN(
        P2_U3199) );
  INV_X1 U12606 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n15061) );
  NAND3_X1 U12607 ( .A1(n10097), .A2(n10096), .A3(n10095), .ZN(n10098) );
  NAND2_X1 U12608 ( .A1(n10098), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10099) );
  INV_X1 U12609 ( .A(n14241), .ZN(n13465) );
  NAND2_X1 U12610 ( .A1(n13484), .A2(n13865), .ZN(n10106) );
  NAND2_X1 U12611 ( .A1(n11726), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n10104) );
  OR2_X1 U12612 ( .A1(n11731), .A2(n9720), .ZN(n10103) );
  XNOR2_X1 U12613 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n10509) );
  OR2_X1 U12614 ( .A1(n11634), .A2(n10509), .ZN(n10102) );
  OR2_X1 U12615 ( .A1(n11730), .A2(n15068), .ZN(n10101) );
  NAND2_X1 U12616 ( .A1(n13483), .A2(n13835), .ZN(n10105) );
  AND2_X1 U12617 ( .A1(n10106), .A2(n10105), .ZN(n14408) );
  AOI22_X1 U12618 ( .A1(n11744), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n11556), 
        .B2(n13524), .ZN(n10110) );
  NAND2_X1 U12619 ( .A1(n10108), .A2(n11743), .ZN(n10109) );
  AOI22_X1 U12620 ( .A1(n14238), .A2(n10243), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10111) );
  OAI21_X1 U12621 ( .B1(n14408), .B2(n13463), .A(n10111), .ZN(n10122) );
  OAI22_X1 U12622 ( .A1(n10221), .A2(n13264), .B1(n14480), .B2(n13367), .ZN(
        n10112) );
  XNOR2_X1 U12623 ( .A(n10112), .B(n13365), .ZN(n10483) );
  OAI22_X1 U12624 ( .A1(n10221), .A2(n13364), .B1(n14480), .B2(n13264), .ZN(
        n10482) );
  XNOR2_X1 U12625 ( .A(n10483), .B(n10482), .ZN(n10120) );
  INV_X1 U12626 ( .A(n10113), .ZN(n10115) );
  AOI211_X1 U12627 ( .C1(n10120), .C2(n10119), .A(n14221), .B(n6478), .ZN(
        n10121) );
  AOI211_X1 U12628 ( .C1(n15061), .C2(n13465), .A(n10122), .B(n10121), .ZN(
        n10123) );
  INV_X1 U12629 ( .A(n10123), .ZN(P1_U3218) );
  INV_X1 U12630 ( .A(n11977), .ZN(n11913) );
  AOI22_X1 U12631 ( .A1(n11979), .A2(n10124), .B1(n11913), .B2(n11996), .ZN(
        n10126) );
  NAND2_X1 U12632 ( .A1(n11373), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10361) );
  NAND2_X1 U12633 ( .A1(n10361), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10125) );
  OAI211_X1 U12634 ( .C1(n11981), .C2(n11798), .A(n10126), .B(n10125), .ZN(
        P3_U3172) );
  INV_X1 U12635 ( .A(n11520), .ZN(n10170) );
  NAND2_X1 U12636 ( .A1(n7295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10128) );
  XNOR2_X1 U12637 ( .A(n10128), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13598) );
  INV_X1 U12638 ( .A(n13598), .ZN(n13593) );
  OAI222_X1 U12639 ( .A1(n13986), .A2(n10170), .B1(n13593), .B2(P1_U3086), 
        .C1(n10129), .C2(n13988), .ZN(P1_U3338) );
  NAND2_X1 U12640 ( .A1(n10130), .A2(n10511), .ZN(n10147) );
  NAND2_X1 U12641 ( .A1(n10132), .A2(n10131), .ZN(n10133) );
  AND2_X1 U12642 ( .A1(n10134), .A2(n10133), .ZN(n10145) );
  NAND2_X1 U12643 ( .A1(n10147), .A2(n10145), .ZN(n10140) );
  MUX2_X1 U12644 ( .A(n11997), .B(n10140), .S(n12531), .Z(n14868) );
  AND2_X1 U12645 ( .A1(P3_U3897), .A2(n12531), .ZN(n14863) );
  MUX2_X1 U12646 ( .A(P3_REG2_REG_0__SCAN_IN), .B(P3_REG1_REG_0__SCAN_IN), .S(
        n14738), .Z(n10135) );
  MUX2_X1 U12647 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n14738), .Z(n10136) );
  NOR2_X1 U12648 ( .A1(n10136), .A2(n6852), .ZN(n10316) );
  AOI21_X1 U12649 ( .B1(n10136), .B2(n6852), .A(n10316), .ZN(n10137) );
  NAND2_X1 U12650 ( .A1(n10137), .A2(n14744), .ZN(n10323) );
  OAI21_X1 U12651 ( .B1(n14744), .B2(n10137), .A(n10323), .ZN(n10152) );
  AOI21_X1 U12652 ( .B1(n10138), .B2(n14932), .A(n10303), .ZN(n10150) );
  OR2_X1 U12653 ( .A1(n10140), .A2(n12168), .ZN(n14741) );
  NAND2_X1 U12654 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n14746), .ZN(n10141) );
  INV_X1 U12655 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n11803) );
  NAND2_X1 U12656 ( .A1(P3_REG1_REG_1__SCAN_IN), .A2(n10143), .ZN(n10308) );
  OAI21_X1 U12657 ( .B1(n10143), .B2(P3_REG1_REG_1__SCAN_IN), .A(n10308), .ZN(
        n10144) );
  NAND2_X1 U12658 ( .A1(n14874), .A2(n10144), .ZN(n10149) );
  INV_X1 U12659 ( .A(n10145), .ZN(n10146) );
  AOI22_X1 U12660 ( .A1(n14871), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10148) );
  OAI211_X1 U12661 ( .C1(n10150), .C2(n14878), .A(n10149), .B(n10148), .ZN(
        n10151) );
  AOI21_X1 U12662 ( .B1(n14863), .B2(n10152), .A(n10151), .ZN(n10153) );
  OAI21_X1 U12663 ( .B1(n6852), .B2(n14868), .A(n10153), .ZN(P3_U3183) );
  AOI21_X1 U12664 ( .B1(n10159), .B2(n10155), .A(n10154), .ZN(n10157) );
  INV_X1 U12665 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U12666 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n11025), .B1(n10186), 
        .B2(n10185), .ZN(n10156) );
  NAND2_X1 U12667 ( .A1(n10156), .A2(n10157), .ZN(n10184) );
  OAI211_X1 U12668 ( .C1(n10157), .C2(n10156), .A(n14370), .B(n10184), .ZN(
        n10165) );
  NAND2_X1 U12669 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13436)
         );
  AOI21_X1 U12670 ( .B1(n10988), .B2(n10159), .A(n10158), .ZN(n10161) );
  INV_X1 U12671 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n11031) );
  MUX2_X1 U12672 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n11031), .S(n11025), .Z(
        n10160) );
  NAND2_X1 U12673 ( .A1(n10161), .A2(n10160), .ZN(n10181) );
  OAI211_X1 U12674 ( .C1(n10161), .C2(n10160), .A(n14367), .B(n10181), .ZN(
        n10162) );
  NAND2_X1 U12675 ( .A1(n13436), .A2(n10162), .ZN(n10163) );
  AOI21_X1 U12676 ( .B1(n14346), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10163), 
        .ZN(n10164) );
  OAI211_X1 U12677 ( .C1(n14375), .C2(n10186), .A(n10165), .B(n10164), .ZN(
        P1_U3256) );
  INV_X1 U12678 ( .A(n10166), .ZN(n10168) );
  OAI222_X1 U12679 ( .A1(n10169), .A2(P3_U3151), .B1(n12528), .B2(n10168), 
        .C1(n10167), .C2(n12521), .ZN(P3_U3275) );
  OAI222_X1 U12680 ( .A1(n13201), .A2(n10171), .B1(n13199), .B2(n10170), .C1(
        n14611), .C2(P2_U3088), .ZN(P2_U3310) );
  INV_X1 U12681 ( .A(n11219), .ZN(n10179) );
  MUX2_X1 U12682 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10172), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n10173) );
  INV_X1 U12683 ( .A(n10173), .ZN(n10175) );
  NOR2_X1 U12684 ( .A1(n10175), .A2(n10174), .ZN(n14356) );
  INV_X1 U12685 ( .A(n14356), .ZN(n11138) );
  OAI222_X1 U12686 ( .A1(n13986), .A2(n10179), .B1(n11138), .B2(P1_U3086), 
        .C1(n10176), .C2(n13988), .ZN(P1_U3340) );
  INV_X1 U12687 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n15093) );
  NAND2_X1 U12688 ( .A1(n11835), .A2(P3_U3897), .ZN(n10177) );
  OAI21_X1 U12689 ( .B1(P3_U3897), .B2(n15093), .A(n10177), .ZN(P3_U3514) );
  OAI222_X1 U12690 ( .A1(P2_U3088), .A2(n10180), .B1(n13199), .B2(n10179), 
        .C1(n10178), .C2(n13201), .ZN(P2_U3312) );
  INV_X1 U12691 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n14291) );
  AOI22_X1 U12692 ( .A1(n11177), .A2(n14291), .B1(P1_REG1_REG_14__SCAN_IN), 
        .B2(n11137), .ZN(n10183) );
  OAI21_X1 U12693 ( .B1(n10186), .B2(n11031), .A(n10181), .ZN(n10182) );
  NOR2_X1 U12694 ( .A1(n10183), .A2(n10182), .ZN(n11136) );
  AOI21_X1 U12695 ( .B1(n10183), .B2(n10182), .A(n11136), .ZN(n10192) );
  INV_X1 U12696 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11128) );
  AOI22_X1 U12697 ( .A1(n11177), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n11128), 
        .B2(n11137), .ZN(n10188) );
  OAI21_X1 U12698 ( .B1(n10186), .B2(n10185), .A(n10184), .ZN(n10187) );
  NAND2_X1 U12699 ( .A1(n10188), .A2(n10187), .ZN(n11127) );
  OAI211_X1 U12700 ( .C1(n10188), .C2(n10187), .A(n14370), .B(n11127), .ZN(
        n10191) );
  INV_X1 U12701 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14027) );
  NAND2_X1 U12702 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14203)
         );
  OAI21_X1 U12703 ( .B1(n14992), .B2(n14027), .A(n14203), .ZN(n10189) );
  AOI21_X1 U12704 ( .B1(n11177), .B2(n14357), .A(n10189), .ZN(n10190) );
  OAI211_X1 U12705 ( .C1(n10192), .C2(n14354), .A(n10191), .B(n10190), .ZN(
        P1_U3257) );
  INV_X1 U12706 ( .A(n10193), .ZN(n10195) );
  OAI222_X1 U12707 ( .A1(n10196), .A2(P3_U3151), .B1(n12528), .B2(n10195), 
        .C1(n10194), .C2(n12521), .ZN(P3_U3274) );
  INV_X1 U12708 ( .A(n10197), .ZN(n10200) );
  OAI22_X1 U12709 ( .A1(n10198), .A2(P3_U3151), .B1(SI_22_), .B2(n12521), .ZN(
        n10199) );
  AOI21_X1 U12710 ( .B1(n10200), .B2(n12515), .A(n10199), .ZN(P3_U3273) );
  XNOR2_X1 U12711 ( .A(n14676), .B(n12576), .ZN(n10202) );
  NOR2_X1 U12712 ( .A1(n10453), .A2(n6438), .ZN(n10201) );
  NAND2_X1 U12713 ( .A1(n10202), .A2(n10201), .ZN(n10529) );
  OAI21_X1 U12714 ( .B1(n10202), .B2(n10201), .A(n10529), .ZN(n10207) );
  AOI211_X1 U12715 ( .C1(n10207), .C2(n10206), .A(n12724), .B(n10530), .ZN(
        n10211) );
  OAI22_X1 U12716 ( .A1(n12658), .A2(n10438), .B1(n14676), .B2(n12653), .ZN(
        n10210) );
  NAND2_X1 U12717 ( .A1(n12685), .A2(n12739), .ZN(n10208) );
  NAND2_X1 U12718 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n12786) );
  OAI211_X1 U12719 ( .C1(n12720), .C2(n10445), .A(n10208), .B(n12786), .ZN(
        n10209) );
  OR3_X1 U12720 ( .A1(n10211), .A2(n10210), .A3(n10209), .ZN(P2_U3211) );
  INV_X1 U12721 ( .A(n10212), .ZN(n10213) );
  NAND2_X1 U12722 ( .A1(n11444), .A2(n10214), .ZN(n10217) );
  NAND2_X1 U12723 ( .A1(n10215), .A2(n9925), .ZN(n10216) );
  NAND2_X1 U12724 ( .A1(n10217), .A2(n10216), .ZN(n14425) );
  NAND2_X1 U12725 ( .A1(n13484), .A2(n11450), .ZN(n10218) );
  NAND2_X1 U12726 ( .A1(n14425), .A2(n10232), .ZN(n10220) );
  NAND2_X1 U12727 ( .A1(n6749), .A2(n11450), .ZN(n10219) );
  NAND2_X1 U12728 ( .A1(n10220), .A2(n10219), .ZN(n14402) );
  NAND2_X1 U12729 ( .A1(n10221), .A2(n10243), .ZN(n11448) );
  NAND2_X1 U12730 ( .A1(n14402), .A2(n14404), .ZN(n10223) );
  NAND2_X1 U12731 ( .A1(n10221), .A2(n14480), .ZN(n10222) );
  NAND2_X1 U12732 ( .A1(n10223), .A2(n10222), .ZN(n10250) );
  NAND2_X1 U12733 ( .A1(n10224), .A2(n11743), .ZN(n10227) );
  AOI22_X1 U12734 ( .A1(n6451), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11556), 
        .B2(n10225), .ZN(n10226) );
  NAND2_X1 U12735 ( .A1(n10227), .A2(n10226), .ZN(n14485) );
  XNOR2_X1 U12736 ( .A(n10250), .B(n11757), .ZN(n14488) );
  INV_X1 U12737 ( .A(n11437), .ZN(n10229) );
  NAND2_X1 U12738 ( .A1(n10229), .A2(n10228), .ZN(n10231) );
  INV_X1 U12739 ( .A(n10232), .ZN(n11441) );
  NAND2_X1 U12740 ( .A1(n14403), .A2(n11448), .ZN(n10281) );
  XNOR2_X1 U12741 ( .A(n10281), .B(n11757), .ZN(n10242) );
  INV_X1 U12742 ( .A(n11634), .ZN(n11621) );
  AOI21_X1 U12743 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10233) );
  AND3_X1 U12744 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n10261) );
  NOR2_X1 U12745 ( .A1(n10233), .A2(n10261), .ZN(n10341) );
  NAND2_X1 U12746 ( .A1(n11621), .A2(n10341), .ZN(n10239) );
  OR2_X1 U12747 ( .A1(n11731), .A2(n10234), .ZN(n10238) );
  INV_X1 U12748 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10235) );
  OR2_X1 U12749 ( .A1(n11044), .A2(n10235), .ZN(n10237) );
  OR2_X1 U12750 ( .A1(n11730), .A2(n14551), .ZN(n10236) );
  AOI22_X1 U12751 ( .A1(n10240), .A2(n13865), .B1(n13835), .B2(n13482), .ZN(
        n10505) );
  INV_X1 U12752 ( .A(n10505), .ZN(n10241) );
  AOI21_X1 U12753 ( .B1(n10242), .B2(n14429), .A(n10241), .ZN(n14486) );
  MUX2_X1 U12754 ( .A(n9720), .B(n14486), .S(n14420), .Z(n10248) );
  INV_X1 U12755 ( .A(n10244), .ZN(n14413) );
  INV_X1 U12756 ( .A(n14485), .ZN(n10245) );
  INV_X1 U12757 ( .A(n10297), .ZN(n10342) );
  AOI211_X1 U12758 ( .C1(n14485), .C2(n14413), .A(n14468), .B(n10342), .ZN(
        n14484) );
  OAI22_X1 U12759 ( .A1(n13876), .A2(n10245), .B1(n14416), .B2(n10509), .ZN(
        n10246) );
  AOI21_X1 U12760 ( .B1(n14484), .B2(n14436), .A(n10246), .ZN(n10247) );
  OAI211_X1 U12761 ( .C1(n13844), .C2(n14488), .A(n10248), .B(n10247), .ZN(
        P1_U3289) );
  INV_X1 U12762 ( .A(n11757), .ZN(n10249) );
  NAND2_X1 U12763 ( .A1(n10250), .A2(n10249), .ZN(n10252) );
  OR2_X1 U12764 ( .A1(n14485), .A2(n13483), .ZN(n10251) );
  NAND2_X1 U12765 ( .A1(n10253), .A2(n11743), .ZN(n10255) );
  AOI22_X1 U12766 ( .A1(n11744), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11556), 
        .B2(n13558), .ZN(n10254) );
  NAND2_X1 U12767 ( .A1(n10255), .A2(n10254), .ZN(n11464) );
  NAND2_X1 U12768 ( .A1(n11464), .A2(n14383), .ZN(n14385) );
  OR2_X1 U12769 ( .A1(n11464), .A2(n14383), .ZN(n10256) );
  NAND2_X1 U12770 ( .A1(n14385), .A2(n10256), .ZN(n11761) );
  INV_X1 U12771 ( .A(n11743), .ZN(n11723) );
  OR2_X1 U12772 ( .A1(n10257), .A2(n11723), .ZN(n10260) );
  AOI22_X1 U12773 ( .A1(n11744), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11556), 
        .B2(n10258), .ZN(n10259) );
  NAND2_X1 U12774 ( .A1(n10260), .A2(n10259), .ZN(n14393) );
  INV_X1 U12775 ( .A(n14393), .ZN(n14499) );
  NAND2_X1 U12776 ( .A1(n11726), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10265) );
  OR2_X1 U12777 ( .A1(n11731), .A2(n9722), .ZN(n10264) );
  NAND2_X1 U12778 ( .A1(n10261), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n10274) );
  OAI21_X1 U12779 ( .B1(n10261), .B2(P1_REG3_REG_6__SCAN_IN), .A(n10274), .ZN(
        n14391) );
  OR2_X1 U12780 ( .A1(n11634), .A2(n14391), .ZN(n10263) );
  OR2_X1 U12781 ( .A1(n6743), .A2(n14553), .ZN(n10262) );
  NAND4_X1 U12782 ( .A1(n10265), .A2(n10264), .A3(n10263), .A4(n10262), .ZN(
        n13481) );
  NAND2_X1 U12783 ( .A1(n14499), .A2(n13481), .ZN(n10266) );
  INV_X1 U12784 ( .A(n13481), .ZN(n10761) );
  NAND2_X1 U12785 ( .A1(n14393), .A2(n10761), .ZN(n10285) );
  NAND2_X1 U12786 ( .A1(n10266), .A2(n10285), .ZN(n14384) );
  OR2_X1 U12787 ( .A1(n14393), .A2(n13481), .ZN(n10267) );
  NAND2_X1 U12788 ( .A1(n10268), .A2(n10267), .ZN(n10409) );
  OR2_X1 U12789 ( .A1(n10269), .A2(n11723), .ZN(n10272) );
  AOI22_X1 U12790 ( .A1(n11744), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11556), 
        .B2(n10270), .ZN(n10271) );
  NAND2_X1 U12791 ( .A1(n11711), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10280) );
  OR2_X1 U12792 ( .A1(n11731), .A2(n10296), .ZN(n10279) );
  AND2_X1 U12793 ( .A1(n10274), .A2(n10273), .ZN(n10275) );
  OR2_X1 U12794 ( .A1(n10275), .A2(n10287), .ZN(n10824) );
  OR2_X1 U12795 ( .A1(n11634), .A2(n10824), .ZN(n10278) );
  INV_X1 U12796 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10276) );
  OR2_X1 U12797 ( .A1(n11044), .A2(n10276), .ZN(n10277) );
  NAND4_X1 U12798 ( .A1(n10280), .A2(n10279), .A3(n10278), .A4(n10277), .ZN(
        n13480) );
  XNOR2_X1 U12799 ( .A(n14506), .B(n13480), .ZN(n11763) );
  XNOR2_X1 U12800 ( .A(n10409), .B(n11763), .ZN(n14510) );
  INV_X1 U12801 ( .A(n13483), .ZN(n10495) );
  NAND2_X1 U12802 ( .A1(n10495), .A2(n14485), .ZN(n10282) );
  INV_X1 U12803 ( .A(n14384), .ZN(n10284) );
  NAND2_X1 U12804 ( .A1(n14388), .A2(n10285), .ZN(n10286) );
  OAI21_X1 U12805 ( .B1(n10286), .B2(n11763), .A(n10388), .ZN(n10295) );
  NAND2_X1 U12806 ( .A1(n13481), .A2(n13865), .ZN(n10294) );
  NAND2_X1 U12807 ( .A1(n11726), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10292) );
  OR2_X1 U12808 ( .A1(n11731), .A2(n9763), .ZN(n10291) );
  NAND2_X1 U12809 ( .A1(n10287), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10399) );
  OR2_X1 U12810 ( .A1(n10287), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10288) );
  NAND2_X1 U12811 ( .A1(n10399), .A2(n10288), .ZN(n11072) );
  OR2_X1 U12812 ( .A1(n11634), .A2(n11072), .ZN(n10290) );
  OR2_X1 U12813 ( .A1(n6743), .A2(n14557), .ZN(n10289) );
  NAND4_X1 U12814 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(n10289), .ZN(
        n13479) );
  NAND2_X1 U12815 ( .A1(n13479), .A2(n13835), .ZN(n10293) );
  NAND2_X1 U12816 ( .A1(n10294), .A2(n10293), .ZN(n10821) );
  AOI21_X1 U12817 ( .B1(n10295), .B2(n14429), .A(n10821), .ZN(n14514) );
  MUX2_X1 U12818 ( .A(n10296), .B(n14514), .S(n14420), .Z(n10302) );
  OR2_X1 U12819 ( .A1(n10297), .A2(n11464), .ZN(n14394) );
  INV_X1 U12820 ( .A(n14506), .ZN(n10299) );
  OAI21_X1 U12821 ( .B1(n14395), .B2(n10299), .A(n14412), .ZN(n10298) );
  AND2_X1 U12822 ( .A1(n14395), .A2(n10299), .ZN(n10411) );
  NOR2_X1 U12823 ( .A1(n10298), .A2(n10411), .ZN(n14508) );
  OAI22_X1 U12824 ( .A1(n10299), .A2(n13876), .B1(n10824), .B2(n14416), .ZN(
        n10300) );
  AOI21_X1 U12825 ( .B1(n14508), .B2(n14436), .A(n10300), .ZN(n10301) );
  OAI211_X1 U12826 ( .C1(n13844), .C2(n14510), .A(n10302), .B(n10301), .ZN(
        P1_U3286) );
  INV_X1 U12827 ( .A(n14868), .ZN(n14828) );
  NOR2_X1 U12828 ( .A1(n10304), .A2(n10303), .ZN(n10306) );
  AOI21_X1 U12829 ( .B1(n10306), .B2(n10305), .A(n10891), .ZN(n10315) );
  INV_X1 U12830 ( .A(n10307), .ZN(n10309) );
  NAND2_X1 U12831 ( .A1(n10309), .A2(n10308), .ZN(n10311) );
  INV_X1 U12832 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15112) );
  XNOR2_X1 U12833 ( .A(n10892), .B(n15112), .ZN(n10310) );
  NAND2_X1 U12834 ( .A1(n10310), .A2(n10311), .ZN(n10838) );
  OAI21_X1 U12835 ( .B1(n10311), .B2(n10310), .A(n10838), .ZN(n10312) );
  NAND2_X1 U12836 ( .A1(n14874), .A2(n10312), .ZN(n10314) );
  AOI22_X1 U12837 ( .A1(n14871), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10313) );
  OAI211_X1 U12838 ( .C1(n10315), .C2(n14878), .A(n10314), .B(n10313), .ZN(
        n10327) );
  INV_X1 U12839 ( .A(n10316), .ZN(n10322) );
  MUX2_X1 U12840 ( .A(n10317), .B(n15112), .S(n14738), .Z(n10318) );
  NAND2_X1 U12841 ( .A1(n10318), .A2(n10839), .ZN(n10850) );
  INV_X1 U12842 ( .A(n10318), .ZN(n10319) );
  NAND2_X1 U12843 ( .A1(n10319), .A2(n10892), .ZN(n10320) );
  NAND2_X1 U12844 ( .A1(n10850), .A2(n10320), .ZN(n10321) );
  INV_X1 U12845 ( .A(n14760), .ZN(n10325) );
  NAND3_X1 U12846 ( .A1(n10323), .A2(n10322), .A3(n10321), .ZN(n10324) );
  INV_X1 U12847 ( .A(n14863), .ZN(n14761) );
  AOI21_X1 U12848 ( .B1(n10325), .B2(n10324), .A(n14761), .ZN(n10326) );
  AOI211_X1 U12849 ( .C1(n14828), .C2(n10839), .A(n10327), .B(n10326), .ZN(
        n10328) );
  INV_X1 U12850 ( .A(n10328), .ZN(P3_U3184) );
  INV_X1 U12851 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n13503) );
  OAI22_X1 U12852 ( .A1(n14420), .A2(n13503), .B1(n9560), .B2(n14416), .ZN(
        n10331) );
  AOI21_X1 U12853 ( .B1(n13857), .B2(n13876), .A(n10329), .ZN(n10330) );
  AOI211_X1 U12854 ( .C1(n10332), .C2(n14420), .A(n10331), .B(n10330), .ZN(
        n10335) );
  NOR2_X1 U12855 ( .A1(n14439), .A2(n14540), .ZN(n13842) );
  OAI21_X1 U12856 ( .B1(n13842), .B2(n14252), .A(n10333), .ZN(n10334) );
  NAND2_X1 U12857 ( .A1(n10335), .A2(n10334), .ZN(P1_U3293) );
  XNOR2_X1 U12858 ( .A(n10336), .B(n7181), .ZN(n14492) );
  OAI21_X1 U12859 ( .B1(n7181), .B2(n10337), .A(n14386), .ZN(n10339) );
  OAI22_X1 U12860 ( .A1(n10495), .A2(n14382), .B1(n10761), .B2(n14380), .ZN(
        n10338) );
  AOI21_X1 U12861 ( .B1(n10339), .B2(n14429), .A(n10338), .ZN(n10340) );
  OAI21_X1 U12862 ( .B1(n14492), .B2(n14509), .A(n10340), .ZN(n14495) );
  NAND2_X1 U12863 ( .A1(n14495), .A2(n14420), .ZN(n10346) );
  INV_X1 U12864 ( .A(n10341), .ZN(n10496) );
  OAI22_X1 U12865 ( .A1(n14420), .A2(n10234), .B1(n10496), .B2(n14416), .ZN(
        n10344) );
  INV_X1 U12866 ( .A(n11464), .ZN(n14494) );
  OAI211_X1 U12867 ( .C1(n10342), .C2(n14494), .A(n14412), .B(n14394), .ZN(
        n14493) );
  NOR2_X1 U12868 ( .A1(n14493), .A2(n13875), .ZN(n10343) );
  AOI211_X1 U12869 ( .C1(n14430), .C2(n11464), .A(n10344), .B(n10343), .ZN(
        n10345) );
  OAI211_X1 U12870 ( .C1(n14492), .C2(n14121), .A(n10346), .B(n10345), .ZN(
        P1_U3288) );
  INV_X1 U12871 ( .A(n14922), .ZN(n10352) );
  NOR3_X1 U12872 ( .A1(n10348), .A2(n10347), .A3(n14917), .ZN(n10350) );
  AOI211_X1 U12873 ( .C1(n10352), .C2(n10351), .A(n10350), .B(n10349), .ZN(
        n10356) );
  AOI22_X1 U12874 ( .A1(n11913), .A2(n14921), .B1(n11940), .B2(n14918), .ZN(
        n10353) );
  OAI21_X1 U12875 ( .B1(n11968), .B2(n14916), .A(n10353), .ZN(n10354) );
  AOI21_X1 U12876 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n10361), .A(n10354), .ZN(
        n10355) );
  OAI21_X1 U12877 ( .B1(n10356), .B2(n11981), .A(n10355), .ZN(P3_U3162) );
  XOR2_X1 U12878 ( .A(n10358), .B(n10357), .Z(n10363) );
  AOI22_X1 U12879 ( .A1(n11913), .A2(n11995), .B1(n11940), .B2(n11996), .ZN(
        n10359) );
  OAI21_X1 U12880 ( .B1(n11968), .B2(n14910), .A(n10359), .ZN(n10360) );
  AOI21_X1 U12881 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10361), .A(n10360), .ZN(
        n10362) );
  OAI21_X1 U12882 ( .B1(n10363), .B2(n11981), .A(n10362), .ZN(P3_U3177) );
  OAI21_X1 U12883 ( .B1(n10365), .B2(n10377), .A(n10364), .ZN(n10366) );
  INV_X1 U12884 ( .A(n10366), .ZN(n14654) );
  INV_X1 U12885 ( .A(n10367), .ZN(n10369) );
  NAND2_X1 U12886 ( .A1(n10369), .A2(n10368), .ZN(n10370) );
  NAND2_X1 U12887 ( .A1(n14689), .A2(n10583), .ZN(n10372) );
  AND2_X1 U12888 ( .A1(n6816), .A2(n10372), .ZN(n10373) );
  NAND3_X1 U12889 ( .A1(n10375), .A2(n10377), .A3(n10376), .ZN(n10378) );
  NAND2_X1 U12890 ( .A1(n10374), .A2(n10378), .ZN(n10379) );
  AOI222_X1 U12891 ( .A1(n13065), .A2(n10379), .B1(n12742), .B2(n13004), .C1(
        n12744), .C2(n13002), .ZN(n14653) );
  MUX2_X1 U12892 ( .A(n10380), .B(n14653), .S(n13038), .Z(n10386) );
  INV_X1 U12893 ( .A(n10429), .ZN(n10381) );
  AOI211_X1 U12894 ( .C1(n14651), .C2(n10663), .A(n10022), .B(n10381), .ZN(
        n14650) );
  OAI22_X1 U12895 ( .A1(n13073), .A2(n10383), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n12998), .ZN(n10384) );
  AOI21_X1 U12896 ( .B1(n14650), .B2(n13085), .A(n10384), .ZN(n10385) );
  OAI211_X1 U12897 ( .C1(n14654), .C2(n13053), .A(n10386), .B(n10385), .ZN(
        P2_U3262) );
  INV_X1 U12898 ( .A(n13480), .ZN(n14381) );
  NAND2_X1 U12899 ( .A1(n14506), .A2(n14381), .ZN(n10387) );
  NAND2_X1 U12900 ( .A1(n10388), .A2(n10387), .ZN(n10395) );
  OR2_X1 U12901 ( .A1(n10389), .A2(n11723), .ZN(n10392) );
  AOI22_X1 U12902 ( .A1(n11744), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11556), 
        .B2(n10390), .ZN(n10391) );
  INV_X1 U12903 ( .A(n13479), .ZN(n10393) );
  OR2_X1 U12904 ( .A1(n14515), .A2(n10393), .ZN(n10539) );
  NAND2_X1 U12905 ( .A1(n14515), .A2(n10393), .ZN(n10394) );
  NAND2_X1 U12906 ( .A1(n10539), .A2(n10394), .ZN(n11762) );
  AOI21_X1 U12907 ( .B1(n10395), .B2(n11762), .A(n14540), .ZN(n10407) );
  INV_X1 U12908 ( .A(n10395), .ZN(n10397) );
  NAND2_X1 U12909 ( .A1(n13480), .A2(n13865), .ZN(n10406) );
  NAND2_X1 U12910 ( .A1(n11726), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10404) );
  OR2_X1 U12911 ( .A1(n11731), .A2(n10608), .ZN(n10403) );
  NAND2_X1 U12912 ( .A1(n10399), .A2(n10398), .ZN(n10400) );
  NAND2_X1 U12913 ( .A1(n10551), .A2(n10400), .ZN(n11267) );
  OR2_X1 U12914 ( .A1(n11634), .A2(n11267), .ZN(n10402) );
  OR2_X1 U12915 ( .A1(n6743), .A2(n14559), .ZN(n10401) );
  NAND4_X1 U12916 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n13478) );
  NAND2_X1 U12917 ( .A1(n13478), .A2(n13835), .ZN(n10405) );
  NAND2_X1 U12918 ( .A1(n10406), .A2(n10405), .ZN(n11075) );
  AOI21_X1 U12919 ( .B1(n10407), .B2(n10540), .A(n11075), .ZN(n14521) );
  MUX2_X1 U12920 ( .A(n9763), .B(n14521), .S(n14420), .Z(n10415) );
  INV_X1 U12921 ( .A(n11763), .ZN(n10408) );
  OR2_X1 U12922 ( .A1(n14506), .A2(n13480), .ZN(n10410) );
  XNOR2_X1 U12923 ( .A(n10576), .B(n11762), .ZN(n14518) );
  INV_X1 U12924 ( .A(n14515), .ZN(n11078) );
  NAND2_X1 U12925 ( .A1(n10411), .A2(n11078), .ZN(n10605) );
  OAI211_X1 U12926 ( .C1(n10411), .C2(n11078), .A(n14412), .B(n10605), .ZN(
        n14517) );
  NOR2_X1 U12927 ( .A1(n14517), .A2(n13875), .ZN(n10413) );
  OAI22_X1 U12928 ( .A1(n11078), .A2(n13876), .B1(n14416), .B2(n11072), .ZN(
        n10412) );
  AOI211_X1 U12929 ( .C1(n14518), .C2(n14252), .A(n10413), .B(n10412), .ZN(
        n10414) );
  NAND2_X1 U12930 ( .A1(n10415), .A2(n10414), .ZN(P1_U3285) );
  OAI21_X1 U12931 ( .B1(n10417), .B2(n10422), .A(n10416), .ZN(n10427) );
  INV_X1 U12932 ( .A(n10427), .ZN(n14663) );
  AND2_X1 U12933 ( .A1(n9186), .A2(n10418), .ZN(n10419) );
  NAND2_X1 U12934 ( .A1(n13038), .A2(n10419), .ZN(n13083) );
  OAI22_X1 U12935 ( .A1(n10438), .A2(n13057), .B1(n10420), .B2(n13055), .ZN(
        n10426) );
  NAND3_X1 U12936 ( .A1(n10374), .A2(n10422), .A3(n10421), .ZN(n10423) );
  AOI21_X1 U12937 ( .B1(n10424), .B2(n10423), .A(n13029), .ZN(n10425) );
  AOI211_X1 U12938 ( .C1(n10427), .C2(n14709), .A(n10426), .B(n10425), .ZN(
        n14662) );
  MUX2_X1 U12939 ( .A(n10428), .B(n14662), .S(n13038), .Z(n10434) );
  AOI211_X1 U12940 ( .C1(n14659), .C2(n10429), .A(n10022), .B(n10468), .ZN(
        n14658) );
  OAI22_X1 U12941 ( .A1(n13073), .A2(n10431), .B1(n10430), .B2(n12998), .ZN(
        n10432) );
  AOI21_X1 U12942 ( .B1(n14658), .B2(n13085), .A(n10432), .ZN(n10433) );
  OAI211_X1 U12943 ( .C1(n14663), .C2(n13083), .A(n10434), .B(n10433), .ZN(
        P2_U3261) );
  XNOR2_X1 U12944 ( .A(n10435), .B(n10437), .ZN(n14674) );
  XNOR2_X1 U12945 ( .A(n10436), .B(n10437), .ZN(n10440) );
  OAI22_X1 U12946 ( .A1(n10438), .A2(n13055), .B1(n10591), .B2(n13057), .ZN(
        n10439) );
  AOI21_X1 U12947 ( .B1(n10440), .B2(n13065), .A(n10439), .ZN(n10441) );
  OAI21_X1 U12948 ( .B1(n14674), .B2(n14689), .A(n10441), .ZN(n14677) );
  INV_X1 U12949 ( .A(n14677), .ZN(n10442) );
  MUX2_X1 U12950 ( .A(n10443), .B(n10442), .S(n13038), .Z(n10449) );
  OAI21_X1 U12951 ( .B1(n10469), .B2(n14676), .A(n6438), .ZN(n10444) );
  OR2_X1 U12952 ( .A1(n10456), .A2(n10444), .ZN(n14675) );
  INV_X1 U12953 ( .A(n14675), .ZN(n10447) );
  OAI22_X1 U12954 ( .A1(n13073), .A2(n14676), .B1(n12998), .B2(n10445), .ZN(
        n10446) );
  AOI21_X1 U12955 ( .B1(n10447), .B2(n13085), .A(n10446), .ZN(n10448) );
  OAI211_X1 U12956 ( .C1(n14674), .C2(n13083), .A(n10449), .B(n10448), .ZN(
        P2_U3259) );
  XNOR2_X1 U12957 ( .A(n10450), .B(n10451), .ZN(n14681) );
  XNOR2_X1 U12958 ( .A(n6783), .B(n10451), .ZN(n10454) );
  OAI22_X1 U12959 ( .A1(n10453), .A2(n13055), .B1(n10741), .B2(n13057), .ZN(
        n10526) );
  AOI21_X1 U12960 ( .B1(n10454), .B2(n13065), .A(n10526), .ZN(n14683) );
  MUX2_X1 U12961 ( .A(n10455), .B(n14683), .S(n13038), .Z(n10461) );
  OAI21_X1 U12962 ( .B1(n10456), .B2(n14684), .A(n6438), .ZN(n10457) );
  OR2_X1 U12963 ( .A1(n10727), .A2(n10457), .ZN(n14682) );
  INV_X1 U12964 ( .A(n14682), .ZN(n10459) );
  OAI22_X1 U12965 ( .A1(n14684), .A2(n13073), .B1(n12998), .B2(n10528), .ZN(
        n10458) );
  AOI21_X1 U12966 ( .B1(n10459), .B2(n13085), .A(n10458), .ZN(n10460) );
  OAI211_X1 U12967 ( .C1(n13053), .C2(n14681), .A(n10461), .B(n10460), .ZN(
        P2_U3258) );
  XNOR2_X1 U12968 ( .A(n10462), .B(n10463), .ZN(n14666) );
  XNOR2_X1 U12969 ( .A(n10464), .B(n10463), .ZN(n10466) );
  AOI21_X1 U12970 ( .B1(n10466), .B2(n13065), .A(n10465), .ZN(n14669) );
  MUX2_X1 U12971 ( .A(n10467), .B(n14669), .S(n13038), .Z(n10475) );
  INV_X1 U12972 ( .A(n10468), .ZN(n10470) );
  AOI211_X1 U12973 ( .C1(n10471), .C2(n10470), .A(n10022), .B(n10469), .ZN(
        n14667) );
  OAI22_X1 U12974 ( .A1(n13073), .A2(n14670), .B1(n12998), .B2(n10472), .ZN(
        n10473) );
  AOI21_X1 U12975 ( .B1(n14667), .B2(n13085), .A(n10473), .ZN(n10474) );
  OAI211_X1 U12976 ( .C1(n13053), .C2(n14666), .A(n10475), .B(n10474), .ZN(
        P2_U3260) );
  INV_X1 U12977 ( .A(n11555), .ZN(n10480) );
  INV_X1 U12978 ( .A(n10476), .ZN(n10477) );
  NAND2_X1 U12979 ( .A1(n10477), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10478) );
  XNOR2_X1 U12980 ( .A(n10478), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13601) );
  INV_X1 U12981 ( .A(n13601), .ZN(n14374) );
  OAI222_X1 U12982 ( .A1(n13988), .A2(n10479), .B1(n13986), .B2(n10480), .C1(
        P1_U3086), .C2(n14374), .ZN(P1_U3337) );
  OAI222_X1 U12983 ( .A1(n13201), .A2(n10481), .B1(n13199), .B2(n10480), .C1(
        P2_U3088), .C2(n14623), .ZN(P2_U3309) );
  NAND2_X1 U12984 ( .A1(n14485), .A2(n6443), .ZN(n10485) );
  NAND2_X1 U12985 ( .A1(n13331), .A2(n13483), .ZN(n10484) );
  NAND2_X1 U12986 ( .A1(n10485), .A2(n10484), .ZN(n10489) );
  AOI22_X1 U12987 ( .A1(n14485), .A2(n7444), .B1(n13483), .B2(n6443), .ZN(
        n10487) );
  XNOR2_X1 U12988 ( .A(n10487), .B(n13365), .ZN(n10503) );
  INV_X1 U12989 ( .A(n10488), .ZN(n10490) );
  AOI22_X1 U12990 ( .A1(n11464), .A2(n7444), .B1(n6443), .B2(n13482), .ZN(
        n10492) );
  XNOR2_X1 U12991 ( .A(n10492), .B(n13365), .ZN(n10757) );
  XNOR2_X1 U12992 ( .A(n10757), .B(n10758), .ZN(n10493) );
  XNOR2_X1 U12993 ( .A(n10759), .B(n10493), .ZN(n10500) );
  INV_X1 U12994 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10494) );
  OAI22_X1 U12995 ( .A1(n14214), .A2(n10495), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10494), .ZN(n10498) );
  OAI22_X1 U12996 ( .A1(n14215), .A2(n10761), .B1(n14241), .B2(n10496), .ZN(
        n10497) );
  AOI211_X1 U12997 ( .C1(n11464), .C2(n14238), .A(n10498), .B(n10497), .ZN(
        n10499) );
  OAI21_X1 U12998 ( .B1(n10500), .B2(n14221), .A(n10499), .ZN(P1_U3227) );
  AOI211_X1 U12999 ( .C1(n10503), .C2(n10502), .A(n14221), .B(n10501), .ZN(
        n10504) );
  INV_X1 U13000 ( .A(n10504), .ZN(n10508) );
  NAND2_X1 U13001 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13532) );
  OAI21_X1 U13002 ( .B1(n10505), .B2(n13463), .A(n13532), .ZN(n10506) );
  AOI21_X1 U13003 ( .B1(n14485), .B2(n14238), .A(n10506), .ZN(n10507) );
  OAI211_X1 U13004 ( .C1(n14241), .C2(n10509), .A(n10508), .B(n10507), .ZN(
        P1_U3230) );
  NAND2_X1 U13005 ( .A1(n10510), .A2(n12515), .ZN(n10512) );
  OAI211_X1 U13006 ( .C1(n10513), .C2(n12521), .A(n10512), .B(n10511), .ZN(
        P3_U3272) );
  AND2_X1 U13007 ( .A1(n10515), .A2(n10514), .ZN(n14641) );
  INV_X1 U13008 ( .A(n14641), .ZN(n10524) );
  INV_X2 U13009 ( .A(n13038), .ZN(n13078) );
  NOR2_X1 U13010 ( .A1(n13083), .A2(n14638), .ZN(n10522) );
  AOI21_X1 U13011 ( .B1(n13029), .B2(n14689), .A(n14638), .ZN(n10518) );
  INV_X1 U13012 ( .A(n10516), .ZN(n10517) );
  NOR2_X1 U13013 ( .A1(n10518), .A2(n10517), .ZN(n14639) );
  INV_X1 U13014 ( .A(n12998), .ZN(n13081) );
  AOI22_X1 U13015 ( .A1(n14641), .A2(n10519), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n13081), .ZN(n10520) );
  AOI21_X1 U13016 ( .B1(n14639), .B2(n10520), .A(n13078), .ZN(n10521) );
  AOI211_X1 U13017 ( .C1(n13078), .C2(P2_REG2_REG_0__SCAN_IN), .A(n10522), .B(
        n10521), .ZN(n10523) );
  OAI21_X1 U13018 ( .B1(n12984), .B2(n10524), .A(n10523), .ZN(P2_U3265) );
  NOR2_X1 U13019 ( .A1(n10525), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12803) );
  AOI21_X1 U13020 ( .B1(n12717), .B2(n10526), .A(n12803), .ZN(n10527) );
  OAI21_X1 U13021 ( .B1(n12720), .B2(n10528), .A(n10527), .ZN(n10536) );
  XNOR2_X1 U13022 ( .A(n14684), .B(n12576), .ZN(n10532) );
  NOR2_X1 U13023 ( .A1(n10591), .A2(n6438), .ZN(n10531) );
  NAND2_X1 U13024 ( .A1(n10532), .A2(n10531), .ZN(n10586) );
  OAI21_X1 U13025 ( .B1(n10532), .B2(n10531), .A(n10586), .ZN(n10533) );
  AOI211_X1 U13026 ( .C1(n10534), .C2(n10533), .A(n12724), .B(n10588), .ZN(
        n10535) );
  AOI211_X1 U13027 ( .C1(n10537), .C2(n12722), .A(n10536), .B(n10535), .ZN(
        n10538) );
  INV_X1 U13028 ( .A(n10538), .ZN(P2_U3185) );
  NAND2_X1 U13029 ( .A1(n10541), .A2(n11743), .ZN(n10544) );
  AOI22_X1 U13030 ( .A1(n11744), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11556), 
        .B2(n10542), .ZN(n10543) );
  XNOR2_X1 U13031 ( .A(n14525), .B(n11346), .ZN(n11766) );
  NAND2_X1 U13032 ( .A1(n14525), .A2(n11346), .ZN(n10545) );
  OR2_X1 U13033 ( .A1(n10546), .A2(n11723), .ZN(n10549) );
  AOI22_X1 U13034 ( .A1(n6451), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n10547), 
        .B2(n11556), .ZN(n10548) );
  NAND2_X1 U13035 ( .A1(n11726), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10557) );
  OR2_X1 U13036 ( .A1(n11731), .A2(n10571), .ZN(n10556) );
  INV_X1 U13037 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n10550) );
  NAND2_X1 U13038 ( .A1(n10551), .A2(n10550), .ZN(n10552) );
  NAND2_X1 U13039 ( .A1(n10563), .A2(n10552), .ZN(n11345) );
  OR2_X1 U13040 ( .A1(n11634), .A2(n11345), .ZN(n10555) );
  OR2_X1 U13041 ( .A1(n6743), .A2(n10553), .ZN(n10554) );
  NAND4_X1 U13042 ( .A1(n10557), .A2(n10556), .A3(n10555), .A4(n10554), .ZN(
        n13477) );
  INV_X1 U13043 ( .A(n13477), .ZN(n14213) );
  OR2_X1 U13044 ( .A1(n14537), .A2(n14213), .ZN(n10993) );
  NAND2_X1 U13045 ( .A1(n14537), .A2(n14213), .ZN(n10558) );
  NAND2_X1 U13046 ( .A1(n10993), .A2(n10558), .ZN(n11768) );
  OAI21_X1 U13047 ( .B1(n10559), .B2(n7184), .A(n10994), .ZN(n14541) );
  INV_X1 U13048 ( .A(n13842), .ZN(n10581) );
  OR2_X2 U13049 ( .A1(n14525), .A2(n10605), .ZN(n10607) );
  NAND2_X1 U13050 ( .A1(n14537), .A2(n10607), .ZN(n10560) );
  NAND2_X1 U13051 ( .A1(n10560), .A2(n14412), .ZN(n10561) );
  OR2_X1 U13052 ( .A1(n11001), .A2(n10561), .ZN(n10570) );
  NAND2_X1 U13053 ( .A1(n11726), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10568) );
  INV_X1 U13054 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10562) );
  AND2_X1 U13055 ( .A1(n10563), .A2(n10562), .ZN(n10564) );
  OR2_X1 U13056 ( .A1(n10564), .A2(n10986), .ZN(n14229) );
  OR2_X1 U13057 ( .A1(n11634), .A2(n14229), .ZN(n10567) );
  OR2_X1 U13058 ( .A1(n11731), .A2(n11002), .ZN(n10566) );
  OR2_X1 U13059 ( .A1(n6743), .A2(n14304), .ZN(n10565) );
  NAND4_X1 U13060 ( .A1(n10568), .A2(n10567), .A3(n10566), .A4(n10565), .ZN(
        n13476) );
  NAND2_X1 U13061 ( .A1(n13476), .A2(n13835), .ZN(n10569) );
  NAND2_X1 U13062 ( .A1(n10570), .A2(n10569), .ZN(n14535) );
  INV_X1 U13063 ( .A(n14537), .ZN(n10574) );
  NOR2_X1 U13064 ( .A1(n11346), .A2(n14382), .ZN(n14536) );
  OAI22_X1 U13065 ( .A1(n14420), .A2(n10571), .B1(n11345), .B2(n14416), .ZN(
        n10572) );
  AOI21_X1 U13066 ( .B1(n14536), .B2(n14420), .A(n10572), .ZN(n10573) );
  OAI21_X1 U13067 ( .B1(n10574), .B2(n13876), .A(n10573), .ZN(n10575) );
  AOI21_X1 U13068 ( .B1(n14535), .B2(n14436), .A(n10575), .ZN(n10580) );
  NAND2_X1 U13069 ( .A1(n10600), .A2(n11766), .ZN(n10578) );
  OR2_X1 U13070 ( .A1(n14525), .A2(n13478), .ZN(n10577) );
  NAND2_X1 U13071 ( .A1(n10578), .A2(n10577), .ZN(n10999) );
  XNOR2_X1 U13072 ( .A(n10999), .B(n11768), .ZN(n14543) );
  NAND2_X1 U13073 ( .A1(n14543), .A2(n14252), .ZN(n10579) );
  OAI211_X1 U13074 ( .C1(n14541), .C2(n10581), .A(n10580), .B(n10579), .ZN(
        P1_U3283) );
  INV_X1 U13075 ( .A(n11533), .ZN(n10584) );
  OAI222_X1 U13076 ( .A1(n13988), .A2(n10582), .B1(n13986), .B2(n10584), .C1(
        n13822), .C2(P1_U3086), .ZN(P1_U3336) );
  OAI222_X1 U13077 ( .A1(n13201), .A2(n10585), .B1(n13199), .B2(n10584), .C1(
        P2_U3088), .C2(n10583), .ZN(P2_U3308) );
  INV_X1 U13078 ( .A(n10586), .ZN(n10587) );
  NOR2_X1 U13079 ( .A1(n10741), .A2(n6438), .ZN(n10790) );
  XNOR2_X1 U13080 ( .A(n10788), .B(n10790), .ZN(n10589) );
  OAI21_X1 U13081 ( .B1(n10590), .B2(n10589), .A(n10789), .ZN(n10598) );
  OR2_X1 U13082 ( .A1(n10591), .A2(n13055), .ZN(n10593) );
  NAND2_X1 U13083 ( .A1(n12736), .A2(n13004), .ZN(n10592) );
  NAND2_X1 U13084 ( .A1(n10593), .A2(n10592), .ZN(n10720) );
  AND2_X1 U13085 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n12818) );
  AOI21_X1 U13086 ( .B1(n12717), .B2(n10720), .A(n12818), .ZN(n10596) );
  INV_X1 U13087 ( .A(n10728), .ZN(n10594) );
  NAND2_X1 U13088 ( .A1(n12708), .A2(n10594), .ZN(n10595) );
  OAI211_X1 U13089 ( .C1(n14692), .C2(n12653), .A(n10596), .B(n10595), .ZN(
        n10597) );
  AOI21_X1 U13090 ( .B1(n10598), .B2(n12689), .A(n10597), .ZN(n10599) );
  INV_X1 U13091 ( .A(n10599), .ZN(P2_U3193) );
  XOR2_X1 U13092 ( .A(n11766), .B(n10600), .Z(n14524) );
  OAI21_X1 U13093 ( .B1(n6579), .B2(n6965), .A(n10601), .ZN(n10604) );
  NAND2_X1 U13094 ( .A1(n13479), .A2(n13865), .ZN(n10603) );
  NAND2_X1 U13095 ( .A1(n13477), .A2(n13835), .ZN(n10602) );
  NAND2_X1 U13096 ( .A1(n10603), .A2(n10602), .ZN(n11264) );
  AOI21_X1 U13097 ( .B1(n10604), .B2(n14429), .A(n11264), .ZN(n14527) );
  INV_X1 U13098 ( .A(n14527), .ZN(n10612) );
  NAND2_X1 U13099 ( .A1(n14525), .A2(n10605), .ZN(n10606) );
  NAND3_X1 U13100 ( .A1(n10607), .A2(n14412), .A3(n10606), .ZN(n14526) );
  OAI22_X1 U13101 ( .A1(n14420), .A2(n10608), .B1(n11267), .B2(n14416), .ZN(
        n10609) );
  AOI21_X1 U13102 ( .B1(n14525), .B2(n14430), .A(n10609), .ZN(n10610) );
  OAI21_X1 U13103 ( .B1(n14526), .B2(n13875), .A(n10610), .ZN(n10611) );
  AOI21_X1 U13104 ( .B1(n10612), .B2(n14420), .A(n10611), .ZN(n10613) );
  OAI21_X1 U13105 ( .B1(n13844), .B2(n14524), .A(n10613), .ZN(P1_U3284) );
  XNOR2_X1 U13106 ( .A(n10614), .B(n10616), .ZN(n14952) );
  NAND2_X1 U13107 ( .A1(n14952), .A2(n14906), .ZN(n10621) );
  NAND2_X1 U13108 ( .A1(n10615), .A2(n10616), .ZN(n10617) );
  NAND2_X1 U13109 ( .A1(n10952), .A2(n10617), .ZN(n10619) );
  OAI22_X1 U13110 ( .A1(n10707), .A2(n14903), .B1(n10920), .B2(n14901), .ZN(
        n10618) );
  AOI21_X1 U13111 ( .B1(n10619), .B2(n14923), .A(n10618), .ZN(n10620) );
  AND2_X1 U13112 ( .A1(n10621), .A2(n10620), .ZN(n14954) );
  NAND2_X1 U13113 ( .A1(n12512), .A2(n10622), .ZN(n10623) );
  OAI21_X1 U13114 ( .B1(n12512), .B2(n10624), .A(n10623), .ZN(n10625) );
  INV_X1 U13115 ( .A(n10625), .ZN(n10626) );
  NAND2_X1 U13116 ( .A1(n10627), .A2(n10626), .ZN(n10629) );
  AND2_X1 U13117 ( .A1(n14911), .A2(n10628), .ZN(n14893) );
  NAND2_X1 U13118 ( .A1(n14933), .A2(n14893), .ZN(n11244) );
  INV_X1 U13119 ( .A(n11244), .ZN(n14930) );
  OR2_X1 U13120 ( .A1(n10629), .A2(n14911), .ZN(n11253) );
  INV_X1 U13121 ( .A(n11253), .ZN(n14896) );
  AND2_X1 U13122 ( .A1(n10630), .A2(n14960), .ZN(n14951) );
  AOI22_X1 U13123 ( .A1(n14896), .A2(n14951), .B1(n14929), .B2(n10811), .ZN(
        n10631) );
  OAI21_X1 U13124 ( .B1(n10862), .B2(n14933), .A(n10631), .ZN(n10632) );
  AOI21_X1 U13125 ( .B1(n14952), .B2(n14930), .A(n10632), .ZN(n10633) );
  OAI21_X1 U13126 ( .B1(n14954), .B2(n14935), .A(n10633), .ZN(P3_U3228) );
  INV_X1 U13127 ( .A(n11974), .ZN(n11916) );
  NAND2_X1 U13128 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n14766) );
  OAI21_X1 U13129 ( .B1(n11916), .B2(n10708), .A(n14766), .ZN(n10634) );
  AOI21_X1 U13130 ( .B1(n11913), .B2(n11994), .A(n10634), .ZN(n10635) );
  OAI21_X1 U13131 ( .B1(n11968), .B2(n10636), .A(n10635), .ZN(n10641) );
  AOI211_X1 U13132 ( .C1(n10639), .C2(n10638), .A(n11981), .B(n10637), .ZN(
        n10640) );
  AOI211_X1 U13133 ( .C1(n10642), .C2(n11972), .A(n10641), .B(n10640), .ZN(
        n10643) );
  INV_X1 U13134 ( .A(n10643), .ZN(P3_U3158) );
  XNOR2_X1 U13135 ( .A(n10645), .B(n10644), .ZN(n14950) );
  INV_X1 U13136 ( .A(n14950), .ZN(n10653) );
  XNOR2_X1 U13137 ( .A(n10647), .B(n10646), .ZN(n10649) );
  AOI22_X1 U13138 ( .A1(n14920), .A2(n10832), .B1(n11995), .B2(n14919), .ZN(
        n10648) );
  OAI21_X1 U13139 ( .B1(n10649), .B2(n14891), .A(n10648), .ZN(n10650) );
  AOI21_X1 U13140 ( .B1(n14950), .B2(n14906), .A(n10650), .ZN(n14947) );
  MUX2_X1 U13141 ( .A(n10896), .B(n14947), .S(n14933), .Z(n10652) );
  AND2_X1 U13142 ( .A1(n10695), .A2(n14960), .ZN(n14949) );
  AOI22_X1 U13143 ( .A1(n14896), .A2(n14949), .B1(n14929), .B2(n10688), .ZN(
        n10651) );
  OAI211_X1 U13144 ( .C1(n10653), .C2(n11244), .A(n10652), .B(n10651), .ZN(
        P3_U3229) );
  NAND3_X1 U13145 ( .A1(n10661), .A2(n10655), .A3(n10654), .ZN(n10656) );
  NAND2_X1 U13146 ( .A1(n10656), .A2(n10375), .ZN(n10657) );
  NAND2_X1 U13147 ( .A1(n10657), .A2(n13065), .ZN(n10659) );
  AOI22_X1 U13148 ( .A1(n12743), .A2(n13004), .B1(n13002), .B2(n12745), .ZN(
        n10658) );
  NAND2_X1 U13149 ( .A1(n10659), .A2(n10658), .ZN(n14646) );
  INV_X1 U13150 ( .A(n14646), .ZN(n10669) );
  INV_X1 U13151 ( .A(n13053), .ZN(n12988) );
  OAI21_X1 U13152 ( .B1(n10662), .B2(n10661), .A(n10660), .ZN(n14648) );
  OAI211_X1 U13153 ( .C1(n10664), .C2(n14645), .A(n6438), .B(n10663), .ZN(
        n14644) );
  OAI22_X1 U13154 ( .A1(n13038), .A2(n9422), .B1(n12760), .B2(n12998), .ZN(
        n10665) );
  AOI21_X1 U13155 ( .B1(n13082), .B2(n12684), .A(n10665), .ZN(n10666) );
  OAI21_X1 U13156 ( .B1(n12984), .B2(n14644), .A(n10666), .ZN(n10667) );
  AOI21_X1 U13157 ( .B1(n12988), .B2(n14648), .A(n10667), .ZN(n10668) );
  OAI21_X1 U13158 ( .B1(n13078), .B2(n10669), .A(n10668), .ZN(P2_U3263) );
  OAI211_X1 U13159 ( .C1(n10671), .C2(n10670), .A(n10768), .B(n13065), .ZN(
        n10675) );
  OR2_X1 U13160 ( .A1(n11288), .A2(n13057), .ZN(n10673) );
  NAND2_X1 U13161 ( .A1(n12736), .A2(n13002), .ZN(n10672) );
  NAND2_X1 U13162 ( .A1(n10673), .A2(n10672), .ZN(n10939) );
  INV_X1 U13163 ( .A(n10939), .ZN(n10674) );
  NAND2_X1 U13164 ( .A1(n10675), .A2(n10674), .ZN(n14708) );
  INV_X1 U13165 ( .A(n14708), .ZN(n10687) );
  OR2_X1 U13166 ( .A1(n10677), .A2(n10676), .ZN(n10678) );
  AND2_X1 U13167 ( .A1(n10679), .A2(n10678), .ZN(n14710) );
  NAND2_X1 U13168 ( .A1(n10933), .A2(n10750), .ZN(n10680) );
  NAND2_X1 U13169 ( .A1(n10680), .A2(n6438), .ZN(n10681) );
  OR2_X1 U13170 ( .A1(n10681), .A2(n10779), .ZN(n14704) );
  OAI22_X1 U13171 ( .A1(n13038), .A2(n10682), .B1(n10937), .B2(n12998), .ZN(
        n10683) );
  AOI21_X1 U13172 ( .B1(n10933), .B2(n13082), .A(n10683), .ZN(n10684) );
  OAI21_X1 U13173 ( .B1(n14704), .B2(n12984), .A(n10684), .ZN(n10685) );
  AOI21_X1 U13174 ( .B1(n14710), .B2(n12988), .A(n10685), .ZN(n10686) );
  OAI21_X1 U13175 ( .B1(n13078), .B2(n10687), .A(n10686), .ZN(P2_U3255) );
  INV_X1 U13176 ( .A(n10688), .ZN(n10698) );
  NAND2_X1 U13177 ( .A1(n10691), .A2(n11963), .ZN(n10697) );
  NOR2_X1 U13178 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10692), .ZN(n14777) );
  AOI21_X1 U13179 ( .B1(n11940), .B2(n11995), .A(n14777), .ZN(n10693) );
  OAI21_X1 U13180 ( .B1(n10948), .B2(n11977), .A(n10693), .ZN(n10694) );
  AOI21_X1 U13181 ( .B1(n11979), .B2(n10695), .A(n10694), .ZN(n10696) );
  OAI211_X1 U13182 ( .C1(n10698), .C2(n11373), .A(n10697), .B(n10696), .ZN(
        P3_U3170) );
  OR2_X1 U13183 ( .A1(n10700), .A2(n10699), .ZN(n10701) );
  NAND2_X1 U13184 ( .A1(n10702), .A2(n10701), .ZN(n14946) );
  NAND2_X1 U13185 ( .A1(n10703), .A2(n14960), .ZN(n14943) );
  OAI22_X1 U13186 ( .A1(n11253), .A2(n14943), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(n12271), .ZN(n10715) );
  NAND2_X1 U13187 ( .A1(n10704), .A2(n14923), .ZN(n10713) );
  AOI21_X1 U13188 ( .B1(n14899), .B2(n10706), .A(n10705), .ZN(n10712) );
  NAND2_X1 U13189 ( .A1(n14946), .A2(n14906), .ZN(n10711) );
  OAI22_X1 U13190 ( .A1(n10708), .A2(n14903), .B1(n10707), .B2(n14901), .ZN(
        n10709) );
  INV_X1 U13191 ( .A(n10709), .ZN(n10710) );
  OAI211_X1 U13192 ( .C1(n10713), .C2(n10712), .A(n10711), .B(n10710), .ZN(
        n14944) );
  MUX2_X1 U13193 ( .A(n14944), .B(P3_REG2_REG_3__SCAN_IN), .S(n14935), .Z(
        n10714) );
  AOI211_X1 U13194 ( .C1(n14930), .C2(n14946), .A(n10715), .B(n10714), .ZN(
        n10716) );
  INV_X1 U13195 ( .A(n10716), .ZN(P3_U3230) );
  XNOR2_X1 U13196 ( .A(n10717), .B(n10718), .ZN(n10719) );
  NAND2_X1 U13197 ( .A1(n10719), .A2(n13065), .ZN(n10722) );
  INV_X1 U13198 ( .A(n10720), .ZN(n10721) );
  NAND2_X1 U13199 ( .A1(n10722), .A2(n10721), .ZN(n14695) );
  INV_X1 U13200 ( .A(n14695), .ZN(n10736) );
  NAND2_X1 U13201 ( .A1(n10724), .A2(n10723), .ZN(n10725) );
  NAND2_X1 U13202 ( .A1(n10726), .A2(n10725), .ZN(n14690) );
  INV_X1 U13203 ( .A(n14690), .ZN(n10734) );
  OAI211_X1 U13204 ( .C1(n10727), .C2(n14692), .A(n6438), .B(n10748), .ZN(
        n14691) );
  OAI22_X1 U13205 ( .A1(n13038), .A2(n10729), .B1(n10728), .B2(n12998), .ZN(
        n10730) );
  AOI21_X1 U13206 ( .B1(n10731), .B2(n13082), .A(n10730), .ZN(n10732) );
  OAI21_X1 U13207 ( .B1(n14691), .B2(n12984), .A(n10732), .ZN(n10733) );
  AOI21_X1 U13208 ( .B1(n10734), .B2(n12988), .A(n10733), .ZN(n10735) );
  OAI21_X1 U13209 ( .B1(n13078), .B2(n10736), .A(n10735), .ZN(P2_U3257) );
  NAND2_X1 U13210 ( .A1(n10737), .A2(n10744), .ZN(n10738) );
  NAND3_X1 U13211 ( .A1(n10739), .A2(n13065), .A3(n10738), .ZN(n10743) );
  NAND2_X1 U13212 ( .A1(n12735), .A2(n13004), .ZN(n10740) );
  OAI21_X1 U13213 ( .B1(n10741), .B2(n13055), .A(n10740), .ZN(n10794) );
  INV_X1 U13214 ( .A(n10794), .ZN(n10742) );
  NAND2_X1 U13215 ( .A1(n10743), .A2(n10742), .ZN(n14699) );
  INV_X1 U13216 ( .A(n14699), .ZN(n10756) );
  OR2_X1 U13217 ( .A1(n10745), .A2(n10744), .ZN(n10746) );
  AND2_X1 U13218 ( .A1(n10747), .A2(n10746), .ZN(n14700) );
  NAND2_X1 U13219 ( .A1(n10748), .A2(n10793), .ZN(n10749) );
  NAND3_X1 U13220 ( .A1(n10750), .A2(n6438), .A3(n10749), .ZN(n14697) );
  OAI22_X1 U13221 ( .A1(n13038), .A2(n10751), .B1(n10797), .B2(n12998), .ZN(
        n10752) );
  AOI21_X1 U13222 ( .B1(n10793), .B2(n13082), .A(n10752), .ZN(n10753) );
  OAI21_X1 U13223 ( .B1(n14697), .B2(n12984), .A(n10753), .ZN(n10754) );
  AOI21_X1 U13224 ( .B1(n14700), .B2(n12988), .A(n10754), .ZN(n10755) );
  OAI21_X1 U13225 ( .B1(n13078), .B2(n10756), .A(n10755), .ZN(P2_U3256) );
  AND2_X1 U13226 ( .A1(n13331), .A2(n13481), .ZN(n10760) );
  AOI21_X1 U13227 ( .B1(n14393), .B2(n6443), .A(n10760), .ZN(n10816) );
  OAI22_X1 U13228 ( .A1(n14499), .A2(n13367), .B1(n10761), .B2(n13264), .ZN(
        n10762) );
  XNOR2_X1 U13229 ( .A(n10762), .B(n13365), .ZN(n10814) );
  XOR2_X1 U13230 ( .A(n10816), .B(n10814), .Z(n10817) );
  XNOR2_X1 U13231 ( .A(n10818), .B(n10817), .ZN(n10767) );
  OAI21_X1 U13232 ( .B1(n14215), .B2(n14381), .A(n10763), .ZN(n10765) );
  OAI22_X1 U13233 ( .A1(n14214), .A2(n14383), .B1(n14241), .B2(n14391), .ZN(
        n10764) );
  AOI211_X1 U13234 ( .C1(n14393), .C2(n14238), .A(n10765), .B(n10764), .ZN(
        n10766) );
  OAI21_X1 U13235 ( .B1(n10767), .B2(n14221), .A(n10766), .ZN(P1_U3239) );
  INV_X1 U13236 ( .A(n10768), .ZN(n10770) );
  OAI21_X1 U13237 ( .B1(n10770), .B2(n10769), .A(n10776), .ZN(n10772) );
  AOI21_X1 U13238 ( .B1(n10772), .B2(n10771), .A(n13029), .ZN(n10774) );
  OAI22_X1 U13239 ( .A1(n10773), .A2(n13055), .B1(n11317), .B2(n13057), .ZN(
        n11086) );
  INV_X1 U13240 ( .A(n14717), .ZN(n10786) );
  OAI21_X1 U13241 ( .B1(n10777), .B2(n10776), .A(n10775), .ZN(n10778) );
  INV_X1 U13242 ( .A(n10778), .ZN(n14720) );
  NOR2_X1 U13243 ( .A1(n14716), .A2(n10779), .ZN(n10780) );
  OR3_X1 U13244 ( .A1(n10971), .A2(n10780), .A3(n10022), .ZN(n14714) );
  OAI22_X1 U13245 ( .A1(n13038), .A2(n10781), .B1(n11089), .B2(n12998), .ZN(
        n10782) );
  AOI21_X1 U13246 ( .B1(n11091), .B2(n13082), .A(n10782), .ZN(n10783) );
  OAI21_X1 U13247 ( .B1(n14714), .B2(n12984), .A(n10783), .ZN(n10784) );
  AOI21_X1 U13248 ( .B1(n14720), .B2(n12988), .A(n10784), .ZN(n10785) );
  OAI21_X1 U13249 ( .B1(n13078), .B2(n10786), .A(n10785), .ZN(P2_U3254) );
  NOR2_X1 U13250 ( .A1(n10787), .A2(n6438), .ZN(n10929) );
  XNOR2_X1 U13251 ( .A(n10793), .B(n6816), .ZN(n10930) );
  XOR2_X1 U13252 ( .A(n10929), .B(n10930), .Z(n10792) );
  OAI21_X1 U13253 ( .B1(n10792), .B2(n10791), .A(n10932), .ZN(n10799) );
  NAND2_X1 U13254 ( .A1(n10793), .A2(n12722), .ZN(n10796) );
  AOI22_X1 U13255 ( .A1(n12717), .A2(n10794), .B1(P2_REG3_REG_9__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10795) );
  OAI211_X1 U13256 ( .C1(n12720), .C2(n10797), .A(n10796), .B(n10795), .ZN(
        n10798) );
  AOI21_X1 U13257 ( .B1(n10799), .B2(n12689), .A(n10798), .ZN(n10800) );
  INV_X1 U13258 ( .A(n10800), .ZN(P2_U3203) );
  INV_X1 U13259 ( .A(n10801), .ZN(n10803) );
  OAI222_X1 U13260 ( .A1(P3_U3151), .A2(n10804), .B1(n12528), .B2(n10803), 
        .C1(n10802), .C2(n12530), .ZN(P3_U3271) );
  XOR2_X1 U13261 ( .A(n10806), .B(n10805), .Z(n10813) );
  AND2_X1 U13262 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n14795) );
  NOR2_X1 U13263 ( .A1(n11977), .A2(n10920), .ZN(n10807) );
  AOI211_X1 U13264 ( .C1(n11940), .C2(n11994), .A(n14795), .B(n10807), .ZN(
        n10808) );
  OAI21_X1 U13265 ( .B1(n11968), .B2(n10809), .A(n10808), .ZN(n10810) );
  AOI21_X1 U13266 ( .B1(n10811), .B2(n11972), .A(n10810), .ZN(n10812) );
  OAI21_X1 U13267 ( .B1(n10813), .B2(n11981), .A(n10812), .ZN(P3_U3167) );
  INV_X1 U13268 ( .A(n10814), .ZN(n10815) );
  AND2_X1 U13269 ( .A1(n13331), .A2(n13480), .ZN(n10819) );
  AOI21_X1 U13270 ( .B1(n14506), .B2(n6443), .A(n10819), .ZN(n11057) );
  AOI22_X1 U13271 ( .A1(n14506), .A2(n7444), .B1(n6443), .B2(n13480), .ZN(
        n10820) );
  XNOR2_X1 U13272 ( .A(n10820), .B(n13365), .ZN(n11058) );
  XOR2_X1 U13273 ( .A(n11057), .B(n11058), .Z(n11061) );
  XNOR2_X1 U13274 ( .A(n11062), .B(n11061), .ZN(n10827) );
  INV_X1 U13275 ( .A(n13463), .ZN(n14235) );
  NAND2_X1 U13276 ( .A1(n14235), .A2(n10821), .ZN(n10823) );
  OAI211_X1 U13277 ( .C1(n14241), .C2(n10824), .A(n10823), .B(n10822), .ZN(
        n10825) );
  AOI21_X1 U13278 ( .B1(n14506), .B2(n14238), .A(n10825), .ZN(n10826) );
  OAI21_X1 U13279 ( .B1(n10827), .B2(n14221), .A(n10826), .ZN(P1_U3213) );
  INV_X1 U13280 ( .A(n10959), .ZN(n10837) );
  OAI211_X1 U13281 ( .C1(n10830), .C2(n10829), .A(n10828), .B(n11963), .ZN(
        n10836) );
  INV_X1 U13282 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10831) );
  NOR2_X1 U13283 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10831), .ZN(n14811) );
  AOI21_X1 U13284 ( .B1(n11974), .B2(n10832), .A(n14811), .ZN(n10833) );
  OAI21_X1 U13285 ( .B1(n10947), .B2(n11977), .A(n10833), .ZN(n10834) );
  AOI21_X1 U13286 ( .B1(n11979), .B2(n10958), .A(n10834), .ZN(n10835) );
  OAI211_X1 U13287 ( .C1(n10837), .C2(n11373), .A(n10836), .B(n10835), .ZN(
        P3_U3179) );
  INV_X1 U13288 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n14988) );
  MUX2_X1 U13289 ( .A(P3_REG1_REG_10__SCAN_IN), .B(n14988), .S(n11098), .Z(
        n10849) );
  INV_X1 U13290 ( .A(n14847), .ZN(n10876) );
  INV_X1 U13291 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n14985) );
  INV_X1 U13292 ( .A(n14809), .ZN(n10866) );
  INV_X1 U13293 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n14982) );
  INV_X1 U13294 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n14979) );
  OAI21_X1 U13295 ( .B1(n10839), .B2(n15112), .A(n10838), .ZN(n10840) );
  NAND2_X1 U13296 ( .A1(n10854), .A2(n10840), .ZN(n10841) );
  XNOR2_X1 U13297 ( .A(n14765), .B(n10840), .ZN(n14754) );
  NAND2_X1 U13298 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n14754), .ZN(n14753) );
  NAND2_X1 U13299 ( .A1(n10841), .A2(n14753), .ZN(n14780) );
  MUX2_X1 U13300 ( .A(n14979), .B(P3_REG1_REG_4__SCAN_IN), .S(n10895), .Z(
        n14779) );
  NAND2_X1 U13301 ( .A1(n14780), .A2(n14779), .ZN(n14778) );
  NAND2_X1 U13302 ( .A1(n14793), .A2(n10842), .ZN(n10843) );
  MUX2_X1 U13303 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n14982), .S(n14809), .Z(
        n14813) );
  NAND2_X1 U13304 ( .A1(n14814), .A2(n14813), .ZN(n14812) );
  OAI21_X1 U13305 ( .B1(n10866), .B2(n14982), .A(n14812), .ZN(n10844) );
  NAND2_X1 U13306 ( .A1(n10900), .A2(n10844), .ZN(n10845) );
  XNOR2_X1 U13307 ( .A(n10844), .B(n14829), .ZN(n14827) );
  NAND2_X1 U13308 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n14827), .ZN(n14826) );
  MUX2_X1 U13309 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n14985), .S(n14847), .Z(
        n14851) );
  NAND2_X1 U13310 ( .A1(n14867), .A2(n10846), .ZN(n10847) );
  NAND2_X1 U13311 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14873), .ZN(n14872) );
  AOI21_X1 U13312 ( .B1(n10849), .B2(n10848), .A(n11097), .ZN(n10916) );
  INV_X1 U13313 ( .A(n10850), .ZN(n14759) );
  INV_X1 U13314 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10851) );
  MUX2_X1 U13315 ( .A(n10852), .B(n10851), .S(n14738), .Z(n10853) );
  NAND2_X1 U13316 ( .A1(n10853), .A2(n14765), .ZN(n14771) );
  INV_X1 U13317 ( .A(n10853), .ZN(n10855) );
  NAND2_X1 U13318 ( .A1(n10855), .A2(n10854), .ZN(n10856) );
  AND2_X1 U13319 ( .A1(n14771), .A2(n10856), .ZN(n14758) );
  OAI21_X1 U13320 ( .B1(n14760), .B2(n14759), .A(n14758), .ZN(n14772) );
  MUX2_X1 U13321 ( .A(n10896), .B(n14979), .S(n14738), .Z(n10857) );
  NAND2_X1 U13322 ( .A1(n10857), .A2(n10895), .ZN(n10860) );
  INV_X1 U13323 ( .A(n10857), .ZN(n10858) );
  NAND2_X1 U13324 ( .A1(n10858), .A2(n14775), .ZN(n10859) );
  NAND2_X1 U13325 ( .A1(n10860), .A2(n10859), .ZN(n14770) );
  INV_X1 U13326 ( .A(n10860), .ZN(n14788) );
  INV_X1 U13327 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n10861) );
  MUX2_X1 U13328 ( .A(n10862), .B(n10861), .S(n14738), .Z(n10863) );
  NAND2_X1 U13329 ( .A1(n10863), .A2(n10898), .ZN(n14805) );
  INV_X1 U13330 ( .A(n10863), .ZN(n10864) );
  NAND2_X1 U13331 ( .A1(n10864), .A2(n14793), .ZN(n10865) );
  AND2_X1 U13332 ( .A1(n14805), .A2(n10865), .ZN(n14787) );
  OAI21_X1 U13333 ( .B1(n14789), .B2(n14788), .A(n14787), .ZN(n14806) );
  MUX2_X1 U13334 ( .A(n10957), .B(n14982), .S(n14738), .Z(n10867) );
  NAND2_X1 U13335 ( .A1(n10867), .A2(n10866), .ZN(n10870) );
  INV_X1 U13336 ( .A(n10867), .ZN(n10868) );
  NAND2_X1 U13337 ( .A1(n10868), .A2(n14809), .ZN(n10869) );
  NAND2_X1 U13338 ( .A1(n10870), .A2(n10869), .ZN(n14804) );
  AOI21_X1 U13339 ( .B1(n14806), .B2(n14805), .A(n14804), .ZN(n14823) );
  INV_X1 U13340 ( .A(n10870), .ZN(n14822) );
  INV_X1 U13341 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n10871) );
  MUX2_X1 U13342 ( .A(n10872), .B(n10871), .S(n14738), .Z(n10873) );
  NAND2_X1 U13343 ( .A1(n10873), .A2(n14829), .ZN(n14843) );
  INV_X1 U13344 ( .A(n10873), .ZN(n10874) );
  NAND2_X1 U13345 ( .A1(n10874), .A2(n10900), .ZN(n10875) );
  AND2_X1 U13346 ( .A1(n14843), .A2(n10875), .ZN(n14821) );
  OAI21_X1 U13347 ( .B1(n14823), .B2(n14822), .A(n14821), .ZN(n14844) );
  INV_X1 U13348 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10903) );
  MUX2_X1 U13349 ( .A(n10903), .B(n14985), .S(n14738), .Z(n10877) );
  NAND2_X1 U13350 ( .A1(n10877), .A2(n10876), .ZN(n10880) );
  INV_X1 U13351 ( .A(n10877), .ZN(n10878) );
  NAND2_X1 U13352 ( .A1(n10878), .A2(n14847), .ZN(n10879) );
  NAND2_X1 U13353 ( .A1(n10880), .A2(n10879), .ZN(n14842) );
  INV_X1 U13354 ( .A(n10880), .ZN(n14861) );
  INV_X1 U13355 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n10881) );
  MUX2_X1 U13356 ( .A(n11272), .B(n10881), .S(n14738), .Z(n10882) );
  NAND2_X1 U13357 ( .A1(n10882), .A2(n10905), .ZN(n10889) );
  INV_X1 U13358 ( .A(n10882), .ZN(n10883) );
  NAND2_X1 U13359 ( .A1(n10883), .A2(n14867), .ZN(n10884) );
  AND2_X1 U13360 ( .A1(n10889), .A2(n10884), .ZN(n14860) );
  OAI21_X1 U13361 ( .B1(n14862), .B2(n14861), .A(n14860), .ZN(n14859) );
  MUX2_X1 U13362 ( .A(n10907), .B(n14988), .S(n14738), .Z(n10885) );
  NAND2_X1 U13363 ( .A1(n10885), .A2(n11098), .ZN(n11102) );
  INV_X1 U13364 ( .A(n10885), .ZN(n10886) );
  NAND2_X1 U13365 ( .A1(n10886), .A2(n11095), .ZN(n10887) );
  NAND2_X1 U13366 ( .A1(n11102), .A2(n10887), .ZN(n10888) );
  AOI21_X1 U13367 ( .B1(n14859), .B2(n10889), .A(n10888), .ZN(n11104) );
  AND3_X1 U13368 ( .A1(n14859), .A2(n10889), .A3(n10888), .ZN(n10890) );
  OAI21_X1 U13369 ( .B1(n11104), .B2(n10890), .A(n14863), .ZN(n10915) );
  MUX2_X1 U13370 ( .A(P3_REG2_REG_4__SCAN_IN), .B(n10896), .S(n10895), .Z(
        n14769) );
  NOR2_X1 U13371 ( .A1(n10898), .A2(n10897), .ZN(n10899) );
  XNOR2_X1 U13372 ( .A(n10898), .B(n10897), .ZN(n14786) );
  MUX2_X1 U13373 ( .A(n10957), .B(P3_REG2_REG_6__SCAN_IN), .S(n14809), .Z(
        n14803) );
  NOR2_X1 U13374 ( .A1(n14829), .A2(n10901), .ZN(n10902) );
  NOR2_X1 U13375 ( .A1(n10872), .A2(n14820), .ZN(n14819) );
  MUX2_X1 U13376 ( .A(n10903), .B(P3_REG2_REG_8__SCAN_IN), .S(n14847), .Z(
        n14840) );
  NOR2_X1 U13377 ( .A1(n10905), .A2(n10904), .ZN(n10906) );
  MUX2_X1 U13378 ( .A(P3_REG2_REG_10__SCAN_IN), .B(n10907), .S(n11098), .Z(
        n10908) );
  AOI21_X1 U13379 ( .B1(n6580), .B2(n10908), .A(n11094), .ZN(n10909) );
  NOR2_X1 U13380 ( .A1(n14878), .A2(n10909), .ZN(n10913) );
  INV_X1 U13381 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n10911) );
  INV_X1 U13382 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15038) );
  NOR2_X1 U13383 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15038), .ZN(n11367) );
  INV_X1 U13384 ( .A(n11367), .ZN(n10910) );
  OAI21_X1 U13385 ( .B1(n14837), .B2(n10911), .A(n10910), .ZN(n10912) );
  AOI211_X1 U13386 ( .C1(n14828), .C2(n11098), .A(n10913), .B(n10912), .ZN(
        n10914) );
  OAI211_X1 U13387 ( .C1(n10916), .C2(n14741), .A(n10915), .B(n10914), .ZN(
        P3_U3192) );
  XNOR2_X1 U13388 ( .A(n10917), .B(n10918), .ZN(n14959) );
  NAND2_X1 U13389 ( .A1(n14959), .A2(n14906), .ZN(n10924) );
  XNOR2_X1 U13390 ( .A(n14882), .B(n10918), .ZN(n10922) );
  NAND2_X1 U13391 ( .A1(n11992), .A2(n14920), .ZN(n10919) );
  OAI21_X1 U13392 ( .B1(n10920), .B2(n14903), .A(n10919), .ZN(n10921) );
  AOI21_X1 U13393 ( .B1(n10922), .B2(n14923), .A(n10921), .ZN(n10923) );
  NAND2_X1 U13394 ( .A1(n10924), .A2(n10923), .ZN(n14964) );
  AOI21_X1 U13395 ( .B1(n14929), .B2(n10977), .A(n14964), .ZN(n10928) );
  OAI22_X1 U13396 ( .A1(n12391), .A2(n10925), .B1(n10872), .B2(n14933), .ZN(
        n10926) );
  AOI21_X1 U13397 ( .B1(n14959), .B2(n14930), .A(n10926), .ZN(n10927) );
  OAI21_X1 U13398 ( .B1(n10928), .B2(n14935), .A(n10927), .ZN(P3_U3226) );
  INV_X1 U13399 ( .A(n10933), .ZN(n14705) );
  NAND2_X1 U13400 ( .A1(n12735), .A2(n10022), .ZN(n11081) );
  XNOR2_X1 U13401 ( .A(n10933), .B(n6816), .ZN(n11079) );
  XOR2_X1 U13402 ( .A(n11081), .B(n11079), .Z(n10935) );
  AOI21_X1 U13403 ( .B1(n10934), .B2(n10935), .A(n12724), .ZN(n10936) );
  NAND2_X1 U13404 ( .A1(n10936), .A2(n11080), .ZN(n10941) );
  AND2_X1 U13405 ( .A1(P2_U3088), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n12839) );
  NOR2_X1 U13406 ( .A1(n12720), .A2(n10937), .ZN(n10938) );
  AOI211_X1 U13407 ( .C1(n12717), .C2(n10939), .A(n12839), .B(n10938), .ZN(
        n10940) );
  OAI211_X1 U13408 ( .C1(n14705), .C2(n12653), .A(n10941), .B(n10940), .ZN(
        P2_U3189) );
  INV_X1 U13409 ( .A(n11579), .ZN(n11008) );
  OAI222_X1 U13410 ( .A1(n13201), .A2(n10943), .B1(n13199), .B2(n11008), .C1(
        n10942), .C2(P2_U3088), .ZN(P2_U3307) );
  OAI21_X1 U13411 ( .B1(n10946), .B2(n10945), .A(n10944), .ZN(n14958) );
  INV_X1 U13412 ( .A(n14958), .ZN(n10962) );
  OAI22_X1 U13413 ( .A1(n10948), .A2(n14903), .B1(n10947), .B2(n14901), .ZN(
        n10956) );
  INV_X1 U13414 ( .A(n10949), .ZN(n10954) );
  AOI21_X1 U13415 ( .B1(n10952), .B2(n10951), .A(n10950), .ZN(n10953) );
  NOR3_X1 U13416 ( .A1(n10954), .A2(n10953), .A3(n14891), .ZN(n10955) );
  AOI211_X1 U13417 ( .C1(n14906), .C2(n14958), .A(n10956), .B(n10955), .ZN(
        n14955) );
  MUX2_X1 U13418 ( .A(n10957), .B(n14955), .S(n14933), .Z(n10961) );
  AND2_X1 U13419 ( .A1(n10958), .A2(n14960), .ZN(n14957) );
  AOI22_X1 U13420 ( .A1(n14896), .A2(n14957), .B1(n14929), .B2(n10959), .ZN(
        n10960) );
  OAI211_X1 U13421 ( .C1(n10962), .C2(n11244), .A(n10961), .B(n10960), .ZN(
        P3_U3227) );
  XNOR2_X1 U13422 ( .A(n10963), .B(n10964), .ZN(n14184) );
  XOR2_X1 U13423 ( .A(n10965), .B(n10964), .Z(n10967) );
  OAI22_X1 U13424 ( .A1(n11288), .A2(n13055), .B1(n11418), .B2(n13057), .ZN(
        n10966) );
  AOI21_X1 U13425 ( .B1(n10967), .B2(n13065), .A(n10966), .ZN(n10968) );
  OAI21_X1 U13426 ( .B1(n14184), .B2(n14689), .A(n10968), .ZN(n14187) );
  NAND2_X1 U13427 ( .A1(n14187), .A2(n13038), .ZN(n10976) );
  OAI22_X1 U13428 ( .A1(n13038), .A2(n10969), .B1(n11287), .B2(n12998), .ZN(
        n10973) );
  INV_X1 U13429 ( .A(n10970), .ZN(n11119) );
  OAI211_X1 U13430 ( .C1(n14186), .C2(n10971), .A(n11119), .B(n6438), .ZN(
        n14185) );
  NOR2_X1 U13431 ( .A1(n14185), .A2(n12984), .ZN(n10972) );
  AOI211_X1 U13432 ( .C1(n13082), .C2(n10974), .A(n10973), .B(n10972), .ZN(
        n10975) );
  OAI211_X1 U13433 ( .C1(n14184), .C2(n13083), .A(n10976), .B(n10975), .ZN(
        P2_U3253) );
  INV_X1 U13434 ( .A(n10977), .ZN(n10985) );
  OAI211_X1 U13435 ( .C1(n10980), .C2(n10979), .A(n10978), .B(n11963), .ZN(
        n10984) );
  NAND2_X1 U13436 ( .A1(n11974), .A2(n11993), .ZN(n10981) );
  NAND2_X1 U13437 ( .A1(P3_REG3_REG_7__SCAN_IN), .A2(P3_U3151), .ZN(n14835) );
  OAI211_X1 U13438 ( .C1(n11977), .C2(n11155), .A(n10981), .B(n14835), .ZN(
        n10982) );
  AOI21_X1 U13439 ( .B1(n11979), .B2(n14961), .A(n10982), .ZN(n10983) );
  OAI211_X1 U13440 ( .C1(n10985), .C2(n11373), .A(n10984), .B(n10983), .ZN(
        P3_U3153) );
  NAND2_X1 U13441 ( .A1(n11726), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10992) );
  OR2_X1 U13442 ( .A1(n11731), .A2(n10155), .ZN(n10991) );
  NAND2_X1 U13443 ( .A1(n10986), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n11029) );
  OR2_X1 U13444 ( .A1(n10986), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10987) );
  NAND2_X1 U13445 ( .A1(n11029), .A2(n10987), .ZN(n13390) );
  OR2_X1 U13446 ( .A1(n11634), .A2(n13390), .ZN(n10990) );
  OR2_X1 U13447 ( .A1(n6743), .A2(n10988), .ZN(n10989) );
  NAND4_X1 U13448 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n13475) );
  NAND2_X1 U13449 ( .A1(n10995), .A2(n11743), .ZN(n10997) );
  AOI22_X1 U13450 ( .A1(n6451), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n13572), 
        .B2(n11556), .ZN(n10996) );
  INV_X1 U13451 ( .A(n13476), .ZN(n11344) );
  XNOR2_X1 U13452 ( .A(n14226), .B(n11344), .ZN(n11767) );
  XNOR2_X1 U13453 ( .A(n11037), .B(n11767), .ZN(n10998) );
  AOI222_X1 U13454 ( .A1(n13477), .A2(n13865), .B1(n13475), .B2(n13835), .C1(
        n14429), .C2(n10998), .ZN(n14300) );
  OR2_X1 U13455 ( .A1(n14537), .A2(n13477), .ZN(n11000) );
  XNOR2_X1 U13456 ( .A(n11017), .B(n11767), .ZN(n14303) );
  INV_X1 U13457 ( .A(n14226), .ZN(n14299) );
  NAND2_X1 U13458 ( .A1(n14299), .A2(n11001), .ZN(n14122) );
  OAI211_X1 U13459 ( .C1(n14299), .C2(n11001), .A(n14412), .B(n14122), .ZN(
        n14298) );
  OAI22_X1 U13460 ( .A1(n14420), .A2(n11002), .B1(n14229), .B2(n14416), .ZN(
        n11003) );
  AOI21_X1 U13461 ( .B1(n14226), .B2(n14430), .A(n11003), .ZN(n11004) );
  OAI21_X1 U13462 ( .B1(n14298), .B2(n13875), .A(n11004), .ZN(n11005) );
  AOI21_X1 U13463 ( .B1(n14303), .B2(n14252), .A(n11005), .ZN(n11006) );
  OAI21_X1 U13464 ( .B1(n14300), .B2(n14439), .A(n11006), .ZN(P1_U3282) );
  OAI222_X1 U13465 ( .A1(n13986), .A2(n11008), .B1(P1_U3086), .B2(n11434), 
        .C1(n11007), .C2(n13988), .ZN(P1_U3335) );
  INV_X1 U13466 ( .A(n11597), .ZN(n11011) );
  OAI222_X1 U13467 ( .A1(n13988), .A2(n11009), .B1(n13986), .B2(n11011), .C1(
        n11433), .C2(P1_U3086), .ZN(P1_U3334) );
  OAI222_X1 U13468 ( .A1(n13201), .A2(n11012), .B1(n13199), .B2(n11011), .C1(
        P2_U3088), .C2(n11010), .ZN(P2_U3306) );
  INV_X1 U13469 ( .A(n11013), .ZN(n11014) );
  OAI222_X1 U13470 ( .A1(n11016), .A2(P3_U3151), .B1(n12530), .B2(n11015), 
        .C1(n12528), .C2(n11014), .ZN(P3_U3270) );
  NAND2_X1 U13471 ( .A1(n11018), .A2(n11743), .ZN(n11021) );
  AOI22_X1 U13472 ( .A1(n11019), .A2(n11556), .B1(n6451), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n11020) );
  XNOR2_X1 U13473 ( .A(n14120), .B(n13475), .ZN(n14114) );
  NAND2_X1 U13474 ( .A1(n14113), .A2(n6957), .ZN(n11023) );
  OR2_X1 U13475 ( .A1(n14120), .A2(n13475), .ZN(n11022) );
  NAND2_X1 U13476 ( .A1(n11023), .A2(n11022), .ZN(n11194) );
  NAND2_X1 U13477 ( .A1(n11024), .A2(n11743), .ZN(n11027) );
  AOI22_X1 U13478 ( .A1(n11025), .A2(n11556), .B1(n11744), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n11026) );
  NAND2_X1 U13479 ( .A1(n11726), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n11035) );
  OR2_X1 U13480 ( .A1(n11731), .A2(n10185), .ZN(n11034) );
  INV_X1 U13481 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11028) );
  NAND2_X1 U13482 ( .A1(n11029), .A2(n11028), .ZN(n11030) );
  NAND2_X1 U13483 ( .A1(n11041), .A2(n11030), .ZN(n11049) );
  OR2_X1 U13484 ( .A1(n11634), .A2(n11049), .ZN(n11033) );
  OR2_X1 U13485 ( .A1(n6743), .A2(n11031), .ZN(n11032) );
  NAND4_X1 U13486 ( .A1(n11035), .A2(n11034), .A3(n11033), .A4(n11032), .ZN(
        n13474) );
  XNOR2_X1 U13487 ( .A(n13433), .B(n13474), .ZN(n11769) );
  XNOR2_X1 U13488 ( .A(n11194), .B(n11769), .ZN(n14294) );
  INV_X1 U13489 ( .A(n11767), .ZN(n11036) );
  INV_X1 U13490 ( .A(n13475), .ZN(n14216) );
  OR2_X1 U13491 ( .A1(n14120), .A2(n14216), .ZN(n11038) );
  XNOR2_X1 U13492 ( .A(n11175), .B(n6982), .ZN(n14297) );
  NAND2_X1 U13493 ( .A1(n14297), .A2(n13842), .ZN(n11056) );
  INV_X1 U13494 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11040) );
  AND2_X1 U13495 ( .A1(n11041), .A2(n11040), .ZN(n11042) );
  OR2_X1 U13496 ( .A1(n11042), .A2(n11223), .ZN(n14205) );
  INV_X1 U13497 ( .A(n14205), .ZN(n11189) );
  NAND2_X1 U13498 ( .A1(n11621), .A2(n11189), .ZN(n11048) );
  OR2_X1 U13499 ( .A1(n11731), .A2(n11128), .ZN(n11047) );
  OR2_X1 U13500 ( .A1(n6743), .A2(n14291), .ZN(n11046) );
  INV_X1 U13501 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11043) );
  OR2_X1 U13502 ( .A1(n11044), .A2(n11043), .ZN(n11045) );
  INV_X1 U13503 ( .A(n13236), .ZN(n13473) );
  AOI22_X1 U13504 ( .A1(n13473), .A2(n13835), .B1(n13865), .B2(n13475), .ZN(
        n14292) );
  INV_X1 U13505 ( .A(n14292), .ZN(n11050) );
  INV_X1 U13506 ( .A(n11049), .ZN(n13438) );
  INV_X1 U13507 ( .A(n14416), .ZN(n14431) );
  AOI22_X1 U13508 ( .A1(n11050), .A2(n14420), .B1(n13438), .B2(n14431), .ZN(
        n11051) );
  OAI21_X1 U13509 ( .B1(n10185), .B2(n14420), .A(n11051), .ZN(n11054) );
  AOI21_X1 U13510 ( .B1(n13433), .B2(n14123), .A(n14468), .ZN(n11052) );
  NAND2_X1 U13511 ( .A1(n11052), .A2(n11187), .ZN(n14293) );
  NOR2_X1 U13512 ( .A1(n14293), .A2(n13875), .ZN(n11053) );
  AOI211_X1 U13513 ( .C1(n14430), .C2(n13433), .A(n11054), .B(n11053), .ZN(
        n11055) );
  OAI211_X1 U13514 ( .C1(n14294), .C2(n13844), .A(n11056), .B(n11055), .ZN(
        P1_U3280) );
  INV_X1 U13515 ( .A(n14238), .ZN(n13469) );
  INV_X1 U13516 ( .A(n11057), .ZN(n11060) );
  INV_X1 U13517 ( .A(n11058), .ZN(n11059) );
  NAND2_X1 U13518 ( .A1(n14515), .A2(n7444), .ZN(n11064) );
  NAND2_X1 U13519 ( .A1(n13479), .A2(n6443), .ZN(n11063) );
  NAND2_X1 U13520 ( .A1(n11064), .A2(n11063), .ZN(n11065) );
  XNOR2_X1 U13521 ( .A(n11065), .B(n13365), .ZN(n11069) );
  NAND2_X1 U13522 ( .A1(n14515), .A2(n6443), .ZN(n11067) );
  NAND2_X1 U13523 ( .A1(n13331), .A2(n13479), .ZN(n11066) );
  NAND2_X1 U13524 ( .A1(n11067), .A2(n11066), .ZN(n11068) );
  OAI21_X1 U13525 ( .B1(n6582), .B2(n6455), .A(n11261), .ZN(n11070) );
  NAND2_X1 U13526 ( .A1(n11070), .A2(n14233), .ZN(n11077) );
  INV_X1 U13527 ( .A(n11071), .ZN(n11074) );
  NOR2_X1 U13528 ( .A1(n14241), .A2(n11072), .ZN(n11073) );
  AOI211_X1 U13529 ( .C1(n14235), .C2(n11075), .A(n11074), .B(n11073), .ZN(
        n11076) );
  OAI211_X1 U13530 ( .C1(n11078), .C2(n13469), .A(n11077), .B(n11076), .ZN(
        P1_U3221) );
  XNOR2_X1 U13531 ( .A(n14716), .B(n6816), .ZN(n11083) );
  OR2_X1 U13532 ( .A1(n11288), .A2(n6438), .ZN(n11082) );
  NOR2_X1 U13533 ( .A1(n11083), .A2(n11082), .ZN(n11281) );
  NAND2_X1 U13534 ( .A1(n11083), .A2(n11082), .ZN(n11282) );
  INV_X1 U13535 ( .A(n11282), .ZN(n11084) );
  NOR2_X1 U13536 ( .A1(n11281), .A2(n11084), .ZN(n11085) );
  XNOR2_X1 U13537 ( .A(n11283), .B(n11085), .ZN(n11093) );
  NAND2_X1 U13538 ( .A1(n12717), .A2(n11086), .ZN(n11087) );
  OAI211_X1 U13539 ( .C1(n12720), .C2(n11089), .A(n11088), .B(n11087), .ZN(
        n11090) );
  AOI21_X1 U13540 ( .B1(n11091), .B2(n12722), .A(n11090), .ZN(n11092) );
  OAI21_X1 U13541 ( .B1(n11093), .B2(n12724), .A(n11092), .ZN(P2_U3208) );
  XNOR2_X1 U13542 ( .A(n12007), .B(n12006), .ZN(n11096) );
  AOI21_X1 U13543 ( .B1(n11384), .B2(n11096), .A(n12008), .ZN(n11112) );
  OAI21_X1 U13544 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11099), .A(n12019), 
        .ZN(n11110) );
  INV_X1 U13545 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n11100) );
  NOR2_X1 U13546 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11100), .ZN(n11939) );
  AOI21_X1 U13547 ( .B1(n14871), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11939), 
        .ZN(n11101) );
  OAI21_X1 U13548 ( .B1(n14868), .B2(n12018), .A(n11101), .ZN(n11109) );
  INV_X1 U13549 ( .A(n11102), .ZN(n11103) );
  NOR2_X1 U13550 ( .A1(n11104), .A2(n11103), .ZN(n11106) );
  MUX2_X1 U13551 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n14738), .Z(n11998) );
  XNOR2_X1 U13552 ( .A(n11998), .B(n12018), .ZN(n11105) );
  AOI21_X1 U13553 ( .B1(n11106), .B2(n11105), .A(n12001), .ZN(n11107) );
  NOR2_X1 U13554 ( .A1(n11107), .A2(n14761), .ZN(n11108) );
  AOI211_X1 U13555 ( .C1(n14874), .C2(n11110), .A(n11109), .B(n11108), .ZN(
        n11111) );
  OAI21_X1 U13556 ( .B1(n11112), .B2(n14878), .A(n11111), .ZN(P3_U3193) );
  XNOR2_X1 U13557 ( .A(n11114), .B(n11113), .ZN(n11326) );
  XNOR2_X1 U13558 ( .A(n11116), .B(n11115), .ZN(n11117) );
  OAI222_X1 U13559 ( .A1(n13057), .A2(n11315), .B1(n13055), .B2(n11317), .C1(
        n11117), .C2(n13029), .ZN(n11322) );
  NAND2_X1 U13560 ( .A1(n11322), .A2(n13038), .ZN(n11124) );
  INV_X1 U13561 ( .A(n11211), .ZN(n11118) );
  AOI211_X1 U13562 ( .C1(n11324), .C2(n11119), .A(n10022), .B(n11118), .ZN(
        n11323) );
  NOR2_X1 U13563 ( .A1(n11314), .A2(n13073), .ZN(n11122) );
  OAI22_X1 U13564 ( .A1(n13038), .A2(n11120), .B1(n11316), .B2(n12998), .ZN(
        n11121) );
  AOI211_X1 U13565 ( .C1(n11323), .C2(n13085), .A(n11122), .B(n11121), .ZN(
        n11123) );
  OAI211_X1 U13566 ( .C1(n11326), .C2(n13053), .A(n11124), .B(n11123), .ZN(
        P2_U3252) );
  NAND2_X1 U13567 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n13585), .ZN(n11131) );
  INV_X1 U13568 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11126) );
  INV_X1 U13569 ( .A(n11131), .ZN(n11125) );
  AOI21_X1 U13570 ( .B1(n11126), .B2(n11142), .A(n11125), .ZN(n13587) );
  OAI21_X1 U13571 ( .B1(n11128), .B2(n11137), .A(n11127), .ZN(n11129) );
  NOR2_X1 U13572 ( .A1(n14356), .A2(n11129), .ZN(n11130) );
  XNOR2_X1 U13573 ( .A(n11129), .B(n14356), .ZN(n14351) );
  NOR2_X1 U13574 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14351), .ZN(n14350) );
  NOR2_X1 U13575 ( .A1(n11130), .A2(n14350), .ZN(n13588) );
  NAND2_X1 U13576 ( .A1(n13587), .A2(n13588), .ZN(n13586) );
  NAND2_X1 U13577 ( .A1(n11131), .A2(n13586), .ZN(n11134) );
  INV_X1 U13578 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n11132) );
  AOI22_X1 U13579 ( .A1(n13598), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n11132), 
        .B2(n13593), .ZN(n11133) );
  NAND2_X1 U13580 ( .A1(n11133), .A2(n11134), .ZN(n13599) );
  OAI211_X1 U13581 ( .C1(n11134), .C2(n11133), .A(n14370), .B(n13599), .ZN(
        n11148) );
  NAND2_X1 U13582 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13410)
         );
  INV_X1 U13583 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n15023) );
  NOR2_X1 U13584 ( .A1(n13593), .A2(n15023), .ZN(n11135) );
  AOI21_X1 U13585 ( .B1(n15023), .B2(n13593), .A(n11135), .ZN(n11144) );
  INV_X1 U13586 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14276) );
  AOI21_X1 U13587 ( .B1(n11137), .B2(n14291), .A(n11136), .ZN(n11139) );
  NOR2_X1 U13588 ( .A1(n14356), .A2(n11139), .ZN(n11140) );
  XOR2_X1 U13589 ( .A(n11139), .B(n11138), .Z(n14353) );
  NOR2_X1 U13590 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n14353), .ZN(n14352) );
  NOR2_X1 U13591 ( .A1(n11140), .A2(n14352), .ZN(n13583) );
  NOR2_X1 U13592 ( .A1(n11142), .A2(n14276), .ZN(n11141) );
  AOI21_X1 U13593 ( .B1(n14276), .B2(n11142), .A(n11141), .ZN(n13582) );
  NAND2_X1 U13594 ( .A1(n13583), .A2(n13582), .ZN(n13581) );
  OAI21_X1 U13595 ( .B1(n14276), .B2(n11142), .A(n13581), .ZN(n11143) );
  NAND2_X1 U13596 ( .A1(n11143), .A2(n11144), .ZN(n13592) );
  OAI211_X1 U13597 ( .C1(n11144), .C2(n11143), .A(n14367), .B(n13592), .ZN(
        n11145) );
  NAND2_X1 U13598 ( .A1(n13410), .A2(n11145), .ZN(n11146) );
  AOI21_X1 U13599 ( .B1(n14346), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n11146), 
        .ZN(n11147) );
  OAI211_X1 U13600 ( .C1(n14375), .C2(n13593), .A(n11148), .B(n11147), .ZN(
        P1_U3260) );
  INV_X1 U13601 ( .A(n11149), .ZN(n11150) );
  OAI222_X1 U13602 ( .A1(n13201), .A2(n11151), .B1(n13199), .B2(n11150), .C1(
        n8194), .C2(P2_U3088), .ZN(P2_U3305) );
  XNOR2_X1 U13603 ( .A(n11152), .B(n7404), .ZN(n11278) );
  INV_X1 U13604 ( .A(n14972), .ZN(n12421) );
  AOI21_X1 U13605 ( .B1(n11154), .B2(n11153), .A(n14891), .ZN(n11158) );
  OAI22_X1 U13606 ( .A1(n11155), .A2(n14903), .B1(n11303), .B2(n14901), .ZN(
        n11156) );
  AOI21_X1 U13607 ( .B1(n11158), .B2(n11157), .A(n11156), .ZN(n11273) );
  OAI21_X1 U13608 ( .B1(n11278), .B2(n12421), .A(n11273), .ZN(n11163) );
  OAI22_X1 U13609 ( .A1(n12459), .A2(n11306), .B1(n14990), .B2(n10881), .ZN(
        n11159) );
  AOI21_X1 U13610 ( .B1(n11163), .B2(n14990), .A(n11159), .ZN(n11160) );
  INV_X1 U13611 ( .A(n11160), .ZN(P3_U3468) );
  INV_X1 U13612 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n11161) );
  OAI22_X1 U13613 ( .A1(n11306), .A2(n12510), .B1(n14974), .B2(n11161), .ZN(
        n11162) );
  AOI21_X1 U13614 ( .B1(n11163), .B2(n14974), .A(n11162), .ZN(n11164) );
  INV_X1 U13615 ( .A(n11164), .ZN(P3_U3417) );
  INV_X1 U13616 ( .A(n14895), .ZN(n11174) );
  OAI211_X1 U13617 ( .C1(n11167), .C2(n11166), .A(n11165), .B(n11963), .ZN(
        n11173) );
  AND2_X1 U13618 ( .A1(P3_U3151), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n14849) );
  AOI21_X1 U13619 ( .B1(n11940), .B2(n14888), .A(n14849), .ZN(n11168) );
  OAI21_X1 U13620 ( .B1(n11169), .B2(n11977), .A(n11168), .ZN(n11170) );
  AOI21_X1 U13621 ( .B1(n11979), .B2(n11171), .A(n11170), .ZN(n11172) );
  OAI211_X1 U13622 ( .C1(n11174), .C2(n11373), .A(n11173), .B(n11172), .ZN(
        P3_U3161) );
  INV_X1 U13623 ( .A(n13474), .ZN(n14194) );
  NAND2_X1 U13624 ( .A1(n11176), .A2(n11743), .ZN(n11179) );
  AOI22_X1 U13625 ( .A1(n11177), .A2(n11556), .B1(n6451), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11178) );
  NAND2_X1 U13626 ( .A1(n14285), .A2(n13236), .ZN(n11502) );
  NAND2_X1 U13627 ( .A1(n11508), .A2(n11502), .ZN(n11771) );
  INV_X1 U13628 ( .A(n11771), .ZN(n11507) );
  XNOR2_X1 U13629 ( .A(n6574), .B(n11507), .ZN(n11186) );
  XNOR2_X1 U13630 ( .A(n11223), .B(P1_REG3_REG_15__SCAN_IN), .ZN(n14240) );
  OR2_X1 U13631 ( .A1(n14240), .A2(n11634), .ZN(n11183) );
  NAND2_X1 U13632 ( .A1(n15191), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n11182) );
  NAND2_X1 U13633 ( .A1(n11711), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n11181) );
  NAND2_X1 U13634 ( .A1(n11726), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n11180) );
  NAND2_X1 U13635 ( .A1(n13474), .A2(n13865), .ZN(n11184) );
  OAI21_X1 U13636 ( .B1(n14208), .B2(n14380), .A(n11184), .ZN(n11185) );
  AOI21_X1 U13637 ( .B1(n11186), .B2(n14429), .A(n11185), .ZN(n14290) );
  INV_X1 U13638 ( .A(n13857), .ZN(n11192) );
  NAND2_X1 U13639 ( .A1(n14285), .A2(n11187), .ZN(n11188) );
  AND2_X1 U13640 ( .A1(n11233), .A2(n11188), .ZN(n14286) );
  AOI22_X1 U13641 ( .A1(n14439), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n11189), 
        .B2(n14431), .ZN(n11190) );
  OAI21_X1 U13642 ( .B1(n6932), .B2(n13876), .A(n11190), .ZN(n11191) );
  AOI21_X1 U13643 ( .B1(n11192), .B2(n14286), .A(n11191), .ZN(n11197) );
  NOR2_X1 U13644 ( .A1(n13433), .A2(n13474), .ZN(n11193) );
  AOI21_X1 U13645 ( .B1(n11194), .B2(n6982), .A(n11193), .ZN(n11195) );
  OR2_X1 U13646 ( .A1(n11195), .A2(n11771), .ZN(n14283) );
  NAND3_X1 U13647 ( .A1(n14283), .A2(n14284), .A3(n14252), .ZN(n11196) );
  OAI211_X1 U13648 ( .C1(n14290), .C2(n14439), .A(n11197), .B(n11196), .ZN(
        P1_U3279) );
  INV_X1 U13649 ( .A(n11198), .ZN(n11199) );
  OAI222_X1 U13650 ( .A1(n11201), .A2(P3_U3151), .B1(n12530), .B2(n11200), 
        .C1(n12528), .C2(n11199), .ZN(P3_U3269) );
  INV_X1 U13651 ( .A(n11627), .ZN(n11206) );
  AOI21_X1 U13652 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n13196), .A(n11202), 
        .ZN(n11203) );
  OAI21_X1 U13653 ( .B1(n11206), .B2(n13199), .A(n11203), .ZN(P2_U3304) );
  INV_X1 U13654 ( .A(n13988), .ZN(n13976) );
  AOI21_X1 U13655 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n13976), .A(n11204), 
        .ZN(n11205) );
  OAI21_X1 U13656 ( .B1(n11206), .B2(n13986), .A(n11205), .ZN(P1_U3332) );
  XNOR2_X1 U13657 ( .A(n11207), .B(n11210), .ZN(n11208) );
  OAI222_X1 U13658 ( .A1(n13055), .A2(n11418), .B1(n13057), .B2(n13056), .C1(
        n11208), .C2(n13029), .ZN(n14181) );
  INV_X1 U13659 ( .A(n14181), .ZN(n11218) );
  XOR2_X1 U13660 ( .A(n11210), .B(n11209), .Z(n14183) );
  AOI21_X1 U13661 ( .B1(n11406), .B2(n11211), .A(n10022), .ZN(n11212) );
  NAND2_X1 U13662 ( .A1(n11212), .A2(n11390), .ZN(n14179) );
  INV_X1 U13663 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11213) );
  OAI22_X1 U13664 ( .A1(n13038), .A2(n11213), .B1(n11417), .B2(n12998), .ZN(
        n11214) );
  AOI21_X1 U13665 ( .B1(n11406), .B2(n13082), .A(n11214), .ZN(n11215) );
  OAI21_X1 U13666 ( .B1(n14179), .B2(n12984), .A(n11215), .ZN(n11216) );
  AOI21_X1 U13667 ( .B1(n14183), .B2(n12988), .A(n11216), .ZN(n11217) );
  OAI21_X1 U13668 ( .B1(n11218), .B2(n13078), .A(n11217), .ZN(P2_U3251) );
  NAND2_X1 U13669 ( .A1(n11219), .A2(n11743), .ZN(n11221) );
  AOI22_X1 U13670 ( .A1(n11744), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11556), 
        .B2(n14356), .ZN(n11220) );
  NAND2_X1 U13671 ( .A1(n14237), .A2(n14208), .ZN(n11510) );
  AOI21_X1 U13672 ( .B1(n6566), .B2(n7206), .A(n14540), .ZN(n11230) );
  OR2_X1 U13673 ( .A1(n13236), .A2(n14382), .ZN(n11229) );
  AND2_X1 U13674 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_16__SCAN_IN), 
        .ZN(n11222) );
  AOI21_X1 U13675 ( .B1(n11223), .B2(P1_REG3_REG_15__SCAN_IN), .A(
        P1_REG3_REG_16__SCAN_IN), .ZN(n11224) );
  OR2_X1 U13676 ( .A1(n11514), .A2(n11224), .ZN(n14244) );
  OAI22_X1 U13677 ( .A1(n14244), .A2(n11634), .B1(n6743), .B2(n14276), .ZN(
        n11227) );
  NAND2_X1 U13678 ( .A1(n11726), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n11225) );
  OAI21_X1 U13679 ( .B1(n11126), .B2(n11731), .A(n11225), .ZN(n11226) );
  NAND2_X1 U13680 ( .A1(n13866), .A2(n13835), .ZN(n11228) );
  NAND2_X1 U13681 ( .A1(n11229), .A2(n11228), .ZN(n14236) );
  AOI21_X1 U13682 ( .B1(n11230), .B2(n13656), .A(n14236), .ZN(n14278) );
  NAND2_X1 U13683 ( .A1(n14285), .A2(n13473), .ZN(n11231) );
  NAND2_X1 U13684 ( .A1(n14284), .A2(n11231), .ZN(n11232) );
  OAI21_X1 U13685 ( .B1(n7207), .B2(n7206), .A(n13630), .ZN(n14281) );
  OAI211_X1 U13686 ( .C1(n6931), .C2(n6442), .A(n14412), .B(n14251), .ZN(
        n14277) );
  INV_X1 U13687 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11234) );
  OAI22_X1 U13688 ( .A1(n14420), .A2(n11234), .B1(n14240), .B2(n14416), .ZN(
        n11235) );
  AOI21_X1 U13689 ( .B1(n14237), .B2(n14430), .A(n11235), .ZN(n11236) );
  OAI21_X1 U13690 ( .B1(n14277), .B2(n13875), .A(n11236), .ZN(n11237) );
  AOI21_X1 U13691 ( .B1(n14281), .B2(n14252), .A(n11237), .ZN(n11238) );
  OAI21_X1 U13692 ( .B1(n14278), .B2(n14439), .A(n11238), .ZN(P1_U3278) );
  INV_X1 U13693 ( .A(n11640), .ZN(n11242) );
  OAI222_X1 U13694 ( .A1(n13201), .A2(n15122), .B1(n13199), .B2(n11242), .C1(
        n11239), .C2(P2_U3088), .ZN(P2_U3303) );
  INV_X1 U13695 ( .A(n11240), .ZN(n11241) );
  OAI222_X1 U13696 ( .A1(n13988), .A2(n15035), .B1(n13986), .B2(n11242), .C1(
        n11241), .C2(P1_U3086), .ZN(P1_U3331) );
  NAND2_X1 U13697 ( .A1(n14933), .A2(n14906), .ZN(n11243) );
  INV_X1 U13698 ( .A(n12393), .ZN(n12327) );
  XNOR2_X1 U13699 ( .A(n11245), .B(n11247), .ZN(n14971) );
  INV_X1 U13700 ( .A(n14971), .ZN(n11257) );
  OAI211_X1 U13701 ( .C1(n11248), .C2(n11247), .A(n11246), .B(n14923), .ZN(
        n11250) );
  AOI22_X1 U13702 ( .A1(n11866), .A2(n14920), .B1(n14919), .B2(n14887), .ZN(
        n11249) );
  NAND2_X1 U13703 ( .A1(n11250), .A2(n11249), .ZN(n14969) );
  NOR2_X1 U13704 ( .A1(n14933), .A2(n10907), .ZN(n11255) );
  AND2_X1 U13705 ( .A1(n11370), .A2(n14960), .ZN(n14970) );
  INV_X1 U13706 ( .A(n14970), .ZN(n11252) );
  INV_X1 U13707 ( .A(n11251), .ZN(n11374) );
  OAI22_X1 U13708 ( .A1(n11253), .A2(n11252), .B1(n11374), .B2(n12271), .ZN(
        n11254) );
  AOI211_X1 U13709 ( .C1(n14969), .C2(n14933), .A(n11255), .B(n11254), .ZN(
        n11256) );
  OAI21_X1 U13710 ( .B1(n12327), .B2(n11257), .A(n11256), .ZN(P3_U3223) );
  INV_X1 U13711 ( .A(n11258), .ZN(n11260) );
  OAI222_X1 U13712 ( .A1(n14738), .A2(P3_U3151), .B1(n12528), .B2(n11260), 
        .C1(n11259), .C2(n12530), .ZN(P3_U3268) );
  AND2_X1 U13713 ( .A1(n13331), .A2(n13478), .ZN(n11262) );
  AOI21_X1 U13714 ( .B1(n14525), .B2(n6443), .A(n11262), .ZN(n11340) );
  AOI22_X1 U13715 ( .A1(n14525), .A2(n7444), .B1(n6443), .B2(n13478), .ZN(
        n11263) );
  XNOR2_X1 U13716 ( .A(n11263), .B(n13365), .ZN(n11341) );
  NAND2_X1 U13717 ( .A1(n14235), .A2(n11264), .ZN(n11266) );
  OAI211_X1 U13718 ( .C1(n14241), .C2(n11267), .A(n11266), .B(n11265), .ZN(
        n11268) );
  AOI21_X1 U13719 ( .B1(n14525), .B2(n14238), .A(n11268), .ZN(n11269) );
  OAI21_X1 U13720 ( .B1(n11270), .B2(n14221), .A(n11269), .ZN(P1_U3231) );
  INV_X1 U13721 ( .A(n12391), .ZN(n12275) );
  INV_X1 U13722 ( .A(n11308), .ZN(n11271) );
  OAI22_X1 U13723 ( .A1(n14933), .A2(n11272), .B1(n11271), .B2(n12271), .ZN(
        n11275) );
  NOR2_X1 U13724 ( .A1(n11273), .A2(n14935), .ZN(n11274) );
  AOI211_X1 U13725 ( .C1(n12275), .C2(n11276), .A(n11275), .B(n11274), .ZN(
        n11277) );
  OAI21_X1 U13726 ( .B1(n12327), .B2(n11278), .A(n11277), .ZN(P3_U3224) );
  NOR2_X1 U13727 ( .A1(n11317), .A2(n6438), .ZN(n11280) );
  XNOR2_X1 U13728 ( .A(n14186), .B(n12576), .ZN(n11279) );
  NOR2_X1 U13729 ( .A1(n11279), .A2(n11280), .ZN(n11311) );
  AOI21_X1 U13730 ( .B1(n11280), .B2(n11279), .A(n11311), .ZN(n11285) );
  OAI21_X1 U13731 ( .B1(n11285), .B2(n11284), .A(n11313), .ZN(n11286) );
  NAND2_X1 U13732 ( .A1(n11286), .A2(n12689), .ZN(n11292) );
  OAI22_X1 U13733 ( .A1(n12658), .A2(n11288), .B1(n11287), .B2(n12720), .ZN(
        n11289) );
  AOI211_X1 U13734 ( .C1(n12685), .C2(n12732), .A(n11290), .B(n11289), .ZN(
        n11291) );
  OAI211_X1 U13735 ( .C1(n14186), .C2(n12653), .A(n11292), .B(n11291), .ZN(
        P2_U3196) );
  INV_X1 U13736 ( .A(n11661), .ZN(n11296) );
  AOI22_X1 U13737 ( .A1(n11293), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n13976), .ZN(n11294) );
  OAI21_X1 U13738 ( .B1(n11296), .B2(n13986), .A(n11294), .ZN(P1_U3330) );
  OAI222_X1 U13739 ( .A1(n13201), .A2(n11297), .B1(n13199), .B2(n11296), .C1(
        n11295), .C2(P2_U3088), .ZN(P2_U3302) );
  INV_X1 U13740 ( .A(n11298), .ZN(n11299) );
  AOI21_X1 U13741 ( .B1(n11301), .B2(n11300), .A(n11299), .ZN(n11310) );
  NOR2_X1 U13742 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11302), .ZN(n14870) );
  NOR2_X1 U13743 ( .A1(n11977), .A2(n11303), .ZN(n11304) );
  AOI211_X1 U13744 ( .C1(n11940), .C2(n11992), .A(n14870), .B(n11304), .ZN(
        n11305) );
  OAI21_X1 U13745 ( .B1(n11968), .B2(n11306), .A(n11305), .ZN(n11307) );
  AOI21_X1 U13746 ( .B1(n11308), .B2(n11972), .A(n11307), .ZN(n11309) );
  OAI21_X1 U13747 ( .B1(n11310), .B2(n11981), .A(n11309), .ZN(P3_U3171) );
  INV_X1 U13748 ( .A(n11311), .ZN(n11312) );
  XNOR2_X1 U13749 ( .A(n11314), .B(n6816), .ZN(n11409) );
  NOR2_X1 U13750 ( .A1(n11418), .A2(n6438), .ZN(n11411) );
  XNOR2_X1 U13751 ( .A(n11409), .B(n11411), .ZN(n11412) );
  XNOR2_X1 U13752 ( .A(n11413), .B(n11412), .ZN(n11321) );
  OAI22_X1 U13753 ( .A1(n12656), .A2(n11315), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10063), .ZN(n11319) );
  OAI22_X1 U13754 ( .A1(n12658), .A2(n11317), .B1(n11316), .B2(n12720), .ZN(
        n11318) );
  AOI211_X1 U13755 ( .C1(n11324), .C2(n12722), .A(n11319), .B(n11318), .ZN(
        n11320) );
  OAI21_X1 U13756 ( .B1(n11321), .B2(n12724), .A(n11320), .ZN(P2_U3206) );
  INV_X1 U13757 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11328) );
  AOI211_X1 U13758 ( .C1(n14660), .C2(n11324), .A(n11323), .B(n11322), .ZN(
        n11325) );
  OAI21_X1 U13759 ( .B1(n14655), .B2(n11326), .A(n11325), .ZN(n11329) );
  NAND2_X1 U13760 ( .A1(n11329), .A2(n14723), .ZN(n11327) );
  OAI21_X1 U13761 ( .B1(n14723), .B2(n11328), .A(n11327), .ZN(P2_U3469) );
  NAND2_X1 U13762 ( .A1(n11329), .A2(n14737), .ZN(n11330) );
  OAI21_X1 U13763 ( .B1(n14737), .B2(n7945), .A(n11330), .ZN(P2_U3512) );
  NAND2_X1 U13764 ( .A1(n14537), .A2(n7444), .ZN(n11332) );
  NAND2_X1 U13765 ( .A1(n13477), .A2(n6443), .ZN(n11331) );
  NAND2_X1 U13766 ( .A1(n11332), .A2(n11331), .ZN(n11333) );
  XNOR2_X1 U13767 ( .A(n11333), .B(n13318), .ZN(n11338) );
  INV_X1 U13768 ( .A(n11338), .ZN(n11336) );
  AND2_X1 U13769 ( .A1(n13331), .A2(n13477), .ZN(n11334) );
  AOI21_X1 U13770 ( .B1(n14537), .B2(n6443), .A(n11334), .ZN(n11337) );
  INV_X1 U13771 ( .A(n11337), .ZN(n11335) );
  NAND2_X1 U13772 ( .A1(n11336), .A2(n11335), .ZN(n14218) );
  NAND2_X1 U13773 ( .A1(n11338), .A2(n11337), .ZN(n13211) );
  NAND2_X1 U13774 ( .A1(n14218), .A2(n13211), .ZN(n11342) );
  XOR2_X1 U13775 ( .A(n11342), .B(n13212), .Z(n11350) );
  OAI21_X1 U13776 ( .B1(n14215), .B2(n11344), .A(n11343), .ZN(n11348) );
  OAI22_X1 U13777 ( .A1(n14214), .A2(n11346), .B1(n14241), .B2(n11345), .ZN(
        n11347) );
  AOI211_X1 U13778 ( .C1(n14537), .C2(n14238), .A(n11348), .B(n11347), .ZN(
        n11349) );
  OAI21_X1 U13779 ( .B1(n11350), .B2(n14221), .A(n11349), .ZN(P1_U3217) );
  OAI211_X1 U13780 ( .C1(n11353), .C2(n11352), .A(n11351), .B(n14923), .ZN(
        n11355) );
  AOI22_X1 U13781 ( .A1(n11866), .A2(n14919), .B1(n14920), .B2(n11920), .ZN(
        n11354) );
  OR2_X1 U13782 ( .A1(n11357), .A2(n11356), .ZN(n11358) );
  NAND2_X1 U13783 ( .A1(n11359), .A2(n11358), .ZN(n14168) );
  AOI22_X1 U13784 ( .A1(n14935), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n14929), 
        .B2(n11870), .ZN(n11360) );
  OAI21_X1 U13785 ( .B1(n12391), .B2(n11868), .A(n11360), .ZN(n11361) );
  AOI21_X1 U13786 ( .B1(n14168), .B2(n12393), .A(n11361), .ZN(n11362) );
  OAI21_X1 U13787 ( .B1(n14169), .B2(n14935), .A(n11362), .ZN(P3_U3221) );
  AOI21_X1 U13788 ( .B1(n11364), .B2(n11363), .A(n11981), .ZN(n11366) );
  NAND2_X1 U13789 ( .A1(n11366), .A2(n11365), .ZN(n11372) );
  AOI21_X1 U13790 ( .B1(n11974), .B2(n14887), .A(n11367), .ZN(n11368) );
  OAI21_X1 U13791 ( .B1(n11945), .B2(n11977), .A(n11368), .ZN(n11369) );
  AOI21_X1 U13792 ( .B1(n11979), .B2(n11370), .A(n11369), .ZN(n11371) );
  OAI211_X1 U13793 ( .C1(n11374), .C2(n11373), .A(n11372), .B(n11371), .ZN(
        P3_U3157) );
  XNOR2_X1 U13794 ( .A(n11375), .B(n11377), .ZN(n14173) );
  OAI211_X1 U13795 ( .C1(n11378), .C2(n11377), .A(n11376), .B(n14923), .ZN(
        n11380) );
  AOI22_X1 U13796 ( .A1(n14920), .A2(n11990), .B1(n11991), .B2(n14919), .ZN(
        n11379) );
  NAND2_X1 U13797 ( .A1(n11380), .A2(n11379), .ZN(n14171) );
  NAND2_X1 U13798 ( .A1(n14171), .A2(n14933), .ZN(n11383) );
  AND2_X1 U13799 ( .A1(n11381), .A2(n14960), .ZN(n14172) );
  AOI22_X1 U13800 ( .A1(n14896), .A2(n14172), .B1(n14929), .B2(n11948), .ZN(
        n11382) );
  OAI211_X1 U13801 ( .C1(n14933), .C2(n11384), .A(n11383), .B(n11382), .ZN(
        n11385) );
  AOI21_X1 U13802 ( .B1(n12393), .B2(n14173), .A(n11385), .ZN(n11386) );
  INV_X1 U13803 ( .A(n11386), .ZN(P3_U3222) );
  XNOR2_X1 U13804 ( .A(n11387), .B(n11394), .ZN(n11389) );
  NAND2_X1 U13805 ( .A1(n12731), .A2(n13002), .ZN(n11388) );
  OAI21_X1 U13806 ( .B1(n12648), .B2(n13057), .A(n11388), .ZN(n12716) );
  AOI21_X1 U13807 ( .B1(n11389), .B2(n13065), .A(n12716), .ZN(n13169) );
  AOI211_X1 U13808 ( .C1(n13167), .C2(n11390), .A(n10022), .B(n6441), .ZN(
        n13166) );
  INV_X1 U13809 ( .A(n12719), .ZN(n11391) );
  AOI22_X1 U13810 ( .A1(n13078), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11391), 
        .B2(n13081), .ZN(n11392) );
  OAI21_X1 U13811 ( .B1(n7014), .B2(n13073), .A(n11392), .ZN(n11396) );
  XOR2_X1 U13812 ( .A(n11394), .B(n11393), .Z(n13170) );
  NOR2_X1 U13813 ( .A1(n13170), .A2(n13053), .ZN(n11395) );
  AOI211_X1 U13814 ( .C1(n13166), .C2(n13085), .A(n11396), .B(n11395), .ZN(
        n11397) );
  OAI21_X1 U13815 ( .B1(n13078), .B2(n13169), .A(n11397), .ZN(P2_U3250) );
  XNOR2_X1 U13816 ( .A(n11398), .B(n11400), .ZN(n11399) );
  AOI222_X1 U13817 ( .A1(n14923), .A2(n11399), .B1(n11990), .B2(n14919), .C1(
        n11989), .C2(n14920), .ZN(n14165) );
  XNOR2_X1 U13818 ( .A(n11401), .B(n11400), .ZN(n14163) );
  INV_X1 U13819 ( .A(n14162), .ZN(n11403) );
  AOI22_X1 U13820 ( .A1(n14935), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n14929), 
        .B2(n11924), .ZN(n11402) );
  OAI21_X1 U13821 ( .B1(n12391), .B2(n11403), .A(n11402), .ZN(n11404) );
  AOI21_X1 U13822 ( .B1(n14163), .B2(n12393), .A(n11404), .ZN(n11405) );
  OAI21_X1 U13823 ( .B1(n14165), .B2(n14935), .A(n11405), .ZN(P3_U3220) );
  AND2_X1 U13824 ( .A1(n12731), .A2(n10022), .ZN(n11408) );
  XNOR2_X1 U13825 ( .A(n11406), .B(n6816), .ZN(n11407) );
  NOR2_X1 U13826 ( .A1(n11407), .A2(n11408), .ZN(n12532) );
  AOI21_X1 U13827 ( .B1(n11408), .B2(n11407), .A(n12532), .ZN(n11415) );
  INV_X1 U13828 ( .A(n11409), .ZN(n11410) );
  OAI21_X1 U13829 ( .B1(n11415), .B2(n11414), .A(n12534), .ZN(n11416) );
  NAND2_X1 U13830 ( .A1(n11416), .A2(n12689), .ZN(n11422) );
  NAND2_X1 U13831 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14574)
         );
  INV_X1 U13832 ( .A(n14574), .ZN(n11420) );
  OAI22_X1 U13833 ( .A1(n12658), .A2(n11418), .B1(n11417), .B2(n12720), .ZN(
        n11419) );
  AOI211_X1 U13834 ( .C1(n12685), .C2(n12730), .A(n11420), .B(n11419), .ZN(
        n11421) );
  OAI211_X1 U13835 ( .C1(n14180), .C2(n12653), .A(n11422), .B(n11421), .ZN(
        P2_U3187) );
  AND2_X1 U13836 ( .A1(n11425), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U13837 ( .A1(n11425), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U13838 ( .A1(n11425), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U13839 ( .A1(n11425), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U13840 ( .A1(n11425), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U13841 ( .A1(n11425), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U13842 ( .A1(n11425), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U13843 ( .A1(n11425), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U13844 ( .A1(n11425), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U13845 ( .A1(n11425), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U13846 ( .A1(n11425), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U13847 ( .A1(n11425), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U13848 ( .A1(n11425), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U13849 ( .A1(n11425), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U13850 ( .A1(n11425), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U13851 ( .A1(n11425), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U13852 ( .A1(n11425), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U13853 ( .A1(n11425), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U13854 ( .A1(n11425), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U13855 ( .A1(n11425), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U13856 ( .A1(n11425), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U13857 ( .A1(n11425), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U13858 ( .A1(n11425), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U13859 ( .A1(n11425), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U13860 ( .A1(n11425), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U13861 ( .A1(n11425), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U13862 ( .A1(n11425), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U13863 ( .A1(n11425), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U13864 ( .A1(n11425), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U13865 ( .A1(n11425), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  OAI222_X1 U13866 ( .A1(n11426), .A2(P2_U3088), .B1(n13199), .B2(n13981), 
        .C1(n11427), .C2(n13201), .ZN(P2_U3297) );
  INV_X1 U13867 ( .A(n11716), .ZN(n13983) );
  OAI222_X1 U13868 ( .A1(n11429), .A2(P2_U3088), .B1(n13199), .B2(n13983), 
        .C1(n11428), .C2(n13201), .ZN(P2_U3298) );
  NAND2_X1 U13869 ( .A1(n14414), .A2(n11430), .ZN(n11432) );
  NAND2_X1 U13870 ( .A1(n11432), .A2(n11431), .ZN(n11435) );
  NAND2_X1 U13871 ( .A1(n11435), .A2(n11433), .ZN(n11736) );
  OR2_X1 U13872 ( .A1(n11435), .A2(n11434), .ZN(n11436) );
  NAND2_X1 U13873 ( .A1(n11736), .A2(n11436), .ZN(n11449) );
  INV_X2 U13874 ( .A(n11449), .ZN(n11738) );
  XNOR2_X1 U13875 ( .A(n11437), .B(n11738), .ZN(n11438) );
  NOR2_X1 U13876 ( .A1(n11438), .A2(n11444), .ZN(n11443) );
  MUX2_X1 U13877 ( .A(n11440), .B(n11439), .S(n11719), .Z(n11442) );
  OAI211_X1 U13878 ( .C1(n11443), .C2(n11442), .A(n11441), .B(n14401), .ZN(
        n11457) );
  NAND4_X1 U13879 ( .A1(n11759), .A2(n11441), .A3(n11446), .A4(n11445), .ZN(
        n11456) );
  MUX2_X1 U13880 ( .A(n11448), .B(n11447), .S(n11719), .Z(n11455) );
  NAND2_X1 U13881 ( .A1(n6748), .A2(n11738), .ZN(n11452) );
  NAND3_X1 U13882 ( .A1(n13484), .A2(n11450), .A3(n11719), .ZN(n11451) );
  OAI21_X1 U13883 ( .B1(n13484), .B2(n11452), .A(n11451), .ZN(n11453) );
  NAND2_X1 U13884 ( .A1(n14401), .A2(n11453), .ZN(n11454) );
  NAND4_X1 U13885 ( .A1(n11457), .A2(n11456), .A3(n11455), .A4(n11454), .ZN(
        n11461) );
  INV_X1 U13886 ( .A(n11458), .ZN(n11460) );
  MUX2_X1 U13887 ( .A(n14485), .B(n13483), .S(n11719), .Z(n11459) );
  OAI21_X1 U13888 ( .B1(n11461), .B2(n11460), .A(n11459), .ZN(n11463) );
  NAND2_X1 U13889 ( .A1(n11461), .A2(n11460), .ZN(n11462) );
  NAND2_X1 U13890 ( .A1(n11463), .A2(n11462), .ZN(n11467) );
  MUX2_X1 U13891 ( .A(n13482), .B(n11464), .S(n11738), .Z(n11466) );
  MUX2_X1 U13892 ( .A(n13482), .B(n11464), .S(n11719), .Z(n11465) );
  MUX2_X1 U13893 ( .A(n13481), .B(n14393), .S(n11719), .Z(n11471) );
  NAND2_X1 U13894 ( .A1(n11470), .A2(n11471), .ZN(n11469) );
  MUX2_X1 U13895 ( .A(n14393), .B(n13481), .S(n11719), .Z(n11468) );
  NAND2_X1 U13896 ( .A1(n11469), .A2(n11468), .ZN(n11475) );
  INV_X1 U13897 ( .A(n11471), .ZN(n11472) );
  NAND2_X1 U13898 ( .A1(n11473), .A2(n11472), .ZN(n11474) );
  MUX2_X1 U13899 ( .A(n13480), .B(n14506), .S(n11738), .Z(n11477) );
  MUX2_X1 U13900 ( .A(n14506), .B(n13480), .S(n11738), .Z(n11476) );
  MUX2_X1 U13901 ( .A(n13479), .B(n14515), .S(n11719), .Z(n11479) );
  MUX2_X1 U13902 ( .A(n13479), .B(n14515), .S(n11738), .Z(n11478) );
  MUX2_X1 U13903 ( .A(n13478), .B(n14525), .S(n11738), .Z(n11483) );
  NAND2_X1 U13904 ( .A1(n11482), .A2(n11483), .ZN(n11481) );
  MUX2_X1 U13905 ( .A(n13478), .B(n14525), .S(n11719), .Z(n11480) );
  NAND2_X1 U13906 ( .A1(n11481), .A2(n11480), .ZN(n11487) );
  INV_X1 U13907 ( .A(n11482), .ZN(n11485) );
  INV_X1 U13908 ( .A(n11483), .ZN(n11484) );
  NAND2_X1 U13909 ( .A1(n11485), .A2(n11484), .ZN(n11486) );
  NAND2_X1 U13910 ( .A1(n11487), .A2(n11486), .ZN(n11489) );
  MUX2_X1 U13911 ( .A(n13477), .B(n14537), .S(n11719), .Z(n11490) );
  MUX2_X1 U13912 ( .A(n13477), .B(n14537), .S(n11738), .Z(n11488) );
  INV_X1 U13913 ( .A(n11490), .ZN(n11491) );
  MUX2_X1 U13914 ( .A(n13476), .B(n14226), .S(n11738), .Z(n11493) );
  MUX2_X1 U13915 ( .A(n13476), .B(n14226), .S(n11449), .Z(n11492) );
  MUX2_X1 U13916 ( .A(n13475), .B(n14120), .S(n11719), .Z(n11498) );
  MUX2_X1 U13917 ( .A(n13475), .B(n14120), .S(n11738), .Z(n11495) );
  NAND2_X1 U13918 ( .A1(n11496), .A2(n11495), .ZN(n11501) );
  INV_X1 U13919 ( .A(n11497), .ZN(n11499) );
  NAND2_X1 U13920 ( .A1(n11499), .A2(n6894), .ZN(n11500) );
  MUX2_X1 U13921 ( .A(n13474), .B(n13433), .S(n11738), .Z(n11504) );
  AND2_X1 U13922 ( .A1(n11510), .A2(n11502), .ZN(n11503) );
  AND2_X1 U13923 ( .A1(n13655), .A2(n13433), .ZN(n11505) );
  MUX2_X1 U13924 ( .A(n13474), .B(n11505), .S(n11719), .Z(n11506) );
  NAND2_X1 U13925 ( .A1(n13655), .A2(n11508), .ZN(n11509) );
  OR2_X1 U13926 ( .A1(n11510), .A2(n11449), .ZN(n11530) );
  NAND2_X1 U13927 ( .A1(n11511), .A2(n11743), .ZN(n11513) );
  AOI22_X1 U13928 ( .A1(n11744), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11556), 
        .B2(n13585), .ZN(n11512) );
  MUX2_X1 U13929 ( .A(n13866), .B(n14271), .S(n11738), .Z(n11550) );
  OR2_X1 U13930 ( .A1(n11514), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n11515) );
  NAND2_X1 U13931 ( .A1(n11559), .A2(n11515), .ZN(n13863) );
  OR2_X1 U13932 ( .A1(n11731), .A2(n11132), .ZN(n11517) );
  OR2_X1 U13933 ( .A1(n6743), .A2(n15023), .ZN(n11516) );
  AND2_X1 U13934 ( .A1(n11517), .A2(n11516), .ZN(n11519) );
  NAND2_X1 U13935 ( .A1(n11726), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11518) );
  OAI211_X1 U13936 ( .C1(n13863), .C2(n11634), .A(n11519), .B(n11518), .ZN(
        n13658) );
  NAND2_X1 U13937 ( .A1(n11550), .A2(n13658), .ZN(n11523) );
  INV_X1 U13938 ( .A(n13866), .ZN(n13411) );
  NAND2_X1 U13939 ( .A1(n13411), .A2(n11738), .ZN(n11525) );
  NAND2_X1 U13940 ( .A1(n11520), .A2(n11743), .ZN(n11522) );
  AOI22_X1 U13941 ( .A1(n11744), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11556), 
        .B2(n13598), .ZN(n11521) );
  AOI21_X1 U13942 ( .B1(n11523), .B2(n11525), .A(n14265), .ZN(n11529) );
  INV_X1 U13943 ( .A(n13658), .ZN(n14209) );
  NAND2_X1 U13944 ( .A1(n11550), .A2(n14209), .ZN(n11524) );
  OR2_X1 U13945 ( .A1(n14271), .A2(n11738), .ZN(n11543) );
  AOI21_X1 U13946 ( .B1(n11524), .B2(n11543), .A(n13659), .ZN(n11528) );
  NAND2_X1 U13947 ( .A1(n13658), .A2(n11719), .ZN(n11545) );
  OR2_X1 U13948 ( .A1(n14271), .A2(n11545), .ZN(n11527) );
  INV_X1 U13949 ( .A(n11525), .ZN(n11549) );
  NAND2_X1 U13950 ( .A1(n11549), .A2(n14209), .ZN(n11526) );
  NAND2_X1 U13951 ( .A1(n11527), .A2(n11526), .ZN(n11547) );
  AOI21_X1 U13952 ( .B1(n11531), .B2(n11530), .A(n7574), .ZN(n11532) );
  INV_X1 U13953 ( .A(n11532), .ZN(n11574) );
  NAND2_X1 U13954 ( .A1(n11533), .A2(n11743), .ZN(n11535) );
  AOI22_X1 U13955 ( .A1(n11744), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14414), 
        .B2(n11556), .ZN(n11534) );
  INV_X1 U13956 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n11537) );
  INV_X1 U13957 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n11536) );
  OAI21_X1 U13958 ( .B1(n11559), .B2(n11537), .A(n11536), .ZN(n11539) );
  NAND2_X1 U13959 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n11538) );
  NAND2_X1 U13960 ( .A1(n11539), .A2(n11575), .ZN(n13837) );
  OR2_X1 U13961 ( .A1(n13837), .A2(n11634), .ZN(n11542) );
  AOI22_X1 U13962 ( .A1(n15191), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n11726), 
        .B2(P1_REG0_REG_19__SCAN_IN), .ZN(n11541) );
  INV_X1 U13963 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n13597) );
  OR2_X1 U13964 ( .A1(n6743), .A2(n13597), .ZN(n11540) );
  NAND2_X1 U13965 ( .A1(n11568), .A2(n13848), .ZN(n13662) );
  INV_X1 U13966 ( .A(n11543), .ZN(n11544) );
  NAND2_X1 U13967 ( .A1(n11550), .A2(n11544), .ZN(n11546) );
  NAND2_X1 U13968 ( .A1(n11546), .A2(n11545), .ZN(n11548) );
  AOI22_X1 U13969 ( .A1(n11548), .A2(n14265), .B1(n11550), .B2(n11547), .ZN(
        n11554) );
  NAND2_X1 U13970 ( .A1(n11550), .A2(n11549), .ZN(n11551) );
  OAI21_X1 U13971 ( .B1(n13658), .B2(n11719), .A(n11551), .ZN(n11552) );
  NAND2_X1 U13972 ( .A1(n11552), .A2(n13659), .ZN(n11553) );
  NAND4_X1 U13973 ( .A1(n11567), .A2(n13662), .A3(n11554), .A4(n11553), .ZN(
        n11566) );
  NAND2_X1 U13974 ( .A1(n11555), .A2(n11743), .ZN(n11558) );
  AOI22_X1 U13975 ( .A1(n6451), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11556), 
        .B2(n13601), .ZN(n11557) );
  XNOR2_X1 U13976 ( .A(n11559), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n13852) );
  NAND2_X1 U13977 ( .A1(n13852), .A2(n11621), .ZN(n11565) );
  INV_X1 U13978 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n11562) );
  NAND2_X1 U13979 ( .A1(n15191), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n11561) );
  NAND2_X1 U13980 ( .A1(n11726), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n11560) );
  OAI211_X1 U13981 ( .C1(n6743), .C2(n11562), .A(n11561), .B(n11560), .ZN(
        n11563) );
  INV_X1 U13982 ( .A(n11563), .ZN(n11564) );
  XNOR2_X1 U13983 ( .A(n13860), .B(n13864), .ZN(n13846) );
  OR2_X1 U13984 ( .A1(n13662), .A2(n11738), .ZN(n11571) );
  NAND4_X1 U13985 ( .A1(n11567), .A2(n13864), .A3(n11719), .A4(n13860), .ZN(
        n11570) );
  OR3_X1 U13986 ( .A1(n11568), .A2(n13848), .A3(n11719), .ZN(n11569) );
  INV_X1 U13987 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13428) );
  AND2_X1 U13988 ( .A1(n11575), .A2(n13428), .ZN(n11576) );
  OR2_X1 U13989 ( .A1(n11576), .A2(n11590), .ZN(n13824) );
  AOI22_X1 U13990 ( .A1(n11711), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n15191), 
        .B2(P1_REG2_REG_20__SCAN_IN), .ZN(n11578) );
  NAND2_X1 U13991 ( .A1(n11726), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11577) );
  OAI211_X1 U13992 ( .C1(n13824), .C2(n11634), .A(n11578), .B(n11577), .ZN(
        n13836) );
  NAND2_X1 U13993 ( .A1(n11744), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n11580) );
  MUX2_X1 U13994 ( .A(n13836), .B(n13950), .S(n11738), .Z(n11584) );
  NAND2_X1 U13995 ( .A1(n11585), .A2(n11584), .ZN(n11583) );
  MUX2_X1 U13996 ( .A(n13836), .B(n13950), .S(n11449), .Z(n11582) );
  NAND2_X1 U13997 ( .A1(n11583), .A2(n11582), .ZN(n11589) );
  INV_X1 U13998 ( .A(n11584), .ZN(n11587) );
  INV_X1 U13999 ( .A(n11585), .ZN(n11586) );
  NAND2_X1 U14000 ( .A1(n11587), .A2(n11586), .ZN(n11588) );
  NOR2_X1 U14001 ( .A1(n11590), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11591) );
  OR2_X1 U14002 ( .A1(n11602), .A2(n11591), .ZN(n13803) );
  INV_X1 U14003 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n11594) );
  NAND2_X1 U14004 ( .A1(n11726), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11593) );
  NAND2_X1 U14005 ( .A1(n15191), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11592) );
  OAI211_X1 U14006 ( .C1(n11594), .C2(n6743), .A(n11593), .B(n11592), .ZN(
        n11595) );
  INV_X1 U14007 ( .A(n11595), .ZN(n11596) );
  OAI21_X1 U14008 ( .B1(n13803), .B2(n11634), .A(n11596), .ZN(n13641) );
  NAND2_X1 U14009 ( .A1(n11597), .A2(n11743), .ZN(n11599) );
  NAND2_X1 U14010 ( .A1(n6451), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n11598) );
  MUX2_X1 U14011 ( .A(n13641), .B(n13945), .S(n11719), .Z(n11601) );
  MUX2_X1 U14012 ( .A(n13945), .B(n13641), .S(n11719), .Z(n11600) );
  NOR2_X1 U14013 ( .A1(n11602), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11603) );
  OR2_X1 U14014 ( .A1(n11619), .A2(n11603), .ZN(n13791) );
  INV_X1 U14015 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n11606) );
  NAND2_X1 U14016 ( .A1(n11726), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11605) );
  NAND2_X1 U14017 ( .A1(n15191), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11604) );
  OAI211_X1 U14018 ( .C1(n11606), .C2(n6743), .A(n11605), .B(n11604), .ZN(
        n11607) );
  INV_X1 U14019 ( .A(n11607), .ZN(n11608) );
  OAI21_X1 U14020 ( .B1(n13791), .B2(n11634), .A(n11608), .ZN(n13666) );
  OR2_X1 U14021 ( .A1(n11610), .A2(n11609), .ZN(n11611) );
  XNOR2_X1 U14022 ( .A(n11611), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n13994) );
  MUX2_X1 U14023 ( .A(n13666), .B(n13793), .S(n11738), .Z(n11613) );
  NAND2_X1 U14024 ( .A1(n11614), .A2(n11613), .ZN(n11616) );
  MUX2_X1 U14025 ( .A(n13666), .B(n13793), .S(n11449), .Z(n11615) );
  NAND2_X1 U14026 ( .A1(n11616), .A2(n11615), .ZN(n11617) );
  OR2_X1 U14027 ( .A1(n11619), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11620) );
  NAND2_X1 U14028 ( .A1(n11619), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11632) );
  AND2_X1 U14029 ( .A1(n11620), .A2(n11632), .ZN(n13777) );
  NAND2_X1 U14030 ( .A1(n13777), .A2(n11621), .ZN(n11626) );
  INV_X1 U14031 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n13775) );
  NAND2_X1 U14032 ( .A1(n11726), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11623) );
  NAND2_X1 U14033 ( .A1(n11711), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n11622) );
  OAI211_X1 U14034 ( .C1(n11731), .C2(n13775), .A(n11623), .B(n11622), .ZN(
        n11624) );
  INV_X1 U14035 ( .A(n11624), .ZN(n11625) );
  NAND2_X1 U14036 ( .A1(n11626), .A2(n11625), .ZN(n13667) );
  NAND2_X1 U14037 ( .A1(n11744), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11628) );
  MUX2_X1 U14038 ( .A(n13667), .B(n13780), .S(n11719), .Z(n11631) );
  MUX2_X1 U14039 ( .A(n13667), .B(n13780), .S(n11738), .Z(n11630) );
  NAND2_X1 U14040 ( .A1(n11726), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11639) );
  INV_X1 U14041 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n13765) );
  OR2_X1 U14042 ( .A1(n11731), .A2(n13765), .ZN(n11638) );
  INV_X1 U14043 ( .A(n11632), .ZN(n11633) );
  NAND2_X1 U14044 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n11633), .ZN(n11654) );
  OAI21_X1 U14045 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11633), .A(n11654), 
        .ZN(n13764) );
  OR2_X1 U14046 ( .A1(n11634), .A2(n13764), .ZN(n11637) );
  INV_X1 U14047 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n11635) );
  OR2_X1 U14048 ( .A1(n6743), .A2(n11635), .ZN(n11636) );
  NAND4_X1 U14049 ( .A1(n11639), .A2(n11638), .A3(n11637), .A4(n11636), .ZN(
        n13645) );
  NAND2_X1 U14050 ( .A1(n11640), .A2(n11743), .ZN(n11642) );
  NAND2_X1 U14051 ( .A1(n6451), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n11641) );
  MUX2_X1 U14052 ( .A(n13645), .B(n13926), .S(n11738), .Z(n11646) );
  NAND2_X1 U14053 ( .A1(n11645), .A2(n11646), .ZN(n11644) );
  MUX2_X1 U14054 ( .A(n13645), .B(n13926), .S(n11719), .Z(n11643) );
  NAND2_X1 U14055 ( .A1(n11644), .A2(n11643), .ZN(n11650) );
  INV_X1 U14056 ( .A(n11645), .ZN(n11648) );
  INV_X1 U14057 ( .A(n11646), .ZN(n11647) );
  NAND2_X1 U14058 ( .A1(n11648), .A2(n11647), .ZN(n11649) );
  NAND2_X1 U14059 ( .A1(n15191), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11660) );
  INV_X1 U14060 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n11651) );
  OR2_X1 U14061 ( .A1(n11044), .A2(n11651), .ZN(n11659) );
  INV_X1 U14062 ( .A(n11654), .ZN(n11652) );
  NAND2_X1 U14063 ( .A1(n11652), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11668) );
  INV_X1 U14064 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n11653) );
  NAND2_X1 U14065 ( .A1(n11654), .A2(n11653), .ZN(n11655) );
  NAND2_X1 U14066 ( .A1(n11668), .A2(n11655), .ZN(n13743) );
  OR2_X1 U14067 ( .A1(n11634), .A2(n13743), .ZN(n11658) );
  INV_X1 U14068 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n11656) );
  OR2_X1 U14069 ( .A1(n6743), .A2(n11656), .ZN(n11657) );
  NAND4_X1 U14070 ( .A1(n11660), .A2(n11659), .A3(n11658), .A4(n11657), .ZN(
        n13654) );
  NAND2_X1 U14071 ( .A1(n11661), .A2(n11743), .ZN(n11663) );
  NAND2_X1 U14072 ( .A1(n6451), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n11662) );
  MUX2_X1 U14073 ( .A(n13654), .B(n13919), .S(n11719), .Z(n11665) );
  MUX2_X1 U14074 ( .A(n13654), .B(n13919), .S(n11738), .Z(n11664) );
  NAND2_X1 U14075 ( .A1(n15191), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n11674) );
  INV_X1 U14076 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n11666) );
  OR2_X1 U14077 ( .A1(n11044), .A2(n11666), .ZN(n11673) );
  INV_X1 U14078 ( .A(n11668), .ZN(n11667) );
  NAND2_X1 U14079 ( .A1(n11667), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11683) );
  INV_X1 U14080 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13462) );
  NAND2_X1 U14081 ( .A1(n11668), .A2(n13462), .ZN(n11669) );
  NAND2_X1 U14082 ( .A1(n11683), .A2(n11669), .ZN(n13730) );
  OR2_X1 U14083 ( .A1(n11634), .A2(n13730), .ZN(n11672) );
  INV_X1 U14084 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n11670) );
  OR2_X1 U14085 ( .A1(n6743), .A2(n11670), .ZN(n11671) );
  NAND4_X1 U14086 ( .A1(n11674), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(
        n13671) );
  NAND2_X1 U14087 ( .A1(n13200), .A2(n11743), .ZN(n11676) );
  NAND2_X1 U14088 ( .A1(n6451), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n11675) );
  MUX2_X1 U14089 ( .A(n13671), .B(n13648), .S(n11738), .Z(n11678) );
  MUX2_X1 U14090 ( .A(n13671), .B(n13648), .S(n11719), .Z(n11677) );
  INV_X1 U14091 ( .A(n11678), .ZN(n11679) );
  NAND2_X1 U14092 ( .A1(n11726), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11689) );
  INV_X1 U14093 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n11680) );
  OR2_X1 U14094 ( .A1(n11731), .A2(n11680), .ZN(n11688) );
  INV_X1 U14095 ( .A(n11683), .ZN(n11681) );
  NAND2_X1 U14096 ( .A1(n11681), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11700) );
  INV_X1 U14097 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11682) );
  NAND2_X1 U14098 ( .A1(n11683), .A2(n11682), .ZN(n11684) );
  NAND2_X1 U14099 ( .A1(n11700), .A2(n11684), .ZN(n13716) );
  OR2_X1 U14100 ( .A1(n11634), .A2(n13716), .ZN(n11687) );
  INV_X1 U14101 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n11685) );
  OR2_X1 U14102 ( .A1(n6743), .A2(n11685), .ZN(n11686) );
  NAND2_X1 U14103 ( .A1(n11744), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11690) );
  MUX2_X1 U14104 ( .A(n13651), .B(n13719), .S(n11738), .Z(n11694) );
  NAND2_X1 U14105 ( .A1(n11693), .A2(n11694), .ZN(n11692) );
  MUX2_X1 U14106 ( .A(n13651), .B(n13719), .S(n11719), .Z(n11691) );
  NAND2_X1 U14107 ( .A1(n11692), .A2(n11691), .ZN(n11698) );
  INV_X1 U14108 ( .A(n11693), .ZN(n11696) );
  INV_X1 U14109 ( .A(n11694), .ZN(n11695) );
  NAND2_X1 U14110 ( .A1(n11696), .A2(n11695), .ZN(n11697) );
  NAND2_X1 U14111 ( .A1(n11726), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11706) );
  INV_X1 U14112 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n13698) );
  OR2_X1 U14113 ( .A1(n11731), .A2(n13698), .ZN(n11705) );
  INV_X1 U14114 ( .A(n11700), .ZN(n11699) );
  NAND2_X1 U14115 ( .A1(n11699), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13678) );
  INV_X1 U14116 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13372) );
  NAND2_X1 U14117 ( .A1(n11700), .A2(n13372), .ZN(n11701) );
  NAND2_X1 U14118 ( .A1(n13678), .A2(n11701), .ZN(n13697) );
  OR2_X1 U14119 ( .A1(n11634), .A2(n13697), .ZN(n11704) );
  INV_X1 U14120 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n11702) );
  OR2_X1 U14121 ( .A1(n6743), .A2(n11702), .ZN(n11703) );
  NAND2_X1 U14122 ( .A1(n13192), .A2(n11743), .ZN(n11708) );
  NAND2_X1 U14123 ( .A1(n6451), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n11707) );
  MUX2_X1 U14124 ( .A(n13675), .B(n13700), .S(n11738), .Z(n11710) );
  MUX2_X1 U14125 ( .A(n13472), .B(n13898), .S(n11719), .Z(n11709) );
  NAND2_X1 U14126 ( .A1(n11726), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n11715) );
  NAND2_X1 U14127 ( .A1(n11711), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11714) );
  INV_X1 U14128 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n15049) );
  OR2_X1 U14129 ( .A1(n11731), .A2(n15049), .ZN(n11713) );
  OR2_X1 U14130 ( .A1(n11634), .A2(n13678), .ZN(n11712) );
  NAND4_X1 U14131 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n13693) );
  NAND2_X1 U14132 ( .A1(n11716), .A2(n11743), .ZN(n11718) );
  NAND2_X1 U14133 ( .A1(n11744), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11717) );
  MUX2_X1 U14134 ( .A(n13693), .B(n13890), .S(n11719), .Z(n11720) );
  MUX2_X1 U14135 ( .A(n13890), .B(n13693), .S(n11719), .Z(n11722) );
  INV_X1 U14136 ( .A(n11720), .ZN(n11721) );
  NAND2_X1 U14137 ( .A1(n6451), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11724) );
  INV_X1 U14138 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U14139 ( .A1(n15191), .A2(P1_REG2_REG_30__SCAN_IN), .B1(n11726), 
        .B2(P1_REG0_REG_30__SCAN_IN), .ZN(n11728) );
  OAI21_X1 U14140 ( .B1(n6743), .B2(n11729), .A(n11728), .ZN(n13471) );
  INV_X1 U14141 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n15094) );
  OR2_X1 U14142 ( .A1(n6743), .A2(n15094), .ZN(n11735) );
  INV_X1 U14143 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n13618) );
  OR2_X1 U14144 ( .A1(n11731), .A2(n13618), .ZN(n11734) );
  INV_X1 U14145 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n11732) );
  OR2_X1 U14146 ( .A1(n11044), .A2(n11732), .ZN(n11733) );
  AND3_X1 U14147 ( .A1(n11735), .A2(n11734), .A3(n11733), .ZN(n13617) );
  OAI21_X1 U14148 ( .B1(n13617), .B2(n11738), .A(n11736), .ZN(n11737) );
  AOI22_X1 U14149 ( .A1(n13626), .A2(n11738), .B1(n13471), .B2(n11737), .ZN(
        n11741) );
  INV_X1 U14150 ( .A(n13617), .ZN(n13470) );
  OAI21_X1 U14151 ( .B1(n13470), .B2(n11739), .A(n13471), .ZN(n11740) );
  MUX2_X1 U14152 ( .A(n11740), .B(n13887), .S(n11719), .Z(n11742) );
  NAND2_X1 U14153 ( .A1(n13187), .A2(n11743), .ZN(n11746) );
  NAND2_X1 U14154 ( .A1(n11744), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n11745) );
  XNOR2_X1 U14155 ( .A(n13881), .B(n13617), .ZN(n11778) );
  NAND2_X1 U14156 ( .A1(n11748), .A2(n11747), .ZN(n11749) );
  NAND2_X1 U14157 ( .A1(n14410), .A2(n11749), .ZN(n11783) );
  NOR3_X1 U14158 ( .A1(n11750), .A2(n11778), .A3(n11783), .ZN(n11791) );
  NOR2_X1 U14159 ( .A1(n13881), .A2(n13617), .ZN(n11752) );
  INV_X1 U14160 ( .A(n13881), .ZN(n13615) );
  NOR2_X1 U14161 ( .A1(n13615), .A2(n13470), .ZN(n11751) );
  MUX2_X1 U14162 ( .A(n11752), .B(n11751), .S(n11719), .Z(n11786) );
  NAND2_X1 U14163 ( .A1(n11783), .A2(n11781), .ZN(n11784) );
  INV_X1 U14164 ( .A(n11784), .ZN(n11753) );
  INV_X1 U14165 ( .A(n13471), .ZN(n13677) );
  XNOR2_X1 U14166 ( .A(n13626), .B(n13677), .ZN(n11777) );
  NAND2_X1 U14167 ( .A1(n13898), .A2(n13472), .ZN(n13652) );
  OR2_X1 U14168 ( .A1(n13898), .A2(n13472), .ZN(n11754) );
  NAND2_X1 U14169 ( .A1(n13906), .A2(n13651), .ZN(n13689) );
  OR2_X1 U14170 ( .A1(n13906), .A2(n13651), .ZN(n11755) );
  NAND2_X1 U14171 ( .A1(n13689), .A2(n11755), .ZN(n13650) );
  INV_X1 U14172 ( .A(n13645), .ZN(n13739) );
  OR2_X1 U14173 ( .A1(n13926), .A2(n13739), .ZN(n13669) );
  NAND2_X1 U14174 ( .A1(n13926), .A2(n13739), .ZN(n11756) );
  NAND2_X1 U14175 ( .A1(n13669), .A2(n11756), .ZN(n13644) );
  INV_X1 U14176 ( .A(n13641), .ZN(n13817) );
  XNOR2_X1 U14177 ( .A(n13945), .B(n13817), .ZN(n13665) );
  XNOR2_X1 U14178 ( .A(n13950), .B(n13836), .ZN(n13663) );
  XNOR2_X1 U14179 ( .A(n14271), .B(n13411), .ZN(n14249) );
  OR2_X1 U14180 ( .A1(n13659), .A2(n13658), .ZN(n13632) );
  NAND2_X1 U14181 ( .A1(n13659), .A2(n13658), .ZN(n13634) );
  NAND2_X1 U14182 ( .A1(n13632), .A2(n13634), .ZN(n13872) );
  NAND4_X1 U14183 ( .A1(n11759), .A2(n11441), .A3(n11758), .A4(n11757), .ZN(
        n11760) );
  NOR4_X1 U14184 ( .A1(n11762), .A2(n11761), .A3(n14384), .A4(n11760), .ZN(
        n11764) );
  NAND2_X1 U14185 ( .A1(n11764), .A2(n11763), .ZN(n11765) );
  NOR4_X1 U14186 ( .A1(n11768), .A2(n11767), .A3(n11766), .A4(n11765), .ZN(
        n11770) );
  NAND4_X1 U14187 ( .A1(n13872), .A2(n11770), .A3(n11769), .A4(n14114), .ZN(
        n11772) );
  NOR4_X1 U14188 ( .A1(n14249), .A2(n7206), .A3(n11772), .A4(n11771), .ZN(
        n11773) );
  INV_X1 U14189 ( .A(n13846), .ZN(n13661) );
  NAND4_X1 U14190 ( .A1(n13663), .A2(n13830), .A3(n11773), .A4(n13661), .ZN(
        n11774) );
  XNOR2_X1 U14191 ( .A(n13939), .B(n13666), .ZN(n13785) );
  NOR4_X1 U14192 ( .A1(n13644), .A2(n13665), .A3(n11774), .A4(n13785), .ZN(
        n11775) );
  XNOR2_X1 U14193 ( .A(n13919), .B(n13654), .ZN(n13747) );
  NAND4_X1 U14194 ( .A1(n11775), .A2(n7172), .A3(n13747), .A4(n13772), .ZN(
        n11776) );
  NOR4_X1 U14195 ( .A1(n11777), .A2(n13704), .A3(n13650), .A4(n11776), .ZN(
        n11779) );
  INV_X1 U14196 ( .A(n11778), .ZN(n11785) );
  NAND3_X1 U14197 ( .A1(n11779), .A2(n11785), .A3(n13672), .ZN(n11780) );
  XNOR2_X1 U14198 ( .A(n11780), .B(n13822), .ZN(n11782) );
  NOR2_X1 U14199 ( .A1(n11782), .A2(n11781), .ZN(n11789) );
  INV_X1 U14200 ( .A(n11783), .ZN(n11788) );
  NOR2_X1 U14201 ( .A1(n11785), .A2(n11784), .ZN(n11787) );
  NOR2_X1 U14202 ( .A1(n11791), .A2(n11790), .ZN(n11796) );
  NOR3_X1 U14203 ( .A1(n11792), .A2(n14344), .A3(n14382), .ZN(n11794) );
  OAI21_X1 U14204 ( .B1(n11795), .B2(n13995), .A(P1_B_REG_SCAN_IN), .ZN(n11793) );
  OAI22_X1 U14205 ( .A1(n11796), .A2(n11795), .B1(n11794), .B2(n11793), .ZN(
        P1_U3242) );
  OR3_X1 U14206 ( .A1(n11798), .A2(n14960), .A3(n11797), .ZN(n11799) );
  OAI21_X1 U14207 ( .B1(n9066), .B2(n14901), .A(n11799), .ZN(n11806) );
  INV_X1 U14208 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n11800) );
  NOR2_X1 U14209 ( .A1(n14974), .A2(n11800), .ZN(n11801) );
  AOI21_X1 U14210 ( .B1(n14974), .B2(n11806), .A(n11801), .ZN(n11802) );
  OAI21_X1 U14211 ( .B1(n11809), .B2(n12510), .A(n11802), .ZN(P3_U3390) );
  NOR2_X1 U14212 ( .A1(n14990), .A2(n11803), .ZN(n11804) );
  AOI21_X1 U14213 ( .B1(n11806), .B2(n14990), .A(n11804), .ZN(n11805) );
  OAI21_X1 U14214 ( .B1(n11809), .B2(n12459), .A(n11805), .ZN(P3_U3459) );
  AOI21_X1 U14215 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n14929), .A(n11806), .ZN(
        n11807) );
  MUX2_X1 U14216 ( .A(n11807), .B(n14739), .S(n14935), .Z(n11808) );
  OAI21_X1 U14217 ( .B1(n11809), .B2(n12391), .A(n11808), .ZN(P3_U3233) );
  XNOR2_X1 U14218 ( .A(n12199), .B(n6435), .ZN(n11816) );
  INV_X1 U14219 ( .A(n11816), .ZN(n11810) );
  NAND2_X1 U14220 ( .A1(n11810), .A2(n11963), .ZN(n11821) );
  INV_X1 U14221 ( .A(n11811), .ZN(n11812) );
  AOI22_X1 U14222 ( .A1(n12201), .A2(n11940), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11814) );
  NAND2_X1 U14223 ( .A1(n12207), .A2(n11972), .ZN(n11813) );
  OAI211_X1 U14224 ( .C1(n12204), .C2(n11977), .A(n11814), .B(n11813), .ZN(
        n11818) );
  NOR4_X1 U14225 ( .A1(n11816), .A2(n11981), .A3(n11815), .A4(n12201), .ZN(
        n11817) );
  AOI211_X1 U14226 ( .C1(n11979), .C2(n11819), .A(n11818), .B(n11817), .ZN(
        n11820) );
  INV_X1 U14227 ( .A(n11822), .ZN(n11823) );
  XNOR2_X1 U14228 ( .A(n11827), .B(n11826), .ZN(n11832) );
  NAND2_X1 U14229 ( .A1(n11972), .A2(n12389), .ZN(n11829) );
  AND2_X1 U14230 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12070) );
  AOI21_X1 U14231 ( .B1(n11940), .B2(n11920), .A(n12070), .ZN(n11828) );
  OAI211_X1 U14232 ( .C1(n12385), .C2(n11977), .A(n11829), .B(n11828), .ZN(
        n11830) );
  AOI21_X1 U14233 ( .B1(n12388), .B2(n11979), .A(n11830), .ZN(n11831) );
  OAI21_X1 U14234 ( .B1(n11832), .B2(n11981), .A(n11831), .ZN(P3_U3155) );
  AOI21_X1 U14235 ( .B1(n11835), .B2(n11834), .A(n11902), .ZN(n11840) );
  AOI22_X1 U14236 ( .A1(n11987), .A2(n11974), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11837) );
  NAND2_X1 U14237 ( .A1(n11972), .A2(n12270), .ZN(n11836) );
  OAI211_X1 U14238 ( .C1(n12266), .C2(n11977), .A(n11837), .B(n11836), .ZN(
        n11838) );
  AOI21_X1 U14239 ( .B1(n12276), .B2(n11979), .A(n11838), .ZN(n11839) );
  OAI21_X1 U14240 ( .B1(n11840), .B2(n11981), .A(n11839), .ZN(P3_U3156) );
  XNOR2_X1 U14241 ( .A(n11842), .B(n11841), .ZN(n11847) );
  NAND2_X1 U14242 ( .A1(n11974), .A2(n12344), .ZN(n11843) );
  NAND2_X1 U14243 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12176)
         );
  OAI211_X1 U14244 ( .C1(n11977), .C2(n12295), .A(n11843), .B(n12176), .ZN(
        n11845) );
  NOR2_X1 U14245 ( .A1(n12496), .A2(n11968), .ZN(n11844) );
  AOI211_X1 U14246 ( .C1(n12322), .C2(n11972), .A(n11845), .B(n11844), .ZN(
        n11846) );
  OAI21_X1 U14247 ( .B1(n11847), .B2(n11981), .A(n11846), .ZN(P3_U3159) );
  NAND2_X1 U14248 ( .A1(n11910), .A2(n11848), .ZN(n11850) );
  AND2_X1 U14249 ( .A1(n11850), .A2(n11849), .ZN(n11853) );
  INV_X1 U14250 ( .A(n11851), .ZN(n11852) );
  AOI21_X1 U14251 ( .B1(n11854), .B2(n11853), .A(n11852), .ZN(n11859) );
  NAND2_X1 U14252 ( .A1(n11972), .A2(n12299), .ZN(n11856) );
  AOI22_X1 U14253 ( .A1(n11940), .A2(n12319), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11855) );
  OAI211_X1 U14254 ( .C1(n12294), .C2(n11977), .A(n11856), .B(n11855), .ZN(
        n11857) );
  AOI21_X1 U14255 ( .B1(n12298), .B2(n11979), .A(n11857), .ZN(n11858) );
  OAI21_X1 U14256 ( .B1(n11859), .B2(n11981), .A(n11858), .ZN(P3_U3163) );
  XNOR2_X1 U14257 ( .A(n11861), .B(n11860), .ZN(n11944) );
  NOR2_X1 U14258 ( .A1(n11944), .A2(n11945), .ZN(n11943) );
  AOI21_X1 U14259 ( .B1(n11861), .B2(n11860), .A(n11943), .ZN(n11864) );
  XNOR2_X1 U14260 ( .A(n11862), .B(n11990), .ZN(n11863) );
  XNOR2_X1 U14261 ( .A(n11864), .B(n11863), .ZN(n11872) );
  AND2_X1 U14262 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n12005) );
  NOR2_X1 U14263 ( .A1(n11977), .A2(n12384), .ZN(n11865) );
  AOI211_X1 U14264 ( .C1(n11974), .C2(n11866), .A(n12005), .B(n11865), .ZN(
        n11867) );
  OAI21_X1 U14265 ( .B1(n11868), .B2(n11968), .A(n11867), .ZN(n11869) );
  AOI21_X1 U14266 ( .B1(n11870), .B2(n11972), .A(n11869), .ZN(n11871) );
  OAI21_X1 U14267 ( .B1(n11872), .B2(n11981), .A(n11871), .ZN(P3_U3164) );
  INV_X1 U14268 ( .A(n11873), .ZN(n11875) );
  NOR3_X1 U14269 ( .A1(n6463), .A2(n11875), .A3(n11874), .ZN(n11878) );
  INV_X1 U14270 ( .A(n11876), .ZN(n11877) );
  OAI21_X1 U14271 ( .B1(n11878), .B2(n11877), .A(n11963), .ZN(n11882) );
  NOR2_X1 U14272 ( .A1(n12266), .A2(n11916), .ZN(n11880) );
  OAI22_X1 U14273 ( .A1(n12215), .A2(n11977), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15102), .ZN(n11879) );
  AOI211_X1 U14274 ( .C1(n12241), .C2(n11972), .A(n11880), .B(n11879), .ZN(
        n11881) );
  OAI211_X1 U14275 ( .C1(n11883), .C2(n11968), .A(n11882), .B(n11881), .ZN(
        P3_U3165) );
  XNOR2_X1 U14276 ( .A(n11884), .B(n12345), .ZN(n11885) );
  XNOR2_X1 U14277 ( .A(n11886), .B(n11885), .ZN(n11891) );
  NAND2_X1 U14278 ( .A1(n11972), .A2(n12362), .ZN(n11888) );
  AND2_X1 U14279 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12118) );
  AOI21_X1 U14280 ( .B1(n11913), .B2(n11952), .A(n12118), .ZN(n11887) );
  OAI211_X1 U14281 ( .C1(n12385), .C2(n11916), .A(n11888), .B(n11887), .ZN(
        n11889) );
  AOI21_X1 U14282 ( .B1(n12361), .B2(n11979), .A(n11889), .ZN(n11890) );
  OAI21_X1 U14283 ( .B1(n11891), .B2(n11981), .A(n11890), .ZN(P3_U3166) );
  XNOR2_X1 U14284 ( .A(n11893), .B(n11892), .ZN(n11898) );
  NAND2_X1 U14285 ( .A1(n11972), .A2(n12350), .ZN(n11895) );
  AND2_X1 U14286 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14154) );
  AOI21_X1 U14287 ( .B1(n11913), .B2(n12344), .A(n14154), .ZN(n11894) );
  OAI211_X1 U14288 ( .C1(n12368), .C2(n11916), .A(n11895), .B(n11894), .ZN(
        n11896) );
  AOI21_X1 U14289 ( .B1(n12444), .B2(n11979), .A(n11896), .ZN(n11897) );
  OAI21_X1 U14290 ( .B1(n11898), .B2(n11981), .A(n11897), .ZN(P3_U3168) );
  INV_X1 U14291 ( .A(n11899), .ZN(n11901) );
  NOR3_X1 U14292 ( .A1(n11902), .A2(n11901), .A3(n11900), .ZN(n11903) );
  OAI21_X1 U14293 ( .B1(n11903), .B2(n6463), .A(n11963), .ZN(n11908) );
  NOR2_X1 U14294 ( .A1(n12282), .A2(n11916), .ZN(n11906) );
  OAI22_X1 U14295 ( .A1(n12249), .A2(n11977), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11904), .ZN(n11905) );
  AOI211_X1 U14296 ( .C1(n12255), .C2(n11972), .A(n11906), .B(n11905), .ZN(
        n11907) );
  OAI211_X1 U14297 ( .C1(n6591), .C2(n11968), .A(n11908), .B(n11907), .ZN(
        P3_U3169) );
  NAND2_X1 U14298 ( .A1(n11910), .A2(n11909), .ZN(n11912) );
  XNOR2_X1 U14299 ( .A(n11912), .B(n11911), .ZN(n11919) );
  AOI22_X1 U14300 ( .A1(n11913), .A2(n12306), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11915) );
  NAND2_X1 U14301 ( .A1(n11972), .A2(n12312), .ZN(n11914) );
  OAI211_X1 U14302 ( .C1(n12332), .C2(n11916), .A(n11915), .B(n11914), .ZN(
        n11917) );
  AOI21_X1 U14303 ( .B1(n12432), .B2(n11979), .A(n11917), .ZN(n11918) );
  OAI21_X1 U14304 ( .B1(n11919), .B2(n11981), .A(n11918), .ZN(P3_U3173) );
  XNOR2_X1 U14305 ( .A(n11921), .B(n11920), .ZN(n11922) );
  XNOR2_X1 U14306 ( .A(n11923), .B(n11922), .ZN(n11930) );
  NAND2_X1 U14307 ( .A1(n11972), .A2(n11924), .ZN(n11927) );
  NOR2_X1 U14308 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11925), .ZN(n12041) );
  AOI21_X1 U14309 ( .B1(n11974), .B2(n11990), .A(n12041), .ZN(n11926) );
  OAI211_X1 U14310 ( .C1(n12369), .C2(n11977), .A(n11927), .B(n11926), .ZN(
        n11928) );
  AOI21_X1 U14311 ( .B1(n14162), .B2(n11979), .A(n11928), .ZN(n11929) );
  OAI21_X1 U14312 ( .B1(n11930), .B2(n11981), .A(n11929), .ZN(P3_U3174) );
  AOI21_X1 U14313 ( .B1(n11987), .B2(n11931), .A(n6467), .ZN(n11936) );
  NAND2_X1 U14314 ( .A1(n11972), .A2(n12287), .ZN(n11933) );
  AOI22_X1 U14315 ( .A1(n11940), .A2(n12306), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11932) );
  OAI211_X1 U14316 ( .C1(n12282), .C2(n11977), .A(n11933), .B(n11932), .ZN(
        n11934) );
  AOI21_X1 U14317 ( .B1(n12286), .B2(n11979), .A(n11934), .ZN(n11935) );
  OAI21_X1 U14318 ( .B1(n11936), .B2(n11981), .A(n11935), .ZN(P3_U3175) );
  NOR2_X1 U14319 ( .A1(n11977), .A2(n11937), .ZN(n11938) );
  AOI211_X1 U14320 ( .C1(n11940), .C2(n11991), .A(n11939), .B(n11938), .ZN(
        n11941) );
  OAI21_X1 U14321 ( .B1(n11968), .B2(n11942), .A(n11941), .ZN(n11947) );
  AOI211_X1 U14322 ( .C1(n11945), .C2(n11944), .A(n11981), .B(n11943), .ZN(
        n11946) );
  AOI211_X1 U14323 ( .C1(n11948), .C2(n11972), .A(n11947), .B(n11946), .ZN(
        n11949) );
  INV_X1 U14324 ( .A(n11949), .ZN(P3_U3176) );
  XNOR2_X1 U14325 ( .A(n11950), .B(n11951), .ZN(n11958) );
  NAND2_X1 U14326 ( .A1(n11974), .A2(n11952), .ZN(n11953) );
  NAND2_X1 U14327 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12134)
         );
  OAI211_X1 U14328 ( .C1(n11977), .C2(n12332), .A(n11953), .B(n12134), .ZN(
        n11956) );
  INV_X1 U14329 ( .A(n11954), .ZN(n12500) );
  NOR2_X1 U14330 ( .A1(n12500), .A2(n11968), .ZN(n11955) );
  AOI211_X1 U14331 ( .C1(n12338), .C2(n11972), .A(n11956), .B(n11955), .ZN(
        n11957) );
  OAI21_X1 U14332 ( .B1(n11958), .B2(n11981), .A(n11957), .ZN(P3_U3178) );
  INV_X1 U14333 ( .A(n11959), .ZN(n12479) );
  OAI21_X1 U14334 ( .B1(n11962), .B2(n11961), .A(n11960), .ZN(n11964) );
  AOI22_X1 U14335 ( .A1(n11986), .A2(n11974), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11965) );
  OAI21_X1 U14336 ( .B1(n12226), .B2(n11977), .A(n11965), .ZN(n11966) );
  AOI21_X1 U14337 ( .B1(n12229), .B2(n11972), .A(n11966), .ZN(n11967) );
  XNOR2_X1 U14338 ( .A(n11970), .B(n11988), .ZN(n11971) );
  XNOR2_X1 U14339 ( .A(n11969), .B(n11971), .ZN(n11982) );
  NAND2_X1 U14340 ( .A1(n11972), .A2(n12376), .ZN(n11976) );
  NOR2_X1 U14341 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11973), .ZN(n12093) );
  AOI21_X1 U14342 ( .B1(n11974), .B2(n11989), .A(n12093), .ZN(n11975) );
  OAI211_X1 U14343 ( .C1(n12368), .C2(n11977), .A(n11976), .B(n11975), .ZN(
        n11978) );
  AOI21_X1 U14344 ( .B1(n12452), .B2(n11979), .A(n11978), .ZN(n11980) );
  OAI21_X1 U14345 ( .B1(n11982), .B2(n11981), .A(n11980), .ZN(P3_U3181) );
  MUX2_X1 U14346 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12183), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14347 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n11983), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14348 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n11984), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14349 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n11985), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14350 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12201), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14351 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12236), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14352 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n11986), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14353 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n6590), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14354 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n11987), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14355 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12306), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14356 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12319), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14357 ( .A(n12305), .B(P3_DATAO_REG_19__SCAN_IN), .S(n11997), .Z(
        P3_U3510) );
  MUX2_X1 U14358 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12344), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14359 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12345), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14360 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n11988), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14361 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n11989), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14362 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n11990), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14363 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n11991), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14364 ( .A(n14887), .B(P3_DATAO_REG_9__SCAN_IN), .S(n11997), .Z(
        P3_U3500) );
  MUX2_X1 U14365 ( .A(n11992), .B(P3_DATAO_REG_8__SCAN_IN), .S(n11997), .Z(
        P3_U3499) );
  MUX2_X1 U14366 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n14888), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14367 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n11993), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14368 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n11994), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14369 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n11995), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14370 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n14921), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14371 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n11996), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14372 ( .A(n14918), .B(P3_DATAO_REG_0__SCAN_IN), .S(n11997), .Z(
        P3_U3491) );
  NOR2_X1 U14373 ( .A1(n11998), .A2(n12018), .ZN(n12000) );
  MUX2_X1 U14374 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n14738), .Z(n12037) );
  XNOR2_X1 U14375 ( .A(n12037), .B(n12036), .ZN(n11999) );
  NOR3_X1 U14376 ( .A1(n12001), .A2(n12000), .A3(n11999), .ZN(n12035) );
  INV_X1 U14377 ( .A(n12035), .ZN(n12003) );
  OAI21_X1 U14378 ( .B1(n12001), .B2(n12000), .A(n11999), .ZN(n12002) );
  NAND3_X1 U14379 ( .A1(n12003), .A2(n14863), .A3(n12002), .ZN(n12028) );
  INV_X1 U14380 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n13999) );
  NOR2_X1 U14381 ( .A1(n14837), .A2(n13999), .ZN(n12004) );
  AOI211_X1 U14382 ( .C1(n14828), .C2(n12033), .A(n12005), .B(n12004), .ZN(
        n12027) );
  NOR2_X1 U14383 ( .A1(n12007), .A2(n12006), .ZN(n12009) );
  INV_X1 U14384 ( .A(n12012), .ZN(n12014) );
  MUX2_X1 U14385 ( .A(n12010), .B(P3_REG2_REG_12__SCAN_IN), .S(n12036), .Z(
        n12011) );
  INV_X1 U14386 ( .A(n12011), .ZN(n12013) );
  OR2_X2 U14387 ( .A1(n12012), .A2(n12011), .ZN(n12030) );
  OAI21_X1 U14388 ( .B1(n12014), .B2(n12013), .A(n12030), .ZN(n12016) );
  INV_X1 U14389 ( .A(n14878), .ZN(n12015) );
  NAND2_X1 U14390 ( .A1(n12016), .A2(n12015), .ZN(n12026) );
  NAND2_X1 U14391 ( .A1(n12018), .A2(n12017), .ZN(n12020) );
  NAND2_X1 U14392 ( .A1(n12020), .A2(n12019), .ZN(n12023) );
  INV_X1 U14393 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12021) );
  MUX2_X1 U14394 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n12021), .S(n12036), .Z(
        n12022) );
  NAND2_X1 U14395 ( .A1(n12023), .A2(n12022), .ZN(n12032) );
  OAI21_X1 U14396 ( .B1(n12023), .B2(n12022), .A(n12032), .ZN(n12024) );
  NAND2_X1 U14397 ( .A1(n12024), .A2(n14874), .ZN(n12025) );
  NAND4_X1 U14398 ( .A1(n12028), .A2(n12027), .A3(n12026), .A4(n12025), .ZN(
        P3_U3194) );
  NAND2_X1 U14399 ( .A1(n12036), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12029) );
  AOI21_X1 U14400 ( .B1(n8579), .B2(n12031), .A(n12049), .ZN(n12047) );
  OAI21_X1 U14401 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n12034), .A(n12056), 
        .ZN(n12045) );
  AOI21_X1 U14402 ( .B1(n12037), .B2(n12036), .A(n12035), .ZN(n12039) );
  MUX2_X1 U14403 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n14738), .Z(n12060) );
  XNOR2_X1 U14404 ( .A(n12060), .B(n12061), .ZN(n12038) );
  NAND2_X1 U14405 ( .A1(n12039), .A2(n12038), .ZN(n12068) );
  OAI21_X1 U14406 ( .B1(n12039), .B2(n12038), .A(n12068), .ZN(n12040) );
  NAND2_X1 U14407 ( .A1(n12040), .A2(n14863), .ZN(n12043) );
  AOI21_X1 U14408 ( .B1(n14871), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n12041), 
        .ZN(n12042) );
  OAI211_X1 U14409 ( .C1(n14868), .C2(n12055), .A(n12043), .B(n12042), .ZN(
        n12044) );
  AOI21_X1 U14410 ( .B1(n14874), .B2(n12045), .A(n12044), .ZN(n12046) );
  OAI21_X1 U14411 ( .B1(n12047), .B2(n14878), .A(n12046), .ZN(P3_U3195) );
  NOR2_X1 U14412 ( .A1(n12061), .A2(n12048), .ZN(n12050) );
  OR2_X1 U14413 ( .A1(n12071), .A2(n12051), .ZN(n12084) );
  NAND2_X1 U14414 ( .A1(n12071), .A2(n12051), .ZN(n12052) );
  NAND2_X1 U14415 ( .A1(n12084), .A2(n12052), .ZN(n12063) );
  NOR2_X2 U14416 ( .A1(n12053), .A2(n12063), .ZN(n12079) );
  AOI21_X1 U14417 ( .B1(n12053), .B2(n12063), .A(n12079), .ZN(n12078) );
  NAND2_X1 U14418 ( .A1(n12055), .A2(n12054), .ZN(n12057) );
  INV_X1 U14419 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n15020) );
  OR2_X1 U14420 ( .A1(n12071), .A2(n15020), .ZN(n12083) );
  NAND2_X1 U14421 ( .A1(n12071), .A2(n15020), .ZN(n12058) );
  AND2_X1 U14422 ( .A1(n12083), .A2(n12058), .ZN(n12064) );
  NAND2_X1 U14423 ( .A1(n12064), .A2(n12059), .ZN(n12081) );
  OAI21_X1 U14424 ( .B1(n12059), .B2(n12064), .A(n12081), .ZN(n12076) );
  INV_X1 U14425 ( .A(n12060), .ZN(n12062) );
  NAND2_X1 U14426 ( .A1(n12062), .A2(n12061), .ZN(n12067) );
  INV_X1 U14427 ( .A(n12063), .ZN(n12065) );
  MUX2_X1 U14428 ( .A(n12065), .B(n12064), .S(n14738), .Z(n12066) );
  NAND3_X1 U14429 ( .A1(n12068), .A2(n12067), .A3(n12066), .ZN(n12086) );
  NAND2_X1 U14430 ( .A1(n12086), .A2(n14863), .ZN(n12074) );
  AOI21_X1 U14431 ( .B1(n12068), .B2(n12067), .A(n12066), .ZN(n12073) );
  INV_X1 U14432 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n13998) );
  NOR2_X1 U14433 ( .A1(n14837), .A2(n13998), .ZN(n12069) );
  AOI211_X1 U14434 ( .C1(n14828), .C2(n12071), .A(n12070), .B(n12069), .ZN(
        n12072) );
  OAI21_X1 U14435 ( .B1(n12074), .B2(n12073), .A(n12072), .ZN(n12075) );
  AOI21_X1 U14436 ( .B1(n14874), .B2(n12076), .A(n12075), .ZN(n12077) );
  OAI21_X1 U14437 ( .B1(n12078), .B2(n14878), .A(n12077), .ZN(P3_U3196) );
  AOI21_X1 U14438 ( .B1(n12089), .B2(n12080), .A(n12103), .ZN(n12099) );
  OAI21_X1 U14439 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12082), .A(n12109), 
        .ZN(n12097) );
  MUX2_X1 U14440 ( .A(n12084), .B(n12083), .S(n14738), .Z(n12085) );
  NAND2_X1 U14441 ( .A1(n12086), .A2(n12085), .ZN(n12113) );
  XNOR2_X1 U14442 ( .A(n12113), .B(n12087), .ZN(n12091) );
  INV_X1 U14443 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12088) );
  MUX2_X1 U14444 ( .A(n12089), .B(n12088), .S(n14738), .Z(n12090) );
  NAND2_X1 U14445 ( .A1(n12091), .A2(n12090), .ZN(n12111) );
  OAI21_X1 U14446 ( .B1(n12091), .B2(n12090), .A(n12111), .ZN(n12092) );
  NAND2_X1 U14447 ( .A1(n12092), .A2(n14863), .ZN(n12095) );
  AOI21_X1 U14448 ( .B1(n14871), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n12093), 
        .ZN(n12094) );
  OAI211_X1 U14449 ( .C1(n14868), .C2(n12112), .A(n12095), .B(n12094), .ZN(
        n12096) );
  AOI21_X1 U14450 ( .B1(n14874), .B2(n12097), .A(n12096), .ZN(n12098) );
  OAI21_X1 U14451 ( .B1(n12099), .B2(n14878), .A(n12098), .ZN(P3_U3197) );
  OR2_X1 U14452 ( .A1(n12126), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12101) );
  NAND2_X1 U14453 ( .A1(n12126), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n12100) );
  AND2_X1 U14454 ( .A1(n12101), .A2(n12100), .ZN(n12107) );
  AND2_X1 U14455 ( .A1(n12112), .A2(n12102), .ZN(n12104) );
  OR2_X2 U14456 ( .A1(n12106), .A2(n12107), .ZN(n12128) );
  INV_X1 U14457 ( .A(n12128), .ZN(n12105) );
  AOI21_X1 U14458 ( .B1(n12107), .B2(n12106), .A(n12105), .ZN(n12124) );
  NAND2_X1 U14459 ( .A1(n12112), .A2(n12108), .ZN(n12110) );
  XNOR2_X1 U14460 ( .A(n12126), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n12137) );
  XNOR2_X1 U14461 ( .A(n12138), .B(n12137), .ZN(n12122) );
  OAI21_X1 U14462 ( .B1(n12113), .B2(n12112), .A(n12111), .ZN(n12148) );
  MUX2_X1 U14463 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n14738), .Z(n12114) );
  NOR2_X1 U14464 ( .A1(n12114), .A2(n12136), .ZN(n12146) );
  INV_X1 U14465 ( .A(n12146), .ZN(n12115) );
  NAND2_X1 U14466 ( .A1(n12114), .A2(n12136), .ZN(n12147) );
  NAND2_X1 U14467 ( .A1(n12115), .A2(n12147), .ZN(n12116) );
  XNOR2_X1 U14468 ( .A(n12148), .B(n12116), .ZN(n12120) );
  INV_X1 U14469 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14089) );
  NOR2_X1 U14470 ( .A1(n14837), .A2(n14089), .ZN(n12117) );
  AOI211_X1 U14471 ( .C1(n14828), .C2(n12126), .A(n12118), .B(n12117), .ZN(
        n12119) );
  OAI21_X1 U14472 ( .B1(n12120), .B2(n14761), .A(n12119), .ZN(n12121) );
  AOI21_X1 U14473 ( .B1(n14874), .B2(n12122), .A(n12121), .ZN(n12123) );
  OAI21_X1 U14474 ( .B1(n12124), .B2(n14878), .A(n12123), .ZN(P3_U3198) );
  OR2_X1 U14475 ( .A1(n12126), .A2(n12125), .ZN(n12127) );
  OR2_X1 U14476 ( .A1(n12165), .A2(n12130), .ZN(n12158) );
  NAND2_X1 U14477 ( .A1(n12165), .A2(n12130), .ZN(n12131) );
  NAND2_X1 U14478 ( .A1(n12158), .A2(n12131), .ZN(n12132) );
  AOI21_X1 U14479 ( .B1(n12133), .B2(n12132), .A(n12160), .ZN(n12157) );
  INV_X1 U14480 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12135) );
  OAI21_X1 U14481 ( .B1(n14837), .B2(n12135), .A(n12134), .ZN(n12145) );
  AOI22_X1 U14482 ( .A1(n12138), .A2(n12137), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n12136), .ZN(n12139) );
  OR2_X1 U14483 ( .A1(n12139), .A2(n12151), .ZN(n12141) );
  XNOR2_X1 U14484 ( .A(n12139), .B(n14157), .ZN(n14150) );
  NAND2_X1 U14485 ( .A1(P3_REG1_REG_17__SCAN_IN), .A2(n14150), .ZN(n14149) );
  INV_X1 U14486 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12442) );
  XNOR2_X1 U14487 ( .A(n12165), .B(n12442), .ZN(n12140) );
  AOI21_X1 U14488 ( .B1(n12141), .B2(n14149), .A(n12140), .ZN(n12172) );
  INV_X1 U14489 ( .A(n12172), .ZN(n12143) );
  NAND3_X1 U14490 ( .A1(n12141), .A2(n14149), .A3(n12140), .ZN(n12142) );
  AOI21_X1 U14491 ( .B1(n12143), .B2(n12142), .A(n14741), .ZN(n12144) );
  AOI211_X1 U14492 ( .C1(n14828), .C2(n12165), .A(n12145), .B(n12144), .ZN(
        n12156) );
  MUX2_X1 U14493 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n14738), .Z(n12149) );
  INV_X1 U14494 ( .A(n12149), .ZN(n12150) );
  AOI21_X1 U14495 ( .B1(n12148), .B2(n12147), .A(n12146), .ZN(n14153) );
  XNOR2_X1 U14496 ( .A(n12149), .B(n12151), .ZN(n14152) );
  NAND2_X1 U14497 ( .A1(n14153), .A2(n14152), .ZN(n14151) );
  MUX2_X1 U14498 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n14738), .Z(n12152) );
  NOR2_X1 U14499 ( .A1(n12153), .A2(n12152), .ZN(n12164) );
  AND2_X1 U14500 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  OAI21_X1 U14501 ( .B1(n12164), .B2(n12154), .A(n14863), .ZN(n12155) );
  OAI211_X1 U14502 ( .C1(n12157), .C2(n14878), .A(n12156), .B(n12155), .ZN(
        P3_U3200) );
  INV_X1 U14503 ( .A(n12158), .ZN(n12159) );
  NOR2_X1 U14504 ( .A1(n12160), .A2(n12159), .ZN(n12162) );
  XNOR2_X1 U14505 ( .A(n12177), .B(n12161), .ZN(n12167) );
  XNOR2_X1 U14506 ( .A(n12162), .B(n12167), .ZN(n12180) );
  INV_X1 U14507 ( .A(n12163), .ZN(n12166) );
  AOI21_X1 U14508 ( .B1(n12166), .B2(n12165), .A(n12164), .ZN(n12171) );
  XNOR2_X1 U14509 ( .A(n12177), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12174) );
  INV_X1 U14510 ( .A(n12167), .ZN(n12169) );
  MUX2_X1 U14511 ( .A(n12174), .B(n12169), .S(n12168), .Z(n12170) );
  XNOR2_X1 U14512 ( .A(n12171), .B(n12170), .ZN(n12179) );
  AOI21_X1 U14513 ( .B1(P3_REG1_REG_18__SCAN_IN), .B2(n6811), .A(n12172), .ZN(
        n12173) );
  NAND2_X1 U14514 ( .A1(n14871), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12175) );
  OAI211_X1 U14515 ( .C1(n14868), .C2(n12177), .A(n12176), .B(n12175), .ZN(
        n12178) );
  NAND2_X1 U14516 ( .A1(n12181), .A2(n12275), .ZN(n12186) );
  NAND2_X1 U14517 ( .A1(n12183), .A2(n12182), .ZN(n12460) );
  INV_X1 U14518 ( .A(n12460), .ZN(n12185) );
  NOR2_X1 U14519 ( .A1(n12184), .A2(n12271), .ZN(n12191) );
  AOI21_X1 U14520 ( .B1(n12185), .B2(n14933), .A(n12191), .ZN(n12189) );
  OAI211_X1 U14521 ( .C1(n14933), .C2(n12187), .A(n12186), .B(n12189), .ZN(
        P3_U3202) );
  NAND2_X1 U14522 ( .A1(n14935), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12188) );
  OAI211_X1 U14523 ( .C1(n12190), .C2(n12391), .A(n12189), .B(n12188), .ZN(
        P3_U3203) );
  AOI21_X1 U14524 ( .B1(n14935), .B2(P3_REG2_REG_29__SCAN_IN), .A(n12191), 
        .ZN(n12192) );
  OAI21_X1 U14525 ( .B1(n12193), .B2(n12391), .A(n12192), .ZN(n12194) );
  AOI21_X1 U14526 ( .B1(n12195), .B2(n12393), .A(n12194), .ZN(n12196) );
  OAI21_X1 U14527 ( .B1(n12197), .B2(n14935), .A(n12196), .ZN(P3_U3204) );
  OAI211_X1 U14528 ( .C1(n12200), .C2(n12199), .A(n12198), .B(n14923), .ZN(
        n12203) );
  NAND2_X1 U14529 ( .A1(n12201), .A2(n14919), .ZN(n12202) );
  OAI211_X1 U14530 ( .C1(n12204), .C2(n14901), .A(n12203), .B(n12202), .ZN(
        n12400) );
  INV_X1 U14531 ( .A(n12400), .ZN(n12211) );
  OAI21_X1 U14532 ( .B1(n12206), .B2(n7384), .A(n12205), .ZN(n12401) );
  AOI22_X1 U14533 ( .A1(n12207), .A2(n14929), .B1(P3_REG2_REG_28__SCAN_IN), 
        .B2(n14935), .ZN(n12208) );
  OAI21_X1 U14534 ( .B1(n12471), .B2(n12391), .A(n12208), .ZN(n12209) );
  AOI21_X1 U14535 ( .B1(n12401), .B2(n12393), .A(n12209), .ZN(n12210) );
  OAI21_X1 U14536 ( .B1(n12211), .B2(n14935), .A(n12210), .ZN(P3_U3205) );
  XNOR2_X1 U14537 ( .A(n12212), .B(n12217), .ZN(n12213) );
  OAI222_X1 U14538 ( .A1(n14903), .A2(n12215), .B1(n14901), .B2(n12214), .C1(
        n12213), .C2(n14891), .ZN(n12404) );
  INV_X1 U14539 ( .A(n12404), .ZN(n12223) );
  OAI21_X1 U14540 ( .B1(n12218), .B2(n12217), .A(n12216), .ZN(n12405) );
  AOI22_X1 U14541 ( .A1(n12219), .A2(n14929), .B1(n14935), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12220) );
  OAI21_X1 U14542 ( .B1(n12475), .B2(n12391), .A(n12220), .ZN(n12221) );
  AOI21_X1 U14543 ( .B1(n12405), .B2(n12393), .A(n12221), .ZN(n12222) );
  OAI21_X1 U14544 ( .B1(n12223), .B2(n14935), .A(n12222), .ZN(P3_U3206) );
  XNOR2_X1 U14545 ( .A(n12224), .B(n12227), .ZN(n12225) );
  OAI222_X1 U14546 ( .A1(n14903), .A2(n12249), .B1(n14901), .B2(n12226), .C1(
        n12225), .C2(n14891), .ZN(n12408) );
  INV_X1 U14547 ( .A(n12408), .ZN(n12233) );
  XNOR2_X1 U14548 ( .A(n12228), .B(n12227), .ZN(n12409) );
  AOI22_X1 U14549 ( .A1(n12229), .A2(n14929), .B1(n14935), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12230) );
  OAI21_X1 U14550 ( .B1(n12479), .B2(n12391), .A(n12230), .ZN(n12231) );
  AOI21_X1 U14551 ( .B1(n12409), .B2(n12393), .A(n12231), .ZN(n12232) );
  OAI21_X1 U14552 ( .B1(n12233), .B2(n14935), .A(n12232), .ZN(P3_U3207) );
  OAI211_X1 U14553 ( .C1(n12235), .C2(n12239), .A(n12234), .B(n14923), .ZN(
        n12238) );
  NAND2_X1 U14554 ( .A1(n12236), .A2(n14920), .ZN(n12237) );
  OAI211_X1 U14555 ( .C1(n12266), .C2(n14903), .A(n12238), .B(n12237), .ZN(
        n12412) );
  XNOR2_X1 U14556 ( .A(n12240), .B(n12239), .ZN(n12415) );
  AOI22_X1 U14557 ( .A1(n14935), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n12241), 
        .B2(n14929), .ZN(n12243) );
  NAND2_X1 U14558 ( .A1(n12413), .A2(n12275), .ZN(n12242) );
  OAI211_X1 U14559 ( .C1(n12415), .C2(n12327), .A(n12243), .B(n12242), .ZN(
        n12244) );
  AOI21_X1 U14560 ( .B1(n12412), .B2(n14933), .A(n12244), .ZN(n12245) );
  INV_X1 U14561 ( .A(n12245), .ZN(P3_U3208) );
  AOI21_X1 U14562 ( .B1(n12247), .B2(n12246), .A(n6517), .ZN(n12248) );
  OAI222_X1 U14563 ( .A1(n14901), .A2(n12249), .B1(n14903), .B2(n12282), .C1(
        n14891), .C2(n12248), .ZN(n12416) );
  INV_X1 U14564 ( .A(n12416), .ZN(n12259) );
  INV_X1 U14565 ( .A(n12262), .ZN(n12252) );
  OAI21_X1 U14566 ( .B1(n12252), .B2(n12251), .A(n12250), .ZN(n12254) );
  NAND2_X1 U14567 ( .A1(n12254), .A2(n12253), .ZN(n12417) );
  AOI22_X1 U14568 ( .A1(n14935), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n14929), 
        .B2(n12255), .ZN(n12256) );
  OAI21_X1 U14569 ( .B1(n6591), .B2(n12391), .A(n12256), .ZN(n12257) );
  AOI21_X1 U14570 ( .B1(n12417), .B2(n12393), .A(n12257), .ZN(n12258) );
  OAI21_X1 U14571 ( .B1(n12259), .B2(n14935), .A(n12258), .ZN(P3_U3209) );
  NAND2_X1 U14572 ( .A1(n12260), .A2(n12263), .ZN(n12261) );
  NAND2_X1 U14573 ( .A1(n12262), .A2(n12261), .ZN(n12422) );
  XNOR2_X1 U14574 ( .A(n12264), .B(n12263), .ZN(n12265) );
  NAND2_X1 U14575 ( .A1(n12265), .A2(n14923), .ZN(n12269) );
  OAI22_X1 U14576 ( .A1(n12266), .A2(n14901), .B1(n12294), .B2(n14903), .ZN(
        n12267) );
  INV_X1 U14577 ( .A(n12267), .ZN(n12268) );
  NAND2_X1 U14578 ( .A1(n12269), .A2(n12268), .ZN(n12424) );
  NAND2_X1 U14579 ( .A1(n12424), .A2(n14933), .ZN(n12278) );
  INV_X1 U14580 ( .A(n12270), .ZN(n12272) );
  OAI22_X1 U14581 ( .A1(n14933), .A2(n12273), .B1(n12272), .B2(n12271), .ZN(
        n12274) );
  AOI21_X1 U14582 ( .B1(n12276), .B2(n12275), .A(n12274), .ZN(n12277) );
  OAI211_X1 U14583 ( .C1(n12327), .C2(n12422), .A(n12278), .B(n12277), .ZN(
        P3_U3210) );
  XNOR2_X1 U14584 ( .A(n12280), .B(n12279), .ZN(n12281) );
  OAI222_X1 U14585 ( .A1(n14903), .A2(n12283), .B1(n14901), .B2(n12282), .C1(
        n14891), .C2(n12281), .ZN(n12425) );
  INV_X1 U14586 ( .A(n12425), .ZN(n12291) );
  XNOR2_X1 U14587 ( .A(n12285), .B(n12284), .ZN(n12426) );
  INV_X1 U14588 ( .A(n12286), .ZN(n12487) );
  AOI22_X1 U14589 ( .A1(n14935), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n14929), 
        .B2(n12287), .ZN(n12288) );
  OAI21_X1 U14590 ( .B1(n12487), .B2(n12391), .A(n12288), .ZN(n12289) );
  AOI21_X1 U14591 ( .B1(n12426), .B2(n12393), .A(n12289), .ZN(n12290) );
  OAI21_X1 U14592 ( .B1(n12291), .B2(n14935), .A(n12290), .ZN(P3_U3211) );
  XNOR2_X1 U14593 ( .A(n12292), .B(n12296), .ZN(n12293) );
  OAI222_X1 U14594 ( .A1(n14903), .A2(n12295), .B1(n14901), .B2(n12294), .C1(
        n12293), .C2(n14891), .ZN(n12428) );
  INV_X1 U14595 ( .A(n12428), .ZN(n12303) );
  XNOR2_X1 U14596 ( .A(n12297), .B(n12296), .ZN(n12429) );
  INV_X1 U14597 ( .A(n12298), .ZN(n12491) );
  AOI22_X1 U14598 ( .A1(n14935), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n14929), 
        .B2(n12299), .ZN(n12300) );
  OAI21_X1 U14599 ( .B1(n12491), .B2(n12391), .A(n12300), .ZN(n12301) );
  AOI21_X1 U14600 ( .B1(n12429), .B2(n12393), .A(n12301), .ZN(n12302) );
  OAI21_X1 U14601 ( .B1(n12303), .B2(n14935), .A(n12302), .ZN(P3_U3212) );
  XOR2_X1 U14602 ( .A(n12304), .B(n12311), .Z(n12307) );
  AOI222_X1 U14603 ( .A1(n14923), .A2(n12307), .B1(n12306), .B2(n14920), .C1(
        n12305), .C2(n14919), .ZN(n12435) );
  INV_X1 U14604 ( .A(n12308), .ZN(n12309) );
  AOI21_X1 U14605 ( .B1(n12311), .B2(n12310), .A(n12309), .ZN(n12433) );
  INV_X1 U14606 ( .A(n12432), .ZN(n12314) );
  AOI22_X1 U14607 ( .A1(n14935), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n14929), 
        .B2(n12312), .ZN(n12313) );
  OAI21_X1 U14608 ( .B1(n12314), .B2(n12391), .A(n12313), .ZN(n12315) );
  AOI21_X1 U14609 ( .B1(n12433), .B2(n12393), .A(n12315), .ZN(n12316) );
  OAI21_X1 U14610 ( .B1(n12435), .B2(n14935), .A(n12316), .ZN(P3_U3213) );
  XNOR2_X1 U14611 ( .A(n12317), .B(n7564), .ZN(n12437) );
  INV_X1 U14612 ( .A(n12437), .ZN(n12326) );
  OAI211_X1 U14613 ( .C1(n6575), .C2(n7564), .A(n14923), .B(n12318), .ZN(
        n12321) );
  AOI22_X1 U14614 ( .A1(n12319), .A2(n14920), .B1(n12344), .B2(n14919), .ZN(
        n12320) );
  NAND2_X1 U14615 ( .A1(n12321), .A2(n12320), .ZN(n12436) );
  AOI22_X1 U14616 ( .A1(n14935), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n14929), 
        .B2(n12322), .ZN(n12323) );
  OAI21_X1 U14617 ( .B1(n12496), .B2(n12391), .A(n12323), .ZN(n12324) );
  AOI21_X1 U14618 ( .B1(n12436), .B2(n14933), .A(n12324), .ZN(n12325) );
  OAI21_X1 U14619 ( .B1(n12327), .B2(n12326), .A(n12325), .ZN(P3_U3214) );
  INV_X1 U14620 ( .A(n12328), .ZN(n12329) );
  AOI21_X1 U14621 ( .B1(n12334), .B2(n12330), .A(n12329), .ZN(n12331) );
  OAI222_X1 U14622 ( .A1(n14903), .A2(n12358), .B1(n14901), .B2(n12332), .C1(
        n14891), .C2(n12331), .ZN(n12440) );
  INV_X1 U14623 ( .A(n12440), .ZN(n12342) );
  INV_X1 U14624 ( .A(n12333), .ZN(n12337) );
  AOI21_X1 U14625 ( .B1(n12347), .B2(n12335), .A(n12334), .ZN(n12336) );
  NOR2_X1 U14626 ( .A1(n12337), .A2(n12336), .ZN(n12441) );
  AOI22_X1 U14627 ( .A1(n14935), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n14929), 
        .B2(n12338), .ZN(n12339) );
  OAI21_X1 U14628 ( .B1(n12500), .B2(n12391), .A(n12339), .ZN(n12340) );
  AOI21_X1 U14629 ( .B1(n12441), .B2(n12393), .A(n12340), .ZN(n12341) );
  OAI21_X1 U14630 ( .B1(n12342), .B2(n14935), .A(n12341), .ZN(P3_U3215) );
  XNOR2_X1 U14631 ( .A(n12343), .B(n12348), .ZN(n12346) );
  AOI222_X1 U14632 ( .A1(n14923), .A2(n12346), .B1(n12345), .B2(n14919), .C1(
        n12344), .C2(n14920), .ZN(n12447) );
  OAI21_X1 U14633 ( .B1(n12349), .B2(n12348), .A(n12347), .ZN(n12445) );
  INV_X1 U14634 ( .A(n12444), .ZN(n12352) );
  AOI22_X1 U14635 ( .A1(n14935), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n14929), 
        .B2(n12350), .ZN(n12351) );
  OAI21_X1 U14636 ( .B1(n12352), .B2(n12391), .A(n12351), .ZN(n12353) );
  AOI21_X1 U14637 ( .B1(n12445), .B2(n12393), .A(n12353), .ZN(n12354) );
  OAI21_X1 U14638 ( .B1(n12447), .B2(n14935), .A(n12354), .ZN(P3_U3216) );
  XNOR2_X1 U14639 ( .A(n12355), .B(n12356), .ZN(n12357) );
  OAI222_X1 U14640 ( .A1(n14903), .A2(n12385), .B1(n14901), .B2(n12358), .C1(
        n12357), .C2(n14891), .ZN(n12448) );
  INV_X1 U14641 ( .A(n12448), .ZN(n12366) );
  XNOR2_X1 U14642 ( .A(n12360), .B(n12359), .ZN(n12449) );
  INV_X1 U14643 ( .A(n12361), .ZN(n12505) );
  AOI22_X1 U14644 ( .A1(n14935), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n14929), 
        .B2(n12362), .ZN(n12363) );
  OAI21_X1 U14645 ( .B1(n12505), .B2(n12391), .A(n12363), .ZN(n12364) );
  AOI21_X1 U14646 ( .B1(n12449), .B2(n12393), .A(n12364), .ZN(n12365) );
  OAI21_X1 U14647 ( .B1(n12366), .B2(n14935), .A(n12365), .ZN(P3_U3217) );
  XNOR2_X1 U14648 ( .A(n12367), .B(n12372), .ZN(n12371) );
  OAI22_X1 U14649 ( .A1(n12369), .A2(n14903), .B1(n12368), .B2(n14901), .ZN(
        n12370) );
  AOI21_X1 U14650 ( .B1(n12371), .B2(n14923), .A(n12370), .ZN(n12455) );
  OR2_X1 U14651 ( .A1(n12373), .A2(n12372), .ZN(n12374) );
  NAND2_X1 U14652 ( .A1(n12375), .A2(n12374), .ZN(n12453) );
  INV_X1 U14653 ( .A(n12452), .ZN(n12378) );
  AOI22_X1 U14654 ( .A1(n14935), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n14929), 
        .B2(n12376), .ZN(n12377) );
  OAI21_X1 U14655 ( .B1(n12378), .B2(n12391), .A(n12377), .ZN(n12379) );
  AOI21_X1 U14656 ( .B1(n12453), .B2(n12393), .A(n12379), .ZN(n12380) );
  OAI21_X1 U14657 ( .B1(n12455), .B2(n14935), .A(n12380), .ZN(P3_U3218) );
  XNOR2_X1 U14658 ( .A(n12381), .B(n12382), .ZN(n12383) );
  OAI222_X1 U14659 ( .A1(n14901), .A2(n12385), .B1(n14903), .B2(n12384), .C1(
        n12383), .C2(n14891), .ZN(n12456) );
  INV_X1 U14660 ( .A(n12456), .ZN(n12395) );
  XNOR2_X1 U14661 ( .A(n12386), .B(n12387), .ZN(n12457) );
  INV_X1 U14662 ( .A(n12388), .ZN(n12511) );
  AOI22_X1 U14663 ( .A1(n14935), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n14929), 
        .B2(n12389), .ZN(n12390) );
  OAI21_X1 U14664 ( .B1(n12511), .B2(n12391), .A(n12390), .ZN(n12392) );
  AOI21_X1 U14665 ( .B1(n12457), .B2(n12393), .A(n12392), .ZN(n12394) );
  OAI21_X1 U14666 ( .B1(n12395), .B2(n14935), .A(n12394), .ZN(P3_U3219) );
  NOR2_X1 U14667 ( .A1(n12460), .A2(n14987), .ZN(n12397) );
  AOI21_X1 U14668 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n14987), .A(n12397), 
        .ZN(n12396) );
  OAI21_X1 U14669 ( .B1(n12462), .B2(n12459), .A(n12396), .ZN(P3_U3490) );
  NAND2_X1 U14670 ( .A1(n12463), .A2(n9055), .ZN(n12399) );
  INV_X1 U14671 ( .A(n12397), .ZN(n12398) );
  OAI211_X1 U14672 ( .C1(n14990), .C2(n8354), .A(n12399), .B(n12398), .ZN(
        P3_U3489) );
  AOI21_X1 U14673 ( .B1(n14972), .B2(n12401), .A(n12400), .ZN(n12468) );
  MUX2_X1 U14674 ( .A(n12402), .B(n12468), .S(n14990), .Z(n12403) );
  OAI21_X1 U14675 ( .B1(n12471), .B2(n12459), .A(n12403), .ZN(P3_U3487) );
  AOI21_X1 U14676 ( .B1(n14972), .B2(n12405), .A(n12404), .ZN(n12472) );
  OAI21_X1 U14677 ( .B1(n12475), .B2(n12459), .A(n12407), .ZN(P3_U3486) );
  INV_X1 U14678 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12410) );
  AOI21_X1 U14679 ( .B1(n12409), .B2(n14972), .A(n12408), .ZN(n12476) );
  MUX2_X1 U14680 ( .A(n12410), .B(n12476), .S(n14990), .Z(n12411) );
  OAI21_X1 U14681 ( .B1(n12479), .B2(n12459), .A(n12411), .ZN(P3_U3485) );
  AOI21_X1 U14682 ( .B1(n14960), .B2(n12413), .A(n12412), .ZN(n12414) );
  OAI21_X1 U14683 ( .B1(n12421), .B2(n12415), .A(n12414), .ZN(n12480) );
  MUX2_X1 U14684 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12480), .S(n14990), .Z(
        P3_U3484) );
  AOI21_X1 U14685 ( .B1(n14972), .B2(n12417), .A(n12416), .ZN(n12481) );
  MUX2_X1 U14686 ( .A(n12418), .B(n12481), .S(n14990), .Z(n12419) );
  OAI21_X1 U14687 ( .B1(n6591), .B2(n12459), .A(n12419), .ZN(P3_U3483) );
  OAI22_X1 U14688 ( .A1(n12422), .A2(n12421), .B1(n12420), .B2(n14915), .ZN(
        n12423) );
  MUX2_X1 U14689 ( .A(n12484), .B(P3_REG1_REG_23__SCAN_IN), .S(n14987), .Z(
        P3_U3482) );
  AOI21_X1 U14690 ( .B1(n14972), .B2(n12426), .A(n12425), .ZN(n12485) );
  MUX2_X1 U14691 ( .A(n15025), .B(n12485), .S(n14990), .Z(n12427) );
  OAI21_X1 U14692 ( .B1(n12487), .B2(n12459), .A(n12427), .ZN(P3_U3481) );
  AOI21_X1 U14693 ( .B1(n14972), .B2(n12429), .A(n12428), .ZN(n12488) );
  MUX2_X1 U14694 ( .A(n12430), .B(n12488), .S(n14990), .Z(n12431) );
  OAI21_X1 U14695 ( .B1(n12491), .B2(n12459), .A(n12431), .ZN(P3_U3480) );
  AOI22_X1 U14696 ( .A1(n12433), .A2(n14972), .B1(n14960), .B2(n12432), .ZN(
        n12434) );
  NAND2_X1 U14697 ( .A1(n12435), .A2(n12434), .ZN(n12492) );
  MUX2_X1 U14698 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12492), .S(n14990), .Z(
        P3_U3479) );
  INV_X1 U14699 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12438) );
  AOI21_X1 U14700 ( .B1(n14972), .B2(n12437), .A(n12436), .ZN(n12493) );
  MUX2_X1 U14701 ( .A(n12438), .B(n12493), .S(n14990), .Z(n12439) );
  OAI21_X1 U14702 ( .B1(n12459), .B2(n12496), .A(n12439), .ZN(P3_U3478) );
  AOI21_X1 U14703 ( .B1(n12441), .B2(n14972), .A(n12440), .ZN(n12497) );
  MUX2_X1 U14704 ( .A(n12442), .B(n12497), .S(n14990), .Z(n12443) );
  OAI21_X1 U14705 ( .B1(n12500), .B2(n12459), .A(n12443), .ZN(P3_U3477) );
  AOI22_X1 U14706 ( .A1(n12445), .A2(n14972), .B1(n14960), .B2(n12444), .ZN(
        n12446) );
  NAND2_X1 U14707 ( .A1(n12447), .A2(n12446), .ZN(n12501) );
  MUX2_X1 U14708 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12501), .S(n14990), .Z(
        P3_U3476) );
  INV_X1 U14709 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12450) );
  AOI21_X1 U14710 ( .B1(n12449), .B2(n14972), .A(n12448), .ZN(n12502) );
  MUX2_X1 U14711 ( .A(n12450), .B(n12502), .S(n14990), .Z(n12451) );
  OAI21_X1 U14712 ( .B1(n12505), .B2(n12459), .A(n12451), .ZN(P3_U3475) );
  AOI22_X1 U14713 ( .A1(n12453), .A2(n14972), .B1(n14960), .B2(n12452), .ZN(
        n12454) );
  NAND2_X1 U14714 ( .A1(n12455), .A2(n12454), .ZN(n12506) );
  MUX2_X1 U14715 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n12506), .S(n14990), .Z(
        P3_U3474) );
  AOI21_X1 U14716 ( .B1(n12457), .B2(n14972), .A(n12456), .ZN(n12507) );
  MUX2_X1 U14717 ( .A(n15020), .B(n12507), .S(n14990), .Z(n12458) );
  OAI21_X1 U14718 ( .B1(n12511), .B2(n12459), .A(n12458), .ZN(P3_U3473) );
  NOR2_X1 U14719 ( .A1(n12460), .A2(n14973), .ZN(n12464) );
  AOI21_X1 U14720 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n14973), .A(n12464), 
        .ZN(n12461) );
  OAI21_X1 U14721 ( .B1(n12462), .B2(n12510), .A(n12461), .ZN(P3_U3458) );
  INV_X1 U14722 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n12467) );
  NAND2_X1 U14723 ( .A1(n12463), .A2(n9184), .ZN(n12466) );
  INV_X1 U14724 ( .A(n12464), .ZN(n12465) );
  OAI211_X1 U14725 ( .C1(n12467), .C2(n14974), .A(n12466), .B(n12465), .ZN(
        P3_U3457) );
  INV_X1 U14726 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12469) );
  MUX2_X1 U14727 ( .A(n12469), .B(n12468), .S(n14974), .Z(n12470) );
  OAI21_X1 U14728 ( .B1(n12471), .B2(n12510), .A(n12470), .ZN(P3_U3455) );
  INV_X1 U14729 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12473) );
  OAI21_X1 U14730 ( .B1(n12475), .B2(n12510), .A(n12474), .ZN(P3_U3454) );
  INV_X1 U14731 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12477) );
  MUX2_X1 U14732 ( .A(n12477), .B(n12476), .S(n14974), .Z(n12478) );
  OAI21_X1 U14733 ( .B1(n12479), .B2(n12510), .A(n12478), .ZN(P3_U3453) );
  MUX2_X1 U14734 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12480), .S(n14974), .Z(
        P3_U3452) );
  INV_X1 U14735 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12482) );
  MUX2_X1 U14736 ( .A(n12482), .B(n12481), .S(n14974), .Z(n12483) );
  OAI21_X1 U14737 ( .B1(n6591), .B2(n12510), .A(n12483), .ZN(P3_U3451) );
  MUX2_X1 U14738 ( .A(n12484), .B(P3_REG0_REG_23__SCAN_IN), .S(n14973), .Z(
        P3_U3450) );
  INV_X1 U14739 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n15022) );
  MUX2_X1 U14740 ( .A(n15022), .B(n12485), .S(n14974), .Z(n12486) );
  OAI21_X1 U14741 ( .B1(n12487), .B2(n12510), .A(n12486), .ZN(P3_U3449) );
  INV_X1 U14742 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12489) );
  MUX2_X1 U14743 ( .A(n12489), .B(n12488), .S(n14974), .Z(n12490) );
  OAI21_X1 U14744 ( .B1(n12491), .B2(n12510), .A(n12490), .ZN(P3_U3448) );
  MUX2_X1 U14745 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n12492), .S(n14974), .Z(
        P3_U3447) );
  INV_X1 U14746 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12494) );
  MUX2_X1 U14747 ( .A(n12494), .B(n12493), .S(n14974), .Z(n12495) );
  OAI21_X1 U14748 ( .B1(n12510), .B2(n12496), .A(n12495), .ZN(P3_U3446) );
  MUX2_X1 U14749 ( .A(n12498), .B(n12497), .S(n14974), .Z(n12499) );
  OAI21_X1 U14750 ( .B1(n12500), .B2(n12510), .A(n12499), .ZN(P3_U3444) );
  MUX2_X1 U14751 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12501), .S(n14974), .Z(
        P3_U3441) );
  MUX2_X1 U14752 ( .A(n12503), .B(n12502), .S(n14974), .Z(n12504) );
  OAI21_X1 U14753 ( .B1(n12505), .B2(n12510), .A(n12504), .ZN(P3_U3438) );
  MUX2_X1 U14754 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n12506), .S(n14974), .Z(
        P3_U3435) );
  MUX2_X1 U14755 ( .A(n12508), .B(n12507), .S(n14974), .Z(n12509) );
  OAI21_X1 U14756 ( .B1(n12511), .B2(n12510), .A(n12509), .ZN(P3_U3432) );
  MUX2_X1 U14757 ( .A(P3_D_REG_1__SCAN_IN), .B(n12512), .S(n12513), .Z(
        P3_U3377) );
  MUX2_X1 U14758 ( .A(P3_D_REG_0__SCAN_IN), .B(n12514), .S(n12513), .Z(
        P3_U3376) );
  NAND2_X1 U14759 ( .A1(n12516), .A2(n12515), .ZN(n12520) );
  NAND4_X1 U14760 ( .A1(n8346), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .A4(n12518), .ZN(n12519) );
  OAI211_X1 U14761 ( .C1(n15060), .C2(n12521), .A(n12520), .B(n12519), .ZN(
        P3_U3264) );
  INV_X1 U14762 ( .A(n12522), .ZN(n12525) );
  OAI222_X1 U14763 ( .A1(n12528), .A2(n12525), .B1(n12524), .B2(P3_U3151), 
        .C1(n12523), .C2(n12530), .ZN(P3_U3266) );
  INV_X1 U14764 ( .A(n12526), .ZN(n12527) );
  OAI222_X1 U14765 ( .A1(P3_U3151), .A2(n12531), .B1(n12530), .B2(n12529), 
        .C1(n12528), .C2(n12527), .ZN(P3_U3267) );
  INV_X1 U14766 ( .A(n12532), .ZN(n12533) );
  NOR2_X1 U14767 ( .A1(n13056), .A2(n6438), .ZN(n12714) );
  NOR2_X1 U14768 ( .A1(n12648), .A2(n6438), .ZN(n12537) );
  XNOR2_X1 U14769 ( .A(n13074), .B(n12576), .ZN(n12536) );
  NOR2_X1 U14770 ( .A1(n12536), .A2(n12537), .ZN(n12538) );
  AOI21_X1 U14771 ( .B1(n12537), .B2(n12536), .A(n12538), .ZN(n12638) );
  INV_X1 U14772 ( .A(n12538), .ZN(n12539) );
  NAND2_X1 U14773 ( .A1(n12636), .A2(n12539), .ZN(n12645) );
  NOR2_X1 U14774 ( .A1(n13058), .A2(n6438), .ZN(n12541) );
  XNOR2_X1 U14775 ( .A(n13045), .B(n12576), .ZN(n12540) );
  NOR2_X1 U14776 ( .A1(n12540), .A2(n12541), .ZN(n12542) );
  AOI21_X1 U14777 ( .B1(n12541), .B2(n12540), .A(n12542), .ZN(n12646) );
  INV_X1 U14778 ( .A(n12542), .ZN(n12543) );
  XNOR2_X1 U14779 ( .A(n13036), .B(n6816), .ZN(n12544) );
  NOR2_X1 U14780 ( .A1(n13014), .A2(n6438), .ZN(n12545) );
  XNOR2_X1 U14781 ( .A(n12544), .B(n12545), .ZN(n12696) );
  INV_X1 U14782 ( .A(n12544), .ZN(n12546) );
  NOR2_X1 U14783 ( .A1(n12697), .A2(n6438), .ZN(n12548) );
  NOR2_X1 U14784 ( .A1(n12547), .A2(n12548), .ZN(n12549) );
  AOI21_X1 U14785 ( .B1(n12548), .B2(n12547), .A(n12549), .ZN(n12589) );
  AND2_X1 U14786 ( .A1(n12976), .A2(n10022), .ZN(n12551) );
  XNOR2_X1 U14787 ( .A(n13142), .B(n6816), .ZN(n12550) );
  NOR2_X1 U14788 ( .A1(n12550), .A2(n12551), .ZN(n12552) );
  AOI21_X1 U14789 ( .B1(n12551), .B2(n12550), .A(n12552), .ZN(n12665) );
  NAND2_X1 U14790 ( .A1(n12664), .A2(n12665), .ZN(n12663) );
  INV_X1 U14791 ( .A(n12552), .ZN(n12553) );
  NAND2_X1 U14792 ( .A1(n13005), .A2(n10022), .ZN(n12555) );
  XNOR2_X1 U14793 ( .A(n13134), .B(n6816), .ZN(n12554) );
  XOR2_X1 U14794 ( .A(n12555), .B(n12554), .Z(n12618) );
  INV_X1 U14795 ( .A(n12554), .ZN(n12556) );
  XNOR2_X1 U14796 ( .A(n13129), .B(n6816), .ZN(n12558) );
  XNOR2_X1 U14797 ( .A(n12557), .B(n12558), .ZN(n12673) );
  NOR2_X1 U14798 ( .A1(n12621), .A2(n6438), .ZN(n12672) );
  XNOR2_X1 U14799 ( .A(n12954), .B(n12576), .ZN(n12561) );
  INV_X1 U14800 ( .A(n12561), .ZN(n12563) );
  NOR2_X1 U14801 ( .A1(n12675), .A2(n6438), .ZN(n12582) );
  NAND2_X1 U14802 ( .A1(n12583), .A2(n12582), .ZN(n12562) );
  OAI21_X1 U14803 ( .B1(n12564), .B2(n12563), .A(n12562), .ZN(n12655) );
  XNOR2_X1 U14804 ( .A(n12939), .B(n6816), .ZN(n12565) );
  NOR2_X1 U14805 ( .A1(n12631), .A2(n6438), .ZN(n12566) );
  XNOR2_X1 U14806 ( .A(n12565), .B(n12566), .ZN(n12654) );
  INV_X1 U14807 ( .A(n12565), .ZN(n12567) );
  NAND2_X1 U14808 ( .A1(n12567), .A2(n12566), .ZN(n12568) );
  XNOR2_X1 U14809 ( .A(n12923), .B(n6816), .ZN(n12569) );
  NOR2_X1 U14810 ( .A1(n12657), .A2(n6438), .ZN(n12570) );
  XNOR2_X1 U14811 ( .A(n12569), .B(n12570), .ZN(n12627) );
  INV_X1 U14812 ( .A(n12569), .ZN(n12571) );
  NAND2_X1 U14813 ( .A1(n12571), .A2(n12570), .ZN(n12572) );
  XNOR2_X1 U14814 ( .A(n12909), .B(n6816), .ZN(n12574) );
  NAND2_X1 U14815 ( .A1(n12918), .A2(n10022), .ZN(n12573) );
  NAND2_X1 U14816 ( .A1(n12574), .A2(n12573), .ZN(n12575) );
  OAI21_X1 U14817 ( .B1(n12574), .B2(n12573), .A(n12575), .ZN(n12706) );
  OR2_X2 U14818 ( .A1(n12707), .A2(n12706), .ZN(n12704) );
  XNOR2_X1 U14819 ( .A(n13103), .B(n12576), .ZN(n12598) );
  NAND2_X1 U14820 ( .A1(n12727), .A2(n10022), .ZN(n12597) );
  XNOR2_X1 U14821 ( .A(n12598), .B(n12597), .ZN(n12600) );
  XNOR2_X1 U14822 ( .A(n12601), .B(n12600), .ZN(n12581) );
  OAI22_X1 U14823 ( .A1(n12602), .A2(n12656), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12577), .ZN(n12579) );
  OAI22_X1 U14824 ( .A1(n12629), .A2(n12658), .B1(n12893), .B2(n12720), .ZN(
        n12578) );
  AOI211_X1 U14825 ( .C1(n13103), .C2(n12722), .A(n12579), .B(n12578), .ZN(
        n12580) );
  OAI21_X1 U14826 ( .B1(n12581), .B2(n12724), .A(n12580), .ZN(P2_U3186) );
  XNOR2_X1 U14827 ( .A(n12583), .B(n12582), .ZN(n12587) );
  OAI22_X1 U14828 ( .A1(n12631), .A2(n13057), .B1(n12621), .B2(n13055), .ZN(
        n13123) );
  AOI22_X1 U14829 ( .A1(n13123), .A2(n12717), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12584) );
  OAI21_X1 U14830 ( .B1(n12950), .B2(n12720), .A(n12584), .ZN(n12585) );
  AOI21_X1 U14831 ( .B1(n13124), .B2(n12722), .A(n12585), .ZN(n12586) );
  OAI21_X1 U14832 ( .B1(n12587), .B2(n12724), .A(n12586), .ZN(P2_U3188) );
  OAI21_X1 U14833 ( .B1(n12590), .B2(n12589), .A(n12588), .ZN(n12591) );
  NAND2_X1 U14834 ( .A1(n12591), .A2(n12689), .ZN(n12596) );
  INV_X1 U14835 ( .A(n13019), .ZN(n12592) );
  OAI22_X1 U14836 ( .A1(n12658), .A2(n13014), .B1(n12592), .B2(n12720), .ZN(
        n12593) );
  AOI211_X1 U14837 ( .C1(n12685), .C2(n12976), .A(n12594), .B(n12593), .ZN(
        n12595) );
  OAI211_X1 U14838 ( .C1(n13022), .C2(n12653), .A(n12596), .B(n12595), .ZN(
        P2_U3191) );
  NOR2_X1 U14839 ( .A1(n12602), .A2(n6438), .ZN(n12603) );
  XOR2_X1 U14840 ( .A(n6816), .B(n12603), .Z(n12605) );
  XNOR2_X1 U14841 ( .A(n13096), .B(n12605), .ZN(n12606) );
  AOI22_X1 U14842 ( .A1(n12869), .A2(n12685), .B1(n12875), .B2(n12708), .ZN(
        n12608) );
  AOI22_X1 U14843 ( .A1(n12727), .A2(n12683), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12607) );
  NAND2_X1 U14844 ( .A1(n12608), .A2(n12607), .ZN(n12609) );
  AOI21_X1 U14845 ( .B1(n13096), .B2(n12722), .A(n12609), .ZN(n12610) );
  AOI22_X1 U14846 ( .A1(n12683), .A2(n12746), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n12682), .ZN(n12617) );
  AOI22_X1 U14847 ( .A1(n12685), .A2(n12744), .B1(n10021), .B2(n12722), .ZN(
        n12616) );
  NOR2_X1 U14848 ( .A1(n12613), .A2(n12612), .ZN(n12614) );
  OAI21_X1 U14849 ( .B1(n12611), .B2(n12614), .A(n12689), .ZN(n12615) );
  NAND3_X1 U14850 ( .A1(n12617), .A2(n12616), .A3(n12615), .ZN(P2_U3194) );
  XNOR2_X1 U14851 ( .A(n12619), .B(n12618), .ZN(n12625) );
  OAI22_X1 U14852 ( .A1(n12656), .A2(n12621), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12620), .ZN(n12623) );
  OAI22_X1 U14853 ( .A1(n12658), .A2(n13015), .B1(n12980), .B2(n12720), .ZN(
        n12622) );
  AOI211_X1 U14854 ( .C1(n13134), .C2(n12722), .A(n12623), .B(n12622), .ZN(
        n12624) );
  OAI21_X1 U14855 ( .B1(n12625), .B2(n12724), .A(n12624), .ZN(P2_U3195) );
  XNOR2_X1 U14856 ( .A(n12626), .B(n12627), .ZN(n12635) );
  OAI22_X1 U14857 ( .A1(n12629), .A2(n12656), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12628), .ZN(n12633) );
  INV_X1 U14858 ( .A(n12921), .ZN(n12630) );
  OAI22_X1 U14859 ( .A1(n12658), .A2(n12631), .B1(n12630), .B2(n12720), .ZN(
        n12632) );
  AOI211_X1 U14860 ( .C1(n13113), .C2(n12722), .A(n12633), .B(n12632), .ZN(
        n12634) );
  OAI21_X1 U14861 ( .B1(n12635), .B2(n12724), .A(n12634), .ZN(P2_U3197) );
  OAI21_X1 U14862 ( .B1(n12638), .B2(n12637), .A(n12636), .ZN(n12639) );
  NAND2_X1 U14863 ( .A1(n12639), .A2(n12689), .ZN(n12643) );
  NAND2_X1 U14864 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n14600)
         );
  INV_X1 U14865 ( .A(n14600), .ZN(n12641) );
  OAI22_X1 U14866 ( .A1(n12658), .A2(n13056), .B1(n13070), .B2(n12720), .ZN(
        n12640) );
  AOI211_X1 U14867 ( .C1(n12685), .C2(n12729), .A(n12641), .B(n12640), .ZN(
        n12642) );
  OAI211_X1 U14868 ( .C1(n13074), .C2(n12653), .A(n12643), .B(n12642), .ZN(
        P2_U3198) );
  OAI21_X1 U14869 ( .B1(n12646), .B2(n12645), .A(n12644), .ZN(n12647) );
  NAND2_X1 U14870 ( .A1(n12647), .A2(n12689), .ZN(n12652) );
  OAI22_X1 U14871 ( .A1(n13014), .A2(n13057), .B1(n12648), .B2(n13055), .ZN(
        n13048) );
  NAND2_X1 U14872 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14613)
         );
  INV_X1 U14873 ( .A(n14613), .ZN(n12650) );
  NOR2_X1 U14874 ( .A1(n12720), .A2(n13042), .ZN(n12649) );
  AOI211_X1 U14875 ( .C1(n12717), .C2(n13048), .A(n12650), .B(n12649), .ZN(
        n12651) );
  OAI211_X1 U14876 ( .C1(n13045), .C2(n12653), .A(n12652), .B(n12651), .ZN(
        P2_U3200) );
  XNOR2_X1 U14877 ( .A(n12655), .B(n12654), .ZN(n12662) );
  OAI22_X1 U14878 ( .A1(n12657), .A2(n12656), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n15051), .ZN(n12660) );
  OAI22_X1 U14879 ( .A1(n12658), .A2(n12675), .B1(n12936), .B2(n12720), .ZN(
        n12659) );
  AOI211_X1 U14880 ( .C1(n13118), .C2(n12722), .A(n12660), .B(n12659), .ZN(
        n12661) );
  OAI21_X1 U14881 ( .B1(n12662), .B2(n12724), .A(n12661), .ZN(P2_U3201) );
  OAI21_X1 U14882 ( .B1(n12665), .B2(n12664), .A(n12663), .ZN(n12666) );
  NAND2_X1 U14883 ( .A1(n12666), .A2(n12689), .ZN(n12671) );
  AOI22_X1 U14884 ( .A1(n12685), .A2(n13005), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12670) );
  INV_X1 U14885 ( .A(n12997), .ZN(n12667) );
  AOI22_X1 U14886 ( .A1(n12683), .A2(n13003), .B1(n12667), .B2(n12708), .ZN(
        n12669) );
  NAND2_X1 U14887 ( .A1(n13142), .A2(n12722), .ZN(n12668) );
  NAND4_X1 U14888 ( .A1(n12671), .A2(n12670), .A3(n12669), .A4(n12668), .ZN(
        P2_U3205) );
  XNOR2_X1 U14889 ( .A(n12673), .B(n12672), .ZN(n12681) );
  INV_X1 U14890 ( .A(n12968), .ZN(n12677) );
  OAI22_X1 U14891 ( .A1(n12675), .A2(n13057), .B1(n12674), .B2(n13055), .ZN(
        n12960) );
  AOI22_X1 U14892 ( .A1(n12960), .A2(n12717), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12676) );
  OAI21_X1 U14893 ( .B1(n12677), .B2(n12720), .A(n12676), .ZN(n12678) );
  AOI21_X1 U14894 ( .B1(n12679), .B2(n12722), .A(n12678), .ZN(n12680) );
  OAI21_X1 U14895 ( .B1(n12681), .B2(n12724), .A(n12680), .ZN(P2_U3207) );
  AOI22_X1 U14896 ( .A1(n12683), .A2(n12745), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n12682), .ZN(n12694) );
  AOI22_X1 U14897 ( .A1(n12685), .A2(n12743), .B1(n12684), .B2(n12722), .ZN(
        n12693) );
  INV_X1 U14898 ( .A(n12686), .ZN(n12691) );
  NOR3_X1 U14899 ( .A1(n12611), .A2(n12688), .A3(n12687), .ZN(n12690) );
  OAI21_X1 U14900 ( .B1(n12691), .B2(n12690), .A(n12689), .ZN(n12692) );
  NAND3_X1 U14901 ( .A1(n12694), .A2(n12693), .A3(n12692), .ZN(P2_U3209) );
  XNOR2_X1 U14902 ( .A(n12695), .B(n12696), .ZN(n12703) );
  OR2_X1 U14903 ( .A1(n12697), .A2(n13057), .ZN(n12699) );
  NAND2_X1 U14904 ( .A1(n12729), .A2(n13002), .ZN(n12698) );
  AND2_X1 U14905 ( .A1(n12699), .A2(n12698), .ZN(n13028) );
  NAND2_X1 U14906 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n14626)
         );
  NAND2_X1 U14907 ( .A1(n12708), .A2(n13033), .ZN(n12700) );
  OAI211_X1 U14908 ( .C1(n12710), .C2(n13028), .A(n14626), .B(n12700), .ZN(
        n12701) );
  AOI21_X1 U14909 ( .B1(n13153), .B2(n12722), .A(n12701), .ZN(n12702) );
  OAI21_X1 U14910 ( .B1(n12703), .B2(n12724), .A(n12702), .ZN(P2_U3210) );
  INV_X1 U14911 ( .A(n12704), .ZN(n12705) );
  AOI21_X1 U14912 ( .B1(n12707), .B2(n12706), .A(n12705), .ZN(n12713) );
  AOI22_X1 U14913 ( .A1(n12727), .A2(n13004), .B1(n13002), .B2(n12932), .ZN(
        n12901) );
  AOI22_X1 U14914 ( .A1(n12907), .A2(n12708), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12709) );
  OAI21_X1 U14915 ( .B1(n12901), .B2(n12710), .A(n12709), .ZN(n12711) );
  AOI21_X1 U14916 ( .B1(n13108), .B2(n12722), .A(n12711), .ZN(n12712) );
  OAI21_X1 U14917 ( .B1(n12713), .B2(n12724), .A(n12712), .ZN(P2_U3212) );
  XNOR2_X1 U14918 ( .A(n12715), .B(n12714), .ZN(n12725) );
  AOI22_X1 U14919 ( .A1(n12717), .A2(n12716), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12718) );
  OAI21_X1 U14920 ( .B1(n12720), .B2(n12719), .A(n12718), .ZN(n12721) );
  AOI21_X1 U14921 ( .B1(n13167), .B2(n12722), .A(n12721), .ZN(n12723) );
  OAI21_X1 U14922 ( .B1(n12725), .B2(n12724), .A(n12723), .ZN(P2_U3213) );
  INV_X2 U14923 ( .A(P2_U3947), .ZN(n12737) );
  MUX2_X1 U14924 ( .A(n12847), .B(P2_DATAO_REG_31__SCAN_IN), .S(n12737), .Z(
        P2_U3562) );
  MUX2_X1 U14925 ( .A(n12726), .B(P2_DATAO_REG_30__SCAN_IN), .S(n12737), .Z(
        P2_U3561) );
  MUX2_X1 U14926 ( .A(n12869), .B(P2_DATAO_REG_29__SCAN_IN), .S(n12737), .Z(
        P2_U3560) );
  MUX2_X1 U14927 ( .A(n12887), .B(P2_DATAO_REG_28__SCAN_IN), .S(n12737), .Z(
        P2_U3559) );
  MUX2_X1 U14928 ( .A(n12727), .B(P2_DATAO_REG_27__SCAN_IN), .S(n12737), .Z(
        P2_U3558) );
  MUX2_X1 U14929 ( .A(n12918), .B(P2_DATAO_REG_26__SCAN_IN), .S(n12737), .Z(
        P2_U3557) );
  MUX2_X1 U14930 ( .A(n12932), .B(P2_DATAO_REG_25__SCAN_IN), .S(n12737), .Z(
        P2_U3556) );
  MUX2_X1 U14931 ( .A(n12917), .B(P2_DATAO_REG_24__SCAN_IN), .S(n12737), .Z(
        P2_U3555) );
  MUX2_X1 U14932 ( .A(n12931), .B(P2_DATAO_REG_23__SCAN_IN), .S(n12737), .Z(
        P2_U3554) );
  MUX2_X1 U14933 ( .A(n12975), .B(P2_DATAO_REG_22__SCAN_IN), .S(n12737), .Z(
        P2_U3553) );
  MUX2_X1 U14934 ( .A(n13005), .B(P2_DATAO_REG_21__SCAN_IN), .S(n12737), .Z(
        P2_U3552) );
  MUX2_X1 U14935 ( .A(n12976), .B(P2_DATAO_REG_20__SCAN_IN), .S(n12737), .Z(
        P2_U3551) );
  MUX2_X1 U14936 ( .A(n13003), .B(P2_DATAO_REG_19__SCAN_IN), .S(n12737), .Z(
        P2_U3550) );
  MUX2_X1 U14937 ( .A(n12728), .B(P2_DATAO_REG_18__SCAN_IN), .S(n12737), .Z(
        P2_U3549) );
  MUX2_X1 U14938 ( .A(n12729), .B(P2_DATAO_REG_17__SCAN_IN), .S(n12737), .Z(
        P2_U3548) );
  MUX2_X1 U14939 ( .A(n7136), .B(P2_DATAO_REG_16__SCAN_IN), .S(n12737), .Z(
        P2_U3547) );
  MUX2_X1 U14940 ( .A(n12730), .B(P2_DATAO_REG_15__SCAN_IN), .S(n12737), .Z(
        P2_U3546) );
  MUX2_X1 U14941 ( .A(n12731), .B(P2_DATAO_REG_14__SCAN_IN), .S(n12737), .Z(
        P2_U3545) );
  MUX2_X1 U14942 ( .A(n12732), .B(P2_DATAO_REG_13__SCAN_IN), .S(n12737), .Z(
        P2_U3544) );
  MUX2_X1 U14943 ( .A(n12733), .B(P2_DATAO_REG_12__SCAN_IN), .S(n12737), .Z(
        P2_U3543) );
  MUX2_X1 U14944 ( .A(n12734), .B(P2_DATAO_REG_11__SCAN_IN), .S(n12737), .Z(
        P2_U3542) );
  MUX2_X1 U14945 ( .A(n12735), .B(P2_DATAO_REG_10__SCAN_IN), .S(n12737), .Z(
        P2_U3541) );
  MUX2_X1 U14946 ( .A(n12736), .B(P2_DATAO_REG_9__SCAN_IN), .S(n12737), .Z(
        P2_U3540) );
  MUX2_X1 U14947 ( .A(n12738), .B(P2_DATAO_REG_8__SCAN_IN), .S(n12737), .Z(
        P2_U3539) );
  MUX2_X1 U14948 ( .A(n12739), .B(P2_DATAO_REG_7__SCAN_IN), .S(n12737), .Z(
        P2_U3538) );
  MUX2_X1 U14949 ( .A(n12740), .B(P2_DATAO_REG_6__SCAN_IN), .S(n12737), .Z(
        P2_U3537) );
  MUX2_X1 U14950 ( .A(n12741), .B(P2_DATAO_REG_5__SCAN_IN), .S(n12737), .Z(
        P2_U3536) );
  MUX2_X1 U14951 ( .A(n12742), .B(P2_DATAO_REG_4__SCAN_IN), .S(n12737), .Z(
        P2_U3535) );
  MUX2_X1 U14952 ( .A(n12743), .B(P2_DATAO_REG_3__SCAN_IN), .S(n12737), .Z(
        P2_U3534) );
  MUX2_X1 U14953 ( .A(n12744), .B(P2_DATAO_REG_2__SCAN_IN), .S(n12737), .Z(
        P2_U3533) );
  MUX2_X1 U14954 ( .A(n12745), .B(P2_DATAO_REG_1__SCAN_IN), .S(n12737), .Z(
        P2_U3532) );
  MUX2_X1 U14955 ( .A(n12746), .B(P2_DATAO_REG_0__SCAN_IN), .S(n12737), .Z(
        P2_U3531) );
  OAI22_X1 U14956 ( .A1(n14624), .A2(n12749), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12747), .ZN(n12748) );
  AOI21_X1 U14957 ( .B1(n14577), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n12748), .ZN(
        n12759) );
  MUX2_X1 U14958 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9459), .S(n12749), .Z(
        n12750) );
  OAI21_X1 U14959 ( .B1(n9836), .B2(n12751), .A(n12750), .ZN(n12752) );
  NAND3_X1 U14960 ( .A1(n14579), .A2(n12753), .A3(n12752), .ZN(n12758) );
  OAI211_X1 U14961 ( .C1(n12756), .C2(n12755), .A(n14582), .B(n12754), .ZN(
        n12757) );
  NAND3_X1 U14962 ( .A1(n12759), .A2(n12758), .A3(n12757), .ZN(P2_U3215) );
  OAI22_X1 U14963 ( .A1(n14624), .A2(n12761), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12760), .ZN(n12762) );
  AOI21_X1 U14964 ( .B1(n14577), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n12762), .ZN(
        n12771) );
  OAI211_X1 U14965 ( .C1(n12765), .C2(n12764), .A(n14579), .B(n12763), .ZN(
        n12770) );
  OAI211_X1 U14966 ( .C1(n12768), .C2(n12767), .A(n14582), .B(n12766), .ZN(
        n12769) );
  NAND3_X1 U14967 ( .A1(n12771), .A2(n12770), .A3(n12769), .ZN(P2_U3216) );
  AOI22_X1 U14968 ( .A1(n14577), .A2(P2_ADDR_REG_4__SCAN_IN), .B1(n14585), 
        .B2(n12777), .ZN(n12785) );
  OAI211_X1 U14969 ( .C1(n12774), .C2(n12773), .A(n14582), .B(n12772), .ZN(
        n12775) );
  AND2_X1 U14970 ( .A1(n12776), .A2(n12775), .ZN(n12784) );
  MUX2_X1 U14971 ( .A(n9469), .B(P2_REG1_REG_4__SCAN_IN), .S(n12777), .Z(
        n12778) );
  NAND3_X1 U14972 ( .A1(n12780), .A2(n12779), .A3(n12778), .ZN(n12781) );
  NAND3_X1 U14973 ( .A1(n14579), .A2(n12782), .A3(n12781), .ZN(n12783) );
  NAND3_X1 U14974 ( .A1(n12785), .A2(n12784), .A3(n12783), .ZN(P2_U3218) );
  OAI21_X1 U14975 ( .B1(n14624), .B2(n12787), .A(n12786), .ZN(n12788) );
  AOI21_X1 U14976 ( .B1(n14577), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n12788), .ZN(
        n12800) );
  MUX2_X1 U14977 ( .A(n10443), .B(P2_REG2_REG_6__SCAN_IN), .S(n12793), .Z(
        n12789) );
  NAND3_X1 U14978 ( .A1(n12791), .A2(n12790), .A3(n12789), .ZN(n12792) );
  NAND3_X1 U14979 ( .A1(n14582), .A2(n12806), .A3(n12792), .ZN(n12799) );
  INV_X1 U14980 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n14729) );
  MUX2_X1 U14981 ( .A(n14729), .B(P2_REG1_REG_6__SCAN_IN), .S(n12793), .Z(
        n12794) );
  NAND3_X1 U14982 ( .A1(n12796), .A2(n12795), .A3(n12794), .ZN(n12797) );
  NAND3_X1 U14983 ( .A1(n14579), .A2(n12811), .A3(n12797), .ZN(n12798) );
  NAND3_X1 U14984 ( .A1(n12800), .A2(n12799), .A3(n12798), .ZN(P2_U3220) );
  NOR2_X1 U14985 ( .A1(n14624), .A2(n12801), .ZN(n12802) );
  AOI211_X1 U14986 ( .C1(n14577), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n12803), .B(
        n12802), .ZN(n12815) );
  MUX2_X1 U14987 ( .A(n10455), .B(P2_REG2_REG_7__SCAN_IN), .S(n12808), .Z(
        n12804) );
  NAND3_X1 U14988 ( .A1(n12806), .A2(n12805), .A3(n12804), .ZN(n12807) );
  NAND3_X1 U14989 ( .A1(n14582), .A2(n12821), .A3(n12807), .ZN(n12814) );
  MUX2_X1 U14990 ( .A(n9477), .B(P2_REG1_REG_7__SCAN_IN), .S(n12808), .Z(
        n12809) );
  NAND3_X1 U14991 ( .A1(n12811), .A2(n12810), .A3(n12809), .ZN(n12812) );
  NAND3_X1 U14992 ( .A1(n14579), .A2(n12827), .A3(n12812), .ZN(n12813) );
  NAND3_X1 U14993 ( .A1(n12815), .A2(n12814), .A3(n12813), .ZN(P2_U3221) );
  NOR2_X1 U14994 ( .A1(n14624), .A2(n12816), .ZN(n12817) );
  AOI211_X1 U14995 ( .C1(n14577), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n12818), .B(
        n12817), .ZN(n12832) );
  MUX2_X1 U14996 ( .A(n10729), .B(P2_REG2_REG_8__SCAN_IN), .S(n12824), .Z(
        n12819) );
  NAND3_X1 U14997 ( .A1(n12821), .A2(n12820), .A3(n12819), .ZN(n12822) );
  NAND3_X1 U14998 ( .A1(n12823), .A2(n14582), .A3(n12822), .ZN(n12831) );
  MUX2_X1 U14999 ( .A(n9480), .B(P2_REG1_REG_8__SCAN_IN), .S(n12824), .Z(
        n12825) );
  NAND3_X1 U15000 ( .A1(n12827), .A2(n12826), .A3(n12825), .ZN(n12828) );
  NAND3_X1 U15001 ( .A1(n12829), .A2(n14579), .A3(n12828), .ZN(n12830) );
  NAND3_X1 U15002 ( .A1(n12832), .A2(n12831), .A3(n12830), .ZN(P2_U3222) );
  OAI211_X1 U15003 ( .C1(n12835), .C2(n12834), .A(n12833), .B(n14582), .ZN(
        n12844) );
  OAI211_X1 U15004 ( .C1(n12838), .C2(n12837), .A(n12836), .B(n14579), .ZN(
        n12843) );
  AOI21_X1 U15005 ( .B1(n14585), .B2(n12840), .A(n12839), .ZN(n12842) );
  NAND2_X1 U15006 ( .A1(n14577), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n12841) );
  NAND4_X1 U15007 ( .A1(n12844), .A2(n12843), .A3(n12842), .A4(n12841), .ZN(
        P2_U3224) );
  NAND2_X1 U15008 ( .A1(n12852), .A2(n13094), .ZN(n12851) );
  INV_X1 U15009 ( .A(n12845), .ZN(n12846) );
  NAND2_X1 U15010 ( .A1(n12847), .A2(n12846), .ZN(n13092) );
  NOR2_X1 U15011 ( .A1(n13078), .A2(n13092), .ZN(n12854) );
  NOR2_X1 U15012 ( .A1(n6837), .A2(n13073), .ZN(n12849) );
  AOI211_X1 U15013 ( .C1(n13078), .C2(P2_REG2_REG_31__SCAN_IN), .A(n12854), 
        .B(n12849), .ZN(n12850) );
  OAI21_X1 U15014 ( .B1(n12984), .B2(n13091), .A(n12850), .ZN(P2_U3234) );
  OAI211_X1 U15015 ( .C1(n12852), .C2(n13094), .A(n12851), .B(n6438), .ZN(
        n13093) );
  NOR2_X1 U15016 ( .A1(n13038), .A2(n12853), .ZN(n12855) );
  AOI211_X1 U15017 ( .C1(n12856), .C2(n13082), .A(n12855), .B(n12854), .ZN(
        n12857) );
  OAI21_X1 U15018 ( .B1(n13093), .B2(n12984), .A(n12857), .ZN(P2_U3235) );
  INV_X1 U15019 ( .A(n12858), .ZN(n12861) );
  AOI22_X1 U15020 ( .A1(n12859), .A2(n13081), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13078), .ZN(n12860) );
  OAI21_X1 U15021 ( .B1(n12861), .B2(n13073), .A(n12860), .ZN(n12863) );
  INV_X1 U15022 ( .A(n12869), .ZN(n12871) );
  OAI22_X1 U15023 ( .A1(n12871), .A2(n13057), .B1(n12870), .B2(n13055), .ZN(
        n12872) );
  AOI21_X1 U15024 ( .B1(n13096), .B2(n12892), .A(n10022), .ZN(n12874) );
  NAND2_X1 U15025 ( .A1(n13096), .A2(n13082), .ZN(n12877) );
  AOI22_X1 U15026 ( .A1(n12875), .A2(n13081), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n13078), .ZN(n12876) );
  NAND2_X1 U15027 ( .A1(n12877), .A2(n12876), .ZN(n12878) );
  AOI21_X1 U15028 ( .B1(n13095), .B2(n13085), .A(n12878), .ZN(n12882) );
  XNOR2_X1 U15029 ( .A(n12880), .B(n12879), .ZN(n13098) );
  OR2_X1 U15030 ( .A1(n13098), .A2(n13053), .ZN(n12881) );
  OAI211_X1 U15031 ( .C1(n13101), .C2(n13078), .A(n12882), .B(n12881), .ZN(
        P2_U3237) );
  XNOR2_X1 U15032 ( .A(n12883), .B(n12884), .ZN(n13106) );
  NAND2_X1 U15033 ( .A1(n12887), .A2(n13004), .ZN(n12889) );
  NAND2_X1 U15034 ( .A1(n12918), .A2(n13002), .ZN(n12888) );
  OR2_X1 U15035 ( .A1(n13105), .A2(n13078), .ZN(n12899) );
  AOI211_X1 U15036 ( .C1(n13103), .C2(n12904), .A(n10022), .B(n6799), .ZN(
        n13102) );
  INV_X1 U15037 ( .A(n12893), .ZN(n12894) );
  AOI22_X1 U15038 ( .A1(n12894), .A2(n13081), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13078), .ZN(n12895) );
  OAI21_X1 U15039 ( .B1(n12896), .B2(n13073), .A(n12895), .ZN(n12897) );
  AOI21_X1 U15040 ( .B1(n13102), .B2(n13085), .A(n12897), .ZN(n12898) );
  OAI211_X1 U15041 ( .C1(n13106), .C2(n13053), .A(n12899), .B(n12898), .ZN(
        P2_U3238) );
  XNOR2_X1 U15042 ( .A(n12900), .B(n12911), .ZN(n12903) );
  INV_X1 U15043 ( .A(n12901), .ZN(n12902) );
  INV_X1 U15044 ( .A(n12920), .ZN(n12906) );
  INV_X1 U15045 ( .A(n12904), .ZN(n12905) );
  AOI211_X1 U15046 ( .C1(n13108), .C2(n12906), .A(n10022), .B(n12905), .ZN(
        n13107) );
  AOI22_X1 U15047 ( .A1(n12907), .A2(n13081), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13078), .ZN(n12908) );
  OAI21_X1 U15048 ( .B1(n12909), .B2(n13073), .A(n12908), .ZN(n12913) );
  XOR2_X1 U15049 ( .A(n12911), .B(n12910), .Z(n13111) );
  NOR2_X1 U15050 ( .A1(n13111), .A2(n13053), .ZN(n12912) );
  AOI211_X1 U15051 ( .C1(n13107), .C2(n13085), .A(n12913), .B(n12912), .ZN(
        n12914) );
  OAI21_X1 U15052 ( .B1(n13110), .B2(n13078), .A(n12914), .ZN(P2_U3239) );
  XNOR2_X1 U15053 ( .A(n12916), .B(n12915), .ZN(n12919) );
  AOI222_X1 U15054 ( .A1(n13065), .A2(n12919), .B1(n12918), .B2(n13004), .C1(
        n12917), .C2(n13002), .ZN(n13115) );
  AOI211_X1 U15055 ( .C1(n13113), .C2(n12934), .A(n10022), .B(n12920), .ZN(
        n13112) );
  AOI22_X1 U15056 ( .A1(n12921), .A2(n13081), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13078), .ZN(n12922) );
  OAI21_X1 U15057 ( .B1(n12923), .B2(n13073), .A(n12922), .ZN(n12927) );
  XNOR2_X1 U15058 ( .A(n12925), .B(n12924), .ZN(n13116) );
  NOR2_X1 U15059 ( .A1(n13116), .A2(n13053), .ZN(n12926) );
  AOI211_X1 U15060 ( .C1(n13112), .C2(n13085), .A(n12927), .B(n12926), .ZN(
        n12928) );
  OAI21_X1 U15061 ( .B1(n13115), .B2(n13078), .A(n12928), .ZN(P2_U3240) );
  XNOR2_X1 U15062 ( .A(n12930), .B(n12929), .ZN(n12933) );
  AOI222_X1 U15063 ( .A1(n13065), .A2(n12933), .B1(n12932), .B2(n13004), .C1(
        n12931), .C2(n13002), .ZN(n13120) );
  INV_X1 U15064 ( .A(n12934), .ZN(n12935) );
  AOI211_X1 U15065 ( .C1(n13118), .C2(n12952), .A(n10022), .B(n12935), .ZN(
        n13117) );
  INV_X1 U15066 ( .A(n12936), .ZN(n12937) );
  AOI22_X1 U15067 ( .A1(n12937), .A2(n13081), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13078), .ZN(n12938) );
  OAI21_X1 U15068 ( .B1(n12939), .B2(n13073), .A(n12938), .ZN(n12943) );
  XNOR2_X1 U15069 ( .A(n12941), .B(n12940), .ZN(n13121) );
  NOR2_X1 U15070 ( .A1(n13121), .A2(n13053), .ZN(n12942) );
  AOI211_X1 U15071 ( .C1(n13117), .C2(n13085), .A(n12943), .B(n12942), .ZN(
        n12944) );
  OAI21_X1 U15072 ( .B1(n13120), .B2(n13078), .A(n12944), .ZN(P2_U3241) );
  XOR2_X1 U15073 ( .A(n12946), .B(n12945), .Z(n13127) );
  XNOR2_X1 U15074 ( .A(n12947), .B(n12946), .ZN(n12948) );
  NAND2_X1 U15075 ( .A1(n12948), .A2(n13065), .ZN(n13126) );
  INV_X1 U15076 ( .A(n13123), .ZN(n12949) );
  OAI211_X1 U15077 ( .C1(n12998), .C2(n12950), .A(n13126), .B(n12949), .ZN(
        n12951) );
  NAND2_X1 U15078 ( .A1(n12951), .A2(n13038), .ZN(n12957) );
  AOI211_X1 U15079 ( .C1(n13124), .C2(n12966), .A(n10022), .B(n7007), .ZN(
        n13122) );
  INV_X1 U15080 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n12953) );
  OAI22_X1 U15081 ( .A1(n12954), .A2(n13073), .B1(n13038), .B2(n12953), .ZN(
        n12955) );
  AOI21_X1 U15082 ( .B1(n13122), .B2(n13085), .A(n12955), .ZN(n12956) );
  OAI211_X1 U15083 ( .C1(n13127), .C2(n13053), .A(n12957), .B(n12956), .ZN(
        P2_U3242) );
  AOI211_X1 U15084 ( .C1(n12963), .C2(n12959), .A(n13029), .B(n12958), .ZN(
        n12961) );
  NOR2_X1 U15085 ( .A1(n12961), .A2(n12960), .ZN(n13133) );
  OAI21_X1 U15086 ( .B1(n12964), .B2(n12963), .A(n12962), .ZN(n12965) );
  INV_X1 U15087 ( .A(n12965), .ZN(n13131) );
  OAI211_X1 U15088 ( .C1(n12967), .C2(n13129), .A(n6438), .B(n12966), .ZN(
        n13128) );
  NOR2_X1 U15089 ( .A1(n13128), .A2(n12984), .ZN(n12971) );
  AOI22_X1 U15090 ( .A1(n13078), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n12968), 
        .B2(n13081), .ZN(n12969) );
  OAI21_X1 U15091 ( .B1(n13129), .B2(n13073), .A(n12969), .ZN(n12970) );
  AOI211_X1 U15092 ( .C1(n13131), .C2(n12988), .A(n12971), .B(n12970), .ZN(
        n12972) );
  OAI21_X1 U15093 ( .B1(n13133), .B2(n13078), .A(n12972), .ZN(P2_U3243) );
  OAI21_X1 U15094 ( .B1(n12974), .B2(n12986), .A(n12973), .ZN(n12977) );
  AOI222_X1 U15095 ( .A1(n13065), .A2(n12977), .B1(n12976), .B2(n13002), .C1(
        n12975), .C2(n13004), .ZN(n13140) );
  NAND2_X1 U15096 ( .A1(n13134), .A2(n12993), .ZN(n12978) );
  NAND3_X1 U15097 ( .A1(n12979), .A2(n6438), .A3(n12978), .ZN(n13137) );
  INV_X1 U15098 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n12981) );
  OAI22_X1 U15099 ( .A1(n13038), .A2(n12981), .B1(n12980), .B2(n12998), .ZN(
        n12982) );
  AOI21_X1 U15100 ( .B1(n13134), .B2(n13082), .A(n12982), .ZN(n12983) );
  OAI21_X1 U15101 ( .B1(n13137), .B2(n12984), .A(n12983), .ZN(n12985) );
  INV_X1 U15102 ( .A(n12985), .ZN(n12990) );
  NAND2_X1 U15103 ( .A1(n12987), .A2(n12986), .ZN(n13135) );
  NAND3_X1 U15104 ( .A1(n13136), .A2(n13135), .A3(n12988), .ZN(n12989) );
  OAI211_X1 U15105 ( .C1(n13140), .C2(n13078), .A(n12990), .B(n12989), .ZN(
        P2_U3244) );
  XNOR2_X1 U15106 ( .A(n12992), .B(n12991), .ZN(n13145) );
  AOI21_X1 U15107 ( .B1(n13142), .B2(n13016), .A(n10022), .ZN(n12994) );
  AND2_X1 U15108 ( .A1(n12994), .A2(n12993), .ZN(n13141) );
  NAND2_X1 U15109 ( .A1(n13142), .A2(n13082), .ZN(n12996) );
  NAND2_X1 U15110 ( .A1(n13078), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n12995) );
  OAI211_X1 U15111 ( .C1(n12998), .C2(n12997), .A(n12996), .B(n12995), .ZN(
        n13008) );
  OAI21_X1 U15112 ( .B1(n13001), .B2(n13000), .A(n12999), .ZN(n13006) );
  AOI222_X1 U15113 ( .A1(n13065), .A2(n13006), .B1(n13005), .B2(n13004), .C1(
        n13003), .C2(n13002), .ZN(n13144) );
  NOR2_X1 U15114 ( .A1(n13144), .A2(n13078), .ZN(n13007) );
  AOI211_X1 U15115 ( .C1(n13141), .C2(n13085), .A(n13008), .B(n13007), .ZN(
        n13009) );
  OAI21_X1 U15116 ( .B1(n13053), .B2(n13145), .A(n13009), .ZN(P2_U3245) );
  XOR2_X1 U15117 ( .A(n13010), .B(n13011), .Z(n13150) );
  XNOR2_X1 U15118 ( .A(n13012), .B(n13011), .ZN(n13013) );
  OAI222_X1 U15119 ( .A1(n13057), .A2(n13015), .B1(n13055), .B2(n13014), .C1(
        n13029), .C2(n13013), .ZN(n13146) );
  INV_X1 U15120 ( .A(n13031), .ZN(n13018) );
  INV_X1 U15121 ( .A(n13016), .ZN(n13017) );
  AOI211_X1 U15122 ( .C1(n13148), .C2(n13018), .A(n10022), .B(n13017), .ZN(
        n13147) );
  NAND2_X1 U15123 ( .A1(n13147), .A2(n13085), .ZN(n13021) );
  AOI22_X1 U15124 ( .A1(n13078), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13019), 
        .B2(n13081), .ZN(n13020) );
  OAI211_X1 U15125 ( .C1(n13022), .C2(n13073), .A(n13021), .B(n13020), .ZN(
        n13023) );
  AOI21_X1 U15126 ( .B1(n13146), .B2(n13038), .A(n13023), .ZN(n13024) );
  OAI21_X1 U15127 ( .B1(n13053), .B2(n13150), .A(n13024), .ZN(P2_U3246) );
  XOR2_X1 U15128 ( .A(n13025), .B(n13026), .Z(n13155) );
  XNOR2_X1 U15129 ( .A(n13027), .B(n13026), .ZN(n13030) );
  OAI21_X1 U15130 ( .B1(n13030), .B2(n13029), .A(n13028), .ZN(n13151) );
  INV_X1 U15131 ( .A(n13041), .ZN(n13032) );
  AOI211_X1 U15132 ( .C1(n13153), .C2(n13032), .A(n10022), .B(n13031), .ZN(
        n13152) );
  NAND2_X1 U15133 ( .A1(n13152), .A2(n13085), .ZN(n13035) );
  AOI22_X1 U15134 ( .A1(n13078), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13033), 
        .B2(n13081), .ZN(n13034) );
  OAI211_X1 U15135 ( .C1(n13036), .C2(n13073), .A(n13035), .B(n13034), .ZN(
        n13037) );
  AOI21_X1 U15136 ( .B1(n13151), .B2(n13038), .A(n13037), .ZN(n13039) );
  OAI21_X1 U15137 ( .B1(n13053), .B2(n13155), .A(n13039), .ZN(P2_U3247) );
  XOR2_X1 U15138 ( .A(n13040), .B(n13046), .Z(n13160) );
  AOI211_X1 U15139 ( .C1(n13157), .C2(n13067), .A(n10022), .B(n13041), .ZN(
        n13156) );
  INV_X1 U15140 ( .A(n13042), .ZN(n13043) );
  AOI22_X1 U15141 ( .A1(n13078), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13043), 
        .B2(n13081), .ZN(n13044) );
  OAI21_X1 U15142 ( .B1(n13045), .B2(n13073), .A(n13044), .ZN(n13051) );
  XNOR2_X1 U15143 ( .A(n13047), .B(n13046), .ZN(n13049) );
  AOI21_X1 U15144 ( .B1(n13049), .B2(n13065), .A(n13048), .ZN(n13159) );
  NOR2_X1 U15145 ( .A1(n13159), .A2(n13078), .ZN(n13050) );
  AOI211_X1 U15146 ( .C1(n13156), .C2(n13085), .A(n13051), .B(n13050), .ZN(
        n13052) );
  OAI21_X1 U15147 ( .B1(n13160), .B2(n13053), .A(n13052), .ZN(P2_U3248) );
  XNOR2_X1 U15148 ( .A(n13054), .B(n13059), .ZN(n13066) );
  OAI22_X1 U15149 ( .A1(n13058), .A2(n13057), .B1(n13056), .B2(n13055), .ZN(
        n13064) );
  NAND2_X1 U15150 ( .A1(n13060), .A2(n13059), .ZN(n13061) );
  NAND2_X1 U15151 ( .A1(n13062), .A2(n13061), .ZN(n13165) );
  NOR2_X1 U15152 ( .A1(n13165), .A2(n14689), .ZN(n13063) );
  AOI211_X1 U15153 ( .C1(n13066), .C2(n13065), .A(n13064), .B(n13063), .ZN(
        n13164) );
  INV_X1 U15154 ( .A(n13067), .ZN(n13068) );
  AOI211_X1 U15155 ( .C1(n13162), .C2(n13069), .A(n10022), .B(n13068), .ZN(
        n13161) );
  INV_X1 U15156 ( .A(n13070), .ZN(n13071) );
  AOI22_X1 U15157 ( .A1(n13078), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n13071), 
        .B2(n13081), .ZN(n13072) );
  OAI21_X1 U15158 ( .B1(n13074), .B2(n13073), .A(n13072), .ZN(n13076) );
  NOR2_X1 U15159 ( .A1(n13165), .A2(n13083), .ZN(n13075) );
  AOI211_X1 U15160 ( .C1(n13161), .C2(n13085), .A(n13076), .B(n13075), .ZN(
        n13077) );
  OAI21_X1 U15161 ( .B1(n13164), .B2(n13078), .A(n13077), .ZN(P2_U3249) );
  MUX2_X1 U15162 ( .A(n13080), .B(n13079), .S(n13038), .Z(n13090) );
  AOI22_X1 U15163 ( .A1(n13082), .A2(n10021), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n13081), .ZN(n13089) );
  INV_X1 U15164 ( .A(n13083), .ZN(n13087) );
  AOI22_X1 U15165 ( .A1(n13087), .A2(n13086), .B1(n13085), .B2(n13084), .ZN(
        n13088) );
  NAND3_X1 U15166 ( .A1(n13090), .A2(n13089), .A3(n13088), .ZN(P2_U3264) );
  MUX2_X1 U15167 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13171), .S(n14737), .Z(
        P2_U3530) );
  OAI211_X1 U15168 ( .C1(n13094), .C2(n14715), .A(n13093), .B(n13092), .ZN(
        n13172) );
  MUX2_X1 U15169 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13172), .S(n14737), .Z(
        P2_U3529) );
  AOI21_X1 U15170 ( .B1(n14660), .B2(n13096), .A(n13095), .ZN(n13097) );
  MUX2_X1 U15171 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13173), .S(n14737), .Z(
        P2_U3527) );
  AOI21_X1 U15172 ( .B1(n14660), .B2(n13103), .A(n13102), .ZN(n13104) );
  OAI211_X1 U15173 ( .C1(n14655), .C2(n13106), .A(n13105), .B(n13104), .ZN(
        n13174) );
  MUX2_X1 U15174 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13174), .S(n14737), .Z(
        P2_U3526) );
  AOI21_X1 U15175 ( .B1(n14660), .B2(n13108), .A(n13107), .ZN(n13109) );
  OAI211_X1 U15176 ( .C1(n14655), .C2(n13111), .A(n13110), .B(n13109), .ZN(
        n13175) );
  MUX2_X1 U15177 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13175), .S(n14737), .Z(
        P2_U3525) );
  AOI21_X1 U15178 ( .B1(n14660), .B2(n13113), .A(n13112), .ZN(n13114) );
  OAI211_X1 U15179 ( .C1(n14655), .C2(n13116), .A(n13115), .B(n13114), .ZN(
        n13176) );
  MUX2_X1 U15180 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13176), .S(n14737), .Z(
        P2_U3524) );
  AOI21_X1 U15181 ( .B1(n14660), .B2(n13118), .A(n13117), .ZN(n13119) );
  OAI211_X1 U15182 ( .C1(n14655), .C2(n13121), .A(n13120), .B(n13119), .ZN(
        n13177) );
  MUX2_X1 U15183 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13177), .S(n14737), .Z(
        P2_U3523) );
  AOI211_X1 U15184 ( .C1(n14660), .C2(n13124), .A(n13123), .B(n13122), .ZN(
        n13125) );
  OAI211_X1 U15185 ( .C1(n14655), .C2(n13127), .A(n13126), .B(n13125), .ZN(
        n13178) );
  MUX2_X1 U15186 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13178), .S(n14737), .Z(
        P2_U3522) );
  INV_X1 U15187 ( .A(n14655), .ZN(n14719) );
  OAI21_X1 U15188 ( .B1(n13129), .B2(n14715), .A(n13128), .ZN(n13130) );
  AOI21_X1 U15189 ( .B1(n13131), .B2(n14719), .A(n13130), .ZN(n13132) );
  NAND2_X1 U15190 ( .A1(n13133), .A2(n13132), .ZN(n13179) );
  MUX2_X1 U15191 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13179), .S(n14737), .Z(
        P2_U3521) );
  NAND2_X1 U15192 ( .A1(n13134), .A2(n14660), .ZN(n13139) );
  NAND3_X1 U15193 ( .A1(n13136), .A2(n13135), .A3(n14719), .ZN(n13138) );
  NAND4_X1 U15194 ( .A1(n13140), .A2(n13139), .A3(n13138), .A4(n13137), .ZN(
        n13180) );
  MUX2_X1 U15195 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13180), .S(n14737), .Z(
        P2_U3520) );
  AOI21_X1 U15196 ( .B1(n14660), .B2(n13142), .A(n13141), .ZN(n13143) );
  OAI211_X1 U15197 ( .C1(n14655), .C2(n13145), .A(n13144), .B(n13143), .ZN(
        n13181) );
  MUX2_X1 U15198 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13181), .S(n14737), .Z(
        P2_U3519) );
  AOI211_X1 U15199 ( .C1(n14660), .C2(n13148), .A(n13147), .B(n13146), .ZN(
        n13149) );
  OAI21_X1 U15200 ( .B1(n14655), .B2(n13150), .A(n13149), .ZN(n13182) );
  MUX2_X1 U15201 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13182), .S(n14737), .Z(
        P2_U3518) );
  AOI211_X1 U15202 ( .C1(n14660), .C2(n13153), .A(n13152), .B(n13151), .ZN(
        n13154) );
  OAI21_X1 U15203 ( .B1(n14655), .B2(n13155), .A(n13154), .ZN(n13183) );
  MUX2_X1 U15204 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13183), .S(n14737), .Z(
        P2_U3517) );
  AOI21_X1 U15205 ( .B1(n14660), .B2(n13157), .A(n13156), .ZN(n13158) );
  OAI211_X1 U15206 ( .C1(n14655), .C2(n13160), .A(n13159), .B(n13158), .ZN(
        n13184) );
  MUX2_X1 U15207 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13184), .S(n14737), .Z(
        P2_U3516) );
  AOI21_X1 U15208 ( .B1(n14660), .B2(n13162), .A(n13161), .ZN(n13163) );
  OAI211_X1 U15209 ( .C1(n14688), .C2(n13165), .A(n13164), .B(n13163), .ZN(
        n13185) );
  MUX2_X1 U15210 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13185), .S(n14737), .Z(
        P2_U3515) );
  AOI21_X1 U15211 ( .B1(n14660), .B2(n13167), .A(n13166), .ZN(n13168) );
  OAI211_X1 U15212 ( .C1(n13170), .C2(n14655), .A(n13169), .B(n13168), .ZN(
        n13186) );
  MUX2_X1 U15213 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13186), .S(n14737), .Z(
        P2_U3514) );
  MUX2_X1 U15214 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13171), .S(n14723), .Z(
        P2_U3498) );
  MUX2_X1 U15215 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13172), .S(n14723), .Z(
        P2_U3497) );
  MUX2_X1 U15216 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13173), .S(n14723), .Z(
        P2_U3495) );
  MUX2_X1 U15217 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13174), .S(n14723), .Z(
        P2_U3494) );
  MUX2_X1 U15218 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13175), .S(n14723), .Z(
        P2_U3493) );
  MUX2_X1 U15219 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13176), .S(n14723), .Z(
        P2_U3492) );
  MUX2_X1 U15220 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13177), .S(n14723), .Z(
        P2_U3491) );
  MUX2_X1 U15221 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13178), .S(n14723), .Z(
        P2_U3490) );
  MUX2_X1 U15222 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13179), .S(n14723), .Z(
        P2_U3489) );
  MUX2_X1 U15223 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13180), .S(n14723), .Z(
        P2_U3488) );
  MUX2_X1 U15224 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13181), .S(n14723), .Z(
        P2_U3487) );
  MUX2_X1 U15225 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13182), .S(n14723), .Z(
        P2_U3486) );
  MUX2_X1 U15226 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13183), .S(n14723), .Z(
        P2_U3484) );
  MUX2_X1 U15227 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13184), .S(n14723), .Z(
        P2_U3481) );
  MUX2_X1 U15228 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13185), .S(n14723), .Z(
        P2_U3478) );
  MUX2_X1 U15229 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13186), .S(n14723), .Z(
        P2_U3475) );
  INV_X1 U15230 ( .A(n13187), .ZN(n13978) );
  NOR4_X1 U15231 ( .A1(n6724), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13189), .A4(
        P2_U3088), .ZN(n13190) );
  AOI21_X1 U15232 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n13196), .A(n13190), 
        .ZN(n13191) );
  OAI21_X1 U15233 ( .B1(n13978), .B2(n13199), .A(n13191), .ZN(P2_U3296) );
  INV_X1 U15234 ( .A(n13192), .ZN(n13985) );
  NAND2_X1 U15235 ( .A1(n13196), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13193) );
  OAI211_X1 U15236 ( .C1(n13985), .C2(n13199), .A(n13194), .B(n13193), .ZN(
        P2_U3299) );
  INV_X1 U15237 ( .A(n13195), .ZN(n13990) );
  NAND2_X1 U15238 ( .A1(n13196), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13198) );
  OAI211_X1 U15239 ( .C1(n13990), .C2(n13199), .A(n13198), .B(n13197), .ZN(
        P2_U3300) );
  INV_X1 U15240 ( .A(n13200), .ZN(n13993) );
  OAI222_X1 U15241 ( .A1(n13203), .A2(P2_U3088), .B1(n13199), .B2(n13993), 
        .C1(n13202), .C2(n13201), .ZN(P2_U3301) );
  MUX2_X1 U15242 ( .A(n13204), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI22_X1 U15243 ( .A1(n13719), .A2(n13367), .B1(n13651), .B2(n13264), .ZN(
        n13205) );
  XNOR2_X1 U15244 ( .A(n13205), .B(n13365), .ZN(n13210) );
  OR2_X1 U15245 ( .A1(n13719), .A2(n13264), .ZN(n13208) );
  OR2_X1 U15246 ( .A1(n13364), .A2(n13651), .ZN(n13207) );
  NAND2_X1 U15247 ( .A1(n13208), .A2(n13207), .ZN(n13209) );
  NOR2_X1 U15248 ( .A1(n13210), .A2(n13209), .ZN(n13362) );
  AOI21_X1 U15249 ( .B1(n13210), .B2(n13209), .A(n13362), .ZN(n13337) );
  NAND2_X1 U15250 ( .A1(n13212), .A2(n13211), .ZN(n14219) );
  NAND2_X1 U15251 ( .A1(n14226), .A2(n7444), .ZN(n13214) );
  NAND2_X1 U15252 ( .A1(n13476), .A2(n6443), .ZN(n13213) );
  NAND2_X1 U15253 ( .A1(n13214), .A2(n13213), .ZN(n13215) );
  XNOR2_X1 U15254 ( .A(n13215), .B(n13365), .ZN(n13220) );
  AND2_X1 U15255 ( .A1(n13331), .A2(n13476), .ZN(n13216) );
  AOI21_X1 U15256 ( .B1(n14226), .B2(n6443), .A(n13216), .ZN(n13218) );
  XNOR2_X1 U15257 ( .A(n13220), .B(n13218), .ZN(n14217) );
  INV_X1 U15258 ( .A(n13218), .ZN(n13219) );
  AND2_X1 U15259 ( .A1(n13331), .A2(n13475), .ZN(n13222) );
  AOI21_X1 U15260 ( .B1(n14120), .B2(n6443), .A(n13222), .ZN(n13227) );
  NAND2_X1 U15261 ( .A1(n14120), .A2(n7444), .ZN(n13224) );
  NAND2_X1 U15262 ( .A1(n13475), .A2(n6443), .ZN(n13223) );
  NAND2_X1 U15263 ( .A1(n13224), .A2(n13223), .ZN(n13225) );
  XNOR2_X1 U15264 ( .A(n13225), .B(n13365), .ZN(n13229) );
  XOR2_X1 U15265 ( .A(n13227), .B(n13229), .Z(n13386) );
  INV_X1 U15266 ( .A(n13386), .ZN(n13226) );
  INV_X1 U15267 ( .A(n13227), .ZN(n13228) );
  NAND2_X1 U15268 ( .A1(n13229), .A2(n13228), .ZN(n13230) );
  AND2_X1 U15269 ( .A1(n13331), .A2(n13474), .ZN(n13231) );
  AOI21_X1 U15270 ( .B1(n13433), .B2(n6443), .A(n13231), .ZN(n13238) );
  AOI22_X1 U15271 ( .A1(n13433), .A2(n7444), .B1(n6443), .B2(n13474), .ZN(
        n13232) );
  XNOR2_X1 U15272 ( .A(n13232), .B(n13365), .ZN(n13239) );
  XOR2_X1 U15273 ( .A(n13238), .B(n13239), .Z(n13435) );
  NAND2_X1 U15274 ( .A1(n14285), .A2(n7444), .ZN(n13234) );
  OR2_X1 U15275 ( .A1(n13236), .A2(n13264), .ZN(n13233) );
  NAND2_X1 U15276 ( .A1(n13234), .A2(n13233), .ZN(n13235) );
  XNOR2_X1 U15277 ( .A(n13235), .B(n13318), .ZN(n13242) );
  NOR2_X1 U15278 ( .A1(n13236), .A2(n13364), .ZN(n13237) );
  AOI21_X1 U15279 ( .B1(n14285), .B2(n6443), .A(n13237), .ZN(n13241) );
  XNOR2_X1 U15280 ( .A(n13242), .B(n13241), .ZN(n14196) );
  NOR2_X1 U15281 ( .A1(n13239), .A2(n13238), .ZN(n14197) );
  NOR2_X1 U15282 ( .A1(n14196), .A2(n14197), .ZN(n13240) );
  NAND2_X1 U15283 ( .A1(n13242), .A2(n13241), .ZN(n13243) );
  NAND2_X1 U15284 ( .A1(n14237), .A2(n7444), .ZN(n13245) );
  OR2_X1 U15285 ( .A1(n14208), .A2(n13264), .ZN(n13244) );
  NAND2_X1 U15286 ( .A1(n13245), .A2(n13244), .ZN(n13246) );
  XNOR2_X1 U15287 ( .A(n13246), .B(n13365), .ZN(n13247) );
  INV_X1 U15288 ( .A(n14208), .ZN(n13628) );
  AOI22_X1 U15289 ( .A1(n14237), .A2(n6443), .B1(n13331), .B2(n13628), .ZN(
        n14232) );
  INV_X1 U15290 ( .A(n13247), .ZN(n13248) );
  NAND2_X1 U15291 ( .A1(n13249), .A2(n13248), .ZN(n13250) );
  NAND2_X1 U15292 ( .A1(n14271), .A2(n7444), .ZN(n13252) );
  NAND2_X1 U15293 ( .A1(n13866), .A2(n6443), .ZN(n13251) );
  NAND2_X1 U15294 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  XNOR2_X1 U15295 ( .A(n13253), .B(n13365), .ZN(n13254) );
  AOI22_X1 U15296 ( .A1(n14271), .A2(n6443), .B1(n13331), .B2(n13866), .ZN(
        n13255) );
  XNOR2_X1 U15297 ( .A(n13254), .B(n13255), .ZN(n14207) );
  INV_X1 U15298 ( .A(n13254), .ZN(n13256) );
  NAND2_X1 U15299 ( .A1(n13256), .A2(n13255), .ZN(n13257) );
  OAI22_X1 U15300 ( .A1(n14265), .A2(n13367), .B1(n14209), .B2(n13264), .ZN(
        n13259) );
  XNOR2_X1 U15301 ( .A(n13259), .B(n13365), .ZN(n13407) );
  OR2_X1 U15302 ( .A1(n14265), .A2(n13264), .ZN(n13261) );
  NAND2_X1 U15303 ( .A1(n13658), .A2(n13331), .ZN(n13260) );
  NAND2_X1 U15304 ( .A1(n13261), .A2(n13260), .ZN(n13406) );
  NOR2_X1 U15305 ( .A1(n13407), .A2(n13406), .ZN(n13263) );
  NAND2_X1 U15306 ( .A1(n13407), .A2(n13406), .ZN(n13262) );
  OAI22_X1 U15307 ( .A1(n14257), .A2(n13367), .B1(n13864), .B2(n13264), .ZN(
        n13265) );
  XNOR2_X1 U15308 ( .A(n13265), .B(n13365), .ZN(n13271) );
  OAI22_X1 U15309 ( .A1(n14257), .A2(n13264), .B1(n13864), .B2(n13364), .ZN(
        n13270) );
  XNOR2_X1 U15310 ( .A(n13271), .B(n13270), .ZN(n13452) );
  NAND2_X1 U15311 ( .A1(n11568), .A2(n7444), .ZN(n13267) );
  INV_X1 U15312 ( .A(n13848), .ZN(n13637) );
  NAND2_X1 U15313 ( .A1(n13637), .A2(n6443), .ZN(n13266) );
  NAND2_X1 U15314 ( .A1(n13267), .A2(n13266), .ZN(n13268) );
  XNOR2_X1 U15315 ( .A(n13268), .B(n13318), .ZN(n13274) );
  NOR2_X1 U15316 ( .A1(n13848), .A2(n13364), .ZN(n13269) );
  AOI21_X1 U15317 ( .B1(n11568), .B2(n6443), .A(n13269), .ZN(n13273) );
  XNOR2_X1 U15318 ( .A(n13274), .B(n13273), .ZN(n13354) );
  NOR2_X1 U15319 ( .A1(n13271), .A2(n13270), .ZN(n13355) );
  NOR2_X1 U15320 ( .A1(n13354), .A2(n13355), .ZN(n13272) );
  NAND2_X1 U15321 ( .A1(n13950), .A2(n7444), .ZN(n13276) );
  NAND2_X1 U15322 ( .A1(n13836), .A2(n6443), .ZN(n13275) );
  NAND2_X1 U15323 ( .A1(n13276), .A2(n13275), .ZN(n13277) );
  XNOR2_X1 U15324 ( .A(n13277), .B(n13365), .ZN(n13280) );
  AOI22_X1 U15325 ( .A1(n13950), .A2(n6443), .B1(n13331), .B2(n13836), .ZN(
        n13278) );
  XNOR2_X1 U15326 ( .A(n13280), .B(n13278), .ZN(n13427) );
  INV_X1 U15327 ( .A(n13278), .ZN(n13279) );
  NAND2_X1 U15328 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  NAND2_X1 U15329 ( .A1(n13945), .A2(n7444), .ZN(n13284) );
  NAND2_X1 U15330 ( .A1(n13641), .A2(n6443), .ZN(n13283) );
  NAND2_X1 U15331 ( .A1(n13284), .A2(n13283), .ZN(n13285) );
  XNOR2_X1 U15332 ( .A(n13285), .B(n13318), .ZN(n13288) );
  AND2_X1 U15333 ( .A1(n13641), .A2(n13331), .ZN(n13286) );
  AOI21_X1 U15334 ( .B1(n13945), .B2(n6443), .A(n13286), .ZN(n13287) );
  NAND2_X1 U15335 ( .A1(n13288), .A2(n13287), .ZN(n13441) );
  OAI21_X1 U15336 ( .B1(n13288), .B2(n13287), .A(n13441), .ZN(n13378) );
  NAND2_X1 U15337 ( .A1(n13793), .A2(n7444), .ZN(n13290) );
  NAND2_X1 U15338 ( .A1(n13666), .A2(n6443), .ZN(n13289) );
  NAND2_X1 U15339 ( .A1(n13290), .A2(n13289), .ZN(n13291) );
  XNOR2_X1 U15340 ( .A(n13291), .B(n13318), .ZN(n13293) );
  AND2_X1 U15341 ( .A1(n13666), .A2(n13331), .ZN(n13292) );
  AOI21_X1 U15342 ( .B1(n13793), .B2(n6443), .A(n13292), .ZN(n13294) );
  NAND2_X1 U15343 ( .A1(n13293), .A2(n13294), .ZN(n13344) );
  INV_X1 U15344 ( .A(n13293), .ZN(n13296) );
  INV_X1 U15345 ( .A(n13294), .ZN(n13295) );
  NAND2_X1 U15346 ( .A1(n13296), .A2(n13295), .ZN(n13297) );
  NAND2_X1 U15347 ( .A1(n13780), .A2(n7444), .ZN(n13299) );
  NAND2_X1 U15348 ( .A1(n13667), .A2(n6443), .ZN(n13298) );
  NAND2_X1 U15349 ( .A1(n13299), .A2(n13298), .ZN(n13300) );
  XNOR2_X1 U15350 ( .A(n13300), .B(n13318), .ZN(n13302) );
  AND2_X1 U15351 ( .A1(n13667), .A2(n13331), .ZN(n13301) );
  AOI21_X1 U15352 ( .B1(n13780), .B2(n6443), .A(n13301), .ZN(n13303) );
  NAND2_X1 U15353 ( .A1(n13302), .A2(n13303), .ZN(n13416) );
  INV_X1 U15354 ( .A(n13302), .ZN(n13305) );
  INV_X1 U15355 ( .A(n13303), .ZN(n13304) );
  NAND2_X1 U15356 ( .A1(n13305), .A2(n13304), .ZN(n13306) );
  NAND2_X1 U15357 ( .A1(n13926), .A2(n7444), .ZN(n13308) );
  NAND2_X1 U15358 ( .A1(n13645), .A2(n6443), .ZN(n13307) );
  NAND2_X1 U15359 ( .A1(n13308), .A2(n13307), .ZN(n13309) );
  XNOR2_X1 U15360 ( .A(n13309), .B(n13318), .ZN(n13311) );
  AND2_X1 U15361 ( .A1(n13331), .A2(n13645), .ZN(n13310) );
  AOI21_X1 U15362 ( .B1(n13926), .B2(n6443), .A(n13310), .ZN(n13312) );
  NAND2_X1 U15363 ( .A1(n13311), .A2(n13312), .ZN(n13396) );
  INV_X1 U15364 ( .A(n13311), .ZN(n13314) );
  INV_X1 U15365 ( .A(n13312), .ZN(n13313) );
  NAND2_X1 U15366 ( .A1(n13314), .A2(n13313), .ZN(n13315) );
  NAND2_X1 U15367 ( .A1(n13395), .A2(n13396), .ZN(n13326) );
  NAND2_X1 U15368 ( .A1(n13919), .A2(n7444), .ZN(n13317) );
  NAND2_X1 U15369 ( .A1(n13654), .A2(n6443), .ZN(n13316) );
  NAND2_X1 U15370 ( .A1(n13317), .A2(n13316), .ZN(n13319) );
  XNOR2_X1 U15371 ( .A(n13319), .B(n13318), .ZN(n13321) );
  AND2_X1 U15372 ( .A1(n13331), .A2(n13654), .ZN(n13320) );
  AOI21_X1 U15373 ( .B1(n13919), .B2(n6443), .A(n13320), .ZN(n13322) );
  INV_X1 U15374 ( .A(n13321), .ZN(n13324) );
  INV_X1 U15375 ( .A(n13322), .ZN(n13323) );
  NAND2_X1 U15376 ( .A1(n13324), .A2(n13323), .ZN(n13325) );
  NAND2_X1 U15377 ( .A1(n13648), .A2(n7444), .ZN(n13329) );
  NAND2_X1 U15378 ( .A1(n13671), .A2(n6443), .ZN(n13328) );
  NAND2_X1 U15379 ( .A1(n13329), .A2(n13328), .ZN(n13330) );
  XNOR2_X1 U15380 ( .A(n13330), .B(n13365), .ZN(n13335) );
  NAND2_X1 U15381 ( .A1(n13648), .A2(n6443), .ZN(n13333) );
  NAND2_X1 U15382 ( .A1(n13331), .A2(n13671), .ZN(n13332) );
  NAND2_X1 U15383 ( .A1(n13333), .A2(n13332), .ZN(n13334) );
  AOI21_X1 U15384 ( .B1(n13335), .B2(n13334), .A(n13336), .ZN(n13460) );
  OR2_X1 U15385 ( .A1(n13675), .A2(n14380), .ZN(n13339) );
  NAND2_X1 U15386 ( .A1(n13671), .A2(n13865), .ZN(n13338) );
  NAND2_X1 U15387 ( .A1(n13339), .A2(n13338), .ZN(n13712) );
  AOI22_X1 U15388 ( .A1(n14235), .A2(n13712), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13341) );
  OR2_X1 U15389 ( .A1(n14241), .A2(n13716), .ZN(n13340) );
  OAI211_X1 U15390 ( .C1(n13719), .C2(n13469), .A(n13341), .B(n13340), .ZN(
        n13342) );
  NOR2_X1 U15391 ( .A1(n13345), .A2(n6632), .ZN(n13348) );
  AOI21_X1 U15392 ( .B1(n13348), .B2(n13347), .A(n6487), .ZN(n13353) );
  AND2_X1 U15393 ( .A1(n13645), .A2(n13835), .ZN(n13349) );
  AOI21_X1 U15394 ( .B1(n13666), .B2(n13865), .A(n13349), .ZN(n13929) );
  AOI22_X1 U15395 ( .A1(n13777), .A2(n13465), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13350) );
  OAI21_X1 U15396 ( .B1(n13929), .B2(n13463), .A(n13350), .ZN(n13351) );
  AOI21_X1 U15397 ( .B1(n13780), .B2(n14238), .A(n13351), .ZN(n13352) );
  OAI21_X1 U15398 ( .B1(n13353), .B2(n14221), .A(n13352), .ZN(P1_U3216) );
  OAI21_X1 U15399 ( .B1(n6488), .B2(n13355), .A(n13354), .ZN(n13357) );
  NAND3_X1 U15400 ( .A1(n13357), .A2(n14233), .A3(n13356), .ZN(n13361) );
  INV_X1 U15401 ( .A(n14215), .ZN(n13359) );
  AND2_X1 U15402 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13612) );
  OAI22_X1 U15403 ( .A1(n14214), .A2(n13864), .B1(n14241), .B2(n13837), .ZN(
        n13358) );
  AOI211_X1 U15404 ( .C1(n13359), .C2(n13836), .A(n13612), .B(n13358), .ZN(
        n13360) );
  OAI211_X1 U15405 ( .C1(n6940), .C2(n13469), .A(n13361), .B(n13360), .ZN(
        P1_U3219) );
  OAI22_X1 U15406 ( .A1(n13700), .A2(n13264), .B1(n13675), .B2(n13364), .ZN(
        n13366) );
  XNOR2_X1 U15407 ( .A(n13366), .B(n13365), .ZN(n13369) );
  OAI22_X1 U15408 ( .A1(n13700), .A2(n13367), .B1(n13675), .B2(n13264), .ZN(
        n13368) );
  XNOR2_X1 U15409 ( .A(n13371), .B(n13370), .ZN(n13377) );
  OAI22_X1 U15410 ( .A1(n14214), .A2(n13651), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13372), .ZN(n13375) );
  INV_X1 U15411 ( .A(n13693), .ZN(n13373) );
  OAI22_X1 U15412 ( .A1(n14215), .A2(n13373), .B1(n14241), .B2(n13697), .ZN(
        n13374) );
  AOI211_X1 U15413 ( .C1(n13898), .C2(n14238), .A(n13375), .B(n13374), .ZN(
        n13376) );
  OAI21_X1 U15414 ( .B1(n13377), .B2(n14221), .A(n13376), .ZN(P1_U3220) );
  AOI21_X1 U15415 ( .B1(n13379), .B2(n13378), .A(n6454), .ZN(n13385) );
  INV_X1 U15416 ( .A(n13666), .ZN(n13381) );
  INV_X1 U15417 ( .A(n13836), .ZN(n13380) );
  OAI22_X1 U15418 ( .A1(n13381), .A2(n14380), .B1(n13380), .B2(n14382), .ZN(
        n13799) );
  AOI22_X1 U15419 ( .A1(n13799), .A2(n14235), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13382) );
  OAI21_X1 U15420 ( .B1(n14241), .B2(n13803), .A(n13382), .ZN(n13383) );
  AOI21_X1 U15421 ( .B1(n13945), .B2(n14238), .A(n13383), .ZN(n13384) );
  OAI21_X1 U15422 ( .B1(n13385), .B2(n14221), .A(n13384), .ZN(P1_U3223) );
  AOI21_X1 U15423 ( .B1(n13387), .B2(n13386), .A(n14221), .ZN(n13389) );
  NAND2_X1 U15424 ( .A1(n13389), .A2(n13388), .ZN(n13394) );
  INV_X1 U15425 ( .A(n13390), .ZN(n14119) );
  AOI22_X1 U15426 ( .A1(n13865), .A2(n13476), .B1(n13474), .B2(n13835), .ZN(
        n14116) );
  OAI22_X1 U15427 ( .A1(n14116), .A2(n13463), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13391), .ZN(n13392) );
  AOI21_X1 U15428 ( .B1(n14119), .B2(n13465), .A(n13392), .ZN(n13393) );
  OAI211_X1 U15429 ( .C1(n6936), .C2(n13469), .A(n13394), .B(n13393), .ZN(
        P1_U3224) );
  INV_X1 U15430 ( .A(n13395), .ZN(n13418) );
  INV_X1 U15431 ( .A(n13396), .ZN(n13398) );
  NOR3_X1 U15432 ( .A1(n13418), .A2(n13398), .A3(n13397), .ZN(n13401) );
  INV_X1 U15433 ( .A(n13399), .ZN(n13400) );
  OAI21_X1 U15434 ( .B1(n13401), .B2(n13400), .A(n14233), .ZN(n13405) );
  INV_X1 U15435 ( .A(n13671), .ZN(n13740) );
  NOR2_X1 U15436 ( .A1(n14215), .A2(n13740), .ZN(n13403) );
  OAI22_X1 U15437 ( .A1(n14241), .A2(n13743), .B1(n14214), .B2(n13739), .ZN(
        n13402) );
  AOI211_X1 U15438 ( .C1(P1_REG3_REG_25__SCAN_IN), .C2(P1_U3086), .A(n13403), 
        .B(n13402), .ZN(n13404) );
  OAI211_X1 U15439 ( .C1(n6945), .C2(n13469), .A(n13405), .B(n13404), .ZN(
        P1_U3225) );
  XNOR2_X1 U15440 ( .A(n13407), .B(n13406), .ZN(n13408) );
  XNOR2_X1 U15441 ( .A(n13409), .B(n13408), .ZN(n13415) );
  OAI21_X1 U15442 ( .B1(n14214), .B2(n13411), .A(n13410), .ZN(n13413) );
  OAI22_X1 U15443 ( .A1(n14215), .A2(n13864), .B1(n14241), .B2(n13863), .ZN(
        n13412) );
  AOI211_X1 U15444 ( .C1(n13659), .C2(n14238), .A(n13413), .B(n13412), .ZN(
        n13414) );
  OAI21_X1 U15445 ( .B1(n13415), .B2(n14221), .A(n13414), .ZN(P1_U3228) );
  NOR3_X1 U15446 ( .A1(n6487), .A2(n6631), .A3(n13417), .ZN(n13419) );
  OAI21_X1 U15447 ( .B1(n13419), .B2(n13418), .A(n14233), .ZN(n13425) );
  NAND2_X1 U15448 ( .A1(n13667), .A2(n13865), .ZN(n13421) );
  NAND2_X1 U15449 ( .A1(n13654), .A2(n13835), .ZN(n13420) );
  NAND2_X1 U15450 ( .A1(n13421), .A2(n13420), .ZN(n13758) );
  INV_X1 U15451 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13422) );
  OAI22_X1 U15452 ( .A1(n14241), .A2(n13764), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13422), .ZN(n13423) );
  AOI21_X1 U15453 ( .B1(n13758), .B2(n14235), .A(n13423), .ZN(n13424) );
  OAI211_X1 U15454 ( .C1(n6946), .C2(n13469), .A(n13425), .B(n13424), .ZN(
        P1_U3229) );
  XNOR2_X1 U15455 ( .A(n13426), .B(n13427), .ZN(n13432) );
  OAI22_X1 U15456 ( .A1(n13817), .A2(n14215), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13428), .ZN(n13430) );
  OAI22_X1 U15457 ( .A1(n14214), .A2(n13848), .B1(n14241), .B2(n13824), .ZN(
        n13429) );
  AOI211_X1 U15458 ( .C1(n13950), .C2(n14238), .A(n13430), .B(n13429), .ZN(
        n13431) );
  OAI21_X1 U15459 ( .B1(n13432), .B2(n14221), .A(n13431), .ZN(P1_U3233) );
  OAI211_X1 U15460 ( .C1(n13435), .C2(n13434), .A(n14195), .B(n14233), .ZN(
        n13440) );
  OAI21_X1 U15461 ( .B1(n14292), .B2(n13463), .A(n13436), .ZN(n13437) );
  AOI21_X1 U15462 ( .B1(n13438), .B2(n13465), .A(n13437), .ZN(n13439) );
  OAI211_X1 U15463 ( .C1(n6934), .C2(n13469), .A(n13440), .B(n13439), .ZN(
        P1_U3234) );
  NOR3_X1 U15464 ( .A1(n6454), .A2(n7475), .A3(n13442), .ZN(n13444) );
  INV_X1 U15465 ( .A(n13347), .ZN(n13443) );
  OAI21_X1 U15466 ( .B1(n13444), .B2(n13443), .A(n14233), .ZN(n13450) );
  NAND2_X1 U15467 ( .A1(n13667), .A2(n13835), .ZN(n13446) );
  NAND2_X1 U15468 ( .A1(n13641), .A2(n13865), .ZN(n13445) );
  NAND2_X1 U15469 ( .A1(n13446), .A2(n13445), .ZN(n13936) );
  INV_X1 U15470 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13447) );
  OAI22_X1 U15471 ( .A1(n13791), .A2(n14241), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13447), .ZN(n13448) );
  AOI21_X1 U15472 ( .B1(n13936), .B2(n14235), .A(n13448), .ZN(n13449) );
  OAI211_X1 U15473 ( .C1(n13469), .C2(n13939), .A(n13450), .B(n13449), .ZN(
        P1_U3235) );
  AOI21_X1 U15474 ( .B1(n13452), .B2(n13451), .A(n6488), .ZN(n13457) );
  AOI22_X1 U15475 ( .A1(n13453), .A2(n13658), .B1(n13465), .B2(n13852), .ZN(
        n13454) );
  NAND2_X1 U15476 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14377)
         );
  OAI211_X1 U15477 ( .C1(n13848), .C2(n14215), .A(n13454), .B(n14377), .ZN(
        n13455) );
  AOI21_X1 U15478 ( .B1(n13860), .B2(n14238), .A(n13455), .ZN(n13456) );
  OAI21_X1 U15479 ( .B1(n13457), .B2(n14221), .A(n13456), .ZN(P1_U3238) );
  OAI21_X1 U15480 ( .B1(n13460), .B2(n13459), .A(n13458), .ZN(n13461) );
  NAND2_X1 U15481 ( .A1(n13461), .A2(n14233), .ZN(n13468) );
  INV_X1 U15482 ( .A(n13730), .ZN(n13466) );
  INV_X1 U15483 ( .A(n13651), .ZN(n13694) );
  AOI22_X1 U15484 ( .A1(n13694), .A2(n13835), .B1(n13865), .B2(n13654), .ZN(
        n13910) );
  OAI22_X1 U15485 ( .A1(n13910), .A2(n13463), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13462), .ZN(n13464) );
  AOI21_X1 U15486 ( .B1(n13466), .B2(n13465), .A(n13464), .ZN(n13467) );
  OAI211_X1 U15487 ( .C1(n13911), .C2(n13469), .A(n13468), .B(n13467), .ZN(
        P1_U3240) );
  MUX2_X1 U15488 ( .A(n13470), .B(P1_DATAO_REG_31__SCAN_IN), .S(n14991), .Z(
        P1_U3591) );
  MUX2_X1 U15489 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13471), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15490 ( .A(n13693), .B(P1_DATAO_REG_29__SCAN_IN), .S(n14991), .Z(
        P1_U3589) );
  MUX2_X1 U15491 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n13472), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15492 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n13694), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15493 ( .A(n13671), .B(P1_DATAO_REG_26__SCAN_IN), .S(n14991), .Z(
        P1_U3586) );
  MUX2_X1 U15494 ( .A(n13654), .B(P1_DATAO_REG_25__SCAN_IN), .S(n14991), .Z(
        P1_U3585) );
  MUX2_X1 U15495 ( .A(n13645), .B(P1_DATAO_REG_24__SCAN_IN), .S(n14991), .Z(
        P1_U3584) );
  MUX2_X1 U15496 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13667), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U15497 ( .A(n13666), .B(P1_DATAO_REG_22__SCAN_IN), .S(n14991), .Z(
        P1_U3582) );
  MUX2_X1 U15498 ( .A(n13641), .B(P1_DATAO_REG_21__SCAN_IN), .S(n14991), .Z(
        P1_U3581) );
  MUX2_X1 U15499 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13836), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15500 ( .A(n13637), .B(P1_DATAO_REG_19__SCAN_IN), .S(n14991), .Z(
        P1_U3579) );
  INV_X1 U15501 ( .A(n13864), .ZN(n13834) );
  MUX2_X1 U15502 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13834), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15503 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n13658), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15504 ( .A(n13866), .B(P1_DATAO_REG_16__SCAN_IN), .S(n14991), .Z(
        P1_U3576) );
  MUX2_X1 U15505 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13628), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15506 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13473), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15507 ( .A(n13474), .B(P1_DATAO_REG_13__SCAN_IN), .S(n14991), .Z(
        P1_U3573) );
  MUX2_X1 U15508 ( .A(n13475), .B(P1_DATAO_REG_12__SCAN_IN), .S(n14991), .Z(
        P1_U3572) );
  MUX2_X1 U15509 ( .A(n13476), .B(P1_DATAO_REG_11__SCAN_IN), .S(n14991), .Z(
        P1_U3571) );
  MUX2_X1 U15510 ( .A(n13477), .B(P1_DATAO_REG_10__SCAN_IN), .S(n14991), .Z(
        P1_U3570) );
  MUX2_X1 U15511 ( .A(n13478), .B(P1_DATAO_REG_9__SCAN_IN), .S(n14991), .Z(
        P1_U3569) );
  MUX2_X1 U15512 ( .A(n13479), .B(P1_DATAO_REG_8__SCAN_IN), .S(n14991), .Z(
        P1_U3568) );
  MUX2_X1 U15513 ( .A(n13480), .B(P1_DATAO_REG_7__SCAN_IN), .S(n14991), .Z(
        P1_U3567) );
  MUX2_X1 U15514 ( .A(n13481), .B(P1_DATAO_REG_6__SCAN_IN), .S(n14991), .Z(
        P1_U3566) );
  MUX2_X1 U15515 ( .A(n13482), .B(P1_DATAO_REG_5__SCAN_IN), .S(n14991), .Z(
        P1_U3565) );
  MUX2_X1 U15516 ( .A(n13483), .B(P1_DATAO_REG_4__SCAN_IN), .S(n14991), .Z(
        P1_U3564) );
  MUX2_X1 U15517 ( .A(n13484), .B(P1_DATAO_REG_2__SCAN_IN), .S(n14991), .Z(
        P1_U3562) );
  MUX2_X1 U15518 ( .A(n13485), .B(P1_DATAO_REG_1__SCAN_IN), .S(n14991), .Z(
        P1_U3561) );
  MUX2_X1 U15519 ( .A(n13486), .B(P1_DATAO_REG_0__SCAN_IN), .S(n14991), .Z(
        P1_U3560) );
  OAI211_X1 U15520 ( .C1(n13489), .C2(n13488), .A(n14367), .B(n13487), .ZN(
        n13500) );
  MUX2_X1 U15521 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n13491), .S(n13490), .Z(
        n13493) );
  INV_X1 U15522 ( .A(n13492), .ZN(n13502) );
  NAND2_X1 U15523 ( .A1(n13493), .A2(n13502), .ZN(n13494) );
  NAND3_X1 U15524 ( .A1(n14370), .A2(n13495), .A3(n13494), .ZN(n13499) );
  AOI22_X1 U15525 ( .A1(n14346), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13498) );
  NAND2_X1 U15526 ( .A1(n14357), .A2(n13496), .ZN(n13497) );
  NAND4_X1 U15527 ( .A1(n13500), .A2(n13499), .A3(n13498), .A4(n13497), .ZN(
        P1_U3244) );
  MUX2_X1 U15528 ( .A(n13502), .B(n13501), .S(n14344), .Z(n13508) );
  NAND2_X1 U15529 ( .A1(n7189), .A2(n13503), .ZN(n13504) );
  NAND2_X1 U15530 ( .A1(n13505), .A2(n13504), .ZN(n14342) );
  AOI21_X1 U15531 ( .B1(n13506), .B2(n14342), .A(n14991), .ZN(n13507) );
  OAI21_X1 U15532 ( .B1(n13508), .B2(n13984), .A(n13507), .ZN(n13550) );
  AOI22_X1 U15533 ( .A1(n14346), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13518) );
  OAI21_X1 U15534 ( .B1(n13510), .B2(n13509), .A(n13522), .ZN(n13511) );
  OAI22_X1 U15535 ( .A1(n13512), .A2(n14375), .B1(n14354), .B2(n13511), .ZN(
        n13513) );
  INV_X1 U15536 ( .A(n13513), .ZN(n13517) );
  OAI211_X1 U15537 ( .C1(n13515), .C2(n13514), .A(n14370), .B(n13527), .ZN(
        n13516) );
  NAND4_X1 U15538 ( .A1(n13550), .A2(n13518), .A3(n13517), .A4(n13516), .ZN(
        P1_U3245) );
  OAI22_X1 U15539 ( .A1(n14992), .A2(n14051), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15061), .ZN(n13519) );
  AOI21_X1 U15540 ( .B1(n13524), .B2(n14357), .A(n13519), .ZN(n13531) );
  MUX2_X1 U15541 ( .A(n9733), .B(P1_REG1_REG_3__SCAN_IN), .S(n13524), .Z(
        n13520) );
  NAND3_X1 U15542 ( .A1(n13522), .A2(n13521), .A3(n13520), .ZN(n13523) );
  NAND3_X1 U15543 ( .A1(n14367), .A2(n13543), .A3(n13523), .ZN(n13530) );
  MUX2_X1 U15544 ( .A(n9717), .B(P1_REG2_REG_3__SCAN_IN), .S(n13524), .Z(
        n13525) );
  NAND3_X1 U15545 ( .A1(n13527), .A2(n13526), .A3(n13525), .ZN(n13528) );
  NAND3_X1 U15546 ( .A1(n14370), .A2(n13538), .A3(n13528), .ZN(n13529) );
  NAND3_X1 U15547 ( .A1(n13531), .A2(n13530), .A3(n13529), .ZN(P1_U3246) );
  NAND2_X1 U15548 ( .A1(n14346), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n13533) );
  OAI211_X1 U15549 ( .C1(n14375), .C2(n13534), .A(n13533), .B(n13532), .ZN(
        n13535) );
  INV_X1 U15550 ( .A(n13535), .ZN(n13549) );
  INV_X1 U15551 ( .A(n13536), .ZN(n13561) );
  NAND3_X1 U15552 ( .A1(n13539), .A2(n13538), .A3(n13537), .ZN(n13540) );
  NAND3_X1 U15553 ( .A1(n14370), .A2(n13561), .A3(n13540), .ZN(n13548) );
  INV_X1 U15554 ( .A(n13541), .ZN(n13546) );
  NAND3_X1 U15555 ( .A1(n13544), .A2(n13543), .A3(n13542), .ZN(n13545) );
  NAND3_X1 U15556 ( .A1(n14367), .A2(n13546), .A3(n13545), .ZN(n13547) );
  NAND4_X1 U15557 ( .A1(n13550), .A2(n13549), .A3(n13548), .A4(n13547), .ZN(
        P1_U3247) );
  INV_X1 U15558 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n15109) );
  NAND2_X1 U15559 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n13551) );
  OAI21_X1 U15560 ( .B1(n14992), .B2(n15109), .A(n13551), .ZN(n13552) );
  AOI21_X1 U15561 ( .B1(n13558), .B2(n14357), .A(n13552), .ZN(n13566) );
  OAI21_X1 U15562 ( .B1(n13555), .B2(n13554), .A(n13553), .ZN(n13556) );
  NAND2_X1 U15563 ( .A1(n14367), .A2(n13556), .ZN(n13565) );
  INV_X1 U15564 ( .A(n13557), .ZN(n13560) );
  MUX2_X1 U15565 ( .A(n10234), .B(P1_REG2_REG_5__SCAN_IN), .S(n13558), .Z(
        n13559) );
  NAND3_X1 U15566 ( .A1(n13561), .A2(n13560), .A3(n13559), .ZN(n13562) );
  NAND3_X1 U15567 ( .A1(n14370), .A2(n13563), .A3(n13562), .ZN(n13564) );
  NAND3_X1 U15568 ( .A1(n13566), .A2(n13565), .A3(n13564), .ZN(P1_U3248) );
  OAI21_X1 U15569 ( .B1(n13569), .B2(n13568), .A(n13567), .ZN(n13570) );
  NAND2_X1 U15570 ( .A1(n13570), .A2(n14367), .ZN(n13580) );
  INV_X1 U15571 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14022) );
  NAND2_X1 U15572 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14227)
         );
  OAI21_X1 U15573 ( .B1(n14992), .B2(n14022), .A(n14227), .ZN(n13571) );
  AOI21_X1 U15574 ( .B1(n14357), .B2(n13572), .A(n13571), .ZN(n13579) );
  OR3_X1 U15575 ( .A1(n13575), .A2(n13574), .A3(n13573), .ZN(n13576) );
  NAND3_X1 U15576 ( .A1(n13577), .A2(n14370), .A3(n13576), .ZN(n13578) );
  NAND3_X1 U15577 ( .A1(n13580), .A2(n13579), .A3(n13578), .ZN(P1_U3254) );
  NAND2_X1 U15578 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14211)
         );
  OAI211_X1 U15579 ( .C1(n13583), .C2(n13582), .A(n13581), .B(n14367), .ZN(
        n13584) );
  AND2_X1 U15580 ( .A1(n14211), .A2(n13584), .ZN(n13591) );
  AOI22_X1 U15581 ( .A1(n14357), .A2(n13585), .B1(n14346), .B2(
        P1_ADDR_REG_16__SCAN_IN), .ZN(n13590) );
  OAI211_X1 U15582 ( .C1(n13588), .C2(n13587), .A(n14370), .B(n13586), .ZN(
        n13589) );
  NAND3_X1 U15583 ( .A1(n13591), .A2(n13590), .A3(n13589), .ZN(P1_U3259) );
  OAI21_X1 U15584 ( .B1(n15023), .B2(n13593), .A(n13592), .ZN(n13594) );
  NAND2_X1 U15585 ( .A1(n13594), .A2(n13601), .ZN(n13595) );
  XOR2_X1 U15586 ( .A(n13601), .B(n13594), .Z(n14368) );
  NAND2_X1 U15587 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n14368), .ZN(n14366) );
  NAND2_X1 U15588 ( .A1(n13595), .A2(n14366), .ZN(n13596) );
  XNOR2_X1 U15589 ( .A(n13597), .B(n13596), .ZN(n13609) );
  NAND2_X1 U15590 ( .A1(n13598), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13600) );
  NAND2_X1 U15591 ( .A1(n13600), .A2(n13599), .ZN(n13602) );
  XOR2_X1 U15592 ( .A(n13601), .B(n13602), .Z(n14371) );
  NAND2_X1 U15593 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14371), .ZN(n14369) );
  NAND2_X1 U15594 ( .A1(n13602), .A2(n13601), .ZN(n13603) );
  NAND2_X1 U15595 ( .A1(n14369), .A2(n13603), .ZN(n13604) );
  XOR2_X1 U15596 ( .A(n13604), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13608) );
  INV_X1 U15597 ( .A(n13608), .ZN(n13605) );
  NAND2_X1 U15598 ( .A1(n13605), .A2(n14370), .ZN(n13606) );
  OAI211_X1 U15599 ( .C1(n13609), .C2(n14354), .A(n13606), .B(n14375), .ZN(
        n13607) );
  INV_X1 U15600 ( .A(n13607), .ZN(n13611) );
  AOI22_X1 U15601 ( .A1(n13609), .A2(n14367), .B1(n14370), .B2(n13608), .ZN(
        n13610) );
  MUX2_X1 U15602 ( .A(n13611), .B(n13610), .S(n13822), .Z(n13614) );
  INV_X1 U15603 ( .A(n13612), .ZN(n13613) );
  OAI211_X1 U15604 ( .C1(n7578), .C2(n14992), .A(n13614), .B(n13613), .ZN(
        P1_U3262) );
  NAND2_X1 U15605 ( .A1(n14250), .A2(n14265), .ZN(n13874) );
  INV_X1 U15606 ( .A(n13780), .ZN(n13931) );
  NAND2_X1 U15607 ( .A1(n13700), .A2(n13714), .ZN(n13699) );
  XNOR2_X1 U15608 ( .A(n13615), .B(n13621), .ZN(n13883) );
  OAI21_X1 U15609 ( .B1(n14344), .B2(n13616), .A(n13835), .ZN(n13676) );
  NOR2_X1 U15610 ( .A1(n13617), .A2(n13676), .ZN(n13884) );
  NAND2_X1 U15611 ( .A1(n14420), .A2(n13884), .ZN(n13623) );
  OAI21_X1 U15612 ( .B1(n14420), .B2(n13618), .A(n13623), .ZN(n13619) );
  AOI21_X1 U15613 ( .B1(n13881), .B2(n14430), .A(n13619), .ZN(n13620) );
  OAI21_X1 U15614 ( .B1(n13883), .B2(n13857), .A(n13620), .ZN(P1_U3263) );
  INV_X1 U15615 ( .A(n13673), .ZN(n13622) );
  INV_X1 U15616 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n13624) );
  OAI21_X1 U15617 ( .B1(n14420), .B2(n13624), .A(n13623), .ZN(n13625) );
  AOI21_X1 U15618 ( .B1(n13626), .B2(n14430), .A(n13625), .ZN(n13627) );
  OAI21_X1 U15619 ( .B1(n13886), .B2(n13875), .A(n13627), .ZN(P1_U3264) );
  OR2_X1 U15620 ( .A1(n14237), .A2(n13628), .ZN(n13629) );
  OR2_X1 U15621 ( .A1(n14271), .A2(n13866), .ZN(n13631) );
  INV_X1 U15622 ( .A(n13632), .ZN(n13633) );
  NAND2_X1 U15623 ( .A1(n13828), .A2(n13636), .ZN(n13639) );
  OR2_X1 U15624 ( .A1(n11568), .A2(n13637), .ZN(n13638) );
  NAND2_X1 U15625 ( .A1(n13639), .A2(n13638), .ZN(n13811) );
  NAND2_X1 U15626 ( .A1(n13950), .A2(n13836), .ZN(n13640) );
  INV_X1 U15627 ( .A(n13665), .ZN(n13807) );
  OR2_X1 U15628 ( .A1(n13793), .A2(n13666), .ZN(n13642) );
  NAND2_X1 U15629 ( .A1(n13780), .A2(n13667), .ZN(n13643) );
  OR2_X1 U15630 ( .A1(n13926), .A2(n13645), .ZN(n13646) );
  NAND2_X1 U15631 ( .A1(n13919), .A2(n13654), .ZN(n13647) );
  NAND2_X1 U15632 ( .A1(n13648), .A2(n13671), .ZN(n13649) );
  INV_X1 U15633 ( .A(n13654), .ZN(n13670) );
  INV_X1 U15634 ( .A(n13950), .ZN(n13664) );
  INV_X1 U15635 ( .A(n14271), .ZN(n13657) );
  NOR2_X1 U15636 ( .A1(n14265), .A2(n13658), .ZN(n13660) );
  NAND2_X1 U15637 ( .A1(n13831), .A2(n13830), .ZN(n13829) );
  INV_X1 U15638 ( .A(n13667), .ZN(n13668) );
  NAND2_X1 U15639 ( .A1(n13780), .A2(n13668), .ZN(n13757) );
  INV_X1 U15640 ( .A(n13747), .ZN(n13738) );
  NOR2_X1 U15641 ( .A1(n13911), .A2(n13671), .ZN(n13709) );
  AOI21_X1 U15642 ( .B1(n13711), .B2(n13689), .A(n13704), .ZN(n13688) );
  INV_X1 U15643 ( .A(n13890), .ZN(n13684) );
  INV_X1 U15644 ( .A(n13699), .ZN(n13674) );
  OAI21_X1 U15645 ( .B1(n13684), .B2(n13674), .A(n13673), .ZN(n13892) );
  NOR2_X1 U15646 ( .A1(n13892), .A2(n13857), .ZN(n13686) );
  NOR2_X1 U15647 ( .A1(n13675), .A2(n14382), .ZN(n13889) );
  NOR2_X1 U15648 ( .A1(n13677), .A2(n13676), .ZN(n13888) );
  INV_X1 U15649 ( .A(n13888), .ZN(n13680) );
  OAI22_X1 U15650 ( .A1(n13680), .A2(n13679), .B1(n13678), .B2(n14416), .ZN(
        n13681) );
  AOI21_X1 U15651 ( .B1(n13889), .B2(n14420), .A(n13681), .ZN(n13683) );
  NAND2_X1 U15652 ( .A1(n14439), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n13682) );
  OAI211_X1 U15653 ( .C1(n13684), .C2(n13876), .A(n13683), .B(n13682), .ZN(
        n13685) );
  AOI211_X1 U15654 ( .C1(n13894), .C2(n13842), .A(n13686), .B(n13685), .ZN(
        n13687) );
  OAI21_X1 U15655 ( .B1(n13895), .B2(n13844), .A(n13687), .ZN(P1_U3356) );
  INV_X1 U15656 ( .A(n13688), .ZN(n13691) );
  NAND3_X1 U15657 ( .A1(n13711), .A2(n13704), .A3(n13689), .ZN(n13690) );
  NAND2_X1 U15658 ( .A1(n13691), .A2(n13690), .ZN(n13692) );
  AOI22_X1 U15659 ( .A1(n13865), .A2(n13694), .B1(n13693), .B2(n13835), .ZN(
        n13695) );
  OAI22_X1 U15660 ( .A1(n14420), .A2(n13698), .B1(n13697), .B2(n14416), .ZN(
        n13702) );
  OAI211_X1 U15661 ( .C1(n13700), .C2(n13714), .A(n13699), .B(n14412), .ZN(
        n13900) );
  NOR2_X1 U15662 ( .A1(n13900), .A2(n13875), .ZN(n13701) );
  AOI211_X1 U15663 ( .C1(n14430), .C2(n13898), .A(n13702), .B(n13701), .ZN(
        n13708) );
  INV_X1 U15664 ( .A(n13703), .ZN(n13706) );
  INV_X1 U15665 ( .A(n13704), .ZN(n13705) );
  NAND2_X1 U15666 ( .A1(n13706), .A2(n13705), .ZN(n13897) );
  NAND3_X1 U15667 ( .A1(n13897), .A2(n14252), .A3(n13896), .ZN(n13707) );
  OAI211_X1 U15668 ( .C1(n13904), .C2(n14439), .A(n13708), .B(n13707), .ZN(
        P1_U3265) );
  NOR2_X1 U15669 ( .A1(n13713), .A2(n13712), .ZN(n13908) );
  INV_X1 U15670 ( .A(n13728), .ZN(n13715) );
  AOI211_X1 U15671 ( .C1(n13906), .C2(n13715), .A(n14468), .B(n13714), .ZN(
        n13905) );
  INV_X1 U15672 ( .A(n13716), .ZN(n13717) );
  AOI22_X1 U15673 ( .A1(n14439), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13717), 
        .B2(n14431), .ZN(n13718) );
  OAI21_X1 U15674 ( .B1(n13719), .B2(n13876), .A(n13718), .ZN(n13723) );
  AOI21_X1 U15675 ( .B1(n13721), .B2(n13720), .A(n6507), .ZN(n13909) );
  NOR2_X1 U15676 ( .A1(n13909), .A2(n13844), .ZN(n13722) );
  AOI211_X1 U15677 ( .C1(n13905), .C2(n14436), .A(n13723), .B(n13722), .ZN(
        n13724) );
  OAI21_X1 U15678 ( .B1(n13908), .B2(n14439), .A(n13724), .ZN(P1_U3266) );
  OAI21_X1 U15679 ( .B1(n13726), .B2(n6481), .A(n13725), .ZN(n13916) );
  OAI21_X1 U15680 ( .B1(n6486), .B2(n13911), .A(n14412), .ZN(n13729) );
  NOR2_X1 U15681 ( .A1(n13729), .A2(n13728), .ZN(n13913) );
  NAND2_X1 U15682 ( .A1(n13913), .A2(n14436), .ZN(n13733) );
  OAI22_X1 U15683 ( .A1(n14439), .A2(n13910), .B1(n13730), .B2(n14416), .ZN(
        n13731) );
  AOI21_X1 U15684 ( .B1(P1_REG2_REG_26__SCAN_IN), .B2(n14439), .A(n13731), 
        .ZN(n13732) );
  OAI211_X1 U15685 ( .C1(n13911), .C2(n13876), .A(n13733), .B(n13732), .ZN(
        n13734) );
  AOI21_X1 U15686 ( .B1(n13914), .B2(n13842), .A(n13734), .ZN(n13735) );
  OAI21_X1 U15687 ( .B1(n13844), .B2(n13916), .A(n13735), .ZN(P1_U3267) );
  INV_X1 U15688 ( .A(n13917), .ZN(n13751) );
  NAND2_X1 U15689 ( .A1(n13762), .A2(n13919), .ZN(n13741) );
  NAND2_X1 U15690 ( .A1(n13741), .A2(n14412), .ZN(n13742) );
  NOR2_X1 U15691 ( .A1(n6486), .A2(n13742), .ZN(n13918) );
  INV_X1 U15692 ( .A(n13743), .ZN(n13744) );
  AOI22_X1 U15693 ( .A1(n14439), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n13744), 
        .B2(n14431), .ZN(n13745) );
  OAI21_X1 U15694 ( .B1(n6945), .B2(n13876), .A(n13745), .ZN(n13746) );
  AOI21_X1 U15695 ( .B1(n13918), .B2(n14436), .A(n13746), .ZN(n13750) );
  NAND2_X1 U15696 ( .A1(n13748), .A2(n13747), .ZN(n13920) );
  NAND3_X1 U15697 ( .A1(n13921), .A2(n13920), .A3(n14252), .ZN(n13749) );
  OAI211_X1 U15698 ( .C1(n13751), .C2(n14439), .A(n13750), .B(n13749), .ZN(
        P1_U3268) );
  INV_X1 U15699 ( .A(n13752), .ZN(n13753) );
  AOI21_X1 U15700 ( .B1(n13756), .B2(n13754), .A(n13753), .ZN(n13928) );
  NAND2_X1 U15701 ( .A1(n13755), .A2(n14429), .ZN(n13761) );
  INV_X1 U15702 ( .A(n13758), .ZN(n13759) );
  OAI21_X1 U15703 ( .B1(n13761), .B2(n13760), .A(n13759), .ZN(n13924) );
  NAND2_X1 U15704 ( .A1(n13924), .A2(n14420), .ZN(n13769) );
  INV_X1 U15705 ( .A(n13762), .ZN(n13763) );
  AOI211_X1 U15706 ( .C1(n13926), .C2(n13774), .A(n14468), .B(n13763), .ZN(
        n13925) );
  NOR2_X1 U15707 ( .A1(n6946), .A2(n13876), .ZN(n13767) );
  OAI22_X1 U15708 ( .A1(n14420), .A2(n13765), .B1(n13764), .B2(n14416), .ZN(
        n13766) );
  AOI211_X1 U15709 ( .C1(n13925), .C2(n14436), .A(n13767), .B(n13766), .ZN(
        n13768) );
  OAI211_X1 U15710 ( .C1(n13844), .C2(n13928), .A(n13769), .B(n13768), .ZN(
        P1_U3269) );
  OAI21_X1 U15711 ( .B1(n6505), .B2(n7241), .A(n13770), .ZN(n13935) );
  OAI21_X1 U15712 ( .B1(n13773), .B2(n13772), .A(n13771), .ZN(n13933) );
  OAI211_X1 U15713 ( .C1(n13787), .C2(n13931), .A(n13774), .B(n14412), .ZN(
        n13930) );
  NOR2_X1 U15714 ( .A1(n14420), .A2(n13775), .ZN(n13776) );
  AOI21_X1 U15715 ( .B1(n13777), .B2(n14431), .A(n13776), .ZN(n13778) );
  OAI21_X1 U15716 ( .B1(n13929), .B2(n14439), .A(n13778), .ZN(n13779) );
  AOI21_X1 U15717 ( .B1(n13780), .B2(n14430), .A(n13779), .ZN(n13781) );
  OAI21_X1 U15718 ( .B1(n13930), .B2(n13875), .A(n13781), .ZN(n13782) );
  AOI21_X1 U15719 ( .B1(n13933), .B2(n13842), .A(n13782), .ZN(n13783) );
  OAI21_X1 U15720 ( .B1(n13844), .B2(n13935), .A(n13783), .ZN(P1_U3270) );
  XOR2_X1 U15721 ( .A(n13785), .B(n13784), .Z(n13943) );
  XNOR2_X1 U15722 ( .A(n13786), .B(n13785), .ZN(n13941) );
  INV_X1 U15723 ( .A(n13787), .ZN(n13789) );
  AOI21_X1 U15724 ( .B1(n13801), .B2(n13793), .A(n14468), .ZN(n13788) );
  NAND2_X1 U15725 ( .A1(n13789), .A2(n13788), .ZN(n13938) );
  INV_X1 U15726 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n13790) );
  OAI22_X1 U15727 ( .A1(n13791), .A2(n14416), .B1(n13790), .B2(n14420), .ZN(
        n13792) );
  AOI21_X1 U15728 ( .B1(n13936), .B2(n14420), .A(n13792), .ZN(n13795) );
  NAND2_X1 U15729 ( .A1(n13793), .A2(n14430), .ZN(n13794) );
  OAI211_X1 U15730 ( .C1(n13938), .C2(n13875), .A(n13795), .B(n13794), .ZN(
        n13796) );
  AOI21_X1 U15731 ( .B1(n13941), .B2(n13842), .A(n13796), .ZN(n13797) );
  OAI21_X1 U15732 ( .B1(n13943), .B2(n13844), .A(n13797), .ZN(P1_U3271) );
  XNOR2_X1 U15733 ( .A(n13798), .B(n13807), .ZN(n13800) );
  AOI21_X1 U15734 ( .B1(n13800), .B2(n14429), .A(n13799), .ZN(n13947) );
  INV_X1 U15735 ( .A(n13801), .ZN(n13802) );
  AOI211_X1 U15736 ( .C1(n13945), .C2(n13820), .A(n14468), .B(n13802), .ZN(
        n13944) );
  INV_X1 U15737 ( .A(n13803), .ZN(n13804) );
  AOI22_X1 U15738 ( .A1(n14439), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n13804), 
        .B2(n14431), .ZN(n13805) );
  OAI21_X1 U15739 ( .B1(n6938), .B2(n13876), .A(n13805), .ZN(n13809) );
  AOI21_X1 U15740 ( .B1(n13807), .B2(n13806), .A(n6515), .ZN(n13948) );
  NOR2_X1 U15741 ( .A1(n13948), .A2(n13844), .ZN(n13808) );
  AOI211_X1 U15742 ( .C1(n13944), .C2(n14436), .A(n13809), .B(n13808), .ZN(
        n13810) );
  OAI21_X1 U15743 ( .B1(n13947), .B2(n14439), .A(n13810), .ZN(P1_U3272) );
  INV_X1 U15744 ( .A(n13811), .ZN(n13813) );
  OAI21_X1 U15745 ( .B1(n13813), .B2(n13816), .A(n13812), .ZN(n13953) );
  AOI211_X1 U15746 ( .C1(n13816), .C2(n13815), .A(n14540), .B(n13814), .ZN(
        n13819) );
  OAI22_X1 U15747 ( .A1(n13817), .A2(n14380), .B1(n13848), .B2(n14382), .ZN(
        n13818) );
  NOR2_X1 U15748 ( .A1(n13819), .A2(n13818), .ZN(n13952) );
  AOI21_X1 U15749 ( .B1(n13950), .B2(n13832), .A(n14468), .ZN(n13821) );
  AND2_X1 U15750 ( .A1(n13821), .A2(n13820), .ZN(n13949) );
  NAND2_X1 U15751 ( .A1(n13949), .A2(n13822), .ZN(n13823) );
  OAI211_X1 U15752 ( .C1(n14416), .C2(n13824), .A(n13952), .B(n13823), .ZN(
        n13825) );
  NAND2_X1 U15753 ( .A1(n13825), .A2(n14420), .ZN(n13827) );
  AOI22_X1 U15754 ( .A1(n13950), .A2(n14430), .B1(P1_REG2_REG_20__SCAN_IN), 
        .B2(n14439), .ZN(n13826) );
  OAI211_X1 U15755 ( .C1(n13953), .C2(n13844), .A(n13827), .B(n13826), .ZN(
        P1_U3273) );
  XNOR2_X1 U15756 ( .A(n13828), .B(n13830), .ZN(n13959) );
  OAI21_X1 U15757 ( .B1(n13831), .B2(n13830), .A(n13829), .ZN(n13957) );
  AOI21_X1 U15758 ( .B1(n11568), .B2(n13856), .A(n14468), .ZN(n13833) );
  NAND2_X1 U15759 ( .A1(n13833), .A2(n13832), .ZN(n13955) );
  AOI22_X1 U15760 ( .A1(n13836), .A2(n13835), .B1(n13865), .B2(n13834), .ZN(
        n13954) );
  OAI22_X1 U15761 ( .A1(n13954), .A2(n14439), .B1(n13837), .B2(n14416), .ZN(
        n13839) );
  NOR2_X1 U15762 ( .A1(n6940), .A2(n13876), .ZN(n13838) );
  AOI211_X1 U15763 ( .C1(n14439), .C2(P1_REG2_REG_19__SCAN_IN), .A(n13839), 
        .B(n13838), .ZN(n13840) );
  OAI21_X1 U15764 ( .B1(n13875), .B2(n13955), .A(n13840), .ZN(n13841) );
  AOI21_X1 U15765 ( .B1(n13957), .B2(n13842), .A(n13841), .ZN(n13843) );
  OAI21_X1 U15766 ( .B1(n13959), .B2(n13844), .A(n13843), .ZN(P1_U3274) );
  XNOR2_X1 U15767 ( .A(n13845), .B(n13846), .ZN(n14256) );
  XNOR2_X1 U15768 ( .A(n13847), .B(n13846), .ZN(n13850) );
  OAI22_X1 U15769 ( .A1(n13848), .A2(n14380), .B1(n14209), .B2(n14382), .ZN(
        n13849) );
  AOI21_X1 U15770 ( .B1(n13850), .B2(n14429), .A(n13849), .ZN(n13851) );
  OAI21_X1 U15771 ( .B1(n14256), .B2(n14509), .A(n13851), .ZN(n14259) );
  NAND2_X1 U15772 ( .A1(n14259), .A2(n14420), .ZN(n13862) );
  INV_X1 U15773 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n13854) );
  INV_X1 U15774 ( .A(n13852), .ZN(n13853) );
  OAI22_X1 U15775 ( .A1(n14420), .A2(n13854), .B1(n13853), .B2(n14416), .ZN(
        n13859) );
  NAND2_X1 U15776 ( .A1(n13860), .A2(n13874), .ZN(n13855) );
  NAND2_X1 U15777 ( .A1(n13856), .A2(n13855), .ZN(n14258) );
  NOR2_X1 U15778 ( .A1(n14258), .A2(n13857), .ZN(n13858) );
  AOI211_X1 U15779 ( .C1(n14430), .C2(n13860), .A(n13859), .B(n13858), .ZN(
        n13861) );
  OAI211_X1 U15780 ( .C1(n14256), .C2(n14121), .A(n13862), .B(n13861), .ZN(
        P1_U3275) );
  INV_X1 U15781 ( .A(n13863), .ZN(n13871) );
  OR2_X1 U15782 ( .A1(n13864), .A2(n14380), .ZN(n13868) );
  NAND2_X1 U15783 ( .A1(n13866), .A2(n13865), .ZN(n13867) );
  NAND2_X1 U15784 ( .A1(n13868), .A2(n13867), .ZN(n14262) );
  XOR2_X1 U15785 ( .A(n13869), .B(n13872), .Z(n13870) );
  NOR2_X1 U15786 ( .A1(n13870), .A2(n14540), .ZN(n14266) );
  AOI211_X1 U15787 ( .C1(n14431), .C2(n13871), .A(n14262), .B(n14266), .ZN(
        n13880) );
  XOR2_X1 U15788 ( .A(n13873), .B(n13872), .Z(n14268) );
  OAI211_X1 U15789 ( .C1(n14250), .C2(n14265), .A(n13874), .B(n14412), .ZN(
        n14264) );
  NOR2_X1 U15790 ( .A1(n14264), .A2(n13875), .ZN(n13878) );
  OAI22_X1 U15791 ( .A1(n14265), .A2(n13876), .B1(n14420), .B2(n11132), .ZN(
        n13877) );
  AOI211_X1 U15792 ( .C1(n14268), .C2(n14252), .A(n13878), .B(n13877), .ZN(
        n13879) );
  OAI21_X1 U15793 ( .B1(n13880), .B2(n14439), .A(n13879), .ZN(P1_U3276) );
  AOI21_X1 U15794 ( .B1(n13881), .B2(n14538), .A(n13884), .ZN(n13882) );
  OAI21_X1 U15795 ( .B1(n13883), .B2(n14468), .A(n13882), .ZN(n13960) );
  MUX2_X1 U15796 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n13960), .S(n14563), .Z(
        P1_U3559) );
  INV_X1 U15797 ( .A(n13884), .ZN(n13885) );
  MUX2_X1 U15798 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n13961), .S(n14563), .Z(
        P1_U3558) );
  AOI211_X1 U15799 ( .C1(n13890), .C2(n14538), .A(n13889), .B(n13888), .ZN(
        n13891) );
  OAI21_X1 U15800 ( .B1(n13892), .B2(n14468), .A(n13891), .ZN(n13893) );
  MUX2_X1 U15801 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n13962), .S(n14563), .Z(
        P1_U3557) );
  NAND3_X1 U15802 ( .A1(n13897), .A2(n14544), .A3(n13896), .ZN(n13902) );
  NAND2_X1 U15803 ( .A1(n13898), .A2(n14538), .ZN(n13899) );
  MUX2_X1 U15804 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n13963), .S(n14563), .Z(
        P1_U3556) );
  AOI21_X1 U15805 ( .B1(n14538), .B2(n13906), .A(n13905), .ZN(n13907) );
  MUX2_X1 U15806 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n13964), .S(n14563), .Z(
        P1_U3555) );
  OAI21_X1 U15807 ( .B1(n13911), .B2(n14528), .A(n13910), .ZN(n13912) );
  AOI211_X1 U15808 ( .C1(n13914), .C2(n14429), .A(n13913), .B(n13912), .ZN(
        n13915) );
  MUX2_X1 U15809 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n13965), .S(n14563), .Z(
        P1_U3554) );
  NAND3_X1 U15810 ( .A1(n13921), .A2(n13920), .A3(n14544), .ZN(n13922) );
  NAND2_X1 U15811 ( .A1(n13923), .A2(n13922), .ZN(n13966) );
  MUX2_X1 U15812 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n13966), .S(n14563), .Z(
        P1_U3553) );
  AOI211_X1 U15813 ( .C1(n14538), .C2(n13926), .A(n13925), .B(n13924), .ZN(
        n13927) );
  MUX2_X1 U15814 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n13967), .S(n14563), .Z(
        P1_U3552) );
  OAI211_X1 U15815 ( .C1(n13931), .C2(n14528), .A(n13930), .B(n13929), .ZN(
        n13932) );
  AOI21_X1 U15816 ( .B1(n13933), .B2(n14429), .A(n13932), .ZN(n13934) );
  OAI21_X1 U15817 ( .B1(n14489), .B2(n13935), .A(n13934), .ZN(n13968) );
  MUX2_X1 U15818 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n13968), .S(n14563), .Z(
        P1_U3551) );
  INV_X1 U15819 ( .A(n13936), .ZN(n13937) );
  OAI211_X1 U15820 ( .C1(n14528), .C2(n13939), .A(n13938), .B(n13937), .ZN(
        n13940) );
  AOI21_X1 U15821 ( .B1(n13941), .B2(n14429), .A(n13940), .ZN(n13942) );
  OAI21_X1 U15822 ( .B1(n14489), .B2(n13943), .A(n13942), .ZN(n13969) );
  MUX2_X1 U15823 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n13969), .S(n14563), .Z(
        P1_U3550) );
  AOI21_X1 U15824 ( .B1(n14538), .B2(n13945), .A(n13944), .ZN(n13946) );
  OAI211_X1 U15825 ( .C1(n14489), .C2(n13948), .A(n13947), .B(n13946), .ZN(
        n13970) );
  MUX2_X1 U15826 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n13970), .S(n14563), .Z(
        P1_U3549) );
  AOI21_X1 U15827 ( .B1(n14538), .B2(n13950), .A(n13949), .ZN(n13951) );
  OAI211_X1 U15828 ( .C1(n14489), .C2(n13953), .A(n13952), .B(n13951), .ZN(
        n13971) );
  MUX2_X1 U15829 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n13971), .S(n14563), .Z(
        P1_U3548) );
  OAI211_X1 U15830 ( .C1(n6940), .C2(n14528), .A(n13955), .B(n13954), .ZN(
        n13956) );
  AOI21_X1 U15831 ( .B1(n13957), .B2(n14429), .A(n13956), .ZN(n13958) );
  OAI21_X1 U15832 ( .B1(n14489), .B2(n13959), .A(n13958), .ZN(n13972) );
  MUX2_X1 U15833 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n13972), .S(n14563), .Z(
        P1_U3547) );
  MUX2_X1 U15834 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n13960), .S(n14546), .Z(
        P1_U3527) );
  MUX2_X1 U15835 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n13961), .S(n14546), .Z(
        P1_U3526) );
  MUX2_X1 U15836 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n13963), .S(n14546), .Z(
        P1_U3524) );
  MUX2_X1 U15837 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n13964), .S(n14546), .Z(
        P1_U3523) );
  MUX2_X1 U15838 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n13966), .S(n14546), .Z(
        P1_U3521) );
  MUX2_X1 U15839 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n13968), .S(n14546), .Z(
        P1_U3519) );
  MUX2_X1 U15840 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n13969), .S(n14546), .Z(
        P1_U3518) );
  MUX2_X1 U15841 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n13970), .S(n14546), .Z(
        P1_U3517) );
  MUX2_X1 U15842 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n13971), .S(n14546), .Z(
        P1_U3516) );
  MUX2_X1 U15843 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n13972), .S(n14546), .Z(
        P1_U3515) );
  NOR4_X1 U15844 ( .A1(n13974), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n13973), .ZN(n13975) );
  AOI21_X1 U15845 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n13976), .A(n13975), 
        .ZN(n13977) );
  OAI21_X1 U15846 ( .B1(n13978), .B2(n13986), .A(n13977), .ZN(P1_U3324) );
  OAI222_X1 U15847 ( .A1(n13986), .A2(n13981), .B1(n13979), .B2(P1_U3086), 
        .C1(n13980), .C2(n13988), .ZN(P1_U3325) );
  OAI222_X1 U15848 ( .A1(n13986), .A2(n13983), .B1(n9558), .B2(P1_U3086), .C1(
        n13982), .C2(n13988), .ZN(P1_U3326) );
  OAI222_X1 U15849 ( .A1(n13988), .A2(n13987), .B1(n13986), .B2(n13985), .C1(
        P1_U3086), .C2(n13984), .ZN(P1_U3327) );
  OAI222_X1 U15850 ( .A1(n13986), .A2(n13990), .B1(n14344), .B2(P1_U3086), 
        .C1(n13989), .C2(n13988), .ZN(P1_U3328) );
  OAI222_X1 U15851 ( .A1(n13986), .A2(n13993), .B1(P1_U3086), .B2(n13992), 
        .C1(n13991), .C2(n13988), .ZN(P1_U3329) );
  MUX2_X1 U15852 ( .A(n13995), .B(n13994), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U15853 ( .A(n13996), .ZN(n13997) );
  MUX2_X1 U15854 ( .A(n13997), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U15855 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14602) );
  NAND2_X1 U15856 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14089), .ZN(n14090) );
  OAI21_X1 U15857 ( .B1(n14089), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n14090), 
        .ZN(n14031) );
  INV_X1 U15858 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14365) );
  NOR2_X1 U15859 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14365), .ZN(n14030) );
  NOR2_X1 U15860 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n13998), .ZN(n14028) );
  INV_X1 U15861 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14026) );
  INV_X1 U15862 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14024) );
  XOR2_X1 U15863 ( .A(n13999), .B(n14024), .Z(n14080) );
  INV_X1 U15864 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14000) );
  XNOR2_X1 U15865 ( .A(n14000), .B(n14022), .ZN(n14034) );
  XNOR2_X1 U15866 ( .A(n15066), .B(P3_ADDR_REG_9__SCAN_IN), .ZN(n14073) );
  XNOR2_X1 U15867 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n14038) );
  NAND2_X1 U15868 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14002), .ZN(n14003) );
  NAND2_X1 U15869 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14004), .ZN(n14007) );
  INV_X1 U15870 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14005) );
  NAND2_X1 U15871 ( .A1(n14040), .A2(n14005), .ZN(n14006) );
  NAND2_X1 U15872 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14008), .ZN(n14010) );
  OR2_X1 U15873 ( .A1(n14012), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14011) );
  INV_X1 U15874 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14838) );
  NAND2_X1 U15875 ( .A1(n14013), .A2(n14838), .ZN(n14015) );
  XNOR2_X1 U15876 ( .A(n14013), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n14064) );
  NAND2_X1 U15877 ( .A1(n14064), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14014) );
  NAND2_X1 U15878 ( .A1(n14015), .A2(n14014), .ZN(n14039) );
  NAND2_X1 U15879 ( .A1(n14038), .A2(n14039), .ZN(n14016) );
  XOR2_X1 U15880 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14020), .Z(n14036) );
  NAND2_X1 U15881 ( .A1(n14037), .A2(n14036), .ZN(n14019) );
  NAND2_X1 U15882 ( .A1(n14034), .A2(n14035), .ZN(n14021) );
  AND2_X1 U15883 ( .A1(n14026), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14025) );
  OAI22_X1 U15884 ( .A1(n14028), .A2(n14083), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n14027), .ZN(n14085) );
  INV_X1 U15885 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14029) );
  OAI22_X1 U15886 ( .A1(n14030), .A2(n14085), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14029), .ZN(n14091) );
  XOR2_X1 U15887 ( .A(n14031), .B(n14091), .Z(n14340) );
  INV_X1 U15888 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14576) );
  INV_X1 U15889 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14329) );
  XOR2_X1 U15890 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .Z(n14032) );
  XNOR2_X1 U15891 ( .A(n14033), .B(n14032), .ZN(n14328) );
  XOR2_X1 U15892 ( .A(n14035), .B(n14034), .Z(n14319) );
  XOR2_X1 U15893 ( .A(n14037), .B(n14036), .Z(n14110) );
  XOR2_X1 U15894 ( .A(n14039), .B(n14038), .Z(n14069) );
  NAND2_X1 U15895 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14041), .ZN(n14054) );
  INV_X1 U15896 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14103) );
  XNOR2_X1 U15897 ( .A(n14043), .B(n14042), .ZN(n14101) );
  XNOR2_X1 U15898 ( .A(n14045), .B(n14044), .ZN(n14046) );
  NAND2_X1 U15899 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14046), .ZN(n14048) );
  AOI21_X1 U15900 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14750), .A(n14045), .ZN(
        n15146) );
  INV_X1 U15901 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15145) );
  NOR2_X1 U15902 ( .A1(n15146), .A2(n15145), .ZN(n15154) );
  XOR2_X1 U15903 ( .A(n14046), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15153) );
  NAND2_X1 U15904 ( .A1(n15154), .A2(n15153), .ZN(n14047) );
  NAND2_X1 U15905 ( .A1(n14048), .A2(n14047), .ZN(n14102) );
  NAND2_X1 U15906 ( .A1(n14101), .A2(n14102), .ZN(n14049) );
  NOR2_X1 U15907 ( .A1(n14101), .A2(n14102), .ZN(n14100) );
  AOI21_X1 U15908 ( .B1(n14103), .B2(n14049), .A(n14100), .ZN(n15150) );
  XNOR2_X1 U15909 ( .A(n14051), .B(n14050), .ZN(n15151) );
  NOR2_X1 U15910 ( .A1(n15150), .A2(n15151), .ZN(n14053) );
  NAND2_X1 U15911 ( .A1(n15150), .A2(n15151), .ZN(n15149) );
  OAI21_X1 U15912 ( .B1(n14053), .B2(n14052), .A(n15149), .ZN(n15142) );
  XNOR2_X1 U15913 ( .A(n15109), .B(n14055), .ZN(n14056) );
  NOR2_X1 U15914 ( .A1(n14057), .A2(n14056), .ZN(n14059) );
  NOR2_X1 U15915 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15144), .ZN(n14058) );
  NAND2_X1 U15916 ( .A1(n14060), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14063) );
  XNOR2_X1 U15917 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14062) );
  XNOR2_X1 U15918 ( .A(n14062), .B(n14061), .ZN(n14105) );
  NAND2_X1 U15919 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14065), .ZN(n14067) );
  XOR2_X1 U15920 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14064), .Z(n15148) );
  NAND2_X1 U15921 ( .A1(n14067), .A2(n14066), .ZN(n14068) );
  NOR2_X1 U15922 ( .A1(n14069), .A2(n14068), .ZN(n14071) );
  XNOR2_X1 U15923 ( .A(n14069), .B(n14068), .ZN(n14107) );
  NOR2_X1 U15924 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n14107), .ZN(n14070) );
  XNOR2_X1 U15925 ( .A(n14073), .B(n14072), .ZN(n14075) );
  NAND2_X1 U15926 ( .A1(n14074), .A2(n14075), .ZN(n14076) );
  NAND2_X1 U15927 ( .A1(n14110), .A2(n14111), .ZN(n14109) );
  NOR2_X1 U15928 ( .A1(n14319), .A2(n14320), .ZN(n14078) );
  INV_X1 U15929 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14077) );
  NAND2_X1 U15930 ( .A1(n14319), .A2(n14320), .ZN(n14318) );
  XNOR2_X1 U15931 ( .A(n14080), .B(n14079), .ZN(n14323) );
  INV_X1 U15932 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14081) );
  NAND2_X1 U15933 ( .A1(n14324), .A2(n14323), .ZN(n14322) );
  XNOR2_X1 U15934 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n14084) );
  XNOR2_X1 U15935 ( .A(n14084), .B(n14083), .ZN(n14333) );
  XNOR2_X1 U15936 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14086) );
  XOR2_X1 U15937 ( .A(n14086), .B(n14085), .Z(n14336) );
  NOR2_X1 U15938 ( .A1(n6482), .A2(n14336), .ZN(n14088) );
  INV_X1 U15939 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14087) );
  NAND2_X1 U15940 ( .A1(n6482), .A2(n14336), .ZN(n14335) );
  NOR2_X1 U15941 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14089), .ZN(n14092) );
  OAI21_X1 U15942 ( .B1(n14092), .B2(n14091), .A(n14090), .ZN(n14093) );
  XOR2_X1 U15943 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14093), .Z(n14094) );
  XNOR2_X1 U15944 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14094), .ZN(n14136) );
  INV_X1 U15945 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15033) );
  NOR2_X1 U15946 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14093), .ZN(n14096) );
  AND2_X1 U15947 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14094), .ZN(n14095) );
  NOR2_X1 U15948 ( .A1(n14096), .A2(n14095), .ZN(n14139) );
  XOR2_X1 U15949 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n14097) );
  XNOR2_X1 U15950 ( .A(n14139), .B(n14097), .ZN(n14144) );
  XNOR2_X1 U15951 ( .A(n14143), .B(n14144), .ZN(n14145) );
  XNOR2_X1 U15952 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14145), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U15953 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14098) );
  OAI21_X1 U15954 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14098), 
        .ZN(U28) );
  AOI21_X1 U15955 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14099) );
  OAI21_X1 U15956 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14099), 
        .ZN(U29) );
  AOI21_X1 U15957 ( .B1(n14102), .B2(n14101), .A(n14100), .ZN(n14104) );
  XNOR2_X1 U15958 ( .A(n14104), .B(n14103), .ZN(SUB_1596_U61) );
  XOR2_X1 U15959 ( .A(n14106), .B(n14105), .Z(SUB_1596_U57) );
  XNOR2_X1 U15960 ( .A(n14107), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U15961 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14108), .Z(SUB_1596_U54) );
  OAI21_X1 U15962 ( .B1(n14111), .B2(n14110), .A(n14109), .ZN(n14112) );
  XNOR2_X1 U15963 ( .A(n14112), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  XNOR2_X1 U15964 ( .A(n14113), .B(n6957), .ZN(n14131) );
  XNOR2_X1 U15965 ( .A(n14115), .B(n14114), .ZN(n14117) );
  OAI21_X1 U15966 ( .B1(n14117), .B2(n14540), .A(n14116), .ZN(n14118) );
  AOI21_X1 U15967 ( .B1(n14532), .B2(n14131), .A(n14118), .ZN(n14128) );
  AOI222_X1 U15968 ( .A1(n14120), .A2(n14430), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n14439), .C1(n14431), .C2(n14119), .ZN(n14126) );
  INV_X1 U15969 ( .A(n14121), .ZN(n14434) );
  OAI211_X1 U15970 ( .C1(n6937), .C2(n6936), .A(n14412), .B(n14123), .ZN(
        n14127) );
  INV_X1 U15971 ( .A(n14127), .ZN(n14124) );
  AOI22_X1 U15972 ( .A1(n14131), .A2(n14434), .B1(n14436), .B2(n14124), .ZN(
        n14125) );
  OAI211_X1 U15973 ( .C1(n14439), .C2(n14128), .A(n14126), .B(n14125), .ZN(
        P1_U3281) );
  INV_X1 U15974 ( .A(n14523), .ZN(n14504) );
  OAI21_X1 U15975 ( .B1(n6936), .B2(n14528), .A(n14127), .ZN(n14130) );
  INV_X1 U15976 ( .A(n14128), .ZN(n14129) );
  AOI211_X1 U15977 ( .C1(n14504), .C2(n14131), .A(n14130), .B(n14129), .ZN(
        n14133) );
  INV_X1 U15978 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14132) );
  AOI22_X1 U15979 ( .A1(n14546), .A2(n14133), .B1(n14132), .B2(n7230), .ZN(
        P1_U3495) );
  AOI22_X1 U15980 ( .A1(n14563), .A2(n14133), .B1(n10988), .B2(n14561), .ZN(
        P1_U3540) );
  OAI21_X1 U15981 ( .B1(n14136), .B2(n14135), .A(n14134), .ZN(n14137) );
  XNOR2_X1 U15982 ( .A(n14137), .B(P2_ADDR_REG_17__SCAN_IN), .ZN(SUB_1596_U63)
         );
  INV_X1 U15983 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15019) );
  NOR2_X1 U15984 ( .A1(P3_ADDR_REG_18__SCAN_IN), .A2(n15019), .ZN(n14138) );
  OAI22_X1 U15985 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n12135), .B1(n14139), 
        .B2(n14138), .ZN(n14142) );
  XNOR2_X1 U15986 ( .A(n14140), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n14141) );
  XNOR2_X1 U15987 ( .A(n14142), .B(n14141), .ZN(n14146) );
  AOI21_X1 U15988 ( .B1(n8639), .B2(n14148), .A(n14147), .ZN(n14161) );
  OAI21_X1 U15989 ( .B1(n14150), .B2(P3_REG1_REG_17__SCAN_IN), .A(n14149), 
        .ZN(n14159) );
  OAI211_X1 U15990 ( .C1(n14153), .C2(n14152), .A(n14151), .B(n14863), .ZN(
        n14156) );
  AOI21_X1 U15991 ( .B1(n14871), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n14154), 
        .ZN(n14155) );
  OAI211_X1 U15992 ( .C1(n14868), .C2(n14157), .A(n14156), .B(n14155), .ZN(
        n14158) );
  AOI21_X1 U15993 ( .B1(n14874), .B2(n14159), .A(n14158), .ZN(n14160) );
  OAI21_X1 U15994 ( .B1(n14161), .B2(n14878), .A(n14160), .ZN(P3_U3199) );
  AOI22_X1 U15995 ( .A1(n14163), .A2(n14972), .B1(n14960), .B2(n14162), .ZN(
        n14164) );
  AND2_X1 U15996 ( .A1(n14165), .A2(n14164), .ZN(n14176) );
  INV_X1 U15997 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14166) );
  AOI22_X1 U15998 ( .A1(n14990), .A2(n14176), .B1(n14166), .B2(n14987), .ZN(
        P3_U3472) );
  AOI22_X1 U15999 ( .A1(n14168), .A2(n14972), .B1(n14960), .B2(n14167), .ZN(
        n14170) );
  AOI22_X1 U16000 ( .A1(n14990), .A2(n14177), .B1(n12021), .B2(n14987), .ZN(
        P3_U3471) );
  AOI211_X1 U16001 ( .C1(n14972), .C2(n14173), .A(n14172), .B(n14171), .ZN(
        n14178) );
  INV_X1 U16002 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14174) );
  AOI22_X1 U16003 ( .A1(n14990), .A2(n14178), .B1(n14174), .B2(n14987), .ZN(
        P3_U3470) );
  INV_X1 U16004 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14175) );
  AOI22_X1 U16005 ( .A1(n14974), .A2(n14176), .B1(n14175), .B2(n14973), .ZN(
        P3_U3429) );
  AOI22_X1 U16006 ( .A1(n14974), .A2(n14177), .B1(n8555), .B2(n14973), .ZN(
        P3_U3426) );
  AOI22_X1 U16007 ( .A1(n14974), .A2(n14178), .B1(n8538), .B2(n14973), .ZN(
        P3_U3423) );
  OAI21_X1 U16008 ( .B1(n14180), .B2(n14715), .A(n14179), .ZN(n14182) );
  AOI211_X1 U16009 ( .C1(n14183), .C2(n14719), .A(n14182), .B(n14181), .ZN(
        n14191) );
  AOI22_X1 U16010 ( .A1(n14737), .A2(n14191), .B1(n7955), .B2(n14735), .ZN(
        P2_U3513) );
  INV_X1 U16011 ( .A(n14688), .ZN(n14707) );
  INV_X1 U16012 ( .A(n14184), .ZN(n14189) );
  OAI21_X1 U16013 ( .B1(n14186), .B2(n14715), .A(n14185), .ZN(n14188) );
  AOI211_X1 U16014 ( .C1(n14707), .C2(n14189), .A(n14188), .B(n14187), .ZN(
        n14193) );
  AOI22_X1 U16015 ( .A1(n14737), .A2(n14193), .B1(n9492), .B2(n14735), .ZN(
        P2_U3511) );
  INV_X1 U16016 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14190) );
  AOI22_X1 U16017 ( .A1(n14723), .A2(n14191), .B1(n14190), .B2(n14721), .ZN(
        P2_U3472) );
  INV_X1 U16018 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14192) );
  AOI22_X1 U16019 ( .A1(n14723), .A2(n14193), .B1(n14192), .B2(n14721), .ZN(
        P2_U3466) );
  OAI22_X1 U16020 ( .A1(n14194), .A2(n14214), .B1(n14215), .B2(n14208), .ZN(
        n14202) );
  INV_X1 U16021 ( .A(n14195), .ZN(n14198) );
  OAI21_X1 U16022 ( .B1(n14198), .B2(n14197), .A(n14196), .ZN(n14200) );
  AOI21_X1 U16023 ( .B1(n14200), .B2(n14199), .A(n14221), .ZN(n14201) );
  AOI211_X1 U16024 ( .C1(n14285), .C2(n14238), .A(n14202), .B(n14201), .ZN(
        n14204) );
  OAI211_X1 U16025 ( .C1(n14241), .C2(n14205), .A(n14204), .B(n14203), .ZN(
        P1_U3215) );
  XNOR2_X1 U16026 ( .A(n14206), .B(n14207), .ZN(n14210) );
  OAI22_X1 U16027 ( .A1(n14209), .A2(n14380), .B1(n14208), .B2(n14382), .ZN(
        n14270) );
  AOI222_X1 U16028 ( .A1(n14238), .A2(n14271), .B1(n14233), .B2(n14210), .C1(
        n14270), .C2(n14235), .ZN(n14212) );
  OAI211_X1 U16029 ( .C1(n14241), .C2(n14244), .A(n14212), .B(n14211), .ZN(
        P1_U3226) );
  OAI22_X1 U16030 ( .A1(n14216), .A2(n14215), .B1(n14214), .B2(n14213), .ZN(
        n14225) );
  AOI21_X1 U16031 ( .B1(n14219), .B2(n14218), .A(n14217), .ZN(n14220) );
  INV_X1 U16032 ( .A(n14220), .ZN(n14223) );
  AOI21_X1 U16033 ( .B1(n14223), .B2(n14222), .A(n14221), .ZN(n14224) );
  AOI211_X1 U16034 ( .C1(n14226), .C2(n14238), .A(n14225), .B(n14224), .ZN(
        n14228) );
  OAI211_X1 U16035 ( .C1(n14241), .C2(n14229), .A(n14228), .B(n14227), .ZN(
        P1_U3236) );
  OAI21_X1 U16036 ( .B1(n14232), .B2(n14231), .A(n14230), .ZN(n14234) );
  AOI222_X1 U16037 ( .A1(n14238), .A2(n14237), .B1(n14236), .B2(n14235), .C1(
        n14234), .C2(n14233), .ZN(n14239) );
  NAND2_X1 U16038 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14363)
         );
  OAI211_X1 U16039 ( .C1(n14241), .C2(n14240), .A(n14239), .B(n14363), .ZN(
        P1_U3241) );
  XNOR2_X1 U16040 ( .A(n14242), .B(n14249), .ZN(n14243) );
  NAND2_X1 U16041 ( .A1(n14243), .A2(n14429), .ZN(n14272) );
  INV_X1 U16042 ( .A(n14244), .ZN(n14245) );
  AOI22_X1 U16043 ( .A1(n14270), .A2(n14420), .B1(n14245), .B2(n14431), .ZN(
        n14246) );
  OAI21_X1 U16044 ( .B1(n11126), .B2(n14420), .A(n14246), .ZN(n14247) );
  AOI21_X1 U16045 ( .B1(n14271), .B2(n14430), .A(n14247), .ZN(n14255) );
  XOR2_X1 U16046 ( .A(n14249), .B(n14248), .Z(n14274) );
  INV_X1 U16047 ( .A(n14274), .ZN(n14253) );
  AOI211_X1 U16048 ( .C1(n14271), .C2(n14251), .A(n14468), .B(n14250), .ZN(
        n14269) );
  AOI22_X1 U16049 ( .A1(n14253), .A2(n14252), .B1(n14436), .B2(n14269), .ZN(
        n14254) );
  OAI211_X1 U16050 ( .C1(n14439), .C2(n14272), .A(n14255), .B(n14254), .ZN(
        P1_U3277) );
  INV_X1 U16051 ( .A(n14256), .ZN(n14261) );
  OAI22_X1 U16052 ( .A1(n14258), .A2(n14468), .B1(n14257), .B2(n14528), .ZN(
        n14260) );
  AOI211_X1 U16053 ( .C1(n14504), .C2(n14261), .A(n14260), .B(n14259), .ZN(
        n14306) );
  AOI22_X1 U16054 ( .A1(n14563), .A2(n14306), .B1(n11562), .B2(n14561), .ZN(
        P1_U3546) );
  INV_X1 U16055 ( .A(n14262), .ZN(n14263) );
  OAI211_X1 U16056 ( .C1(n14265), .C2(n14528), .A(n14264), .B(n14263), .ZN(
        n14267) );
  AOI211_X1 U16057 ( .C1(n14268), .C2(n14544), .A(n14267), .B(n14266), .ZN(
        n14308) );
  AOI22_X1 U16058 ( .A1(n14563), .A2(n14308), .B1(n15023), .B2(n14561), .ZN(
        P1_U3545) );
  AOI211_X1 U16059 ( .C1(n14538), .C2(n14271), .A(n14270), .B(n14269), .ZN(
        n14273) );
  OAI211_X1 U16060 ( .C1(n14489), .C2(n14274), .A(n14273), .B(n14272), .ZN(
        n14275) );
  INV_X1 U16061 ( .A(n14275), .ZN(n14310) );
  AOI22_X1 U16062 ( .A1(n14563), .A2(n14310), .B1(n14276), .B2(n14561), .ZN(
        P1_U3544) );
  OAI21_X1 U16063 ( .B1(n6931), .B2(n14528), .A(n14277), .ZN(n14280) );
  INV_X1 U16064 ( .A(n14278), .ZN(n14279) );
  AOI211_X1 U16065 ( .C1(n14544), .C2(n14281), .A(n14280), .B(n14279), .ZN(
        n14312) );
  INV_X1 U16066 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14282) );
  AOI22_X1 U16067 ( .A1(n14563), .A2(n14312), .B1(n14282), .B2(n14561), .ZN(
        P1_U3543) );
  NAND3_X1 U16068 ( .A1(n14284), .A2(n14283), .A3(n14544), .ZN(n14288) );
  AOI22_X1 U16069 ( .A1(n14286), .A2(n14412), .B1(n14538), .B2(n14285), .ZN(
        n14287) );
  AND2_X1 U16070 ( .A1(n14288), .A2(n14287), .ZN(n14289) );
  AOI22_X1 U16071 ( .A1(n14563), .A2(n14313), .B1(n14291), .B2(n14561), .ZN(
        P1_U3542) );
  OAI211_X1 U16072 ( .C1(n6934), .C2(n14528), .A(n14293), .B(n14292), .ZN(
        n14296) );
  NOR2_X1 U16073 ( .A1(n14294), .A2(n14489), .ZN(n14295) );
  AOI211_X1 U16074 ( .C1(n14297), .C2(n14429), .A(n14296), .B(n14295), .ZN(
        n14315) );
  AOI22_X1 U16075 ( .A1(n14563), .A2(n14315), .B1(n11031), .B2(n14561), .ZN(
        P1_U3541) );
  OAI21_X1 U16076 ( .B1(n14299), .B2(n14528), .A(n14298), .ZN(n14302) );
  INV_X1 U16077 ( .A(n14300), .ZN(n14301) );
  AOI211_X1 U16078 ( .C1(n14303), .C2(n14544), .A(n14302), .B(n14301), .ZN(
        n14317) );
  AOI22_X1 U16079 ( .A1(n14563), .A2(n14317), .B1(n14304), .B2(n14561), .ZN(
        P1_U3539) );
  INV_X1 U16080 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14305) );
  AOI22_X1 U16081 ( .A1(n14546), .A2(n14306), .B1(n14305), .B2(n7230), .ZN(
        P1_U3513) );
  INV_X1 U16082 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14307) );
  AOI22_X1 U16083 ( .A1(n14546), .A2(n14308), .B1(n14307), .B2(n7230), .ZN(
        P1_U3510) );
  INV_X1 U16084 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14309) );
  AOI22_X1 U16085 ( .A1(n14546), .A2(n14310), .B1(n14309), .B2(n7230), .ZN(
        P1_U3507) );
  INV_X1 U16086 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14311) );
  AOI22_X1 U16087 ( .A1(n14546), .A2(n14312), .B1(n14311), .B2(n7230), .ZN(
        P1_U3504) );
  AOI22_X1 U16088 ( .A1(n14546), .A2(n14313), .B1(n11043), .B2(n7230), .ZN(
        P1_U3501) );
  INV_X1 U16089 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14314) );
  AOI22_X1 U16090 ( .A1(n14546), .A2(n14315), .B1(n14314), .B2(n7230), .ZN(
        P1_U3498) );
  INV_X1 U16091 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14316) );
  AOI22_X1 U16092 ( .A1(n14546), .A2(n14317), .B1(n14316), .B2(n7230), .ZN(
        P1_U3492) );
  OAI21_X1 U16093 ( .B1(n14320), .B2(n14319), .A(n14318), .ZN(n14321) );
  XNOR2_X1 U16094 ( .A(n14321), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16095 ( .B1(n14324), .B2(n14323), .A(n14322), .ZN(n14325) );
  XNOR2_X1 U16096 ( .A(n14325), .B(P2_ADDR_REG_12__SCAN_IN), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U16097 ( .B1(n14328), .B2(n14327), .A(n14326), .ZN(n14330) );
  XNOR2_X1 U16098 ( .A(n14330), .B(n14329), .ZN(SUB_1596_U67) );
  AOI21_X1 U16099 ( .B1(n14333), .B2(n14332), .A(n14331), .ZN(n14334) );
  XNOR2_X1 U16100 ( .A(n14334), .B(n14576), .ZN(SUB_1596_U66) );
  OAI21_X1 U16101 ( .B1(n14336), .B2(n6482), .A(n14335), .ZN(n14337) );
  XNOR2_X1 U16102 ( .A(n14337), .B(P2_ADDR_REG_15__SCAN_IN), .ZN(SUB_1596_U65)
         );
  AOI21_X1 U16103 ( .B1(n14340), .B2(n14339), .A(n14338), .ZN(n14341) );
  XNOR2_X1 U16104 ( .A(n14341), .B(n14602), .ZN(SUB_1596_U64) );
  AOI21_X1 U16105 ( .B1(n14344), .B2(n14343), .A(n14342), .ZN(n14345) );
  XNOR2_X1 U16106 ( .A(n14345), .B(P1_IR_REG_0__SCAN_IN), .ZN(n14349) );
  AOI22_X1 U16107 ( .A1(n14346), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14347) );
  OAI21_X1 U16108 ( .B1(n14349), .B2(n14348), .A(n14347), .ZN(P1_U3243) );
  AOI21_X1 U16109 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14351), .A(n14350), 
        .ZN(n14361) );
  AOI21_X1 U16110 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n14353), .A(n14352), 
        .ZN(n14355) );
  OR2_X1 U16111 ( .A1(n14355), .A2(n14354), .ZN(n14359) );
  NAND2_X1 U16112 ( .A1(n14357), .A2(n14356), .ZN(n14358) );
  OAI211_X1 U16113 ( .C1(n14361), .C2(n14360), .A(n14359), .B(n14358), .ZN(
        n14362) );
  INV_X1 U16114 ( .A(n14362), .ZN(n14364) );
  OAI211_X1 U16115 ( .C1(n14365), .C2(n14992), .A(n14364), .B(n14363), .ZN(
        P1_U3258) );
  OAI211_X1 U16116 ( .C1(n14368), .C2(P1_REG1_REG_18__SCAN_IN), .A(n14367), 
        .B(n14366), .ZN(n14373) );
  OAI211_X1 U16117 ( .C1(n14371), .C2(P1_REG2_REG_18__SCAN_IN), .A(n14370), 
        .B(n14369), .ZN(n14372) );
  OAI211_X1 U16118 ( .C1(n14375), .C2(n14374), .A(n14373), .B(n14372), .ZN(
        n14376) );
  INV_X1 U16119 ( .A(n14376), .ZN(n14378) );
  OAI211_X1 U16120 ( .C1(n15019), .C2(n14992), .A(n14378), .B(n14377), .ZN(
        P1_U3261) );
  XNOR2_X1 U16121 ( .A(n14379), .B(n14384), .ZN(n14503) );
  OAI22_X1 U16122 ( .A1(n14383), .A2(n14382), .B1(n14381), .B2(n14380), .ZN(
        n14390) );
  NAND3_X1 U16123 ( .A1(n14386), .A2(n14385), .A3(n14384), .ZN(n14387) );
  AOI21_X1 U16124 ( .B1(n14388), .B2(n14387), .A(n14540), .ZN(n14389) );
  AOI211_X1 U16125 ( .C1(n14532), .C2(n14503), .A(n14390), .B(n14389), .ZN(
        n14500) );
  INV_X1 U16126 ( .A(n14391), .ZN(n14392) );
  AOI222_X1 U16127 ( .A1(n14393), .A2(n14430), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n14439), .C1(n14431), .C2(n14392), .ZN(n14400) );
  INV_X1 U16128 ( .A(n14394), .ZN(n14397) );
  INV_X1 U16129 ( .A(n14395), .ZN(n14396) );
  OAI211_X1 U16130 ( .C1(n14499), .C2(n14397), .A(n14396), .B(n14412), .ZN(
        n14498) );
  INV_X1 U16131 ( .A(n14498), .ZN(n14398) );
  AOI22_X1 U16132 ( .A1(n14503), .A2(n14434), .B1(n14436), .B2(n14398), .ZN(
        n14399) );
  OAI211_X1 U16133 ( .C1(n14439), .C2(n14500), .A(n14400), .B(n14399), .ZN(
        P1_U3287) );
  XNOR2_X1 U16134 ( .A(n14402), .B(n14401), .ZN(n14478) );
  INV_X1 U16135 ( .A(n14403), .ZN(n14407) );
  AND3_X1 U16136 ( .A1(n14422), .A2(n14405), .A3(n14404), .ZN(n14406) );
  OAI21_X1 U16137 ( .B1(n14407), .B2(n14406), .A(n14429), .ZN(n14409) );
  OAI211_X1 U16138 ( .C1(n14478), .C2(n14509), .A(n14409), .B(n14408), .ZN(
        n14481) );
  NOR2_X1 U16139 ( .A1(n14478), .A2(n14410), .ZN(n14419) );
  INV_X1 U16140 ( .A(n14411), .ZN(n14432) );
  OAI211_X1 U16141 ( .C1(n14480), .C2(n14432), .A(n14413), .B(n14412), .ZN(
        n14479) );
  NOR2_X1 U16142 ( .A1(n14479), .A2(n14414), .ZN(n14418) );
  OAI22_X1 U16143 ( .A1(n14416), .A2(P1_REG3_REG_3__SCAN_IN), .B1(n14480), 
        .B2(n14415), .ZN(n14417) );
  NOR4_X1 U16144 ( .A1(n14481), .A2(n14419), .A3(n14418), .A4(n14417), .ZN(
        n14421) );
  AOI22_X1 U16145 ( .A1(n14439), .A2(n9717), .B1(n14421), .B2(n14420), .ZN(
        P1_U3290) );
  OAI21_X1 U16146 ( .B1(n11441), .B2(n14423), .A(n14422), .ZN(n14428) );
  INV_X1 U16147 ( .A(n14424), .ZN(n14427) );
  XNOR2_X1 U16148 ( .A(n14425), .B(n11441), .ZN(n14476) );
  NOR2_X1 U16149 ( .A1(n14476), .A2(n14509), .ZN(n14426) );
  AOI211_X1 U16150 ( .C1(n14429), .C2(n14428), .A(n14427), .B(n14426), .ZN(
        n14475) );
  AOI222_X1 U16151 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n14439), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14431), .C1(n6748), .C2(n14430), .ZN(
        n14438) );
  AOI211_X1 U16152 ( .C1(n6748), .C2(n14433), .A(n14468), .B(n14432), .ZN(
        n14473) );
  INV_X1 U16153 ( .A(n14476), .ZN(n14435) );
  AOI22_X1 U16154 ( .A1(n14436), .A2(n14473), .B1(n14435), .B2(n14434), .ZN(
        n14437) );
  OAI211_X1 U16155 ( .C1(n14439), .C2(n14475), .A(n14438), .B(n14437), .ZN(
        P1_U3291) );
  INV_X1 U16156 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14440) );
  NOR2_X1 U16157 ( .A1(n14467), .A2(n14440), .ZN(P1_U3294) );
  INV_X1 U16158 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14441) );
  NOR2_X1 U16159 ( .A1(n14467), .A2(n14441), .ZN(P1_U3295) );
  INV_X1 U16160 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14442) );
  NOR2_X1 U16161 ( .A1(n14467), .A2(n14442), .ZN(P1_U3296) );
  INV_X1 U16162 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14443) );
  NOR2_X1 U16163 ( .A1(n14467), .A2(n14443), .ZN(P1_U3297) );
  INV_X1 U16164 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14444) );
  NOR2_X1 U16165 ( .A1(n14467), .A2(n14444), .ZN(P1_U3298) );
  INV_X1 U16166 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14445) );
  NOR2_X1 U16167 ( .A1(n14467), .A2(n14445), .ZN(P1_U3299) );
  INV_X1 U16168 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n14446) );
  NOR2_X1 U16169 ( .A1(n14467), .A2(n14446), .ZN(P1_U3300) );
  INV_X1 U16170 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14447) );
  NOR2_X1 U16171 ( .A1(n14467), .A2(n14447), .ZN(P1_U3301) );
  INV_X1 U16172 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14448) );
  NOR2_X1 U16173 ( .A1(n14467), .A2(n14448), .ZN(P1_U3302) );
  INV_X1 U16174 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14449) );
  NOR2_X1 U16175 ( .A1(n14467), .A2(n14449), .ZN(P1_U3303) );
  INV_X1 U16176 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14450) );
  NOR2_X1 U16177 ( .A1(n14467), .A2(n14450), .ZN(P1_U3304) );
  NOR2_X1 U16178 ( .A1(n14467), .A2(n15108), .ZN(P1_U3305) );
  INV_X1 U16179 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14451) );
  NOR2_X1 U16180 ( .A1(n14467), .A2(n14451), .ZN(P1_U3306) );
  NOR2_X1 U16181 ( .A1(n14467), .A2(n15086), .ZN(P1_U3307) );
  INV_X1 U16182 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14452) );
  NOR2_X1 U16183 ( .A1(n14467), .A2(n14452), .ZN(P1_U3308) );
  INV_X1 U16184 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14453) );
  NOR2_X1 U16185 ( .A1(n14467), .A2(n14453), .ZN(P1_U3309) );
  INV_X1 U16186 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14454) );
  NOR2_X1 U16187 ( .A1(n14467), .A2(n14454), .ZN(P1_U3310) );
  INV_X1 U16188 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14455) );
  NOR2_X1 U16189 ( .A1(n14467), .A2(n14455), .ZN(P1_U3311) );
  INV_X1 U16190 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14456) );
  NOR2_X1 U16191 ( .A1(n14467), .A2(n14456), .ZN(P1_U3312) );
  INV_X1 U16192 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14457) );
  NOR2_X1 U16193 ( .A1(n14467), .A2(n14457), .ZN(P1_U3313) );
  INV_X1 U16194 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14458) );
  NOR2_X1 U16195 ( .A1(n14467), .A2(n14458), .ZN(P1_U3314) );
  INV_X1 U16196 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14459) );
  NOR2_X1 U16197 ( .A1(n14467), .A2(n14459), .ZN(P1_U3315) );
  INV_X1 U16198 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14460) );
  NOR2_X1 U16199 ( .A1(n14467), .A2(n14460), .ZN(P1_U3316) );
  NOR2_X1 U16200 ( .A1(n14467), .A2(n15125), .ZN(P1_U3317) );
  INV_X1 U16201 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14461) );
  NOR2_X1 U16202 ( .A1(n14467), .A2(n14461), .ZN(P1_U3318) );
  INV_X1 U16203 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14462) );
  NOR2_X1 U16204 ( .A1(n14467), .A2(n14462), .ZN(P1_U3319) );
  INV_X1 U16205 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14463) );
  NOR2_X1 U16206 ( .A1(n14467), .A2(n14463), .ZN(P1_U3320) );
  INV_X1 U16207 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14464) );
  NOR2_X1 U16208 ( .A1(n14467), .A2(n14464), .ZN(P1_U3321) );
  INV_X1 U16209 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14465) );
  NOR2_X1 U16210 ( .A1(n14467), .A2(n14465), .ZN(P1_U3322) );
  NOR2_X1 U16211 ( .A1(n14467), .A2(n14466), .ZN(P1_U3323) );
  OAI22_X1 U16212 ( .A1(n14469), .A2(n14468), .B1(n9925), .B2(n14528), .ZN(
        n14471) );
  AOI211_X1 U16213 ( .C1(n14504), .C2(n14472), .A(n14471), .B(n14470), .ZN(
        n14547) );
  AOI22_X1 U16214 ( .A1(n14546), .A2(n14547), .B1(n9559), .B2(n7230), .ZN(
        P1_U3462) );
  AOI21_X1 U16215 ( .B1(n14538), .B2(n6748), .A(n14473), .ZN(n14474) );
  OAI211_X1 U16216 ( .C1(n14476), .C2(n14523), .A(n14475), .B(n14474), .ZN(
        n14477) );
  INV_X1 U16217 ( .A(n14477), .ZN(n14548) );
  AOI22_X1 U16218 ( .A1(n14546), .A2(n14548), .B1(n9581), .B2(n7230), .ZN(
        P1_U3465) );
  INV_X1 U16219 ( .A(n14478), .ZN(n14483) );
  OAI21_X1 U16220 ( .B1(n14480), .B2(n14528), .A(n14479), .ZN(n14482) );
  AOI211_X1 U16221 ( .C1(n14504), .C2(n14483), .A(n14482), .B(n14481), .ZN(
        n14549) );
  AOI22_X1 U16222 ( .A1(n14546), .A2(n14549), .B1(n9706), .B2(n7230), .ZN(
        P1_U3468) );
  AOI21_X1 U16223 ( .B1(n14538), .B2(n14485), .A(n14484), .ZN(n14487) );
  OAI211_X1 U16224 ( .C1(n14489), .C2(n14488), .A(n14487), .B(n14486), .ZN(
        n14490) );
  INV_X1 U16225 ( .A(n14490), .ZN(n14550) );
  INV_X1 U16226 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14491) );
  AOI22_X1 U16227 ( .A1(n14546), .A2(n14550), .B1(n14491), .B2(n7230), .ZN(
        P1_U3471) );
  INV_X1 U16228 ( .A(n14492), .ZN(n14497) );
  OAI21_X1 U16229 ( .B1(n14494), .B2(n14528), .A(n14493), .ZN(n14496) );
  AOI211_X1 U16230 ( .C1(n14504), .C2(n14497), .A(n14496), .B(n14495), .ZN(
        n14552) );
  AOI22_X1 U16231 ( .A1(n14546), .A2(n14552), .B1(n10235), .B2(n7230), .ZN(
        P1_U3474) );
  OAI21_X1 U16232 ( .B1(n14499), .B2(n14528), .A(n14498), .ZN(n14502) );
  INV_X1 U16233 ( .A(n14500), .ZN(n14501) );
  AOI211_X1 U16234 ( .C1(n14504), .C2(n14503), .A(n14502), .B(n14501), .ZN(
        n14554) );
  INV_X1 U16235 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14505) );
  AOI22_X1 U16236 ( .A1(n14546), .A2(n14554), .B1(n14505), .B2(n7230), .ZN(
        P1_U3477) );
  AND2_X1 U16237 ( .A1(n14506), .A2(n14538), .ZN(n14507) );
  NOR2_X1 U16238 ( .A1(n14508), .A2(n14507), .ZN(n14513) );
  OR2_X1 U16239 ( .A1(n14510), .A2(n14523), .ZN(n14512) );
  OR2_X1 U16240 ( .A1(n14510), .A2(n14509), .ZN(n14511) );
  AND4_X1 U16241 ( .A1(n14514), .A2(n14513), .A3(n14512), .A4(n14511), .ZN(
        n14556) );
  AOI22_X1 U16242 ( .A1(n14546), .A2(n14556), .B1(n10276), .B2(n7230), .ZN(
        P1_U3480) );
  NAND2_X1 U16243 ( .A1(n14515), .A2(n14538), .ZN(n14516) );
  AND2_X1 U16244 ( .A1(n14517), .A2(n14516), .ZN(n14520) );
  NAND2_X1 U16245 ( .A1(n14518), .A2(n14544), .ZN(n14519) );
  AND3_X1 U16246 ( .A1(n14521), .A2(n14520), .A3(n14519), .ZN(n14558) );
  INV_X1 U16247 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14522) );
  AOI22_X1 U16248 ( .A1(n14546), .A2(n14558), .B1(n14522), .B2(n7230), .ZN(
        P1_U3483) );
  INV_X1 U16249 ( .A(n14524), .ZN(n14533) );
  NOR2_X1 U16250 ( .A1(n14524), .A2(n14523), .ZN(n14531) );
  INV_X1 U16251 ( .A(n14525), .ZN(n14529) );
  OAI211_X1 U16252 ( .C1(n14529), .C2(n14528), .A(n14527), .B(n14526), .ZN(
        n14530) );
  AOI211_X1 U16253 ( .C1(n14533), .C2(n14532), .A(n14531), .B(n14530), .ZN(
        n14560) );
  INV_X1 U16254 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14534) );
  AOI22_X1 U16255 ( .A1(n14546), .A2(n14560), .B1(n14534), .B2(n7230), .ZN(
        P1_U3486) );
  AOI211_X1 U16256 ( .C1(n14538), .C2(n14537), .A(n14536), .B(n14535), .ZN(
        n14539) );
  OAI21_X1 U16257 ( .B1(n14541), .B2(n14540), .A(n14539), .ZN(n14542) );
  AOI21_X1 U16258 ( .B1(n14544), .B2(n14543), .A(n14542), .ZN(n14562) );
  INV_X1 U16259 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14545) );
  AOI22_X1 U16260 ( .A1(n14546), .A2(n14562), .B1(n14545), .B2(n7230), .ZN(
        P1_U3489) );
  AOI22_X1 U16261 ( .A1(n14563), .A2(n14547), .B1(n9732), .B2(n14561), .ZN(
        P1_U3529) );
  AOI22_X1 U16262 ( .A1(n14563), .A2(n14548), .B1(n9731), .B2(n14561), .ZN(
        P1_U3530) );
  AOI22_X1 U16263 ( .A1(n14563), .A2(n14549), .B1(n9733), .B2(n14561), .ZN(
        P1_U3531) );
  AOI22_X1 U16264 ( .A1(n14563), .A2(n14550), .B1(n15068), .B2(n14561), .ZN(
        P1_U3532) );
  AOI22_X1 U16265 ( .A1(n14563), .A2(n14552), .B1(n14551), .B2(n14561), .ZN(
        P1_U3533) );
  AOI22_X1 U16266 ( .A1(n14563), .A2(n14554), .B1(n14553), .B2(n14561), .ZN(
        P1_U3534) );
  AOI22_X1 U16267 ( .A1(n14563), .A2(n14556), .B1(n14555), .B2(n14561), .ZN(
        P1_U3535) );
  AOI22_X1 U16268 ( .A1(n14563), .A2(n14558), .B1(n14557), .B2(n14561), .ZN(
        P1_U3536) );
  AOI22_X1 U16269 ( .A1(n14563), .A2(n14560), .B1(n14559), .B2(n14561), .ZN(
        P1_U3537) );
  AOI22_X1 U16270 ( .A1(n14563), .A2(n14562), .B1(n10553), .B2(n14561), .ZN(
        P1_U3538) );
  NOR2_X1 U16271 ( .A1(n14577), .A2(P2_U3947), .ZN(P2_U3087) );
  XNOR2_X1 U16272 ( .A(n14564), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n14573) );
  AOI21_X1 U16273 ( .B1(n14571), .B2(P2_REG1_REG_14__SCAN_IN), .A(n14565), 
        .ZN(n14566) );
  OAI21_X1 U16274 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n14571), .A(n14566), 
        .ZN(n14568) );
  OAI211_X1 U16275 ( .C1(n14569), .C2(n14568), .A(n14567), .B(n14579), .ZN(
        n14570) );
  OAI21_X1 U16276 ( .B1(n14624), .B2(n14571), .A(n14570), .ZN(n14572) );
  AOI21_X1 U16277 ( .B1(n14573), .B2(n14582), .A(n14572), .ZN(n14575) );
  OAI211_X1 U16278 ( .C1(n14576), .C2(n14628), .A(n14575), .B(n14574), .ZN(
        P2_U3228) );
  AOI22_X1 U16279 ( .A1(n14577), .A2(P2_ADDR_REG_15__SCAN_IN), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(P2_U3088), .ZN(n14589) );
  OAI211_X1 U16280 ( .C1(n14580), .C2(P2_REG1_REG_15__SCAN_IN), .A(n14579), 
        .B(n14578), .ZN(n14588) );
  OAI211_X1 U16281 ( .C1(n14583), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14582), 
        .B(n14581), .ZN(n14587) );
  NAND2_X1 U16282 ( .A1(n14585), .A2(n14584), .ZN(n14586) );
  NAND4_X1 U16283 ( .A1(n14589), .A2(n14588), .A3(n14587), .A4(n14586), .ZN(
        P2_U3229) );
  OAI21_X1 U16284 ( .B1(n14592), .B2(n14591), .A(n14590), .ZN(n14597) );
  OAI21_X1 U16285 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(n14596) );
  OAI222_X1 U16286 ( .A1(n14624), .A2(n14598), .B1(n14622), .B2(n14597), .C1(
        n14620), .C2(n14596), .ZN(n14599) );
  INV_X1 U16287 ( .A(n14599), .ZN(n14601) );
  OAI211_X1 U16288 ( .C1(n14602), .C2(n14628), .A(n14601), .B(n14600), .ZN(
        P2_U3230) );
  OAI21_X1 U16289 ( .B1(n14605), .B2(n14604), .A(n14603), .ZN(n14610) );
  OAI21_X1 U16290 ( .B1(n14608), .B2(n14607), .A(n14606), .ZN(n14609) );
  OAI222_X1 U16291 ( .A1(n14624), .A2(n14611), .B1(n14622), .B2(n14610), .C1(
        n14620), .C2(n14609), .ZN(n14612) );
  INV_X1 U16292 ( .A(n14612), .ZN(n14614) );
  OAI211_X1 U16293 ( .C1(n15033), .C2(n14628), .A(n14614), .B(n14613), .ZN(
        P2_U3231) );
  INV_X1 U16294 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n14629) );
  AOI21_X1 U16295 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n14616), .A(n14615), 
        .ZN(n14621) );
  OAI21_X1 U16296 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n14618), .A(n14617), 
        .ZN(n14619) );
  OAI222_X1 U16297 ( .A1(n14624), .A2(n14623), .B1(n14622), .B2(n14621), .C1(
        n14620), .C2(n14619), .ZN(n14625) );
  INV_X1 U16298 ( .A(n14625), .ZN(n14627) );
  OAI211_X1 U16299 ( .C1(n14629), .C2(n14628), .A(n14627), .B(n14626), .ZN(
        P2_U3232) );
  NOR2_X1 U16300 ( .A1(n14635), .A2(n14630), .ZN(n14631) );
  AND2_X1 U16301 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14632), .ZN(P2_U3266) );
  INV_X1 U16302 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15121) );
  NOR2_X1 U16303 ( .A1(n14631), .A2(n15121), .ZN(P2_U3267) );
  AND2_X1 U16304 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14632), .ZN(P2_U3268) );
  INV_X1 U16305 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15096) );
  NOR2_X1 U16306 ( .A1(n14631), .A2(n15096), .ZN(P2_U3269) );
  AND2_X1 U16307 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14632), .ZN(P2_U3270) );
  AND2_X1 U16308 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14632), .ZN(P2_U3271) );
  AND2_X1 U16309 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14632), .ZN(P2_U3272) );
  AND2_X1 U16310 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14632), .ZN(P2_U3273) );
  AND2_X1 U16311 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14632), .ZN(P2_U3274) );
  AND2_X1 U16312 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14632), .ZN(P2_U3275) );
  AND2_X1 U16313 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14632), .ZN(P2_U3276) );
  AND2_X1 U16314 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14632), .ZN(P2_U3277) );
  AND2_X1 U16315 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14632), .ZN(P2_U3278) );
  AND2_X1 U16316 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14632), .ZN(P2_U3279) );
  AND2_X1 U16317 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14632), .ZN(P2_U3280) );
  INV_X1 U16318 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15087) );
  NOR2_X1 U16319 ( .A1(n14631), .A2(n15087), .ZN(P2_U3281) );
  AND2_X1 U16320 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14632), .ZN(P2_U3282) );
  AND2_X1 U16321 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14632), .ZN(P2_U3283) );
  AND2_X1 U16322 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14632), .ZN(P2_U3284) );
  AND2_X1 U16323 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14632), .ZN(P2_U3285) );
  AND2_X1 U16324 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14632), .ZN(P2_U3286) );
  AND2_X1 U16325 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14632), .ZN(P2_U3287) );
  AND2_X1 U16326 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14632), .ZN(P2_U3288) );
  AND2_X1 U16327 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14632), .ZN(P2_U3289) );
  AND2_X1 U16328 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14632), .ZN(P2_U3290) );
  AND2_X1 U16329 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14632), .ZN(P2_U3291) );
  AND2_X1 U16330 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14632), .ZN(P2_U3292) );
  AND2_X1 U16331 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14632), .ZN(P2_U3293) );
  AND2_X1 U16332 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14632), .ZN(P2_U3294) );
  AND2_X1 U16333 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14632), .ZN(P2_U3295) );
  OAI21_X1 U16334 ( .B1(n14637), .B2(n14634), .A(n14633), .ZN(P2_U3416) );
  AOI22_X1 U16335 ( .A1(n14637), .A2(n14636), .B1(n15046), .B2(n14635), .ZN(
        P2_U3417) );
  INV_X1 U16336 ( .A(n14638), .ZN(n14642) );
  INV_X1 U16337 ( .A(n14639), .ZN(n14640) );
  AOI211_X1 U16338 ( .C1(n14642), .C2(n14707), .A(n14641), .B(n14640), .ZN(
        n14724) );
  INV_X1 U16339 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14643) );
  AOI22_X1 U16340 ( .A1(n14723), .A2(n14724), .B1(n14643), .B2(n14721), .ZN(
        P2_U3430) );
  OAI21_X1 U16341 ( .B1(n14645), .B2(n14715), .A(n14644), .ZN(n14647) );
  AOI211_X1 U16342 ( .C1(n14719), .C2(n14648), .A(n14647), .B(n14646), .ZN(
        n14725) );
  INV_X1 U16343 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14649) );
  AOI22_X1 U16344 ( .A1(n14723), .A2(n14725), .B1(n14649), .B2(n14721), .ZN(
        P2_U3436) );
  AOI21_X1 U16345 ( .B1(n14660), .B2(n14651), .A(n14650), .ZN(n14652) );
  OAI211_X1 U16346 ( .C1(n14655), .C2(n14654), .A(n14653), .B(n14652), .ZN(
        n14656) );
  INV_X1 U16347 ( .A(n14656), .ZN(n14726) );
  INV_X1 U16348 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14657) );
  AOI22_X1 U16349 ( .A1(n14723), .A2(n14726), .B1(n14657), .B2(n14721), .ZN(
        P2_U3439) );
  AOI21_X1 U16350 ( .B1(n14660), .B2(n14659), .A(n14658), .ZN(n14661) );
  OAI211_X1 U16351 ( .C1(n14663), .C2(n14688), .A(n14662), .B(n14661), .ZN(
        n14664) );
  INV_X1 U16352 ( .A(n14664), .ZN(n14727) );
  INV_X1 U16353 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14665) );
  AOI22_X1 U16354 ( .A1(n14723), .A2(n14727), .B1(n14665), .B2(n14721), .ZN(
        P2_U3442) );
  AOI21_X1 U16355 ( .B1(n14689), .B2(n14688), .A(n14666), .ZN(n14672) );
  INV_X1 U16356 ( .A(n14667), .ZN(n14668) );
  OAI211_X1 U16357 ( .C1(n14670), .C2(n14715), .A(n14669), .B(n14668), .ZN(
        n14671) );
  NOR2_X1 U16358 ( .A1(n14672), .A2(n14671), .ZN(n14728) );
  INV_X1 U16359 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14673) );
  AOI22_X1 U16360 ( .A1(n14723), .A2(n14728), .B1(n14673), .B2(n14721), .ZN(
        P2_U3445) );
  INV_X1 U16361 ( .A(n14674), .ZN(n14679) );
  OAI21_X1 U16362 ( .B1(n14676), .B2(n14715), .A(n14675), .ZN(n14678) );
  AOI211_X1 U16363 ( .C1(n14707), .C2(n14679), .A(n14678), .B(n14677), .ZN(
        n14730) );
  INV_X1 U16364 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14680) );
  AOI22_X1 U16365 ( .A1(n14723), .A2(n14730), .B1(n14680), .B2(n14721), .ZN(
        P2_U3448) );
  INV_X1 U16366 ( .A(n14681), .ZN(n14686) );
  OAI211_X1 U16367 ( .C1(n14684), .C2(n14715), .A(n14683), .B(n14682), .ZN(
        n14685) );
  AOI21_X1 U16368 ( .B1(n14686), .B2(n14719), .A(n14685), .ZN(n14731) );
  INV_X1 U16369 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14687) );
  AOI22_X1 U16370 ( .A1(n14723), .A2(n14731), .B1(n14687), .B2(n14721), .ZN(
        P2_U3451) );
  NOR2_X1 U16371 ( .A1(n14690), .A2(n14688), .ZN(n14696) );
  NOR2_X1 U16372 ( .A1(n14690), .A2(n14689), .ZN(n14694) );
  OAI21_X1 U16373 ( .B1(n14692), .B2(n14715), .A(n14691), .ZN(n14693) );
  NOR4_X1 U16374 ( .A1(n14696), .A2(n14695), .A3(n14694), .A4(n14693), .ZN(
        n14732) );
  AOI22_X1 U16375 ( .A1(n14723), .A2(n14732), .B1(n7871), .B2(n14721), .ZN(
        P2_U3454) );
  OAI21_X1 U16376 ( .B1(n6802), .B2(n14715), .A(n14697), .ZN(n14698) );
  AOI21_X1 U16377 ( .B1(n14700), .B2(n14707), .A(n14698), .ZN(n14702) );
  AOI21_X1 U16378 ( .B1(n14700), .B2(n14709), .A(n14699), .ZN(n14701) );
  AND2_X1 U16379 ( .A1(n14702), .A2(n14701), .ZN(n14733) );
  INV_X1 U16380 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n14703) );
  AOI22_X1 U16381 ( .A1(n14723), .A2(n14733), .B1(n14703), .B2(n14721), .ZN(
        P2_U3457) );
  OAI21_X1 U16382 ( .B1(n14705), .B2(n14715), .A(n14704), .ZN(n14706) );
  AOI21_X1 U16383 ( .B1(n14710), .B2(n14707), .A(n14706), .ZN(n14712) );
  AOI21_X1 U16384 ( .B1(n14710), .B2(n14709), .A(n14708), .ZN(n14711) );
  AND2_X1 U16385 ( .A1(n14712), .A2(n14711), .ZN(n14734) );
  INV_X1 U16386 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14713) );
  AOI22_X1 U16387 ( .A1(n14723), .A2(n14734), .B1(n14713), .B2(n14721), .ZN(
        P2_U3460) );
  OAI21_X1 U16388 ( .B1(n14716), .B2(n14715), .A(n14714), .ZN(n14718) );
  AOI211_X1 U16389 ( .C1(n14720), .C2(n14719), .A(n14718), .B(n14717), .ZN(
        n14736) );
  INV_X1 U16390 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14722) );
  AOI22_X1 U16391 ( .A1(n14723), .A2(n14736), .B1(n14722), .B2(n14721), .ZN(
        P2_U3463) );
  AOI22_X1 U16392 ( .A1(n14737), .A2(n14724), .B1(n9836), .B2(n14735), .ZN(
        P2_U3499) );
  AOI22_X1 U16393 ( .A1(n14737), .A2(n14725), .B1(n9464), .B2(n14735), .ZN(
        P2_U3501) );
  AOI22_X1 U16394 ( .A1(n14737), .A2(n14726), .B1(n9466), .B2(n14735), .ZN(
        P2_U3502) );
  AOI22_X1 U16395 ( .A1(n14737), .A2(n14727), .B1(n9469), .B2(n14735), .ZN(
        P2_U3503) );
  AOI22_X1 U16396 ( .A1(n14737), .A2(n14728), .B1(n9472), .B2(n14735), .ZN(
        P2_U3504) );
  AOI22_X1 U16397 ( .A1(n14737), .A2(n14730), .B1(n14729), .B2(n14735), .ZN(
        P2_U3505) );
  AOI22_X1 U16398 ( .A1(n14737), .A2(n14731), .B1(n9477), .B2(n14735), .ZN(
        P2_U3506) );
  AOI22_X1 U16399 ( .A1(n14737), .A2(n14732), .B1(n9480), .B2(n14735), .ZN(
        P2_U3507) );
  AOI22_X1 U16400 ( .A1(n14737), .A2(n14733), .B1(n9518), .B2(n14735), .ZN(
        P2_U3508) );
  AOI22_X1 U16401 ( .A1(n14737), .A2(n14734), .B1(n9487), .B2(n14735), .ZN(
        P2_U3509) );
  AOI22_X1 U16402 ( .A1(n14737), .A2(n14736), .B1(n9488), .B2(n14735), .ZN(
        P2_U3510) );
  NOR2_X1 U16403 ( .A1(P3_U3897), .A2(n14871), .ZN(P3_U3150) );
  MUX2_X1 U16404 ( .A(n14739), .B(n11803), .S(n14738), .Z(n14740) );
  NOR2_X1 U16405 ( .A1(n14740), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14743) );
  NAND3_X1 U16406 ( .A1(n14878), .A2(n14741), .A3(n14761), .ZN(n14742) );
  OAI21_X1 U16407 ( .B1(n14744), .B2(n14743), .A(n14742), .ZN(n14749) );
  INV_X1 U16408 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n14745) );
  OAI22_X1 U16409 ( .A1(n14868), .A2(n14746), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14745), .ZN(n14747) );
  INV_X1 U16410 ( .A(n14747), .ZN(n14748) );
  OAI211_X1 U16411 ( .C1(n14750), .C2(n14837), .A(n14749), .B(n14748), .ZN(
        P3_U3182) );
  AOI21_X1 U16412 ( .B1(n14752), .B2(n10852), .A(n14751), .ZN(n14757) );
  OAI21_X1 U16413 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n14754), .A(n14753), .ZN(
        n14755) );
  NAND2_X1 U16414 ( .A1(n14874), .A2(n14755), .ZN(n14756) );
  OAI21_X1 U16415 ( .B1(n14757), .B2(n14878), .A(n14756), .ZN(n14764) );
  OR3_X1 U16416 ( .A1(n14760), .A2(n14759), .A3(n14758), .ZN(n14762) );
  AOI21_X1 U16417 ( .B1(n14772), .B2(n14762), .A(n14761), .ZN(n14763) );
  AOI211_X1 U16418 ( .C1(n14828), .C2(n14765), .A(n14764), .B(n14763), .ZN(
        n14767) );
  OAI211_X1 U16419 ( .C1(n7079), .C2(n14837), .A(n14767), .B(n14766), .ZN(
        P3_U3185) );
  AOI21_X1 U16420 ( .B1(n6588), .B2(n14769), .A(n14768), .ZN(n14784) );
  AND3_X1 U16421 ( .A1(n14772), .A2(n14771), .A3(n14770), .ZN(n14773) );
  OAI21_X1 U16422 ( .B1(n14789), .B2(n14773), .A(n14863), .ZN(n14774) );
  OAI21_X1 U16423 ( .B1(n14868), .B2(n14775), .A(n14774), .ZN(n14776) );
  AOI211_X1 U16424 ( .C1(P3_ADDR_REG_4__SCAN_IN), .C2(n14871), .A(n14777), .B(
        n14776), .ZN(n14783) );
  OAI21_X1 U16425 ( .B1(n14780), .B2(n14779), .A(n14778), .ZN(n14781) );
  NAND2_X1 U16426 ( .A1(n14874), .A2(n14781), .ZN(n14782) );
  OAI211_X1 U16427 ( .C1(n14784), .C2(n14878), .A(n14783), .B(n14782), .ZN(
        P3_U3186) );
  AOI21_X1 U16428 ( .B1(n10862), .B2(n14786), .A(n14785), .ZN(n14801) );
  INV_X1 U16429 ( .A(n14806), .ZN(n14791) );
  NOR3_X1 U16430 ( .A1(n14789), .A2(n14788), .A3(n14787), .ZN(n14790) );
  OAI21_X1 U16431 ( .B1(n14791), .B2(n14790), .A(n14863), .ZN(n14792) );
  OAI21_X1 U16432 ( .B1(n14868), .B2(n14793), .A(n14792), .ZN(n14794) );
  AOI211_X1 U16433 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n14871), .A(n14795), .B(
        n14794), .ZN(n14800) );
  OAI21_X1 U16434 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n14797), .A(n14796), .ZN(
        n14798) );
  NAND2_X1 U16435 ( .A1(n14874), .A2(n14798), .ZN(n14799) );
  OAI211_X1 U16436 ( .C1(n14801), .C2(n14878), .A(n14800), .B(n14799), .ZN(
        P3_U3187) );
  AOI21_X1 U16437 ( .B1(n6587), .B2(n14803), .A(n14802), .ZN(n14818) );
  AND3_X1 U16438 ( .A1(n14806), .A2(n14805), .A3(n14804), .ZN(n14807) );
  OAI21_X1 U16439 ( .B1(n14823), .B2(n14807), .A(n14863), .ZN(n14808) );
  OAI21_X1 U16440 ( .B1(n14868), .B2(n14809), .A(n14808), .ZN(n14810) );
  AOI211_X1 U16441 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n14871), .A(n14811), .B(
        n14810), .ZN(n14817) );
  OAI21_X1 U16442 ( .B1(n14814), .B2(n14813), .A(n14812), .ZN(n14815) );
  NAND2_X1 U16443 ( .A1(n14874), .A2(n14815), .ZN(n14816) );
  OAI211_X1 U16444 ( .C1(n14818), .C2(n14878), .A(n14817), .B(n14816), .ZN(
        P3_U3188) );
  AOI21_X1 U16445 ( .B1(n14820), .B2(n10872), .A(n14819), .ZN(n14833) );
  INV_X1 U16446 ( .A(n14844), .ZN(n14825) );
  NOR3_X1 U16447 ( .A1(n14823), .A2(n14822), .A3(n14821), .ZN(n14824) );
  OAI21_X1 U16448 ( .B1(n14825), .B2(n14824), .A(n14863), .ZN(n14832) );
  OAI21_X1 U16449 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n14827), .A(n14826), .ZN(
        n14830) );
  AOI22_X1 U16450 ( .A1(n14830), .A2(n14874), .B1(n14829), .B2(n14828), .ZN(
        n14831) );
  OAI211_X1 U16451 ( .C1(n14833), .C2(n14878), .A(n14832), .B(n14831), .ZN(
        n14834) );
  INV_X1 U16452 ( .A(n14834), .ZN(n14836) );
  OAI211_X1 U16453 ( .C1(n14838), .C2(n14837), .A(n14836), .B(n14835), .ZN(
        P3_U3189) );
  AOI21_X1 U16454 ( .B1(n14841), .B2(n14840), .A(n14839), .ZN(n14856) );
  AND3_X1 U16455 ( .A1(n14844), .A2(n14843), .A3(n14842), .ZN(n14845) );
  OAI21_X1 U16456 ( .B1(n14862), .B2(n14845), .A(n14863), .ZN(n14846) );
  OAI21_X1 U16457 ( .B1(n14868), .B2(n14847), .A(n14846), .ZN(n14848) );
  AOI211_X1 U16458 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n14871), .A(n14849), .B(
        n14848), .ZN(n14855) );
  OAI21_X1 U16459 ( .B1(n14852), .B2(n14851), .A(n14850), .ZN(n14853) );
  NAND2_X1 U16460 ( .A1(n14853), .A2(n14874), .ZN(n14854) );
  OAI211_X1 U16461 ( .C1(n14856), .C2(n14878), .A(n14855), .B(n14854), .ZN(
        P3_U3190) );
  AOI21_X1 U16462 ( .B1(n11272), .B2(n14858), .A(n14857), .ZN(n14879) );
  INV_X1 U16463 ( .A(n14859), .ZN(n14865) );
  NOR3_X1 U16464 ( .A1(n14862), .A2(n14861), .A3(n14860), .ZN(n14864) );
  OAI21_X1 U16465 ( .B1(n14865), .B2(n14864), .A(n14863), .ZN(n14866) );
  OAI21_X1 U16466 ( .B1(n14868), .B2(n14867), .A(n14866), .ZN(n14869) );
  AOI211_X1 U16467 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n14871), .A(n14870), .B(
        n14869), .ZN(n14877) );
  OAI21_X1 U16468 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n14873), .A(n14872), .ZN(
        n14875) );
  NAND2_X1 U16469 ( .A1(n14875), .A2(n14874), .ZN(n14876) );
  OAI211_X1 U16470 ( .C1(n14879), .C2(n14878), .A(n14877), .B(n14876), .ZN(
        P3_U3191) );
  XNOR2_X1 U16471 ( .A(n14880), .B(n14886), .ZN(n14967) );
  NAND2_X1 U16472 ( .A1(n14882), .A2(n14881), .ZN(n14884) );
  NAND2_X1 U16473 ( .A1(n14884), .A2(n14883), .ZN(n14885) );
  XOR2_X1 U16474 ( .A(n14886), .B(n14885), .Z(n14892) );
  AOI22_X1 U16475 ( .A1(n14888), .A2(n14919), .B1(n14920), .B2(n14887), .ZN(
        n14890) );
  NAND2_X1 U16476 ( .A1(n14967), .A2(n14906), .ZN(n14889) );
  OAI211_X1 U16477 ( .C1(n14892), .C2(n14891), .A(n14890), .B(n14889), .ZN(
        n14965) );
  AOI21_X1 U16478 ( .B1(n14893), .B2(n14967), .A(n14965), .ZN(n14898) );
  NOR2_X1 U16479 ( .A1(n14894), .A2(n14915), .ZN(n14966) );
  AOI22_X1 U16480 ( .A1(n14896), .A2(n14966), .B1(n14929), .B2(n14895), .ZN(
        n14897) );
  OAI221_X1 U16481 ( .B1(n14935), .B2(n14898), .C1(n14933), .C2(n10903), .A(
        n14897), .ZN(P3_U3225) );
  OAI21_X1 U16482 ( .B1(n14900), .B2(n14905), .A(n14899), .ZN(n14909) );
  OAI22_X1 U16483 ( .A1(n9066), .A2(n14903), .B1(n14902), .B2(n14901), .ZN(
        n14908) );
  XNOR2_X1 U16484 ( .A(n14904), .B(n14905), .ZN(n14912) );
  INV_X1 U16485 ( .A(n14906), .ZN(n14927) );
  NOR2_X1 U16486 ( .A1(n14912), .A2(n14927), .ZN(n14907) );
  AOI211_X1 U16487 ( .C1(n14923), .C2(n14909), .A(n14908), .B(n14907), .ZN(
        n14939) );
  NOR2_X1 U16488 ( .A1(n14910), .A2(n14915), .ZN(n14941) );
  AOI22_X1 U16489 ( .A1(n14941), .A2(n7109), .B1(P3_REG3_REG_2__SCAN_IN), .B2(
        n14929), .ZN(n14914) );
  INV_X1 U16490 ( .A(n14912), .ZN(n14942) );
  AOI22_X1 U16491 ( .A1(n14942), .A2(n14930), .B1(P3_REG2_REG_2__SCAN_IN), 
        .B2(n14935), .ZN(n14913) );
  OAI221_X1 U16492 ( .B1(n14935), .B2(n14939), .C1(n14935), .C2(n14914), .A(
        n14913), .ZN(P3_U3231) );
  NOR2_X1 U16493 ( .A1(n14916), .A2(n14915), .ZN(n14937) );
  XNOR2_X1 U16494 ( .A(n8982), .B(n14917), .ZN(n14928) );
  AOI22_X1 U16495 ( .A1(n14921), .A2(n14920), .B1(n14919), .B2(n14918), .ZN(
        n14926) );
  XNOR2_X1 U16496 ( .A(n8982), .B(n14922), .ZN(n14924) );
  NAND2_X1 U16497 ( .A1(n14924), .A2(n14923), .ZN(n14925) );
  OAI211_X1 U16498 ( .C1(n14928), .C2(n14927), .A(n14926), .B(n14925), .ZN(
        n14936) );
  AOI21_X1 U16499 ( .B1(n14937), .B2(n7109), .A(n14936), .ZN(n14934) );
  INV_X1 U16500 ( .A(n14928), .ZN(n14938) );
  AOI22_X1 U16501 ( .A1(n14930), .A2(n14938), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n14929), .ZN(n14931) );
  OAI221_X1 U16502 ( .B1(n14935), .B2(n14934), .C1(n14933), .C2(n14932), .A(
        n14931), .ZN(P3_U3232) );
  AOI211_X1 U16503 ( .C1(n14968), .C2(n14938), .A(n14937), .B(n14936), .ZN(
        n14976) );
  AOI22_X1 U16504 ( .A1(n14974), .A2(n14976), .B1(n8391), .B2(n14973), .ZN(
        P3_U3393) );
  INV_X1 U16505 ( .A(n14939), .ZN(n14940) );
  AOI211_X1 U16506 ( .C1(n14942), .C2(n14968), .A(n14941), .B(n14940), .ZN(
        n14977) );
  AOI22_X1 U16507 ( .A1(n14974), .A2(n14977), .B1(n8368), .B2(n14973), .ZN(
        P3_U3396) );
  INV_X1 U16508 ( .A(n14943), .ZN(n14945) );
  AOI211_X1 U16509 ( .C1(n14968), .C2(n14946), .A(n14945), .B(n14944), .ZN(
        n14978) );
  AOI22_X1 U16510 ( .A1(n14974), .A2(n14978), .B1(n8406), .B2(n14973), .ZN(
        P3_U3399) );
  INV_X1 U16511 ( .A(n14947), .ZN(n14948) );
  AOI211_X1 U16512 ( .C1(n14950), .C2(n14968), .A(n14949), .B(n14948), .ZN(
        n14980) );
  AOI22_X1 U16513 ( .A1(n14974), .A2(n14980), .B1(n8423), .B2(n14973), .ZN(
        P3_U3402) );
  AOI21_X1 U16514 ( .B1(n14952), .B2(n14968), .A(n14951), .ZN(n14953) );
  AND2_X1 U16515 ( .A1(n14954), .A2(n14953), .ZN(n14981) );
  AOI22_X1 U16516 ( .A1(n14974), .A2(n14981), .B1(n8441), .B2(n14973), .ZN(
        P3_U3405) );
  INV_X1 U16517 ( .A(n14955), .ZN(n14956) );
  AOI211_X1 U16518 ( .C1(n14968), .C2(n14958), .A(n14957), .B(n14956), .ZN(
        n14983) );
  AOI22_X1 U16519 ( .A1(n14974), .A2(n14983), .B1(n8455), .B2(n14973), .ZN(
        P3_U3408) );
  AND2_X1 U16520 ( .A1(n14959), .A2(n14968), .ZN(n14963) );
  AND2_X1 U16521 ( .A1(n14961), .A2(n14960), .ZN(n14962) );
  NOR3_X1 U16522 ( .A1(n14964), .A2(n14963), .A3(n14962), .ZN(n14984) );
  AOI22_X1 U16523 ( .A1(n14974), .A2(n14984), .B1(n8468), .B2(n14973), .ZN(
        P3_U3411) );
  AOI211_X1 U16524 ( .C1(n14968), .C2(n14967), .A(n14966), .B(n14965), .ZN(
        n14986) );
  AOI22_X1 U16525 ( .A1(n14974), .A2(n14986), .B1(n8485), .B2(n14973), .ZN(
        P3_U3414) );
  AOI211_X1 U16526 ( .C1(n14972), .C2(n14971), .A(n14970), .B(n14969), .ZN(
        n14989) );
  AOI22_X1 U16527 ( .A1(n14974), .A2(n14989), .B1(n8520), .B2(n14973), .ZN(
        P3_U3420) );
  INV_X1 U16528 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n14975) );
  AOI22_X1 U16529 ( .A1(n14990), .A2(n14976), .B1(n14975), .B2(n14987), .ZN(
        P3_U3460) );
  AOI22_X1 U16530 ( .A1(n14990), .A2(n14977), .B1(n15112), .B2(n14987), .ZN(
        P3_U3461) );
  AOI22_X1 U16531 ( .A1(n14990), .A2(n14978), .B1(n10851), .B2(n14987), .ZN(
        P3_U3462) );
  AOI22_X1 U16532 ( .A1(n14990), .A2(n14980), .B1(n14979), .B2(n14987), .ZN(
        P3_U3463) );
  AOI22_X1 U16533 ( .A1(n14990), .A2(n14981), .B1(n10861), .B2(n14987), .ZN(
        P3_U3464) );
  AOI22_X1 U16534 ( .A1(n14990), .A2(n14983), .B1(n14982), .B2(n14987), .ZN(
        P3_U3465) );
  AOI22_X1 U16535 ( .A1(n14990), .A2(n14984), .B1(n10871), .B2(n14987), .ZN(
        P3_U3466) );
  AOI22_X1 U16536 ( .A1(n14990), .A2(n14986), .B1(n14985), .B2(n14987), .ZN(
        P3_U3467) );
  AOI22_X1 U16537 ( .A1(n14990), .A2(n14989), .B1(n14988), .B2(n14987), .ZN(
        P3_U3469) );
  NAND2_X1 U16538 ( .A1(n14992), .A2(n14991), .ZN(n15141) );
  NAND2_X1 U16539 ( .A1(keyinput30), .A2(keyinput29), .ZN(n14993) );
  NOR3_X1 U16540 ( .A1(keyinput43), .A2(keyinput23), .A3(n14993), .ZN(n14998)
         );
  NOR3_X1 U16541 ( .A1(keyinput61), .A2(keyinput42), .A3(keyinput18), .ZN(
        n14997) );
  NAND4_X1 U16542 ( .A1(keyinput51), .A2(keyinput39), .A3(keyinput57), .A4(
        keyinput37), .ZN(n14995) );
  NAND2_X1 U16543 ( .A1(keyinput28), .A2(keyinput36), .ZN(n14994) );
  NOR4_X1 U16544 ( .A1(keyinput1), .A2(keyinput33), .A3(n14995), .A4(n14994), 
        .ZN(n14996) );
  NAND4_X1 U16545 ( .A1(n14998), .A2(keyinput63), .A3(n14997), .A4(n14996), 
        .ZN(n15005) );
  NOR2_X1 U16546 ( .A1(keyinput17), .A2(keyinput55), .ZN(n14999) );
  NAND3_X1 U16547 ( .A1(keyinput49), .A2(keyinput22), .A3(n14999), .ZN(n15004)
         );
  NAND4_X1 U16548 ( .A1(keyinput50), .A2(keyinput47), .A3(keyinput15), .A4(
        keyinput16), .ZN(n15003) );
  NOR3_X1 U16549 ( .A1(keyinput59), .A2(keyinput5), .A3(keyinput0), .ZN(n15001) );
  NOR3_X1 U16550 ( .A1(keyinput41), .A2(keyinput31), .A3(keyinput38), .ZN(
        n15000) );
  NAND4_X1 U16551 ( .A1(keyinput44), .A2(n15001), .A3(keyinput54), .A4(n15000), 
        .ZN(n15002) );
  NOR4_X1 U16552 ( .A1(n15005), .A2(n15004), .A3(n15003), .A4(n15002), .ZN(
        n15139) );
  NAND4_X1 U16553 ( .A1(keyinput11), .A2(keyinput4), .A3(keyinput26), .A4(
        keyinput19), .ZN(n15017) );
  NOR3_X1 U16554 ( .A1(keyinput21), .A2(keyinput14), .A3(keyinput45), .ZN(
        n15009) );
  NAND3_X1 U16555 ( .A1(keyinput25), .A2(keyinput10), .A3(keyinput27), .ZN(
        n15007) );
  NAND3_X1 U16556 ( .A1(keyinput2), .A2(keyinput40), .A3(keyinput24), .ZN(
        n15006) );
  NOR4_X1 U16557 ( .A1(keyinput35), .A2(keyinput9), .A3(n15007), .A4(n15006), 
        .ZN(n15008) );
  NAND3_X1 U16558 ( .A1(keyinput34), .A2(n15009), .A3(n15008), .ZN(n15016) );
  NAND4_X1 U16559 ( .A1(keyinput48), .A2(keyinput7), .A3(keyinput62), .A4(
        keyinput3), .ZN(n15015) );
  NOR2_X1 U16560 ( .A1(keyinput8), .A2(keyinput6), .ZN(n15013) );
  NAND3_X1 U16561 ( .A1(keyinput56), .A2(keyinput13), .A3(keyinput60), .ZN(
        n15011) );
  NAND3_X1 U16562 ( .A1(keyinput20), .A2(keyinput58), .A3(keyinput53), .ZN(
        n15010) );
  NOR4_X1 U16563 ( .A1(keyinput52), .A2(keyinput46), .A3(n15011), .A4(n15010), 
        .ZN(n15012) );
  NAND4_X1 U16564 ( .A1(keyinput12), .A2(keyinput32), .A3(n15013), .A4(n15012), 
        .ZN(n15014) );
  NOR4_X1 U16565 ( .A1(n15017), .A2(n15016), .A3(n15015), .A4(n15014), .ZN(
        n15138) );
  AOI22_X1 U16566 ( .A1(n15020), .A2(keyinput34), .B1(keyinput21), .B2(n15019), 
        .ZN(n15018) );
  OAI221_X1 U16567 ( .B1(n15020), .B2(keyinput34), .C1(n15019), .C2(keyinput21), .A(n15018), .ZN(n15031) );
  AOI22_X1 U16568 ( .A1(n15023), .A2(keyinput14), .B1(n15022), .B2(keyinput45), 
        .ZN(n15021) );
  OAI221_X1 U16569 ( .B1(n15023), .B2(keyinput14), .C1(n15022), .C2(keyinput45), .A(n15021), .ZN(n15030) );
  AOI22_X1 U16570 ( .A1(n15025), .A2(keyinput25), .B1(keyinput35), .B2(n7294), 
        .ZN(n15024) );
  OAI221_X1 U16571 ( .B1(n15025), .B2(keyinput25), .C1(n7294), .C2(keyinput35), 
        .A(n15024), .ZN(n15029) );
  AOI22_X1 U16572 ( .A1(n15027), .A2(keyinput10), .B1(n8745), .B2(keyinput27), 
        .ZN(n15026) );
  OAI221_X1 U16573 ( .B1(n15027), .B2(keyinput10), .C1(n8745), .C2(keyinput27), 
        .A(n15026), .ZN(n15028) );
  NOR4_X1 U16574 ( .A1(n15031), .A2(n15030), .A3(n15029), .A4(n15028), .ZN(
        n15076) );
  AOI22_X1 U16575 ( .A1(n9715), .A2(keyinput2), .B1(keyinput40), .B2(n15033), 
        .ZN(n15032) );
  OAI221_X1 U16576 ( .B1(n9715), .B2(keyinput2), .C1(n15033), .C2(keyinput40), 
        .A(n15032), .ZN(n15044) );
  AOI22_X1 U16577 ( .A1(n9567), .A2(keyinput9), .B1(n15035), .B2(keyinput24), 
        .ZN(n15034) );
  OAI221_X1 U16578 ( .B1(n9567), .B2(keyinput9), .C1(n15035), .C2(keyinput24), 
        .A(n15034), .ZN(n15043) );
  AOI22_X1 U16579 ( .A1(n15038), .A2(keyinput11), .B1(keyinput4), .B2(n15037), 
        .ZN(n15036) );
  OAI221_X1 U16580 ( .B1(n15038), .B2(keyinput11), .C1(n15037), .C2(keyinput4), 
        .A(n15036), .ZN(n15042) );
  AOI22_X1 U16581 ( .A1(n10729), .A2(keyinput26), .B1(keyinput19), .B2(n15040), 
        .ZN(n15039) );
  OAI221_X1 U16582 ( .B1(n10729), .B2(keyinput26), .C1(n15040), .C2(keyinput19), .A(n15039), .ZN(n15041) );
  NOR4_X1 U16583 ( .A1(n15044), .A2(n15043), .A3(n15042), .A4(n15041), .ZN(
        n15075) );
  AOI22_X1 U16584 ( .A1(n15046), .A2(keyinput62), .B1(keyinput3), .B2(n13775), 
        .ZN(n15045) );
  OAI221_X1 U16585 ( .B1(n15046), .B2(keyinput62), .C1(n13775), .C2(keyinput3), 
        .A(n15045), .ZN(n15058) );
  AOI22_X1 U16586 ( .A1(n15049), .A2(keyinput12), .B1(n15048), .B2(keyinput32), 
        .ZN(n15047) );
  OAI221_X1 U16587 ( .B1(n15049), .B2(keyinput12), .C1(n15048), .C2(keyinput32), .A(n15047), .ZN(n15057) );
  AOI22_X1 U16588 ( .A1(n15052), .A2(keyinput48), .B1(n15051), .B2(keyinput7), 
        .ZN(n15050) );
  OAI221_X1 U16589 ( .B1(n15052), .B2(keyinput48), .C1(n15051), .C2(keyinput7), 
        .A(n15050), .ZN(n15056) );
  XOR2_X1 U16590 ( .A(n9965), .B(keyinput8), .Z(n15054) );
  XNOR2_X1 U16591 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput6), .ZN(n15053) );
  NAND2_X1 U16592 ( .A1(n15054), .A2(n15053), .ZN(n15055) );
  NOR4_X1 U16593 ( .A1(n15058), .A2(n15057), .A3(n15056), .A4(n15055), .ZN(
        n15074) );
  INV_X1 U16594 ( .A(SI_31_), .ZN(n15060) );
  AOI22_X1 U16595 ( .A1(n15061), .A2(keyinput56), .B1(n15060), .B2(keyinput52), 
        .ZN(n15059) );
  OAI221_X1 U16596 ( .B1(n15061), .B2(keyinput56), .C1(n15060), .C2(keyinput52), .A(n15059), .ZN(n15072) );
  INV_X1 U16597 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15064) );
  INV_X1 U16598 ( .A(keyinput13), .ZN(n15063) );
  AOI22_X1 U16599 ( .A1(n15064), .A2(keyinput60), .B1(P2_WR_REG_SCAN_IN), .B2(
        n15063), .ZN(n15062) );
  OAI221_X1 U16600 ( .B1(n15064), .B2(keyinput60), .C1(n15063), .C2(
        P2_WR_REG_SCAN_IN), .A(n15062), .ZN(n15071) );
  AOI22_X1 U16601 ( .A1(n11043), .A2(keyinput20), .B1(keyinput46), .B2(n15066), 
        .ZN(n15065) );
  OAI221_X1 U16602 ( .B1(n11043), .B2(keyinput20), .C1(n15066), .C2(keyinput46), .A(n15065), .ZN(n15070) );
  AOI22_X1 U16603 ( .A1(n15068), .A2(keyinput58), .B1(n7674), .B2(keyinput53), 
        .ZN(n15067) );
  OAI221_X1 U16604 ( .B1(n15068), .B2(keyinput58), .C1(n7674), .C2(keyinput53), 
        .A(n15067), .ZN(n15069) );
  NOR4_X1 U16605 ( .A1(n15072), .A2(n15071), .A3(n15070), .A4(n15069), .ZN(
        n15073) );
  NAND4_X1 U16606 ( .A1(n15076), .A2(n15075), .A3(n15074), .A4(n15073), .ZN(
        n15137) );
  INV_X1 U16607 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n15078) );
  AOI22_X1 U16608 ( .A1(n15079), .A2(keyinput33), .B1(keyinput28), .B2(n15078), 
        .ZN(n15077) );
  OAI221_X1 U16609 ( .B1(n15079), .B2(keyinput33), .C1(n15078), .C2(keyinput28), .A(n15077), .ZN(n15084) );
  XOR2_X1 U16610 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput1), .Z(n15083) );
  XOR2_X1 U16611 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput39), .Z(n15082) );
  XNOR2_X1 U16612 ( .A(n15080), .B(keyinput57), .ZN(n15081) );
  OR4_X1 U16613 ( .A1(n15084), .A2(n15083), .A3(n15082), .A4(n15081), .ZN(
        n15091) );
  INV_X1 U16614 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n15085) );
  XNOR2_X1 U16615 ( .A(n15085), .B(keyinput36), .ZN(n15090) );
  XNOR2_X1 U16616 ( .A(n15086), .B(keyinput37), .ZN(n15089) );
  XNOR2_X1 U16617 ( .A(n15087), .B(keyinput51), .ZN(n15088) );
  NOR4_X1 U16618 ( .A1(n15091), .A2(n15090), .A3(n15089), .A4(n15088), .ZN(
        n15135) );
  AOI22_X1 U16619 ( .A1(n15094), .A2(keyinput29), .B1(keyinput30), .B2(n15093), 
        .ZN(n15092) );
  OAI221_X1 U16620 ( .B1(n15094), .B2(keyinput29), .C1(n15093), .C2(keyinput30), .A(n15092), .ZN(n15106) );
  AOI22_X1 U16621 ( .A1(n15097), .A2(keyinput43), .B1(keyinput23), .B2(n15096), 
        .ZN(n15095) );
  OAI221_X1 U16622 ( .B1(n15097), .B2(keyinput43), .C1(n15096), .C2(keyinput23), .A(n15095), .ZN(n15105) );
  INV_X1 U16623 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n15100) );
  INV_X1 U16624 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n15099) );
  AOI22_X1 U16625 ( .A1(n15100), .A2(keyinput42), .B1(n15099), .B2(keyinput18), 
        .ZN(n15098) );
  OAI221_X1 U16626 ( .B1(n15100), .B2(keyinput42), .C1(n15099), .C2(keyinput18), .A(n15098), .ZN(n15104) );
  AOI22_X1 U16627 ( .A1(n7077), .A2(keyinput63), .B1(n15102), .B2(keyinput61), 
        .ZN(n15101) );
  OAI221_X1 U16628 ( .B1(n7077), .B2(keyinput63), .C1(n15102), .C2(keyinput61), 
        .A(n15101), .ZN(n15103) );
  NOR4_X1 U16629 ( .A1(n15106), .A2(n15105), .A3(n15104), .A4(n15103), .ZN(
        n15134) );
  AOI22_X1 U16630 ( .A1(n15109), .A2(keyinput41), .B1(n15108), .B2(keyinput31), 
        .ZN(n15107) );
  OAI221_X1 U16631 ( .B1(n15109), .B2(keyinput41), .C1(n15108), .C2(keyinput31), .A(n15107), .ZN(n15118) );
  AOI22_X1 U16632 ( .A1(n12273), .A2(keyinput50), .B1(keyinput47), .B2(n7685), 
        .ZN(n15110) );
  OAI221_X1 U16633 ( .B1(n12273), .B2(keyinput50), .C1(n7685), .C2(keyinput47), 
        .A(n15110), .ZN(n15117) );
  AOI22_X1 U16634 ( .A1(n7666), .A2(keyinput15), .B1(n15112), .B2(keyinput16), 
        .ZN(n15111) );
  OAI221_X1 U16635 ( .B1(n7666), .B2(keyinput15), .C1(n15112), .C2(keyinput16), 
        .A(n15111), .ZN(n15116) );
  XNOR2_X1 U16636 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput38), .ZN(n15114) );
  XNOR2_X1 U16637 ( .A(SI_4_), .B(keyinput54), .ZN(n15113) );
  NAND2_X1 U16638 ( .A1(n15114), .A2(n15113), .ZN(n15115) );
  NOR4_X1 U16639 ( .A1(n15118), .A2(n15117), .A3(n15116), .A4(n15115), .ZN(
        n15133) );
  AOI22_X1 U16640 ( .A1(n10862), .A2(keyinput17), .B1(keyinput22), .B2(n9459), 
        .ZN(n15119) );
  OAI221_X1 U16641 ( .B1(n10862), .B2(keyinput17), .C1(n9459), .C2(keyinput22), 
        .A(n15119), .ZN(n15131) );
  AOI22_X1 U16642 ( .A1(n15122), .A2(keyinput49), .B1(keyinput55), .B2(n15121), 
        .ZN(n15120) );
  OAI221_X1 U16643 ( .B1(n15122), .B2(keyinput49), .C1(n15121), .C2(keyinput55), .A(n15120), .ZN(n15130) );
  AOI22_X1 U16644 ( .A1(n15125), .A2(keyinput44), .B1(n15124), .B2(keyinput0), 
        .ZN(n15123) );
  OAI221_X1 U16645 ( .B1(n15125), .B2(keyinput44), .C1(n15124), .C2(keyinput0), 
        .A(n15123), .ZN(n15129) );
  AOI22_X1 U16646 ( .A1(n11031), .A2(keyinput59), .B1(keyinput5), .B2(n15127), 
        .ZN(n15126) );
  OAI221_X1 U16647 ( .B1(n11031), .B2(keyinput59), .C1(n15127), .C2(keyinput5), 
        .A(n15126), .ZN(n15128) );
  NOR4_X1 U16648 ( .A1(n15131), .A2(n15130), .A3(n15129), .A4(n15128), .ZN(
        n15132) );
  NAND4_X1 U16649 ( .A1(n15135), .A2(n15134), .A3(n15133), .A4(n15132), .ZN(
        n15136) );
  AOI211_X1 U16650 ( .C1(n15139), .C2(n15138), .A(n15137), .B(n15136), .ZN(
        n15140) );
  XNOR2_X1 U16651 ( .A(n15141), .B(n15140), .ZN(P1_U3085) );
  XOR2_X1 U16652 ( .A(n15143), .B(n15142), .Z(SUB_1596_U59) );
  XNOR2_X1 U16653 ( .A(n15144), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16654 ( .B1(n15146), .B2(n15145), .A(n15154), .ZN(SUB_1596_U53) );
  XOR2_X1 U16655 ( .A(n15148), .B(n15147), .Z(SUB_1596_U56) );
  OAI21_X1 U16656 ( .B1(n15151), .B2(n15150), .A(n15149), .ZN(n15152) );
  XNOR2_X1 U16657 ( .A(n15152), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U16658 ( .A(n15154), .B(n15153), .Z(SUB_1596_U5) );
  INV_X1 U7492 ( .A(n13206), .ZN(n13264) );
  CLKBUF_X1 U7209 ( .A(n10107), .Z(n6451) );
  CLKBUF_X1 U7244 ( .A(n7762), .Z(n6770) );
  XNOR2_X1 U7255 ( .A(n9556), .B(n9555), .ZN(n9558) );
  XNOR2_X1 U7603 ( .A(n9568), .B(n9567), .ZN(n11434) );
  AND2_X2 U9296 ( .A1(n6968), .A2(n9558), .ZN(n15191) );
endmodule

